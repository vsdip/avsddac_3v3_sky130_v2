magic
tech sky130A
timestamp 1633152104
<< nwell >>
rect 748 5533 1559 5757
rect 1796 5529 2607 5753
rect 748 4854 1559 5078
rect 3243 4849 4054 5073
rect 748 4086 1559 4310
rect 1796 4082 2607 4306
rect 748 3407 1559 3631
rect 3286 3404 4097 3628
rect 749 2566 1560 2790
rect 1797 2562 2608 2786
rect 749 1887 1560 2111
rect 3244 1882 4055 2106
rect 749 1119 1560 1343
rect 1797 1115 2608 1339
rect 749 440 1560 664
<< nmos >>
rect 812 5432 862 5474
rect 1025 5432 1075 5474
rect 1233 5432 1283 5474
rect 1441 5432 1491 5474
rect 1860 5428 1910 5470
rect 2073 5428 2123 5470
rect 2281 5428 2331 5470
rect 2489 5428 2539 5470
rect 812 4753 862 4795
rect 1025 4753 1075 4795
rect 1233 4753 1283 4795
rect 1441 4753 1491 4795
rect 3307 4748 3357 4790
rect 3520 4748 3570 4790
rect 3728 4748 3778 4790
rect 3936 4748 3986 4790
rect 812 3985 862 4027
rect 1025 3985 1075 4027
rect 1233 3985 1283 4027
rect 1441 3985 1491 4027
rect 1860 3981 1910 4023
rect 2073 3981 2123 4023
rect 2281 3981 2331 4023
rect 2489 3981 2539 4023
rect 812 3306 862 3348
rect 1025 3306 1075 3348
rect 1233 3306 1283 3348
rect 1441 3306 1491 3348
rect 3350 3303 3400 3345
rect 3563 3303 3613 3345
rect 3771 3303 3821 3345
rect 3979 3303 4029 3345
rect 813 2465 863 2507
rect 1026 2465 1076 2507
rect 1234 2465 1284 2507
rect 1442 2465 1492 2507
rect 1861 2461 1911 2503
rect 2074 2461 2124 2503
rect 2282 2461 2332 2503
rect 2490 2461 2540 2503
rect 813 1786 863 1828
rect 1026 1786 1076 1828
rect 1234 1786 1284 1828
rect 1442 1786 1492 1828
rect 3308 1781 3358 1823
rect 3521 1781 3571 1823
rect 3729 1781 3779 1823
rect 3937 1781 3987 1823
rect 813 1018 863 1060
rect 1026 1018 1076 1060
rect 1234 1018 1284 1060
rect 1442 1018 1492 1060
rect 1861 1014 1911 1056
rect 2074 1014 2124 1056
rect 2282 1014 2332 1056
rect 2490 1014 2540 1056
rect 813 339 863 381
rect 1026 339 1076 381
rect 1234 339 1284 381
rect 1442 339 1492 381
<< pmos >>
rect 812 5551 862 5651
rect 1025 5551 1075 5651
rect 1233 5551 1283 5651
rect 1441 5551 1491 5651
rect 1860 5547 1910 5647
rect 2073 5547 2123 5647
rect 2281 5547 2331 5647
rect 2489 5547 2539 5647
rect 812 4872 862 4972
rect 1025 4872 1075 4972
rect 1233 4872 1283 4972
rect 1441 4872 1491 4972
rect 3307 4867 3357 4967
rect 3520 4867 3570 4967
rect 3728 4867 3778 4967
rect 3936 4867 3986 4967
rect 812 4104 862 4204
rect 1025 4104 1075 4204
rect 1233 4104 1283 4204
rect 1441 4104 1491 4204
rect 1860 4100 1910 4200
rect 2073 4100 2123 4200
rect 2281 4100 2331 4200
rect 2489 4100 2539 4200
rect 812 3425 862 3525
rect 1025 3425 1075 3525
rect 1233 3425 1283 3525
rect 1441 3425 1491 3525
rect 3350 3422 3400 3522
rect 3563 3422 3613 3522
rect 3771 3422 3821 3522
rect 3979 3422 4029 3522
rect 813 2584 863 2684
rect 1026 2584 1076 2684
rect 1234 2584 1284 2684
rect 1442 2584 1492 2684
rect 1861 2580 1911 2680
rect 2074 2580 2124 2680
rect 2282 2580 2332 2680
rect 2490 2580 2540 2680
rect 813 1905 863 2005
rect 1026 1905 1076 2005
rect 1234 1905 1284 2005
rect 1442 1905 1492 2005
rect 3308 1900 3358 2000
rect 3521 1900 3571 2000
rect 3729 1900 3779 2000
rect 3937 1900 3987 2000
rect 813 1137 863 1237
rect 1026 1137 1076 1237
rect 1234 1137 1284 1237
rect 1442 1137 1492 1237
rect 1861 1133 1911 1233
rect 2074 1133 2124 1233
rect 2282 1133 2332 1233
rect 2490 1133 2540 1233
rect 813 458 863 558
rect 1026 458 1076 558
rect 1234 458 1284 558
rect 1442 458 1492 558
<< ndiff >>
rect 763 5464 812 5474
rect 763 5444 774 5464
rect 794 5444 812 5464
rect 763 5432 812 5444
rect 862 5468 906 5474
rect 862 5448 877 5468
rect 897 5448 906 5468
rect 862 5432 906 5448
rect 976 5464 1025 5474
rect 976 5444 987 5464
rect 1007 5444 1025 5464
rect 976 5432 1025 5444
rect 1075 5468 1119 5474
rect 1075 5448 1090 5468
rect 1110 5448 1119 5468
rect 1075 5432 1119 5448
rect 1184 5464 1233 5474
rect 1184 5444 1195 5464
rect 1215 5444 1233 5464
rect 1184 5432 1233 5444
rect 1283 5468 1327 5474
rect 1283 5448 1298 5468
rect 1318 5448 1327 5468
rect 1283 5432 1327 5448
rect 1397 5468 1441 5474
rect 1397 5448 1406 5468
rect 1426 5448 1441 5468
rect 1397 5432 1441 5448
rect 1491 5464 1540 5474
rect 1491 5444 1509 5464
rect 1529 5444 1540 5464
rect 1491 5432 1540 5444
rect 1811 5460 1860 5470
rect 1811 5440 1822 5460
rect 1842 5440 1860 5460
rect 1811 5428 1860 5440
rect 1910 5464 1954 5470
rect 1910 5444 1925 5464
rect 1945 5444 1954 5464
rect 1910 5428 1954 5444
rect 2024 5460 2073 5470
rect 2024 5440 2035 5460
rect 2055 5440 2073 5460
rect 2024 5428 2073 5440
rect 2123 5464 2167 5470
rect 2123 5444 2138 5464
rect 2158 5444 2167 5464
rect 2123 5428 2167 5444
rect 2232 5460 2281 5470
rect 2232 5440 2243 5460
rect 2263 5440 2281 5460
rect 2232 5428 2281 5440
rect 2331 5464 2375 5470
rect 2331 5444 2346 5464
rect 2366 5444 2375 5464
rect 2331 5428 2375 5444
rect 2445 5464 2489 5470
rect 2445 5444 2454 5464
rect 2474 5444 2489 5464
rect 2445 5428 2489 5444
rect 2539 5460 2588 5470
rect 2539 5440 2557 5460
rect 2577 5440 2588 5460
rect 2539 5428 2588 5440
rect 763 4785 812 4795
rect 763 4765 774 4785
rect 794 4765 812 4785
rect 763 4753 812 4765
rect 862 4789 906 4795
rect 862 4769 877 4789
rect 897 4769 906 4789
rect 862 4753 906 4769
rect 976 4785 1025 4795
rect 976 4765 987 4785
rect 1007 4765 1025 4785
rect 976 4753 1025 4765
rect 1075 4789 1119 4795
rect 1075 4769 1090 4789
rect 1110 4769 1119 4789
rect 1075 4753 1119 4769
rect 1184 4785 1233 4795
rect 1184 4765 1195 4785
rect 1215 4765 1233 4785
rect 1184 4753 1233 4765
rect 1283 4789 1327 4795
rect 1283 4769 1298 4789
rect 1318 4769 1327 4789
rect 1283 4753 1327 4769
rect 1397 4789 1441 4795
rect 1397 4769 1406 4789
rect 1426 4769 1441 4789
rect 1397 4753 1441 4769
rect 1491 4785 1540 4795
rect 1491 4765 1509 4785
rect 1529 4765 1540 4785
rect 1491 4753 1540 4765
rect 3258 4780 3307 4790
rect 3258 4760 3269 4780
rect 3289 4760 3307 4780
rect 3258 4748 3307 4760
rect 3357 4784 3401 4790
rect 3357 4764 3372 4784
rect 3392 4764 3401 4784
rect 3357 4748 3401 4764
rect 3471 4780 3520 4790
rect 3471 4760 3482 4780
rect 3502 4760 3520 4780
rect 3471 4748 3520 4760
rect 3570 4784 3614 4790
rect 3570 4764 3585 4784
rect 3605 4764 3614 4784
rect 3570 4748 3614 4764
rect 3679 4780 3728 4790
rect 3679 4760 3690 4780
rect 3710 4760 3728 4780
rect 3679 4748 3728 4760
rect 3778 4784 3822 4790
rect 3778 4764 3793 4784
rect 3813 4764 3822 4784
rect 3778 4748 3822 4764
rect 3892 4784 3936 4790
rect 3892 4764 3901 4784
rect 3921 4764 3936 4784
rect 3892 4748 3936 4764
rect 3986 4780 4035 4790
rect 3986 4760 4004 4780
rect 4024 4760 4035 4780
rect 3986 4748 4035 4760
rect 763 4017 812 4027
rect 763 3997 774 4017
rect 794 3997 812 4017
rect 763 3985 812 3997
rect 862 4021 906 4027
rect 862 4001 877 4021
rect 897 4001 906 4021
rect 862 3985 906 4001
rect 976 4017 1025 4027
rect 976 3997 987 4017
rect 1007 3997 1025 4017
rect 976 3985 1025 3997
rect 1075 4021 1119 4027
rect 1075 4001 1090 4021
rect 1110 4001 1119 4021
rect 1075 3985 1119 4001
rect 1184 4017 1233 4027
rect 1184 3997 1195 4017
rect 1215 3997 1233 4017
rect 1184 3985 1233 3997
rect 1283 4021 1327 4027
rect 1283 4001 1298 4021
rect 1318 4001 1327 4021
rect 1283 3985 1327 4001
rect 1397 4021 1441 4027
rect 1397 4001 1406 4021
rect 1426 4001 1441 4021
rect 1397 3985 1441 4001
rect 1491 4017 1540 4027
rect 1491 3997 1509 4017
rect 1529 3997 1540 4017
rect 1491 3985 1540 3997
rect 1811 4013 1860 4023
rect 1811 3993 1822 4013
rect 1842 3993 1860 4013
rect 1811 3981 1860 3993
rect 1910 4017 1954 4023
rect 1910 3997 1925 4017
rect 1945 3997 1954 4017
rect 1910 3981 1954 3997
rect 2024 4013 2073 4023
rect 2024 3993 2035 4013
rect 2055 3993 2073 4013
rect 2024 3981 2073 3993
rect 2123 4017 2167 4023
rect 2123 3997 2138 4017
rect 2158 3997 2167 4017
rect 2123 3981 2167 3997
rect 2232 4013 2281 4023
rect 2232 3993 2243 4013
rect 2263 3993 2281 4013
rect 2232 3981 2281 3993
rect 2331 4017 2375 4023
rect 2331 3997 2346 4017
rect 2366 3997 2375 4017
rect 2331 3981 2375 3997
rect 2445 4017 2489 4023
rect 2445 3997 2454 4017
rect 2474 3997 2489 4017
rect 2445 3981 2489 3997
rect 2539 4013 2588 4023
rect 2539 3993 2557 4013
rect 2577 3993 2588 4013
rect 2539 3981 2588 3993
rect 763 3338 812 3348
rect 763 3318 774 3338
rect 794 3318 812 3338
rect 763 3306 812 3318
rect 862 3342 906 3348
rect 862 3322 877 3342
rect 897 3322 906 3342
rect 862 3306 906 3322
rect 976 3338 1025 3348
rect 976 3318 987 3338
rect 1007 3318 1025 3338
rect 976 3306 1025 3318
rect 1075 3342 1119 3348
rect 1075 3322 1090 3342
rect 1110 3322 1119 3342
rect 1075 3306 1119 3322
rect 1184 3338 1233 3348
rect 1184 3318 1195 3338
rect 1215 3318 1233 3338
rect 1184 3306 1233 3318
rect 1283 3342 1327 3348
rect 1283 3322 1298 3342
rect 1318 3322 1327 3342
rect 1283 3306 1327 3322
rect 1397 3342 1441 3348
rect 1397 3322 1406 3342
rect 1426 3322 1441 3342
rect 1397 3306 1441 3322
rect 1491 3338 1540 3348
rect 1491 3318 1509 3338
rect 1529 3318 1540 3338
rect 1491 3306 1540 3318
rect 3301 3335 3350 3345
rect 3301 3315 3312 3335
rect 3332 3315 3350 3335
rect 3301 3303 3350 3315
rect 3400 3339 3444 3345
rect 3400 3319 3415 3339
rect 3435 3319 3444 3339
rect 3400 3303 3444 3319
rect 3514 3335 3563 3345
rect 3514 3315 3525 3335
rect 3545 3315 3563 3335
rect 3514 3303 3563 3315
rect 3613 3339 3657 3345
rect 3613 3319 3628 3339
rect 3648 3319 3657 3339
rect 3613 3303 3657 3319
rect 3722 3335 3771 3345
rect 3722 3315 3733 3335
rect 3753 3315 3771 3335
rect 3722 3303 3771 3315
rect 3821 3339 3865 3345
rect 3821 3319 3836 3339
rect 3856 3319 3865 3339
rect 3821 3303 3865 3319
rect 3935 3339 3979 3345
rect 3935 3319 3944 3339
rect 3964 3319 3979 3339
rect 3935 3303 3979 3319
rect 4029 3335 4078 3345
rect 4029 3315 4047 3335
rect 4067 3315 4078 3335
rect 4029 3303 4078 3315
rect 764 2497 813 2507
rect 764 2477 775 2497
rect 795 2477 813 2497
rect 764 2465 813 2477
rect 863 2501 907 2507
rect 863 2481 878 2501
rect 898 2481 907 2501
rect 863 2465 907 2481
rect 977 2497 1026 2507
rect 977 2477 988 2497
rect 1008 2477 1026 2497
rect 977 2465 1026 2477
rect 1076 2501 1120 2507
rect 1076 2481 1091 2501
rect 1111 2481 1120 2501
rect 1076 2465 1120 2481
rect 1185 2497 1234 2507
rect 1185 2477 1196 2497
rect 1216 2477 1234 2497
rect 1185 2465 1234 2477
rect 1284 2501 1328 2507
rect 1284 2481 1299 2501
rect 1319 2481 1328 2501
rect 1284 2465 1328 2481
rect 1398 2501 1442 2507
rect 1398 2481 1407 2501
rect 1427 2481 1442 2501
rect 1398 2465 1442 2481
rect 1492 2497 1541 2507
rect 1492 2477 1510 2497
rect 1530 2477 1541 2497
rect 1492 2465 1541 2477
rect 1812 2493 1861 2503
rect 1812 2473 1823 2493
rect 1843 2473 1861 2493
rect 1812 2461 1861 2473
rect 1911 2497 1955 2503
rect 1911 2477 1926 2497
rect 1946 2477 1955 2497
rect 1911 2461 1955 2477
rect 2025 2493 2074 2503
rect 2025 2473 2036 2493
rect 2056 2473 2074 2493
rect 2025 2461 2074 2473
rect 2124 2497 2168 2503
rect 2124 2477 2139 2497
rect 2159 2477 2168 2497
rect 2124 2461 2168 2477
rect 2233 2493 2282 2503
rect 2233 2473 2244 2493
rect 2264 2473 2282 2493
rect 2233 2461 2282 2473
rect 2332 2497 2376 2503
rect 2332 2477 2347 2497
rect 2367 2477 2376 2497
rect 2332 2461 2376 2477
rect 2446 2497 2490 2503
rect 2446 2477 2455 2497
rect 2475 2477 2490 2497
rect 2446 2461 2490 2477
rect 2540 2493 2589 2503
rect 2540 2473 2558 2493
rect 2578 2473 2589 2493
rect 2540 2461 2589 2473
rect 764 1818 813 1828
rect 764 1798 775 1818
rect 795 1798 813 1818
rect 764 1786 813 1798
rect 863 1822 907 1828
rect 863 1802 878 1822
rect 898 1802 907 1822
rect 863 1786 907 1802
rect 977 1818 1026 1828
rect 977 1798 988 1818
rect 1008 1798 1026 1818
rect 977 1786 1026 1798
rect 1076 1822 1120 1828
rect 1076 1802 1091 1822
rect 1111 1802 1120 1822
rect 1076 1786 1120 1802
rect 1185 1818 1234 1828
rect 1185 1798 1196 1818
rect 1216 1798 1234 1818
rect 1185 1786 1234 1798
rect 1284 1822 1328 1828
rect 1284 1802 1299 1822
rect 1319 1802 1328 1822
rect 1284 1786 1328 1802
rect 1398 1822 1442 1828
rect 1398 1802 1407 1822
rect 1427 1802 1442 1822
rect 1398 1786 1442 1802
rect 1492 1818 1541 1828
rect 1492 1798 1510 1818
rect 1530 1798 1541 1818
rect 1492 1786 1541 1798
rect 3259 1813 3308 1823
rect 3259 1793 3270 1813
rect 3290 1793 3308 1813
rect 3259 1781 3308 1793
rect 3358 1817 3402 1823
rect 3358 1797 3373 1817
rect 3393 1797 3402 1817
rect 3358 1781 3402 1797
rect 3472 1813 3521 1823
rect 3472 1793 3483 1813
rect 3503 1793 3521 1813
rect 3472 1781 3521 1793
rect 3571 1817 3615 1823
rect 3571 1797 3586 1817
rect 3606 1797 3615 1817
rect 3571 1781 3615 1797
rect 3680 1813 3729 1823
rect 3680 1793 3691 1813
rect 3711 1793 3729 1813
rect 3680 1781 3729 1793
rect 3779 1817 3823 1823
rect 3779 1797 3794 1817
rect 3814 1797 3823 1817
rect 3779 1781 3823 1797
rect 3893 1817 3937 1823
rect 3893 1797 3902 1817
rect 3922 1797 3937 1817
rect 3893 1781 3937 1797
rect 3987 1813 4036 1823
rect 3987 1793 4005 1813
rect 4025 1793 4036 1813
rect 3987 1781 4036 1793
rect 764 1050 813 1060
rect 764 1030 775 1050
rect 795 1030 813 1050
rect 764 1018 813 1030
rect 863 1054 907 1060
rect 863 1034 878 1054
rect 898 1034 907 1054
rect 863 1018 907 1034
rect 977 1050 1026 1060
rect 977 1030 988 1050
rect 1008 1030 1026 1050
rect 977 1018 1026 1030
rect 1076 1054 1120 1060
rect 1076 1034 1091 1054
rect 1111 1034 1120 1054
rect 1076 1018 1120 1034
rect 1185 1050 1234 1060
rect 1185 1030 1196 1050
rect 1216 1030 1234 1050
rect 1185 1018 1234 1030
rect 1284 1054 1328 1060
rect 1284 1034 1299 1054
rect 1319 1034 1328 1054
rect 1284 1018 1328 1034
rect 1398 1054 1442 1060
rect 1398 1034 1407 1054
rect 1427 1034 1442 1054
rect 1398 1018 1442 1034
rect 1492 1050 1541 1060
rect 1492 1030 1510 1050
rect 1530 1030 1541 1050
rect 1492 1018 1541 1030
rect 1812 1046 1861 1056
rect 1812 1026 1823 1046
rect 1843 1026 1861 1046
rect 1812 1014 1861 1026
rect 1911 1050 1955 1056
rect 1911 1030 1926 1050
rect 1946 1030 1955 1050
rect 1911 1014 1955 1030
rect 2025 1046 2074 1056
rect 2025 1026 2036 1046
rect 2056 1026 2074 1046
rect 2025 1014 2074 1026
rect 2124 1050 2168 1056
rect 2124 1030 2139 1050
rect 2159 1030 2168 1050
rect 2124 1014 2168 1030
rect 2233 1046 2282 1056
rect 2233 1026 2244 1046
rect 2264 1026 2282 1046
rect 2233 1014 2282 1026
rect 2332 1050 2376 1056
rect 2332 1030 2347 1050
rect 2367 1030 2376 1050
rect 2332 1014 2376 1030
rect 2446 1050 2490 1056
rect 2446 1030 2455 1050
rect 2475 1030 2490 1050
rect 2446 1014 2490 1030
rect 2540 1046 2589 1056
rect 2540 1026 2558 1046
rect 2578 1026 2589 1046
rect 2540 1014 2589 1026
rect 764 371 813 381
rect 764 351 775 371
rect 795 351 813 371
rect 764 339 813 351
rect 863 375 907 381
rect 863 355 878 375
rect 898 355 907 375
rect 863 339 907 355
rect 977 371 1026 381
rect 977 351 988 371
rect 1008 351 1026 371
rect 977 339 1026 351
rect 1076 375 1120 381
rect 1076 355 1091 375
rect 1111 355 1120 375
rect 1076 339 1120 355
rect 1185 371 1234 381
rect 1185 351 1196 371
rect 1216 351 1234 371
rect 1185 339 1234 351
rect 1284 375 1328 381
rect 1284 355 1299 375
rect 1319 355 1328 375
rect 1284 339 1328 355
rect 1398 375 1442 381
rect 1398 355 1407 375
rect 1427 355 1442 375
rect 1398 339 1442 355
rect 1492 371 1541 381
rect 1492 351 1510 371
rect 1530 351 1541 371
rect 1492 339 1541 351
<< pdiff >>
rect 768 5613 812 5651
rect 768 5593 780 5613
rect 800 5593 812 5613
rect 768 5551 812 5593
rect 862 5613 904 5651
rect 862 5593 876 5613
rect 896 5593 904 5613
rect 862 5551 904 5593
rect 981 5613 1025 5651
rect 981 5593 993 5613
rect 1013 5593 1025 5613
rect 981 5551 1025 5593
rect 1075 5613 1117 5651
rect 1075 5593 1089 5613
rect 1109 5593 1117 5613
rect 1075 5551 1117 5593
rect 1189 5613 1233 5651
rect 1189 5593 1201 5613
rect 1221 5593 1233 5613
rect 1189 5551 1233 5593
rect 1283 5613 1325 5651
rect 1283 5593 1297 5613
rect 1317 5593 1325 5613
rect 1283 5551 1325 5593
rect 1399 5613 1441 5651
rect 1399 5593 1407 5613
rect 1427 5593 1441 5613
rect 1399 5551 1441 5593
rect 1491 5620 1536 5651
rect 1491 5613 1535 5620
rect 1491 5593 1503 5613
rect 1523 5593 1535 5613
rect 1491 5551 1535 5593
rect 1816 5609 1860 5647
rect 1816 5589 1828 5609
rect 1848 5589 1860 5609
rect 1816 5547 1860 5589
rect 1910 5609 1952 5647
rect 1910 5589 1924 5609
rect 1944 5589 1952 5609
rect 1910 5547 1952 5589
rect 2029 5609 2073 5647
rect 2029 5589 2041 5609
rect 2061 5589 2073 5609
rect 2029 5547 2073 5589
rect 2123 5609 2165 5647
rect 2123 5589 2137 5609
rect 2157 5589 2165 5609
rect 2123 5547 2165 5589
rect 2237 5609 2281 5647
rect 2237 5589 2249 5609
rect 2269 5589 2281 5609
rect 2237 5547 2281 5589
rect 2331 5609 2373 5647
rect 2331 5589 2345 5609
rect 2365 5589 2373 5609
rect 2331 5547 2373 5589
rect 2447 5609 2489 5647
rect 2447 5589 2455 5609
rect 2475 5589 2489 5609
rect 2447 5547 2489 5589
rect 2539 5616 2584 5647
rect 2539 5609 2583 5616
rect 2539 5589 2551 5609
rect 2571 5589 2583 5609
rect 2539 5547 2583 5589
rect 768 4934 812 4972
rect 768 4914 780 4934
rect 800 4914 812 4934
rect 768 4872 812 4914
rect 862 4934 904 4972
rect 862 4914 876 4934
rect 896 4914 904 4934
rect 862 4872 904 4914
rect 981 4934 1025 4972
rect 981 4914 993 4934
rect 1013 4914 1025 4934
rect 981 4872 1025 4914
rect 1075 4934 1117 4972
rect 1075 4914 1089 4934
rect 1109 4914 1117 4934
rect 1075 4872 1117 4914
rect 1189 4934 1233 4972
rect 1189 4914 1201 4934
rect 1221 4914 1233 4934
rect 1189 4872 1233 4914
rect 1283 4934 1325 4972
rect 1283 4914 1297 4934
rect 1317 4914 1325 4934
rect 1283 4872 1325 4914
rect 1399 4934 1441 4972
rect 1399 4914 1407 4934
rect 1427 4914 1441 4934
rect 1399 4872 1441 4914
rect 1491 4941 1536 4972
rect 1491 4934 1535 4941
rect 1491 4914 1503 4934
rect 1523 4914 1535 4934
rect 1491 4872 1535 4914
rect 3263 4929 3307 4967
rect 3263 4909 3275 4929
rect 3295 4909 3307 4929
rect 3263 4867 3307 4909
rect 3357 4929 3399 4967
rect 3357 4909 3371 4929
rect 3391 4909 3399 4929
rect 3357 4867 3399 4909
rect 3476 4929 3520 4967
rect 3476 4909 3488 4929
rect 3508 4909 3520 4929
rect 3476 4867 3520 4909
rect 3570 4929 3612 4967
rect 3570 4909 3584 4929
rect 3604 4909 3612 4929
rect 3570 4867 3612 4909
rect 3684 4929 3728 4967
rect 3684 4909 3696 4929
rect 3716 4909 3728 4929
rect 3684 4867 3728 4909
rect 3778 4929 3820 4967
rect 3778 4909 3792 4929
rect 3812 4909 3820 4929
rect 3778 4867 3820 4909
rect 3894 4929 3936 4967
rect 3894 4909 3902 4929
rect 3922 4909 3936 4929
rect 3894 4867 3936 4909
rect 3986 4936 4031 4967
rect 3986 4929 4030 4936
rect 3986 4909 3998 4929
rect 4018 4909 4030 4929
rect 3986 4867 4030 4909
rect 768 4166 812 4204
rect 768 4146 780 4166
rect 800 4146 812 4166
rect 768 4104 812 4146
rect 862 4166 904 4204
rect 862 4146 876 4166
rect 896 4146 904 4166
rect 862 4104 904 4146
rect 981 4166 1025 4204
rect 981 4146 993 4166
rect 1013 4146 1025 4166
rect 981 4104 1025 4146
rect 1075 4166 1117 4204
rect 1075 4146 1089 4166
rect 1109 4146 1117 4166
rect 1075 4104 1117 4146
rect 1189 4166 1233 4204
rect 1189 4146 1201 4166
rect 1221 4146 1233 4166
rect 1189 4104 1233 4146
rect 1283 4166 1325 4204
rect 1283 4146 1297 4166
rect 1317 4146 1325 4166
rect 1283 4104 1325 4146
rect 1399 4166 1441 4204
rect 1399 4146 1407 4166
rect 1427 4146 1441 4166
rect 1399 4104 1441 4146
rect 1491 4173 1536 4204
rect 1491 4166 1535 4173
rect 1491 4146 1503 4166
rect 1523 4146 1535 4166
rect 1491 4104 1535 4146
rect 1816 4162 1860 4200
rect 1816 4142 1828 4162
rect 1848 4142 1860 4162
rect 1816 4100 1860 4142
rect 1910 4162 1952 4200
rect 1910 4142 1924 4162
rect 1944 4142 1952 4162
rect 1910 4100 1952 4142
rect 2029 4162 2073 4200
rect 2029 4142 2041 4162
rect 2061 4142 2073 4162
rect 2029 4100 2073 4142
rect 2123 4162 2165 4200
rect 2123 4142 2137 4162
rect 2157 4142 2165 4162
rect 2123 4100 2165 4142
rect 2237 4162 2281 4200
rect 2237 4142 2249 4162
rect 2269 4142 2281 4162
rect 2237 4100 2281 4142
rect 2331 4162 2373 4200
rect 2331 4142 2345 4162
rect 2365 4142 2373 4162
rect 2331 4100 2373 4142
rect 2447 4162 2489 4200
rect 2447 4142 2455 4162
rect 2475 4142 2489 4162
rect 2447 4100 2489 4142
rect 2539 4169 2584 4200
rect 2539 4162 2583 4169
rect 2539 4142 2551 4162
rect 2571 4142 2583 4162
rect 2539 4100 2583 4142
rect 768 3487 812 3525
rect 768 3467 780 3487
rect 800 3467 812 3487
rect 768 3425 812 3467
rect 862 3487 904 3525
rect 862 3467 876 3487
rect 896 3467 904 3487
rect 862 3425 904 3467
rect 981 3487 1025 3525
rect 981 3467 993 3487
rect 1013 3467 1025 3487
rect 981 3425 1025 3467
rect 1075 3487 1117 3525
rect 1075 3467 1089 3487
rect 1109 3467 1117 3487
rect 1075 3425 1117 3467
rect 1189 3487 1233 3525
rect 1189 3467 1201 3487
rect 1221 3467 1233 3487
rect 1189 3425 1233 3467
rect 1283 3487 1325 3525
rect 1283 3467 1297 3487
rect 1317 3467 1325 3487
rect 1283 3425 1325 3467
rect 1399 3487 1441 3525
rect 1399 3467 1407 3487
rect 1427 3467 1441 3487
rect 1399 3425 1441 3467
rect 1491 3494 1536 3525
rect 1491 3487 1535 3494
rect 1491 3467 1503 3487
rect 1523 3467 1535 3487
rect 1491 3425 1535 3467
rect 3306 3484 3350 3522
rect 3306 3464 3318 3484
rect 3338 3464 3350 3484
rect 3306 3422 3350 3464
rect 3400 3484 3442 3522
rect 3400 3464 3414 3484
rect 3434 3464 3442 3484
rect 3400 3422 3442 3464
rect 3519 3484 3563 3522
rect 3519 3464 3531 3484
rect 3551 3464 3563 3484
rect 3519 3422 3563 3464
rect 3613 3484 3655 3522
rect 3613 3464 3627 3484
rect 3647 3464 3655 3484
rect 3613 3422 3655 3464
rect 3727 3484 3771 3522
rect 3727 3464 3739 3484
rect 3759 3464 3771 3484
rect 3727 3422 3771 3464
rect 3821 3484 3863 3522
rect 3821 3464 3835 3484
rect 3855 3464 3863 3484
rect 3821 3422 3863 3464
rect 3937 3484 3979 3522
rect 3937 3464 3945 3484
rect 3965 3464 3979 3484
rect 3937 3422 3979 3464
rect 4029 3491 4074 3522
rect 4029 3484 4073 3491
rect 4029 3464 4041 3484
rect 4061 3464 4073 3484
rect 4029 3422 4073 3464
rect 769 2646 813 2684
rect 769 2626 781 2646
rect 801 2626 813 2646
rect 769 2584 813 2626
rect 863 2646 905 2684
rect 863 2626 877 2646
rect 897 2626 905 2646
rect 863 2584 905 2626
rect 982 2646 1026 2684
rect 982 2626 994 2646
rect 1014 2626 1026 2646
rect 982 2584 1026 2626
rect 1076 2646 1118 2684
rect 1076 2626 1090 2646
rect 1110 2626 1118 2646
rect 1076 2584 1118 2626
rect 1190 2646 1234 2684
rect 1190 2626 1202 2646
rect 1222 2626 1234 2646
rect 1190 2584 1234 2626
rect 1284 2646 1326 2684
rect 1284 2626 1298 2646
rect 1318 2626 1326 2646
rect 1284 2584 1326 2626
rect 1400 2646 1442 2684
rect 1400 2626 1408 2646
rect 1428 2626 1442 2646
rect 1400 2584 1442 2626
rect 1492 2653 1537 2684
rect 1492 2646 1536 2653
rect 1492 2626 1504 2646
rect 1524 2626 1536 2646
rect 1492 2584 1536 2626
rect 1817 2642 1861 2680
rect 1817 2622 1829 2642
rect 1849 2622 1861 2642
rect 1817 2580 1861 2622
rect 1911 2642 1953 2680
rect 1911 2622 1925 2642
rect 1945 2622 1953 2642
rect 1911 2580 1953 2622
rect 2030 2642 2074 2680
rect 2030 2622 2042 2642
rect 2062 2622 2074 2642
rect 2030 2580 2074 2622
rect 2124 2642 2166 2680
rect 2124 2622 2138 2642
rect 2158 2622 2166 2642
rect 2124 2580 2166 2622
rect 2238 2642 2282 2680
rect 2238 2622 2250 2642
rect 2270 2622 2282 2642
rect 2238 2580 2282 2622
rect 2332 2642 2374 2680
rect 2332 2622 2346 2642
rect 2366 2622 2374 2642
rect 2332 2580 2374 2622
rect 2448 2642 2490 2680
rect 2448 2622 2456 2642
rect 2476 2622 2490 2642
rect 2448 2580 2490 2622
rect 2540 2649 2585 2680
rect 2540 2642 2584 2649
rect 2540 2622 2552 2642
rect 2572 2622 2584 2642
rect 2540 2580 2584 2622
rect 769 1967 813 2005
rect 769 1947 781 1967
rect 801 1947 813 1967
rect 769 1905 813 1947
rect 863 1967 905 2005
rect 863 1947 877 1967
rect 897 1947 905 1967
rect 863 1905 905 1947
rect 982 1967 1026 2005
rect 982 1947 994 1967
rect 1014 1947 1026 1967
rect 982 1905 1026 1947
rect 1076 1967 1118 2005
rect 1076 1947 1090 1967
rect 1110 1947 1118 1967
rect 1076 1905 1118 1947
rect 1190 1967 1234 2005
rect 1190 1947 1202 1967
rect 1222 1947 1234 1967
rect 1190 1905 1234 1947
rect 1284 1967 1326 2005
rect 1284 1947 1298 1967
rect 1318 1947 1326 1967
rect 1284 1905 1326 1947
rect 1400 1967 1442 2005
rect 1400 1947 1408 1967
rect 1428 1947 1442 1967
rect 1400 1905 1442 1947
rect 1492 1974 1537 2005
rect 1492 1967 1536 1974
rect 1492 1947 1504 1967
rect 1524 1947 1536 1967
rect 1492 1905 1536 1947
rect 3264 1962 3308 2000
rect 3264 1942 3276 1962
rect 3296 1942 3308 1962
rect 3264 1900 3308 1942
rect 3358 1962 3400 2000
rect 3358 1942 3372 1962
rect 3392 1942 3400 1962
rect 3358 1900 3400 1942
rect 3477 1962 3521 2000
rect 3477 1942 3489 1962
rect 3509 1942 3521 1962
rect 3477 1900 3521 1942
rect 3571 1962 3613 2000
rect 3571 1942 3585 1962
rect 3605 1942 3613 1962
rect 3571 1900 3613 1942
rect 3685 1962 3729 2000
rect 3685 1942 3697 1962
rect 3717 1942 3729 1962
rect 3685 1900 3729 1942
rect 3779 1962 3821 2000
rect 3779 1942 3793 1962
rect 3813 1942 3821 1962
rect 3779 1900 3821 1942
rect 3895 1962 3937 2000
rect 3895 1942 3903 1962
rect 3923 1942 3937 1962
rect 3895 1900 3937 1942
rect 3987 1969 4032 2000
rect 3987 1962 4031 1969
rect 3987 1942 3999 1962
rect 4019 1942 4031 1962
rect 3987 1900 4031 1942
rect 769 1199 813 1237
rect 769 1179 781 1199
rect 801 1179 813 1199
rect 769 1137 813 1179
rect 863 1199 905 1237
rect 863 1179 877 1199
rect 897 1179 905 1199
rect 863 1137 905 1179
rect 982 1199 1026 1237
rect 982 1179 994 1199
rect 1014 1179 1026 1199
rect 982 1137 1026 1179
rect 1076 1199 1118 1237
rect 1076 1179 1090 1199
rect 1110 1179 1118 1199
rect 1076 1137 1118 1179
rect 1190 1199 1234 1237
rect 1190 1179 1202 1199
rect 1222 1179 1234 1199
rect 1190 1137 1234 1179
rect 1284 1199 1326 1237
rect 1284 1179 1298 1199
rect 1318 1179 1326 1199
rect 1284 1137 1326 1179
rect 1400 1199 1442 1237
rect 1400 1179 1408 1199
rect 1428 1179 1442 1199
rect 1400 1137 1442 1179
rect 1492 1206 1537 1237
rect 1492 1199 1536 1206
rect 1492 1179 1504 1199
rect 1524 1179 1536 1199
rect 1492 1137 1536 1179
rect 1817 1195 1861 1233
rect 1817 1175 1829 1195
rect 1849 1175 1861 1195
rect 1817 1133 1861 1175
rect 1911 1195 1953 1233
rect 1911 1175 1925 1195
rect 1945 1175 1953 1195
rect 1911 1133 1953 1175
rect 2030 1195 2074 1233
rect 2030 1175 2042 1195
rect 2062 1175 2074 1195
rect 2030 1133 2074 1175
rect 2124 1195 2166 1233
rect 2124 1175 2138 1195
rect 2158 1175 2166 1195
rect 2124 1133 2166 1175
rect 2238 1195 2282 1233
rect 2238 1175 2250 1195
rect 2270 1175 2282 1195
rect 2238 1133 2282 1175
rect 2332 1195 2374 1233
rect 2332 1175 2346 1195
rect 2366 1175 2374 1195
rect 2332 1133 2374 1175
rect 2448 1195 2490 1233
rect 2448 1175 2456 1195
rect 2476 1175 2490 1195
rect 2448 1133 2490 1175
rect 2540 1202 2585 1233
rect 2540 1195 2584 1202
rect 2540 1175 2552 1195
rect 2572 1175 2584 1195
rect 2540 1133 2584 1175
rect 769 520 813 558
rect 769 500 781 520
rect 801 500 813 520
rect 769 458 813 500
rect 863 520 905 558
rect 863 500 877 520
rect 897 500 905 520
rect 863 458 905 500
rect 982 520 1026 558
rect 982 500 994 520
rect 1014 500 1026 520
rect 982 458 1026 500
rect 1076 520 1118 558
rect 1076 500 1090 520
rect 1110 500 1118 520
rect 1076 458 1118 500
rect 1190 520 1234 558
rect 1190 500 1202 520
rect 1222 500 1234 520
rect 1190 458 1234 500
rect 1284 520 1326 558
rect 1284 500 1298 520
rect 1318 500 1326 520
rect 1284 458 1326 500
rect 1400 520 1442 558
rect 1400 500 1408 520
rect 1428 500 1442 520
rect 1400 458 1442 500
rect 1492 527 1537 558
rect 1492 520 1536 527
rect 1492 500 1504 520
rect 1524 500 1536 520
rect 1492 458 1536 500
<< ndiffc >>
rect 454 5767 472 5785
rect 456 5668 474 5686
rect 454 5511 472 5529
rect 774 5444 794 5464
rect 877 5448 897 5468
rect 987 5444 1007 5464
rect 1090 5448 1110 5468
rect 1195 5444 1215 5464
rect 1298 5448 1318 5468
rect 1406 5448 1426 5468
rect 1509 5444 1529 5464
rect 1822 5440 1842 5460
rect 456 5412 474 5430
rect 1925 5444 1945 5464
rect 2035 5440 2055 5460
rect 2138 5444 2158 5464
rect 2243 5440 2263 5460
rect 2346 5444 2366 5464
rect 2454 5444 2474 5464
rect 2557 5440 2577 5460
rect 454 5116 472 5134
rect 456 5017 474 5035
rect 454 4861 472 4879
rect 456 4762 474 4780
rect 774 4765 794 4785
rect 877 4769 897 4789
rect 987 4765 1007 4785
rect 1090 4769 1110 4789
rect 1195 4765 1215 4785
rect 1298 4769 1318 4789
rect 1406 4769 1426 4789
rect 1509 4765 1529 4785
rect 3269 4760 3289 4780
rect 3372 4764 3392 4784
rect 3482 4760 3502 4780
rect 3585 4764 3605 4784
rect 3690 4760 3710 4780
rect 3793 4764 3813 4784
rect 3901 4764 3921 4784
rect 4004 4760 4024 4780
rect 454 4320 472 4338
rect 456 4221 474 4239
rect 454 4064 472 4082
rect 774 3997 794 4017
rect 877 4001 897 4021
rect 987 3997 1007 4017
rect 1090 4001 1110 4021
rect 1195 3997 1215 4017
rect 1298 4001 1318 4021
rect 1406 4001 1426 4021
rect 1509 3997 1529 4017
rect 1822 3993 1842 4013
rect 456 3965 474 3983
rect 1925 3997 1945 4017
rect 2035 3993 2055 4013
rect 2138 3997 2158 4017
rect 2243 3993 2263 4013
rect 2346 3997 2366 4017
rect 2454 3997 2474 4017
rect 2557 3993 2577 4013
rect 454 3669 472 3687
rect 456 3570 474 3588
rect 454 3414 472 3432
rect 456 3315 474 3333
rect 774 3318 794 3338
rect 877 3322 897 3342
rect 987 3318 1007 3338
rect 1090 3322 1110 3342
rect 1195 3318 1215 3338
rect 1298 3322 1318 3342
rect 1406 3322 1426 3342
rect 1509 3318 1529 3338
rect 3312 3315 3332 3335
rect 3415 3319 3435 3339
rect 3525 3315 3545 3335
rect 3628 3319 3648 3339
rect 3733 3315 3753 3335
rect 3836 3319 3856 3339
rect 3944 3319 3964 3339
rect 4047 3315 4067 3335
rect 455 2800 473 2818
rect 457 2701 475 2719
rect 455 2544 473 2562
rect 775 2477 795 2497
rect 878 2481 898 2501
rect 988 2477 1008 2497
rect 1091 2481 1111 2501
rect 1196 2477 1216 2497
rect 1299 2481 1319 2501
rect 1407 2481 1427 2501
rect 1510 2477 1530 2497
rect 1823 2473 1843 2493
rect 457 2445 475 2463
rect 1926 2477 1946 2497
rect 2036 2473 2056 2493
rect 2139 2477 2159 2497
rect 2244 2473 2264 2493
rect 2347 2477 2367 2497
rect 2455 2477 2475 2497
rect 2558 2473 2578 2493
rect 455 2149 473 2167
rect 457 2050 475 2068
rect 455 1894 473 1912
rect 457 1795 475 1813
rect 775 1798 795 1818
rect 878 1802 898 1822
rect 988 1798 1008 1818
rect 1091 1802 1111 1822
rect 1196 1798 1216 1818
rect 1299 1802 1319 1822
rect 1407 1802 1427 1822
rect 1510 1798 1530 1818
rect 3270 1793 3290 1813
rect 3373 1797 3393 1817
rect 3483 1793 3503 1813
rect 3586 1797 3606 1817
rect 3691 1793 3711 1813
rect 3794 1797 3814 1817
rect 3902 1797 3922 1817
rect 4005 1793 4025 1813
rect 455 1353 473 1371
rect 457 1254 475 1272
rect 455 1097 473 1115
rect 775 1030 795 1050
rect 878 1034 898 1054
rect 988 1030 1008 1050
rect 1091 1034 1111 1054
rect 1196 1030 1216 1050
rect 1299 1034 1319 1054
rect 1407 1034 1427 1054
rect 1510 1030 1530 1050
rect 1823 1026 1843 1046
rect 457 998 475 1016
rect 1926 1030 1946 1050
rect 2036 1026 2056 1046
rect 2139 1030 2159 1050
rect 2244 1026 2264 1046
rect 2347 1030 2367 1050
rect 2455 1030 2475 1050
rect 2558 1026 2578 1046
rect 455 702 473 720
rect 457 603 475 621
rect 455 447 473 465
rect 457 348 475 366
rect 775 351 795 371
rect 878 355 898 375
rect 988 351 1008 371
rect 1091 355 1111 375
rect 1196 351 1216 371
rect 1299 355 1319 375
rect 1407 355 1427 375
rect 1510 351 1530 371
<< pdiffc >>
rect 780 5593 800 5613
rect 876 5593 896 5613
rect 993 5593 1013 5613
rect 1089 5593 1109 5613
rect 1201 5593 1221 5613
rect 1297 5593 1317 5613
rect 1407 5593 1427 5613
rect 1503 5593 1523 5613
rect 1828 5589 1848 5609
rect 1924 5589 1944 5609
rect 2041 5589 2061 5609
rect 2137 5589 2157 5609
rect 2249 5589 2269 5609
rect 2345 5589 2365 5609
rect 2455 5589 2475 5609
rect 2551 5589 2571 5609
rect 780 4914 800 4934
rect 876 4914 896 4934
rect 993 4914 1013 4934
rect 1089 4914 1109 4934
rect 1201 4914 1221 4934
rect 1297 4914 1317 4934
rect 1407 4914 1427 4934
rect 1503 4914 1523 4934
rect 3275 4909 3295 4929
rect 3371 4909 3391 4929
rect 3488 4909 3508 4929
rect 3584 4909 3604 4929
rect 3696 4909 3716 4929
rect 3792 4909 3812 4929
rect 3902 4909 3922 4929
rect 3998 4909 4018 4929
rect 780 4146 800 4166
rect 876 4146 896 4166
rect 993 4146 1013 4166
rect 1089 4146 1109 4166
rect 1201 4146 1221 4166
rect 1297 4146 1317 4166
rect 1407 4146 1427 4166
rect 1503 4146 1523 4166
rect 1828 4142 1848 4162
rect 1924 4142 1944 4162
rect 2041 4142 2061 4162
rect 2137 4142 2157 4162
rect 2249 4142 2269 4162
rect 2345 4142 2365 4162
rect 2455 4142 2475 4162
rect 2551 4142 2571 4162
rect 780 3467 800 3487
rect 876 3467 896 3487
rect 993 3467 1013 3487
rect 1089 3467 1109 3487
rect 1201 3467 1221 3487
rect 1297 3467 1317 3487
rect 1407 3467 1427 3487
rect 1503 3467 1523 3487
rect 3318 3464 3338 3484
rect 3414 3464 3434 3484
rect 3531 3464 3551 3484
rect 3627 3464 3647 3484
rect 3739 3464 3759 3484
rect 3835 3464 3855 3484
rect 3945 3464 3965 3484
rect 4041 3464 4061 3484
rect 781 2626 801 2646
rect 877 2626 897 2646
rect 994 2626 1014 2646
rect 1090 2626 1110 2646
rect 1202 2626 1222 2646
rect 1298 2626 1318 2646
rect 1408 2626 1428 2646
rect 1504 2626 1524 2646
rect 1829 2622 1849 2642
rect 1925 2622 1945 2642
rect 2042 2622 2062 2642
rect 2138 2622 2158 2642
rect 2250 2622 2270 2642
rect 2346 2622 2366 2642
rect 2456 2622 2476 2642
rect 2552 2622 2572 2642
rect 781 1947 801 1967
rect 877 1947 897 1967
rect 994 1947 1014 1967
rect 1090 1947 1110 1967
rect 1202 1947 1222 1967
rect 1298 1947 1318 1967
rect 1408 1947 1428 1967
rect 1504 1947 1524 1967
rect 3276 1942 3296 1962
rect 3372 1942 3392 1962
rect 3489 1942 3509 1962
rect 3585 1942 3605 1962
rect 3697 1942 3717 1962
rect 3793 1942 3813 1962
rect 3903 1942 3923 1962
rect 3999 1942 4019 1962
rect 781 1179 801 1199
rect 877 1179 897 1199
rect 994 1179 1014 1199
rect 1090 1179 1110 1199
rect 1202 1179 1222 1199
rect 1298 1179 1318 1199
rect 1408 1179 1428 1199
rect 1504 1179 1524 1199
rect 1829 1175 1849 1195
rect 1925 1175 1945 1195
rect 2042 1175 2062 1195
rect 2138 1175 2158 1195
rect 2250 1175 2270 1195
rect 2346 1175 2366 1195
rect 2456 1175 2476 1195
rect 2552 1175 2572 1195
rect 781 500 801 520
rect 877 500 897 520
rect 994 500 1014 520
rect 1090 500 1110 520
rect 1202 500 1222 520
rect 1298 500 1318 520
rect 1408 500 1428 520
rect 1504 500 1524 520
<< psubdiff >>
rect 848 5377 959 5391
rect 848 5347 889 5377
rect 917 5347 959 5377
rect 848 5332 959 5347
rect 1896 5373 2007 5387
rect 1896 5343 1937 5373
rect 1965 5343 2007 5373
rect 1896 5328 2007 5343
rect 848 4698 959 4712
rect 848 4668 889 4698
rect 917 4668 959 4698
rect 848 4655 959 4668
rect 3343 4693 3454 4707
rect 3343 4663 3384 4693
rect 3412 4663 3454 4693
rect 3343 4648 3454 4663
rect 848 3930 959 3944
rect 848 3900 889 3930
rect 917 3900 959 3930
rect 848 3885 959 3900
rect 1896 3926 2007 3940
rect 1896 3896 1937 3926
rect 1965 3896 2007 3926
rect 1896 3881 2007 3896
rect 848 3251 959 3265
rect 848 3221 889 3251
rect 917 3221 959 3251
rect 848 3206 959 3221
rect 3386 3248 3497 3262
rect 3386 3218 3427 3248
rect 3455 3218 3497 3248
rect 3386 3203 3497 3218
rect 849 2410 960 2424
rect 849 2380 890 2410
rect 918 2380 960 2410
rect 849 2365 960 2380
rect 1897 2406 2008 2420
rect 1897 2376 1938 2406
rect 1966 2376 2008 2406
rect 1897 2361 2008 2376
rect 849 1731 960 1745
rect 849 1701 890 1731
rect 918 1701 960 1731
rect 849 1688 960 1701
rect 3344 1726 3455 1740
rect 3344 1696 3385 1726
rect 3413 1696 3455 1726
rect 3344 1681 3455 1696
rect 849 963 960 977
rect 849 933 890 963
rect 918 933 960 963
rect 849 918 960 933
rect 1897 959 2008 973
rect 1897 929 1938 959
rect 1966 929 2008 959
rect 1897 914 2008 929
rect 849 284 960 298
rect 849 254 890 284
rect 918 254 960 284
rect 849 239 960 254
<< nsubdiff >>
rect 849 5724 959 5738
rect 849 5694 892 5724
rect 920 5694 959 5724
rect 849 5679 959 5694
rect 1897 5720 2007 5734
rect 1897 5690 1940 5720
rect 1968 5690 2007 5720
rect 1897 5675 2007 5690
rect 849 5045 959 5059
rect 849 5015 892 5045
rect 920 5015 959 5045
rect 849 5000 959 5015
rect 3344 5040 3454 5054
rect 3344 5010 3387 5040
rect 3415 5010 3454 5040
rect 3344 4995 3454 5010
rect 849 4277 959 4291
rect 849 4247 892 4277
rect 920 4247 959 4277
rect 849 4232 959 4247
rect 1897 4273 2007 4287
rect 1897 4243 1940 4273
rect 1968 4243 2007 4273
rect 1897 4228 2007 4243
rect 849 3598 959 3612
rect 849 3568 892 3598
rect 920 3568 959 3598
rect 849 3553 959 3568
rect 3387 3595 3497 3609
rect 3387 3565 3430 3595
rect 3458 3565 3497 3595
rect 3387 3550 3497 3565
rect 850 2757 960 2771
rect 850 2727 893 2757
rect 921 2727 960 2757
rect 850 2712 960 2727
rect 1898 2753 2008 2767
rect 1898 2723 1941 2753
rect 1969 2723 2008 2753
rect 1898 2708 2008 2723
rect 850 2078 960 2092
rect 850 2048 893 2078
rect 921 2048 960 2078
rect 850 2033 960 2048
rect 3345 2073 3455 2087
rect 3345 2043 3388 2073
rect 3416 2043 3455 2073
rect 3345 2028 3455 2043
rect 850 1310 960 1324
rect 850 1280 893 1310
rect 921 1280 960 1310
rect 850 1265 960 1280
rect 1898 1306 2008 1320
rect 1898 1276 1941 1306
rect 1969 1276 2008 1306
rect 1898 1261 2008 1276
rect 850 631 960 645
rect 850 601 893 631
rect 921 601 960 631
rect 850 586 960 601
<< psubdiffcont >>
rect 889 5347 917 5377
rect 1937 5343 1965 5373
rect 889 4668 917 4698
rect 3384 4663 3412 4693
rect 889 3900 917 3930
rect 1937 3896 1965 3926
rect 889 3221 917 3251
rect 3427 3218 3455 3248
rect 890 2380 918 2410
rect 1938 2376 1966 2406
rect 890 1701 918 1731
rect 3385 1696 3413 1726
rect 890 933 918 963
rect 1938 929 1966 959
rect 890 254 918 284
<< nsubdiffcont >>
rect 892 5694 920 5724
rect 1940 5690 1968 5720
rect 892 5015 920 5045
rect 3387 5010 3415 5040
rect 892 4247 920 4277
rect 1940 4243 1968 4273
rect 892 3568 920 3598
rect 3430 3565 3458 3595
rect 893 2727 921 2757
rect 1941 2723 1969 2753
rect 893 2048 921 2078
rect 3388 2043 3416 2073
rect 893 1280 921 1310
rect 1941 1276 1969 1306
rect 893 601 921 631
<< poly >>
rect 812 5651 862 5664
rect 1025 5651 1075 5664
rect 1233 5651 1283 5664
rect 1441 5651 1491 5664
rect 1860 5647 1910 5660
rect 2073 5647 2123 5660
rect 2281 5647 2331 5660
rect 2489 5647 2539 5660
rect 812 5523 862 5551
rect 812 5503 825 5523
rect 845 5503 862 5523
rect 812 5474 862 5503
rect 1025 5522 1075 5551
rect 1025 5498 1036 5522
rect 1060 5498 1075 5522
rect 1025 5474 1075 5498
rect 1233 5527 1283 5551
rect 1233 5503 1245 5527
rect 1269 5503 1283 5527
rect 1233 5474 1283 5503
rect 1441 5525 1491 5551
rect 1441 5499 1459 5525
rect 1485 5499 1491 5525
rect 1441 5474 1491 5499
rect 1860 5519 1910 5547
rect 1860 5499 1873 5519
rect 1893 5499 1910 5519
rect 1860 5470 1910 5499
rect 2073 5518 2123 5547
rect 2073 5494 2084 5518
rect 2108 5494 2123 5518
rect 2073 5470 2123 5494
rect 2281 5523 2331 5547
rect 2281 5499 2293 5523
rect 2317 5499 2331 5523
rect 2281 5470 2331 5499
rect 2489 5521 2539 5547
rect 2489 5495 2507 5521
rect 2533 5495 2539 5521
rect 2489 5470 2539 5495
rect 812 5416 862 5432
rect 1025 5416 1075 5432
rect 1233 5416 1283 5432
rect 1441 5416 1491 5432
rect 1860 5412 1910 5428
rect 2073 5412 2123 5428
rect 2281 5412 2331 5428
rect 2489 5412 2539 5428
rect 812 4972 862 4985
rect 1025 4972 1075 4985
rect 1233 4972 1283 4985
rect 1441 4972 1491 4985
rect 3307 4967 3357 4980
rect 3520 4967 3570 4980
rect 3728 4967 3778 4980
rect 3936 4967 3986 4980
rect 812 4844 862 4872
rect 812 4824 825 4844
rect 845 4824 862 4844
rect 812 4795 862 4824
rect 1025 4843 1075 4872
rect 1025 4819 1036 4843
rect 1060 4819 1075 4843
rect 1025 4795 1075 4819
rect 1233 4848 1283 4872
rect 1233 4824 1245 4848
rect 1269 4824 1283 4848
rect 1233 4795 1283 4824
rect 1441 4846 1491 4872
rect 1441 4820 1459 4846
rect 1485 4820 1491 4846
rect 1441 4795 1491 4820
rect 3307 4839 3357 4867
rect 3307 4819 3320 4839
rect 3340 4819 3357 4839
rect 3307 4790 3357 4819
rect 3520 4838 3570 4867
rect 3520 4814 3531 4838
rect 3555 4814 3570 4838
rect 3520 4790 3570 4814
rect 3728 4843 3778 4867
rect 3728 4819 3740 4843
rect 3764 4819 3778 4843
rect 3728 4790 3778 4819
rect 3936 4841 3986 4867
rect 3936 4815 3954 4841
rect 3980 4815 3986 4841
rect 3936 4790 3986 4815
rect 812 4737 862 4753
rect 1025 4737 1075 4753
rect 1233 4737 1283 4753
rect 1441 4737 1491 4753
rect 3307 4732 3357 4748
rect 3520 4732 3570 4748
rect 3728 4732 3778 4748
rect 3936 4732 3986 4748
rect 812 4204 862 4217
rect 1025 4204 1075 4217
rect 1233 4204 1283 4217
rect 1441 4204 1491 4217
rect 1860 4200 1910 4213
rect 2073 4200 2123 4213
rect 2281 4200 2331 4213
rect 2489 4200 2539 4213
rect 812 4076 862 4104
rect 812 4056 825 4076
rect 845 4056 862 4076
rect 812 4027 862 4056
rect 1025 4075 1075 4104
rect 1025 4051 1036 4075
rect 1060 4051 1075 4075
rect 1025 4027 1075 4051
rect 1233 4080 1283 4104
rect 1233 4056 1245 4080
rect 1269 4056 1283 4080
rect 1233 4027 1283 4056
rect 1441 4078 1491 4104
rect 1441 4052 1459 4078
rect 1485 4052 1491 4078
rect 1441 4027 1491 4052
rect 1860 4072 1910 4100
rect 1860 4052 1873 4072
rect 1893 4052 1910 4072
rect 1860 4023 1910 4052
rect 2073 4071 2123 4100
rect 2073 4047 2084 4071
rect 2108 4047 2123 4071
rect 2073 4023 2123 4047
rect 2281 4076 2331 4100
rect 2281 4052 2293 4076
rect 2317 4052 2331 4076
rect 2281 4023 2331 4052
rect 2489 4074 2539 4100
rect 2489 4048 2507 4074
rect 2533 4048 2539 4074
rect 2489 4023 2539 4048
rect 812 3969 862 3985
rect 1025 3969 1075 3985
rect 1233 3969 1283 3985
rect 1441 3969 1491 3985
rect 1860 3965 1910 3981
rect 2073 3965 2123 3981
rect 2281 3965 2331 3981
rect 2489 3965 2539 3981
rect 812 3525 862 3538
rect 1025 3525 1075 3538
rect 1233 3525 1283 3538
rect 1441 3525 1491 3538
rect 3350 3522 3400 3535
rect 3563 3522 3613 3535
rect 3771 3522 3821 3535
rect 3979 3522 4029 3535
rect 812 3397 862 3425
rect 812 3377 825 3397
rect 845 3377 862 3397
rect 812 3348 862 3377
rect 1025 3396 1075 3425
rect 1025 3372 1036 3396
rect 1060 3372 1075 3396
rect 1025 3348 1075 3372
rect 1233 3401 1283 3425
rect 1233 3377 1245 3401
rect 1269 3377 1283 3401
rect 1233 3348 1283 3377
rect 1441 3399 1491 3425
rect 1441 3373 1459 3399
rect 1485 3373 1491 3399
rect 1441 3348 1491 3373
rect 3350 3394 3400 3422
rect 3350 3374 3363 3394
rect 3383 3374 3400 3394
rect 3350 3345 3400 3374
rect 3563 3393 3613 3422
rect 3563 3369 3574 3393
rect 3598 3369 3613 3393
rect 3563 3345 3613 3369
rect 3771 3398 3821 3422
rect 3771 3374 3783 3398
rect 3807 3374 3821 3398
rect 3771 3345 3821 3374
rect 3979 3396 4029 3422
rect 3979 3370 3997 3396
rect 4023 3370 4029 3396
rect 3979 3345 4029 3370
rect 812 3290 862 3306
rect 1025 3290 1075 3306
rect 1233 3290 1283 3306
rect 1441 3290 1491 3306
rect 3350 3287 3400 3303
rect 3563 3287 3613 3303
rect 3771 3287 3821 3303
rect 3979 3287 4029 3303
rect 813 2684 863 2697
rect 1026 2684 1076 2697
rect 1234 2684 1284 2697
rect 1442 2684 1492 2697
rect 1861 2680 1911 2693
rect 2074 2680 2124 2693
rect 2282 2680 2332 2693
rect 2490 2680 2540 2693
rect 813 2556 863 2584
rect 813 2536 826 2556
rect 846 2536 863 2556
rect 813 2507 863 2536
rect 1026 2555 1076 2584
rect 1026 2531 1037 2555
rect 1061 2531 1076 2555
rect 1026 2507 1076 2531
rect 1234 2560 1284 2584
rect 1234 2536 1246 2560
rect 1270 2536 1284 2560
rect 1234 2507 1284 2536
rect 1442 2558 1492 2584
rect 1442 2532 1460 2558
rect 1486 2532 1492 2558
rect 1442 2507 1492 2532
rect 1861 2552 1911 2580
rect 1861 2532 1874 2552
rect 1894 2532 1911 2552
rect 1861 2503 1911 2532
rect 2074 2551 2124 2580
rect 2074 2527 2085 2551
rect 2109 2527 2124 2551
rect 2074 2503 2124 2527
rect 2282 2556 2332 2580
rect 2282 2532 2294 2556
rect 2318 2532 2332 2556
rect 2282 2503 2332 2532
rect 2490 2554 2540 2580
rect 2490 2528 2508 2554
rect 2534 2528 2540 2554
rect 2490 2503 2540 2528
rect 813 2449 863 2465
rect 1026 2449 1076 2465
rect 1234 2449 1284 2465
rect 1442 2449 1492 2465
rect 1861 2445 1911 2461
rect 2074 2445 2124 2461
rect 2282 2445 2332 2461
rect 2490 2445 2540 2461
rect 813 2005 863 2018
rect 1026 2005 1076 2018
rect 1234 2005 1284 2018
rect 1442 2005 1492 2018
rect 3308 2000 3358 2013
rect 3521 2000 3571 2013
rect 3729 2000 3779 2013
rect 3937 2000 3987 2013
rect 813 1877 863 1905
rect 813 1857 826 1877
rect 846 1857 863 1877
rect 813 1828 863 1857
rect 1026 1876 1076 1905
rect 1026 1852 1037 1876
rect 1061 1852 1076 1876
rect 1026 1828 1076 1852
rect 1234 1881 1284 1905
rect 1234 1857 1246 1881
rect 1270 1857 1284 1881
rect 1234 1828 1284 1857
rect 1442 1879 1492 1905
rect 1442 1853 1460 1879
rect 1486 1853 1492 1879
rect 1442 1828 1492 1853
rect 3308 1872 3358 1900
rect 3308 1852 3321 1872
rect 3341 1852 3358 1872
rect 3308 1823 3358 1852
rect 3521 1871 3571 1900
rect 3521 1847 3532 1871
rect 3556 1847 3571 1871
rect 3521 1823 3571 1847
rect 3729 1876 3779 1900
rect 3729 1852 3741 1876
rect 3765 1852 3779 1876
rect 3729 1823 3779 1852
rect 3937 1874 3987 1900
rect 3937 1848 3955 1874
rect 3981 1848 3987 1874
rect 3937 1823 3987 1848
rect 813 1770 863 1786
rect 1026 1770 1076 1786
rect 1234 1770 1284 1786
rect 1442 1770 1492 1786
rect 3308 1765 3358 1781
rect 3521 1765 3571 1781
rect 3729 1765 3779 1781
rect 3937 1765 3987 1781
rect 813 1237 863 1250
rect 1026 1237 1076 1250
rect 1234 1237 1284 1250
rect 1442 1237 1492 1250
rect 1861 1233 1911 1246
rect 2074 1233 2124 1246
rect 2282 1233 2332 1246
rect 2490 1233 2540 1246
rect 813 1109 863 1137
rect 813 1089 826 1109
rect 846 1089 863 1109
rect 813 1060 863 1089
rect 1026 1108 1076 1137
rect 1026 1084 1037 1108
rect 1061 1084 1076 1108
rect 1026 1060 1076 1084
rect 1234 1113 1284 1137
rect 1234 1089 1246 1113
rect 1270 1089 1284 1113
rect 1234 1060 1284 1089
rect 1442 1111 1492 1137
rect 1442 1085 1460 1111
rect 1486 1085 1492 1111
rect 1442 1060 1492 1085
rect 1861 1105 1911 1133
rect 1861 1085 1874 1105
rect 1894 1085 1911 1105
rect 1861 1056 1911 1085
rect 2074 1104 2124 1133
rect 2074 1080 2085 1104
rect 2109 1080 2124 1104
rect 2074 1056 2124 1080
rect 2282 1109 2332 1133
rect 2282 1085 2294 1109
rect 2318 1085 2332 1109
rect 2282 1056 2332 1085
rect 2490 1107 2540 1133
rect 2490 1081 2508 1107
rect 2534 1081 2540 1107
rect 2490 1056 2540 1081
rect 813 1002 863 1018
rect 1026 1002 1076 1018
rect 1234 1002 1284 1018
rect 1442 1002 1492 1018
rect 1861 998 1911 1014
rect 2074 998 2124 1014
rect 2282 998 2332 1014
rect 2490 998 2540 1014
rect 813 558 863 571
rect 1026 558 1076 571
rect 1234 558 1284 571
rect 1442 558 1492 571
rect 813 430 863 458
rect 813 410 826 430
rect 846 410 863 430
rect 813 381 863 410
rect 1026 429 1076 458
rect 1026 405 1037 429
rect 1061 405 1076 429
rect 1026 381 1076 405
rect 1234 434 1284 458
rect 1234 410 1246 434
rect 1270 410 1284 434
rect 1234 381 1284 410
rect 1442 432 1492 458
rect 1442 406 1460 432
rect 1486 406 1492 432
rect 1442 381 1492 406
rect 813 323 863 339
rect 1026 323 1076 339
rect 1234 323 1284 339
rect 1442 323 1492 339
<< polycont >>
rect 825 5503 845 5523
rect 1036 5498 1060 5522
rect 1245 5503 1269 5527
rect 1459 5499 1485 5525
rect 1873 5499 1893 5519
rect 2084 5494 2108 5518
rect 2293 5499 2317 5523
rect 2507 5495 2533 5521
rect 825 4824 845 4844
rect 1036 4819 1060 4843
rect 1245 4824 1269 4848
rect 1459 4820 1485 4846
rect 3320 4819 3340 4839
rect 3531 4814 3555 4838
rect 3740 4819 3764 4843
rect 3954 4815 3980 4841
rect 825 4056 845 4076
rect 1036 4051 1060 4075
rect 1245 4056 1269 4080
rect 1459 4052 1485 4078
rect 1873 4052 1893 4072
rect 2084 4047 2108 4071
rect 2293 4052 2317 4076
rect 2507 4048 2533 4074
rect 825 3377 845 3397
rect 1036 3372 1060 3396
rect 1245 3377 1269 3401
rect 1459 3373 1485 3399
rect 3363 3374 3383 3394
rect 3574 3369 3598 3393
rect 3783 3374 3807 3398
rect 3997 3370 4023 3396
rect 826 2536 846 2556
rect 1037 2531 1061 2555
rect 1246 2536 1270 2560
rect 1460 2532 1486 2558
rect 1874 2532 1894 2552
rect 2085 2527 2109 2551
rect 2294 2532 2318 2556
rect 2508 2528 2534 2554
rect 826 1857 846 1877
rect 1037 1852 1061 1876
rect 1246 1857 1270 1881
rect 1460 1853 1486 1879
rect 3321 1852 3341 1872
rect 3532 1847 3556 1871
rect 3741 1852 3765 1876
rect 3955 1848 3981 1874
rect 826 1089 846 1109
rect 1037 1084 1061 1108
rect 1246 1089 1270 1113
rect 1460 1085 1486 1111
rect 1874 1085 1894 1105
rect 2085 1080 2109 1104
rect 2294 1085 2318 1109
rect 2508 1081 2534 1107
rect 826 410 846 430
rect 1037 405 1061 429
rect 1246 410 1270 434
rect 1460 406 1486 432
<< ndiffres >>
rect 433 5785 490 5804
rect 433 5782 454 5785
rect 339 5767 454 5782
rect 472 5767 490 5785
rect 339 5744 490 5767
rect 339 5708 381 5744
rect 338 5707 438 5708
rect 338 5686 494 5707
rect 338 5668 456 5686
rect 474 5668 494 5686
rect 338 5664 494 5668
rect 433 5648 494 5664
rect 433 5529 490 5548
rect 433 5526 454 5529
rect 339 5511 454 5526
rect 472 5511 490 5529
rect 339 5488 490 5511
rect 339 5452 381 5488
rect 338 5451 438 5452
rect 338 5430 494 5451
rect 338 5412 456 5430
rect 474 5412 494 5430
rect 338 5408 494 5412
rect 433 5392 494 5408
rect 433 5134 490 5153
rect 433 5131 454 5134
rect 339 5116 454 5131
rect 472 5116 490 5134
rect 339 5093 490 5116
rect 339 5057 381 5093
rect 338 5056 438 5057
rect 338 5035 494 5056
rect 338 5017 456 5035
rect 474 5017 494 5035
rect 338 5013 494 5017
rect 433 4997 494 5013
rect 433 4879 490 4898
rect 433 4876 454 4879
rect 339 4861 454 4876
rect 472 4861 490 4879
rect 339 4838 490 4861
rect 339 4802 381 4838
rect 338 4801 438 4802
rect 338 4780 494 4801
rect 338 4762 456 4780
rect 474 4762 494 4780
rect 338 4758 494 4762
rect 433 4742 494 4758
rect 433 4338 490 4357
rect 433 4335 454 4338
rect 339 4320 454 4335
rect 472 4320 490 4338
rect 339 4297 490 4320
rect 339 4261 381 4297
rect 338 4260 438 4261
rect 338 4239 494 4260
rect 338 4221 456 4239
rect 474 4221 494 4239
rect 338 4217 494 4221
rect 433 4201 494 4217
rect 433 4082 490 4101
rect 433 4079 454 4082
rect 339 4064 454 4079
rect 472 4064 490 4082
rect 339 4041 490 4064
rect 339 4005 381 4041
rect 338 4004 438 4005
rect 338 3983 494 4004
rect 338 3965 456 3983
rect 474 3965 494 3983
rect 338 3961 494 3965
rect 433 3945 494 3961
rect 433 3687 490 3706
rect 433 3684 454 3687
rect 339 3669 454 3684
rect 472 3669 490 3687
rect 339 3646 490 3669
rect 339 3610 381 3646
rect 338 3609 438 3610
rect 338 3588 494 3609
rect 338 3570 456 3588
rect 474 3570 494 3588
rect 338 3566 494 3570
rect 433 3550 494 3566
rect 433 3432 490 3451
rect 433 3429 454 3432
rect 339 3414 454 3429
rect 472 3414 490 3432
rect 339 3391 490 3414
rect 339 3355 381 3391
rect 338 3354 438 3355
rect 338 3333 494 3354
rect 338 3315 456 3333
rect 474 3315 494 3333
rect 338 3311 494 3315
rect 433 3295 494 3311
rect 434 2818 491 2837
rect 434 2815 455 2818
rect 340 2800 455 2815
rect 473 2800 491 2818
rect 340 2777 491 2800
rect 340 2741 382 2777
rect 339 2740 439 2741
rect 339 2719 495 2740
rect 339 2701 457 2719
rect 475 2701 495 2719
rect 339 2697 495 2701
rect 434 2681 495 2697
rect 434 2562 491 2581
rect 434 2559 455 2562
rect 340 2544 455 2559
rect 473 2544 491 2562
rect 340 2521 491 2544
rect 340 2485 382 2521
rect 339 2484 439 2485
rect 339 2463 495 2484
rect 339 2445 457 2463
rect 475 2445 495 2463
rect 339 2441 495 2445
rect 434 2425 495 2441
rect 434 2167 491 2186
rect 434 2164 455 2167
rect 340 2149 455 2164
rect 473 2149 491 2167
rect 340 2126 491 2149
rect 340 2090 382 2126
rect 339 2089 439 2090
rect 339 2068 495 2089
rect 339 2050 457 2068
rect 475 2050 495 2068
rect 339 2046 495 2050
rect 434 2030 495 2046
rect 434 1912 491 1931
rect 434 1909 455 1912
rect 340 1894 455 1909
rect 473 1894 491 1912
rect 340 1871 491 1894
rect 340 1835 382 1871
rect 339 1834 439 1835
rect 339 1813 495 1834
rect 339 1795 457 1813
rect 475 1795 495 1813
rect 339 1791 495 1795
rect 434 1775 495 1791
rect 434 1371 491 1390
rect 434 1368 455 1371
rect 340 1353 455 1368
rect 473 1353 491 1371
rect 340 1330 491 1353
rect 340 1294 382 1330
rect 339 1293 439 1294
rect 339 1272 495 1293
rect 339 1254 457 1272
rect 475 1254 495 1272
rect 339 1250 495 1254
rect 434 1234 495 1250
rect 434 1115 491 1134
rect 434 1112 455 1115
rect 340 1097 455 1112
rect 473 1097 491 1115
rect 340 1074 491 1097
rect 340 1038 382 1074
rect 339 1037 439 1038
rect 339 1016 495 1037
rect 339 998 457 1016
rect 475 998 495 1016
rect 339 994 495 998
rect 434 978 495 994
rect 434 720 491 739
rect 434 717 455 720
rect 340 702 455 717
rect 473 702 491 720
rect 340 679 491 702
rect 340 643 382 679
rect 339 642 439 643
rect 339 621 495 642
rect 339 603 457 621
rect 475 603 495 621
rect 339 599 495 603
rect 434 583 495 599
rect 434 465 491 484
rect 434 462 455 465
rect 340 447 455 462
rect 473 447 491 465
rect 340 424 491 447
rect 340 388 382 424
rect 339 387 439 388
rect 339 366 495 387
rect 339 348 457 366
rect 475 348 495 366
rect 339 344 495 348
rect 434 328 495 344
<< locali >>
rect 432 5785 491 5975
rect 2809 5966 2874 5977
rect 2809 5918 2822 5966
rect 2859 5918 2874 5966
rect 2809 5905 2874 5918
rect 3022 5868 3733 5870
rect 2395 5867 3733 5868
rect 1345 5866 1417 5867
rect 1344 5858 1443 5866
rect 1344 5855 1396 5858
rect 1344 5820 1352 5855
rect 1377 5820 1396 5855
rect 1421 5847 1443 5858
rect 2394 5859 3733 5867
rect 2394 5856 2446 5859
rect 1421 5846 2288 5847
rect 1421 5820 2289 5846
rect 1344 5810 2289 5820
rect 1344 5808 1443 5810
rect 432 5767 454 5785
rect 472 5767 491 5785
rect 432 5745 491 5767
rect 699 5781 1231 5786
rect 699 5761 1585 5781
rect 1605 5761 1608 5781
rect 2244 5777 2289 5810
rect 2394 5821 2402 5856
rect 2427 5821 2446 5856
rect 2471 5821 3733 5859
rect 2394 5812 3733 5821
rect 2394 5809 2483 5812
rect 3022 5810 3733 5812
rect 699 5757 1608 5761
rect 699 5710 742 5757
rect 1192 5756 1608 5757
rect 2240 5757 2633 5777
rect 2653 5757 2656 5777
rect 1192 5755 1533 5756
rect 849 5724 959 5738
rect 849 5721 892 5724
rect 849 5716 853 5721
rect 687 5709 742 5710
rect 431 5686 742 5709
rect 431 5668 456 5686
rect 474 5674 742 5686
rect 771 5694 853 5716
rect 882 5694 892 5721
rect 920 5697 927 5724
rect 956 5716 959 5724
rect 956 5697 1021 5716
rect 920 5694 1021 5697
rect 771 5692 1021 5694
rect 474 5668 496 5674
rect 431 5529 496 5668
rect 771 5613 808 5692
rect 849 5679 959 5692
rect 923 5623 954 5624
rect 771 5593 780 5613
rect 800 5593 808 5613
rect 431 5511 454 5529
rect 472 5511 496 5529
rect 431 5494 496 5511
rect 651 5575 719 5588
rect 771 5583 808 5593
rect 867 5613 954 5623
rect 867 5593 876 5613
rect 896 5593 954 5613
rect 867 5584 954 5593
rect 867 5583 904 5584
rect 651 5533 658 5575
rect 707 5533 719 5575
rect 651 5530 719 5533
rect 923 5531 954 5584
rect 984 5613 1021 5692
rect 1136 5623 1167 5624
rect 984 5593 993 5613
rect 1013 5593 1021 5613
rect 984 5583 1021 5593
rect 1080 5616 1167 5623
rect 1080 5613 1141 5616
rect 1080 5593 1089 5613
rect 1109 5596 1141 5613
rect 1162 5596 1167 5616
rect 1109 5593 1167 5596
rect 1080 5586 1167 5593
rect 1192 5613 1229 5755
rect 1495 5754 1532 5755
rect 2240 5752 2656 5757
rect 2240 5751 2581 5752
rect 1897 5720 2007 5734
rect 1897 5717 1940 5720
rect 1897 5712 1901 5717
rect 1819 5690 1901 5712
rect 1930 5690 1940 5717
rect 1968 5693 1975 5720
rect 2004 5712 2007 5720
rect 2004 5693 2069 5712
rect 1968 5690 2069 5693
rect 1819 5688 2069 5690
rect 1344 5623 1380 5624
rect 1192 5593 1201 5613
rect 1221 5593 1229 5613
rect 1080 5584 1136 5586
rect 1080 5583 1117 5584
rect 1192 5583 1229 5593
rect 1288 5613 1436 5623
rect 1536 5620 1632 5622
rect 1288 5593 1297 5613
rect 1317 5593 1407 5613
rect 1427 5593 1436 5613
rect 1288 5587 1436 5593
rect 1288 5584 1352 5587
rect 1288 5583 1325 5584
rect 1344 5557 1352 5584
rect 1373 5584 1436 5587
rect 1494 5613 1632 5620
rect 1494 5593 1503 5613
rect 1523 5593 1632 5613
rect 1494 5584 1632 5593
rect 1819 5609 1856 5688
rect 1897 5675 2007 5688
rect 1971 5619 2002 5620
rect 1819 5589 1828 5609
rect 1848 5589 1856 5609
rect 1373 5557 1380 5584
rect 1399 5583 1436 5584
rect 1495 5583 1532 5584
rect 1344 5532 1380 5557
rect 815 5530 856 5531
rect 651 5523 856 5530
rect 651 5512 825 5523
rect 651 5479 659 5512
rect 652 5470 659 5479
rect 708 5503 825 5512
rect 845 5503 856 5523
rect 708 5495 856 5503
rect 923 5527 1282 5531
rect 923 5522 1245 5527
rect 923 5498 1036 5522
rect 1060 5503 1245 5522
rect 1269 5503 1282 5527
rect 1060 5498 1282 5503
rect 923 5495 1282 5498
rect 1344 5495 1379 5532
rect 1447 5529 1547 5532
rect 1447 5525 1514 5529
rect 1447 5499 1459 5525
rect 1485 5503 1514 5525
rect 1540 5503 1547 5529
rect 1485 5499 1547 5503
rect 1447 5495 1547 5499
rect 708 5479 719 5495
rect 708 5470 716 5479
rect 923 5474 954 5495
rect 1344 5474 1380 5495
rect 766 5473 803 5474
rect 431 5430 496 5449
rect 431 5412 456 5430
rect 474 5412 496 5430
rect 431 5211 496 5412
rect 652 5286 716 5470
rect 765 5464 803 5473
rect 765 5444 774 5464
rect 794 5444 803 5464
rect 765 5436 803 5444
rect 869 5468 954 5474
rect 979 5473 1016 5474
rect 869 5448 877 5468
rect 897 5448 954 5468
rect 869 5440 954 5448
rect 978 5464 1016 5473
rect 978 5444 987 5464
rect 1007 5444 1016 5464
rect 869 5439 905 5440
rect 978 5436 1016 5444
rect 1082 5468 1167 5474
rect 1187 5473 1224 5474
rect 1082 5448 1090 5468
rect 1110 5467 1167 5468
rect 1110 5448 1139 5467
rect 1082 5447 1139 5448
rect 1160 5447 1167 5467
rect 1082 5440 1167 5447
rect 1186 5464 1224 5473
rect 1186 5444 1195 5464
rect 1215 5444 1224 5464
rect 1082 5439 1118 5440
rect 1186 5436 1224 5444
rect 1290 5468 1434 5474
rect 1290 5448 1298 5468
rect 1318 5448 1406 5468
rect 1426 5448 1434 5468
rect 1290 5440 1434 5448
rect 1290 5439 1326 5440
rect 1398 5439 1434 5440
rect 1500 5473 1537 5474
rect 1500 5472 1538 5473
rect 1500 5464 1564 5472
rect 1500 5444 1509 5464
rect 1529 5450 1564 5464
rect 1584 5450 1587 5470
rect 1529 5445 1587 5450
rect 1529 5444 1564 5445
rect 766 5407 803 5436
rect 767 5405 803 5407
rect 979 5405 1016 5436
rect 767 5383 1016 5405
rect 848 5377 959 5383
rect 848 5369 889 5377
rect 848 5349 856 5369
rect 875 5349 889 5369
rect 848 5347 889 5349
rect 917 5369 959 5377
rect 917 5349 933 5369
rect 952 5349 959 5369
rect 917 5347 959 5349
rect 848 5332 959 5347
rect 652 5276 720 5286
rect 652 5243 669 5276
rect 709 5243 720 5276
rect 652 5231 720 5243
rect 652 5229 716 5231
rect 1187 5212 1224 5436
rect 1500 5432 1564 5444
rect 1604 5214 1631 5584
rect 1819 5579 1856 5589
rect 1915 5609 2002 5619
rect 1915 5589 1924 5609
rect 1944 5589 2002 5609
rect 1915 5580 2002 5589
rect 1915 5579 1952 5580
rect 1695 5566 1765 5571
rect 1690 5560 1765 5566
rect 1690 5527 1698 5560
rect 1751 5527 1765 5560
rect 1971 5527 2002 5580
rect 2032 5609 2069 5688
rect 2184 5619 2215 5620
rect 2032 5589 2041 5609
rect 2061 5589 2069 5609
rect 2032 5579 2069 5589
rect 2128 5612 2215 5619
rect 2128 5609 2189 5612
rect 2128 5589 2137 5609
rect 2157 5592 2189 5609
rect 2210 5592 2215 5612
rect 2157 5589 2215 5592
rect 2128 5582 2215 5589
rect 2240 5609 2277 5751
rect 2543 5750 2580 5751
rect 2392 5619 2428 5620
rect 2240 5589 2249 5609
rect 2269 5589 2277 5609
rect 2128 5580 2184 5582
rect 2128 5579 2165 5580
rect 2240 5579 2277 5589
rect 2336 5609 2484 5619
rect 2584 5616 2680 5618
rect 2336 5589 2345 5609
rect 2365 5589 2455 5609
rect 2475 5589 2484 5609
rect 2336 5583 2484 5589
rect 2336 5580 2400 5583
rect 2336 5579 2373 5580
rect 2392 5553 2400 5580
rect 2421 5580 2484 5583
rect 2542 5609 2680 5616
rect 2542 5589 2551 5609
rect 2571 5589 2680 5609
rect 2542 5580 2680 5589
rect 2421 5553 2428 5580
rect 2447 5579 2484 5580
rect 2543 5579 2580 5580
rect 2392 5528 2428 5553
rect 1690 5526 1773 5527
rect 1863 5526 1904 5527
rect 1690 5519 1904 5526
rect 1690 5502 1873 5519
rect 1690 5469 1703 5502
rect 1756 5499 1873 5502
rect 1893 5499 1904 5519
rect 1756 5491 1904 5499
rect 1971 5523 2330 5527
rect 1971 5518 2293 5523
rect 1971 5494 2084 5518
rect 2108 5499 2293 5518
rect 2317 5499 2330 5523
rect 2108 5494 2330 5499
rect 1971 5491 2330 5494
rect 2392 5491 2427 5528
rect 2495 5525 2595 5528
rect 2495 5521 2562 5525
rect 2495 5495 2507 5521
rect 2533 5499 2562 5521
rect 2588 5499 2595 5525
rect 2533 5495 2595 5499
rect 2495 5491 2595 5495
rect 1756 5469 1773 5491
rect 1971 5470 2002 5491
rect 2392 5470 2428 5491
rect 1814 5469 1851 5470
rect 1690 5455 1773 5469
rect 1463 5212 1631 5214
rect 1187 5211 1631 5212
rect 431 5181 1631 5211
rect 1701 5245 1773 5455
rect 1813 5460 1851 5469
rect 1813 5440 1822 5460
rect 1842 5440 1851 5460
rect 1813 5432 1851 5440
rect 1917 5464 2002 5470
rect 2027 5469 2064 5470
rect 1917 5444 1925 5464
rect 1945 5444 2002 5464
rect 1917 5436 2002 5444
rect 2026 5460 2064 5469
rect 2026 5440 2035 5460
rect 2055 5440 2064 5460
rect 1917 5435 1953 5436
rect 2026 5432 2064 5440
rect 2130 5464 2215 5470
rect 2235 5469 2272 5470
rect 2130 5444 2138 5464
rect 2158 5463 2215 5464
rect 2158 5444 2187 5463
rect 2130 5443 2187 5444
rect 2208 5443 2215 5463
rect 2130 5436 2215 5443
rect 2234 5460 2272 5469
rect 2234 5440 2243 5460
rect 2263 5440 2272 5460
rect 2130 5435 2166 5436
rect 2234 5432 2272 5440
rect 2338 5464 2482 5470
rect 2338 5444 2346 5464
rect 2366 5444 2454 5464
rect 2474 5444 2482 5464
rect 2338 5436 2482 5444
rect 2338 5435 2374 5436
rect 2446 5435 2482 5436
rect 2548 5469 2585 5470
rect 2548 5468 2586 5469
rect 2548 5460 2612 5468
rect 2548 5440 2557 5460
rect 2577 5446 2612 5460
rect 2632 5446 2635 5466
rect 2577 5441 2635 5446
rect 2577 5440 2612 5441
rect 1814 5403 1851 5432
rect 1815 5401 1851 5403
rect 2027 5401 2064 5432
rect 1815 5379 2064 5401
rect 1896 5373 2007 5379
rect 1896 5365 1937 5373
rect 1896 5345 1904 5365
rect 1923 5345 1937 5365
rect 1896 5343 1937 5345
rect 1965 5365 2007 5373
rect 1965 5345 1981 5365
rect 2000 5345 2007 5365
rect 1965 5343 2007 5345
rect 1896 5328 2007 5343
rect 1701 5206 1720 5245
rect 1765 5206 1773 5245
rect 1701 5189 1773 5206
rect 2235 5233 2272 5432
rect 2548 5428 2612 5440
rect 2235 5227 2276 5233
rect 2652 5229 2679 5580
rect 2974 5567 3069 5593
rect 2810 5545 2874 5564
rect 2810 5506 2823 5545
rect 2857 5506 2874 5545
rect 2810 5487 2874 5506
rect 2511 5227 2679 5229
rect 2235 5201 2679 5227
rect 431 5134 496 5181
rect 431 5116 454 5134
rect 472 5116 496 5134
rect 1344 5161 1379 5163
rect 1344 5159 1448 5161
rect 2237 5159 2276 5201
rect 2511 5200 2679 5201
rect 1344 5152 2278 5159
rect 1344 5151 1395 5152
rect 1344 5131 1347 5151
rect 1372 5132 1395 5151
rect 1427 5132 2278 5152
rect 1372 5131 2278 5132
rect 1344 5124 2278 5131
rect 1617 5123 2278 5124
rect 431 5095 496 5116
rect 708 5106 748 5109
rect 708 5102 1611 5106
rect 708 5082 1585 5102
rect 1605 5082 1611 5102
rect 708 5079 1611 5082
rect 432 5035 497 5055
rect 432 5017 456 5035
rect 474 5017 497 5035
rect 432 4990 497 5017
rect 708 4990 748 5079
rect 1192 5077 1608 5079
rect 1192 5076 1533 5077
rect 849 5045 959 5059
rect 849 5042 892 5045
rect 849 5037 853 5042
rect 431 4955 748 4990
rect 771 5015 853 5037
rect 882 5015 892 5042
rect 920 5018 927 5045
rect 956 5037 959 5045
rect 956 5018 1021 5037
rect 920 5015 1021 5018
rect 771 5013 1021 5015
rect 432 4879 497 4955
rect 771 4934 808 5013
rect 849 5000 959 5013
rect 923 4944 954 4945
rect 771 4914 780 4934
rect 800 4914 808 4934
rect 771 4904 808 4914
rect 867 4934 954 4944
rect 867 4914 876 4934
rect 896 4914 954 4934
rect 867 4905 954 4914
rect 867 4904 904 4905
rect 432 4861 454 4879
rect 472 4861 497 4879
rect 432 4840 497 4861
rect 645 4859 710 4868
rect 645 4822 655 4859
rect 695 4851 710 4859
rect 923 4852 954 4905
rect 984 4934 1021 5013
rect 1136 4944 1167 4945
rect 984 4914 993 4934
rect 1013 4914 1021 4934
rect 984 4904 1021 4914
rect 1080 4937 1167 4944
rect 1080 4934 1141 4937
rect 1080 4914 1089 4934
rect 1109 4917 1141 4934
rect 1162 4917 1167 4937
rect 1109 4914 1167 4917
rect 1080 4907 1167 4914
rect 1192 4934 1229 5076
rect 1495 5075 1532 5076
rect 2812 5016 2874 5487
rect 2974 5526 3000 5567
rect 3036 5526 3069 5567
rect 2974 5230 3069 5526
rect 2974 5186 2989 5230
rect 3049 5186 3069 5230
rect 2974 5166 3069 5186
rect 3686 5097 3729 5810
rect 3686 5077 4080 5097
rect 4100 5077 4103 5097
rect 3687 5072 4103 5077
rect 3687 5071 4028 5072
rect 3344 5040 3454 5054
rect 3344 5037 3387 5040
rect 3344 5032 3348 5037
rect 2807 4964 2882 5016
rect 3266 5010 3348 5032
rect 3377 5010 3387 5037
rect 3415 5013 3422 5040
rect 3451 5032 3454 5040
rect 3451 5013 3516 5032
rect 3415 5010 3516 5013
rect 3266 5008 3516 5010
rect 3176 4964 3222 4965
rect 1344 4944 1380 4945
rect 1192 4914 1201 4934
rect 1221 4914 1229 4934
rect 1080 4905 1136 4907
rect 1080 4904 1117 4905
rect 1192 4904 1229 4914
rect 1288 4934 1436 4944
rect 1536 4941 1632 4943
rect 1288 4914 1297 4934
rect 1317 4914 1407 4934
rect 1427 4914 1436 4934
rect 1288 4908 1436 4914
rect 1288 4905 1352 4908
rect 1288 4904 1325 4905
rect 1344 4878 1352 4905
rect 1373 4905 1436 4908
rect 1494 4934 1632 4941
rect 1494 4914 1503 4934
rect 1523 4914 1632 4934
rect 1494 4905 1632 4914
rect 2807 4929 3222 4964
rect 1373 4878 1380 4905
rect 1399 4904 1436 4905
rect 1495 4904 1532 4905
rect 1344 4853 1380 4878
rect 815 4851 856 4852
rect 695 4844 856 4851
rect 695 4824 825 4844
rect 845 4824 856 4844
rect 695 4822 856 4824
rect 645 4816 856 4822
rect 923 4848 1282 4852
rect 923 4843 1245 4848
rect 923 4819 1036 4843
rect 1060 4824 1245 4843
rect 1269 4824 1282 4848
rect 1060 4819 1282 4824
rect 923 4816 1282 4819
rect 1344 4816 1379 4853
rect 1447 4850 1547 4853
rect 1447 4846 1514 4850
rect 1447 4820 1459 4846
rect 1485 4824 1514 4846
rect 1540 4824 1547 4850
rect 1485 4820 1547 4824
rect 1447 4816 1547 4820
rect 645 4803 712 4816
rect 437 4780 493 4800
rect 437 4762 456 4780
rect 474 4762 493 4780
rect 437 4649 493 4762
rect 645 4782 659 4803
rect 695 4782 712 4803
rect 923 4795 954 4816
rect 1344 4795 1380 4816
rect 766 4794 803 4795
rect 645 4775 712 4782
rect 765 4785 803 4794
rect 437 4511 492 4649
rect 645 4623 710 4775
rect 765 4765 774 4785
rect 794 4765 803 4785
rect 765 4757 803 4765
rect 869 4789 954 4795
rect 979 4794 1016 4795
rect 869 4769 877 4789
rect 897 4769 954 4789
rect 869 4761 954 4769
rect 978 4785 1016 4794
rect 978 4765 987 4785
rect 1007 4765 1016 4785
rect 869 4760 905 4761
rect 978 4757 1016 4765
rect 1082 4789 1167 4795
rect 1187 4794 1224 4795
rect 1082 4769 1090 4789
rect 1110 4788 1167 4789
rect 1110 4769 1139 4788
rect 1082 4768 1139 4769
rect 1160 4768 1167 4788
rect 1082 4761 1167 4768
rect 1186 4785 1224 4794
rect 1186 4765 1195 4785
rect 1215 4765 1224 4785
rect 1082 4760 1118 4761
rect 1186 4757 1224 4765
rect 1290 4789 1434 4795
rect 1290 4769 1298 4789
rect 1318 4769 1406 4789
rect 1426 4769 1434 4789
rect 1290 4761 1434 4769
rect 1290 4760 1326 4761
rect 1398 4760 1434 4761
rect 1500 4794 1537 4795
rect 1500 4793 1538 4794
rect 1500 4785 1564 4793
rect 1500 4765 1509 4785
rect 1529 4771 1564 4785
rect 1584 4771 1587 4791
rect 1529 4766 1587 4771
rect 1529 4765 1564 4766
rect 766 4728 803 4757
rect 767 4726 803 4728
rect 979 4726 1016 4757
rect 767 4704 1016 4726
rect 848 4698 959 4704
rect 848 4690 889 4698
rect 848 4670 856 4690
rect 875 4670 889 4690
rect 848 4668 889 4670
rect 917 4690 959 4698
rect 917 4670 933 4690
rect 952 4670 959 4690
rect 917 4668 959 4670
rect 848 4655 959 4668
rect 1187 4658 1224 4757
rect 1500 4753 1564 4765
rect 638 4613 759 4623
rect 638 4611 707 4613
rect 638 4570 651 4611
rect 688 4572 707 4611
rect 744 4572 759 4613
rect 688 4570 759 4572
rect 638 4552 759 4570
rect 430 4508 494 4511
rect 850 4508 954 4514
rect 1185 4508 1226 4658
rect 1604 4650 1631 4905
rect 1693 4895 1773 4906
rect 1693 4869 1710 4895
rect 1750 4869 1773 4895
rect 1693 4842 1773 4869
rect 1693 4816 1714 4842
rect 1754 4816 1773 4842
rect 1693 4797 1773 4816
rect 1693 4771 1717 4797
rect 1757 4771 1773 4797
rect 1693 4720 1773 4771
rect 430 4505 1226 4508
rect 1605 4519 1631 4650
rect 1605 4505 1633 4519
rect 430 4470 1633 4505
rect 1695 4512 1765 4720
rect 2807 4645 2882 4929
rect 3176 4846 3222 4929
rect 3266 4929 3303 5008
rect 3344 4995 3454 5008
rect 3418 4939 3449 4940
rect 3266 4909 3275 4929
rect 3295 4909 3303 4929
rect 3266 4899 3303 4909
rect 3362 4929 3449 4939
rect 3362 4909 3371 4929
rect 3391 4909 3449 4929
rect 3362 4900 3449 4909
rect 3362 4899 3399 4900
rect 3418 4847 3449 4900
rect 3479 4929 3516 5008
rect 3631 4939 3662 4940
rect 3479 4909 3488 4929
rect 3508 4909 3516 4929
rect 3479 4899 3516 4909
rect 3575 4932 3662 4939
rect 3575 4929 3636 4932
rect 3575 4909 3584 4929
rect 3604 4912 3636 4929
rect 3657 4912 3662 4932
rect 3604 4909 3662 4912
rect 3575 4902 3662 4909
rect 3687 4929 3724 5071
rect 3990 5070 4027 5071
rect 3839 4939 3875 4940
rect 3687 4909 3696 4929
rect 3716 4909 3724 4929
rect 3575 4900 3631 4902
rect 3575 4899 3612 4900
rect 3687 4899 3724 4909
rect 3783 4929 3931 4939
rect 4031 4936 4127 4938
rect 3783 4909 3792 4929
rect 3812 4909 3902 4929
rect 3922 4909 3931 4929
rect 3783 4903 3931 4909
rect 3783 4900 3847 4903
rect 3783 4899 3820 4900
rect 3839 4873 3847 4900
rect 3868 4900 3931 4903
rect 3989 4929 4127 4936
rect 3989 4909 3998 4929
rect 4018 4909 4127 4929
rect 3989 4900 4127 4909
rect 3868 4873 3875 4900
rect 3894 4899 3931 4900
rect 3990 4899 4027 4900
rect 3839 4848 3875 4873
rect 3310 4846 3351 4847
rect 3176 4839 3351 4846
rect 2974 4813 3060 4832
rect 2974 4772 2989 4813
rect 3043 4772 3060 4813
rect 3176 4819 3320 4839
rect 3340 4819 3351 4839
rect 3176 4811 3351 4819
rect 3418 4843 3777 4847
rect 3418 4838 3740 4843
rect 3418 4814 3531 4838
rect 3555 4819 3740 4838
rect 3764 4819 3777 4843
rect 3555 4814 3777 4819
rect 3418 4811 3777 4814
rect 3839 4811 3874 4848
rect 3942 4845 4042 4848
rect 3942 4841 4009 4845
rect 3942 4815 3954 4841
rect 3980 4819 4009 4841
rect 4035 4819 4042 4845
rect 3980 4815 4042 4819
rect 3942 4811 4042 4815
rect 3176 4807 3222 4811
rect 3418 4790 3449 4811
rect 3839 4790 3875 4811
rect 3261 4789 3298 4790
rect 2974 4736 3060 4772
rect 3260 4780 3298 4789
rect 3260 4760 3269 4780
rect 3289 4760 3298 4780
rect 3260 4752 3298 4760
rect 3364 4784 3449 4790
rect 3474 4789 3511 4790
rect 3364 4764 3372 4784
rect 3392 4764 3449 4784
rect 3364 4756 3449 4764
rect 3473 4780 3511 4789
rect 3473 4760 3482 4780
rect 3502 4760 3511 4780
rect 3364 4755 3400 4756
rect 3473 4752 3511 4760
rect 3577 4784 3662 4790
rect 3682 4789 3719 4790
rect 3577 4764 3585 4784
rect 3605 4783 3662 4784
rect 3605 4764 3634 4783
rect 3577 4763 3634 4764
rect 3655 4763 3662 4783
rect 3577 4756 3662 4763
rect 3681 4780 3719 4789
rect 3681 4760 3690 4780
rect 3710 4760 3719 4780
rect 3577 4755 3613 4756
rect 3681 4752 3719 4760
rect 3785 4784 3929 4790
rect 3785 4764 3793 4784
rect 3813 4764 3901 4784
rect 3921 4764 3929 4784
rect 3785 4756 3929 4764
rect 3785 4755 3821 4756
rect 430 4409 494 4470
rect 850 4468 954 4470
rect 1185 4468 1226 4470
rect 1695 4467 1716 4512
rect 1696 4446 1716 4467
rect 1746 4467 1765 4512
rect 2802 4603 2882 4645
rect 1746 4446 1763 4467
rect 1696 4427 1763 4446
rect 1345 4419 1417 4420
rect 1344 4411 1443 4419
rect 432 4338 491 4409
rect 1344 4408 1396 4411
rect 1344 4373 1352 4408
rect 1377 4373 1396 4408
rect 1421 4400 1443 4411
rect 1421 4399 2288 4400
rect 1421 4373 2289 4399
rect 1344 4363 2289 4373
rect 1344 4361 1443 4363
rect 432 4320 454 4338
rect 472 4320 491 4338
rect 432 4298 491 4320
rect 699 4334 1231 4339
rect 699 4314 1585 4334
rect 1605 4314 1608 4334
rect 2244 4330 2289 4363
rect 699 4310 1608 4314
rect 699 4263 742 4310
rect 1192 4309 1608 4310
rect 2240 4310 2633 4330
rect 2653 4310 2656 4330
rect 1192 4308 1533 4309
rect 849 4277 959 4291
rect 849 4274 892 4277
rect 849 4269 853 4274
rect 687 4262 742 4263
rect 431 4239 742 4262
rect 431 4221 456 4239
rect 474 4227 742 4239
rect 771 4247 853 4269
rect 882 4247 892 4274
rect 920 4250 927 4277
rect 956 4269 959 4277
rect 956 4250 1021 4269
rect 920 4247 1021 4250
rect 771 4245 1021 4247
rect 474 4221 496 4227
rect 431 4082 496 4221
rect 771 4166 808 4245
rect 849 4232 959 4245
rect 923 4176 954 4177
rect 771 4146 780 4166
rect 800 4146 808 4166
rect 431 4064 454 4082
rect 472 4064 496 4082
rect 431 4047 496 4064
rect 651 4128 719 4141
rect 771 4136 808 4146
rect 867 4166 954 4176
rect 867 4146 876 4166
rect 896 4146 954 4166
rect 867 4137 954 4146
rect 867 4136 904 4137
rect 651 4086 658 4128
rect 707 4086 719 4128
rect 651 4083 719 4086
rect 923 4084 954 4137
rect 984 4166 1021 4245
rect 1136 4176 1167 4177
rect 984 4146 993 4166
rect 1013 4146 1021 4166
rect 984 4136 1021 4146
rect 1080 4169 1167 4176
rect 1080 4166 1141 4169
rect 1080 4146 1089 4166
rect 1109 4149 1141 4166
rect 1162 4149 1167 4169
rect 1109 4146 1167 4149
rect 1080 4139 1167 4146
rect 1192 4166 1229 4308
rect 1495 4307 1532 4308
rect 2240 4305 2656 4310
rect 2240 4304 2581 4305
rect 1897 4273 2007 4287
rect 1897 4270 1940 4273
rect 1897 4265 1901 4270
rect 1819 4243 1901 4265
rect 1930 4243 1940 4270
rect 1968 4246 1975 4273
rect 2004 4265 2007 4273
rect 2004 4246 2069 4265
rect 1968 4243 2069 4246
rect 1819 4241 2069 4243
rect 1344 4176 1380 4177
rect 1192 4146 1201 4166
rect 1221 4146 1229 4166
rect 1080 4137 1136 4139
rect 1080 4136 1117 4137
rect 1192 4136 1229 4146
rect 1288 4166 1436 4176
rect 1536 4173 1632 4175
rect 1288 4146 1297 4166
rect 1317 4146 1407 4166
rect 1427 4146 1436 4166
rect 1288 4140 1436 4146
rect 1288 4137 1352 4140
rect 1288 4136 1325 4137
rect 1344 4110 1352 4137
rect 1373 4137 1436 4140
rect 1494 4166 1632 4173
rect 1494 4146 1503 4166
rect 1523 4146 1632 4166
rect 1494 4137 1632 4146
rect 1819 4162 1856 4241
rect 1897 4228 2007 4241
rect 1971 4172 2002 4173
rect 1819 4142 1828 4162
rect 1848 4142 1856 4162
rect 1373 4110 1380 4137
rect 1399 4136 1436 4137
rect 1495 4136 1532 4137
rect 1344 4085 1380 4110
rect 815 4083 856 4084
rect 651 4076 856 4083
rect 651 4065 825 4076
rect 651 4032 659 4065
rect 652 4023 659 4032
rect 708 4056 825 4065
rect 845 4056 856 4076
rect 708 4048 856 4056
rect 923 4080 1282 4084
rect 923 4075 1245 4080
rect 923 4051 1036 4075
rect 1060 4056 1245 4075
rect 1269 4056 1282 4080
rect 1060 4051 1282 4056
rect 923 4048 1282 4051
rect 1344 4048 1379 4085
rect 1447 4082 1547 4085
rect 1447 4078 1514 4082
rect 1447 4052 1459 4078
rect 1485 4056 1514 4078
rect 1540 4056 1547 4082
rect 1485 4052 1547 4056
rect 1447 4048 1547 4052
rect 708 4032 719 4048
rect 708 4023 716 4032
rect 923 4027 954 4048
rect 1344 4027 1380 4048
rect 766 4026 803 4027
rect 431 3983 496 4002
rect 431 3965 456 3983
rect 474 3965 496 3983
rect 431 3764 496 3965
rect 652 3839 716 4023
rect 765 4017 803 4026
rect 765 3997 774 4017
rect 794 3997 803 4017
rect 765 3989 803 3997
rect 869 4021 954 4027
rect 979 4026 1016 4027
rect 869 4001 877 4021
rect 897 4001 954 4021
rect 869 3993 954 4001
rect 978 4017 1016 4026
rect 978 3997 987 4017
rect 1007 3997 1016 4017
rect 869 3992 905 3993
rect 978 3989 1016 3997
rect 1082 4021 1167 4027
rect 1187 4026 1224 4027
rect 1082 4001 1090 4021
rect 1110 4020 1167 4021
rect 1110 4001 1139 4020
rect 1082 4000 1139 4001
rect 1160 4000 1167 4020
rect 1082 3993 1167 4000
rect 1186 4017 1224 4026
rect 1186 3997 1195 4017
rect 1215 3997 1224 4017
rect 1082 3992 1118 3993
rect 1186 3989 1224 3997
rect 1290 4021 1434 4027
rect 1290 4001 1298 4021
rect 1318 4001 1406 4021
rect 1426 4001 1434 4021
rect 1290 3993 1434 4001
rect 1290 3992 1326 3993
rect 1398 3992 1434 3993
rect 1500 4026 1537 4027
rect 1500 4025 1538 4026
rect 1500 4017 1564 4025
rect 1500 3997 1509 4017
rect 1529 4003 1564 4017
rect 1584 4003 1587 4023
rect 1529 3998 1587 4003
rect 1529 3997 1564 3998
rect 766 3960 803 3989
rect 767 3958 803 3960
rect 979 3958 1016 3989
rect 767 3936 1016 3958
rect 848 3930 959 3936
rect 848 3922 889 3930
rect 848 3902 856 3922
rect 875 3902 889 3922
rect 848 3900 889 3902
rect 917 3922 959 3930
rect 917 3902 933 3922
rect 952 3902 959 3922
rect 917 3900 959 3902
rect 848 3885 959 3900
rect 652 3829 720 3839
rect 652 3796 669 3829
rect 709 3796 720 3829
rect 652 3784 720 3796
rect 652 3782 716 3784
rect 1187 3765 1224 3989
rect 1500 3985 1564 3997
rect 1604 3767 1631 4137
rect 1819 4132 1856 4142
rect 1915 4162 2002 4172
rect 1915 4142 1924 4162
rect 1944 4142 2002 4162
rect 1915 4133 2002 4142
rect 1915 4132 1952 4133
rect 1695 4119 1765 4124
rect 1690 4113 1765 4119
rect 1690 4080 1698 4113
rect 1751 4080 1765 4113
rect 1971 4080 2002 4133
rect 2032 4162 2069 4241
rect 2184 4172 2215 4173
rect 2032 4142 2041 4162
rect 2061 4142 2069 4162
rect 2032 4132 2069 4142
rect 2128 4165 2215 4172
rect 2128 4162 2189 4165
rect 2128 4142 2137 4162
rect 2157 4145 2189 4162
rect 2210 4145 2215 4165
rect 2157 4142 2215 4145
rect 2128 4135 2215 4142
rect 2240 4162 2277 4304
rect 2543 4303 2580 4304
rect 2392 4172 2428 4173
rect 2240 4142 2249 4162
rect 2269 4142 2277 4162
rect 2128 4133 2184 4135
rect 2128 4132 2165 4133
rect 2240 4132 2277 4142
rect 2336 4162 2484 4172
rect 2584 4169 2680 4171
rect 2336 4142 2345 4162
rect 2365 4142 2455 4162
rect 2475 4142 2484 4162
rect 2336 4136 2484 4142
rect 2336 4133 2400 4136
rect 2336 4132 2373 4133
rect 2392 4106 2400 4133
rect 2421 4133 2484 4136
rect 2542 4162 2680 4169
rect 2542 4142 2551 4162
rect 2571 4142 2680 4162
rect 2542 4133 2680 4142
rect 2421 4106 2428 4133
rect 2447 4132 2484 4133
rect 2543 4132 2580 4133
rect 2392 4081 2428 4106
rect 1690 4079 1773 4080
rect 1863 4079 1904 4080
rect 1690 4072 1904 4079
rect 1690 4055 1873 4072
rect 1690 4022 1703 4055
rect 1756 4052 1873 4055
rect 1893 4052 1904 4072
rect 1756 4044 1904 4052
rect 1971 4076 2330 4080
rect 1971 4071 2293 4076
rect 1971 4047 2084 4071
rect 2108 4052 2293 4071
rect 2317 4052 2330 4076
rect 2108 4047 2330 4052
rect 1971 4044 2330 4047
rect 2392 4044 2427 4081
rect 2495 4078 2595 4081
rect 2495 4074 2562 4078
rect 2495 4048 2507 4074
rect 2533 4052 2562 4074
rect 2588 4052 2595 4078
rect 2533 4048 2595 4052
rect 2495 4044 2595 4048
rect 1756 4022 1773 4044
rect 1971 4023 2002 4044
rect 2392 4023 2428 4044
rect 1814 4022 1851 4023
rect 1690 4008 1773 4022
rect 1463 3765 1631 3767
rect 1187 3764 1631 3765
rect 431 3734 1631 3764
rect 1701 3798 1773 4008
rect 1813 4013 1851 4022
rect 1813 3993 1822 4013
rect 1842 3993 1851 4013
rect 1813 3985 1851 3993
rect 1917 4017 2002 4023
rect 2027 4022 2064 4023
rect 1917 3997 1925 4017
rect 1945 3997 2002 4017
rect 1917 3989 2002 3997
rect 2026 4013 2064 4022
rect 2026 3993 2035 4013
rect 2055 3993 2064 4013
rect 1917 3988 1953 3989
rect 2026 3985 2064 3993
rect 2130 4017 2215 4023
rect 2235 4022 2272 4023
rect 2130 3997 2138 4017
rect 2158 4016 2215 4017
rect 2158 3997 2187 4016
rect 2130 3996 2187 3997
rect 2208 3996 2215 4016
rect 2130 3989 2215 3996
rect 2234 4013 2272 4022
rect 2234 3993 2243 4013
rect 2263 3993 2272 4013
rect 2130 3988 2166 3989
rect 2234 3985 2272 3993
rect 2338 4017 2482 4023
rect 2338 3997 2346 4017
rect 2366 3997 2454 4017
rect 2474 3997 2482 4017
rect 2338 3989 2482 3997
rect 2338 3988 2374 3989
rect 2446 3988 2482 3989
rect 2548 4022 2585 4023
rect 2548 4021 2586 4022
rect 2548 4013 2612 4021
rect 2548 3993 2557 4013
rect 2577 3999 2612 4013
rect 2632 3999 2635 4019
rect 2577 3994 2635 3999
rect 2577 3993 2612 3994
rect 1814 3956 1851 3985
rect 1815 3954 1851 3956
rect 2027 3954 2064 3985
rect 1815 3932 2064 3954
rect 1896 3926 2007 3932
rect 1896 3918 1937 3926
rect 1896 3898 1904 3918
rect 1923 3898 1937 3918
rect 1896 3896 1937 3898
rect 1965 3918 2007 3926
rect 1965 3898 1981 3918
rect 2000 3898 2007 3918
rect 1965 3896 2007 3898
rect 1896 3881 2007 3896
rect 1701 3759 1720 3798
rect 1765 3759 1773 3798
rect 1701 3742 1773 3759
rect 2235 3786 2272 3985
rect 2548 3981 2612 3993
rect 2235 3780 2276 3786
rect 2652 3782 2679 4133
rect 2802 4003 2881 4603
rect 2978 4151 3057 4736
rect 3261 4723 3298 4752
rect 3262 4721 3298 4723
rect 3474 4721 3511 4752
rect 3262 4699 3511 4721
rect 3343 4693 3454 4699
rect 3343 4685 3384 4693
rect 3343 4665 3351 4685
rect 3370 4665 3384 4685
rect 3343 4663 3384 4665
rect 3412 4685 3454 4693
rect 3412 4665 3428 4685
rect 3447 4665 3454 4685
rect 3412 4663 3454 4665
rect 3343 4648 3454 4663
rect 3682 4637 3719 4752
rect 3675 4525 3722 4637
rect 3843 4597 3873 4756
rect 3893 4755 3929 4756
rect 3995 4789 4032 4790
rect 3995 4788 4033 4789
rect 3995 4780 4059 4788
rect 3995 4760 4004 4780
rect 4024 4766 4059 4780
rect 4079 4766 4082 4786
rect 4024 4761 4082 4766
rect 4024 4760 4059 4761
rect 3995 4748 4059 4760
rect 3843 4593 3929 4597
rect 3843 4575 3858 4593
rect 3910 4575 3929 4593
rect 3843 4566 3929 4575
rect 4099 4527 4126 4900
rect 3958 4525 4126 4527
rect 3675 4499 4126 4525
rect 3675 4421 3722 4499
rect 3958 4498 4126 4499
rect 3620 4420 3722 4421
rect 3619 4412 3722 4420
rect 3619 4409 3671 4412
rect 3619 4374 3627 4409
rect 3652 4374 3671 4409
rect 3696 4374 3722 4412
rect 3619 4368 3722 4374
rect 3882 4413 3918 4417
rect 3882 4390 3890 4413
rect 3914 4390 3918 4413
rect 3882 4369 3918 4390
rect 3619 4364 3718 4368
rect 3882 4346 3890 4369
rect 3914 4346 3918 4369
rect 2511 3780 2679 3782
rect 2235 3754 2679 3780
rect 431 3687 496 3734
rect 431 3669 454 3687
rect 472 3669 496 3687
rect 1344 3714 1379 3716
rect 1344 3712 1448 3714
rect 2237 3712 2276 3754
rect 2511 3753 2679 3754
rect 1344 3705 2278 3712
rect 1344 3704 1395 3705
rect 1344 3684 1347 3704
rect 1372 3685 1395 3704
rect 1427 3685 2278 3705
rect 1372 3684 2278 3685
rect 1344 3677 2278 3684
rect 1617 3676 2278 3677
rect 431 3648 496 3669
rect 708 3659 748 3662
rect 708 3655 1611 3659
rect 708 3635 1585 3655
rect 1605 3635 1611 3655
rect 708 3632 1611 3635
rect 432 3588 497 3608
rect 432 3570 456 3588
rect 474 3570 497 3588
rect 432 3543 497 3570
rect 708 3543 748 3632
rect 1192 3630 1608 3632
rect 1192 3629 1533 3630
rect 849 3598 959 3612
rect 849 3595 892 3598
rect 849 3590 853 3595
rect 431 3508 748 3543
rect 771 3568 853 3590
rect 882 3568 892 3595
rect 920 3571 927 3598
rect 956 3590 959 3598
rect 956 3571 1021 3590
rect 920 3568 1021 3571
rect 771 3566 1021 3568
rect 432 3432 497 3508
rect 771 3487 808 3566
rect 849 3553 959 3566
rect 923 3497 954 3498
rect 771 3467 780 3487
rect 800 3467 808 3487
rect 771 3457 808 3467
rect 867 3487 954 3497
rect 867 3467 876 3487
rect 896 3467 954 3487
rect 867 3458 954 3467
rect 867 3457 904 3458
rect 432 3414 454 3432
rect 472 3414 497 3432
rect 432 3393 497 3414
rect 645 3412 710 3421
rect 645 3375 655 3412
rect 695 3404 710 3412
rect 923 3405 954 3458
rect 984 3487 1021 3566
rect 1136 3497 1167 3498
rect 984 3467 993 3487
rect 1013 3467 1021 3487
rect 984 3457 1021 3467
rect 1080 3490 1167 3497
rect 1080 3487 1141 3490
rect 1080 3467 1089 3487
rect 1109 3470 1141 3487
rect 1162 3470 1167 3490
rect 1109 3467 1167 3470
rect 1080 3460 1167 3467
rect 1192 3487 1229 3629
rect 1495 3628 1532 3629
rect 1344 3497 1380 3498
rect 1192 3467 1201 3487
rect 1221 3467 1229 3487
rect 1080 3458 1136 3460
rect 1080 3457 1117 3458
rect 1192 3457 1229 3467
rect 1288 3487 1436 3497
rect 1536 3494 1632 3496
rect 1288 3467 1297 3487
rect 1317 3467 1407 3487
rect 1427 3467 1436 3487
rect 1288 3461 1436 3467
rect 1288 3458 1352 3461
rect 1288 3457 1325 3458
rect 1344 3431 1352 3458
rect 1373 3458 1436 3461
rect 1494 3487 1632 3494
rect 1494 3467 1503 3487
rect 1523 3467 1632 3487
rect 1494 3458 1632 3467
rect 1373 3431 1380 3458
rect 1399 3457 1436 3458
rect 1495 3457 1532 3458
rect 1344 3406 1380 3431
rect 815 3404 856 3405
rect 695 3397 856 3404
rect 695 3377 825 3397
rect 845 3377 856 3397
rect 695 3375 856 3377
rect 645 3369 856 3375
rect 923 3401 1282 3405
rect 923 3396 1245 3401
rect 923 3372 1036 3396
rect 1060 3377 1245 3396
rect 1269 3377 1282 3401
rect 1060 3372 1282 3377
rect 923 3369 1282 3372
rect 1344 3369 1379 3406
rect 1447 3403 1547 3406
rect 1447 3399 1514 3403
rect 1447 3373 1459 3399
rect 1485 3377 1514 3399
rect 1540 3377 1547 3403
rect 1485 3373 1547 3377
rect 1447 3369 1547 3373
rect 645 3356 712 3369
rect 437 3333 493 3353
rect 437 3315 456 3333
rect 474 3315 493 3333
rect 437 3202 493 3315
rect 645 3335 659 3356
rect 695 3335 712 3356
rect 923 3348 954 3369
rect 1344 3348 1380 3369
rect 766 3347 803 3348
rect 645 3328 712 3335
rect 765 3338 803 3347
rect 437 3073 492 3202
rect 645 3176 710 3328
rect 765 3318 774 3338
rect 794 3318 803 3338
rect 765 3310 803 3318
rect 869 3342 954 3348
rect 979 3347 1016 3348
rect 869 3322 877 3342
rect 897 3322 954 3342
rect 869 3314 954 3322
rect 978 3338 1016 3347
rect 978 3318 987 3338
rect 1007 3318 1016 3338
rect 869 3313 905 3314
rect 978 3310 1016 3318
rect 1082 3342 1167 3348
rect 1187 3347 1224 3348
rect 1082 3322 1090 3342
rect 1110 3341 1167 3342
rect 1110 3322 1139 3341
rect 1082 3321 1139 3322
rect 1160 3321 1167 3341
rect 1082 3314 1167 3321
rect 1186 3338 1224 3347
rect 1186 3318 1195 3338
rect 1215 3318 1224 3338
rect 1082 3313 1118 3314
rect 1186 3310 1224 3318
rect 1290 3342 1434 3348
rect 1290 3322 1298 3342
rect 1318 3322 1406 3342
rect 1426 3322 1434 3342
rect 1290 3314 1434 3322
rect 1290 3313 1326 3314
rect 1398 3313 1434 3314
rect 1500 3347 1537 3348
rect 1500 3346 1538 3347
rect 1500 3338 1564 3346
rect 1500 3318 1509 3338
rect 1529 3324 1564 3338
rect 1584 3324 1587 3344
rect 1529 3319 1587 3324
rect 1529 3318 1564 3319
rect 766 3281 803 3310
rect 767 3279 803 3281
rect 979 3279 1016 3310
rect 767 3257 1016 3279
rect 848 3251 959 3257
rect 848 3243 889 3251
rect 848 3223 856 3243
rect 875 3223 889 3243
rect 848 3221 889 3223
rect 917 3243 959 3251
rect 917 3223 933 3243
rect 952 3223 959 3243
rect 917 3221 959 3223
rect 848 3206 959 3221
rect 1187 3211 1224 3310
rect 1500 3306 1564 3318
rect 850 3197 954 3206
rect 638 3166 759 3176
rect 638 3164 707 3166
rect 638 3123 651 3164
rect 688 3125 707 3164
rect 744 3125 759 3166
rect 688 3123 759 3125
rect 638 3105 759 3123
rect 431 3061 492 3073
rect 1185 3061 1226 3211
rect 1604 3203 1631 3458
rect 1693 3448 1773 3459
rect 1693 3422 1710 3448
rect 1750 3422 1773 3448
rect 1693 3395 1773 3422
rect 1693 3369 1714 3395
rect 1754 3369 1773 3395
rect 1693 3350 1773 3369
rect 1693 3324 1717 3350
rect 1757 3324 1773 3350
rect 1693 3273 1773 3324
rect 431 3058 1226 3061
rect 1605 3072 1631 3203
rect 1695 3117 1765 3273
rect 1694 3101 1770 3117
rect 1605 3058 1633 3072
rect 431 3023 1633 3058
rect 1694 3064 1709 3101
rect 1753 3064 1770 3101
rect 1694 3044 1770 3064
rect 2808 3094 2878 4003
rect 2977 3402 3058 4151
rect 3882 3848 3918 4346
rect 3806 3819 3919 3848
rect 3806 3652 3837 3819
rect 3730 3632 4123 3652
rect 4143 3632 4146 3652
rect 3730 3627 4146 3632
rect 3730 3626 4071 3627
rect 3387 3595 3497 3609
rect 3387 3592 3430 3595
rect 3387 3587 3391 3592
rect 3309 3565 3391 3587
rect 3420 3565 3430 3592
rect 3458 3568 3465 3595
rect 3494 3587 3497 3595
rect 3494 3568 3559 3587
rect 3458 3565 3559 3568
rect 3309 3563 3559 3565
rect 3309 3484 3346 3563
rect 3387 3550 3497 3563
rect 3461 3494 3492 3495
rect 3309 3464 3318 3484
rect 3338 3464 3346 3484
rect 3309 3454 3346 3464
rect 3405 3484 3492 3494
rect 3405 3464 3414 3484
rect 3434 3464 3492 3484
rect 3405 3455 3492 3464
rect 3405 3454 3442 3455
rect 3461 3402 3492 3455
rect 3522 3484 3559 3563
rect 3674 3494 3705 3495
rect 3522 3464 3531 3484
rect 3551 3464 3559 3484
rect 3522 3454 3559 3464
rect 3618 3487 3705 3494
rect 3618 3484 3679 3487
rect 3618 3464 3627 3484
rect 3647 3467 3679 3484
rect 3700 3467 3705 3487
rect 3647 3464 3705 3467
rect 3618 3457 3705 3464
rect 3730 3484 3767 3626
rect 4033 3625 4070 3626
rect 3882 3494 3918 3495
rect 3730 3464 3739 3484
rect 3759 3464 3767 3484
rect 3618 3455 3674 3457
rect 3618 3454 3655 3455
rect 3730 3454 3767 3464
rect 3826 3484 3974 3494
rect 4074 3491 4170 3493
rect 3826 3464 3835 3484
rect 3855 3464 3945 3484
rect 3965 3464 3974 3484
rect 3826 3458 3974 3464
rect 3826 3455 3890 3458
rect 3826 3454 3863 3455
rect 3882 3428 3890 3455
rect 3911 3455 3974 3458
rect 4032 3484 4170 3491
rect 4032 3464 4041 3484
rect 4061 3464 4170 3484
rect 4032 3455 4170 3464
rect 3911 3428 3918 3455
rect 3937 3454 3974 3455
rect 4033 3454 4070 3455
rect 3882 3403 3918 3428
rect 2977 3401 3311 3402
rect 3353 3401 3394 3402
rect 2977 3394 3394 3401
rect 2977 3374 3363 3394
rect 3383 3374 3394 3394
rect 2977 3366 3394 3374
rect 3461 3398 3820 3402
rect 3461 3393 3783 3398
rect 3461 3369 3574 3393
rect 3598 3374 3783 3393
rect 3807 3374 3820 3398
rect 3598 3369 3820 3374
rect 3461 3366 3820 3369
rect 3882 3366 3917 3403
rect 3985 3400 4085 3403
rect 3985 3396 4052 3400
rect 3985 3370 3997 3396
rect 4023 3374 4052 3396
rect 4078 3374 4085 3400
rect 4023 3370 4085 3374
rect 3985 3366 4085 3370
rect 2977 3362 3311 3366
rect 3461 3345 3492 3366
rect 3882 3345 3918 3366
rect 3304 3344 3341 3345
rect 3303 3335 3341 3344
rect 3303 3315 3312 3335
rect 3332 3315 3341 3335
rect 3303 3307 3341 3315
rect 3407 3339 3492 3345
rect 3517 3344 3554 3345
rect 3407 3319 3415 3339
rect 3435 3319 3492 3339
rect 3407 3311 3492 3319
rect 3516 3335 3554 3344
rect 3516 3315 3525 3335
rect 3545 3315 3554 3335
rect 3407 3310 3443 3311
rect 3516 3307 3554 3315
rect 3620 3339 3705 3345
rect 3725 3344 3762 3345
rect 3620 3319 3628 3339
rect 3648 3338 3705 3339
rect 3648 3319 3677 3338
rect 3620 3318 3677 3319
rect 3698 3318 3705 3338
rect 3620 3311 3705 3318
rect 3724 3335 3762 3344
rect 3724 3315 3733 3335
rect 3753 3315 3762 3335
rect 3620 3310 3656 3311
rect 3724 3307 3762 3315
rect 3828 3339 3972 3345
rect 3828 3319 3836 3339
rect 3856 3319 3944 3339
rect 3964 3319 3972 3339
rect 3828 3311 3972 3319
rect 3828 3310 3864 3311
rect 3936 3310 3972 3311
rect 4038 3344 4075 3345
rect 4038 3343 4076 3344
rect 4038 3335 4102 3343
rect 4038 3315 4047 3335
rect 4067 3321 4102 3335
rect 4122 3321 4125 3341
rect 4067 3316 4125 3321
rect 4067 3315 4102 3316
rect 3304 3278 3341 3307
rect 3305 3276 3341 3278
rect 3517 3276 3554 3307
rect 3305 3254 3554 3276
rect 3386 3248 3497 3254
rect 3386 3240 3427 3248
rect 3386 3220 3394 3240
rect 3413 3220 3427 3240
rect 3386 3218 3427 3220
rect 3455 3240 3497 3248
rect 3455 3220 3471 3240
rect 3490 3220 3497 3240
rect 3455 3218 3497 3220
rect 3386 3203 3497 3218
rect 3725 3186 3762 3307
rect 4038 3303 4102 3315
rect 3843 3186 3872 3190
rect 4142 3188 4169 3455
rect 4001 3186 4169 3188
rect 3725 3160 4169 3186
rect 2808 3044 2880 3094
rect 431 2948 492 3023
rect 850 3021 954 3023
rect 1185 3021 1226 3023
rect 1694 2978 1704 3044
rect 1758 2978 1770 3044
rect 1694 2954 1770 2978
rect 433 2818 492 2948
rect 1346 2899 1418 2900
rect 1345 2891 1444 2899
rect 1345 2888 1397 2891
rect 1345 2853 1353 2888
rect 1378 2853 1397 2888
rect 1422 2880 1444 2891
rect 1422 2879 2289 2880
rect 1422 2853 2290 2879
rect 1345 2843 2290 2853
rect 1345 2841 1444 2843
rect 433 2800 455 2818
rect 473 2800 492 2818
rect 433 2778 492 2800
rect 700 2814 1232 2819
rect 700 2794 1586 2814
rect 1606 2794 1609 2814
rect 2245 2810 2290 2843
rect 700 2790 1609 2794
rect 700 2743 743 2790
rect 1193 2789 1609 2790
rect 2241 2790 2634 2810
rect 2654 2790 2657 2810
rect 1193 2788 1534 2789
rect 850 2757 960 2771
rect 850 2754 893 2757
rect 850 2749 854 2754
rect 688 2742 743 2743
rect 432 2719 743 2742
rect 432 2701 457 2719
rect 475 2707 743 2719
rect 772 2727 854 2749
rect 883 2727 893 2754
rect 921 2730 928 2757
rect 957 2749 960 2757
rect 957 2730 1022 2749
rect 921 2727 1022 2730
rect 772 2725 1022 2727
rect 475 2701 497 2707
rect 432 2562 497 2701
rect 772 2646 809 2725
rect 850 2712 960 2725
rect 924 2656 955 2657
rect 772 2626 781 2646
rect 801 2626 809 2646
rect 432 2544 455 2562
rect 473 2544 497 2562
rect 432 2527 497 2544
rect 652 2608 720 2621
rect 772 2616 809 2626
rect 868 2646 955 2656
rect 868 2626 877 2646
rect 897 2626 955 2646
rect 868 2617 955 2626
rect 868 2616 905 2617
rect 652 2566 659 2608
rect 708 2566 720 2608
rect 652 2563 720 2566
rect 924 2564 955 2617
rect 985 2646 1022 2725
rect 1137 2656 1168 2657
rect 985 2626 994 2646
rect 1014 2626 1022 2646
rect 985 2616 1022 2626
rect 1081 2649 1168 2656
rect 1081 2646 1142 2649
rect 1081 2626 1090 2646
rect 1110 2629 1142 2646
rect 1163 2629 1168 2649
rect 1110 2626 1168 2629
rect 1081 2619 1168 2626
rect 1193 2646 1230 2788
rect 1496 2787 1533 2788
rect 2241 2785 2657 2790
rect 2241 2784 2582 2785
rect 1898 2753 2008 2767
rect 1898 2750 1941 2753
rect 1898 2745 1902 2750
rect 1820 2723 1902 2745
rect 1931 2723 1941 2750
rect 1969 2726 1976 2753
rect 2005 2745 2008 2753
rect 2005 2726 2070 2745
rect 1969 2723 2070 2726
rect 1820 2721 2070 2723
rect 1345 2656 1381 2657
rect 1193 2626 1202 2646
rect 1222 2626 1230 2646
rect 1081 2617 1137 2619
rect 1081 2616 1118 2617
rect 1193 2616 1230 2626
rect 1289 2646 1437 2656
rect 1537 2653 1633 2655
rect 1289 2626 1298 2646
rect 1318 2626 1408 2646
rect 1428 2626 1437 2646
rect 1289 2620 1437 2626
rect 1289 2617 1353 2620
rect 1289 2616 1326 2617
rect 1345 2590 1353 2617
rect 1374 2617 1437 2620
rect 1495 2646 1633 2653
rect 1495 2626 1504 2646
rect 1524 2626 1633 2646
rect 1495 2617 1633 2626
rect 1820 2642 1857 2721
rect 1898 2708 2008 2721
rect 1972 2652 2003 2653
rect 1820 2622 1829 2642
rect 1849 2622 1857 2642
rect 1374 2590 1381 2617
rect 1400 2616 1437 2617
rect 1496 2616 1533 2617
rect 1345 2565 1381 2590
rect 816 2563 857 2564
rect 652 2556 857 2563
rect 652 2545 826 2556
rect 652 2512 660 2545
rect 653 2503 660 2512
rect 709 2536 826 2545
rect 846 2536 857 2556
rect 709 2528 857 2536
rect 924 2560 1283 2564
rect 924 2555 1246 2560
rect 924 2531 1037 2555
rect 1061 2536 1246 2555
rect 1270 2536 1283 2560
rect 1061 2531 1283 2536
rect 924 2528 1283 2531
rect 1345 2528 1380 2565
rect 1448 2562 1548 2565
rect 1448 2558 1515 2562
rect 1448 2532 1460 2558
rect 1486 2536 1515 2558
rect 1541 2536 1548 2562
rect 1486 2532 1548 2536
rect 1448 2528 1548 2532
rect 709 2512 720 2528
rect 709 2503 717 2512
rect 924 2507 955 2528
rect 1345 2507 1381 2528
rect 767 2506 804 2507
rect 432 2463 497 2482
rect 432 2445 457 2463
rect 475 2445 497 2463
rect 432 2244 497 2445
rect 653 2319 717 2503
rect 766 2497 804 2506
rect 766 2477 775 2497
rect 795 2477 804 2497
rect 766 2469 804 2477
rect 870 2501 955 2507
rect 980 2506 1017 2507
rect 870 2481 878 2501
rect 898 2481 955 2501
rect 870 2473 955 2481
rect 979 2497 1017 2506
rect 979 2477 988 2497
rect 1008 2477 1017 2497
rect 870 2472 906 2473
rect 979 2469 1017 2477
rect 1083 2501 1168 2507
rect 1188 2506 1225 2507
rect 1083 2481 1091 2501
rect 1111 2500 1168 2501
rect 1111 2481 1140 2500
rect 1083 2480 1140 2481
rect 1161 2480 1168 2500
rect 1083 2473 1168 2480
rect 1187 2497 1225 2506
rect 1187 2477 1196 2497
rect 1216 2477 1225 2497
rect 1083 2472 1119 2473
rect 1187 2469 1225 2477
rect 1291 2501 1435 2507
rect 1291 2481 1299 2501
rect 1319 2481 1407 2501
rect 1427 2481 1435 2501
rect 1291 2473 1435 2481
rect 1291 2472 1327 2473
rect 1399 2472 1435 2473
rect 1501 2506 1538 2507
rect 1501 2505 1539 2506
rect 1501 2497 1565 2505
rect 1501 2477 1510 2497
rect 1530 2483 1565 2497
rect 1585 2483 1588 2503
rect 1530 2478 1588 2483
rect 1530 2477 1565 2478
rect 767 2440 804 2469
rect 768 2438 804 2440
rect 980 2438 1017 2469
rect 768 2416 1017 2438
rect 849 2410 960 2416
rect 849 2402 890 2410
rect 849 2382 857 2402
rect 876 2382 890 2402
rect 849 2380 890 2382
rect 918 2402 960 2410
rect 918 2382 934 2402
rect 953 2382 960 2402
rect 918 2380 960 2382
rect 849 2365 960 2380
rect 653 2309 721 2319
rect 653 2276 670 2309
rect 710 2276 721 2309
rect 653 2264 721 2276
rect 653 2262 717 2264
rect 1188 2245 1225 2469
rect 1501 2465 1565 2477
rect 1605 2247 1632 2617
rect 1820 2612 1857 2622
rect 1916 2642 2003 2652
rect 1916 2622 1925 2642
rect 1945 2622 2003 2642
rect 1916 2613 2003 2622
rect 1916 2612 1953 2613
rect 1696 2599 1766 2604
rect 1691 2593 1766 2599
rect 1691 2560 1699 2593
rect 1752 2560 1766 2593
rect 1972 2560 2003 2613
rect 2033 2642 2070 2721
rect 2185 2652 2216 2653
rect 2033 2622 2042 2642
rect 2062 2622 2070 2642
rect 2033 2612 2070 2622
rect 2129 2645 2216 2652
rect 2129 2642 2190 2645
rect 2129 2622 2138 2642
rect 2158 2625 2190 2642
rect 2211 2625 2216 2645
rect 2158 2622 2216 2625
rect 2129 2615 2216 2622
rect 2241 2642 2278 2784
rect 2544 2783 2581 2784
rect 2393 2652 2429 2653
rect 2241 2622 2250 2642
rect 2270 2622 2278 2642
rect 2129 2613 2185 2615
rect 2129 2612 2166 2613
rect 2241 2612 2278 2622
rect 2337 2642 2485 2652
rect 2585 2649 2681 2651
rect 2337 2622 2346 2642
rect 2366 2622 2456 2642
rect 2476 2622 2485 2642
rect 2337 2616 2485 2622
rect 2337 2613 2401 2616
rect 2337 2612 2374 2613
rect 2393 2586 2401 2613
rect 2422 2613 2485 2616
rect 2543 2642 2681 2649
rect 2543 2622 2552 2642
rect 2572 2622 2681 2642
rect 2543 2613 2681 2622
rect 2422 2586 2429 2613
rect 2448 2612 2485 2613
rect 2544 2612 2581 2613
rect 2393 2561 2429 2586
rect 1691 2559 1774 2560
rect 1864 2559 1905 2560
rect 1691 2552 1905 2559
rect 1691 2535 1874 2552
rect 1691 2502 1704 2535
rect 1757 2532 1874 2535
rect 1894 2532 1905 2552
rect 1757 2524 1905 2532
rect 1972 2556 2331 2560
rect 1972 2551 2294 2556
rect 1972 2527 2085 2551
rect 2109 2532 2294 2551
rect 2318 2532 2331 2556
rect 2109 2527 2331 2532
rect 1972 2524 2331 2527
rect 2393 2524 2428 2561
rect 2496 2558 2596 2561
rect 2496 2554 2563 2558
rect 2496 2528 2508 2554
rect 2534 2532 2563 2554
rect 2589 2532 2596 2558
rect 2534 2528 2596 2532
rect 2496 2524 2596 2528
rect 1757 2502 1774 2524
rect 1972 2503 2003 2524
rect 2393 2503 2429 2524
rect 1815 2502 1852 2503
rect 1691 2488 1774 2502
rect 1464 2245 1632 2247
rect 1188 2244 1632 2245
rect 432 2214 1632 2244
rect 1702 2278 1774 2488
rect 1814 2493 1852 2502
rect 1814 2473 1823 2493
rect 1843 2473 1852 2493
rect 1814 2465 1852 2473
rect 1918 2497 2003 2503
rect 2028 2502 2065 2503
rect 1918 2477 1926 2497
rect 1946 2477 2003 2497
rect 1918 2469 2003 2477
rect 2027 2493 2065 2502
rect 2027 2473 2036 2493
rect 2056 2473 2065 2493
rect 1918 2468 1954 2469
rect 2027 2465 2065 2473
rect 2131 2497 2216 2503
rect 2236 2502 2273 2503
rect 2131 2477 2139 2497
rect 2159 2496 2216 2497
rect 2159 2477 2188 2496
rect 2131 2476 2188 2477
rect 2209 2476 2216 2496
rect 2131 2469 2216 2476
rect 2235 2493 2273 2502
rect 2235 2473 2244 2493
rect 2264 2473 2273 2493
rect 2131 2468 2167 2469
rect 2235 2465 2273 2473
rect 2339 2497 2483 2503
rect 2339 2477 2347 2497
rect 2367 2477 2455 2497
rect 2475 2477 2483 2497
rect 2339 2469 2483 2477
rect 2339 2468 2375 2469
rect 2447 2468 2483 2469
rect 2549 2502 2586 2503
rect 2549 2501 2587 2502
rect 2549 2493 2613 2501
rect 2549 2473 2558 2493
rect 2578 2479 2613 2493
rect 2633 2479 2636 2499
rect 2578 2474 2636 2479
rect 2578 2473 2613 2474
rect 1815 2436 1852 2465
rect 1816 2434 1852 2436
rect 2028 2434 2065 2465
rect 1816 2412 2065 2434
rect 1897 2406 2008 2412
rect 1897 2398 1938 2406
rect 1897 2378 1905 2398
rect 1924 2378 1938 2398
rect 1897 2376 1938 2378
rect 1966 2398 2008 2406
rect 1966 2378 1982 2398
rect 2001 2378 2008 2398
rect 1966 2376 2008 2378
rect 1897 2361 2008 2376
rect 1702 2239 1721 2278
rect 1766 2239 1774 2278
rect 1702 2222 1774 2239
rect 2236 2266 2273 2465
rect 2549 2461 2613 2473
rect 2236 2260 2277 2266
rect 2653 2262 2680 2613
rect 2809 2565 2880 3044
rect 3684 2892 3729 2901
rect 3684 2854 3694 2892
rect 3719 2854 3729 2892
rect 3684 2843 3729 2854
rect 3687 2835 3729 2843
rect 2809 2481 2878 2565
rect 2512 2260 2680 2262
rect 2236 2234 2680 2260
rect 432 2167 497 2214
rect 432 2149 455 2167
rect 473 2149 497 2167
rect 1345 2194 1380 2196
rect 1345 2192 1449 2194
rect 2238 2192 2277 2234
rect 2512 2233 2680 2234
rect 1345 2185 2279 2192
rect 1345 2184 1396 2185
rect 1345 2164 1348 2184
rect 1373 2165 1396 2184
rect 1428 2165 2279 2185
rect 1373 2164 2279 2165
rect 1345 2157 2279 2164
rect 1618 2156 2279 2157
rect 432 2128 497 2149
rect 709 2139 749 2142
rect 709 2135 1612 2139
rect 709 2115 1586 2135
rect 1606 2115 1612 2135
rect 709 2112 1612 2115
rect 433 2068 498 2088
rect 433 2050 457 2068
rect 475 2050 498 2068
rect 433 2023 498 2050
rect 709 2023 749 2112
rect 1193 2110 1609 2112
rect 1193 2109 1534 2110
rect 850 2078 960 2092
rect 850 2075 893 2078
rect 850 2070 854 2075
rect 432 1988 749 2023
rect 772 2048 854 2070
rect 883 2048 893 2075
rect 921 2051 928 2078
rect 957 2070 960 2078
rect 957 2051 1022 2070
rect 921 2048 1022 2051
rect 772 2046 1022 2048
rect 433 1912 498 1988
rect 772 1967 809 2046
rect 850 2033 960 2046
rect 924 1977 955 1978
rect 772 1947 781 1967
rect 801 1947 809 1967
rect 772 1937 809 1947
rect 868 1967 955 1977
rect 868 1947 877 1967
rect 897 1947 955 1967
rect 868 1938 955 1947
rect 868 1937 905 1938
rect 433 1894 455 1912
rect 473 1894 498 1912
rect 433 1873 498 1894
rect 646 1892 711 1901
rect 646 1855 656 1892
rect 696 1884 711 1892
rect 924 1885 955 1938
rect 985 1967 1022 2046
rect 1137 1977 1168 1978
rect 985 1947 994 1967
rect 1014 1947 1022 1967
rect 985 1937 1022 1947
rect 1081 1970 1168 1977
rect 1081 1967 1142 1970
rect 1081 1947 1090 1967
rect 1110 1950 1142 1967
rect 1163 1950 1168 1970
rect 1110 1947 1168 1950
rect 1081 1940 1168 1947
rect 1193 1967 1230 2109
rect 1496 2108 1533 2109
rect 1345 1977 1381 1978
rect 1193 1947 1202 1967
rect 1222 1947 1230 1967
rect 1081 1938 1137 1940
rect 1081 1937 1118 1938
rect 1193 1937 1230 1947
rect 1289 1967 1437 1977
rect 1537 1974 1633 1976
rect 1289 1947 1298 1967
rect 1318 1947 1408 1967
rect 1428 1947 1437 1967
rect 1289 1941 1437 1947
rect 1289 1938 1353 1941
rect 1289 1937 1326 1938
rect 1345 1911 1353 1938
rect 1374 1938 1437 1941
rect 1495 1967 1633 1974
rect 1495 1947 1504 1967
rect 1524 1947 1633 1967
rect 1495 1938 1633 1947
rect 1374 1911 1381 1938
rect 1400 1937 1437 1938
rect 1496 1937 1533 1938
rect 1345 1886 1381 1911
rect 816 1884 857 1885
rect 696 1877 857 1884
rect 696 1857 826 1877
rect 846 1857 857 1877
rect 696 1855 857 1857
rect 646 1849 857 1855
rect 924 1881 1283 1885
rect 924 1876 1246 1881
rect 924 1852 1037 1876
rect 1061 1857 1246 1876
rect 1270 1857 1283 1881
rect 1061 1852 1283 1857
rect 924 1849 1283 1852
rect 1345 1849 1380 1886
rect 1448 1883 1548 1886
rect 1448 1879 1515 1883
rect 1448 1853 1460 1879
rect 1486 1857 1515 1879
rect 1541 1857 1548 1883
rect 1486 1853 1548 1857
rect 1448 1849 1548 1853
rect 646 1836 713 1849
rect 438 1813 494 1833
rect 438 1795 457 1813
rect 475 1795 494 1813
rect 438 1682 494 1795
rect 646 1815 660 1836
rect 696 1815 713 1836
rect 924 1828 955 1849
rect 1345 1828 1381 1849
rect 767 1827 804 1828
rect 646 1808 713 1815
rect 766 1818 804 1827
rect 438 1544 493 1682
rect 646 1656 711 1808
rect 766 1798 775 1818
rect 795 1798 804 1818
rect 766 1790 804 1798
rect 870 1822 955 1828
rect 980 1827 1017 1828
rect 870 1802 878 1822
rect 898 1802 955 1822
rect 870 1794 955 1802
rect 979 1818 1017 1827
rect 979 1798 988 1818
rect 1008 1798 1017 1818
rect 870 1793 906 1794
rect 979 1790 1017 1798
rect 1083 1822 1168 1828
rect 1188 1827 1225 1828
rect 1083 1802 1091 1822
rect 1111 1821 1168 1822
rect 1111 1802 1140 1821
rect 1083 1801 1140 1802
rect 1161 1801 1168 1821
rect 1083 1794 1168 1801
rect 1187 1818 1225 1827
rect 1187 1798 1196 1818
rect 1216 1798 1225 1818
rect 1083 1793 1119 1794
rect 1187 1790 1225 1798
rect 1291 1822 1435 1828
rect 1291 1802 1299 1822
rect 1319 1802 1407 1822
rect 1427 1802 1435 1822
rect 1291 1794 1435 1802
rect 1291 1793 1327 1794
rect 1399 1793 1435 1794
rect 1501 1827 1538 1828
rect 1501 1826 1539 1827
rect 1501 1818 1565 1826
rect 1501 1798 1510 1818
rect 1530 1804 1565 1818
rect 1585 1804 1588 1824
rect 1530 1799 1588 1804
rect 1530 1798 1565 1799
rect 767 1761 804 1790
rect 768 1759 804 1761
rect 980 1759 1017 1790
rect 768 1737 1017 1759
rect 849 1731 960 1737
rect 849 1723 890 1731
rect 849 1703 857 1723
rect 876 1703 890 1723
rect 849 1701 890 1703
rect 918 1723 960 1731
rect 918 1703 934 1723
rect 953 1703 960 1723
rect 918 1701 960 1703
rect 849 1688 960 1701
rect 1188 1691 1225 1790
rect 1501 1786 1565 1798
rect 639 1646 760 1656
rect 639 1644 708 1646
rect 639 1603 652 1644
rect 689 1605 708 1644
rect 745 1605 760 1646
rect 689 1603 760 1605
rect 639 1585 760 1603
rect 431 1541 495 1544
rect 851 1541 955 1547
rect 1186 1541 1227 1691
rect 1605 1683 1632 1938
rect 1694 1928 1774 1939
rect 2813 1930 2875 2481
rect 3687 2130 3730 2835
rect 3843 2221 3872 3160
rect 4001 3159 4169 3160
rect 3841 2200 3878 2221
rect 3841 2163 3852 2200
rect 3869 2163 3878 2200
rect 3841 2153 3878 2163
rect 3687 2110 4081 2130
rect 4101 2110 4104 2130
rect 3688 2105 4104 2110
rect 3688 2104 4029 2105
rect 3345 2073 3455 2087
rect 3345 2070 3388 2073
rect 3345 2065 3349 2070
rect 3267 2043 3349 2065
rect 3378 2043 3388 2070
rect 3416 2046 3423 2073
rect 3452 2065 3455 2073
rect 3452 2046 3517 2065
rect 3416 2043 3517 2046
rect 3267 2041 3517 2043
rect 3267 1962 3304 2041
rect 3345 2028 3455 2041
rect 3419 1972 3450 1973
rect 3267 1942 3276 1962
rect 3296 1942 3304 1962
rect 3267 1932 3304 1942
rect 3363 1962 3450 1972
rect 3363 1942 3372 1962
rect 3392 1942 3450 1962
rect 3363 1933 3450 1942
rect 3363 1932 3400 1933
rect 1694 1902 1711 1928
rect 1751 1902 1774 1928
rect 1694 1875 1774 1902
rect 1694 1849 1715 1875
rect 1755 1849 1774 1875
rect 1694 1830 1774 1849
rect 1694 1804 1718 1830
rect 1758 1804 1774 1830
rect 2807 1868 2879 1930
rect 3419 1880 3450 1933
rect 3480 1962 3517 2041
rect 3632 1972 3663 1973
rect 3480 1942 3489 1962
rect 3509 1942 3517 1962
rect 3480 1932 3517 1942
rect 3576 1965 3663 1972
rect 3576 1962 3637 1965
rect 3576 1942 3585 1962
rect 3605 1945 3637 1962
rect 3658 1945 3663 1965
rect 3605 1942 3663 1945
rect 3576 1935 3663 1942
rect 3688 1962 3725 2104
rect 3991 2103 4028 2104
rect 3840 1972 3876 1973
rect 3688 1942 3697 1962
rect 3717 1942 3725 1962
rect 3576 1933 3632 1935
rect 3576 1932 3613 1933
rect 3688 1932 3725 1942
rect 3784 1962 3932 1972
rect 4032 1969 4128 1971
rect 3784 1942 3793 1962
rect 3813 1942 3903 1962
rect 3923 1942 3932 1962
rect 3784 1936 3932 1942
rect 3784 1933 3848 1936
rect 3784 1932 3821 1933
rect 3840 1906 3848 1933
rect 3869 1933 3932 1936
rect 3990 1962 4128 1969
rect 3990 1942 3999 1962
rect 4019 1942 4128 1962
rect 3990 1933 4128 1942
rect 3869 1906 3876 1933
rect 3895 1932 3932 1933
rect 3991 1932 4028 1933
rect 3840 1881 3876 1906
rect 3311 1879 3352 1880
rect 3231 1874 3352 1879
rect 2807 1845 2825 1868
rect 2851 1845 2879 1868
rect 2807 1825 2879 1845
rect 3182 1872 3352 1874
rect 3182 1861 3321 1872
rect 3182 1838 3205 1861
rect 3231 1852 3321 1861
rect 3341 1852 3352 1872
rect 3231 1844 3352 1852
rect 3419 1876 3778 1880
rect 3419 1871 3741 1876
rect 3419 1847 3532 1871
rect 3556 1852 3741 1871
rect 3765 1852 3778 1876
rect 3556 1847 3778 1852
rect 3419 1844 3778 1847
rect 3840 1844 3875 1881
rect 3943 1878 4043 1881
rect 3943 1874 4010 1878
rect 3943 1848 3955 1874
rect 3981 1852 4010 1874
rect 4036 1852 4043 1878
rect 3981 1848 4043 1852
rect 3943 1844 4043 1848
rect 3231 1838 3239 1844
rect 3182 1830 3239 1838
rect 3419 1823 3450 1844
rect 3840 1823 3876 1844
rect 3262 1822 3299 1823
rect 1694 1753 1774 1804
rect 3261 1813 3299 1822
rect 3261 1793 3270 1813
rect 3290 1793 3299 1813
rect 3261 1785 3299 1793
rect 3365 1817 3450 1823
rect 3475 1822 3512 1823
rect 3365 1797 3373 1817
rect 3393 1797 3450 1817
rect 3365 1789 3450 1797
rect 3474 1813 3512 1822
rect 3474 1793 3483 1813
rect 3503 1793 3512 1813
rect 3365 1788 3401 1789
rect 3474 1785 3512 1793
rect 3578 1817 3663 1823
rect 3683 1822 3720 1823
rect 3578 1797 3586 1817
rect 3606 1816 3663 1817
rect 3606 1797 3635 1816
rect 3578 1796 3635 1797
rect 3656 1796 3663 1816
rect 3578 1789 3663 1796
rect 3682 1813 3720 1822
rect 3682 1793 3691 1813
rect 3711 1793 3720 1813
rect 3578 1788 3614 1789
rect 3682 1785 3720 1793
rect 3786 1817 3930 1823
rect 3786 1797 3794 1817
rect 3814 1797 3902 1817
rect 3922 1797 3930 1817
rect 3786 1789 3930 1797
rect 3786 1788 3822 1789
rect 3894 1788 3930 1789
rect 3996 1822 4033 1823
rect 3996 1821 4034 1822
rect 3996 1813 4060 1821
rect 3996 1793 4005 1813
rect 4025 1799 4060 1813
rect 4080 1799 4083 1819
rect 4025 1794 4083 1799
rect 4025 1793 4060 1794
rect 3262 1756 3299 1785
rect 3263 1754 3299 1756
rect 3475 1754 3512 1785
rect 431 1538 1227 1541
rect 1606 1552 1632 1683
rect 1606 1538 1634 1552
rect 431 1503 1634 1538
rect 1696 1545 1766 1753
rect 3263 1732 3512 1754
rect 3344 1726 3455 1732
rect 3344 1718 3385 1726
rect 3344 1698 3352 1718
rect 3371 1698 3385 1718
rect 3344 1696 3385 1698
rect 3413 1718 3455 1726
rect 3413 1698 3429 1718
rect 3448 1698 3455 1718
rect 3413 1696 3455 1698
rect 3344 1681 3455 1696
rect 3683 1670 3720 1785
rect 3996 1781 4060 1793
rect 431 1442 495 1503
rect 851 1501 955 1503
rect 1186 1501 1227 1503
rect 1696 1500 1717 1545
rect 1697 1479 1717 1500
rect 1747 1500 1766 1545
rect 3676 1664 3723 1670
rect 4100 1666 4127 1933
rect 3959 1664 4127 1666
rect 3676 1638 4127 1664
rect 3676 1503 3723 1638
rect 3959 1637 4127 1638
rect 1747 1479 1764 1500
rect 1697 1460 1764 1479
rect 3674 1454 3733 1503
rect 1346 1452 1418 1453
rect 1345 1444 1444 1452
rect 433 1371 492 1442
rect 1345 1441 1397 1444
rect 1345 1406 1353 1441
rect 1378 1406 1397 1441
rect 1422 1433 1444 1444
rect 1422 1432 2289 1433
rect 1422 1406 2290 1432
rect 3674 1426 3692 1454
rect 3720 1426 3733 1454
rect 3674 1416 3733 1426
rect 1345 1396 2290 1406
rect 1345 1394 1444 1396
rect 433 1353 455 1371
rect 473 1353 492 1371
rect 433 1331 492 1353
rect 700 1367 1232 1372
rect 700 1347 1586 1367
rect 1606 1347 1609 1367
rect 2245 1363 2290 1396
rect 700 1343 1609 1347
rect 700 1296 743 1343
rect 1193 1342 1609 1343
rect 2241 1343 2634 1363
rect 2654 1343 2657 1363
rect 1193 1341 1534 1342
rect 850 1310 960 1324
rect 850 1307 893 1310
rect 850 1302 854 1307
rect 688 1295 743 1296
rect 432 1272 743 1295
rect 432 1254 457 1272
rect 475 1260 743 1272
rect 772 1280 854 1302
rect 883 1280 893 1307
rect 921 1283 928 1310
rect 957 1302 960 1310
rect 957 1283 1022 1302
rect 921 1280 1022 1283
rect 772 1278 1022 1280
rect 475 1254 497 1260
rect 432 1115 497 1254
rect 772 1199 809 1278
rect 850 1265 960 1278
rect 924 1209 955 1210
rect 772 1179 781 1199
rect 801 1179 809 1199
rect 432 1097 455 1115
rect 473 1097 497 1115
rect 432 1080 497 1097
rect 652 1161 720 1174
rect 772 1169 809 1179
rect 868 1199 955 1209
rect 868 1179 877 1199
rect 897 1179 955 1199
rect 868 1170 955 1179
rect 868 1169 905 1170
rect 652 1119 659 1161
rect 708 1119 720 1161
rect 652 1116 720 1119
rect 924 1117 955 1170
rect 985 1199 1022 1278
rect 1137 1209 1168 1210
rect 985 1179 994 1199
rect 1014 1179 1022 1199
rect 985 1169 1022 1179
rect 1081 1202 1168 1209
rect 1081 1199 1142 1202
rect 1081 1179 1090 1199
rect 1110 1182 1142 1199
rect 1163 1182 1168 1202
rect 1110 1179 1168 1182
rect 1081 1172 1168 1179
rect 1193 1199 1230 1341
rect 1496 1340 1533 1341
rect 2241 1338 2657 1343
rect 2241 1337 2582 1338
rect 1898 1306 2008 1320
rect 1898 1303 1941 1306
rect 1898 1298 1902 1303
rect 1820 1276 1902 1298
rect 1931 1276 1941 1303
rect 1969 1279 1976 1306
rect 2005 1298 2008 1306
rect 2005 1279 2070 1298
rect 1969 1276 2070 1279
rect 1820 1274 2070 1276
rect 1345 1209 1381 1210
rect 1193 1179 1202 1199
rect 1222 1179 1230 1199
rect 1081 1170 1137 1172
rect 1081 1169 1118 1170
rect 1193 1169 1230 1179
rect 1289 1199 1437 1209
rect 1537 1206 1633 1208
rect 1289 1179 1298 1199
rect 1318 1179 1408 1199
rect 1428 1179 1437 1199
rect 1289 1173 1437 1179
rect 1289 1170 1353 1173
rect 1289 1169 1326 1170
rect 1345 1143 1353 1170
rect 1374 1170 1437 1173
rect 1495 1199 1633 1206
rect 1495 1179 1504 1199
rect 1524 1179 1633 1199
rect 1495 1170 1633 1179
rect 1820 1195 1857 1274
rect 1898 1261 2008 1274
rect 1972 1205 2003 1206
rect 1820 1175 1829 1195
rect 1849 1175 1857 1195
rect 1374 1143 1381 1170
rect 1400 1169 1437 1170
rect 1496 1169 1533 1170
rect 1345 1118 1381 1143
rect 816 1116 857 1117
rect 652 1109 857 1116
rect 652 1098 826 1109
rect 652 1065 660 1098
rect 653 1056 660 1065
rect 709 1089 826 1098
rect 846 1089 857 1109
rect 709 1081 857 1089
rect 924 1113 1283 1117
rect 924 1108 1246 1113
rect 924 1084 1037 1108
rect 1061 1089 1246 1108
rect 1270 1089 1283 1113
rect 1061 1084 1283 1089
rect 924 1081 1283 1084
rect 1345 1081 1380 1118
rect 1448 1115 1548 1118
rect 1448 1111 1515 1115
rect 1448 1085 1460 1111
rect 1486 1089 1515 1111
rect 1541 1089 1548 1115
rect 1486 1085 1548 1089
rect 1448 1081 1548 1085
rect 709 1065 720 1081
rect 709 1056 717 1065
rect 924 1060 955 1081
rect 1345 1060 1381 1081
rect 767 1059 804 1060
rect 432 1016 497 1035
rect 432 998 457 1016
rect 475 998 497 1016
rect 432 797 497 998
rect 653 872 717 1056
rect 766 1050 804 1059
rect 766 1030 775 1050
rect 795 1030 804 1050
rect 766 1022 804 1030
rect 870 1054 955 1060
rect 980 1059 1017 1060
rect 870 1034 878 1054
rect 898 1034 955 1054
rect 870 1026 955 1034
rect 979 1050 1017 1059
rect 979 1030 988 1050
rect 1008 1030 1017 1050
rect 870 1025 906 1026
rect 979 1022 1017 1030
rect 1083 1054 1168 1060
rect 1188 1059 1225 1060
rect 1083 1034 1091 1054
rect 1111 1053 1168 1054
rect 1111 1034 1140 1053
rect 1083 1033 1140 1034
rect 1161 1033 1168 1053
rect 1083 1026 1168 1033
rect 1187 1050 1225 1059
rect 1187 1030 1196 1050
rect 1216 1030 1225 1050
rect 1083 1025 1119 1026
rect 1187 1022 1225 1030
rect 1291 1054 1435 1060
rect 1291 1034 1299 1054
rect 1319 1034 1407 1054
rect 1427 1034 1435 1054
rect 1291 1026 1435 1034
rect 1291 1025 1327 1026
rect 1399 1025 1435 1026
rect 1501 1059 1538 1060
rect 1501 1058 1539 1059
rect 1501 1050 1565 1058
rect 1501 1030 1510 1050
rect 1530 1036 1565 1050
rect 1585 1036 1588 1056
rect 1530 1031 1588 1036
rect 1530 1030 1565 1031
rect 767 993 804 1022
rect 768 991 804 993
rect 980 991 1017 1022
rect 768 969 1017 991
rect 849 963 960 969
rect 849 955 890 963
rect 849 935 857 955
rect 876 935 890 955
rect 849 933 890 935
rect 918 955 960 963
rect 918 935 934 955
rect 953 935 960 955
rect 918 933 960 935
rect 849 918 960 933
rect 653 862 721 872
rect 653 829 670 862
rect 710 829 721 862
rect 653 817 721 829
rect 653 815 717 817
rect 1188 798 1225 1022
rect 1501 1018 1565 1030
rect 1605 800 1632 1170
rect 1820 1165 1857 1175
rect 1916 1195 2003 1205
rect 1916 1175 1925 1195
rect 1945 1175 2003 1195
rect 1916 1166 2003 1175
rect 1916 1165 1953 1166
rect 1696 1152 1766 1157
rect 1691 1146 1766 1152
rect 1691 1113 1699 1146
rect 1752 1113 1766 1146
rect 1972 1113 2003 1166
rect 2033 1195 2070 1274
rect 2185 1205 2216 1206
rect 2033 1175 2042 1195
rect 2062 1175 2070 1195
rect 2033 1165 2070 1175
rect 2129 1198 2216 1205
rect 2129 1195 2190 1198
rect 2129 1175 2138 1195
rect 2158 1178 2190 1195
rect 2211 1178 2216 1198
rect 2158 1175 2216 1178
rect 2129 1168 2216 1175
rect 2241 1195 2278 1337
rect 2544 1336 2581 1337
rect 2393 1205 2429 1206
rect 2241 1175 2250 1195
rect 2270 1175 2278 1195
rect 2129 1166 2185 1168
rect 2129 1165 2166 1166
rect 2241 1165 2278 1175
rect 2337 1195 2485 1205
rect 2585 1202 2681 1204
rect 2337 1175 2346 1195
rect 2366 1175 2456 1195
rect 2476 1175 2485 1195
rect 2337 1169 2485 1175
rect 2337 1166 2401 1169
rect 2337 1165 2374 1166
rect 2393 1139 2401 1166
rect 2422 1166 2485 1169
rect 2543 1195 2681 1202
rect 2543 1175 2552 1195
rect 2572 1175 2681 1195
rect 2543 1166 2681 1175
rect 2422 1139 2429 1166
rect 2448 1165 2485 1166
rect 2544 1165 2581 1166
rect 2393 1114 2429 1139
rect 1691 1112 1774 1113
rect 1864 1112 1905 1113
rect 1691 1105 1905 1112
rect 1691 1088 1874 1105
rect 1691 1055 1704 1088
rect 1757 1085 1874 1088
rect 1894 1085 1905 1105
rect 1757 1077 1905 1085
rect 1972 1109 2331 1113
rect 1972 1104 2294 1109
rect 1972 1080 2085 1104
rect 2109 1085 2294 1104
rect 2318 1085 2331 1109
rect 2109 1080 2331 1085
rect 1972 1077 2331 1080
rect 2393 1077 2428 1114
rect 2496 1111 2596 1114
rect 2496 1107 2563 1111
rect 2496 1081 2508 1107
rect 2534 1085 2563 1107
rect 2589 1085 2596 1111
rect 2534 1081 2596 1085
rect 2496 1077 2596 1081
rect 1757 1055 1774 1077
rect 1972 1056 2003 1077
rect 2393 1056 2429 1077
rect 1815 1055 1852 1056
rect 1691 1041 1774 1055
rect 1464 798 1632 800
rect 1188 797 1632 798
rect 432 767 1632 797
rect 1702 831 1774 1041
rect 1814 1046 1852 1055
rect 1814 1026 1823 1046
rect 1843 1026 1852 1046
rect 1814 1018 1852 1026
rect 1918 1050 2003 1056
rect 2028 1055 2065 1056
rect 1918 1030 1926 1050
rect 1946 1030 2003 1050
rect 1918 1022 2003 1030
rect 2027 1046 2065 1055
rect 2027 1026 2036 1046
rect 2056 1026 2065 1046
rect 1918 1021 1954 1022
rect 2027 1018 2065 1026
rect 2131 1050 2216 1056
rect 2236 1055 2273 1056
rect 2131 1030 2139 1050
rect 2159 1049 2216 1050
rect 2159 1030 2188 1049
rect 2131 1029 2188 1030
rect 2209 1029 2216 1049
rect 2131 1022 2216 1029
rect 2235 1046 2273 1055
rect 2235 1026 2244 1046
rect 2264 1026 2273 1046
rect 2131 1021 2167 1022
rect 2235 1018 2273 1026
rect 2339 1050 2483 1056
rect 2339 1030 2347 1050
rect 2367 1030 2455 1050
rect 2475 1030 2483 1050
rect 2339 1022 2483 1030
rect 2339 1021 2375 1022
rect 2447 1021 2483 1022
rect 2549 1055 2586 1056
rect 2549 1054 2587 1055
rect 2549 1046 2613 1054
rect 2549 1026 2558 1046
rect 2578 1032 2613 1046
rect 2633 1032 2636 1052
rect 2578 1027 2636 1032
rect 2578 1026 2613 1027
rect 1815 989 1852 1018
rect 1816 987 1852 989
rect 2028 987 2065 1018
rect 1816 965 2065 987
rect 1897 959 2008 965
rect 1897 951 1938 959
rect 1897 931 1905 951
rect 1924 931 1938 951
rect 1897 929 1938 931
rect 1966 951 2008 959
rect 1966 931 1982 951
rect 2001 931 2008 951
rect 1966 929 2008 931
rect 1897 914 2008 929
rect 1702 792 1721 831
rect 1766 792 1774 831
rect 1702 775 1774 792
rect 2236 819 2273 1018
rect 2549 1014 2613 1026
rect 2236 813 2277 819
rect 2653 815 2680 1166
rect 2512 813 2680 815
rect 2236 787 2680 813
rect 432 720 497 767
rect 432 702 455 720
rect 473 702 497 720
rect 1345 747 1380 749
rect 1345 745 1449 747
rect 2238 745 2277 787
rect 2512 786 2680 787
rect 1345 738 2279 745
rect 1345 737 1396 738
rect 1345 717 1348 737
rect 1373 718 1396 737
rect 1428 718 2279 738
rect 1373 717 2279 718
rect 1345 710 2279 717
rect 1618 709 2279 710
rect 432 681 497 702
rect 709 692 749 695
rect 709 688 1612 692
rect 709 668 1586 688
rect 1606 668 1612 688
rect 709 665 1612 668
rect 433 621 498 641
rect 433 603 457 621
rect 475 603 498 621
rect 433 576 498 603
rect 709 576 749 665
rect 1193 663 1609 665
rect 1193 662 1534 663
rect 850 631 960 645
rect 850 628 893 631
rect 850 623 854 628
rect 432 541 749 576
rect 772 601 854 623
rect 883 601 893 628
rect 921 604 928 631
rect 957 623 960 631
rect 957 604 1022 623
rect 921 601 1022 604
rect 772 599 1022 601
rect 433 465 498 541
rect 772 520 809 599
rect 850 586 960 599
rect 924 530 955 531
rect 772 500 781 520
rect 801 500 809 520
rect 772 490 809 500
rect 868 520 955 530
rect 868 500 877 520
rect 897 500 955 520
rect 868 491 955 500
rect 868 490 905 491
rect 433 447 455 465
rect 473 447 498 465
rect 433 426 498 447
rect 646 445 711 454
rect 646 408 656 445
rect 696 437 711 445
rect 924 438 955 491
rect 985 520 1022 599
rect 1137 530 1168 531
rect 985 500 994 520
rect 1014 500 1022 520
rect 985 490 1022 500
rect 1081 523 1168 530
rect 1081 520 1142 523
rect 1081 500 1090 520
rect 1110 503 1142 520
rect 1163 503 1168 523
rect 1110 500 1168 503
rect 1081 493 1168 500
rect 1193 520 1230 662
rect 1496 661 1533 662
rect 1345 530 1381 531
rect 1193 500 1202 520
rect 1222 500 1230 520
rect 1081 491 1137 493
rect 1081 490 1118 491
rect 1193 490 1230 500
rect 1289 520 1437 530
rect 1537 527 1633 529
rect 1289 500 1298 520
rect 1318 500 1408 520
rect 1428 500 1437 520
rect 1289 494 1437 500
rect 1289 491 1353 494
rect 1289 490 1326 491
rect 1345 464 1353 491
rect 1374 491 1437 494
rect 1495 520 1633 527
rect 1495 500 1504 520
rect 1524 500 1633 520
rect 1495 491 1633 500
rect 1374 464 1381 491
rect 1400 490 1437 491
rect 1496 490 1533 491
rect 1345 439 1381 464
rect 816 437 857 438
rect 696 430 857 437
rect 696 410 826 430
rect 846 410 857 430
rect 696 408 857 410
rect 646 402 857 408
rect 924 434 1283 438
rect 924 429 1246 434
rect 924 405 1037 429
rect 1061 410 1246 429
rect 1270 410 1283 434
rect 1061 405 1283 410
rect 924 402 1283 405
rect 1345 402 1380 439
rect 1448 436 1548 439
rect 1448 432 1515 436
rect 1448 406 1460 432
rect 1486 410 1515 432
rect 1541 410 1548 436
rect 1486 406 1548 410
rect 1448 402 1548 406
rect 646 389 713 402
rect 438 366 494 386
rect 438 348 457 366
rect 475 348 494 366
rect 438 235 494 348
rect 646 368 660 389
rect 696 368 713 389
rect 924 381 955 402
rect 1345 381 1381 402
rect 767 380 804 381
rect 646 361 713 368
rect 766 371 804 380
rect 438 94 493 235
rect 646 209 711 361
rect 766 351 775 371
rect 795 351 804 371
rect 766 343 804 351
rect 870 375 955 381
rect 980 380 1017 381
rect 870 355 878 375
rect 898 355 955 375
rect 870 347 955 355
rect 979 371 1017 380
rect 979 351 988 371
rect 1008 351 1017 371
rect 870 346 906 347
rect 979 343 1017 351
rect 1083 375 1168 381
rect 1188 380 1225 381
rect 1083 355 1091 375
rect 1111 374 1168 375
rect 1111 355 1140 374
rect 1083 354 1140 355
rect 1161 354 1168 374
rect 1083 347 1168 354
rect 1187 371 1225 380
rect 1187 351 1196 371
rect 1216 351 1225 371
rect 1083 346 1119 347
rect 1187 343 1225 351
rect 1291 375 1435 381
rect 1291 355 1299 375
rect 1319 355 1407 375
rect 1427 355 1435 375
rect 1291 347 1435 355
rect 1291 346 1327 347
rect 1399 346 1435 347
rect 1501 380 1538 381
rect 1501 379 1539 380
rect 1501 371 1565 379
rect 1501 351 1510 371
rect 1530 357 1565 371
rect 1585 357 1588 377
rect 1530 352 1588 357
rect 1530 351 1565 352
rect 767 314 804 343
rect 768 312 804 314
rect 980 312 1017 343
rect 768 290 1017 312
rect 849 284 960 290
rect 849 276 890 284
rect 849 256 857 276
rect 876 256 890 276
rect 849 254 890 256
rect 918 276 960 284
rect 918 256 934 276
rect 953 256 960 276
rect 918 254 960 256
rect 849 239 960 254
rect 1188 244 1225 343
rect 1501 339 1565 351
rect 639 199 760 209
rect 639 197 708 199
rect 639 156 652 197
rect 689 158 708 197
rect 745 158 760 199
rect 689 156 760 158
rect 639 138 760 156
rect 851 94 955 239
rect 1186 94 1227 244
rect 1605 236 1632 491
rect 1694 481 1774 492
rect 1694 455 1711 481
rect 1751 455 1774 481
rect 1694 428 1774 455
rect 1694 402 1715 428
rect 1755 402 1774 428
rect 1694 383 1774 402
rect 1694 357 1718 383
rect 1758 357 1774 383
rect 1694 306 1774 357
rect 438 91 1227 94
rect 1606 105 1632 236
rect 1606 91 1634 105
rect 438 58 1634 91
rect 440 56 1634 58
rect 851 54 955 56
rect 1186 54 1227 56
rect 1696 53 1766 306
<< viali >>
rect 2822 5918 2859 5966
rect 1352 5820 1377 5855
rect 1396 5820 1421 5858
rect 1585 5761 1605 5781
rect 2402 5821 2427 5856
rect 2446 5821 2471 5859
rect 2633 5757 2653 5777
rect 853 5694 882 5721
rect 927 5697 956 5724
rect 658 5533 707 5575
rect 1141 5596 1162 5616
rect 1901 5690 1930 5717
rect 1975 5693 2004 5720
rect 1352 5557 1373 5587
rect 659 5470 708 5512
rect 1514 5503 1540 5529
rect 1139 5447 1160 5467
rect 1564 5450 1584 5470
rect 856 5349 875 5369
rect 933 5349 952 5369
rect 669 5243 709 5276
rect 1698 5527 1751 5560
rect 2189 5592 2210 5612
rect 2400 5553 2421 5583
rect 1703 5469 1756 5502
rect 2562 5499 2588 5525
rect 2187 5443 2208 5463
rect 2612 5446 2632 5466
rect 1904 5345 1923 5365
rect 1981 5345 2000 5365
rect 1720 5206 1765 5245
rect 2823 5506 2857 5545
rect 1347 5131 1372 5151
rect 1395 5132 1427 5152
rect 1585 5082 1605 5102
rect 853 5015 882 5042
rect 927 5018 956 5045
rect 655 4822 695 4859
rect 1141 4917 1162 4937
rect 3000 5526 3036 5567
rect 2989 5186 3049 5230
rect 4080 5077 4100 5097
rect 3348 5010 3377 5037
rect 3422 5013 3451 5040
rect 1352 4878 1373 4908
rect 1514 4824 1540 4850
rect 659 4782 695 4803
rect 1139 4768 1160 4788
rect 1564 4771 1584 4791
rect 856 4670 875 4690
rect 933 4670 952 4690
rect 651 4570 688 4611
rect 707 4572 744 4613
rect 1710 4869 1750 4895
rect 1714 4816 1754 4842
rect 1717 4771 1757 4797
rect 3636 4912 3657 4932
rect 3847 4873 3868 4903
rect 2989 4772 3043 4813
rect 4009 4819 4035 4845
rect 3634 4763 3655 4783
rect 1716 4446 1746 4512
rect 1352 4373 1377 4408
rect 1396 4373 1421 4411
rect 1585 4314 1605 4334
rect 2633 4310 2653 4330
rect 853 4247 882 4274
rect 927 4250 956 4277
rect 658 4086 707 4128
rect 1141 4149 1162 4169
rect 1901 4243 1930 4270
rect 1975 4246 2004 4273
rect 1352 4110 1373 4140
rect 659 4023 708 4065
rect 1514 4056 1540 4082
rect 1139 4000 1160 4020
rect 1564 4003 1584 4023
rect 856 3902 875 3922
rect 933 3902 952 3922
rect 669 3796 709 3829
rect 1698 4080 1751 4113
rect 2189 4145 2210 4165
rect 2400 4106 2421 4136
rect 1703 4022 1756 4055
rect 2562 4052 2588 4078
rect 2187 3996 2208 4016
rect 2612 3999 2632 4019
rect 1904 3898 1923 3918
rect 1981 3898 2000 3918
rect 1720 3759 1765 3798
rect 3351 4665 3370 4685
rect 3428 4665 3447 4685
rect 4059 4766 4079 4786
rect 3858 4575 3910 4593
rect 3627 4374 3652 4409
rect 3671 4374 3696 4412
rect 3890 4390 3914 4413
rect 3890 4346 3914 4369
rect 1347 3684 1372 3704
rect 1395 3685 1427 3705
rect 1585 3635 1605 3655
rect 853 3568 882 3595
rect 927 3571 956 3598
rect 655 3375 695 3412
rect 1141 3470 1162 3490
rect 1352 3431 1373 3461
rect 1514 3377 1540 3403
rect 659 3335 695 3356
rect 1139 3321 1160 3341
rect 1564 3324 1584 3344
rect 856 3223 875 3243
rect 933 3223 952 3243
rect 651 3123 688 3164
rect 707 3125 744 3166
rect 1710 3422 1750 3448
rect 1714 3369 1754 3395
rect 1717 3324 1757 3350
rect 1709 3064 1753 3101
rect 4123 3632 4143 3652
rect 3391 3565 3420 3592
rect 3465 3568 3494 3595
rect 3679 3467 3700 3487
rect 3890 3428 3911 3458
rect 4052 3374 4078 3400
rect 3677 3318 3698 3338
rect 4102 3321 4122 3341
rect 3394 3220 3413 3240
rect 3471 3220 3490 3240
rect 1704 2978 1758 3044
rect 1353 2853 1378 2888
rect 1397 2853 1422 2891
rect 1586 2794 1606 2814
rect 2634 2790 2654 2810
rect 854 2727 883 2754
rect 928 2730 957 2757
rect 659 2566 708 2608
rect 1142 2629 1163 2649
rect 1902 2723 1931 2750
rect 1976 2726 2005 2753
rect 1353 2590 1374 2620
rect 660 2503 709 2545
rect 1515 2536 1541 2562
rect 1140 2480 1161 2500
rect 1565 2483 1585 2503
rect 857 2382 876 2402
rect 934 2382 953 2402
rect 670 2276 710 2309
rect 1699 2560 1752 2593
rect 2190 2625 2211 2645
rect 2401 2586 2422 2616
rect 1704 2502 1757 2535
rect 2563 2532 2589 2558
rect 2188 2476 2209 2496
rect 2613 2479 2633 2499
rect 1905 2378 1924 2398
rect 1982 2378 2001 2398
rect 1721 2239 1766 2278
rect 3694 2854 3719 2892
rect 1348 2164 1373 2184
rect 1396 2165 1428 2185
rect 1586 2115 1606 2135
rect 854 2048 883 2075
rect 928 2051 957 2078
rect 656 1855 696 1892
rect 1142 1950 1163 1970
rect 1353 1911 1374 1941
rect 1515 1857 1541 1883
rect 660 1815 696 1836
rect 1140 1801 1161 1821
rect 1565 1804 1585 1824
rect 857 1703 876 1723
rect 934 1703 953 1723
rect 652 1603 689 1644
rect 708 1605 745 1646
rect 3852 2163 3869 2200
rect 4081 2110 4101 2130
rect 3349 2043 3378 2070
rect 3423 2046 3452 2073
rect 1711 1902 1751 1928
rect 1715 1849 1755 1875
rect 1718 1804 1758 1830
rect 3637 1945 3658 1965
rect 3848 1906 3869 1936
rect 2825 1845 2851 1868
rect 3205 1838 3231 1861
rect 4010 1852 4036 1878
rect 3635 1796 3656 1816
rect 4060 1799 4080 1819
rect 3352 1698 3371 1718
rect 3429 1698 3448 1718
rect 1717 1479 1747 1545
rect 1353 1406 1378 1441
rect 1397 1406 1422 1444
rect 3692 1426 3720 1454
rect 1586 1347 1606 1367
rect 2634 1343 2654 1363
rect 854 1280 883 1307
rect 928 1283 957 1310
rect 659 1119 708 1161
rect 1142 1182 1163 1202
rect 1902 1276 1931 1303
rect 1976 1279 2005 1306
rect 1353 1143 1374 1173
rect 660 1056 709 1098
rect 1515 1089 1541 1115
rect 1140 1033 1161 1053
rect 1565 1036 1585 1056
rect 857 935 876 955
rect 934 935 953 955
rect 670 829 710 862
rect 1699 1113 1752 1146
rect 2190 1178 2211 1198
rect 2401 1139 2422 1169
rect 1704 1055 1757 1088
rect 2563 1085 2589 1111
rect 2188 1029 2209 1049
rect 2613 1032 2633 1052
rect 1905 931 1924 951
rect 1982 931 2001 951
rect 1721 792 1766 831
rect 1348 717 1373 737
rect 1396 718 1428 738
rect 1586 668 1606 688
rect 854 601 883 628
rect 928 604 957 631
rect 656 408 696 445
rect 1142 503 1163 523
rect 1353 464 1374 494
rect 1515 410 1541 436
rect 660 368 696 389
rect 1140 354 1161 374
rect 1565 357 1585 377
rect 857 256 876 276
rect 934 256 953 276
rect 652 156 689 197
rect 708 158 745 199
rect 1711 455 1751 481
rect 1715 402 1755 428
rect 1718 357 1758 383
<< metal1 >>
rect 170 5387 277 5984
rect 649 5575 721 5975
rect 1345 5866 1417 5867
rect 1344 5858 1443 5866
rect 1344 5855 1396 5858
rect 1344 5820 1352 5855
rect 1377 5820 1396 5855
rect 1421 5820 1443 5858
rect 1344 5808 1443 5820
rect 1345 5789 1413 5808
rect 1346 5786 1379 5789
rect 1581 5786 1613 5787
rect 756 5725 959 5738
rect 756 5692 780 5725
rect 816 5724 959 5725
rect 816 5721 927 5724
rect 816 5694 853 5721
rect 882 5697 927 5721
rect 956 5697 959 5724
rect 882 5694 959 5697
rect 816 5692 959 5694
rect 756 5679 959 5692
rect 756 5678 857 5679
rect 649 5533 658 5575
rect 707 5533 721 5575
rect 649 5512 721 5533
rect 649 5470 659 5512
rect 708 5470 721 5512
rect 649 5452 721 5470
rect 1134 5616 1166 5623
rect 1134 5596 1141 5616
rect 1162 5596 1166 5616
rect 1134 5531 1166 5596
rect 1346 5587 1377 5786
rect 1578 5781 1613 5786
rect 1578 5761 1585 5781
rect 1605 5761 1613 5781
rect 1578 5753 1613 5761
rect 1346 5557 1352 5587
rect 1373 5557 1377 5587
rect 1346 5549 1377 5557
rect 1504 5531 1544 5532
rect 1134 5529 1546 5531
rect 1134 5503 1514 5529
rect 1540 5503 1546 5529
rect 1134 5495 1546 5503
rect 1134 5467 1166 5495
rect 1579 5475 1613 5753
rect 1695 5566 1765 5976
rect 2809 5966 2874 6001
rect 2809 5962 2822 5966
rect 2810 5918 2822 5962
rect 2859 5962 2874 5966
rect 2859 5918 2872 5962
rect 2395 5867 2467 5868
rect 2394 5859 2483 5867
rect 2394 5856 2446 5859
rect 2394 5821 2402 5856
rect 2427 5821 2446 5856
rect 2471 5821 2483 5859
rect 2394 5809 2483 5821
rect 2394 5808 2463 5809
rect 2394 5790 2430 5808
rect 1804 5721 2007 5734
rect 1804 5688 1828 5721
rect 1864 5720 2007 5721
rect 1864 5717 1975 5720
rect 1864 5690 1901 5717
rect 1930 5693 1975 5717
rect 2004 5693 2007 5720
rect 1930 5690 2007 5693
rect 1864 5688 2007 5690
rect 1804 5675 2007 5688
rect 1804 5674 1905 5675
rect 1134 5447 1139 5467
rect 1160 5447 1166 5467
rect 1134 5440 1166 5447
rect 1557 5470 1613 5475
rect 1557 5450 1564 5470
rect 1584 5450 1613 5470
rect 1690 5560 1765 5566
rect 1690 5527 1698 5560
rect 1751 5527 1765 5560
rect 1690 5502 1765 5527
rect 1690 5469 1703 5502
rect 1756 5469 1765 5502
rect 1690 5460 1765 5469
rect 2182 5612 2214 5619
rect 2182 5592 2189 5612
rect 2210 5592 2214 5612
rect 2182 5527 2214 5592
rect 2394 5583 2425 5790
rect 2629 5782 2661 5783
rect 2626 5777 2661 5782
rect 2626 5757 2633 5777
rect 2653 5757 2661 5777
rect 2626 5749 2661 5757
rect 2394 5553 2400 5583
rect 2421 5553 2425 5583
rect 2394 5545 2425 5553
rect 2552 5527 2592 5528
rect 2182 5525 2594 5527
rect 2182 5499 2562 5525
rect 2588 5499 2594 5525
rect 2182 5491 2594 5499
rect 2182 5463 2214 5491
rect 2627 5471 2661 5749
rect 2810 5564 2872 5918
rect 2979 5567 3061 5996
rect 2810 5545 2874 5564
rect 2810 5506 2823 5545
rect 2857 5506 2874 5545
rect 2810 5487 2874 5506
rect 2979 5526 3000 5567
rect 3036 5526 3061 5567
rect 2979 5497 3061 5526
rect 1690 5455 1748 5460
rect 1557 5443 1613 5450
rect 2182 5443 2187 5463
rect 2208 5443 2214 5463
rect 1557 5442 1592 5443
rect 2182 5436 2214 5443
rect 2605 5466 2661 5471
rect 2605 5446 2612 5466
rect 2632 5446 2661 5466
rect 2605 5439 2661 5446
rect 2605 5438 2640 5439
rect 848 5387 959 5391
rect 2631 5387 4201 5388
rect 170 5369 4201 5387
rect 170 5349 856 5369
rect 875 5349 933 5369
rect 952 5365 4201 5369
rect 952 5349 1904 5365
rect 170 5345 1904 5349
rect 1923 5345 1981 5365
rect 2000 5345 4201 5365
rect 170 5331 4201 5345
rect 170 4708 277 5331
rect 1896 5328 2007 5331
rect 656 5282 720 5286
rect 652 5276 720 5282
rect 652 5243 669 5276
rect 709 5243 720 5276
rect 652 5231 720 5243
rect 1703 5245 1768 5267
rect 652 5229 709 5231
rect 656 4868 707 5229
rect 1703 5206 1720 5245
rect 1765 5206 1768 5245
rect 1344 5161 1379 5163
rect 1344 5152 1448 5161
rect 1344 5151 1395 5152
rect 1344 5131 1347 5151
rect 1372 5132 1395 5151
rect 1427 5132 1448 5152
rect 1372 5131 1448 5132
rect 1344 5124 1448 5131
rect 1344 5112 1379 5124
rect 756 5046 959 5059
rect 756 5013 780 5046
rect 816 5045 959 5046
rect 816 5042 927 5045
rect 816 5015 853 5042
rect 882 5018 927 5042
rect 956 5018 959 5045
rect 882 5015 959 5018
rect 816 5013 959 5015
rect 756 5000 959 5013
rect 756 4999 857 5000
rect 1134 4937 1166 4944
rect 1134 4917 1141 4937
rect 1162 4917 1166 4937
rect 645 4859 710 4868
rect 645 4822 655 4859
rect 695 4825 710 4859
rect 1134 4852 1166 4917
rect 1346 4908 1377 5112
rect 1581 5107 1613 5108
rect 1578 5102 1613 5107
rect 1578 5082 1585 5102
rect 1605 5082 1613 5102
rect 1578 5074 1613 5082
rect 1346 4878 1352 4908
rect 1373 4878 1377 4908
rect 1346 4870 1377 4878
rect 1504 4852 1544 4853
rect 1134 4850 1546 4852
rect 695 4822 712 4825
rect 645 4803 712 4822
rect 645 4782 659 4803
rect 695 4782 712 4803
rect 645 4775 712 4782
rect 1134 4824 1514 4850
rect 1540 4824 1546 4850
rect 1134 4816 1546 4824
rect 1134 4788 1166 4816
rect 1579 4796 1613 5074
rect 1703 4906 1768 5206
rect 2974 5230 3067 5245
rect 2974 5186 2989 5230
rect 3049 5186 3067 5230
rect 1134 4768 1139 4788
rect 1160 4768 1166 4788
rect 1134 4761 1166 4768
rect 1557 4791 1613 4796
rect 1557 4771 1564 4791
rect 1584 4771 1613 4791
rect 1557 4764 1613 4771
rect 1693 4895 1773 4906
rect 1693 4869 1710 4895
rect 1750 4869 1773 4895
rect 1693 4842 1773 4869
rect 1693 4816 1714 4842
rect 1754 4816 1773 4842
rect 1693 4797 1773 4816
rect 1693 4771 1717 4797
rect 1757 4771 1773 4797
rect 1557 4763 1592 4764
rect 1693 4759 1773 4771
rect 2974 4813 3067 5186
rect 3251 5041 3454 5054
rect 3251 5008 3275 5041
rect 3311 5040 3454 5041
rect 3311 5037 3422 5040
rect 3311 5010 3348 5037
rect 3377 5013 3422 5037
rect 3451 5013 3454 5040
rect 3377 5010 3454 5013
rect 3311 5008 3454 5010
rect 3251 4995 3454 5008
rect 3251 4994 3352 4995
rect 2974 4772 2989 4813
rect 3043 4772 3067 4813
rect 2974 4765 3067 4772
rect 3629 4932 3661 4939
rect 3629 4912 3636 4932
rect 3657 4912 3661 4932
rect 3629 4847 3661 4912
rect 3841 4903 3872 5104
rect 4076 5102 4108 5103
rect 4073 5097 4108 5102
rect 4073 5077 4080 5097
rect 4100 5077 4108 5097
rect 4073 5069 4108 5077
rect 3841 4873 3847 4903
rect 3868 4873 3872 4903
rect 3841 4865 3872 4873
rect 3999 4847 4039 4848
rect 3629 4845 4041 4847
rect 3629 4819 4009 4845
rect 4035 4819 4041 4845
rect 3629 4811 4041 4819
rect 3629 4783 3661 4811
rect 4074 4791 4108 5069
rect 3629 4763 3634 4783
rect 3655 4763 3661 4783
rect 3629 4756 3661 4763
rect 4052 4786 4108 4791
rect 4052 4766 4059 4786
rect 4079 4766 4108 4786
rect 4052 4759 4108 4766
rect 4052 4758 4087 4759
rect 848 4708 959 4712
rect 2590 4708 4234 4711
rect 168 4690 4234 4708
rect 168 4670 856 4690
rect 875 4670 933 4690
rect 952 4685 4234 4690
rect 952 4670 3351 4685
rect 168 4665 3351 4670
rect 3370 4665 3428 4685
rect 3447 4665 4234 4685
rect 168 4655 4234 4665
rect 168 4652 793 4655
rect 980 4652 4234 4655
rect 170 4424 277 4652
rect 2590 4651 4234 4652
rect 3343 4648 3454 4651
rect 638 4613 759 4623
rect 638 4611 707 4613
rect 638 4570 651 4611
rect 688 4572 707 4611
rect 744 4572 759 4613
rect 688 4570 759 4572
rect 638 4552 759 4570
rect 3843 4593 3929 4597
rect 3843 4575 3858 4593
rect 3910 4575 3929 4593
rect 3843 4566 3929 4575
rect 644 4450 723 4552
rect 1696 4512 1763 4531
rect 1696 4492 1716 4512
rect 170 4369 278 4424
rect 645 4369 723 4450
rect 1695 4446 1716 4492
rect 1746 4492 1763 4512
rect 1746 4462 1765 4492
rect 1746 4446 1766 4462
rect 1695 4430 1766 4446
rect 1345 4419 1417 4420
rect 1344 4411 1443 4419
rect 1344 4408 1396 4411
rect 1344 4373 1352 4408
rect 1377 4373 1396 4408
rect 1421 4373 1443 4411
rect 170 3940 277 4369
rect 649 4128 721 4369
rect 1344 4361 1443 4373
rect 1345 4342 1413 4361
rect 1346 4339 1379 4342
rect 1581 4339 1613 4340
rect 756 4278 959 4291
rect 756 4245 780 4278
rect 816 4277 959 4278
rect 816 4274 927 4277
rect 816 4247 853 4274
rect 882 4250 927 4274
rect 956 4250 959 4277
rect 882 4247 959 4250
rect 816 4245 959 4247
rect 756 4232 959 4245
rect 756 4231 857 4232
rect 649 4086 658 4128
rect 707 4086 721 4128
rect 649 4065 721 4086
rect 649 4023 659 4065
rect 708 4023 721 4065
rect 649 4005 721 4023
rect 1134 4169 1166 4176
rect 1134 4149 1141 4169
rect 1162 4149 1166 4169
rect 1134 4084 1166 4149
rect 1346 4140 1377 4339
rect 1578 4334 1613 4339
rect 1578 4314 1585 4334
rect 1605 4314 1613 4334
rect 1578 4306 1613 4314
rect 1346 4110 1352 4140
rect 1373 4110 1377 4140
rect 1346 4102 1377 4110
rect 1504 4084 1544 4085
rect 1134 4082 1546 4084
rect 1134 4056 1514 4082
rect 1540 4056 1546 4082
rect 1134 4048 1546 4056
rect 1134 4020 1166 4048
rect 1579 4028 1613 4306
rect 1695 4119 1765 4430
rect 3620 4420 3692 4421
rect 3619 4417 3708 4420
rect 2391 4415 3708 4417
rect 2388 4412 3708 4415
rect 2388 4409 3671 4412
rect 2388 4374 3627 4409
rect 3652 4374 3671 4409
rect 3696 4374 3708 4412
rect 2388 4364 3708 4374
rect 3884 4413 3920 4566
rect 3884 4390 3890 4413
rect 3914 4390 3920 4413
rect 3884 4369 3920 4390
rect 2388 4362 3673 4364
rect 2388 4352 2485 4362
rect 2394 4343 2430 4352
rect 3884 4346 3890 4369
rect 3914 4346 3920 4369
rect 1804 4274 2007 4287
rect 1804 4241 1828 4274
rect 1864 4273 2007 4274
rect 1864 4270 1975 4273
rect 1864 4243 1901 4270
rect 1930 4246 1975 4270
rect 2004 4246 2007 4273
rect 1930 4243 2007 4246
rect 1864 4241 2007 4243
rect 1804 4228 2007 4241
rect 1804 4227 1905 4228
rect 1134 4000 1139 4020
rect 1160 4000 1166 4020
rect 1134 3993 1166 4000
rect 1557 4023 1613 4028
rect 1557 4003 1564 4023
rect 1584 4003 1613 4023
rect 1690 4113 1765 4119
rect 1690 4080 1698 4113
rect 1751 4080 1765 4113
rect 1690 4055 1765 4080
rect 1690 4022 1703 4055
rect 1756 4022 1765 4055
rect 1690 4013 1765 4022
rect 2182 4165 2214 4172
rect 2182 4145 2189 4165
rect 2210 4145 2214 4165
rect 2182 4080 2214 4145
rect 2394 4136 2425 4343
rect 2629 4335 2661 4336
rect 3884 4335 3920 4346
rect 2626 4330 2661 4335
rect 2626 4310 2633 4330
rect 2653 4310 2661 4330
rect 2626 4302 2661 4310
rect 2394 4106 2400 4136
rect 2421 4106 2425 4136
rect 2394 4098 2425 4106
rect 2552 4080 2592 4081
rect 2182 4078 2594 4080
rect 2182 4052 2562 4078
rect 2588 4052 2594 4078
rect 2182 4044 2594 4052
rect 2182 4016 2214 4044
rect 2627 4024 2661 4302
rect 1690 4008 1748 4013
rect 1557 3996 1613 4003
rect 2182 3996 2187 4016
rect 2208 3996 2214 4016
rect 1557 3995 1592 3996
rect 2182 3989 2214 3996
rect 2605 4019 2661 4024
rect 2605 3999 2612 4019
rect 2632 3999 2661 4019
rect 2605 3992 2661 3999
rect 2605 3991 2640 3992
rect 848 3940 959 3944
rect 2723 3940 4234 3941
rect 170 3922 4234 3940
rect 170 3902 856 3922
rect 875 3902 933 3922
rect 952 3918 4234 3922
rect 952 3902 1904 3918
rect 170 3898 1904 3902
rect 1923 3898 1981 3918
rect 2000 3898 4234 3918
rect 170 3884 4234 3898
rect 170 3261 277 3884
rect 1896 3881 2007 3884
rect 656 3835 720 3839
rect 652 3829 720 3835
rect 652 3796 669 3829
rect 709 3796 720 3829
rect 652 3784 720 3796
rect 1703 3798 1768 3820
rect 652 3782 709 3784
rect 656 3421 707 3782
rect 1703 3759 1720 3798
rect 1765 3759 1768 3798
rect 1344 3714 1379 3716
rect 1344 3705 1448 3714
rect 1344 3704 1395 3705
rect 1344 3684 1347 3704
rect 1372 3685 1395 3704
rect 1427 3685 1448 3705
rect 1372 3684 1448 3685
rect 1344 3677 1448 3684
rect 1344 3665 1379 3677
rect 756 3599 959 3612
rect 756 3566 780 3599
rect 816 3598 959 3599
rect 816 3595 927 3598
rect 816 3568 853 3595
rect 882 3571 927 3595
rect 956 3571 959 3598
rect 882 3568 959 3571
rect 816 3566 959 3568
rect 756 3553 959 3566
rect 756 3552 857 3553
rect 1134 3490 1166 3497
rect 1134 3470 1141 3490
rect 1162 3470 1166 3490
rect 645 3412 710 3421
rect 645 3375 655 3412
rect 695 3378 710 3412
rect 1134 3405 1166 3470
rect 1346 3461 1377 3665
rect 1581 3660 1613 3661
rect 1578 3655 1613 3660
rect 1578 3635 1585 3655
rect 1605 3635 1613 3655
rect 1578 3627 1613 3635
rect 1346 3431 1352 3461
rect 1373 3431 1377 3461
rect 1346 3423 1377 3431
rect 1504 3405 1544 3406
rect 1134 3403 1546 3405
rect 695 3375 712 3378
rect 645 3356 712 3375
rect 645 3335 659 3356
rect 695 3335 712 3356
rect 645 3328 712 3335
rect 1134 3377 1514 3403
rect 1540 3377 1546 3403
rect 1134 3369 1546 3377
rect 1134 3341 1166 3369
rect 1579 3349 1613 3627
rect 1703 3459 1768 3759
rect 3294 3596 3497 3609
rect 3294 3563 3318 3596
rect 3354 3595 3497 3596
rect 3354 3592 3465 3595
rect 3354 3565 3391 3592
rect 3420 3568 3465 3592
rect 3494 3568 3497 3595
rect 3420 3565 3497 3568
rect 3354 3563 3497 3565
rect 3294 3550 3497 3563
rect 3294 3549 3395 3550
rect 3672 3487 3704 3494
rect 3672 3467 3679 3487
rect 3700 3467 3704 3487
rect 1134 3321 1139 3341
rect 1160 3321 1166 3341
rect 1134 3314 1166 3321
rect 1557 3344 1613 3349
rect 1557 3324 1564 3344
rect 1584 3324 1613 3344
rect 1557 3317 1613 3324
rect 1693 3448 1773 3459
rect 1693 3422 1710 3448
rect 1750 3422 1773 3448
rect 1693 3395 1773 3422
rect 1693 3369 1714 3395
rect 1754 3369 1773 3395
rect 1693 3350 1773 3369
rect 1693 3324 1717 3350
rect 1757 3324 1773 3350
rect 1557 3316 1592 3317
rect 1693 3312 1773 3324
rect 3672 3402 3704 3467
rect 3884 3458 3915 3728
rect 4119 3657 4151 3658
rect 4116 3652 4151 3657
rect 4116 3632 4123 3652
rect 4143 3632 4151 3652
rect 4116 3624 4151 3632
rect 3884 3428 3890 3458
rect 3911 3428 3915 3458
rect 3884 3420 3915 3428
rect 4042 3402 4082 3403
rect 3672 3400 4084 3402
rect 3672 3374 4052 3400
rect 4078 3374 4084 3400
rect 3672 3366 4084 3374
rect 3672 3338 3704 3366
rect 4117 3346 4151 3624
rect 3672 3318 3677 3338
rect 3698 3318 3704 3338
rect 3672 3311 3704 3318
rect 4095 3341 4151 3346
rect 4095 3321 4102 3341
rect 4122 3321 4151 3341
rect 4095 3314 4151 3321
rect 4095 3313 4130 3314
rect 848 3261 959 3265
rect 2603 3261 2810 3262
rect 3386 3261 3497 3262
rect 168 3243 4234 3261
rect 168 3223 856 3243
rect 875 3223 933 3243
rect 952 3240 4234 3243
rect 952 3223 3394 3240
rect 168 3220 3394 3223
rect 3413 3220 3471 3240
rect 3490 3220 4234 3240
rect 168 3205 4234 3220
rect 170 3017 277 3205
rect 2765 3203 4234 3205
rect 638 3166 759 3176
rect 638 3164 707 3166
rect 638 3123 651 3164
rect 688 3125 707 3164
rect 744 3125 759 3166
rect 688 3123 759 3125
rect 638 3105 759 3123
rect 170 3013 278 3017
rect 644 3013 721 3105
rect 1694 3101 1770 3117
rect 1694 3078 1709 3101
rect 171 2420 278 3013
rect 646 2962 721 3013
rect 1687 3064 1709 3078
rect 1753 3064 1770 3101
rect 1687 3044 1770 3064
rect 1687 2978 1704 3044
rect 1758 2978 1770 3044
rect 646 2919 722 2962
rect 650 2608 722 2919
rect 1687 2954 1770 2978
rect 1687 2934 1763 2954
rect 1687 2915 1766 2934
rect 1346 2899 1418 2900
rect 1345 2891 1444 2899
rect 1345 2888 1397 2891
rect 1345 2853 1353 2888
rect 1378 2853 1397 2888
rect 1422 2853 1444 2891
rect 1345 2841 1444 2853
rect 1346 2822 1414 2841
rect 1347 2819 1380 2822
rect 1582 2819 1614 2820
rect 757 2758 960 2771
rect 757 2725 781 2758
rect 817 2757 960 2758
rect 817 2754 928 2757
rect 817 2727 854 2754
rect 883 2730 928 2754
rect 957 2730 960 2757
rect 883 2727 960 2730
rect 817 2725 960 2727
rect 757 2712 960 2725
rect 757 2711 858 2712
rect 650 2566 659 2608
rect 708 2566 722 2608
rect 650 2545 722 2566
rect 650 2503 660 2545
rect 709 2503 722 2545
rect 650 2485 722 2503
rect 1135 2649 1167 2656
rect 1135 2629 1142 2649
rect 1163 2629 1167 2649
rect 1135 2564 1167 2629
rect 1347 2620 1378 2819
rect 1579 2814 1614 2819
rect 1579 2794 1586 2814
rect 1606 2794 1614 2814
rect 1579 2786 1614 2794
rect 1347 2590 1353 2620
rect 1374 2590 1378 2620
rect 1347 2582 1378 2590
rect 1505 2564 1545 2565
rect 1135 2562 1547 2564
rect 1135 2536 1515 2562
rect 1541 2536 1547 2562
rect 1135 2528 1547 2536
rect 1135 2500 1167 2528
rect 1580 2508 1614 2786
rect 1696 2599 1766 2915
rect 3684 2900 3715 2901
rect 3684 2892 3729 2900
rect 2764 2869 2928 2876
rect 3684 2869 3694 2892
rect 2390 2854 3694 2869
rect 3719 2854 3729 2892
rect 2390 2836 3729 2854
rect 2395 2823 2431 2836
rect 2764 2833 2928 2836
rect 1805 2754 2008 2767
rect 1805 2721 1829 2754
rect 1865 2753 2008 2754
rect 1865 2750 1976 2753
rect 1865 2723 1902 2750
rect 1931 2726 1976 2750
rect 2005 2726 2008 2753
rect 1931 2723 2008 2726
rect 1865 2721 2008 2723
rect 1805 2708 2008 2721
rect 1805 2707 1906 2708
rect 1135 2480 1140 2500
rect 1161 2480 1167 2500
rect 1135 2473 1167 2480
rect 1558 2503 1614 2508
rect 1558 2483 1565 2503
rect 1585 2483 1614 2503
rect 1691 2593 1766 2599
rect 1691 2560 1699 2593
rect 1752 2560 1766 2593
rect 1691 2535 1766 2560
rect 1691 2502 1704 2535
rect 1757 2502 1766 2535
rect 1691 2493 1766 2502
rect 2183 2645 2215 2652
rect 2183 2625 2190 2645
rect 2211 2625 2215 2645
rect 2183 2560 2215 2625
rect 2395 2616 2426 2823
rect 2630 2815 2662 2816
rect 2627 2810 2662 2815
rect 2627 2790 2634 2810
rect 2654 2790 2662 2810
rect 2627 2782 2662 2790
rect 2395 2586 2401 2616
rect 2422 2586 2426 2616
rect 2395 2578 2426 2586
rect 2553 2560 2593 2561
rect 2183 2558 2595 2560
rect 2183 2532 2563 2558
rect 2589 2532 2595 2558
rect 2183 2524 2595 2532
rect 2183 2496 2215 2524
rect 2628 2504 2662 2782
rect 1691 2488 1749 2493
rect 1558 2476 1614 2483
rect 2183 2476 2188 2496
rect 2209 2476 2215 2496
rect 1558 2475 1593 2476
rect 2183 2469 2215 2476
rect 2606 2499 2662 2504
rect 2606 2479 2613 2499
rect 2633 2479 2662 2499
rect 2606 2472 2662 2479
rect 2606 2471 2641 2472
rect 849 2420 960 2424
rect 2632 2420 4202 2421
rect 171 2402 4202 2420
rect 171 2382 857 2402
rect 876 2382 934 2402
rect 953 2398 4202 2402
rect 953 2382 1905 2398
rect 171 2378 1905 2382
rect 1924 2378 1982 2398
rect 2001 2378 4202 2398
rect 171 2364 4202 2378
rect 171 1741 278 2364
rect 1897 2361 2008 2364
rect 657 2315 721 2319
rect 653 2309 721 2315
rect 653 2276 670 2309
rect 710 2276 721 2309
rect 653 2264 721 2276
rect 1704 2278 1769 2300
rect 653 2262 710 2264
rect 657 1901 708 2262
rect 1704 2239 1721 2278
rect 1766 2239 1769 2278
rect 1345 2194 1380 2196
rect 1345 2185 1449 2194
rect 1345 2184 1396 2185
rect 1345 2164 1348 2184
rect 1373 2165 1396 2184
rect 1428 2165 1449 2185
rect 1373 2164 1449 2165
rect 1345 2157 1449 2164
rect 1345 2145 1380 2157
rect 757 2079 960 2092
rect 757 2046 781 2079
rect 817 2078 960 2079
rect 817 2075 928 2078
rect 817 2048 854 2075
rect 883 2051 928 2075
rect 957 2051 960 2078
rect 883 2048 960 2051
rect 817 2046 960 2048
rect 757 2033 960 2046
rect 757 2032 858 2033
rect 1135 1970 1167 1977
rect 1135 1950 1142 1970
rect 1163 1950 1167 1970
rect 646 1892 711 1901
rect 646 1855 656 1892
rect 696 1858 711 1892
rect 1135 1885 1167 1950
rect 1347 1941 1378 2145
rect 1582 2140 1614 2141
rect 1579 2135 1614 2140
rect 1579 2115 1586 2135
rect 1606 2115 1614 2135
rect 1579 2107 1614 2115
rect 1347 1911 1353 1941
rect 1374 1911 1378 1941
rect 1347 1903 1378 1911
rect 1505 1885 1545 1886
rect 1135 1883 1547 1885
rect 696 1855 713 1858
rect 646 1836 713 1855
rect 646 1815 660 1836
rect 696 1815 713 1836
rect 646 1808 713 1815
rect 1135 1857 1515 1883
rect 1541 1857 1547 1883
rect 1135 1849 1547 1857
rect 1135 1821 1167 1849
rect 1580 1829 1614 2107
rect 1704 1939 1769 2239
rect 3841 2200 3878 2221
rect 3841 2163 3852 2200
rect 3869 2176 3878 2200
rect 3869 2163 3879 2176
rect 3841 2153 3879 2163
rect 3842 2149 3879 2153
rect 3842 2143 3875 2149
rect 3252 2074 3455 2087
rect 3252 2041 3276 2074
rect 3312 2073 3455 2074
rect 3312 2070 3423 2073
rect 3312 2043 3349 2070
rect 3378 2046 3423 2070
rect 3452 2046 3455 2073
rect 3378 2043 3455 2046
rect 3312 2041 3455 2043
rect 3252 2028 3455 2041
rect 3252 2027 3353 2028
rect 3630 1965 3662 1972
rect 3630 1945 3637 1965
rect 3658 1945 3662 1965
rect 1135 1801 1140 1821
rect 1161 1801 1167 1821
rect 1135 1794 1167 1801
rect 1558 1824 1614 1829
rect 1558 1804 1565 1824
rect 1585 1804 1614 1824
rect 1558 1797 1614 1804
rect 1694 1928 1774 1939
rect 1694 1902 1711 1928
rect 1751 1902 1774 1928
rect 1694 1875 1774 1902
rect 1694 1849 1715 1875
rect 1755 1849 1774 1875
rect 3630 1880 3662 1945
rect 3842 1936 3873 2143
rect 4077 2135 4109 2136
rect 4074 2130 4109 2135
rect 4074 2110 4081 2130
rect 4101 2110 4109 2130
rect 4074 2102 4109 2110
rect 3842 1906 3848 1936
rect 3869 1906 3873 1936
rect 3842 1898 3873 1906
rect 4000 1880 4040 1881
rect 3630 1878 4042 1880
rect 1694 1830 1774 1849
rect 1694 1804 1718 1830
rect 1758 1804 1774 1830
rect 2807 1868 3244 1874
rect 2807 1845 2825 1868
rect 2851 1861 3244 1868
rect 2851 1845 3205 1861
rect 2807 1838 3205 1845
rect 3231 1838 3244 1861
rect 2807 1825 3244 1838
rect 3630 1852 4010 1878
rect 4036 1852 4042 1878
rect 3630 1844 4042 1852
rect 1558 1796 1593 1797
rect 1694 1792 1774 1804
rect 3630 1816 3662 1844
rect 4075 1824 4109 2102
rect 3630 1796 3635 1816
rect 3656 1796 3662 1816
rect 3630 1789 3662 1796
rect 4053 1819 4109 1824
rect 4053 1799 4060 1819
rect 4080 1799 4109 1819
rect 4053 1792 4109 1799
rect 4053 1791 4088 1792
rect 849 1741 960 1745
rect 2591 1741 4244 1744
rect 169 1723 4244 1741
rect 169 1703 857 1723
rect 876 1703 934 1723
rect 953 1718 4244 1723
rect 953 1703 3352 1718
rect 169 1698 3352 1703
rect 3371 1698 3429 1718
rect 3448 1698 4244 1718
rect 169 1688 4244 1698
rect 169 1685 794 1688
rect 981 1685 4244 1688
rect 171 1457 278 1685
rect 2591 1684 4244 1685
rect 3344 1681 3455 1684
rect 639 1646 760 1656
rect 639 1644 708 1646
rect 639 1603 652 1644
rect 689 1605 708 1644
rect 745 1605 760 1646
rect 689 1603 760 1605
rect 639 1585 760 1603
rect 645 1483 724 1585
rect 1697 1545 1764 1564
rect 1697 1525 1717 1545
rect 171 1402 279 1457
rect 646 1402 724 1483
rect 1696 1479 1717 1525
rect 1747 1525 1764 1545
rect 1747 1495 1766 1525
rect 1747 1479 1767 1495
rect 1696 1463 1767 1479
rect 1346 1452 1418 1453
rect 1345 1444 1444 1452
rect 1345 1441 1397 1444
rect 1345 1406 1353 1441
rect 1378 1406 1397 1441
rect 1422 1406 1444 1444
rect 171 973 278 1402
rect 650 1161 722 1402
rect 1345 1394 1444 1406
rect 1346 1375 1414 1394
rect 1347 1372 1380 1375
rect 1582 1372 1614 1373
rect 757 1311 960 1324
rect 757 1278 781 1311
rect 817 1310 960 1311
rect 817 1307 928 1310
rect 817 1280 854 1307
rect 883 1283 928 1307
rect 957 1283 960 1310
rect 883 1280 960 1283
rect 817 1278 960 1280
rect 757 1265 960 1278
rect 757 1264 858 1265
rect 650 1119 659 1161
rect 708 1119 722 1161
rect 650 1098 722 1119
rect 650 1056 660 1098
rect 709 1056 722 1098
rect 650 1038 722 1056
rect 1135 1202 1167 1209
rect 1135 1182 1142 1202
rect 1163 1182 1167 1202
rect 1135 1117 1167 1182
rect 1347 1173 1378 1372
rect 1579 1367 1614 1372
rect 1579 1347 1586 1367
rect 1606 1347 1614 1367
rect 1579 1339 1614 1347
rect 1347 1143 1353 1173
rect 1374 1143 1378 1173
rect 1347 1135 1378 1143
rect 1505 1117 1545 1118
rect 1135 1115 1547 1117
rect 1135 1089 1515 1115
rect 1541 1089 1547 1115
rect 1135 1081 1547 1089
rect 1135 1053 1167 1081
rect 1580 1061 1614 1339
rect 1696 1152 1766 1463
rect 2393 1454 3735 1459
rect 2393 1452 3692 1454
rect 2390 1426 3692 1452
rect 3720 1426 3735 1454
rect 2390 1418 3735 1426
rect 2390 1393 2429 1418
rect 2390 1376 2431 1393
rect 2390 1369 2429 1376
rect 1805 1307 2008 1320
rect 1805 1274 1829 1307
rect 1865 1306 2008 1307
rect 1865 1303 1976 1306
rect 1865 1276 1902 1303
rect 1931 1279 1976 1303
rect 2005 1279 2008 1306
rect 1931 1276 2008 1279
rect 1865 1274 2008 1276
rect 1805 1261 2008 1274
rect 1805 1260 1906 1261
rect 1135 1033 1140 1053
rect 1161 1033 1167 1053
rect 1135 1026 1167 1033
rect 1558 1056 1614 1061
rect 1558 1036 1565 1056
rect 1585 1036 1614 1056
rect 1691 1146 1766 1152
rect 1691 1113 1699 1146
rect 1752 1113 1766 1146
rect 1691 1088 1766 1113
rect 1691 1055 1704 1088
rect 1757 1055 1766 1088
rect 1691 1046 1766 1055
rect 2183 1198 2215 1205
rect 2183 1178 2190 1198
rect 2211 1178 2215 1198
rect 2183 1113 2215 1178
rect 2395 1169 2426 1369
rect 2630 1368 2662 1369
rect 2627 1363 2662 1368
rect 2627 1343 2634 1363
rect 2654 1343 2662 1363
rect 2627 1335 2662 1343
rect 2395 1139 2401 1169
rect 2422 1139 2426 1169
rect 2395 1131 2426 1139
rect 2553 1113 2593 1114
rect 2183 1111 2595 1113
rect 2183 1085 2563 1111
rect 2589 1085 2595 1111
rect 2183 1077 2595 1085
rect 2183 1049 2215 1077
rect 2628 1057 2662 1335
rect 1691 1041 1749 1046
rect 1558 1029 1614 1036
rect 2183 1029 2188 1049
rect 2209 1029 2215 1049
rect 1558 1028 1593 1029
rect 2183 1022 2215 1029
rect 2606 1052 2662 1057
rect 2606 1032 2613 1052
rect 2633 1032 2662 1052
rect 2606 1025 2662 1032
rect 2606 1024 2641 1025
rect 849 973 960 977
rect 2724 973 4244 974
rect 171 955 4244 973
rect 171 935 857 955
rect 876 935 934 955
rect 953 951 4244 955
rect 953 935 1905 951
rect 171 931 1905 935
rect 1924 931 1982 951
rect 2001 931 4244 951
rect 171 917 4244 931
rect 171 294 278 917
rect 1897 914 2008 917
rect 657 868 721 872
rect 653 862 721 868
rect 653 829 670 862
rect 710 829 721 862
rect 653 817 721 829
rect 1704 831 1769 853
rect 653 815 710 817
rect 657 454 708 815
rect 1704 792 1721 831
rect 1766 792 1769 831
rect 1345 747 1380 749
rect 1345 738 1449 747
rect 1345 737 1396 738
rect 1345 717 1348 737
rect 1373 718 1396 737
rect 1428 718 1449 738
rect 1373 717 1449 718
rect 1345 710 1449 717
rect 1345 698 1380 710
rect 757 632 960 645
rect 757 599 781 632
rect 817 631 960 632
rect 817 628 928 631
rect 817 601 854 628
rect 883 604 928 628
rect 957 604 960 631
rect 883 601 960 604
rect 817 599 960 601
rect 757 586 960 599
rect 757 585 858 586
rect 1135 523 1167 530
rect 1135 503 1142 523
rect 1163 503 1167 523
rect 646 445 711 454
rect 646 408 656 445
rect 696 411 711 445
rect 1135 438 1167 503
rect 1347 494 1378 698
rect 1582 693 1614 694
rect 1579 688 1614 693
rect 1579 668 1586 688
rect 1606 668 1614 688
rect 1579 660 1614 668
rect 1347 464 1353 494
rect 1374 464 1378 494
rect 1347 456 1378 464
rect 1505 438 1545 439
rect 1135 436 1547 438
rect 696 408 713 411
rect 646 389 713 408
rect 646 368 660 389
rect 696 368 713 389
rect 646 361 713 368
rect 1135 410 1515 436
rect 1541 410 1547 436
rect 1135 402 1547 410
rect 1135 374 1167 402
rect 1580 382 1614 660
rect 1704 492 1769 792
rect 1135 354 1140 374
rect 1161 354 1167 374
rect 1135 347 1167 354
rect 1558 377 1614 382
rect 1558 357 1565 377
rect 1585 357 1614 377
rect 1558 350 1614 357
rect 1694 481 1774 492
rect 1694 455 1711 481
rect 1751 455 1774 481
rect 1694 428 1774 455
rect 1694 402 1715 428
rect 1755 402 1774 428
rect 1694 383 1774 402
rect 1694 357 1718 383
rect 1758 357 1774 383
rect 1558 349 1593 350
rect 1694 345 1774 357
rect 849 294 960 298
rect 2604 294 2811 295
rect 169 276 4244 294
rect 169 256 857 276
rect 876 256 934 276
rect 953 256 4244 276
rect 169 238 4244 256
rect 171 38 278 238
rect 2766 236 4244 238
rect 639 199 760 209
rect 639 197 708 199
rect 639 156 652 197
rect 689 158 708 197
rect 745 158 760 199
rect 689 156 760 158
rect 639 138 760 156
rect 645 0 710 138
<< via1 >>
rect 780 5692 816 5725
rect 1828 5688 1864 5721
rect 780 5013 816 5046
rect 3275 5008 3311 5041
rect 780 4245 816 4278
rect 1828 4241 1864 4274
rect 780 3566 816 3599
rect 3318 3563 3354 3596
rect 781 2725 817 2758
rect 1829 2721 1865 2754
rect 781 2046 817 2079
rect 3276 2041 3312 2074
rect 781 1278 817 1311
rect 1829 1274 1865 1307
rect 781 599 817 632
<< metal2 >>
rect -1 5740 106 5981
rect -1 5725 4178 5740
rect -1 5692 780 5725
rect 816 5721 4178 5725
rect 816 5692 1828 5721
rect -1 5688 1828 5692
rect 1864 5688 4178 5721
rect -1 5671 4178 5688
rect -1 5065 106 5671
rect 2606 5669 4178 5671
rect -1 5046 4234 5065
rect -1 5013 780 5046
rect 816 5041 4234 5046
rect 816 5013 3275 5041
rect -1 5008 3275 5013
rect 3311 5008 4234 5041
rect -1 4996 4234 5008
rect -1 4293 106 4996
rect 2527 4995 4234 4996
rect 2756 4296 2999 4301
rect 2704 4293 4234 4296
rect -1 4278 4234 4293
rect -1 4245 780 4278
rect 816 4274 4234 4278
rect 816 4245 1828 4274
rect -1 4241 1828 4245
rect 1864 4241 4234 4274
rect -1 4224 4234 4241
rect -1 3618 106 4224
rect 2756 4215 2999 4224
rect 2738 3618 4234 3620
rect -1 3599 4234 3618
rect -1 3566 780 3599
rect 816 3596 4234 3599
rect 816 3566 3318 3596
rect -1 3563 3318 3566
rect 3354 3563 4234 3596
rect -1 3549 4234 3563
rect -1 3014 106 3549
rect 2738 3548 4234 3549
rect -1 3013 107 3014
rect 0 2990 107 3013
rect -2 2946 107 2990
rect 0 2773 107 2946
rect 2748 2773 2936 2775
rect 0 2758 4179 2773
rect 0 2725 781 2758
rect 817 2754 4179 2758
rect 817 2725 1829 2754
rect 0 2721 1829 2725
rect 1865 2721 4179 2754
rect 0 2704 4179 2721
rect 0 2098 107 2704
rect 2607 2702 4179 2704
rect 0 2079 4243 2098
rect 0 2046 781 2079
rect 817 2074 4243 2079
rect 817 2046 3276 2074
rect 0 2041 3276 2046
rect 3312 2041 4243 2074
rect 0 2029 4243 2041
rect 0 1326 107 2029
rect 2528 2028 4243 2029
rect 2705 1326 4244 1329
rect 0 1311 4244 1326
rect 0 1278 781 1311
rect 817 1307 4244 1311
rect 817 1278 1829 1307
rect 0 1274 1829 1278
rect 1865 1274 4244 1307
rect 0 1257 4244 1274
rect 0 651 107 1257
rect 2739 651 4244 653
rect 0 632 4244 651
rect 0 599 781 632
rect 817 599 4244 632
rect 0 582 4244 599
rect 0 36 107 582
rect 2739 581 4244 582
<< labels >>
rlabel locali 442 5932 486 5954 1 vref
rlabel metal1 178 5921 274 5954 1 gnd
rlabel metal2 2 5921 98 5954 1 vdd
rlabel metal1 657 5936 719 5963 1 d0
rlabel metal1 1703 5918 1756 5940 1 d1
rlabel metal1 2813 5981 2863 5994 1 d2
rlabel metal1 3899 3681 3908 3711 1 vout
rlabel metal1 2989 5964 3041 5983 1 d3
<< end >>
