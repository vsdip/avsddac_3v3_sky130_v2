magic
tech sky130A
timestamp 1614953301
<< nwell >>
rect 0 139 1310 288
rect 5 -291 650 -142
<< pwell >>
rect 470 383 628 394
rect 1135 383 1293 394
rect 470 288 645 383
rect 1135 288 1310 383
rect 0 33 493 139
rect 665 33 1158 139
rect 188 0 454 33
rect 853 0 1119 33
rect 475 -47 633 -36
rect 475 -142 650 -47
rect 5 -397 498 -291
rect 193 -430 459 -397
<< nmos >>
rect 548 326 598 368
rect 1213 326 1263 368
rect 47 59 97 101
rect 194 59 244 101
rect 369 59 419 101
rect 712 59 762 101
rect 859 59 909 101
rect 1034 59 1084 101
rect 553 -104 603 -62
rect 52 -371 102 -329
rect 199 -371 249 -329
rect 374 -371 424 -329
<< pmos >>
rect 47 162 97 264
rect 194 162 244 264
rect 369 162 419 264
rect 548 163 598 265
rect 712 162 762 264
rect 859 162 909 264
rect 1034 162 1084 264
rect 1213 163 1263 265
rect 52 -268 102 -166
rect 199 -268 249 -166
rect 374 -268 424 -166
rect 553 -267 603 -165
<< ndiff >>
rect 517 360 548 368
rect 517 343 523 360
rect 540 343 548 360
rect 517 326 548 343
rect 598 360 629 368
rect 598 343 604 360
rect 621 343 629 360
rect 598 326 629 343
rect 1182 360 1213 368
rect 1182 343 1188 360
rect 1205 343 1213 360
rect 1182 326 1213 343
rect 1263 360 1294 368
rect 1263 343 1269 360
rect 1286 343 1294 360
rect 1263 326 1294 343
rect 16 84 47 101
rect 16 67 24 84
rect 41 67 47 84
rect 16 59 47 67
rect 97 84 128 101
rect 97 67 105 84
rect 122 67 128 84
rect 97 59 128 67
rect 163 84 194 101
rect 163 67 171 84
rect 188 67 194 84
rect 163 59 194 67
rect 244 84 275 101
rect 244 67 252 84
rect 269 67 275 84
rect 244 59 275 67
rect 338 84 369 101
rect 338 67 346 84
rect 363 67 369 84
rect 338 59 369 67
rect 419 84 450 101
rect 419 67 427 84
rect 444 67 450 84
rect 419 59 450 67
rect 681 84 712 101
rect 681 67 689 84
rect 706 67 712 84
rect 681 59 712 67
rect 762 84 793 101
rect 762 67 770 84
rect 787 67 793 84
rect 762 59 793 67
rect 828 84 859 101
rect 828 67 836 84
rect 853 67 859 84
rect 828 59 859 67
rect 909 84 940 101
rect 909 67 917 84
rect 934 67 940 84
rect 909 59 940 67
rect 1003 84 1034 101
rect 1003 67 1011 84
rect 1028 67 1034 84
rect 1003 59 1034 67
rect 1084 84 1115 101
rect 1084 67 1092 84
rect 1109 67 1115 84
rect 1084 59 1115 67
rect 522 -70 553 -62
rect 522 -87 528 -70
rect 545 -87 553 -70
rect 522 -104 553 -87
rect 603 -70 634 -62
rect 603 -87 609 -70
rect 626 -87 634 -70
rect 603 -104 634 -87
rect 21 -346 52 -329
rect 21 -363 29 -346
rect 46 -363 52 -346
rect 21 -371 52 -363
rect 102 -346 133 -329
rect 102 -363 110 -346
rect 127 -363 133 -346
rect 102 -371 133 -363
rect 168 -346 199 -329
rect 168 -363 176 -346
rect 193 -363 199 -346
rect 168 -371 199 -363
rect 249 -346 280 -329
rect 249 -363 257 -346
rect 274 -363 280 -346
rect 249 -371 280 -363
rect 343 -346 374 -329
rect 343 -363 351 -346
rect 368 -363 374 -346
rect 343 -371 374 -363
rect 424 -346 455 -329
rect 424 -363 432 -346
rect 449 -363 455 -346
rect 424 -371 455 -363
<< pdiff >>
rect 22 213 47 264
rect 20 205 47 213
rect 20 188 24 205
rect 41 188 47 205
rect 20 162 47 188
rect 97 212 122 264
rect 169 213 194 264
rect 97 204 126 212
rect 97 187 103 204
rect 120 187 126 204
rect 97 162 126 187
rect 167 205 194 213
rect 167 188 171 205
rect 188 188 194 205
rect 167 162 194 188
rect 244 212 269 264
rect 344 213 369 264
rect 244 204 273 212
rect 244 187 250 204
rect 267 187 273 204
rect 244 162 273 187
rect 342 205 369 213
rect 342 188 346 205
rect 363 188 369 205
rect 342 162 369 188
rect 419 212 444 264
rect 519 240 548 265
rect 519 223 525 240
rect 542 223 548 240
rect 519 215 548 223
rect 419 204 448 212
rect 419 187 425 204
rect 442 187 448 204
rect 419 162 448 187
rect 523 163 548 215
rect 598 239 625 265
rect 598 222 604 239
rect 621 222 625 239
rect 598 214 625 222
rect 598 163 623 214
rect 687 213 712 264
rect 685 205 712 213
rect 685 188 689 205
rect 706 188 712 205
rect 685 162 712 188
rect 762 212 787 264
rect 834 213 859 264
rect 762 204 791 212
rect 762 187 768 204
rect 785 187 791 204
rect 762 162 791 187
rect 832 205 859 213
rect 832 188 836 205
rect 853 188 859 205
rect 832 162 859 188
rect 909 212 934 264
rect 1009 213 1034 264
rect 909 204 938 212
rect 909 187 915 204
rect 932 187 938 204
rect 909 162 938 187
rect 1007 205 1034 213
rect 1007 188 1011 205
rect 1028 188 1034 205
rect 1007 162 1034 188
rect 1084 212 1109 264
rect 1184 240 1213 265
rect 1184 223 1190 240
rect 1207 223 1213 240
rect 1184 215 1213 223
rect 1084 204 1113 212
rect 1084 187 1090 204
rect 1107 187 1113 204
rect 1084 162 1113 187
rect 1188 163 1213 215
rect 1263 239 1290 265
rect 1263 222 1269 239
rect 1286 222 1290 239
rect 1263 214 1290 222
rect 1263 163 1288 214
rect 27 -217 52 -166
rect 25 -225 52 -217
rect 25 -242 29 -225
rect 46 -242 52 -225
rect 25 -268 52 -242
rect 102 -218 127 -166
rect 174 -217 199 -166
rect 102 -226 131 -218
rect 102 -243 108 -226
rect 125 -243 131 -226
rect 102 -268 131 -243
rect 172 -225 199 -217
rect 172 -242 176 -225
rect 193 -242 199 -225
rect 172 -268 199 -242
rect 249 -218 274 -166
rect 349 -217 374 -166
rect 249 -226 278 -218
rect 249 -243 255 -226
rect 272 -243 278 -226
rect 249 -268 278 -243
rect 347 -225 374 -217
rect 347 -242 351 -225
rect 368 -242 374 -225
rect 347 -268 374 -242
rect 424 -218 449 -166
rect 524 -190 553 -165
rect 524 -207 530 -190
rect 547 -207 553 -190
rect 524 -215 553 -207
rect 424 -226 453 -218
rect 424 -243 430 -226
rect 447 -243 453 -226
rect 424 -268 453 -243
rect 528 -267 553 -215
rect 603 -191 630 -165
rect 603 -208 609 -191
rect 626 -208 630 -191
rect 603 -216 630 -208
rect 603 -267 628 -216
<< ndiffc >>
rect 523 343 540 360
rect 604 343 621 360
rect 1188 343 1205 360
rect 1269 343 1286 360
rect 24 67 41 84
rect 105 67 122 84
rect 171 67 188 84
rect 252 67 269 84
rect 346 67 363 84
rect 427 67 444 84
rect 689 67 706 84
rect 770 67 787 84
rect 836 67 853 84
rect 917 67 934 84
rect 1011 67 1028 84
rect 1092 67 1109 84
rect 528 -87 545 -70
rect 609 -87 626 -70
rect 29 -363 46 -346
rect 110 -363 127 -346
rect 176 -363 193 -346
rect 257 -363 274 -346
rect 351 -363 368 -346
rect 432 -363 449 -346
<< pdiffc >>
rect 24 188 41 205
rect 103 187 120 204
rect 171 188 188 205
rect 250 187 267 204
rect 346 188 363 205
rect 525 223 542 240
rect 425 187 442 204
rect 604 222 621 239
rect 689 188 706 205
rect 768 187 785 204
rect 836 188 853 205
rect 915 187 932 204
rect 1011 188 1028 205
rect 1190 223 1207 240
rect 1090 187 1107 204
rect 1269 222 1286 239
rect 29 -242 46 -225
rect 108 -243 125 -226
rect 176 -242 193 -225
rect 255 -243 272 -226
rect 351 -242 368 -225
rect 530 -207 547 -190
rect 430 -243 447 -226
rect 609 -208 626 -191
<< poly >>
rect 548 368 598 387
rect 1213 368 1263 387
rect 548 307 598 326
rect 548 289 563 307
rect 581 289 598 307
rect 47 264 97 278
rect 194 264 244 278
rect 369 264 419 278
rect 548 265 598 289
rect 1213 307 1263 326
rect 1213 289 1228 307
rect 1246 289 1263 307
rect 712 264 762 278
rect 859 264 909 278
rect 1034 264 1084 278
rect 1213 265 1263 289
rect 47 138 97 162
rect 47 120 64 138
rect 82 120 97 138
rect 47 101 97 120
rect 194 138 244 162
rect 194 120 211 138
rect 229 120 244 138
rect 194 101 244 120
rect 369 138 419 162
rect 548 149 598 163
rect 369 120 386 138
rect 404 120 419 138
rect 369 101 419 120
rect 712 138 762 162
rect 712 120 729 138
rect 747 120 762 138
rect 712 101 762 120
rect 859 138 909 162
rect 859 120 876 138
rect 894 120 909 138
rect 859 101 909 120
rect 1034 138 1084 162
rect 1213 149 1263 163
rect 1034 120 1051 138
rect 1069 120 1084 138
rect 1034 101 1084 120
rect 47 40 97 59
rect 194 40 244 59
rect 369 40 419 59
rect 712 40 762 59
rect 859 40 909 59
rect 1034 40 1084 59
rect 553 -62 603 -43
rect 553 -123 603 -104
rect 553 -141 568 -123
rect 586 -141 603 -123
rect 52 -166 102 -152
rect 199 -166 249 -152
rect 374 -166 424 -152
rect 553 -165 603 -141
rect 52 -292 102 -268
rect 52 -310 69 -292
rect 87 -310 102 -292
rect 52 -329 102 -310
rect 199 -292 249 -268
rect 199 -310 216 -292
rect 234 -310 249 -292
rect 199 -329 249 -310
rect 374 -292 424 -268
rect 553 -281 603 -267
rect 374 -310 391 -292
rect 409 -310 424 -292
rect 374 -329 424 -310
rect 52 -390 102 -371
rect 199 -390 249 -371
rect 374 -390 424 -371
<< polycont >>
rect 563 289 581 307
rect 1228 289 1246 307
rect 64 120 82 138
rect 211 120 229 138
rect 386 120 404 138
rect 729 120 747 138
rect 876 120 894 138
rect 1051 120 1069 138
rect 568 -141 586 -123
rect 69 -310 87 -292
rect 216 -310 234 -292
rect 391 -310 409 -292
<< locali >>
rect 338 395 629 419
rect 338 374 367 395
rect 17 288 193 304
rect 339 288 367 374
rect 500 360 548 368
rect 500 343 523 360
rect 540 343 548 360
rect 500 335 548 343
rect 597 360 629 395
rect 1003 395 1294 419
rect 1003 374 1032 395
rect 597 343 604 360
rect 621 343 629 360
rect 597 335 629 343
rect 1004 352 1032 374
rect 17 282 194 288
rect 17 213 47 282
rect 164 213 194 282
rect 339 213 369 288
rect 500 248 517 335
rect 1004 331 1008 352
rect 1029 331 1032 352
rect 557 311 645 315
rect 557 307 615 311
rect 557 289 563 307
rect 581 290 615 307
rect 636 290 645 311
rect 581 289 645 290
rect 557 281 645 289
rect 682 288 858 304
rect 1004 288 1032 331
rect 1165 360 1213 368
rect 1165 343 1188 360
rect 1205 343 1213 360
rect 1165 335 1213 343
rect 1262 360 1294 395
rect 1262 343 1269 360
rect 1286 343 1294 360
rect 1262 335 1294 343
rect 682 282 859 288
rect 500 240 548 248
rect 464 234 525 240
rect 16 205 47 213
rect 16 188 24 205
rect 41 188 47 205
rect 16 180 47 188
rect 17 178 47 180
rect 97 204 145 212
rect 97 187 103 204
rect 120 187 145 204
rect 97 179 145 187
rect 163 205 194 213
rect 163 188 171 205
rect 188 188 194 205
rect 163 180 194 188
rect 128 146 145 179
rect 164 178 194 180
rect 244 211 292 212
rect 244 206 318 211
rect 244 204 286 206
rect 244 187 250 204
rect 267 187 286 204
rect 244 185 286 187
rect 307 185 318 206
rect 244 179 318 185
rect 338 205 369 213
rect 449 213 474 234
rect 495 223 525 234
rect 542 234 548 240
rect 598 247 628 249
rect 598 239 629 247
rect 542 223 549 234
rect 495 213 549 223
rect 449 212 549 213
rect 598 222 604 239
rect 621 222 629 239
rect 598 214 629 222
rect 338 188 346 205
rect 363 188 369 205
rect 338 180 369 188
rect 0 138 88 146
rect 0 120 64 138
rect 82 120 88 138
rect 0 112 88 120
rect 128 139 235 146
rect 128 119 161 139
rect 181 138 235 139
rect 181 120 211 138
rect 229 120 235 138
rect 181 119 235 120
rect 128 112 235 119
rect 128 92 145 112
rect 275 92 292 179
rect 339 178 369 180
rect 419 207 505 212
rect 419 204 467 207
rect 419 187 425 204
rect 442 187 467 204
rect 419 179 467 187
rect 322 140 410 146
rect 322 120 336 140
rect 356 138 410 140
rect 356 120 386 138
rect 404 120 410 138
rect 322 112 410 120
rect 450 92 467 179
rect 598 139 628 214
rect 682 213 712 282
rect 829 213 859 282
rect 1004 213 1034 288
rect 1165 248 1182 335
rect 1222 311 1310 315
rect 1222 307 1280 311
rect 1222 289 1228 307
rect 1246 290 1280 307
rect 1301 290 1310 311
rect 1246 289 1310 290
rect 1222 281 1310 289
rect 1165 240 1213 248
rect 1165 234 1190 240
rect 681 205 712 213
rect 681 188 689 205
rect 706 188 712 205
rect 681 180 712 188
rect 682 178 712 180
rect 762 204 810 212
rect 762 187 768 204
rect 785 187 810 204
rect 762 179 810 187
rect 828 205 859 213
rect 828 188 836 205
rect 853 188 859 205
rect 828 180 859 188
rect 793 146 810 179
rect 829 178 859 180
rect 909 211 957 212
rect 909 206 983 211
rect 909 204 951 206
rect 909 187 915 204
rect 932 187 951 204
rect 909 185 951 187
rect 972 185 983 206
rect 909 179 983 185
rect 1003 205 1034 213
rect 1114 223 1190 234
rect 1207 234 1213 240
rect 1263 247 1293 249
rect 1263 239 1294 247
rect 1207 223 1214 234
rect 1114 212 1214 223
rect 1263 222 1269 239
rect 1286 222 1294 239
rect 1263 214 1294 222
rect 1003 188 1011 205
rect 1028 188 1034 205
rect 1003 180 1034 188
rect 16 84 48 92
rect 16 67 24 84
rect 41 67 48 84
rect 16 59 48 67
rect 97 84 145 92
rect 97 67 105 84
rect 122 67 145 84
rect 97 59 145 67
rect 163 84 195 92
rect 163 67 171 84
rect 188 67 195 84
rect 163 59 195 67
rect 244 84 292 92
rect 244 67 252 84
rect 269 67 292 84
rect 244 59 292 67
rect 338 84 370 92
rect 338 67 346 84
rect 363 67 370 84
rect 338 59 370 67
rect 419 84 467 92
rect 419 67 427 84
rect 444 67 467 84
rect 419 59 467 67
rect 17 39 48 59
rect 164 39 195 59
rect 16 15 196 39
rect 339 33 370 59
rect 605 33 625 139
rect 665 138 753 146
rect 665 120 729 138
rect 747 120 753 138
rect 665 112 753 120
rect 793 139 900 146
rect 793 119 826 139
rect 846 138 900 139
rect 846 120 876 138
rect 894 120 900 138
rect 846 119 900 120
rect 793 112 900 119
rect 793 92 810 112
rect 940 92 957 179
rect 1004 178 1034 180
rect 1084 204 1132 212
rect 1084 187 1090 204
rect 1107 187 1132 204
rect 1084 179 1132 187
rect 987 140 1075 146
rect 987 120 1001 140
rect 1021 138 1075 140
rect 1021 120 1051 138
rect 1069 120 1075 138
rect 987 112 1075 120
rect 1115 92 1132 179
rect 1263 139 1293 214
rect 681 84 713 92
rect 681 67 689 84
rect 706 67 713 84
rect 681 59 713 67
rect 762 84 810 92
rect 762 67 770 84
rect 787 67 810 84
rect 762 59 810 67
rect 828 84 860 92
rect 828 67 836 84
rect 853 67 860 84
rect 828 59 860 67
rect 909 84 957 92
rect 909 67 917 84
rect 934 67 957 84
rect 909 59 957 67
rect 1003 84 1035 92
rect 1003 67 1011 84
rect 1028 67 1035 84
rect 1003 59 1035 67
rect 1084 84 1132 92
rect 1084 67 1092 84
rect 1109 67 1132 84
rect 1084 59 1132 67
rect 682 39 713 59
rect 829 39 860 59
rect 338 13 625 33
rect 681 15 861 39
rect 1004 33 1035 59
rect 1121 33 1159 38
rect 1270 33 1290 139
rect 1003 30 1290 33
rect 1003 13 1128 30
rect 605 12 625 13
rect 1121 7 1128 13
rect 1151 13 1290 30
rect 1151 7 1159 13
rect 1270 12 1290 13
rect 1121 -2 1159 7
rect 343 -35 634 -11
rect 343 -56 372 -35
rect 22 -142 198 -126
rect 344 -142 372 -56
rect 505 -70 553 -62
rect 505 -87 528 -70
rect 545 -87 553 -70
rect 505 -95 553 -87
rect 602 -70 634 -35
rect 602 -87 609 -70
rect 626 -87 634 -70
rect 602 -95 634 -87
rect 22 -148 199 -142
rect 22 -217 52 -148
rect 169 -217 199 -148
rect 344 -217 374 -142
rect 505 -182 522 -95
rect 562 -119 650 -115
rect 562 -123 620 -119
rect 562 -141 568 -123
rect 586 -140 620 -123
rect 641 -140 650 -119
rect 586 -141 650 -140
rect 562 -149 650 -141
rect 505 -187 553 -182
rect 471 -190 553 -187
rect 471 -193 530 -190
rect 471 -196 481 -193
rect 21 -225 52 -217
rect 21 -242 29 -225
rect 46 -242 52 -225
rect 21 -250 52 -242
rect 22 -252 52 -250
rect 102 -226 150 -218
rect 102 -243 108 -226
rect 125 -243 150 -226
rect 102 -251 150 -243
rect 168 -225 199 -217
rect 168 -242 176 -225
rect 193 -242 199 -225
rect 168 -250 199 -242
rect 133 -284 150 -251
rect 169 -252 199 -250
rect 249 -219 297 -218
rect 249 -224 323 -219
rect 249 -226 291 -224
rect 249 -243 255 -226
rect 272 -243 291 -226
rect 249 -245 291 -243
rect 312 -245 323 -224
rect 249 -251 323 -245
rect 343 -225 374 -217
rect 454 -214 481 -196
rect 502 -207 530 -193
rect 547 -196 553 -190
rect 603 -183 633 -181
rect 603 -191 634 -183
rect 547 -207 554 -196
rect 502 -214 554 -207
rect 454 -218 554 -214
rect 603 -208 609 -191
rect 626 -208 634 -191
rect 603 -216 634 -208
rect 343 -242 351 -225
rect 368 -242 374 -225
rect 343 -250 374 -242
rect 5 -292 93 -284
rect 5 -310 69 -292
rect 87 -310 93 -292
rect 5 -318 93 -310
rect 133 -291 240 -284
rect 133 -311 166 -291
rect 186 -292 240 -291
rect 186 -310 216 -292
rect 234 -310 240 -292
rect 186 -311 240 -310
rect 133 -318 240 -311
rect 133 -338 150 -318
rect 280 -338 297 -251
rect 344 -252 374 -250
rect 424 -220 512 -218
rect 424 -226 472 -220
rect 424 -243 430 -226
rect 447 -243 472 -226
rect 424 -251 472 -243
rect 327 -290 415 -284
rect 327 -310 341 -290
rect 361 -292 415 -290
rect 361 -310 391 -292
rect 409 -310 415 -292
rect 327 -318 415 -310
rect 455 -338 472 -251
rect 603 -291 633 -216
rect 21 -346 53 -338
rect 21 -363 29 -346
rect 46 -363 53 -346
rect 21 -371 53 -363
rect 102 -346 150 -338
rect 102 -363 110 -346
rect 127 -363 150 -346
rect 102 -371 150 -363
rect 168 -346 200 -338
rect 168 -363 176 -346
rect 193 -363 200 -346
rect 168 -371 200 -363
rect 249 -346 297 -338
rect 249 -363 257 -346
rect 274 -363 297 -346
rect 249 -371 297 -363
rect 343 -346 375 -338
rect 343 -363 351 -346
rect 368 -363 375 -346
rect 343 -371 375 -363
rect 424 -346 472 -338
rect 424 -363 432 -346
rect 449 -363 472 -346
rect 424 -371 472 -363
rect 22 -391 53 -371
rect 169 -391 200 -371
rect 21 -415 201 -391
rect 344 -397 375 -371
rect 610 -397 630 -291
rect 343 -417 630 -397
rect 610 -418 630 -417
<< viali >>
rect 1008 331 1029 352
rect 615 290 636 311
rect 286 185 307 206
rect 474 213 495 234
rect 161 119 181 139
rect 336 120 356 140
rect 1280 290 1301 311
rect 951 185 972 206
rect 826 119 846 139
rect 1001 120 1021 140
rect 1128 7 1151 30
rect 620 -140 641 -119
rect 291 -245 312 -224
rect 481 -214 502 -193
rect 166 -311 186 -291
rect 341 -310 361 -290
<< metal1 >>
rect 1004 353 1038 362
rect 857 352 1038 353
rect 857 331 1008 352
rect 1029 331 1038 352
rect 857 328 1038 331
rect 599 312 643 316
rect 282 311 643 312
rect 282 290 615 311
rect 636 290 643 311
rect 282 288 643 290
rect 282 212 311 288
rect 599 283 643 288
rect 464 238 505 240
rect 859 238 892 328
rect 1004 326 1038 328
rect 1264 312 1308 316
rect 464 234 892 238
rect 464 213 474 234
rect 495 214 892 234
rect 947 311 1308 312
rect 947 290 1280 311
rect 1301 290 1308 311
rect 947 288 1308 290
rect 495 213 891 214
rect 464 212 891 213
rect 947 212 976 288
rect 1264 283 1308 288
rect 275 206 319 212
rect 464 207 505 212
rect 275 185 286 206
rect 307 185 319 206
rect 275 179 319 185
rect 940 206 984 212
rect 940 185 951 206
rect 972 185 984 206
rect 940 179 984 185
rect 150 139 192 146
rect 150 119 161 139
rect 181 138 192 139
rect 323 140 365 146
rect 323 138 336 140
rect 181 124 336 138
rect 181 119 192 124
rect 150 112 192 119
rect 323 120 336 124
rect 356 120 365 140
rect 323 112 365 120
rect 815 139 857 146
rect 815 119 826 139
rect 846 138 857 139
rect 988 140 1030 146
rect 988 138 1001 140
rect 846 124 1001 138
rect 846 119 857 124
rect 815 112 857 119
rect 988 120 1001 124
rect 1021 120 1030 140
rect 988 112 1030 120
rect 1123 30 1157 36
rect 1123 7 1128 30
rect 1151 7 1157 30
rect 1123 0 1157 7
rect 604 -118 648 -114
rect 287 -119 648 -118
rect 287 -140 620 -119
rect 641 -140 648 -119
rect 287 -142 648 -140
rect 287 -218 316 -142
rect 604 -147 648 -142
rect 471 -193 512 -187
rect 471 -214 481 -193
rect 502 -194 512 -193
rect 1126 -194 1155 0
rect 502 -214 1155 -194
rect 280 -224 324 -218
rect 471 -220 1155 -214
rect 472 -222 1155 -220
rect 280 -245 291 -224
rect 312 -245 324 -224
rect 280 -251 324 -245
rect 155 -291 197 -284
rect 155 -311 166 -291
rect 186 -292 197 -291
rect 328 -290 370 -284
rect 328 -292 341 -290
rect 186 -306 341 -292
rect 186 -311 197 -306
rect 155 -318 197 -311
rect 328 -310 341 -306
rect 361 -310 370 -290
rect 328 -318 370 -310
<< labels >>
rlabel nwell 30 277 30 277 1 vdd
rlabel pwell 32 43 32 43 1 Gnd
rlabel pwell 179 43 179 43 1 Gnd
rlabel nwell 177 277 177 277 1 vdd
rlabel locali 352 277 352 277 1 vin1
rlabel locali 354 43 354 43 1 vin2
rlabel pwell 274 20 274 20 1 Gnd
rlabel nwell 465 272 465 272 1 vdd
rlabel pwell 495 383 495 383 1 Gnd
rlabel pwell 500 -47 500 -47 1 Gnd
rlabel nwell 470 -158 470 -158 1 vdd
rlabel pwell 279 -410 279 -410 1 Gnd
rlabel nwell 182 -153 182 -153 1 vdd
rlabel pwell 184 -387 184 -387 1 Gnd
rlabel pwell 37 -387 37 -387 1 Gnd
rlabel nwell 35 -153 35 -153 1 vdd
rlabel nwell 695 277 695 277 1 vdd
rlabel pwell 697 43 697 43 1 Gnd
rlabel pwell 844 43 844 43 1 Gnd
rlabel nwell 842 277 842 277 1 vdd
rlabel locali 1172 227 1172 227 5 out
rlabel pwell 939 20 939 20 1 Gnd
rlabel nwell 1130 272 1130 272 1 vdd
rlabel pwell 1160 383 1160 383 1 Gnd
rlabel locali 6 127 6 127 1 d0
rlabel locali 11 -303 11 -303 1 d0
rlabel locali 356 -80 356 -80 1 vin3
rlabel locali 359 -387 359 -387 1 vin4
rlabel locali 671 127 671 127 1 d1
rlabel metal1 606 297 606 297 1 d0
rlabel metal1 614 -131 614 -131 1 d0
rlabel metal1 1267 297 1267 297 1 d1
<< end >>
