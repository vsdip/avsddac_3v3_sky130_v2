* SPICE3 file created from 3bit_DAC.ext - technology: sky130A

.option scale=10000u

X0 a_431_177# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1 a_117_n262# a_646_n372# a_854_n372# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2 a_852_177# a_1583_487# a_1791_487# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3 a_1791_487# a_1370_487# a_853_731# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4 a_646_n372# a_433_n372# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5 a_645_n926# a_432_n926# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6 a_116_841# a_116_612# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7 a_432_731# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8 a_1370_487# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9 a_117_n75# a_117_n262# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X10 a_433_n372# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X11 a_432_n926# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X12 a_1583_487# a_1370_487# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X13 a_431_177# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X14 a_1584_n616# a_1371_n616# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X15 a_1791_487# a_1724_n105# vout gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X16 a_1371_n616# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X17 vout a_1511_n105# a_1792_n616# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X18 a_853_n926# a_432_n926# a_117_n721# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X19 a_116_382# a_117_n75# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X20 a_1792_n616# a_1371_n616# a_853_n926# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X21 a_646_n372# a_433_n372# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X22 a_117_n491# a_117_n721# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X23 a_432_731# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X24 a_433_n372# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X25 a_1511_n105# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X26 a_853_n926# a_1584_n616# a_1792_n616# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X27 vout a_1511_n105# a_1791_487# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X28 a_116_612# a_116_382# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X29 a_852_177# a_431_177# a_117_n75# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X30 a_116_382# a_644_177# a_852_177# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X31 a_854_n372# a_433_n372# a_117_n262# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X32 a_117_n721# gnd gnd sky130_fd_pr__res_generic_nd w=17 l=81
X33 a_853_n926# a_432_n926# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X34 a_644_177# a_431_177# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X35 a_853_731# a_1583_487# a_1791_487# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X36 gnd a_645_n926# a_853_n926# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X37 vref a_116_841# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X38 a_853_731# a_432_731# a_116_612# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X39 a_1583_487# a_1370_487# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X40 a_1370_487# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X41 a_1791_487# a_1370_487# a_852_177# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X42 a_852_177# a_431_177# a_116_382# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X43 a_1792_n616# a_1724_n105# vout vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X44 a_117_n262# a_117_n491# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X45 a_645_731# a_432_731# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X46 a_116_841# a_645_731# a_853_731# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X47 a_117_n75# a_644_177# a_852_177# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X48 a_1724_n105# a_1511_n105# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X49 a_1724_n105# a_1511_n105# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X50 a_644_177# a_431_177# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X51 a_1511_n105# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X52 a_854_n372# a_433_n372# a_117_n491# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X53 a_1371_n616# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X54 a_1584_n616# a_1371_n616# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X55 a_117_n721# a_645_n926# a_853_n926# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X56 a_117_n491# a_646_n372# a_854_n372# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X57 a_1792_n616# a_1371_n616# a_854_n372# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X58 a_853_731# a_432_731# a_116_841# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X59 a_645_731# a_432_731# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X60 a_116_612# a_645_731# a_853_731# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X61 a_854_n372# a_1584_n616# a_1792_n616# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X62 a_645_n926# a_432_n926# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X63 a_432_n926# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
C0 a_117_n721# gnd 2.75fF
C1 a_853_n926# gnd 2.79fF
C2 a_117_n491# gnd 2.38fF
C3 a_854_n372# gnd 2.18fF
C4 a_117_n262# gnd 2.28fF
C5 a_117_n75# gnd 2.49fF
C6 a_116_382# gnd 2.23fF
C7 a_852_177# gnd 2.52fF
C8 a_116_612# gnd 2.38fF
C9 a_853_731# gnd 2.38fF
C10 a_116_841# gnd 2.22fF
C11 vdd gnd 11.40fF
