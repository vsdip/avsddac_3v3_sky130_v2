magic
tech sky130A
timestamp 1633277651
<< nwell >>
rect 749 1119 1560 1343
rect 1797 1115 2608 1339
rect 749 440 1560 664
<< nmos >>
rect 813 1018 863 1060
rect 1026 1018 1076 1060
rect 1234 1018 1284 1060
rect 1442 1018 1492 1060
rect 1861 1014 1911 1056
rect 2074 1014 2124 1056
rect 2282 1014 2332 1056
rect 2490 1014 2540 1056
rect 813 339 863 381
rect 1026 339 1076 381
rect 1234 339 1284 381
rect 1442 339 1492 381
<< pmos >>
rect 813 1137 863 1237
rect 1026 1137 1076 1237
rect 1234 1137 1284 1237
rect 1442 1137 1492 1237
rect 1861 1133 1911 1233
rect 2074 1133 2124 1233
rect 2282 1133 2332 1233
rect 2490 1133 2540 1233
rect 813 458 863 558
rect 1026 458 1076 558
rect 1234 458 1284 558
rect 1442 458 1492 558
<< ndiff >>
rect 764 1050 813 1060
rect 764 1030 775 1050
rect 795 1030 813 1050
rect 764 1018 813 1030
rect 863 1054 907 1060
rect 863 1034 878 1054
rect 898 1034 907 1054
rect 863 1018 907 1034
rect 977 1050 1026 1060
rect 977 1030 988 1050
rect 1008 1030 1026 1050
rect 977 1018 1026 1030
rect 1076 1054 1120 1060
rect 1076 1034 1091 1054
rect 1111 1034 1120 1054
rect 1076 1018 1120 1034
rect 1185 1050 1234 1060
rect 1185 1030 1196 1050
rect 1216 1030 1234 1050
rect 1185 1018 1234 1030
rect 1284 1054 1328 1060
rect 1284 1034 1299 1054
rect 1319 1034 1328 1054
rect 1284 1018 1328 1034
rect 1398 1054 1442 1060
rect 1398 1034 1407 1054
rect 1427 1034 1442 1054
rect 1398 1018 1442 1034
rect 1492 1050 1541 1060
rect 1492 1030 1510 1050
rect 1530 1030 1541 1050
rect 1492 1018 1541 1030
rect 1812 1046 1861 1056
rect 1812 1026 1823 1046
rect 1843 1026 1861 1046
rect 1812 1014 1861 1026
rect 1911 1050 1955 1056
rect 1911 1030 1926 1050
rect 1946 1030 1955 1050
rect 1911 1014 1955 1030
rect 2025 1046 2074 1056
rect 2025 1026 2036 1046
rect 2056 1026 2074 1046
rect 2025 1014 2074 1026
rect 2124 1050 2168 1056
rect 2124 1030 2139 1050
rect 2159 1030 2168 1050
rect 2124 1014 2168 1030
rect 2233 1046 2282 1056
rect 2233 1026 2244 1046
rect 2264 1026 2282 1046
rect 2233 1014 2282 1026
rect 2332 1050 2376 1056
rect 2332 1030 2347 1050
rect 2367 1030 2376 1050
rect 2332 1014 2376 1030
rect 2446 1050 2490 1056
rect 2446 1030 2455 1050
rect 2475 1030 2490 1050
rect 2446 1014 2490 1030
rect 2540 1046 2589 1056
rect 2540 1026 2558 1046
rect 2578 1026 2589 1046
rect 2540 1014 2589 1026
rect 764 371 813 381
rect 764 351 775 371
rect 795 351 813 371
rect 764 339 813 351
rect 863 375 907 381
rect 863 355 878 375
rect 898 355 907 375
rect 863 339 907 355
rect 977 371 1026 381
rect 977 351 988 371
rect 1008 351 1026 371
rect 977 339 1026 351
rect 1076 375 1120 381
rect 1076 355 1091 375
rect 1111 355 1120 375
rect 1076 339 1120 355
rect 1185 371 1234 381
rect 1185 351 1196 371
rect 1216 351 1234 371
rect 1185 339 1234 351
rect 1284 375 1328 381
rect 1284 355 1299 375
rect 1319 355 1328 375
rect 1284 339 1328 355
rect 1398 375 1442 381
rect 1398 355 1407 375
rect 1427 355 1442 375
rect 1398 339 1442 355
rect 1492 371 1541 381
rect 1492 351 1510 371
rect 1530 351 1541 371
rect 1492 339 1541 351
<< pdiff >>
rect 769 1199 813 1237
rect 769 1179 781 1199
rect 801 1179 813 1199
rect 769 1137 813 1179
rect 863 1199 905 1237
rect 863 1179 877 1199
rect 897 1179 905 1199
rect 863 1137 905 1179
rect 982 1199 1026 1237
rect 982 1179 994 1199
rect 1014 1179 1026 1199
rect 982 1137 1026 1179
rect 1076 1199 1118 1237
rect 1076 1179 1090 1199
rect 1110 1179 1118 1199
rect 1076 1137 1118 1179
rect 1190 1199 1234 1237
rect 1190 1179 1202 1199
rect 1222 1179 1234 1199
rect 1190 1137 1234 1179
rect 1284 1199 1326 1237
rect 1284 1179 1298 1199
rect 1318 1179 1326 1199
rect 1284 1137 1326 1179
rect 1400 1199 1442 1237
rect 1400 1179 1408 1199
rect 1428 1179 1442 1199
rect 1400 1137 1442 1179
rect 1492 1206 1537 1237
rect 1492 1199 1536 1206
rect 1492 1179 1504 1199
rect 1524 1179 1536 1199
rect 1492 1137 1536 1179
rect 1817 1195 1861 1233
rect 1817 1175 1829 1195
rect 1849 1175 1861 1195
rect 1817 1133 1861 1175
rect 1911 1195 1953 1233
rect 1911 1175 1925 1195
rect 1945 1175 1953 1195
rect 1911 1133 1953 1175
rect 2030 1195 2074 1233
rect 2030 1175 2042 1195
rect 2062 1175 2074 1195
rect 2030 1133 2074 1175
rect 2124 1195 2166 1233
rect 2124 1175 2138 1195
rect 2158 1175 2166 1195
rect 2124 1133 2166 1175
rect 2238 1195 2282 1233
rect 2238 1175 2250 1195
rect 2270 1175 2282 1195
rect 2238 1133 2282 1175
rect 2332 1195 2374 1233
rect 2332 1175 2346 1195
rect 2366 1175 2374 1195
rect 2332 1133 2374 1175
rect 2448 1195 2490 1233
rect 2448 1175 2456 1195
rect 2476 1175 2490 1195
rect 2448 1133 2490 1175
rect 2540 1202 2585 1233
rect 2540 1195 2584 1202
rect 2540 1175 2552 1195
rect 2572 1175 2584 1195
rect 2540 1133 2584 1175
rect 769 520 813 558
rect 769 500 781 520
rect 801 500 813 520
rect 769 458 813 500
rect 863 520 905 558
rect 863 500 877 520
rect 897 500 905 520
rect 863 458 905 500
rect 982 520 1026 558
rect 982 500 994 520
rect 1014 500 1026 520
rect 982 458 1026 500
rect 1076 520 1118 558
rect 1076 500 1090 520
rect 1110 500 1118 520
rect 1076 458 1118 500
rect 1190 520 1234 558
rect 1190 500 1202 520
rect 1222 500 1234 520
rect 1190 458 1234 500
rect 1284 520 1326 558
rect 1284 500 1298 520
rect 1318 500 1326 520
rect 1284 458 1326 500
rect 1400 520 1442 558
rect 1400 500 1408 520
rect 1428 500 1442 520
rect 1400 458 1442 500
rect 1492 527 1537 558
rect 1492 520 1536 527
rect 1492 500 1504 520
rect 1524 500 1536 520
rect 1492 458 1536 500
<< ndiffc >>
rect 455 1353 473 1371
rect 457 1254 475 1272
rect 455 1097 473 1115
rect 775 1030 795 1050
rect 878 1034 898 1054
rect 988 1030 1008 1050
rect 1091 1034 1111 1054
rect 1196 1030 1216 1050
rect 1299 1034 1319 1054
rect 1407 1034 1427 1054
rect 1510 1030 1530 1050
rect 1823 1026 1843 1046
rect 457 998 475 1016
rect 1926 1030 1946 1050
rect 2036 1026 2056 1046
rect 2139 1030 2159 1050
rect 2244 1026 2264 1046
rect 2347 1030 2367 1050
rect 2455 1030 2475 1050
rect 2558 1026 2578 1046
rect 455 702 473 720
rect 457 603 475 621
rect 455 447 473 465
rect 457 348 475 366
rect 775 351 795 371
rect 878 355 898 375
rect 988 351 1008 371
rect 1091 355 1111 375
rect 1196 351 1216 371
rect 1299 355 1319 375
rect 1407 355 1427 375
rect 1510 351 1530 371
<< pdiffc >>
rect 781 1179 801 1199
rect 877 1179 897 1199
rect 994 1179 1014 1199
rect 1090 1179 1110 1199
rect 1202 1179 1222 1199
rect 1298 1179 1318 1199
rect 1408 1179 1428 1199
rect 1504 1179 1524 1199
rect 1829 1175 1849 1195
rect 1925 1175 1945 1195
rect 2042 1175 2062 1195
rect 2138 1175 2158 1195
rect 2250 1175 2270 1195
rect 2346 1175 2366 1195
rect 2456 1175 2476 1195
rect 2552 1175 2572 1195
rect 781 500 801 520
rect 877 500 897 520
rect 994 500 1014 520
rect 1090 500 1110 520
rect 1202 500 1222 520
rect 1298 500 1318 520
rect 1408 500 1428 520
rect 1504 500 1524 520
<< psubdiff >>
rect 849 963 960 977
rect 849 933 890 963
rect 918 933 960 963
rect 849 918 960 933
rect 1897 959 2008 973
rect 1897 929 1938 959
rect 1966 929 2008 959
rect 1897 914 2008 929
rect 849 284 960 298
rect 849 254 890 284
rect 918 254 960 284
rect 849 239 960 254
<< nsubdiff >>
rect 850 1310 960 1324
rect 850 1280 893 1310
rect 921 1280 960 1310
rect 850 1265 960 1280
rect 1898 1306 2008 1320
rect 1898 1276 1941 1306
rect 1969 1276 2008 1306
rect 1898 1261 2008 1276
rect 850 631 960 645
rect 850 601 893 631
rect 921 601 960 631
rect 850 586 960 601
<< psubdiffcont >>
rect 890 933 918 963
rect 1938 929 1966 959
rect 890 254 918 284
<< nsubdiffcont >>
rect 893 1280 921 1310
rect 1941 1276 1969 1306
rect 893 601 921 631
<< poly >>
rect 813 1237 863 1250
rect 1026 1237 1076 1250
rect 1234 1237 1284 1250
rect 1442 1237 1492 1250
rect 1861 1233 1911 1246
rect 2074 1233 2124 1246
rect 2282 1233 2332 1246
rect 2490 1233 2540 1246
rect 813 1109 863 1137
rect 813 1089 826 1109
rect 846 1089 863 1109
rect 813 1060 863 1089
rect 1026 1108 1076 1137
rect 1026 1084 1037 1108
rect 1061 1084 1076 1108
rect 1026 1060 1076 1084
rect 1234 1113 1284 1137
rect 1234 1089 1246 1113
rect 1270 1089 1284 1113
rect 1234 1060 1284 1089
rect 1442 1111 1492 1137
rect 1442 1085 1460 1111
rect 1486 1085 1492 1111
rect 1442 1060 1492 1085
rect 1861 1105 1911 1133
rect 1861 1085 1874 1105
rect 1894 1085 1911 1105
rect 1861 1056 1911 1085
rect 2074 1104 2124 1133
rect 2074 1080 2085 1104
rect 2109 1080 2124 1104
rect 2074 1056 2124 1080
rect 2282 1109 2332 1133
rect 2282 1085 2294 1109
rect 2318 1085 2332 1109
rect 2282 1056 2332 1085
rect 2490 1107 2540 1133
rect 2490 1081 2508 1107
rect 2534 1081 2540 1107
rect 2490 1056 2540 1081
rect 813 1002 863 1018
rect 1026 1002 1076 1018
rect 1234 1002 1284 1018
rect 1442 1002 1492 1018
rect 1861 998 1911 1014
rect 2074 998 2124 1014
rect 2282 998 2332 1014
rect 2490 998 2540 1014
rect 813 558 863 571
rect 1026 558 1076 571
rect 1234 558 1284 571
rect 1442 558 1492 571
rect 813 430 863 458
rect 813 410 826 430
rect 846 410 863 430
rect 813 381 863 410
rect 1026 429 1076 458
rect 1026 405 1037 429
rect 1061 405 1076 429
rect 1026 381 1076 405
rect 1234 434 1284 458
rect 1234 410 1246 434
rect 1270 410 1284 434
rect 1234 381 1284 410
rect 1442 432 1492 458
rect 1442 406 1460 432
rect 1486 406 1492 432
rect 1442 381 1492 406
rect 813 323 863 339
rect 1026 323 1076 339
rect 1234 323 1284 339
rect 1442 323 1492 339
<< polycont >>
rect 826 1089 846 1109
rect 1037 1084 1061 1108
rect 1246 1089 1270 1113
rect 1460 1085 1486 1111
rect 1874 1085 1894 1105
rect 2085 1080 2109 1104
rect 2294 1085 2318 1109
rect 2508 1081 2534 1107
rect 826 410 846 430
rect 1037 405 1061 429
rect 1246 410 1270 434
rect 1460 406 1486 432
<< ndiffres >>
rect 434 1371 491 1390
rect 434 1368 455 1371
rect 340 1353 455 1368
rect 473 1353 491 1371
rect 340 1330 491 1353
rect 340 1294 382 1330
rect 339 1293 439 1294
rect 339 1272 495 1293
rect 339 1254 457 1272
rect 475 1254 495 1272
rect 339 1250 495 1254
rect 434 1234 495 1250
rect 434 1115 491 1134
rect 434 1112 455 1115
rect 340 1097 455 1112
rect 473 1097 491 1115
rect 340 1074 491 1097
rect 340 1038 382 1074
rect 339 1037 439 1038
rect 339 1016 495 1037
rect 339 998 457 1016
rect 475 998 495 1016
rect 339 994 495 998
rect 434 978 495 994
rect 434 720 491 739
rect 434 717 455 720
rect 340 702 455 717
rect 473 702 491 720
rect 340 679 491 702
rect 340 643 382 679
rect 339 642 439 643
rect 339 621 495 642
rect 339 603 457 621
rect 475 603 495 621
rect 339 599 495 603
rect 434 583 495 599
rect 434 465 491 484
rect 434 462 455 465
rect 340 447 455 462
rect 473 447 491 465
rect 340 424 491 447
rect 340 388 382 424
rect 339 387 439 388
rect 339 366 495 387
rect 339 348 457 366
rect 475 348 495 366
rect 339 344 495 348
rect 434 328 495 344
<< locali >>
rect 433 1371 492 1477
rect 2396 1453 2468 1454
rect 1346 1452 1418 1453
rect 1345 1444 1444 1452
rect 1345 1441 1397 1444
rect 1345 1406 1353 1441
rect 1378 1406 1397 1441
rect 1422 1433 1444 1444
rect 2395 1445 2494 1453
rect 2395 1442 2447 1445
rect 1422 1432 2289 1433
rect 1422 1406 2290 1432
rect 1345 1396 2290 1406
rect 1345 1394 1444 1396
rect 433 1353 455 1371
rect 473 1353 492 1371
rect 433 1331 492 1353
rect 700 1367 1232 1372
rect 700 1347 1586 1367
rect 1606 1347 1609 1367
rect 2245 1363 2290 1396
rect 2395 1407 2403 1442
rect 2428 1407 2447 1442
rect 2472 1407 2494 1445
rect 2395 1395 2494 1407
rect 700 1343 1609 1347
rect 700 1296 743 1343
rect 1193 1342 1609 1343
rect 2241 1343 2634 1363
rect 2654 1343 2657 1363
rect 1193 1341 1534 1342
rect 850 1310 960 1324
rect 850 1307 893 1310
rect 850 1302 854 1307
rect 688 1295 743 1296
rect 432 1272 743 1295
rect 432 1254 457 1272
rect 475 1260 743 1272
rect 772 1280 854 1302
rect 883 1280 893 1307
rect 921 1283 928 1310
rect 957 1302 960 1310
rect 957 1283 1022 1302
rect 921 1280 1022 1283
rect 772 1278 1022 1280
rect 475 1254 497 1260
rect 432 1115 497 1254
rect 772 1199 809 1278
rect 850 1265 960 1278
rect 924 1209 955 1210
rect 772 1179 781 1199
rect 801 1179 809 1199
rect 432 1097 455 1115
rect 473 1097 497 1115
rect 432 1080 497 1097
rect 652 1161 720 1174
rect 772 1169 809 1179
rect 868 1199 955 1209
rect 868 1179 877 1199
rect 897 1179 955 1199
rect 868 1170 955 1179
rect 868 1169 905 1170
rect 652 1119 659 1161
rect 708 1119 720 1161
rect 652 1116 720 1119
rect 924 1117 955 1170
rect 985 1199 1022 1278
rect 1137 1209 1168 1210
rect 985 1179 994 1199
rect 1014 1179 1022 1199
rect 985 1169 1022 1179
rect 1081 1202 1168 1209
rect 1081 1199 1142 1202
rect 1081 1179 1090 1199
rect 1110 1182 1142 1199
rect 1163 1182 1168 1202
rect 1110 1179 1168 1182
rect 1081 1172 1168 1179
rect 1193 1199 1230 1341
rect 1496 1340 1533 1341
rect 2241 1338 2657 1343
rect 2241 1337 2582 1338
rect 1898 1306 2008 1320
rect 1898 1303 1941 1306
rect 1898 1298 1902 1303
rect 1820 1276 1902 1298
rect 1931 1276 1941 1303
rect 1969 1279 1976 1306
rect 2005 1298 2008 1306
rect 2005 1279 2070 1298
rect 1969 1276 2070 1279
rect 1820 1274 2070 1276
rect 1345 1209 1381 1210
rect 1193 1179 1202 1199
rect 1222 1179 1230 1199
rect 1081 1170 1137 1172
rect 1081 1169 1118 1170
rect 1193 1169 1230 1179
rect 1289 1199 1437 1209
rect 1537 1206 1633 1208
rect 1289 1179 1298 1199
rect 1318 1179 1408 1199
rect 1428 1179 1437 1199
rect 1289 1173 1437 1179
rect 1289 1170 1353 1173
rect 1289 1169 1326 1170
rect 1345 1143 1353 1170
rect 1374 1170 1437 1173
rect 1495 1199 1633 1206
rect 1495 1179 1504 1199
rect 1524 1179 1633 1199
rect 1495 1170 1633 1179
rect 1820 1195 1857 1274
rect 1898 1261 2008 1274
rect 1972 1205 2003 1206
rect 1820 1175 1829 1195
rect 1849 1175 1857 1195
rect 1374 1143 1381 1170
rect 1400 1169 1437 1170
rect 1496 1169 1533 1170
rect 1345 1118 1381 1143
rect 816 1116 857 1117
rect 652 1109 857 1116
rect 652 1098 826 1109
rect 652 1065 660 1098
rect 653 1056 660 1065
rect 709 1089 826 1098
rect 846 1089 857 1109
rect 709 1081 857 1089
rect 924 1113 1283 1117
rect 924 1108 1246 1113
rect 924 1084 1037 1108
rect 1061 1089 1246 1108
rect 1270 1089 1283 1113
rect 1061 1084 1283 1089
rect 924 1081 1283 1084
rect 1345 1081 1380 1118
rect 1448 1115 1548 1118
rect 1448 1111 1515 1115
rect 1448 1085 1460 1111
rect 1486 1089 1515 1111
rect 1541 1089 1548 1115
rect 1486 1085 1548 1089
rect 1448 1081 1548 1085
rect 709 1065 720 1081
rect 709 1056 717 1065
rect 924 1060 955 1081
rect 1345 1060 1381 1081
rect 767 1059 804 1060
rect 432 1016 497 1035
rect 432 998 457 1016
rect 475 998 497 1016
rect 432 797 497 998
rect 653 872 717 1056
rect 766 1050 804 1059
rect 766 1030 775 1050
rect 795 1030 804 1050
rect 766 1022 804 1030
rect 870 1054 955 1060
rect 980 1059 1017 1060
rect 870 1034 878 1054
rect 898 1034 955 1054
rect 870 1026 955 1034
rect 979 1050 1017 1059
rect 979 1030 988 1050
rect 1008 1030 1017 1050
rect 870 1025 906 1026
rect 979 1022 1017 1030
rect 1083 1054 1168 1060
rect 1188 1059 1225 1060
rect 1083 1034 1091 1054
rect 1111 1053 1168 1054
rect 1111 1034 1140 1053
rect 1083 1033 1140 1034
rect 1161 1033 1168 1053
rect 1083 1026 1168 1033
rect 1187 1050 1225 1059
rect 1187 1030 1196 1050
rect 1216 1030 1225 1050
rect 1083 1025 1119 1026
rect 1187 1022 1225 1030
rect 1291 1054 1435 1060
rect 1291 1034 1299 1054
rect 1319 1034 1407 1054
rect 1427 1034 1435 1054
rect 1291 1026 1435 1034
rect 1291 1025 1327 1026
rect 1399 1025 1435 1026
rect 1501 1059 1538 1060
rect 1501 1058 1539 1059
rect 1501 1050 1565 1058
rect 1501 1030 1510 1050
rect 1530 1036 1565 1050
rect 1585 1036 1588 1056
rect 1530 1031 1588 1036
rect 1530 1030 1565 1031
rect 767 993 804 1022
rect 768 991 804 993
rect 980 991 1017 1022
rect 768 969 1017 991
rect 849 963 960 969
rect 849 955 890 963
rect 849 935 857 955
rect 876 935 890 955
rect 849 933 890 935
rect 918 955 960 963
rect 918 935 934 955
rect 953 935 960 955
rect 918 933 960 935
rect 849 918 960 933
rect 653 862 721 872
rect 653 829 670 862
rect 710 829 721 862
rect 653 817 721 829
rect 653 815 717 817
rect 1188 798 1225 1022
rect 1501 1018 1565 1030
rect 1605 800 1632 1170
rect 1820 1165 1857 1175
rect 1916 1195 2003 1205
rect 1916 1175 1925 1195
rect 1945 1175 2003 1195
rect 1916 1166 2003 1175
rect 1916 1165 1953 1166
rect 1696 1152 1766 1157
rect 1691 1146 1766 1152
rect 1691 1113 1699 1146
rect 1752 1113 1766 1146
rect 1972 1113 2003 1166
rect 2033 1195 2070 1274
rect 2185 1205 2216 1206
rect 2033 1175 2042 1195
rect 2062 1175 2070 1195
rect 2033 1165 2070 1175
rect 2129 1198 2216 1205
rect 2129 1195 2190 1198
rect 2129 1175 2138 1195
rect 2158 1178 2190 1195
rect 2211 1178 2216 1198
rect 2158 1175 2216 1178
rect 2129 1168 2216 1175
rect 2241 1195 2278 1337
rect 2544 1336 2581 1337
rect 2393 1205 2429 1206
rect 2241 1175 2250 1195
rect 2270 1175 2278 1195
rect 2129 1166 2185 1168
rect 2129 1165 2166 1166
rect 2241 1165 2278 1175
rect 2337 1195 2485 1205
rect 2585 1202 2681 1204
rect 2337 1175 2346 1195
rect 2366 1175 2456 1195
rect 2476 1175 2485 1195
rect 2337 1169 2485 1175
rect 2337 1166 2401 1169
rect 2337 1165 2374 1166
rect 2393 1139 2401 1166
rect 2422 1166 2485 1169
rect 2543 1195 2681 1202
rect 2543 1175 2552 1195
rect 2572 1175 2681 1195
rect 2543 1166 2681 1175
rect 2422 1139 2429 1166
rect 2448 1165 2485 1166
rect 2544 1165 2581 1166
rect 2393 1114 2429 1139
rect 1691 1112 1774 1113
rect 1864 1112 1905 1113
rect 1691 1105 1905 1112
rect 1691 1088 1874 1105
rect 1691 1055 1704 1088
rect 1757 1085 1874 1088
rect 1894 1085 1905 1105
rect 1757 1077 1905 1085
rect 1972 1109 2331 1113
rect 1972 1104 2294 1109
rect 1972 1080 2085 1104
rect 2109 1085 2294 1104
rect 2318 1085 2331 1109
rect 2109 1080 2331 1085
rect 1972 1077 2331 1080
rect 2393 1077 2428 1114
rect 2496 1111 2596 1114
rect 2496 1107 2563 1111
rect 2496 1081 2508 1107
rect 2534 1085 2563 1107
rect 2589 1085 2596 1111
rect 2534 1081 2596 1085
rect 2496 1077 2596 1081
rect 1757 1055 1774 1077
rect 1972 1056 2003 1077
rect 2393 1056 2429 1077
rect 1815 1055 1852 1056
rect 1691 1041 1774 1055
rect 1464 798 1632 800
rect 1188 797 1632 798
rect 432 767 1632 797
rect 1702 831 1774 1041
rect 1814 1046 1852 1055
rect 1814 1026 1823 1046
rect 1843 1026 1852 1046
rect 1814 1018 1852 1026
rect 1918 1050 2003 1056
rect 2028 1055 2065 1056
rect 1918 1030 1926 1050
rect 1946 1030 2003 1050
rect 1918 1022 2003 1030
rect 2027 1046 2065 1055
rect 2027 1026 2036 1046
rect 2056 1026 2065 1046
rect 1918 1021 1954 1022
rect 2027 1018 2065 1026
rect 2131 1050 2216 1056
rect 2236 1055 2273 1056
rect 2131 1030 2139 1050
rect 2159 1049 2216 1050
rect 2159 1030 2188 1049
rect 2131 1029 2188 1030
rect 2209 1029 2216 1049
rect 2131 1022 2216 1029
rect 2235 1046 2273 1055
rect 2235 1026 2244 1046
rect 2264 1026 2273 1046
rect 2131 1021 2167 1022
rect 2235 1018 2273 1026
rect 2339 1050 2483 1056
rect 2339 1030 2347 1050
rect 2367 1030 2455 1050
rect 2475 1030 2483 1050
rect 2339 1022 2483 1030
rect 2339 1021 2375 1022
rect 2447 1021 2483 1022
rect 2549 1055 2586 1056
rect 2549 1054 2587 1055
rect 2549 1046 2613 1054
rect 2549 1026 2558 1046
rect 2578 1032 2613 1046
rect 2633 1032 2636 1052
rect 2578 1027 2636 1032
rect 2578 1026 2613 1027
rect 1815 989 1852 1018
rect 1816 987 1852 989
rect 2028 987 2065 1018
rect 1816 965 2065 987
rect 1897 959 2008 965
rect 1897 951 1938 959
rect 1897 931 1905 951
rect 1924 931 1938 951
rect 1897 929 1938 931
rect 1966 951 2008 959
rect 1966 931 1982 951
rect 2001 931 2008 951
rect 1966 929 2008 931
rect 1897 914 2008 929
rect 1702 792 1721 831
rect 1766 792 1774 831
rect 1702 775 1774 792
rect 2236 819 2273 1018
rect 2549 1014 2613 1026
rect 2236 813 2277 819
rect 2653 815 2680 1166
rect 2512 813 2680 815
rect 2236 787 2680 813
rect 432 720 497 767
rect 432 702 455 720
rect 473 702 497 720
rect 1345 747 1380 749
rect 1345 745 1449 747
rect 2238 745 2277 787
rect 2512 786 2680 787
rect 1345 738 2279 745
rect 1345 737 1396 738
rect 1345 717 1348 737
rect 1373 718 1396 737
rect 1428 718 2279 738
rect 1373 717 2279 718
rect 1345 710 2279 717
rect 1618 709 2279 710
rect 432 681 497 702
rect 709 692 749 695
rect 709 688 1612 692
rect 709 668 1586 688
rect 1606 668 1612 688
rect 709 665 1612 668
rect 433 621 498 641
rect 433 603 457 621
rect 475 603 498 621
rect 433 576 498 603
rect 709 576 749 665
rect 1193 663 1609 665
rect 1193 662 1534 663
rect 850 631 960 645
rect 850 628 893 631
rect 850 623 854 628
rect 432 541 749 576
rect 772 601 854 623
rect 883 601 893 628
rect 921 604 928 631
rect 957 623 960 631
rect 957 604 1022 623
rect 921 601 1022 604
rect 772 599 1022 601
rect 433 465 498 541
rect 772 520 809 599
rect 850 586 960 599
rect 924 530 955 531
rect 772 500 781 520
rect 801 500 809 520
rect 772 490 809 500
rect 868 520 955 530
rect 868 500 877 520
rect 897 500 955 520
rect 868 491 955 500
rect 868 490 905 491
rect 433 447 455 465
rect 473 447 498 465
rect 433 426 498 447
rect 646 445 711 454
rect 646 408 656 445
rect 696 437 711 445
rect 924 438 955 491
rect 985 520 1022 599
rect 1137 530 1168 531
rect 985 500 994 520
rect 1014 500 1022 520
rect 985 490 1022 500
rect 1081 523 1168 530
rect 1081 520 1142 523
rect 1081 500 1090 520
rect 1110 503 1142 520
rect 1163 503 1168 523
rect 1110 500 1168 503
rect 1081 493 1168 500
rect 1193 520 1230 662
rect 1496 661 1533 662
rect 1345 530 1381 531
rect 1193 500 1202 520
rect 1222 500 1230 520
rect 1081 491 1137 493
rect 1081 490 1118 491
rect 1193 490 1230 500
rect 1289 520 1437 530
rect 1537 527 1633 529
rect 1289 500 1298 520
rect 1318 500 1408 520
rect 1428 500 1437 520
rect 1289 494 1437 500
rect 1289 491 1353 494
rect 1289 490 1326 491
rect 1345 464 1353 491
rect 1374 491 1437 494
rect 1495 520 1633 527
rect 1495 500 1504 520
rect 1524 500 1633 520
rect 1495 491 1633 500
rect 1374 464 1381 491
rect 1400 490 1437 491
rect 1496 490 1533 491
rect 1345 439 1381 464
rect 816 437 857 438
rect 696 430 857 437
rect 696 410 826 430
rect 846 410 857 430
rect 696 408 857 410
rect 646 402 857 408
rect 924 434 1283 438
rect 924 429 1246 434
rect 924 405 1037 429
rect 1061 410 1246 429
rect 1270 410 1283 434
rect 1061 405 1283 410
rect 924 402 1283 405
rect 1345 402 1380 439
rect 1448 436 1548 439
rect 1448 432 1515 436
rect 1448 406 1460 432
rect 1486 410 1515 432
rect 1541 410 1548 436
rect 1486 406 1548 410
rect 1448 402 1548 406
rect 646 389 713 402
rect 438 366 494 386
rect 438 348 457 366
rect 475 348 494 366
rect 438 235 494 348
rect 646 368 660 389
rect 696 368 713 389
rect 924 381 955 402
rect 1345 381 1381 402
rect 767 380 804 381
rect 646 361 713 368
rect 766 371 804 380
rect 438 94 493 235
rect 646 209 711 361
rect 766 351 775 371
rect 795 351 804 371
rect 766 343 804 351
rect 870 375 955 381
rect 980 380 1017 381
rect 870 355 878 375
rect 898 355 955 375
rect 870 347 955 355
rect 979 371 1017 380
rect 979 351 988 371
rect 1008 351 1017 371
rect 870 346 906 347
rect 979 343 1017 351
rect 1083 375 1168 381
rect 1188 380 1225 381
rect 1083 355 1091 375
rect 1111 374 1168 375
rect 1111 355 1140 374
rect 1083 354 1140 355
rect 1161 354 1168 374
rect 1083 347 1168 354
rect 1187 371 1225 380
rect 1187 351 1196 371
rect 1216 351 1225 371
rect 1083 346 1119 347
rect 1187 343 1225 351
rect 1291 375 1435 381
rect 1291 355 1299 375
rect 1319 355 1407 375
rect 1427 355 1435 375
rect 1291 347 1435 355
rect 1291 346 1327 347
rect 1399 346 1435 347
rect 1501 380 1538 381
rect 1501 379 1539 380
rect 1501 371 1565 379
rect 1501 351 1510 371
rect 1530 357 1565 371
rect 1585 357 1588 377
rect 1530 352 1588 357
rect 1530 351 1565 352
rect 767 314 804 343
rect 768 312 804 314
rect 980 312 1017 343
rect 768 290 1017 312
rect 849 284 960 290
rect 849 276 890 284
rect 849 256 857 276
rect 876 256 890 276
rect 849 254 890 256
rect 918 276 960 284
rect 918 256 934 276
rect 953 256 960 276
rect 918 254 960 256
rect 849 239 960 254
rect 1188 244 1225 343
rect 1501 339 1565 351
rect 639 199 760 209
rect 639 197 708 199
rect 639 156 652 197
rect 689 158 708 197
rect 745 158 760 199
rect 689 156 760 158
rect 639 138 760 156
rect 851 94 955 239
rect 1186 94 1227 244
rect 1605 236 1632 491
rect 1694 481 1774 492
rect 1694 455 1711 481
rect 1751 455 1774 481
rect 1694 428 1774 455
rect 1694 402 1715 428
rect 1755 402 1774 428
rect 1694 383 1774 402
rect 1694 357 1718 383
rect 1758 357 1774 383
rect 1694 306 1774 357
rect 438 91 1227 94
rect 1606 105 1632 236
rect 1606 91 1634 105
rect 438 58 1634 91
rect 440 56 1634 58
rect 851 54 955 56
rect 1186 54 1227 56
rect 1696 53 1766 306
<< viali >>
rect 1353 1406 1378 1441
rect 1397 1406 1422 1444
rect 1586 1347 1606 1367
rect 2403 1407 2428 1442
rect 2447 1407 2472 1445
rect 2634 1343 2654 1363
rect 854 1280 883 1307
rect 928 1283 957 1310
rect 659 1119 708 1161
rect 1142 1182 1163 1202
rect 1902 1276 1931 1303
rect 1976 1279 2005 1306
rect 1353 1143 1374 1173
rect 660 1056 709 1098
rect 1515 1089 1541 1115
rect 1140 1033 1161 1053
rect 1565 1036 1585 1056
rect 857 935 876 955
rect 934 935 953 955
rect 670 829 710 862
rect 1699 1113 1752 1146
rect 2190 1178 2211 1198
rect 2401 1139 2422 1169
rect 1704 1055 1757 1088
rect 2563 1085 2589 1111
rect 2188 1029 2209 1049
rect 2613 1032 2633 1052
rect 1905 931 1924 951
rect 1982 931 2001 951
rect 1721 792 1766 831
rect 1348 717 1373 737
rect 1396 718 1428 738
rect 1586 668 1606 688
rect 854 601 883 628
rect 928 604 957 631
rect 656 408 696 445
rect 1142 503 1163 523
rect 1353 464 1374 494
rect 1515 410 1541 436
rect 660 368 696 389
rect 1140 354 1161 374
rect 1565 357 1585 377
rect 857 256 876 276
rect 934 256 953 276
rect 652 156 689 197
rect 708 158 745 199
rect 1711 455 1751 481
rect 1715 402 1755 428
rect 1718 357 1758 383
<< metal1 >>
rect 3024 13745 3512 13777
rect 3024 13146 16418 13745
rect 171 973 278 1486
rect 650 1161 722 1477
rect 1346 1452 1418 1453
rect 1345 1444 1444 1452
rect 1345 1441 1397 1444
rect 1345 1406 1353 1441
rect 1378 1406 1397 1441
rect 1422 1406 1444 1444
rect 1345 1394 1444 1406
rect 1346 1375 1414 1394
rect 1347 1372 1380 1375
rect 1582 1372 1614 1373
rect 757 1311 960 1324
rect 757 1278 781 1311
rect 817 1310 960 1311
rect 817 1307 928 1310
rect 817 1280 854 1307
rect 883 1283 928 1307
rect 957 1283 960 1310
rect 883 1280 960 1283
rect 817 1278 960 1280
rect 757 1265 960 1278
rect 757 1264 858 1265
rect 650 1119 659 1161
rect 708 1119 722 1161
rect 650 1098 722 1119
rect 650 1056 660 1098
rect 709 1056 722 1098
rect 650 1038 722 1056
rect 1135 1202 1167 1209
rect 1135 1182 1142 1202
rect 1163 1182 1167 1202
rect 1135 1117 1167 1182
rect 1347 1173 1378 1372
rect 1579 1367 1614 1372
rect 1579 1347 1586 1367
rect 1606 1347 1614 1367
rect 1579 1339 1614 1347
rect 1347 1143 1353 1173
rect 1374 1143 1378 1173
rect 1347 1135 1378 1143
rect 1505 1117 1545 1118
rect 1135 1115 1547 1117
rect 1135 1089 1515 1115
rect 1541 1089 1547 1115
rect 1135 1081 1547 1089
rect 1135 1053 1167 1081
rect 1580 1061 1614 1339
rect 1696 1152 1766 1525
rect 2396 1453 2468 1454
rect 2395 1450 2494 1453
rect 3024 1450 16383 13146
rect 2395 1445 16383 1450
rect 2395 1442 2447 1445
rect 2395 1407 2403 1442
rect 2428 1407 2447 1442
rect 2472 1407 16383 1445
rect 2395 1395 16383 1407
rect 2395 1394 2464 1395
rect 2395 1376 2431 1394
rect 1805 1307 2008 1320
rect 1805 1274 1829 1307
rect 1865 1306 2008 1307
rect 1865 1303 1976 1306
rect 1865 1276 1902 1303
rect 1931 1279 1976 1303
rect 2005 1279 2008 1306
rect 1931 1276 2008 1279
rect 1865 1274 2008 1276
rect 1805 1261 2008 1274
rect 1805 1260 1906 1261
rect 1135 1033 1140 1053
rect 1161 1033 1167 1053
rect 1135 1026 1167 1033
rect 1558 1056 1614 1061
rect 1558 1036 1565 1056
rect 1585 1036 1614 1056
rect 1691 1146 1766 1152
rect 1691 1113 1699 1146
rect 1752 1113 1766 1146
rect 1691 1088 1766 1113
rect 1691 1055 1704 1088
rect 1757 1055 1766 1088
rect 1691 1046 1766 1055
rect 2183 1198 2215 1205
rect 2183 1178 2190 1198
rect 2211 1178 2215 1198
rect 2183 1113 2215 1178
rect 2395 1169 2426 1376
rect 2630 1368 2662 1369
rect 2627 1363 2662 1368
rect 2627 1343 2634 1363
rect 2654 1343 2662 1363
rect 2627 1335 2662 1343
rect 2395 1139 2401 1169
rect 2422 1139 2426 1169
rect 2395 1131 2426 1139
rect 2553 1113 2593 1114
rect 2183 1111 2595 1113
rect 2183 1085 2563 1111
rect 2589 1085 2595 1111
rect 2183 1077 2595 1085
rect 2183 1049 2215 1077
rect 2628 1057 2662 1335
rect 1691 1041 1749 1046
rect 1558 1029 1614 1036
rect 2183 1029 2188 1049
rect 2209 1029 2215 1049
rect 1558 1028 1593 1029
rect 2183 1022 2215 1029
rect 2606 1052 2662 1057
rect 2606 1032 2613 1052
rect 2633 1032 2662 1052
rect 2606 1025 2662 1032
rect 2606 1024 2641 1025
rect 849 973 960 977
rect 171 955 2847 973
rect 171 935 857 955
rect 876 935 934 955
rect 953 951 2847 955
rect 953 935 1905 951
rect 171 931 1905 935
rect 1924 931 1982 951
rect 2001 931 2847 951
rect 171 917 2847 931
rect 171 294 278 917
rect 1897 914 2008 917
rect 657 868 721 872
rect 653 862 721 868
rect 653 829 670 862
rect 710 829 721 862
rect 653 817 721 829
rect 1704 831 1769 853
rect 653 815 710 817
rect 657 454 708 815
rect 1704 792 1721 831
rect 1766 792 1769 831
rect 1345 747 1380 749
rect 1345 738 1449 747
rect 1345 737 1396 738
rect 1345 717 1348 737
rect 1373 718 1396 737
rect 1428 718 1449 738
rect 1373 717 1449 718
rect 1345 710 1449 717
rect 1345 698 1380 710
rect 757 632 960 645
rect 757 599 781 632
rect 817 631 960 632
rect 817 628 928 631
rect 817 601 854 628
rect 883 604 928 628
rect 957 604 960 631
rect 883 601 960 604
rect 817 599 960 601
rect 757 586 960 599
rect 757 585 858 586
rect 1135 523 1167 530
rect 1135 503 1142 523
rect 1163 503 1167 523
rect 646 445 711 454
rect 646 408 656 445
rect 696 411 711 445
rect 1135 438 1167 503
rect 1347 494 1378 698
rect 1582 693 1614 694
rect 1579 688 1614 693
rect 1579 668 1586 688
rect 1606 668 1614 688
rect 1579 660 1614 668
rect 1347 464 1353 494
rect 1374 464 1378 494
rect 1347 456 1378 464
rect 1505 438 1545 439
rect 1135 436 1547 438
rect 696 408 713 411
rect 646 389 713 408
rect 646 368 660 389
rect 696 368 713 389
rect 646 361 713 368
rect 1135 410 1515 436
rect 1541 410 1547 436
rect 1135 402 1547 410
rect 1135 374 1167 402
rect 1580 382 1614 660
rect 1704 492 1769 792
rect 1135 354 1140 374
rect 1161 354 1167 374
rect 1135 347 1167 354
rect 1558 377 1614 382
rect 1558 357 1565 377
rect 1585 357 1614 377
rect 1558 350 1614 357
rect 1694 481 1774 492
rect 1694 455 1711 481
rect 1751 455 1774 481
rect 1694 428 1774 455
rect 1694 402 1715 428
rect 1755 402 1774 428
rect 1694 383 1774 402
rect 1694 357 1718 383
rect 1758 357 1774 383
rect 1558 349 1593 350
rect 1694 345 1774 357
rect 849 294 960 298
rect 2604 294 2839 295
rect 169 276 2839 294
rect 169 256 857 276
rect 876 256 934 276
rect 953 256 2839 276
rect 169 238 2839 256
rect 171 38 278 238
rect 639 199 760 209
rect 639 197 708 199
rect 639 156 652 197
rect 689 158 708 197
rect 745 158 760 199
rect 689 156 760 158
rect 639 138 760 156
rect 3024 165 16383 1395
rect 645 0 710 138
rect 3024 102 3544 165
rect 15863 102 16383 165
<< via1 >>
rect 781 1278 817 1311
rect 1829 1274 1865 1307
rect 781 599 817 632
<< metal2 >>
rect 0 1326 107 1483
rect 0 1311 2879 1326
rect 0 1278 781 1311
rect 817 1307 2879 1311
rect 817 1278 1829 1307
rect 0 1274 1829 1278
rect 1865 1274 2879 1307
rect 0 1257 2879 1274
rect 0 651 107 1257
rect 0 632 2887 651
rect 0 599 781 632
rect 817 599 2887 632
rect 0 582 2887 599
rect 0 36 107 582
<< metal3 >>
rect 3024 13745 3512 13777
rect 3024 13146 16418 13745
rect 3024 165 16383 13146
rect 3024 102 3544 165
rect 15863 102 16383 165
<< mimcap >>
rect 3748 886 15811 13034
<< labels >>
rlabel metal1 2486 1404 2494 1444 1 vout
rlabel locali 443 1434 487 1456 1 vref
rlabel metal1 179 1423 275 1456 1 gnd
rlabel metal2 3 1423 99 1456 1 vdd
rlabel metal1 658 1438 720 1465 1 d0
rlabel metal1 1704 1467 1757 1489 1 d1
<< end >>
