magic
tech sky130A
timestamp 1620547697
<< nwell >>
rect 41 351 368 425
rect 41 201 852 351
rect 979 107 1306 181
rect 979 -43 1790 107
rect 40 -203 367 -129
rect 40 -353 851 -203
<< nmos >>
rect 105 100 155 142
rect 318 100 368 142
rect 526 100 576 142
rect 734 100 784 142
rect 1043 -144 1093 -102
rect 1256 -144 1306 -102
rect 1464 -144 1514 -102
rect 1672 -144 1722 -102
rect 104 -454 154 -412
rect 317 -454 367 -412
rect 525 -454 575 -412
rect 733 -454 783 -412
<< pmos >>
rect 105 219 155 319
rect 318 219 368 319
rect 526 219 576 319
rect 734 219 784 319
rect 1043 -25 1093 75
rect 1256 -25 1306 75
rect 1464 -25 1514 75
rect 1672 -25 1722 75
rect 104 -335 154 -235
rect 317 -335 367 -235
rect 525 -335 575 -235
rect 733 -335 783 -235
<< ndiff >>
rect 56 132 105 142
rect 56 112 67 132
rect 87 112 105 132
rect 56 100 105 112
rect 155 136 199 142
rect 155 116 170 136
rect 190 116 199 136
rect 155 100 199 116
rect 269 132 318 142
rect 269 112 280 132
rect 300 112 318 132
rect 269 100 318 112
rect 368 136 412 142
rect 368 116 383 136
rect 403 116 412 136
rect 368 100 412 116
rect 477 132 526 142
rect 477 112 488 132
rect 508 112 526 132
rect 477 100 526 112
rect 576 136 620 142
rect 576 116 591 136
rect 611 116 620 136
rect 576 100 620 116
rect 690 136 734 142
rect 690 116 699 136
rect 719 116 734 136
rect 690 100 734 116
rect 784 132 833 142
rect 784 112 802 132
rect 822 112 833 132
rect 784 100 833 112
rect 994 -112 1043 -102
rect 994 -132 1005 -112
rect 1025 -132 1043 -112
rect 994 -144 1043 -132
rect 1093 -108 1137 -102
rect 1093 -128 1108 -108
rect 1128 -128 1137 -108
rect 1093 -144 1137 -128
rect 1207 -112 1256 -102
rect 1207 -132 1218 -112
rect 1238 -132 1256 -112
rect 1207 -144 1256 -132
rect 1306 -108 1350 -102
rect 1306 -128 1321 -108
rect 1341 -128 1350 -108
rect 1306 -144 1350 -128
rect 1415 -112 1464 -102
rect 1415 -132 1426 -112
rect 1446 -132 1464 -112
rect 1415 -144 1464 -132
rect 1514 -108 1558 -102
rect 1514 -128 1529 -108
rect 1549 -128 1558 -108
rect 1514 -144 1558 -128
rect 1628 -108 1672 -102
rect 1628 -128 1637 -108
rect 1657 -128 1672 -108
rect 1628 -144 1672 -128
rect 1722 -112 1771 -102
rect 1722 -132 1740 -112
rect 1760 -132 1771 -112
rect 1722 -144 1771 -132
rect 55 -422 104 -412
rect 55 -442 66 -422
rect 86 -442 104 -422
rect 55 -454 104 -442
rect 154 -418 198 -412
rect 154 -438 169 -418
rect 189 -438 198 -418
rect 154 -454 198 -438
rect 268 -422 317 -412
rect 268 -442 279 -422
rect 299 -442 317 -422
rect 268 -454 317 -442
rect 367 -418 411 -412
rect 367 -438 382 -418
rect 402 -438 411 -418
rect 367 -454 411 -438
rect 476 -422 525 -412
rect 476 -442 487 -422
rect 507 -442 525 -422
rect 476 -454 525 -442
rect 575 -418 619 -412
rect 575 -438 590 -418
rect 610 -438 619 -418
rect 575 -454 619 -438
rect 689 -418 733 -412
rect 689 -438 698 -418
rect 718 -438 733 -418
rect 689 -454 733 -438
rect 783 -422 832 -412
rect 783 -442 801 -422
rect 821 -442 832 -422
rect 783 -454 832 -442
<< pdiff >>
rect 61 281 105 319
rect 61 261 73 281
rect 93 261 105 281
rect 61 219 105 261
rect 155 281 197 319
rect 155 261 169 281
rect 189 261 197 281
rect 155 219 197 261
rect 274 281 318 319
rect 274 261 286 281
rect 306 261 318 281
rect 274 219 318 261
rect 368 281 410 319
rect 368 261 382 281
rect 402 261 410 281
rect 368 219 410 261
rect 482 281 526 319
rect 482 261 494 281
rect 514 261 526 281
rect 482 219 526 261
rect 576 281 618 319
rect 576 261 590 281
rect 610 261 618 281
rect 576 219 618 261
rect 692 281 734 319
rect 692 261 700 281
rect 720 261 734 281
rect 692 219 734 261
rect 784 288 829 319
rect 784 281 828 288
rect 784 261 796 281
rect 816 261 828 281
rect 784 219 828 261
rect 999 37 1043 75
rect 999 17 1011 37
rect 1031 17 1043 37
rect 999 -25 1043 17
rect 1093 37 1135 75
rect 1093 17 1107 37
rect 1127 17 1135 37
rect 1093 -25 1135 17
rect 1212 37 1256 75
rect 1212 17 1224 37
rect 1244 17 1256 37
rect 1212 -25 1256 17
rect 1306 37 1348 75
rect 1306 17 1320 37
rect 1340 17 1348 37
rect 1306 -25 1348 17
rect 1420 37 1464 75
rect 1420 17 1432 37
rect 1452 17 1464 37
rect 1420 -25 1464 17
rect 1514 37 1556 75
rect 1514 17 1528 37
rect 1548 17 1556 37
rect 1514 -25 1556 17
rect 1630 37 1672 75
rect 1630 17 1638 37
rect 1658 17 1672 37
rect 1630 -25 1672 17
rect 1722 44 1767 75
rect 1722 37 1766 44
rect 1722 17 1734 37
rect 1754 17 1766 37
rect 1722 -25 1766 17
rect 60 -273 104 -235
rect 60 -293 72 -273
rect 92 -293 104 -273
rect 60 -335 104 -293
rect 154 -273 196 -235
rect 154 -293 168 -273
rect 188 -293 196 -273
rect 154 -335 196 -293
rect 273 -273 317 -235
rect 273 -293 285 -273
rect 305 -293 317 -273
rect 273 -335 317 -293
rect 367 -273 409 -235
rect 367 -293 381 -273
rect 401 -293 409 -273
rect 367 -335 409 -293
rect 481 -273 525 -235
rect 481 -293 493 -273
rect 513 -293 525 -273
rect 481 -335 525 -293
rect 575 -273 617 -235
rect 575 -293 589 -273
rect 609 -293 617 -273
rect 575 -335 617 -293
rect 691 -273 733 -235
rect 691 -293 699 -273
rect 719 -293 733 -273
rect 691 -335 733 -293
rect 783 -266 828 -235
rect 783 -273 827 -266
rect 783 -293 795 -273
rect 815 -293 827 -273
rect 783 -335 827 -293
<< ndiffc >>
rect -161 397 -143 415
rect -159 298 -141 316
rect -161 210 -143 228
rect -159 111 -141 129
rect 67 112 87 132
rect 170 116 190 136
rect 280 112 300 132
rect 383 116 403 136
rect 488 112 508 132
rect 591 116 611 136
rect 699 116 719 136
rect 802 112 822 132
rect -161 -19 -143 -1
rect -159 -118 -141 -100
rect 1005 -132 1025 -112
rect 1108 -128 1128 -108
rect 1218 -132 1238 -112
rect 1321 -128 1341 -108
rect 1426 -132 1446 -112
rect 1529 -128 1549 -108
rect 1637 -128 1657 -108
rect 1740 -132 1760 -112
rect -161 -249 -143 -231
rect -159 -348 -141 -330
rect 66 -442 86 -422
rect 169 -438 189 -418
rect 279 -442 299 -422
rect 382 -438 402 -418
rect 487 -442 507 -422
rect 590 -438 610 -418
rect 698 -438 718 -418
rect 801 -442 821 -422
<< pdiffc >>
rect 73 261 93 281
rect 169 261 189 281
rect 286 261 306 281
rect 382 261 402 281
rect 494 261 514 281
rect 590 261 610 281
rect 700 261 720 281
rect 796 261 816 281
rect 1011 17 1031 37
rect 1107 17 1127 37
rect 1224 17 1244 37
rect 1320 17 1340 37
rect 1432 17 1452 37
rect 1528 17 1548 37
rect 1638 17 1658 37
rect 1734 17 1754 37
rect 72 -293 92 -273
rect 168 -293 188 -273
rect 285 -293 305 -273
rect 381 -293 401 -273
rect 493 -293 513 -273
rect 589 -293 609 -273
rect 699 -293 719 -273
rect 795 -293 815 -273
<< psubdiff >>
rect 141 45 252 59
rect 141 15 182 45
rect 210 15 252 45
rect 141 0 252 15
rect 1079 -199 1190 -185
rect 1079 -229 1120 -199
rect 1148 -229 1190 -199
rect 1079 -244 1190 -229
rect 140 -509 251 -495
rect 140 -539 181 -509
rect 209 -539 251 -509
rect 140 -554 251 -539
<< nsubdiff >>
rect 142 392 252 406
rect 142 362 185 392
rect 213 362 252 392
rect 142 347 252 362
rect 1080 148 1190 162
rect 1080 118 1123 148
rect 1151 118 1190 148
rect 1080 103 1190 118
rect 141 -162 251 -148
rect 141 -192 184 -162
rect 212 -192 251 -162
rect 141 -207 251 -192
<< psubdiffcont >>
rect 182 15 210 45
rect 1120 -229 1148 -199
rect 181 -539 209 -509
<< nsubdiffcont >>
rect 185 362 213 392
rect 1123 118 1151 148
rect 184 -192 212 -162
<< poly >>
rect 105 319 155 332
rect 318 319 368 332
rect 526 319 576 332
rect 734 319 784 332
rect 105 191 155 219
rect 105 171 118 191
rect 138 171 155 191
rect 105 142 155 171
rect 318 190 368 219
rect 318 166 329 190
rect 353 166 368 190
rect 318 142 368 166
rect 526 195 576 219
rect 526 171 538 195
rect 562 171 576 195
rect 526 142 576 171
rect 734 193 784 219
rect 734 167 752 193
rect 778 167 784 193
rect 734 142 784 167
rect 105 84 155 100
rect 318 84 368 100
rect 526 84 576 100
rect 734 84 784 100
rect 1043 75 1093 88
rect 1256 75 1306 88
rect 1464 75 1514 88
rect 1672 75 1722 88
rect 1043 -53 1093 -25
rect 1043 -73 1056 -53
rect 1076 -73 1093 -53
rect 1043 -102 1093 -73
rect 1256 -54 1306 -25
rect 1256 -78 1267 -54
rect 1291 -78 1306 -54
rect 1256 -102 1306 -78
rect 1464 -49 1514 -25
rect 1464 -73 1476 -49
rect 1500 -73 1514 -49
rect 1464 -102 1514 -73
rect 1672 -51 1722 -25
rect 1672 -77 1690 -51
rect 1716 -77 1722 -51
rect 1672 -102 1722 -77
rect 1043 -160 1093 -144
rect 1256 -160 1306 -144
rect 1464 -160 1514 -144
rect 1672 -160 1722 -144
rect 104 -235 154 -222
rect 317 -235 367 -222
rect 525 -235 575 -222
rect 733 -235 783 -222
rect 104 -363 154 -335
rect 104 -383 117 -363
rect 137 -383 154 -363
rect 104 -412 154 -383
rect 317 -364 367 -335
rect 317 -388 328 -364
rect 352 -388 367 -364
rect 317 -412 367 -388
rect 525 -359 575 -335
rect 525 -383 537 -359
rect 561 -383 575 -359
rect 525 -412 575 -383
rect 733 -361 783 -335
rect 733 -387 751 -361
rect 777 -387 783 -361
rect 733 -412 783 -387
rect 104 -470 154 -454
rect 317 -470 367 -454
rect 525 -470 575 -454
rect 733 -470 783 -454
<< polycont >>
rect 118 171 138 191
rect 329 166 353 190
rect 538 171 562 195
rect 752 167 778 193
rect 1056 -73 1076 -53
rect 1267 -78 1291 -54
rect 1476 -73 1500 -49
rect 1690 -77 1716 -51
rect 117 -383 137 -363
rect 328 -388 352 -364
rect 537 -383 561 -359
rect 751 -387 777 -361
<< ndiffres >>
rect -182 415 -125 434
rect -182 412 -161 415
rect -276 397 -161 412
rect -143 397 -125 415
rect -276 374 -125 397
rect -276 338 -234 374
rect -277 337 -177 338
rect -277 316 -121 337
rect -277 298 -159 316
rect -141 298 -121 316
rect -277 294 -121 298
rect -182 278 -121 294
rect -182 228 -125 247
rect -182 225 -161 228
rect -276 210 -161 225
rect -143 210 -125 228
rect -276 187 -125 210
rect -276 151 -234 187
rect -277 150 -177 151
rect -277 129 -121 150
rect -277 111 -159 129
rect -141 111 -121 129
rect -277 107 -121 111
rect -182 91 -121 107
rect -182 -1 -125 18
rect -182 -4 -161 -1
rect -276 -19 -161 -4
rect -143 -19 -125 -1
rect -276 -42 -125 -19
rect -276 -78 -234 -42
rect -277 -79 -177 -78
rect -277 -100 -121 -79
rect -277 -118 -159 -100
rect -141 -118 -121 -100
rect -277 -122 -121 -118
rect -182 -138 -121 -122
rect -182 -231 -125 -212
rect -182 -234 -161 -231
rect -276 -249 -161 -234
rect -143 -249 -125 -231
rect -276 -272 -125 -249
rect -276 -308 -234 -272
rect -277 -309 -177 -308
rect -277 -330 -121 -309
rect -277 -348 -159 -330
rect -141 -348 -121 -330
rect -277 -352 -121 -348
rect -182 -368 -121 -352
<< locali >>
rect -172 417 -133 474
rect -172 415 -124 417
rect -172 397 -161 415
rect -143 397 -124 415
rect -172 388 -124 397
rect -171 387 -124 388
rect 142 392 252 406
rect 142 389 185 392
rect 142 384 146 389
rect 64 362 146 384
rect 175 362 185 389
rect 213 365 220 392
rect 249 384 252 392
rect 249 365 314 384
rect 213 362 314 365
rect 64 360 314 362
rect -168 324 -131 325
rect -172 321 -131 324
rect -172 316 -130 321
rect -172 298 -159 316
rect -141 298 -130 316
rect -172 284 -130 298
rect -92 284 -45 288
rect -172 278 -45 284
rect -172 249 -84 278
rect -55 249 -45 278
rect 64 281 101 360
rect 142 347 252 360
rect 216 291 247 292
rect 64 261 73 281
rect 93 261 101 281
rect 64 251 101 261
rect 160 281 247 291
rect 160 261 169 281
rect 189 261 247 281
rect 160 252 247 261
rect 160 251 197 252
rect -172 245 -45 249
rect -172 228 -133 245
rect -92 244 -45 245
rect -172 210 -161 228
rect -143 210 -133 228
rect -172 201 -133 210
rect -171 200 -134 201
rect 216 199 247 252
rect 277 281 314 360
rect 485 357 878 377
rect 898 357 901 377
rect 485 352 901 357
rect 485 351 826 352
rect 429 291 460 292
rect 277 261 286 281
rect 306 261 314 281
rect 277 251 314 261
rect 373 284 460 291
rect 373 281 434 284
rect 373 261 382 281
rect 402 264 434 281
rect 455 264 460 284
rect 402 261 460 264
rect 373 254 460 261
rect 485 281 522 351
rect 788 350 825 351
rect 637 291 673 292
rect 485 261 494 281
rect 514 261 522 281
rect 373 252 429 254
rect 373 251 410 252
rect 485 251 522 261
rect 581 281 729 291
rect 829 288 925 290
rect 581 261 590 281
rect 610 261 700 281
rect 720 261 729 281
rect 581 252 729 261
rect 787 281 925 288
rect 787 261 796 281
rect 816 261 925 281
rect 787 252 925 261
rect 581 251 618 252
rect 637 200 673 252
rect 692 251 729 252
rect 788 251 825 252
rect 108 198 149 199
rect 0 191 149 198
rect 0 171 118 191
rect 138 171 149 191
rect 0 163 149 171
rect 216 195 575 199
rect 216 190 538 195
rect 216 166 329 190
rect 353 171 538 190
rect 562 171 575 195
rect 353 166 575 171
rect 216 163 575 166
rect 637 163 672 200
rect 740 197 840 200
rect 740 193 807 197
rect 740 167 752 193
rect 778 171 807 193
rect 833 171 840 197
rect 778 167 840 171
rect 740 163 840 167
rect 216 142 247 163
rect 637 142 673 163
rect 59 141 96 142
rect -167 138 -133 139
rect -168 129 -131 138
rect -168 111 -159 129
rect -141 111 -131 129
rect -168 101 -131 111
rect 58 132 96 141
rect 58 112 67 132
rect 87 112 96 132
rect 58 104 96 112
rect 162 136 247 142
rect 272 141 309 142
rect 162 116 170 136
rect 190 116 247 136
rect 162 108 247 116
rect 271 132 309 141
rect 271 112 280 132
rect 300 112 309 132
rect 162 107 198 108
rect 271 104 309 112
rect 375 136 460 142
rect 480 141 517 142
rect 375 116 383 136
rect 403 135 460 136
rect 403 116 432 135
rect 375 115 432 116
rect 453 115 460 135
rect 375 108 460 115
rect 479 132 517 141
rect 479 112 488 132
rect 508 112 517 132
rect 375 107 411 108
rect 479 104 517 112
rect 583 136 727 142
rect 583 116 591 136
rect 611 135 699 136
rect 611 116 642 135
rect 583 115 642 116
rect 667 116 699 135
rect 719 116 727 136
rect 667 115 727 116
rect 583 108 727 115
rect 583 107 619 108
rect 691 107 727 108
rect 793 141 830 142
rect 793 140 831 141
rect 793 132 857 140
rect 793 112 802 132
rect 822 118 857 132
rect 877 118 880 138
rect 822 113 880 118
rect 822 112 857 113
rect -167 73 -133 101
rect 59 75 96 104
rect 60 73 96 75
rect 272 73 309 104
rect -167 72 5 73
rect -167 40 19 72
rect 60 51 309 73
rect 480 72 517 104
rect 793 100 857 112
rect 897 74 924 252
rect 1080 148 1190 162
rect 1080 145 1123 148
rect 1080 140 1084 145
rect 756 72 924 74
rect 480 66 924 72
rect -167 8 -133 40
rect -171 -1 -133 8
rect -171 -19 -161 -1
rect -143 -19 -133 -1
rect -171 -25 -133 -19
rect -15 -23 19 40
rect 141 45 252 51
rect 141 37 182 45
rect 141 17 149 37
rect 168 17 182 37
rect 141 15 182 17
rect 210 37 252 45
rect 210 17 226 37
rect 245 17 252 37
rect 210 15 252 17
rect 141 0 252 15
rect 479 46 924 66
rect 479 -23 517 46
rect 756 45 924 46
rect 1002 118 1084 140
rect 1113 118 1123 145
rect 1151 121 1158 148
rect 1187 140 1190 148
rect 1187 121 1252 140
rect 1151 118 1252 121
rect 1002 116 1252 118
rect 1002 37 1039 116
rect 1080 103 1190 116
rect 1154 47 1185 48
rect 1002 17 1011 37
rect 1031 17 1039 37
rect 1002 7 1039 17
rect 1098 37 1185 47
rect 1098 17 1107 37
rect 1127 17 1185 37
rect 1098 8 1185 17
rect 1098 7 1135 8
rect -171 -29 -134 -25
rect -15 -34 517 -23
rect -16 -50 517 -34
rect 1154 -45 1185 8
rect 1215 37 1252 116
rect 1423 113 1816 133
rect 1836 113 1839 133
rect 1423 108 1839 113
rect 1423 107 1764 108
rect 1367 47 1398 48
rect 1215 17 1224 37
rect 1244 17 1252 37
rect 1215 7 1252 17
rect 1311 40 1398 47
rect 1311 37 1372 40
rect 1311 17 1320 37
rect 1340 20 1372 37
rect 1393 20 1398 40
rect 1340 17 1398 20
rect 1311 10 1398 17
rect 1423 37 1460 107
rect 1726 106 1763 107
rect 1575 47 1611 48
rect 1423 17 1432 37
rect 1452 17 1460 37
rect 1311 8 1367 10
rect 1311 7 1348 8
rect 1423 7 1460 17
rect 1519 37 1667 47
rect 1767 44 1863 46
rect 1519 17 1528 37
rect 1548 17 1638 37
rect 1658 17 1667 37
rect 1519 8 1667 17
rect 1725 37 1863 44
rect 1725 17 1734 37
rect 1754 17 1863 37
rect 1725 8 1863 17
rect 1519 7 1556 8
rect 1575 -44 1611 8
rect 1630 7 1667 8
rect 1726 7 1763 8
rect 1046 -46 1087 -45
rect -16 -51 498 -50
rect 938 -53 1087 -46
rect 938 -73 1056 -53
rect 1076 -73 1087 -53
rect 938 -81 1087 -73
rect 1154 -49 1513 -45
rect 1154 -54 1476 -49
rect 1154 -78 1267 -54
rect 1291 -73 1476 -54
rect 1500 -73 1513 -49
rect 1291 -78 1513 -73
rect 1154 -81 1513 -78
rect 1575 -81 1610 -44
rect 1678 -47 1778 -44
rect 1678 -51 1745 -47
rect 1678 -77 1690 -51
rect 1716 -73 1745 -51
rect 1771 -73 1778 -47
rect 1716 -77 1778 -73
rect 1678 -81 1778 -77
rect -168 -92 -131 -91
rect -170 -100 -130 -92
rect -170 -118 -159 -100
rect -141 -118 -130 -100
rect 1154 -102 1185 -81
rect 1575 -102 1611 -81
rect 997 -103 1034 -102
rect -170 -166 -130 -118
rect 996 -112 1034 -103
rect 996 -132 1005 -112
rect 1025 -132 1034 -112
rect 996 -140 1034 -132
rect 1100 -108 1185 -102
rect 1210 -103 1247 -102
rect 1100 -128 1108 -108
rect 1128 -128 1185 -108
rect 1100 -136 1185 -128
rect 1209 -112 1247 -103
rect 1209 -132 1218 -112
rect 1238 -132 1247 -112
rect 1100 -137 1136 -136
rect 1209 -140 1247 -132
rect 1313 -108 1398 -102
rect 1418 -103 1455 -102
rect 1313 -128 1321 -108
rect 1341 -109 1398 -108
rect 1341 -128 1370 -109
rect 1313 -129 1370 -128
rect 1391 -129 1398 -109
rect 1313 -136 1398 -129
rect 1417 -112 1455 -103
rect 1417 -132 1426 -112
rect 1446 -132 1455 -112
rect 1313 -137 1349 -136
rect 1417 -140 1455 -132
rect 1521 -108 1665 -102
rect 1521 -128 1529 -108
rect 1549 -128 1637 -108
rect 1657 -128 1665 -108
rect 1521 -136 1665 -128
rect 1521 -137 1557 -136
rect 1629 -137 1665 -136
rect 1731 -103 1768 -102
rect 1731 -104 1769 -103
rect 1731 -112 1795 -104
rect 1731 -132 1740 -112
rect 1760 -126 1795 -112
rect 1815 -126 1818 -106
rect 1760 -131 1818 -126
rect 1760 -132 1795 -131
rect 141 -162 251 -148
rect 141 -165 184 -162
rect -170 -173 -45 -166
rect 141 -170 145 -165
rect -170 -192 -78 -173
rect -53 -192 -45 -173
rect -170 -202 -45 -192
rect 63 -192 145 -170
rect 174 -192 184 -165
rect 212 -189 219 -162
rect 248 -170 251 -162
rect 997 -169 1034 -140
rect 248 -189 313 -170
rect 998 -171 1034 -169
rect 1210 -171 1247 -140
rect 1418 -167 1455 -140
rect 1731 -144 1795 -132
rect 212 -192 313 -189
rect 63 -194 313 -192
rect -170 -222 -130 -202
rect -171 -231 -130 -222
rect -171 -249 -161 -231
rect -143 -249 -130 -231
rect -171 -258 -130 -249
rect -171 -259 -134 -258
rect 63 -273 100 -194
rect 141 -207 251 -194
rect 215 -263 246 -262
rect 63 -293 72 -273
rect 92 -293 100 -273
rect 63 -303 100 -293
rect 159 -273 246 -263
rect 159 -293 168 -273
rect 188 -293 246 -273
rect 159 -302 246 -293
rect 159 -303 196 -302
rect -168 -325 -131 -321
rect -171 -330 -131 -325
rect -171 -348 -159 -330
rect -141 -348 -131 -330
rect -171 -528 -131 -348
rect 215 -355 246 -302
rect 276 -273 313 -194
rect 484 -197 877 -177
rect 897 -197 900 -177
rect 998 -193 1247 -171
rect 1416 -172 1457 -167
rect 1835 -170 1862 8
rect 1694 -172 1862 -170
rect 1416 -178 1862 -172
rect 484 -202 900 -197
rect 1079 -199 1190 -193
rect 484 -203 825 -202
rect 428 -263 459 -262
rect 276 -293 285 -273
rect 305 -293 313 -273
rect 276 -303 313 -293
rect 372 -270 459 -263
rect 372 -273 433 -270
rect 372 -293 381 -273
rect 401 -290 433 -273
rect 454 -290 459 -270
rect 401 -293 459 -290
rect 372 -300 459 -293
rect 484 -273 521 -203
rect 787 -204 824 -203
rect 1079 -207 1120 -199
rect 1079 -227 1087 -207
rect 1106 -227 1120 -207
rect 1079 -229 1120 -227
rect 1148 -207 1190 -199
rect 1148 -227 1164 -207
rect 1183 -227 1190 -207
rect 1416 -200 1422 -178
rect 1448 -198 1862 -178
rect 1448 -200 1457 -198
rect 1694 -199 1862 -198
rect 1416 -209 1457 -200
rect 1148 -229 1190 -227
rect 1079 -244 1190 -229
rect 636 -263 672 -262
rect 484 -293 493 -273
rect 513 -293 521 -273
rect 372 -302 428 -300
rect 372 -303 409 -302
rect 484 -303 521 -293
rect 580 -273 728 -263
rect 828 -266 924 -264
rect 580 -293 589 -273
rect 609 -293 699 -273
rect 719 -293 728 -273
rect 580 -302 728 -293
rect 786 -273 924 -266
rect 786 -293 795 -273
rect 815 -293 924 -273
rect 786 -302 924 -293
rect 580 -303 617 -302
rect 636 -354 672 -302
rect 691 -303 728 -302
rect 787 -303 824 -302
rect 107 -356 148 -355
rect -1 -363 148 -356
rect -1 -383 117 -363
rect 137 -383 148 -363
rect -1 -391 148 -383
rect 215 -359 574 -355
rect 215 -364 537 -359
rect 215 -388 328 -364
rect 352 -383 537 -364
rect 561 -383 574 -359
rect 352 -388 574 -383
rect 215 -391 574 -388
rect 636 -391 671 -354
rect 739 -357 839 -354
rect 739 -361 806 -357
rect 739 -387 751 -361
rect 777 -383 806 -361
rect 832 -383 839 -357
rect 777 -387 839 -383
rect 739 -391 839 -387
rect 215 -412 246 -391
rect 636 -412 672 -391
rect 58 -413 95 -412
rect 57 -422 95 -413
rect 57 -442 66 -422
rect 86 -442 95 -422
rect 57 -450 95 -442
rect 161 -418 246 -412
rect 271 -413 308 -412
rect 161 -438 169 -418
rect 189 -438 246 -418
rect 161 -446 246 -438
rect 270 -422 308 -413
rect 270 -442 279 -422
rect 299 -442 308 -422
rect 161 -447 197 -446
rect 270 -450 308 -442
rect 374 -418 459 -412
rect 479 -413 516 -412
rect 374 -438 382 -418
rect 402 -419 459 -418
rect 402 -438 431 -419
rect 374 -439 431 -438
rect 452 -439 459 -419
rect 374 -446 459 -439
rect 478 -422 516 -413
rect 478 -442 487 -422
rect 507 -442 516 -422
rect 374 -447 410 -446
rect 478 -450 516 -442
rect 582 -418 726 -412
rect 582 -438 590 -418
rect 610 -421 698 -418
rect 610 -438 641 -421
rect 582 -441 641 -438
rect 664 -438 698 -421
rect 718 -438 726 -418
rect 664 -441 726 -438
rect 582 -446 726 -441
rect 582 -447 618 -446
rect 690 -447 726 -446
rect 792 -413 829 -412
rect 792 -414 830 -413
rect 792 -422 856 -414
rect 792 -442 801 -422
rect 821 -436 856 -422
rect 876 -436 879 -416
rect 821 -441 879 -436
rect 821 -442 856 -441
rect 58 -479 95 -450
rect 59 -481 95 -479
rect 271 -481 308 -450
rect 59 -503 308 -481
rect 479 -482 516 -450
rect 792 -454 856 -442
rect 896 -480 923 -302
rect 755 -482 923 -480
rect 479 -485 923 -482
rect 140 -509 251 -503
rect 140 -517 181 -509
rect -171 -572 -132 -528
rect 140 -537 148 -517
rect 167 -537 181 -517
rect 140 -539 181 -537
rect 209 -517 251 -509
rect 209 -537 225 -517
rect 244 -537 251 -517
rect 209 -538 251 -537
rect 477 -508 923 -485
rect 209 -539 252 -538
rect -171 -596 -131 -572
rect 140 -578 252 -539
rect 169 -596 216 -578
rect 477 -596 515 -508
rect 755 -509 923 -508
rect -171 -629 515 -596
rect 477 -631 515 -629
<< viali >>
rect 146 362 175 389
rect 220 365 249 392
rect -84 249 -55 278
rect 878 357 898 377
rect 434 264 455 284
rect 807 171 833 197
rect 432 115 453 135
rect 642 115 667 135
rect 857 118 877 138
rect 149 17 168 37
rect 226 17 245 37
rect 1084 118 1113 145
rect 1158 121 1187 148
rect 1816 113 1836 133
rect 1372 20 1393 40
rect 1745 -73 1771 -47
rect 1370 -129 1391 -109
rect 1795 -126 1815 -106
rect -78 -192 -53 -173
rect 145 -192 174 -165
rect 219 -189 248 -162
rect 877 -197 897 -177
rect 433 -290 454 -270
rect 1087 -227 1106 -207
rect 1164 -227 1183 -207
rect 1422 -200 1448 -178
rect 806 -383 832 -357
rect 431 -439 452 -419
rect 641 -441 664 -421
rect 856 -436 876 -416
rect 148 -537 167 -517
rect 225 -537 244 -517
<< metal1 >>
rect 873 460 908 462
rect -91 457 908 460
rect -92 433 908 457
rect -92 278 -44 433
rect 142 392 252 406
rect 142 389 220 392
rect 142 362 146 389
rect 175 365 220 389
rect 249 365 252 392
rect 873 382 908 433
rect 175 362 252 365
rect 142 347 252 362
rect 871 377 908 382
rect 871 357 878 377
rect 898 357 908 377
rect 871 350 908 357
rect 871 349 906 350
rect -92 249 -84 278
rect -55 249 -44 278
rect -92 244 -44 249
rect 427 284 459 291
rect 427 264 434 284
rect 455 264 459 284
rect 427 199 459 264
rect 797 199 837 200
rect 427 197 839 199
rect 427 171 807 197
rect 833 171 839 197
rect 427 163 839 171
rect 427 135 459 163
rect 872 143 906 349
rect 1810 216 1844 217
rect 941 181 1845 216
rect 427 115 432 135
rect 453 115 459 135
rect 427 108 459 115
rect 634 135 673 141
rect 634 115 642 135
rect 667 115 673 135
rect 634 108 673 115
rect 850 138 906 143
rect 850 118 857 138
rect 877 118 906 138
rect 850 111 906 118
rect 850 110 885 111
rect 642 62 673 108
rect 141 37 252 59
rect 141 17 149 37
rect 168 17 226 37
rect 245 17 252 37
rect 641 45 673 62
rect 942 45 979 181
rect 1080 148 1190 162
rect 1080 145 1158 148
rect 1080 118 1084 145
rect 1113 121 1158 145
rect 1187 121 1190 148
rect 1810 138 1844 181
rect 1113 118 1190 121
rect 1080 103 1190 118
rect 1809 133 1844 138
rect 1809 113 1816 133
rect 1836 113 1844 133
rect 1809 105 1844 113
rect 641 32 979 45
rect 141 0 252 17
rect 642 13 979 32
rect 921 12 979 13
rect 1365 40 1397 47
rect 1365 20 1372 40
rect 1393 20 1397 40
rect 1365 -45 1397 20
rect 1735 -45 1775 -44
rect 1365 -47 1777 -45
rect 1365 -73 1745 -47
rect 1771 -73 1777 -47
rect 1365 -81 1777 -73
rect -89 -120 907 -94
rect 1365 -109 1397 -81
rect 1810 -101 1844 105
rect -87 -173 -45 -120
rect -87 -192 -78 -173
rect -53 -192 -45 -173
rect -87 -202 -45 -192
rect 141 -162 251 -148
rect 141 -165 219 -162
rect 141 -192 145 -165
rect 174 -189 219 -165
rect 248 -189 251 -162
rect 871 -172 905 -120
rect 1365 -129 1370 -109
rect 1391 -129 1397 -109
rect 1365 -136 1397 -129
rect 1788 -106 1844 -101
rect 1788 -126 1795 -106
rect 1815 -126 1844 -106
rect 1788 -133 1844 -126
rect 1788 -134 1823 -133
rect 1416 -168 1457 -167
rect 174 -192 251 -189
rect 141 -207 251 -192
rect 870 -177 905 -172
rect 870 -197 877 -177
rect 897 -197 905 -177
rect 1415 -178 1457 -168
rect 870 -205 905 -197
rect 426 -270 458 -263
rect 426 -290 433 -270
rect 454 -290 458 -270
rect 426 -355 458 -290
rect 796 -355 836 -354
rect 426 -357 838 -355
rect 426 -383 806 -357
rect 832 -383 838 -357
rect 426 -391 838 -383
rect 426 -419 458 -391
rect 871 -411 905 -205
rect 1079 -207 1190 -185
rect 1079 -227 1087 -207
rect 1106 -227 1164 -207
rect 1183 -227 1190 -207
rect 1079 -244 1190 -227
rect 1415 -200 1422 -178
rect 1448 -200 1457 -178
rect 1415 -209 1457 -200
rect 632 -414 675 -412
rect 426 -439 431 -419
rect 452 -439 458 -419
rect 426 -446 458 -439
rect 631 -421 675 -414
rect 631 -441 641 -421
rect 664 -441 675 -421
rect 631 -445 675 -441
rect 849 -416 905 -411
rect 849 -436 856 -416
rect 876 -436 905 -416
rect 849 -443 905 -436
rect 961 -275 994 -274
rect 1415 -275 1452 -209
rect 961 -304 1452 -275
rect 849 -444 884 -443
rect 140 -517 251 -495
rect 140 -537 148 -517
rect 167 -537 225 -517
rect 244 -537 251 -517
rect 140 -554 251 -537
rect 631 -526 673 -445
rect 961 -524 994 -304
rect 1415 -306 1452 -304
rect 933 -526 994 -524
rect 631 -555 994 -526
rect 631 -557 933 -555
<< labels >>
rlabel locali 13 173 35 188 1 d0
rlabel metal1 182 396 210 401 1 vdd
rlabel metal1 179 3 213 9 1 gnd
rlabel locali 950 -75 978 -54 1 d1
rlabel metal1 1117 -241 1151 -235 1 gnd
rlabel metal1 1120 152 1148 157 1 vdd
rlabel locali 1581 -36 1603 -21 1 vout
rlabel locali 12 -381 34 -366 1 d0
rlabel metal1 181 -158 209 -153 1 vdd
rlabel metal1 178 -551 212 -545 1 gnd
rlabel locali -167 458 -139 466 1 vref
<< end >>
