magic
tech sky130A
timestamp 1616157205
<< nwell >>
rect -19 0 792 150
<< nmos >>
rect 45 -101 95 -59
rect 258 -101 308 -59
rect 466 -101 516 -59
rect 674 -101 724 -59
<< pmos >>
rect 45 18 95 118
rect 258 18 308 118
rect 466 18 516 118
rect 674 18 724 118
<< ndiff >>
rect -4 -69 45 -59
rect -4 -89 7 -69
rect 27 -89 45 -69
rect -4 -101 45 -89
rect 95 -65 139 -59
rect 95 -85 110 -65
rect 130 -85 139 -65
rect 95 -101 139 -85
rect 209 -69 258 -59
rect 209 -89 220 -69
rect 240 -89 258 -69
rect 209 -101 258 -89
rect 308 -65 352 -59
rect 308 -85 323 -65
rect 343 -85 352 -65
rect 308 -101 352 -85
rect 417 -69 466 -59
rect 417 -89 428 -69
rect 448 -89 466 -69
rect 417 -101 466 -89
rect 516 -65 560 -59
rect 516 -85 531 -65
rect 551 -85 560 -65
rect 516 -101 560 -85
rect 630 -65 674 -59
rect 630 -85 639 -65
rect 659 -85 674 -65
rect 630 -101 674 -85
rect 724 -69 773 -59
rect 724 -89 742 -69
rect 762 -89 773 -69
rect 724 -101 773 -89
<< pdiff >>
rect 1 80 45 118
rect 1 60 13 80
rect 33 60 45 80
rect 1 18 45 60
rect 95 80 137 118
rect 95 60 109 80
rect 129 60 137 80
rect 95 18 137 60
rect 214 80 258 118
rect 214 60 226 80
rect 246 60 258 80
rect 214 18 258 60
rect 308 80 350 118
rect 308 60 322 80
rect 342 60 350 80
rect 308 18 350 60
rect 422 80 466 118
rect 422 60 434 80
rect 454 60 466 80
rect 422 18 466 60
rect 516 80 558 118
rect 516 60 530 80
rect 550 60 558 80
rect 516 18 558 60
rect 632 80 674 118
rect 632 60 640 80
rect 660 60 674 80
rect 632 18 674 60
rect 724 87 769 118
rect 724 80 768 87
rect 724 60 736 80
rect 756 60 768 80
rect 724 18 768 60
<< ndiffc >>
rect 7 -89 27 -69
rect 110 -85 130 -65
rect 220 -89 240 -69
rect 323 -85 343 -65
rect 428 -89 448 -69
rect 531 -85 551 -65
rect 639 -85 659 -65
rect 742 -89 762 -69
<< pdiffc >>
rect 13 60 33 80
rect 109 60 129 80
rect 226 60 246 80
rect 322 60 342 80
rect 434 60 454 80
rect 530 60 550 80
rect 640 60 660 80
rect 736 60 756 80
<< poly >>
rect 45 118 95 131
rect 258 118 308 131
rect 466 118 516 131
rect 674 118 724 131
rect 45 -10 95 18
rect 45 -30 58 -10
rect 78 -30 95 -10
rect 45 -59 95 -30
rect 258 -11 308 18
rect 258 -35 269 -11
rect 293 -35 308 -11
rect 258 -59 308 -35
rect 466 -6 516 18
rect 466 -30 478 -6
rect 502 -30 516 -6
rect 466 -59 516 -30
rect 674 -8 724 18
rect 674 -34 692 -8
rect 718 -34 724 -8
rect 674 -59 724 -34
rect 45 -117 95 -101
rect 258 -117 308 -101
rect 466 -117 516 -101
rect 674 -117 724 -101
<< polycont >>
rect 58 -30 78 -10
rect 269 -35 293 -11
rect 478 -30 502 -6
rect 692 -34 718 -8
<< locali >>
rect 4 151 254 175
rect 4 80 41 151
rect 156 90 187 91
rect 4 60 13 80
rect 33 60 41 80
rect 4 50 41 60
rect 100 80 187 90
rect 100 60 109 80
rect 129 60 187 80
rect 100 51 187 60
rect 100 50 137 51
rect 156 -2 187 51
rect 217 80 254 151
rect 425 156 818 176
rect 838 156 841 176
rect 425 151 841 156
rect 425 150 766 151
rect 369 90 400 91
rect 217 60 226 80
rect 246 60 254 80
rect 217 50 254 60
rect 313 83 400 90
rect 313 80 374 83
rect 313 60 322 80
rect 342 63 374 80
rect 395 63 400 83
rect 342 60 400 63
rect 313 53 400 60
rect 425 80 462 150
rect 728 149 765 150
rect 577 90 613 91
rect 425 60 434 80
rect 454 60 462 80
rect 313 51 369 53
rect 313 50 350 51
rect 425 50 462 60
rect 521 80 669 90
rect 769 87 865 89
rect 521 60 530 80
rect 550 60 640 80
rect 660 60 669 80
rect 521 51 669 60
rect 727 80 865 87
rect 727 60 736 80
rect 756 60 865 80
rect 727 51 865 60
rect 521 50 558 51
rect 577 -1 613 51
rect 632 50 669 51
rect 728 50 765 51
rect 48 -3 89 -2
rect -60 -10 89 -3
rect -60 -30 58 -10
rect 78 -30 89 -10
rect -60 -38 89 -30
rect 156 -6 515 -2
rect 156 -11 478 -6
rect 156 -35 269 -11
rect 293 -30 478 -11
rect 502 -30 515 -6
rect 293 -35 515 -30
rect 156 -38 515 -35
rect 577 -38 612 -1
rect 680 -4 780 -1
rect 680 -8 747 -4
rect 680 -34 692 -8
rect 718 -30 747 -8
rect 773 -30 780 -4
rect 718 -34 780 -30
rect 680 -38 780 -34
rect 156 -59 187 -38
rect 577 -59 613 -38
rect -1 -60 36 -59
rect -2 -69 36 -60
rect -2 -89 7 -69
rect 27 -89 36 -69
rect -2 -97 36 -89
rect 102 -65 187 -59
rect 212 -60 249 -59
rect 102 -85 110 -65
rect 130 -85 187 -65
rect 102 -93 187 -85
rect 211 -69 249 -60
rect 211 -89 220 -69
rect 240 -89 249 -69
rect 102 -94 138 -93
rect 211 -97 249 -89
rect 315 -65 400 -59
rect 420 -60 457 -59
rect 315 -85 323 -65
rect 343 -66 400 -65
rect 343 -85 372 -66
rect 315 -86 372 -85
rect 393 -86 400 -66
rect 315 -93 400 -86
rect 419 -69 457 -60
rect 419 -89 428 -69
rect 448 -89 457 -69
rect 315 -94 351 -93
rect 419 -97 457 -89
rect 523 -65 667 -59
rect 523 -85 531 -65
rect 551 -85 639 -65
rect 659 -85 667 -65
rect 523 -93 667 -85
rect 523 -94 559 -93
rect 631 -94 667 -93
rect 733 -60 770 -59
rect 733 -61 771 -60
rect 733 -69 797 -61
rect 733 -89 742 -69
rect 762 -83 797 -69
rect 817 -83 820 -63
rect 762 -88 820 -83
rect 762 -89 797 -88
rect -1 -126 36 -97
rect 0 -128 36 -126
rect 212 -128 249 -97
rect 0 -150 249 -128
rect 420 -129 457 -97
rect 733 -101 797 -89
rect 837 -127 864 51
rect 696 -129 864 -127
rect 420 -155 864 -129
rect 696 -156 864 -155
<< viali >>
rect 818 156 838 176
rect 374 63 395 83
rect 747 -30 773 -4
rect 372 -86 393 -66
rect 797 -83 817 -63
<< metal1 >>
rect 814 181 846 182
rect 811 176 846 181
rect 811 156 818 176
rect 838 156 846 176
rect 811 148 846 156
rect 367 83 399 90
rect 367 63 374 83
rect 395 63 399 83
rect 367 -2 399 63
rect 737 -2 777 -1
rect 367 -4 779 -2
rect 367 -30 747 -4
rect 773 -30 779 -4
rect 367 -38 779 -30
rect 367 -66 399 -38
rect 812 -58 846 148
rect 367 -86 372 -66
rect 393 -86 399 -66
rect 367 -93 399 -86
rect 790 -63 846 -58
rect 790 -83 797 -63
rect 817 -83 846 -63
rect 790 -90 846 -83
rect 790 -91 825 -90
<< labels >>
rlabel locali 7 160 36 166 1 vdd
rlabel locali 220 157 249 163 1 vdd
rlabel locali 583 7 605 22 1 vout
rlabel locali -47 -28 -25 -13 1 d0
rlabel nwell 374 127 397 130 1 vdd
rlabel locali 4 -139 33 -133 1 gnd
rlabel locali 217 -139 246 -133 1 gnd
rlabel space 314 -144 343 -135 1 gnd
<< end >>
