magic
tech sky130A
timestamp 1620565581
<< nwell >>
rect 318 8703 645 8777
rect 318 8553 1129 8703
rect 1256 8459 1583 8533
rect 3801 8483 4612 8633
rect 1256 8309 2067 8459
rect 4285 8409 4612 8483
rect 317 8149 644 8223
rect 2862 8173 3673 8323
rect 317 7999 1128 8149
rect 3346 8099 3673 8173
rect 1397 7867 1724 7941
rect 3800 7929 4611 8079
rect 1397 7717 2208 7867
rect 4284 7855 4611 7929
rect 319 7600 646 7674
rect 2722 7662 3533 7812
rect 319 7450 1130 7600
rect 3206 7588 3533 7662
rect 1257 7356 1584 7430
rect 3802 7380 4613 7530
rect 1257 7206 2068 7356
rect 4286 7306 4613 7380
rect 318 7046 645 7120
rect 2863 7070 3674 7220
rect 318 6896 1129 7046
rect 3347 6996 3674 7070
rect 1367 6777 1694 6851
rect 3801 6826 4612 6976
rect 1367 6627 2178 6777
rect 4285 6752 4612 6826
rect 319 6497 646 6571
rect 2753 6546 3564 6696
rect 319 6347 1130 6497
rect 3237 6472 3564 6546
rect 1257 6253 1584 6327
rect 3802 6277 4613 6427
rect 1257 6103 2068 6253
rect 4286 6203 4613 6277
rect 318 5943 645 6017
rect 2863 5967 3674 6117
rect 318 5793 1129 5943
rect 3347 5893 3674 5967
rect 1398 5661 1725 5735
rect 3801 5723 4612 5873
rect 1398 5511 2209 5661
rect 4285 5649 4612 5723
rect 320 5394 647 5468
rect 2723 5456 3534 5606
rect 320 5244 1131 5394
rect 3207 5382 3534 5456
rect 1258 5150 1585 5224
rect 3803 5174 4614 5324
rect 1258 5000 2069 5150
rect 4287 5100 4614 5174
rect 319 4840 646 4914
rect 2864 4864 3675 5014
rect 319 4690 1130 4840
rect 3348 4790 3675 4864
rect 1367 4577 1694 4651
rect 3802 4620 4613 4770
rect 1367 4427 2178 4577
rect 4286 4546 4613 4620
rect 320 4291 647 4365
rect 2755 4334 3566 4484
rect 320 4141 1131 4291
rect 3239 4260 3566 4334
rect 1258 4047 1585 4121
rect 3803 4071 4614 4221
rect 1258 3897 2069 4047
rect 4287 3997 4614 4071
rect 319 3737 646 3811
rect 2864 3761 3675 3911
rect 319 3587 1130 3737
rect 3348 3687 3675 3761
rect 1399 3455 1726 3529
rect 3802 3517 4613 3667
rect 1399 3305 2210 3455
rect 4286 3443 4613 3517
rect 321 3188 648 3262
rect 2724 3250 3535 3400
rect 321 3038 1132 3188
rect 3208 3176 3535 3250
rect 1259 2944 1586 3018
rect 3804 2968 4615 3118
rect 1259 2794 2070 2944
rect 4288 2894 4615 2968
rect 320 2634 647 2708
rect 2865 2658 3676 2808
rect 320 2484 1131 2634
rect 3349 2584 3676 2658
rect 1369 2365 1696 2439
rect 3803 2414 4614 2564
rect 1369 2215 2180 2365
rect 4287 2340 4614 2414
rect 321 2085 648 2159
rect 2755 2134 3566 2284
rect 321 1935 1132 2085
rect 3239 2060 3566 2134
rect 1259 1841 1586 1915
rect 3804 1865 4615 2015
rect 1259 1691 2070 1841
rect 4288 1791 4615 1865
rect 320 1531 647 1605
rect 2865 1555 3676 1705
rect 320 1381 1131 1531
rect 3349 1481 3676 1555
rect 1400 1249 1727 1323
rect 3803 1311 4614 1461
rect 1400 1099 2211 1249
rect 4287 1237 4614 1311
rect 322 982 649 1056
rect 2725 1044 3536 1194
rect 322 832 1133 982
rect 3209 970 3536 1044
rect 1260 738 1587 812
rect 3805 762 4616 912
rect 1260 588 2071 738
rect 4289 688 4616 762
rect 321 428 648 502
rect 2866 452 3677 602
rect 321 278 1132 428
rect 3350 378 3677 452
rect 3804 208 4615 358
rect 4288 134 4615 208
rect 1568 -131 1895 -57
rect 1568 -281 2379 -131
<< nmos >>
rect 3869 8692 3919 8734
rect 4077 8692 4127 8734
rect 4285 8692 4335 8734
rect 4498 8692 4548 8734
rect 382 8452 432 8494
rect 595 8452 645 8494
rect 803 8452 853 8494
rect 1011 8452 1061 8494
rect 2930 8382 2980 8424
rect 3138 8382 3188 8424
rect 3346 8382 3396 8424
rect 3559 8382 3609 8424
rect 1320 8208 1370 8250
rect 1533 8208 1583 8250
rect 1741 8208 1791 8250
rect 1949 8208 1999 8250
rect 3868 8138 3918 8180
rect 4076 8138 4126 8180
rect 4284 8138 4334 8180
rect 4497 8138 4547 8180
rect 381 7898 431 7940
rect 594 7898 644 7940
rect 802 7898 852 7940
rect 1010 7898 1060 7940
rect 2790 7871 2840 7913
rect 2998 7871 3048 7913
rect 3206 7871 3256 7913
rect 3419 7871 3469 7913
rect 1461 7616 1511 7658
rect 1674 7616 1724 7658
rect 1882 7616 1932 7658
rect 2090 7616 2140 7658
rect 3870 7589 3920 7631
rect 4078 7589 4128 7631
rect 4286 7589 4336 7631
rect 4499 7589 4549 7631
rect 383 7349 433 7391
rect 596 7349 646 7391
rect 804 7349 854 7391
rect 1012 7349 1062 7391
rect 2931 7279 2981 7321
rect 3139 7279 3189 7321
rect 3347 7279 3397 7321
rect 3560 7279 3610 7321
rect 1321 7105 1371 7147
rect 1534 7105 1584 7147
rect 1742 7105 1792 7147
rect 1950 7105 2000 7147
rect 3869 7035 3919 7077
rect 4077 7035 4127 7077
rect 4285 7035 4335 7077
rect 4498 7035 4548 7077
rect 382 6795 432 6837
rect 595 6795 645 6837
rect 803 6795 853 6837
rect 1011 6795 1061 6837
rect 2821 6755 2871 6797
rect 3029 6755 3079 6797
rect 3237 6755 3287 6797
rect 3450 6755 3500 6797
rect 1431 6526 1481 6568
rect 1644 6526 1694 6568
rect 1852 6526 1902 6568
rect 2060 6526 2110 6568
rect 3870 6486 3920 6528
rect 4078 6486 4128 6528
rect 4286 6486 4336 6528
rect 4499 6486 4549 6528
rect 383 6246 433 6288
rect 596 6246 646 6288
rect 804 6246 854 6288
rect 1012 6246 1062 6288
rect 2931 6176 2981 6218
rect 3139 6176 3189 6218
rect 3347 6176 3397 6218
rect 3560 6176 3610 6218
rect 1321 6002 1371 6044
rect 1534 6002 1584 6044
rect 1742 6002 1792 6044
rect 1950 6002 2000 6044
rect 3869 5932 3919 5974
rect 4077 5932 4127 5974
rect 4285 5932 4335 5974
rect 4498 5932 4548 5974
rect 382 5692 432 5734
rect 595 5692 645 5734
rect 803 5692 853 5734
rect 1011 5692 1061 5734
rect 2791 5665 2841 5707
rect 2999 5665 3049 5707
rect 3207 5665 3257 5707
rect 3420 5665 3470 5707
rect 1462 5410 1512 5452
rect 1675 5410 1725 5452
rect 1883 5410 1933 5452
rect 2091 5410 2141 5452
rect 3871 5383 3921 5425
rect 4079 5383 4129 5425
rect 4287 5383 4337 5425
rect 4500 5383 4550 5425
rect 384 5143 434 5185
rect 597 5143 647 5185
rect 805 5143 855 5185
rect 1013 5143 1063 5185
rect 2932 5073 2982 5115
rect 3140 5073 3190 5115
rect 3348 5073 3398 5115
rect 3561 5073 3611 5115
rect 1322 4899 1372 4941
rect 1535 4899 1585 4941
rect 1743 4899 1793 4941
rect 1951 4899 2001 4941
rect 3870 4829 3920 4871
rect 4078 4829 4128 4871
rect 4286 4829 4336 4871
rect 4499 4829 4549 4871
rect 383 4589 433 4631
rect 596 4589 646 4631
rect 804 4589 854 4631
rect 1012 4589 1062 4631
rect 2823 4543 2873 4585
rect 3031 4543 3081 4585
rect 3239 4543 3289 4585
rect 3452 4543 3502 4585
rect 1431 4326 1481 4368
rect 1644 4326 1694 4368
rect 1852 4326 1902 4368
rect 2060 4326 2110 4368
rect 3871 4280 3921 4322
rect 4079 4280 4129 4322
rect 4287 4280 4337 4322
rect 4500 4280 4550 4322
rect 384 4040 434 4082
rect 597 4040 647 4082
rect 805 4040 855 4082
rect 1013 4040 1063 4082
rect 2932 3970 2982 4012
rect 3140 3970 3190 4012
rect 3348 3970 3398 4012
rect 3561 3970 3611 4012
rect 1322 3796 1372 3838
rect 1535 3796 1585 3838
rect 1743 3796 1793 3838
rect 1951 3796 2001 3838
rect 3870 3726 3920 3768
rect 4078 3726 4128 3768
rect 4286 3726 4336 3768
rect 4499 3726 4549 3768
rect 383 3486 433 3528
rect 596 3486 646 3528
rect 804 3486 854 3528
rect 1012 3486 1062 3528
rect 2792 3459 2842 3501
rect 3000 3459 3050 3501
rect 3208 3459 3258 3501
rect 3421 3459 3471 3501
rect 1463 3204 1513 3246
rect 1676 3204 1726 3246
rect 1884 3204 1934 3246
rect 2092 3204 2142 3246
rect 3872 3177 3922 3219
rect 4080 3177 4130 3219
rect 4288 3177 4338 3219
rect 4501 3177 4551 3219
rect 385 2937 435 2979
rect 598 2937 648 2979
rect 806 2937 856 2979
rect 1014 2937 1064 2979
rect 2933 2867 2983 2909
rect 3141 2867 3191 2909
rect 3349 2867 3399 2909
rect 3562 2867 3612 2909
rect 1323 2693 1373 2735
rect 1536 2693 1586 2735
rect 1744 2693 1794 2735
rect 1952 2693 2002 2735
rect 3871 2623 3921 2665
rect 4079 2623 4129 2665
rect 4287 2623 4337 2665
rect 4500 2623 4550 2665
rect 384 2383 434 2425
rect 597 2383 647 2425
rect 805 2383 855 2425
rect 1013 2383 1063 2425
rect 2823 2343 2873 2385
rect 3031 2343 3081 2385
rect 3239 2343 3289 2385
rect 3452 2343 3502 2385
rect 1433 2114 1483 2156
rect 1646 2114 1696 2156
rect 1854 2114 1904 2156
rect 2062 2114 2112 2156
rect 3872 2074 3922 2116
rect 4080 2074 4130 2116
rect 4288 2074 4338 2116
rect 4501 2074 4551 2116
rect 385 1834 435 1876
rect 598 1834 648 1876
rect 806 1834 856 1876
rect 1014 1834 1064 1876
rect 2933 1764 2983 1806
rect 3141 1764 3191 1806
rect 3349 1764 3399 1806
rect 3562 1764 3612 1806
rect 1323 1590 1373 1632
rect 1536 1590 1586 1632
rect 1744 1590 1794 1632
rect 1952 1590 2002 1632
rect 3871 1520 3921 1562
rect 4079 1520 4129 1562
rect 4287 1520 4337 1562
rect 4500 1520 4550 1562
rect 384 1280 434 1322
rect 597 1280 647 1322
rect 805 1280 855 1322
rect 1013 1280 1063 1322
rect 2793 1253 2843 1295
rect 3001 1253 3051 1295
rect 3209 1253 3259 1295
rect 3422 1253 3472 1295
rect 1464 998 1514 1040
rect 1677 998 1727 1040
rect 1885 998 1935 1040
rect 2093 998 2143 1040
rect 3873 971 3923 1013
rect 4081 971 4131 1013
rect 4289 971 4339 1013
rect 4502 971 4552 1013
rect 386 731 436 773
rect 599 731 649 773
rect 807 731 857 773
rect 1015 731 1065 773
rect 2934 661 2984 703
rect 3142 661 3192 703
rect 3350 661 3400 703
rect 3563 661 3613 703
rect 1324 487 1374 529
rect 1537 487 1587 529
rect 1745 487 1795 529
rect 1953 487 2003 529
rect 3872 417 3922 459
rect 4080 417 4130 459
rect 4288 417 4338 459
rect 4501 417 4551 459
rect 385 177 435 219
rect 598 177 648 219
rect 806 177 856 219
rect 1014 177 1064 219
rect 1632 -382 1682 -340
rect 1845 -382 1895 -340
rect 2053 -382 2103 -340
rect 2261 -382 2311 -340
<< pmos >>
rect 382 8571 432 8671
rect 595 8571 645 8671
rect 803 8571 853 8671
rect 1011 8571 1061 8671
rect 3869 8515 3919 8615
rect 4077 8515 4127 8615
rect 4285 8515 4335 8615
rect 4498 8515 4548 8615
rect 1320 8327 1370 8427
rect 1533 8327 1583 8427
rect 1741 8327 1791 8427
rect 1949 8327 1999 8427
rect 2930 8205 2980 8305
rect 3138 8205 3188 8305
rect 3346 8205 3396 8305
rect 3559 8205 3609 8305
rect 381 8017 431 8117
rect 594 8017 644 8117
rect 802 8017 852 8117
rect 1010 8017 1060 8117
rect 3868 7961 3918 8061
rect 4076 7961 4126 8061
rect 4284 7961 4334 8061
rect 4497 7961 4547 8061
rect 1461 7735 1511 7835
rect 1674 7735 1724 7835
rect 1882 7735 1932 7835
rect 2090 7735 2140 7835
rect 2790 7694 2840 7794
rect 2998 7694 3048 7794
rect 3206 7694 3256 7794
rect 3419 7694 3469 7794
rect 383 7468 433 7568
rect 596 7468 646 7568
rect 804 7468 854 7568
rect 1012 7468 1062 7568
rect 3870 7412 3920 7512
rect 4078 7412 4128 7512
rect 4286 7412 4336 7512
rect 4499 7412 4549 7512
rect 1321 7224 1371 7324
rect 1534 7224 1584 7324
rect 1742 7224 1792 7324
rect 1950 7224 2000 7324
rect 2931 7102 2981 7202
rect 3139 7102 3189 7202
rect 3347 7102 3397 7202
rect 3560 7102 3610 7202
rect 382 6914 432 7014
rect 595 6914 645 7014
rect 803 6914 853 7014
rect 1011 6914 1061 7014
rect 3869 6858 3919 6958
rect 4077 6858 4127 6958
rect 4285 6858 4335 6958
rect 4498 6858 4548 6958
rect 1431 6645 1481 6745
rect 1644 6645 1694 6745
rect 1852 6645 1902 6745
rect 2060 6645 2110 6745
rect 2821 6578 2871 6678
rect 3029 6578 3079 6678
rect 3237 6578 3287 6678
rect 3450 6578 3500 6678
rect 383 6365 433 6465
rect 596 6365 646 6465
rect 804 6365 854 6465
rect 1012 6365 1062 6465
rect 3870 6309 3920 6409
rect 4078 6309 4128 6409
rect 4286 6309 4336 6409
rect 4499 6309 4549 6409
rect 1321 6121 1371 6221
rect 1534 6121 1584 6221
rect 1742 6121 1792 6221
rect 1950 6121 2000 6221
rect 2931 5999 2981 6099
rect 3139 5999 3189 6099
rect 3347 5999 3397 6099
rect 3560 5999 3610 6099
rect 382 5811 432 5911
rect 595 5811 645 5911
rect 803 5811 853 5911
rect 1011 5811 1061 5911
rect 3869 5755 3919 5855
rect 4077 5755 4127 5855
rect 4285 5755 4335 5855
rect 4498 5755 4548 5855
rect 1462 5529 1512 5629
rect 1675 5529 1725 5629
rect 1883 5529 1933 5629
rect 2091 5529 2141 5629
rect 2791 5488 2841 5588
rect 2999 5488 3049 5588
rect 3207 5488 3257 5588
rect 3420 5488 3470 5588
rect 384 5262 434 5362
rect 597 5262 647 5362
rect 805 5262 855 5362
rect 1013 5262 1063 5362
rect 3871 5206 3921 5306
rect 4079 5206 4129 5306
rect 4287 5206 4337 5306
rect 4500 5206 4550 5306
rect 1322 5018 1372 5118
rect 1535 5018 1585 5118
rect 1743 5018 1793 5118
rect 1951 5018 2001 5118
rect 2932 4896 2982 4996
rect 3140 4896 3190 4996
rect 3348 4896 3398 4996
rect 3561 4896 3611 4996
rect 383 4708 433 4808
rect 596 4708 646 4808
rect 804 4708 854 4808
rect 1012 4708 1062 4808
rect 3870 4652 3920 4752
rect 4078 4652 4128 4752
rect 4286 4652 4336 4752
rect 4499 4652 4549 4752
rect 1431 4445 1481 4545
rect 1644 4445 1694 4545
rect 1852 4445 1902 4545
rect 2060 4445 2110 4545
rect 2823 4366 2873 4466
rect 3031 4366 3081 4466
rect 3239 4366 3289 4466
rect 3452 4366 3502 4466
rect 384 4159 434 4259
rect 597 4159 647 4259
rect 805 4159 855 4259
rect 1013 4159 1063 4259
rect 3871 4103 3921 4203
rect 4079 4103 4129 4203
rect 4287 4103 4337 4203
rect 4500 4103 4550 4203
rect 1322 3915 1372 4015
rect 1535 3915 1585 4015
rect 1743 3915 1793 4015
rect 1951 3915 2001 4015
rect 2932 3793 2982 3893
rect 3140 3793 3190 3893
rect 3348 3793 3398 3893
rect 3561 3793 3611 3893
rect 383 3605 433 3705
rect 596 3605 646 3705
rect 804 3605 854 3705
rect 1012 3605 1062 3705
rect 3870 3549 3920 3649
rect 4078 3549 4128 3649
rect 4286 3549 4336 3649
rect 4499 3549 4549 3649
rect 1463 3323 1513 3423
rect 1676 3323 1726 3423
rect 1884 3323 1934 3423
rect 2092 3323 2142 3423
rect 2792 3282 2842 3382
rect 3000 3282 3050 3382
rect 3208 3282 3258 3382
rect 3421 3282 3471 3382
rect 385 3056 435 3156
rect 598 3056 648 3156
rect 806 3056 856 3156
rect 1014 3056 1064 3156
rect 3872 3000 3922 3100
rect 4080 3000 4130 3100
rect 4288 3000 4338 3100
rect 4501 3000 4551 3100
rect 1323 2812 1373 2912
rect 1536 2812 1586 2912
rect 1744 2812 1794 2912
rect 1952 2812 2002 2912
rect 2933 2690 2983 2790
rect 3141 2690 3191 2790
rect 3349 2690 3399 2790
rect 3562 2690 3612 2790
rect 384 2502 434 2602
rect 597 2502 647 2602
rect 805 2502 855 2602
rect 1013 2502 1063 2602
rect 3871 2446 3921 2546
rect 4079 2446 4129 2546
rect 4287 2446 4337 2546
rect 4500 2446 4550 2546
rect 1433 2233 1483 2333
rect 1646 2233 1696 2333
rect 1854 2233 1904 2333
rect 2062 2233 2112 2333
rect 2823 2166 2873 2266
rect 3031 2166 3081 2266
rect 3239 2166 3289 2266
rect 3452 2166 3502 2266
rect 385 1953 435 2053
rect 598 1953 648 2053
rect 806 1953 856 2053
rect 1014 1953 1064 2053
rect 3872 1897 3922 1997
rect 4080 1897 4130 1997
rect 4288 1897 4338 1997
rect 4501 1897 4551 1997
rect 1323 1709 1373 1809
rect 1536 1709 1586 1809
rect 1744 1709 1794 1809
rect 1952 1709 2002 1809
rect 2933 1587 2983 1687
rect 3141 1587 3191 1687
rect 3349 1587 3399 1687
rect 3562 1587 3612 1687
rect 384 1399 434 1499
rect 597 1399 647 1499
rect 805 1399 855 1499
rect 1013 1399 1063 1499
rect 3871 1343 3921 1443
rect 4079 1343 4129 1443
rect 4287 1343 4337 1443
rect 4500 1343 4550 1443
rect 1464 1117 1514 1217
rect 1677 1117 1727 1217
rect 1885 1117 1935 1217
rect 2093 1117 2143 1217
rect 2793 1076 2843 1176
rect 3001 1076 3051 1176
rect 3209 1076 3259 1176
rect 3422 1076 3472 1176
rect 386 850 436 950
rect 599 850 649 950
rect 807 850 857 950
rect 1015 850 1065 950
rect 3873 794 3923 894
rect 4081 794 4131 894
rect 4289 794 4339 894
rect 4502 794 4552 894
rect 1324 606 1374 706
rect 1537 606 1587 706
rect 1745 606 1795 706
rect 1953 606 2003 706
rect 2934 484 2984 584
rect 3142 484 3192 584
rect 3350 484 3400 584
rect 3563 484 3613 584
rect 385 296 435 396
rect 598 296 648 396
rect 806 296 856 396
rect 1014 296 1064 396
rect 3872 240 3922 340
rect 4080 240 4130 340
rect 4288 240 4338 340
rect 4501 240 4551 340
rect 1632 -263 1682 -163
rect 1845 -263 1895 -163
rect 2053 -263 2103 -163
rect 2261 -263 2311 -163
<< ndiff >>
rect 3820 8722 3869 8734
rect 3820 8702 3831 8722
rect 3851 8702 3869 8722
rect 3820 8692 3869 8702
rect 3919 8718 3963 8734
rect 3919 8698 3934 8718
rect 3954 8698 3963 8718
rect 3919 8692 3963 8698
rect 4033 8718 4077 8734
rect 4033 8698 4042 8718
rect 4062 8698 4077 8718
rect 4033 8692 4077 8698
rect 4127 8722 4176 8734
rect 4127 8702 4145 8722
rect 4165 8702 4176 8722
rect 4127 8692 4176 8702
rect 4241 8718 4285 8734
rect 4241 8698 4250 8718
rect 4270 8698 4285 8718
rect 4241 8692 4285 8698
rect 4335 8722 4384 8734
rect 4335 8702 4353 8722
rect 4373 8702 4384 8722
rect 4335 8692 4384 8702
rect 4454 8718 4498 8734
rect 4454 8698 4463 8718
rect 4483 8698 4498 8718
rect 4454 8692 4498 8698
rect 4548 8722 4597 8734
rect 4548 8702 4566 8722
rect 4586 8702 4597 8722
rect 4548 8692 4597 8702
rect 333 8484 382 8494
rect 333 8464 344 8484
rect 364 8464 382 8484
rect 333 8452 382 8464
rect 432 8488 476 8494
rect 432 8468 447 8488
rect 467 8468 476 8488
rect 432 8452 476 8468
rect 546 8484 595 8494
rect 546 8464 557 8484
rect 577 8464 595 8484
rect 546 8452 595 8464
rect 645 8488 689 8494
rect 645 8468 660 8488
rect 680 8468 689 8488
rect 645 8452 689 8468
rect 754 8484 803 8494
rect 754 8464 765 8484
rect 785 8464 803 8484
rect 754 8452 803 8464
rect 853 8488 897 8494
rect 853 8468 868 8488
rect 888 8468 897 8488
rect 853 8452 897 8468
rect 967 8488 1011 8494
rect 967 8468 976 8488
rect 996 8468 1011 8488
rect 967 8452 1011 8468
rect 1061 8484 1110 8494
rect 1061 8464 1079 8484
rect 1099 8464 1110 8484
rect 1061 8452 1110 8464
rect 2881 8412 2930 8424
rect 2881 8392 2892 8412
rect 2912 8392 2930 8412
rect 2881 8382 2930 8392
rect 2980 8408 3024 8424
rect 2980 8388 2995 8408
rect 3015 8388 3024 8408
rect 2980 8382 3024 8388
rect 3094 8408 3138 8424
rect 3094 8388 3103 8408
rect 3123 8388 3138 8408
rect 3094 8382 3138 8388
rect 3188 8412 3237 8424
rect 3188 8392 3206 8412
rect 3226 8392 3237 8412
rect 3188 8382 3237 8392
rect 3302 8408 3346 8424
rect 3302 8388 3311 8408
rect 3331 8388 3346 8408
rect 3302 8382 3346 8388
rect 3396 8412 3445 8424
rect 3396 8392 3414 8412
rect 3434 8392 3445 8412
rect 3396 8382 3445 8392
rect 3515 8408 3559 8424
rect 3515 8388 3524 8408
rect 3544 8388 3559 8408
rect 3515 8382 3559 8388
rect 3609 8412 3658 8424
rect 3609 8392 3627 8412
rect 3647 8392 3658 8412
rect 3609 8382 3658 8392
rect 1271 8240 1320 8250
rect 1271 8220 1282 8240
rect 1302 8220 1320 8240
rect 1271 8208 1320 8220
rect 1370 8244 1414 8250
rect 1370 8224 1385 8244
rect 1405 8224 1414 8244
rect 1370 8208 1414 8224
rect 1484 8240 1533 8250
rect 1484 8220 1495 8240
rect 1515 8220 1533 8240
rect 1484 8208 1533 8220
rect 1583 8244 1627 8250
rect 1583 8224 1598 8244
rect 1618 8224 1627 8244
rect 1583 8208 1627 8224
rect 1692 8240 1741 8250
rect 1692 8220 1703 8240
rect 1723 8220 1741 8240
rect 1692 8208 1741 8220
rect 1791 8244 1835 8250
rect 1791 8224 1806 8244
rect 1826 8224 1835 8244
rect 1791 8208 1835 8224
rect 1905 8244 1949 8250
rect 1905 8224 1914 8244
rect 1934 8224 1949 8244
rect 1905 8208 1949 8224
rect 1999 8240 2048 8250
rect 1999 8220 2017 8240
rect 2037 8220 2048 8240
rect 1999 8208 2048 8220
rect 3819 8168 3868 8180
rect 3819 8148 3830 8168
rect 3850 8148 3868 8168
rect 3819 8138 3868 8148
rect 3918 8164 3962 8180
rect 3918 8144 3933 8164
rect 3953 8144 3962 8164
rect 3918 8138 3962 8144
rect 4032 8164 4076 8180
rect 4032 8144 4041 8164
rect 4061 8144 4076 8164
rect 4032 8138 4076 8144
rect 4126 8168 4175 8180
rect 4126 8148 4144 8168
rect 4164 8148 4175 8168
rect 4126 8138 4175 8148
rect 4240 8164 4284 8180
rect 4240 8144 4249 8164
rect 4269 8144 4284 8164
rect 4240 8138 4284 8144
rect 4334 8168 4383 8180
rect 4334 8148 4352 8168
rect 4372 8148 4383 8168
rect 4334 8138 4383 8148
rect 4453 8164 4497 8180
rect 4453 8144 4462 8164
rect 4482 8144 4497 8164
rect 4453 8138 4497 8144
rect 4547 8168 4596 8180
rect 4547 8148 4565 8168
rect 4585 8148 4596 8168
rect 4547 8138 4596 8148
rect 332 7930 381 7940
rect 332 7910 343 7930
rect 363 7910 381 7930
rect 332 7898 381 7910
rect 431 7934 475 7940
rect 431 7914 446 7934
rect 466 7914 475 7934
rect 431 7898 475 7914
rect 545 7930 594 7940
rect 545 7910 556 7930
rect 576 7910 594 7930
rect 545 7898 594 7910
rect 644 7934 688 7940
rect 644 7914 659 7934
rect 679 7914 688 7934
rect 644 7898 688 7914
rect 753 7930 802 7940
rect 753 7910 764 7930
rect 784 7910 802 7930
rect 753 7898 802 7910
rect 852 7934 896 7940
rect 852 7914 867 7934
rect 887 7914 896 7934
rect 852 7898 896 7914
rect 966 7934 1010 7940
rect 966 7914 975 7934
rect 995 7914 1010 7934
rect 966 7898 1010 7914
rect 1060 7930 1109 7940
rect 1060 7910 1078 7930
rect 1098 7910 1109 7930
rect 1060 7898 1109 7910
rect 2741 7901 2790 7913
rect 2741 7881 2752 7901
rect 2772 7881 2790 7901
rect 2741 7871 2790 7881
rect 2840 7897 2884 7913
rect 2840 7877 2855 7897
rect 2875 7877 2884 7897
rect 2840 7871 2884 7877
rect 2954 7897 2998 7913
rect 2954 7877 2963 7897
rect 2983 7877 2998 7897
rect 2954 7871 2998 7877
rect 3048 7901 3097 7913
rect 3048 7881 3066 7901
rect 3086 7881 3097 7901
rect 3048 7871 3097 7881
rect 3162 7897 3206 7913
rect 3162 7877 3171 7897
rect 3191 7877 3206 7897
rect 3162 7871 3206 7877
rect 3256 7901 3305 7913
rect 3256 7881 3274 7901
rect 3294 7881 3305 7901
rect 3256 7871 3305 7881
rect 3375 7897 3419 7913
rect 3375 7877 3384 7897
rect 3404 7877 3419 7897
rect 3375 7871 3419 7877
rect 3469 7901 3518 7913
rect 3469 7881 3487 7901
rect 3507 7881 3518 7901
rect 3469 7871 3518 7881
rect 1412 7648 1461 7658
rect 1412 7628 1423 7648
rect 1443 7628 1461 7648
rect 1412 7616 1461 7628
rect 1511 7652 1555 7658
rect 1511 7632 1526 7652
rect 1546 7632 1555 7652
rect 1511 7616 1555 7632
rect 1625 7648 1674 7658
rect 1625 7628 1636 7648
rect 1656 7628 1674 7648
rect 1625 7616 1674 7628
rect 1724 7652 1768 7658
rect 1724 7632 1739 7652
rect 1759 7632 1768 7652
rect 1724 7616 1768 7632
rect 1833 7648 1882 7658
rect 1833 7628 1844 7648
rect 1864 7628 1882 7648
rect 1833 7616 1882 7628
rect 1932 7652 1976 7658
rect 1932 7632 1947 7652
rect 1967 7632 1976 7652
rect 1932 7616 1976 7632
rect 2046 7652 2090 7658
rect 2046 7632 2055 7652
rect 2075 7632 2090 7652
rect 2046 7616 2090 7632
rect 2140 7648 2189 7658
rect 2140 7628 2158 7648
rect 2178 7628 2189 7648
rect 2140 7616 2189 7628
rect 3821 7619 3870 7631
rect 3821 7599 3832 7619
rect 3852 7599 3870 7619
rect 3821 7589 3870 7599
rect 3920 7615 3964 7631
rect 3920 7595 3935 7615
rect 3955 7595 3964 7615
rect 3920 7589 3964 7595
rect 4034 7615 4078 7631
rect 4034 7595 4043 7615
rect 4063 7595 4078 7615
rect 4034 7589 4078 7595
rect 4128 7619 4177 7631
rect 4128 7599 4146 7619
rect 4166 7599 4177 7619
rect 4128 7589 4177 7599
rect 4242 7615 4286 7631
rect 4242 7595 4251 7615
rect 4271 7595 4286 7615
rect 4242 7589 4286 7595
rect 4336 7619 4385 7631
rect 4336 7599 4354 7619
rect 4374 7599 4385 7619
rect 4336 7589 4385 7599
rect 4455 7615 4499 7631
rect 4455 7595 4464 7615
rect 4484 7595 4499 7615
rect 4455 7589 4499 7595
rect 4549 7619 4598 7631
rect 4549 7599 4567 7619
rect 4587 7599 4598 7619
rect 4549 7589 4598 7599
rect 334 7381 383 7391
rect 334 7361 345 7381
rect 365 7361 383 7381
rect 334 7349 383 7361
rect 433 7385 477 7391
rect 433 7365 448 7385
rect 468 7365 477 7385
rect 433 7349 477 7365
rect 547 7381 596 7391
rect 547 7361 558 7381
rect 578 7361 596 7381
rect 547 7349 596 7361
rect 646 7385 690 7391
rect 646 7365 661 7385
rect 681 7365 690 7385
rect 646 7349 690 7365
rect 755 7381 804 7391
rect 755 7361 766 7381
rect 786 7361 804 7381
rect 755 7349 804 7361
rect 854 7385 898 7391
rect 854 7365 869 7385
rect 889 7365 898 7385
rect 854 7349 898 7365
rect 968 7385 1012 7391
rect 968 7365 977 7385
rect 997 7365 1012 7385
rect 968 7349 1012 7365
rect 1062 7381 1111 7391
rect 1062 7361 1080 7381
rect 1100 7361 1111 7381
rect 1062 7349 1111 7361
rect 2882 7309 2931 7321
rect 2882 7289 2893 7309
rect 2913 7289 2931 7309
rect 2882 7279 2931 7289
rect 2981 7305 3025 7321
rect 2981 7285 2996 7305
rect 3016 7285 3025 7305
rect 2981 7279 3025 7285
rect 3095 7305 3139 7321
rect 3095 7285 3104 7305
rect 3124 7285 3139 7305
rect 3095 7279 3139 7285
rect 3189 7309 3238 7321
rect 3189 7289 3207 7309
rect 3227 7289 3238 7309
rect 3189 7279 3238 7289
rect 3303 7305 3347 7321
rect 3303 7285 3312 7305
rect 3332 7285 3347 7305
rect 3303 7279 3347 7285
rect 3397 7309 3446 7321
rect 3397 7289 3415 7309
rect 3435 7289 3446 7309
rect 3397 7279 3446 7289
rect 3516 7305 3560 7321
rect 3516 7285 3525 7305
rect 3545 7285 3560 7305
rect 3516 7279 3560 7285
rect 3610 7309 3659 7321
rect 3610 7289 3628 7309
rect 3648 7289 3659 7309
rect 3610 7279 3659 7289
rect 1272 7137 1321 7147
rect 1272 7117 1283 7137
rect 1303 7117 1321 7137
rect 1272 7105 1321 7117
rect 1371 7141 1415 7147
rect 1371 7121 1386 7141
rect 1406 7121 1415 7141
rect 1371 7105 1415 7121
rect 1485 7137 1534 7147
rect 1485 7117 1496 7137
rect 1516 7117 1534 7137
rect 1485 7105 1534 7117
rect 1584 7141 1628 7147
rect 1584 7121 1599 7141
rect 1619 7121 1628 7141
rect 1584 7105 1628 7121
rect 1693 7137 1742 7147
rect 1693 7117 1704 7137
rect 1724 7117 1742 7137
rect 1693 7105 1742 7117
rect 1792 7141 1836 7147
rect 1792 7121 1807 7141
rect 1827 7121 1836 7141
rect 1792 7105 1836 7121
rect 1906 7141 1950 7147
rect 1906 7121 1915 7141
rect 1935 7121 1950 7141
rect 1906 7105 1950 7121
rect 2000 7137 2049 7147
rect 2000 7117 2018 7137
rect 2038 7117 2049 7137
rect 2000 7105 2049 7117
rect 3820 7065 3869 7077
rect 3820 7045 3831 7065
rect 3851 7045 3869 7065
rect 3820 7035 3869 7045
rect 3919 7061 3963 7077
rect 3919 7041 3934 7061
rect 3954 7041 3963 7061
rect 3919 7035 3963 7041
rect 4033 7061 4077 7077
rect 4033 7041 4042 7061
rect 4062 7041 4077 7061
rect 4033 7035 4077 7041
rect 4127 7065 4176 7077
rect 4127 7045 4145 7065
rect 4165 7045 4176 7065
rect 4127 7035 4176 7045
rect 4241 7061 4285 7077
rect 4241 7041 4250 7061
rect 4270 7041 4285 7061
rect 4241 7035 4285 7041
rect 4335 7065 4384 7077
rect 4335 7045 4353 7065
rect 4373 7045 4384 7065
rect 4335 7035 4384 7045
rect 4454 7061 4498 7077
rect 4454 7041 4463 7061
rect 4483 7041 4498 7061
rect 4454 7035 4498 7041
rect 4548 7065 4597 7077
rect 4548 7045 4566 7065
rect 4586 7045 4597 7065
rect 4548 7035 4597 7045
rect 333 6827 382 6837
rect 333 6807 344 6827
rect 364 6807 382 6827
rect 333 6795 382 6807
rect 432 6831 476 6837
rect 432 6811 447 6831
rect 467 6811 476 6831
rect 432 6795 476 6811
rect 546 6827 595 6837
rect 546 6807 557 6827
rect 577 6807 595 6827
rect 546 6795 595 6807
rect 645 6831 689 6837
rect 645 6811 660 6831
rect 680 6811 689 6831
rect 645 6795 689 6811
rect 754 6827 803 6837
rect 754 6807 765 6827
rect 785 6807 803 6827
rect 754 6795 803 6807
rect 853 6831 897 6837
rect 853 6811 868 6831
rect 888 6811 897 6831
rect 853 6795 897 6811
rect 967 6831 1011 6837
rect 967 6811 976 6831
rect 996 6811 1011 6831
rect 967 6795 1011 6811
rect 1061 6827 1110 6837
rect 1061 6807 1079 6827
rect 1099 6807 1110 6827
rect 1061 6795 1110 6807
rect 2772 6785 2821 6797
rect 2772 6765 2783 6785
rect 2803 6765 2821 6785
rect 2772 6755 2821 6765
rect 2871 6781 2915 6797
rect 2871 6761 2886 6781
rect 2906 6761 2915 6781
rect 2871 6755 2915 6761
rect 2985 6781 3029 6797
rect 2985 6761 2994 6781
rect 3014 6761 3029 6781
rect 2985 6755 3029 6761
rect 3079 6785 3128 6797
rect 3079 6765 3097 6785
rect 3117 6765 3128 6785
rect 3079 6755 3128 6765
rect 3193 6781 3237 6797
rect 3193 6761 3202 6781
rect 3222 6761 3237 6781
rect 3193 6755 3237 6761
rect 3287 6785 3336 6797
rect 3287 6765 3305 6785
rect 3325 6765 3336 6785
rect 3287 6755 3336 6765
rect 3406 6781 3450 6797
rect 3406 6761 3415 6781
rect 3435 6761 3450 6781
rect 3406 6755 3450 6761
rect 3500 6785 3549 6797
rect 3500 6765 3518 6785
rect 3538 6765 3549 6785
rect 3500 6755 3549 6765
rect 1382 6558 1431 6568
rect 1382 6538 1393 6558
rect 1413 6538 1431 6558
rect 1382 6526 1431 6538
rect 1481 6562 1525 6568
rect 1481 6542 1496 6562
rect 1516 6542 1525 6562
rect 1481 6526 1525 6542
rect 1595 6558 1644 6568
rect 1595 6538 1606 6558
rect 1626 6538 1644 6558
rect 1595 6526 1644 6538
rect 1694 6562 1738 6568
rect 1694 6542 1709 6562
rect 1729 6542 1738 6562
rect 1694 6526 1738 6542
rect 1803 6558 1852 6568
rect 1803 6538 1814 6558
rect 1834 6538 1852 6558
rect 1803 6526 1852 6538
rect 1902 6562 1946 6568
rect 1902 6542 1917 6562
rect 1937 6542 1946 6562
rect 1902 6526 1946 6542
rect 2016 6562 2060 6568
rect 2016 6542 2025 6562
rect 2045 6542 2060 6562
rect 2016 6526 2060 6542
rect 2110 6558 2159 6568
rect 2110 6538 2128 6558
rect 2148 6538 2159 6558
rect 2110 6526 2159 6538
rect 3821 6516 3870 6528
rect 3821 6496 3832 6516
rect 3852 6496 3870 6516
rect 3821 6486 3870 6496
rect 3920 6512 3964 6528
rect 3920 6492 3935 6512
rect 3955 6492 3964 6512
rect 3920 6486 3964 6492
rect 4034 6512 4078 6528
rect 4034 6492 4043 6512
rect 4063 6492 4078 6512
rect 4034 6486 4078 6492
rect 4128 6516 4177 6528
rect 4128 6496 4146 6516
rect 4166 6496 4177 6516
rect 4128 6486 4177 6496
rect 4242 6512 4286 6528
rect 4242 6492 4251 6512
rect 4271 6492 4286 6512
rect 4242 6486 4286 6492
rect 4336 6516 4385 6528
rect 4336 6496 4354 6516
rect 4374 6496 4385 6516
rect 4336 6486 4385 6496
rect 4455 6512 4499 6528
rect 4455 6492 4464 6512
rect 4484 6492 4499 6512
rect 4455 6486 4499 6492
rect 4549 6516 4598 6528
rect 4549 6496 4567 6516
rect 4587 6496 4598 6516
rect 4549 6486 4598 6496
rect 334 6278 383 6288
rect 334 6258 345 6278
rect 365 6258 383 6278
rect 334 6246 383 6258
rect 433 6282 477 6288
rect 433 6262 448 6282
rect 468 6262 477 6282
rect 433 6246 477 6262
rect 547 6278 596 6288
rect 547 6258 558 6278
rect 578 6258 596 6278
rect 547 6246 596 6258
rect 646 6282 690 6288
rect 646 6262 661 6282
rect 681 6262 690 6282
rect 646 6246 690 6262
rect 755 6278 804 6288
rect 755 6258 766 6278
rect 786 6258 804 6278
rect 755 6246 804 6258
rect 854 6282 898 6288
rect 854 6262 869 6282
rect 889 6262 898 6282
rect 854 6246 898 6262
rect 968 6282 1012 6288
rect 968 6262 977 6282
rect 997 6262 1012 6282
rect 968 6246 1012 6262
rect 1062 6278 1111 6288
rect 1062 6258 1080 6278
rect 1100 6258 1111 6278
rect 1062 6246 1111 6258
rect 2882 6206 2931 6218
rect 2882 6186 2893 6206
rect 2913 6186 2931 6206
rect 2882 6176 2931 6186
rect 2981 6202 3025 6218
rect 2981 6182 2996 6202
rect 3016 6182 3025 6202
rect 2981 6176 3025 6182
rect 3095 6202 3139 6218
rect 3095 6182 3104 6202
rect 3124 6182 3139 6202
rect 3095 6176 3139 6182
rect 3189 6206 3238 6218
rect 3189 6186 3207 6206
rect 3227 6186 3238 6206
rect 3189 6176 3238 6186
rect 3303 6202 3347 6218
rect 3303 6182 3312 6202
rect 3332 6182 3347 6202
rect 3303 6176 3347 6182
rect 3397 6206 3446 6218
rect 3397 6186 3415 6206
rect 3435 6186 3446 6206
rect 3397 6176 3446 6186
rect 3516 6202 3560 6218
rect 3516 6182 3525 6202
rect 3545 6182 3560 6202
rect 3516 6176 3560 6182
rect 3610 6206 3659 6218
rect 3610 6186 3628 6206
rect 3648 6186 3659 6206
rect 3610 6176 3659 6186
rect 1272 6034 1321 6044
rect 1272 6014 1283 6034
rect 1303 6014 1321 6034
rect 1272 6002 1321 6014
rect 1371 6038 1415 6044
rect 1371 6018 1386 6038
rect 1406 6018 1415 6038
rect 1371 6002 1415 6018
rect 1485 6034 1534 6044
rect 1485 6014 1496 6034
rect 1516 6014 1534 6034
rect 1485 6002 1534 6014
rect 1584 6038 1628 6044
rect 1584 6018 1599 6038
rect 1619 6018 1628 6038
rect 1584 6002 1628 6018
rect 1693 6034 1742 6044
rect 1693 6014 1704 6034
rect 1724 6014 1742 6034
rect 1693 6002 1742 6014
rect 1792 6038 1836 6044
rect 1792 6018 1807 6038
rect 1827 6018 1836 6038
rect 1792 6002 1836 6018
rect 1906 6038 1950 6044
rect 1906 6018 1915 6038
rect 1935 6018 1950 6038
rect 1906 6002 1950 6018
rect 2000 6034 2049 6044
rect 2000 6014 2018 6034
rect 2038 6014 2049 6034
rect 2000 6002 2049 6014
rect 3820 5962 3869 5974
rect 3820 5942 3831 5962
rect 3851 5942 3869 5962
rect 3820 5932 3869 5942
rect 3919 5958 3963 5974
rect 3919 5938 3934 5958
rect 3954 5938 3963 5958
rect 3919 5932 3963 5938
rect 4033 5958 4077 5974
rect 4033 5938 4042 5958
rect 4062 5938 4077 5958
rect 4033 5932 4077 5938
rect 4127 5962 4176 5974
rect 4127 5942 4145 5962
rect 4165 5942 4176 5962
rect 4127 5932 4176 5942
rect 4241 5958 4285 5974
rect 4241 5938 4250 5958
rect 4270 5938 4285 5958
rect 4241 5932 4285 5938
rect 4335 5962 4384 5974
rect 4335 5942 4353 5962
rect 4373 5942 4384 5962
rect 4335 5932 4384 5942
rect 4454 5958 4498 5974
rect 4454 5938 4463 5958
rect 4483 5938 4498 5958
rect 4454 5932 4498 5938
rect 4548 5962 4597 5974
rect 4548 5942 4566 5962
rect 4586 5942 4597 5962
rect 4548 5932 4597 5942
rect 333 5724 382 5734
rect 333 5704 344 5724
rect 364 5704 382 5724
rect 333 5692 382 5704
rect 432 5728 476 5734
rect 432 5708 447 5728
rect 467 5708 476 5728
rect 432 5692 476 5708
rect 546 5724 595 5734
rect 546 5704 557 5724
rect 577 5704 595 5724
rect 546 5692 595 5704
rect 645 5728 689 5734
rect 645 5708 660 5728
rect 680 5708 689 5728
rect 645 5692 689 5708
rect 754 5724 803 5734
rect 754 5704 765 5724
rect 785 5704 803 5724
rect 754 5692 803 5704
rect 853 5728 897 5734
rect 853 5708 868 5728
rect 888 5708 897 5728
rect 853 5692 897 5708
rect 967 5728 1011 5734
rect 967 5708 976 5728
rect 996 5708 1011 5728
rect 967 5692 1011 5708
rect 1061 5724 1110 5734
rect 1061 5704 1079 5724
rect 1099 5704 1110 5724
rect 1061 5692 1110 5704
rect 2742 5695 2791 5707
rect 2742 5675 2753 5695
rect 2773 5675 2791 5695
rect 2742 5665 2791 5675
rect 2841 5691 2885 5707
rect 2841 5671 2856 5691
rect 2876 5671 2885 5691
rect 2841 5665 2885 5671
rect 2955 5691 2999 5707
rect 2955 5671 2964 5691
rect 2984 5671 2999 5691
rect 2955 5665 2999 5671
rect 3049 5695 3098 5707
rect 3049 5675 3067 5695
rect 3087 5675 3098 5695
rect 3049 5665 3098 5675
rect 3163 5691 3207 5707
rect 3163 5671 3172 5691
rect 3192 5671 3207 5691
rect 3163 5665 3207 5671
rect 3257 5695 3306 5707
rect 3257 5675 3275 5695
rect 3295 5675 3306 5695
rect 3257 5665 3306 5675
rect 3376 5691 3420 5707
rect 3376 5671 3385 5691
rect 3405 5671 3420 5691
rect 3376 5665 3420 5671
rect 3470 5695 3519 5707
rect 3470 5675 3488 5695
rect 3508 5675 3519 5695
rect 3470 5665 3519 5675
rect 1413 5442 1462 5452
rect 1413 5422 1424 5442
rect 1444 5422 1462 5442
rect 1413 5410 1462 5422
rect 1512 5446 1556 5452
rect 1512 5426 1527 5446
rect 1547 5426 1556 5446
rect 1512 5410 1556 5426
rect 1626 5442 1675 5452
rect 1626 5422 1637 5442
rect 1657 5422 1675 5442
rect 1626 5410 1675 5422
rect 1725 5446 1769 5452
rect 1725 5426 1740 5446
rect 1760 5426 1769 5446
rect 1725 5410 1769 5426
rect 1834 5442 1883 5452
rect 1834 5422 1845 5442
rect 1865 5422 1883 5442
rect 1834 5410 1883 5422
rect 1933 5446 1977 5452
rect 1933 5426 1948 5446
rect 1968 5426 1977 5446
rect 1933 5410 1977 5426
rect 2047 5446 2091 5452
rect 2047 5426 2056 5446
rect 2076 5426 2091 5446
rect 2047 5410 2091 5426
rect 2141 5442 2190 5452
rect 2141 5422 2159 5442
rect 2179 5422 2190 5442
rect 2141 5410 2190 5422
rect 3822 5413 3871 5425
rect 3822 5393 3833 5413
rect 3853 5393 3871 5413
rect 3822 5383 3871 5393
rect 3921 5409 3965 5425
rect 3921 5389 3936 5409
rect 3956 5389 3965 5409
rect 3921 5383 3965 5389
rect 4035 5409 4079 5425
rect 4035 5389 4044 5409
rect 4064 5389 4079 5409
rect 4035 5383 4079 5389
rect 4129 5413 4178 5425
rect 4129 5393 4147 5413
rect 4167 5393 4178 5413
rect 4129 5383 4178 5393
rect 4243 5409 4287 5425
rect 4243 5389 4252 5409
rect 4272 5389 4287 5409
rect 4243 5383 4287 5389
rect 4337 5413 4386 5425
rect 4337 5393 4355 5413
rect 4375 5393 4386 5413
rect 4337 5383 4386 5393
rect 4456 5409 4500 5425
rect 4456 5389 4465 5409
rect 4485 5389 4500 5409
rect 4456 5383 4500 5389
rect 4550 5413 4599 5425
rect 4550 5393 4568 5413
rect 4588 5393 4599 5413
rect 4550 5383 4599 5393
rect 335 5175 384 5185
rect 335 5155 346 5175
rect 366 5155 384 5175
rect 335 5143 384 5155
rect 434 5179 478 5185
rect 434 5159 449 5179
rect 469 5159 478 5179
rect 434 5143 478 5159
rect 548 5175 597 5185
rect 548 5155 559 5175
rect 579 5155 597 5175
rect 548 5143 597 5155
rect 647 5179 691 5185
rect 647 5159 662 5179
rect 682 5159 691 5179
rect 647 5143 691 5159
rect 756 5175 805 5185
rect 756 5155 767 5175
rect 787 5155 805 5175
rect 756 5143 805 5155
rect 855 5179 899 5185
rect 855 5159 870 5179
rect 890 5159 899 5179
rect 855 5143 899 5159
rect 969 5179 1013 5185
rect 969 5159 978 5179
rect 998 5159 1013 5179
rect 969 5143 1013 5159
rect 1063 5175 1112 5185
rect 1063 5155 1081 5175
rect 1101 5155 1112 5175
rect 1063 5143 1112 5155
rect 2883 5103 2932 5115
rect 2883 5083 2894 5103
rect 2914 5083 2932 5103
rect 2883 5073 2932 5083
rect 2982 5099 3026 5115
rect 2982 5079 2997 5099
rect 3017 5079 3026 5099
rect 2982 5073 3026 5079
rect 3096 5099 3140 5115
rect 3096 5079 3105 5099
rect 3125 5079 3140 5099
rect 3096 5073 3140 5079
rect 3190 5103 3239 5115
rect 3190 5083 3208 5103
rect 3228 5083 3239 5103
rect 3190 5073 3239 5083
rect 3304 5099 3348 5115
rect 3304 5079 3313 5099
rect 3333 5079 3348 5099
rect 3304 5073 3348 5079
rect 3398 5103 3447 5115
rect 3398 5083 3416 5103
rect 3436 5083 3447 5103
rect 3398 5073 3447 5083
rect 3517 5099 3561 5115
rect 3517 5079 3526 5099
rect 3546 5079 3561 5099
rect 3517 5073 3561 5079
rect 3611 5103 3660 5115
rect 3611 5083 3629 5103
rect 3649 5083 3660 5103
rect 3611 5073 3660 5083
rect 1273 4931 1322 4941
rect 1273 4911 1284 4931
rect 1304 4911 1322 4931
rect 1273 4899 1322 4911
rect 1372 4935 1416 4941
rect 1372 4915 1387 4935
rect 1407 4915 1416 4935
rect 1372 4899 1416 4915
rect 1486 4931 1535 4941
rect 1486 4911 1497 4931
rect 1517 4911 1535 4931
rect 1486 4899 1535 4911
rect 1585 4935 1629 4941
rect 1585 4915 1600 4935
rect 1620 4915 1629 4935
rect 1585 4899 1629 4915
rect 1694 4931 1743 4941
rect 1694 4911 1705 4931
rect 1725 4911 1743 4931
rect 1694 4899 1743 4911
rect 1793 4935 1837 4941
rect 1793 4915 1808 4935
rect 1828 4915 1837 4935
rect 1793 4899 1837 4915
rect 1907 4935 1951 4941
rect 1907 4915 1916 4935
rect 1936 4915 1951 4935
rect 1907 4899 1951 4915
rect 2001 4931 2050 4941
rect 2001 4911 2019 4931
rect 2039 4911 2050 4931
rect 2001 4899 2050 4911
rect 3821 4859 3870 4871
rect 3821 4839 3832 4859
rect 3852 4839 3870 4859
rect 3821 4829 3870 4839
rect 3920 4855 3964 4871
rect 3920 4835 3935 4855
rect 3955 4835 3964 4855
rect 3920 4829 3964 4835
rect 4034 4855 4078 4871
rect 4034 4835 4043 4855
rect 4063 4835 4078 4855
rect 4034 4829 4078 4835
rect 4128 4859 4177 4871
rect 4128 4839 4146 4859
rect 4166 4839 4177 4859
rect 4128 4829 4177 4839
rect 4242 4855 4286 4871
rect 4242 4835 4251 4855
rect 4271 4835 4286 4855
rect 4242 4829 4286 4835
rect 4336 4859 4385 4871
rect 4336 4839 4354 4859
rect 4374 4839 4385 4859
rect 4336 4829 4385 4839
rect 4455 4855 4499 4871
rect 4455 4835 4464 4855
rect 4484 4835 4499 4855
rect 4455 4829 4499 4835
rect 4549 4859 4598 4871
rect 4549 4839 4567 4859
rect 4587 4839 4598 4859
rect 4549 4829 4598 4839
rect 334 4621 383 4631
rect 334 4601 345 4621
rect 365 4601 383 4621
rect 334 4589 383 4601
rect 433 4625 477 4631
rect 433 4605 448 4625
rect 468 4605 477 4625
rect 433 4589 477 4605
rect 547 4621 596 4631
rect 547 4601 558 4621
rect 578 4601 596 4621
rect 547 4589 596 4601
rect 646 4625 690 4631
rect 646 4605 661 4625
rect 681 4605 690 4625
rect 646 4589 690 4605
rect 755 4621 804 4631
rect 755 4601 766 4621
rect 786 4601 804 4621
rect 755 4589 804 4601
rect 854 4625 898 4631
rect 854 4605 869 4625
rect 889 4605 898 4625
rect 854 4589 898 4605
rect 968 4625 1012 4631
rect 968 4605 977 4625
rect 997 4605 1012 4625
rect 968 4589 1012 4605
rect 1062 4621 1111 4631
rect 1062 4601 1080 4621
rect 1100 4601 1111 4621
rect 1062 4589 1111 4601
rect 2774 4573 2823 4585
rect 2774 4553 2785 4573
rect 2805 4553 2823 4573
rect 2774 4543 2823 4553
rect 2873 4569 2917 4585
rect 2873 4549 2888 4569
rect 2908 4549 2917 4569
rect 2873 4543 2917 4549
rect 2987 4569 3031 4585
rect 2987 4549 2996 4569
rect 3016 4549 3031 4569
rect 2987 4543 3031 4549
rect 3081 4573 3130 4585
rect 3081 4553 3099 4573
rect 3119 4553 3130 4573
rect 3081 4543 3130 4553
rect 3195 4569 3239 4585
rect 3195 4549 3204 4569
rect 3224 4549 3239 4569
rect 3195 4543 3239 4549
rect 3289 4573 3338 4585
rect 3289 4553 3307 4573
rect 3327 4553 3338 4573
rect 3289 4543 3338 4553
rect 3408 4569 3452 4585
rect 3408 4549 3417 4569
rect 3437 4549 3452 4569
rect 3408 4543 3452 4549
rect 3502 4573 3551 4585
rect 3502 4553 3520 4573
rect 3540 4553 3551 4573
rect 3502 4543 3551 4553
rect 1382 4358 1431 4368
rect 1382 4338 1393 4358
rect 1413 4338 1431 4358
rect 1382 4326 1431 4338
rect 1481 4362 1525 4368
rect 1481 4342 1496 4362
rect 1516 4342 1525 4362
rect 1481 4326 1525 4342
rect 1595 4358 1644 4368
rect 1595 4338 1606 4358
rect 1626 4338 1644 4358
rect 1595 4326 1644 4338
rect 1694 4362 1738 4368
rect 1694 4342 1709 4362
rect 1729 4342 1738 4362
rect 1694 4326 1738 4342
rect 1803 4358 1852 4368
rect 1803 4338 1814 4358
rect 1834 4338 1852 4358
rect 1803 4326 1852 4338
rect 1902 4362 1946 4368
rect 1902 4342 1917 4362
rect 1937 4342 1946 4362
rect 1902 4326 1946 4342
rect 2016 4362 2060 4368
rect 2016 4342 2025 4362
rect 2045 4342 2060 4362
rect 2016 4326 2060 4342
rect 2110 4358 2159 4368
rect 2110 4338 2128 4358
rect 2148 4338 2159 4358
rect 2110 4326 2159 4338
rect 3822 4310 3871 4322
rect 3822 4290 3833 4310
rect 3853 4290 3871 4310
rect 3822 4280 3871 4290
rect 3921 4306 3965 4322
rect 3921 4286 3936 4306
rect 3956 4286 3965 4306
rect 3921 4280 3965 4286
rect 4035 4306 4079 4322
rect 4035 4286 4044 4306
rect 4064 4286 4079 4306
rect 4035 4280 4079 4286
rect 4129 4310 4178 4322
rect 4129 4290 4147 4310
rect 4167 4290 4178 4310
rect 4129 4280 4178 4290
rect 4243 4306 4287 4322
rect 4243 4286 4252 4306
rect 4272 4286 4287 4306
rect 4243 4280 4287 4286
rect 4337 4310 4386 4322
rect 4337 4290 4355 4310
rect 4375 4290 4386 4310
rect 4337 4280 4386 4290
rect 4456 4306 4500 4322
rect 4456 4286 4465 4306
rect 4485 4286 4500 4306
rect 4456 4280 4500 4286
rect 4550 4310 4599 4322
rect 4550 4290 4568 4310
rect 4588 4290 4599 4310
rect 4550 4280 4599 4290
rect 335 4072 384 4082
rect 335 4052 346 4072
rect 366 4052 384 4072
rect 335 4040 384 4052
rect 434 4076 478 4082
rect 434 4056 449 4076
rect 469 4056 478 4076
rect 434 4040 478 4056
rect 548 4072 597 4082
rect 548 4052 559 4072
rect 579 4052 597 4072
rect 548 4040 597 4052
rect 647 4076 691 4082
rect 647 4056 662 4076
rect 682 4056 691 4076
rect 647 4040 691 4056
rect 756 4072 805 4082
rect 756 4052 767 4072
rect 787 4052 805 4072
rect 756 4040 805 4052
rect 855 4076 899 4082
rect 855 4056 870 4076
rect 890 4056 899 4076
rect 855 4040 899 4056
rect 969 4076 1013 4082
rect 969 4056 978 4076
rect 998 4056 1013 4076
rect 969 4040 1013 4056
rect 1063 4072 1112 4082
rect 1063 4052 1081 4072
rect 1101 4052 1112 4072
rect 1063 4040 1112 4052
rect 2883 4000 2932 4012
rect 2883 3980 2894 4000
rect 2914 3980 2932 4000
rect 2883 3970 2932 3980
rect 2982 3996 3026 4012
rect 2982 3976 2997 3996
rect 3017 3976 3026 3996
rect 2982 3970 3026 3976
rect 3096 3996 3140 4012
rect 3096 3976 3105 3996
rect 3125 3976 3140 3996
rect 3096 3970 3140 3976
rect 3190 4000 3239 4012
rect 3190 3980 3208 4000
rect 3228 3980 3239 4000
rect 3190 3970 3239 3980
rect 3304 3996 3348 4012
rect 3304 3976 3313 3996
rect 3333 3976 3348 3996
rect 3304 3970 3348 3976
rect 3398 4000 3447 4012
rect 3398 3980 3416 4000
rect 3436 3980 3447 4000
rect 3398 3970 3447 3980
rect 3517 3996 3561 4012
rect 3517 3976 3526 3996
rect 3546 3976 3561 3996
rect 3517 3970 3561 3976
rect 3611 4000 3660 4012
rect 3611 3980 3629 4000
rect 3649 3980 3660 4000
rect 3611 3970 3660 3980
rect 1273 3828 1322 3838
rect 1273 3808 1284 3828
rect 1304 3808 1322 3828
rect 1273 3796 1322 3808
rect 1372 3832 1416 3838
rect 1372 3812 1387 3832
rect 1407 3812 1416 3832
rect 1372 3796 1416 3812
rect 1486 3828 1535 3838
rect 1486 3808 1497 3828
rect 1517 3808 1535 3828
rect 1486 3796 1535 3808
rect 1585 3832 1629 3838
rect 1585 3812 1600 3832
rect 1620 3812 1629 3832
rect 1585 3796 1629 3812
rect 1694 3828 1743 3838
rect 1694 3808 1705 3828
rect 1725 3808 1743 3828
rect 1694 3796 1743 3808
rect 1793 3832 1837 3838
rect 1793 3812 1808 3832
rect 1828 3812 1837 3832
rect 1793 3796 1837 3812
rect 1907 3832 1951 3838
rect 1907 3812 1916 3832
rect 1936 3812 1951 3832
rect 1907 3796 1951 3812
rect 2001 3828 2050 3838
rect 2001 3808 2019 3828
rect 2039 3808 2050 3828
rect 2001 3796 2050 3808
rect 3821 3756 3870 3768
rect 3821 3736 3832 3756
rect 3852 3736 3870 3756
rect 3821 3726 3870 3736
rect 3920 3752 3964 3768
rect 3920 3732 3935 3752
rect 3955 3732 3964 3752
rect 3920 3726 3964 3732
rect 4034 3752 4078 3768
rect 4034 3732 4043 3752
rect 4063 3732 4078 3752
rect 4034 3726 4078 3732
rect 4128 3756 4177 3768
rect 4128 3736 4146 3756
rect 4166 3736 4177 3756
rect 4128 3726 4177 3736
rect 4242 3752 4286 3768
rect 4242 3732 4251 3752
rect 4271 3732 4286 3752
rect 4242 3726 4286 3732
rect 4336 3756 4385 3768
rect 4336 3736 4354 3756
rect 4374 3736 4385 3756
rect 4336 3726 4385 3736
rect 4455 3752 4499 3768
rect 4455 3732 4464 3752
rect 4484 3732 4499 3752
rect 4455 3726 4499 3732
rect 4549 3756 4598 3768
rect 4549 3736 4567 3756
rect 4587 3736 4598 3756
rect 4549 3726 4598 3736
rect 334 3518 383 3528
rect 334 3498 345 3518
rect 365 3498 383 3518
rect 334 3486 383 3498
rect 433 3522 477 3528
rect 433 3502 448 3522
rect 468 3502 477 3522
rect 433 3486 477 3502
rect 547 3518 596 3528
rect 547 3498 558 3518
rect 578 3498 596 3518
rect 547 3486 596 3498
rect 646 3522 690 3528
rect 646 3502 661 3522
rect 681 3502 690 3522
rect 646 3486 690 3502
rect 755 3518 804 3528
rect 755 3498 766 3518
rect 786 3498 804 3518
rect 755 3486 804 3498
rect 854 3522 898 3528
rect 854 3502 869 3522
rect 889 3502 898 3522
rect 854 3486 898 3502
rect 968 3522 1012 3528
rect 968 3502 977 3522
rect 997 3502 1012 3522
rect 968 3486 1012 3502
rect 1062 3518 1111 3528
rect 1062 3498 1080 3518
rect 1100 3498 1111 3518
rect 1062 3486 1111 3498
rect 2743 3489 2792 3501
rect 2743 3469 2754 3489
rect 2774 3469 2792 3489
rect 2743 3459 2792 3469
rect 2842 3485 2886 3501
rect 2842 3465 2857 3485
rect 2877 3465 2886 3485
rect 2842 3459 2886 3465
rect 2956 3485 3000 3501
rect 2956 3465 2965 3485
rect 2985 3465 3000 3485
rect 2956 3459 3000 3465
rect 3050 3489 3099 3501
rect 3050 3469 3068 3489
rect 3088 3469 3099 3489
rect 3050 3459 3099 3469
rect 3164 3485 3208 3501
rect 3164 3465 3173 3485
rect 3193 3465 3208 3485
rect 3164 3459 3208 3465
rect 3258 3489 3307 3501
rect 3258 3469 3276 3489
rect 3296 3469 3307 3489
rect 3258 3459 3307 3469
rect 3377 3485 3421 3501
rect 3377 3465 3386 3485
rect 3406 3465 3421 3485
rect 3377 3459 3421 3465
rect 3471 3489 3520 3501
rect 3471 3469 3489 3489
rect 3509 3469 3520 3489
rect 3471 3459 3520 3469
rect 1414 3236 1463 3246
rect 1414 3216 1425 3236
rect 1445 3216 1463 3236
rect 1414 3204 1463 3216
rect 1513 3240 1557 3246
rect 1513 3220 1528 3240
rect 1548 3220 1557 3240
rect 1513 3204 1557 3220
rect 1627 3236 1676 3246
rect 1627 3216 1638 3236
rect 1658 3216 1676 3236
rect 1627 3204 1676 3216
rect 1726 3240 1770 3246
rect 1726 3220 1741 3240
rect 1761 3220 1770 3240
rect 1726 3204 1770 3220
rect 1835 3236 1884 3246
rect 1835 3216 1846 3236
rect 1866 3216 1884 3236
rect 1835 3204 1884 3216
rect 1934 3240 1978 3246
rect 1934 3220 1949 3240
rect 1969 3220 1978 3240
rect 1934 3204 1978 3220
rect 2048 3240 2092 3246
rect 2048 3220 2057 3240
rect 2077 3220 2092 3240
rect 2048 3204 2092 3220
rect 2142 3236 2191 3246
rect 2142 3216 2160 3236
rect 2180 3216 2191 3236
rect 2142 3204 2191 3216
rect 3823 3207 3872 3219
rect 3823 3187 3834 3207
rect 3854 3187 3872 3207
rect 3823 3177 3872 3187
rect 3922 3203 3966 3219
rect 3922 3183 3937 3203
rect 3957 3183 3966 3203
rect 3922 3177 3966 3183
rect 4036 3203 4080 3219
rect 4036 3183 4045 3203
rect 4065 3183 4080 3203
rect 4036 3177 4080 3183
rect 4130 3207 4179 3219
rect 4130 3187 4148 3207
rect 4168 3187 4179 3207
rect 4130 3177 4179 3187
rect 4244 3203 4288 3219
rect 4244 3183 4253 3203
rect 4273 3183 4288 3203
rect 4244 3177 4288 3183
rect 4338 3207 4387 3219
rect 4338 3187 4356 3207
rect 4376 3187 4387 3207
rect 4338 3177 4387 3187
rect 4457 3203 4501 3219
rect 4457 3183 4466 3203
rect 4486 3183 4501 3203
rect 4457 3177 4501 3183
rect 4551 3207 4600 3219
rect 4551 3187 4569 3207
rect 4589 3187 4600 3207
rect 4551 3177 4600 3187
rect 336 2969 385 2979
rect 336 2949 347 2969
rect 367 2949 385 2969
rect 336 2937 385 2949
rect 435 2973 479 2979
rect 435 2953 450 2973
rect 470 2953 479 2973
rect 435 2937 479 2953
rect 549 2969 598 2979
rect 549 2949 560 2969
rect 580 2949 598 2969
rect 549 2937 598 2949
rect 648 2973 692 2979
rect 648 2953 663 2973
rect 683 2953 692 2973
rect 648 2937 692 2953
rect 757 2969 806 2979
rect 757 2949 768 2969
rect 788 2949 806 2969
rect 757 2937 806 2949
rect 856 2973 900 2979
rect 856 2953 871 2973
rect 891 2953 900 2973
rect 856 2937 900 2953
rect 970 2973 1014 2979
rect 970 2953 979 2973
rect 999 2953 1014 2973
rect 970 2937 1014 2953
rect 1064 2969 1113 2979
rect 1064 2949 1082 2969
rect 1102 2949 1113 2969
rect 1064 2937 1113 2949
rect 2884 2897 2933 2909
rect 2884 2877 2895 2897
rect 2915 2877 2933 2897
rect 2884 2867 2933 2877
rect 2983 2893 3027 2909
rect 2983 2873 2998 2893
rect 3018 2873 3027 2893
rect 2983 2867 3027 2873
rect 3097 2893 3141 2909
rect 3097 2873 3106 2893
rect 3126 2873 3141 2893
rect 3097 2867 3141 2873
rect 3191 2897 3240 2909
rect 3191 2877 3209 2897
rect 3229 2877 3240 2897
rect 3191 2867 3240 2877
rect 3305 2893 3349 2909
rect 3305 2873 3314 2893
rect 3334 2873 3349 2893
rect 3305 2867 3349 2873
rect 3399 2897 3448 2909
rect 3399 2877 3417 2897
rect 3437 2877 3448 2897
rect 3399 2867 3448 2877
rect 3518 2893 3562 2909
rect 3518 2873 3527 2893
rect 3547 2873 3562 2893
rect 3518 2867 3562 2873
rect 3612 2897 3661 2909
rect 3612 2877 3630 2897
rect 3650 2877 3661 2897
rect 3612 2867 3661 2877
rect 1274 2725 1323 2735
rect 1274 2705 1285 2725
rect 1305 2705 1323 2725
rect 1274 2693 1323 2705
rect 1373 2729 1417 2735
rect 1373 2709 1388 2729
rect 1408 2709 1417 2729
rect 1373 2693 1417 2709
rect 1487 2725 1536 2735
rect 1487 2705 1498 2725
rect 1518 2705 1536 2725
rect 1487 2693 1536 2705
rect 1586 2729 1630 2735
rect 1586 2709 1601 2729
rect 1621 2709 1630 2729
rect 1586 2693 1630 2709
rect 1695 2725 1744 2735
rect 1695 2705 1706 2725
rect 1726 2705 1744 2725
rect 1695 2693 1744 2705
rect 1794 2729 1838 2735
rect 1794 2709 1809 2729
rect 1829 2709 1838 2729
rect 1794 2693 1838 2709
rect 1908 2729 1952 2735
rect 1908 2709 1917 2729
rect 1937 2709 1952 2729
rect 1908 2693 1952 2709
rect 2002 2725 2051 2735
rect 2002 2705 2020 2725
rect 2040 2705 2051 2725
rect 2002 2693 2051 2705
rect 3822 2653 3871 2665
rect 3822 2633 3833 2653
rect 3853 2633 3871 2653
rect 3822 2623 3871 2633
rect 3921 2649 3965 2665
rect 3921 2629 3936 2649
rect 3956 2629 3965 2649
rect 3921 2623 3965 2629
rect 4035 2649 4079 2665
rect 4035 2629 4044 2649
rect 4064 2629 4079 2649
rect 4035 2623 4079 2629
rect 4129 2653 4178 2665
rect 4129 2633 4147 2653
rect 4167 2633 4178 2653
rect 4129 2623 4178 2633
rect 4243 2649 4287 2665
rect 4243 2629 4252 2649
rect 4272 2629 4287 2649
rect 4243 2623 4287 2629
rect 4337 2653 4386 2665
rect 4337 2633 4355 2653
rect 4375 2633 4386 2653
rect 4337 2623 4386 2633
rect 4456 2649 4500 2665
rect 4456 2629 4465 2649
rect 4485 2629 4500 2649
rect 4456 2623 4500 2629
rect 4550 2653 4599 2665
rect 4550 2633 4568 2653
rect 4588 2633 4599 2653
rect 4550 2623 4599 2633
rect 335 2415 384 2425
rect 335 2395 346 2415
rect 366 2395 384 2415
rect 335 2383 384 2395
rect 434 2419 478 2425
rect 434 2399 449 2419
rect 469 2399 478 2419
rect 434 2383 478 2399
rect 548 2415 597 2425
rect 548 2395 559 2415
rect 579 2395 597 2415
rect 548 2383 597 2395
rect 647 2419 691 2425
rect 647 2399 662 2419
rect 682 2399 691 2419
rect 647 2383 691 2399
rect 756 2415 805 2425
rect 756 2395 767 2415
rect 787 2395 805 2415
rect 756 2383 805 2395
rect 855 2419 899 2425
rect 855 2399 870 2419
rect 890 2399 899 2419
rect 855 2383 899 2399
rect 969 2419 1013 2425
rect 969 2399 978 2419
rect 998 2399 1013 2419
rect 969 2383 1013 2399
rect 1063 2415 1112 2425
rect 1063 2395 1081 2415
rect 1101 2395 1112 2415
rect 1063 2383 1112 2395
rect 2774 2373 2823 2385
rect 2774 2353 2785 2373
rect 2805 2353 2823 2373
rect 2774 2343 2823 2353
rect 2873 2369 2917 2385
rect 2873 2349 2888 2369
rect 2908 2349 2917 2369
rect 2873 2343 2917 2349
rect 2987 2369 3031 2385
rect 2987 2349 2996 2369
rect 3016 2349 3031 2369
rect 2987 2343 3031 2349
rect 3081 2373 3130 2385
rect 3081 2353 3099 2373
rect 3119 2353 3130 2373
rect 3081 2343 3130 2353
rect 3195 2369 3239 2385
rect 3195 2349 3204 2369
rect 3224 2349 3239 2369
rect 3195 2343 3239 2349
rect 3289 2373 3338 2385
rect 3289 2353 3307 2373
rect 3327 2353 3338 2373
rect 3289 2343 3338 2353
rect 3408 2369 3452 2385
rect 3408 2349 3417 2369
rect 3437 2349 3452 2369
rect 3408 2343 3452 2349
rect 3502 2373 3551 2385
rect 3502 2353 3520 2373
rect 3540 2353 3551 2373
rect 3502 2343 3551 2353
rect 1384 2146 1433 2156
rect 1384 2126 1395 2146
rect 1415 2126 1433 2146
rect 1384 2114 1433 2126
rect 1483 2150 1527 2156
rect 1483 2130 1498 2150
rect 1518 2130 1527 2150
rect 1483 2114 1527 2130
rect 1597 2146 1646 2156
rect 1597 2126 1608 2146
rect 1628 2126 1646 2146
rect 1597 2114 1646 2126
rect 1696 2150 1740 2156
rect 1696 2130 1711 2150
rect 1731 2130 1740 2150
rect 1696 2114 1740 2130
rect 1805 2146 1854 2156
rect 1805 2126 1816 2146
rect 1836 2126 1854 2146
rect 1805 2114 1854 2126
rect 1904 2150 1948 2156
rect 1904 2130 1919 2150
rect 1939 2130 1948 2150
rect 1904 2114 1948 2130
rect 2018 2150 2062 2156
rect 2018 2130 2027 2150
rect 2047 2130 2062 2150
rect 2018 2114 2062 2130
rect 2112 2146 2161 2156
rect 2112 2126 2130 2146
rect 2150 2126 2161 2146
rect 2112 2114 2161 2126
rect 3823 2104 3872 2116
rect 3823 2084 3834 2104
rect 3854 2084 3872 2104
rect 3823 2074 3872 2084
rect 3922 2100 3966 2116
rect 3922 2080 3937 2100
rect 3957 2080 3966 2100
rect 3922 2074 3966 2080
rect 4036 2100 4080 2116
rect 4036 2080 4045 2100
rect 4065 2080 4080 2100
rect 4036 2074 4080 2080
rect 4130 2104 4179 2116
rect 4130 2084 4148 2104
rect 4168 2084 4179 2104
rect 4130 2074 4179 2084
rect 4244 2100 4288 2116
rect 4244 2080 4253 2100
rect 4273 2080 4288 2100
rect 4244 2074 4288 2080
rect 4338 2104 4387 2116
rect 4338 2084 4356 2104
rect 4376 2084 4387 2104
rect 4338 2074 4387 2084
rect 4457 2100 4501 2116
rect 4457 2080 4466 2100
rect 4486 2080 4501 2100
rect 4457 2074 4501 2080
rect 4551 2104 4600 2116
rect 4551 2084 4569 2104
rect 4589 2084 4600 2104
rect 4551 2074 4600 2084
rect 336 1866 385 1876
rect 336 1846 347 1866
rect 367 1846 385 1866
rect 336 1834 385 1846
rect 435 1870 479 1876
rect 435 1850 450 1870
rect 470 1850 479 1870
rect 435 1834 479 1850
rect 549 1866 598 1876
rect 549 1846 560 1866
rect 580 1846 598 1866
rect 549 1834 598 1846
rect 648 1870 692 1876
rect 648 1850 663 1870
rect 683 1850 692 1870
rect 648 1834 692 1850
rect 757 1866 806 1876
rect 757 1846 768 1866
rect 788 1846 806 1866
rect 757 1834 806 1846
rect 856 1870 900 1876
rect 856 1850 871 1870
rect 891 1850 900 1870
rect 856 1834 900 1850
rect 970 1870 1014 1876
rect 970 1850 979 1870
rect 999 1850 1014 1870
rect 970 1834 1014 1850
rect 1064 1866 1113 1876
rect 1064 1846 1082 1866
rect 1102 1846 1113 1866
rect 1064 1834 1113 1846
rect 2884 1794 2933 1806
rect 2884 1774 2895 1794
rect 2915 1774 2933 1794
rect 2884 1764 2933 1774
rect 2983 1790 3027 1806
rect 2983 1770 2998 1790
rect 3018 1770 3027 1790
rect 2983 1764 3027 1770
rect 3097 1790 3141 1806
rect 3097 1770 3106 1790
rect 3126 1770 3141 1790
rect 3097 1764 3141 1770
rect 3191 1794 3240 1806
rect 3191 1774 3209 1794
rect 3229 1774 3240 1794
rect 3191 1764 3240 1774
rect 3305 1790 3349 1806
rect 3305 1770 3314 1790
rect 3334 1770 3349 1790
rect 3305 1764 3349 1770
rect 3399 1794 3448 1806
rect 3399 1774 3417 1794
rect 3437 1774 3448 1794
rect 3399 1764 3448 1774
rect 3518 1790 3562 1806
rect 3518 1770 3527 1790
rect 3547 1770 3562 1790
rect 3518 1764 3562 1770
rect 3612 1794 3661 1806
rect 3612 1774 3630 1794
rect 3650 1774 3661 1794
rect 3612 1764 3661 1774
rect 1274 1622 1323 1632
rect 1274 1602 1285 1622
rect 1305 1602 1323 1622
rect 1274 1590 1323 1602
rect 1373 1626 1417 1632
rect 1373 1606 1388 1626
rect 1408 1606 1417 1626
rect 1373 1590 1417 1606
rect 1487 1622 1536 1632
rect 1487 1602 1498 1622
rect 1518 1602 1536 1622
rect 1487 1590 1536 1602
rect 1586 1626 1630 1632
rect 1586 1606 1601 1626
rect 1621 1606 1630 1626
rect 1586 1590 1630 1606
rect 1695 1622 1744 1632
rect 1695 1602 1706 1622
rect 1726 1602 1744 1622
rect 1695 1590 1744 1602
rect 1794 1626 1838 1632
rect 1794 1606 1809 1626
rect 1829 1606 1838 1626
rect 1794 1590 1838 1606
rect 1908 1626 1952 1632
rect 1908 1606 1917 1626
rect 1937 1606 1952 1626
rect 1908 1590 1952 1606
rect 2002 1622 2051 1632
rect 2002 1602 2020 1622
rect 2040 1602 2051 1622
rect 2002 1590 2051 1602
rect 3822 1550 3871 1562
rect 3822 1530 3833 1550
rect 3853 1530 3871 1550
rect 3822 1520 3871 1530
rect 3921 1546 3965 1562
rect 3921 1526 3936 1546
rect 3956 1526 3965 1546
rect 3921 1520 3965 1526
rect 4035 1546 4079 1562
rect 4035 1526 4044 1546
rect 4064 1526 4079 1546
rect 4035 1520 4079 1526
rect 4129 1550 4178 1562
rect 4129 1530 4147 1550
rect 4167 1530 4178 1550
rect 4129 1520 4178 1530
rect 4243 1546 4287 1562
rect 4243 1526 4252 1546
rect 4272 1526 4287 1546
rect 4243 1520 4287 1526
rect 4337 1550 4386 1562
rect 4337 1530 4355 1550
rect 4375 1530 4386 1550
rect 4337 1520 4386 1530
rect 4456 1546 4500 1562
rect 4456 1526 4465 1546
rect 4485 1526 4500 1546
rect 4456 1520 4500 1526
rect 4550 1550 4599 1562
rect 4550 1530 4568 1550
rect 4588 1530 4599 1550
rect 4550 1520 4599 1530
rect 335 1312 384 1322
rect 335 1292 346 1312
rect 366 1292 384 1312
rect 335 1280 384 1292
rect 434 1316 478 1322
rect 434 1296 449 1316
rect 469 1296 478 1316
rect 434 1280 478 1296
rect 548 1312 597 1322
rect 548 1292 559 1312
rect 579 1292 597 1312
rect 548 1280 597 1292
rect 647 1316 691 1322
rect 647 1296 662 1316
rect 682 1296 691 1316
rect 647 1280 691 1296
rect 756 1312 805 1322
rect 756 1292 767 1312
rect 787 1292 805 1312
rect 756 1280 805 1292
rect 855 1316 899 1322
rect 855 1296 870 1316
rect 890 1296 899 1316
rect 855 1280 899 1296
rect 969 1316 1013 1322
rect 969 1296 978 1316
rect 998 1296 1013 1316
rect 969 1280 1013 1296
rect 1063 1312 1112 1322
rect 1063 1292 1081 1312
rect 1101 1292 1112 1312
rect 1063 1280 1112 1292
rect 2744 1283 2793 1295
rect 2744 1263 2755 1283
rect 2775 1263 2793 1283
rect 2744 1253 2793 1263
rect 2843 1279 2887 1295
rect 2843 1259 2858 1279
rect 2878 1259 2887 1279
rect 2843 1253 2887 1259
rect 2957 1279 3001 1295
rect 2957 1259 2966 1279
rect 2986 1259 3001 1279
rect 2957 1253 3001 1259
rect 3051 1283 3100 1295
rect 3051 1263 3069 1283
rect 3089 1263 3100 1283
rect 3051 1253 3100 1263
rect 3165 1279 3209 1295
rect 3165 1259 3174 1279
rect 3194 1259 3209 1279
rect 3165 1253 3209 1259
rect 3259 1283 3308 1295
rect 3259 1263 3277 1283
rect 3297 1263 3308 1283
rect 3259 1253 3308 1263
rect 3378 1279 3422 1295
rect 3378 1259 3387 1279
rect 3407 1259 3422 1279
rect 3378 1253 3422 1259
rect 3472 1283 3521 1295
rect 3472 1263 3490 1283
rect 3510 1263 3521 1283
rect 3472 1253 3521 1263
rect 1415 1030 1464 1040
rect 1415 1010 1426 1030
rect 1446 1010 1464 1030
rect 1415 998 1464 1010
rect 1514 1034 1558 1040
rect 1514 1014 1529 1034
rect 1549 1014 1558 1034
rect 1514 998 1558 1014
rect 1628 1030 1677 1040
rect 1628 1010 1639 1030
rect 1659 1010 1677 1030
rect 1628 998 1677 1010
rect 1727 1034 1771 1040
rect 1727 1014 1742 1034
rect 1762 1014 1771 1034
rect 1727 998 1771 1014
rect 1836 1030 1885 1040
rect 1836 1010 1847 1030
rect 1867 1010 1885 1030
rect 1836 998 1885 1010
rect 1935 1034 1979 1040
rect 1935 1014 1950 1034
rect 1970 1014 1979 1034
rect 1935 998 1979 1014
rect 2049 1034 2093 1040
rect 2049 1014 2058 1034
rect 2078 1014 2093 1034
rect 2049 998 2093 1014
rect 2143 1030 2192 1040
rect 2143 1010 2161 1030
rect 2181 1010 2192 1030
rect 2143 998 2192 1010
rect 3824 1001 3873 1013
rect 3824 981 3835 1001
rect 3855 981 3873 1001
rect 3824 971 3873 981
rect 3923 997 3967 1013
rect 3923 977 3938 997
rect 3958 977 3967 997
rect 3923 971 3967 977
rect 4037 997 4081 1013
rect 4037 977 4046 997
rect 4066 977 4081 997
rect 4037 971 4081 977
rect 4131 1001 4180 1013
rect 4131 981 4149 1001
rect 4169 981 4180 1001
rect 4131 971 4180 981
rect 4245 997 4289 1013
rect 4245 977 4254 997
rect 4274 977 4289 997
rect 4245 971 4289 977
rect 4339 1001 4388 1013
rect 4339 981 4357 1001
rect 4377 981 4388 1001
rect 4339 971 4388 981
rect 4458 997 4502 1013
rect 4458 977 4467 997
rect 4487 977 4502 997
rect 4458 971 4502 977
rect 4552 1001 4601 1013
rect 4552 981 4570 1001
rect 4590 981 4601 1001
rect 4552 971 4601 981
rect 337 763 386 773
rect 337 743 348 763
rect 368 743 386 763
rect 337 731 386 743
rect 436 767 480 773
rect 436 747 451 767
rect 471 747 480 767
rect 436 731 480 747
rect 550 763 599 773
rect 550 743 561 763
rect 581 743 599 763
rect 550 731 599 743
rect 649 767 693 773
rect 649 747 664 767
rect 684 747 693 767
rect 649 731 693 747
rect 758 763 807 773
rect 758 743 769 763
rect 789 743 807 763
rect 758 731 807 743
rect 857 767 901 773
rect 857 747 872 767
rect 892 747 901 767
rect 857 731 901 747
rect 971 767 1015 773
rect 971 747 980 767
rect 1000 747 1015 767
rect 971 731 1015 747
rect 1065 763 1114 773
rect 1065 743 1083 763
rect 1103 743 1114 763
rect 1065 731 1114 743
rect 2885 691 2934 703
rect 2885 671 2896 691
rect 2916 671 2934 691
rect 2885 661 2934 671
rect 2984 687 3028 703
rect 2984 667 2999 687
rect 3019 667 3028 687
rect 2984 661 3028 667
rect 3098 687 3142 703
rect 3098 667 3107 687
rect 3127 667 3142 687
rect 3098 661 3142 667
rect 3192 691 3241 703
rect 3192 671 3210 691
rect 3230 671 3241 691
rect 3192 661 3241 671
rect 3306 687 3350 703
rect 3306 667 3315 687
rect 3335 667 3350 687
rect 3306 661 3350 667
rect 3400 691 3449 703
rect 3400 671 3418 691
rect 3438 671 3449 691
rect 3400 661 3449 671
rect 3519 687 3563 703
rect 3519 667 3528 687
rect 3548 667 3563 687
rect 3519 661 3563 667
rect 3613 691 3662 703
rect 3613 671 3631 691
rect 3651 671 3662 691
rect 3613 661 3662 671
rect 1275 519 1324 529
rect 1275 499 1286 519
rect 1306 499 1324 519
rect 1275 487 1324 499
rect 1374 523 1418 529
rect 1374 503 1389 523
rect 1409 503 1418 523
rect 1374 487 1418 503
rect 1488 519 1537 529
rect 1488 499 1499 519
rect 1519 499 1537 519
rect 1488 487 1537 499
rect 1587 523 1631 529
rect 1587 503 1602 523
rect 1622 503 1631 523
rect 1587 487 1631 503
rect 1696 519 1745 529
rect 1696 499 1707 519
rect 1727 499 1745 519
rect 1696 487 1745 499
rect 1795 523 1839 529
rect 1795 503 1810 523
rect 1830 503 1839 523
rect 1795 487 1839 503
rect 1909 523 1953 529
rect 1909 503 1918 523
rect 1938 503 1953 523
rect 1909 487 1953 503
rect 2003 519 2052 529
rect 2003 499 2021 519
rect 2041 499 2052 519
rect 2003 487 2052 499
rect 3823 447 3872 459
rect 3823 427 3834 447
rect 3854 427 3872 447
rect 3823 417 3872 427
rect 3922 443 3966 459
rect 3922 423 3937 443
rect 3957 423 3966 443
rect 3922 417 3966 423
rect 4036 443 4080 459
rect 4036 423 4045 443
rect 4065 423 4080 443
rect 4036 417 4080 423
rect 4130 447 4179 459
rect 4130 427 4148 447
rect 4168 427 4179 447
rect 4130 417 4179 427
rect 4244 443 4288 459
rect 4244 423 4253 443
rect 4273 423 4288 443
rect 4244 417 4288 423
rect 4338 447 4387 459
rect 4338 427 4356 447
rect 4376 427 4387 447
rect 4338 417 4387 427
rect 4457 443 4501 459
rect 4457 423 4466 443
rect 4486 423 4501 443
rect 4457 417 4501 423
rect 4551 447 4600 459
rect 4551 427 4569 447
rect 4589 427 4600 447
rect 4551 417 4600 427
rect 336 209 385 219
rect 336 189 347 209
rect 367 189 385 209
rect 336 177 385 189
rect 435 213 479 219
rect 435 193 450 213
rect 470 193 479 213
rect 435 177 479 193
rect 549 209 598 219
rect 549 189 560 209
rect 580 189 598 209
rect 549 177 598 189
rect 648 213 692 219
rect 648 193 663 213
rect 683 193 692 213
rect 648 177 692 193
rect 757 209 806 219
rect 757 189 768 209
rect 788 189 806 209
rect 757 177 806 189
rect 856 213 900 219
rect 856 193 871 213
rect 891 193 900 213
rect 856 177 900 193
rect 970 213 1014 219
rect 970 193 979 213
rect 999 193 1014 213
rect 970 177 1014 193
rect 1064 209 1113 219
rect 1064 189 1082 209
rect 1102 189 1113 209
rect 1064 177 1113 189
rect 1583 -350 1632 -340
rect 1583 -370 1594 -350
rect 1614 -370 1632 -350
rect 1583 -382 1632 -370
rect 1682 -346 1726 -340
rect 1682 -366 1697 -346
rect 1717 -366 1726 -346
rect 1682 -382 1726 -366
rect 1796 -350 1845 -340
rect 1796 -370 1807 -350
rect 1827 -370 1845 -350
rect 1796 -382 1845 -370
rect 1895 -346 1939 -340
rect 1895 -366 1910 -346
rect 1930 -366 1939 -346
rect 1895 -382 1939 -366
rect 2004 -350 2053 -340
rect 2004 -370 2015 -350
rect 2035 -370 2053 -350
rect 2004 -382 2053 -370
rect 2103 -346 2147 -340
rect 2103 -366 2118 -346
rect 2138 -366 2147 -346
rect 2103 -382 2147 -366
rect 2217 -346 2261 -340
rect 2217 -366 2226 -346
rect 2246 -366 2261 -346
rect 2217 -382 2261 -366
rect 2311 -350 2360 -340
rect 2311 -370 2329 -350
rect 2349 -370 2360 -350
rect 2311 -382 2360 -370
<< pdiff >>
rect 338 8633 382 8671
rect 338 8613 350 8633
rect 370 8613 382 8633
rect 338 8571 382 8613
rect 432 8633 474 8671
rect 432 8613 446 8633
rect 466 8613 474 8633
rect 432 8571 474 8613
rect 551 8633 595 8671
rect 551 8613 563 8633
rect 583 8613 595 8633
rect 551 8571 595 8613
rect 645 8633 687 8671
rect 645 8613 659 8633
rect 679 8613 687 8633
rect 645 8571 687 8613
rect 759 8633 803 8671
rect 759 8613 771 8633
rect 791 8613 803 8633
rect 759 8571 803 8613
rect 853 8633 895 8671
rect 853 8613 867 8633
rect 887 8613 895 8633
rect 853 8571 895 8613
rect 969 8633 1011 8671
rect 969 8613 977 8633
rect 997 8613 1011 8633
rect 969 8571 1011 8613
rect 1061 8640 1106 8671
rect 1061 8633 1105 8640
rect 1061 8613 1073 8633
rect 1093 8613 1105 8633
rect 1061 8571 1105 8613
rect 3825 8573 3869 8615
rect 3825 8553 3837 8573
rect 3857 8553 3869 8573
rect 3825 8546 3869 8553
rect 3824 8515 3869 8546
rect 3919 8573 3961 8615
rect 3919 8553 3933 8573
rect 3953 8553 3961 8573
rect 3919 8515 3961 8553
rect 4035 8573 4077 8615
rect 4035 8553 4043 8573
rect 4063 8553 4077 8573
rect 4035 8515 4077 8553
rect 4127 8573 4171 8615
rect 4127 8553 4139 8573
rect 4159 8553 4171 8573
rect 4127 8515 4171 8553
rect 4243 8573 4285 8615
rect 4243 8553 4251 8573
rect 4271 8553 4285 8573
rect 4243 8515 4285 8553
rect 4335 8573 4379 8615
rect 4335 8553 4347 8573
rect 4367 8553 4379 8573
rect 4335 8515 4379 8553
rect 4456 8573 4498 8615
rect 4456 8553 4464 8573
rect 4484 8553 4498 8573
rect 4456 8515 4498 8553
rect 4548 8573 4592 8615
rect 4548 8553 4560 8573
rect 4580 8553 4592 8573
rect 4548 8515 4592 8553
rect 1276 8389 1320 8427
rect 1276 8369 1288 8389
rect 1308 8369 1320 8389
rect 1276 8327 1320 8369
rect 1370 8389 1412 8427
rect 1370 8369 1384 8389
rect 1404 8369 1412 8389
rect 1370 8327 1412 8369
rect 1489 8389 1533 8427
rect 1489 8369 1501 8389
rect 1521 8369 1533 8389
rect 1489 8327 1533 8369
rect 1583 8389 1625 8427
rect 1583 8369 1597 8389
rect 1617 8369 1625 8389
rect 1583 8327 1625 8369
rect 1697 8389 1741 8427
rect 1697 8369 1709 8389
rect 1729 8369 1741 8389
rect 1697 8327 1741 8369
rect 1791 8389 1833 8427
rect 1791 8369 1805 8389
rect 1825 8369 1833 8389
rect 1791 8327 1833 8369
rect 1907 8389 1949 8427
rect 1907 8369 1915 8389
rect 1935 8369 1949 8389
rect 1907 8327 1949 8369
rect 1999 8396 2044 8427
rect 1999 8389 2043 8396
rect 1999 8369 2011 8389
rect 2031 8369 2043 8389
rect 1999 8327 2043 8369
rect 2886 8263 2930 8305
rect 2886 8243 2898 8263
rect 2918 8243 2930 8263
rect 2886 8236 2930 8243
rect 2885 8205 2930 8236
rect 2980 8263 3022 8305
rect 2980 8243 2994 8263
rect 3014 8243 3022 8263
rect 2980 8205 3022 8243
rect 3096 8263 3138 8305
rect 3096 8243 3104 8263
rect 3124 8243 3138 8263
rect 3096 8205 3138 8243
rect 3188 8263 3232 8305
rect 3188 8243 3200 8263
rect 3220 8243 3232 8263
rect 3188 8205 3232 8243
rect 3304 8263 3346 8305
rect 3304 8243 3312 8263
rect 3332 8243 3346 8263
rect 3304 8205 3346 8243
rect 3396 8263 3440 8305
rect 3396 8243 3408 8263
rect 3428 8243 3440 8263
rect 3396 8205 3440 8243
rect 3517 8263 3559 8305
rect 3517 8243 3525 8263
rect 3545 8243 3559 8263
rect 3517 8205 3559 8243
rect 3609 8263 3653 8305
rect 3609 8243 3621 8263
rect 3641 8243 3653 8263
rect 3609 8205 3653 8243
rect 337 8079 381 8117
rect 337 8059 349 8079
rect 369 8059 381 8079
rect 337 8017 381 8059
rect 431 8079 473 8117
rect 431 8059 445 8079
rect 465 8059 473 8079
rect 431 8017 473 8059
rect 550 8079 594 8117
rect 550 8059 562 8079
rect 582 8059 594 8079
rect 550 8017 594 8059
rect 644 8079 686 8117
rect 644 8059 658 8079
rect 678 8059 686 8079
rect 644 8017 686 8059
rect 758 8079 802 8117
rect 758 8059 770 8079
rect 790 8059 802 8079
rect 758 8017 802 8059
rect 852 8079 894 8117
rect 852 8059 866 8079
rect 886 8059 894 8079
rect 852 8017 894 8059
rect 968 8079 1010 8117
rect 968 8059 976 8079
rect 996 8059 1010 8079
rect 968 8017 1010 8059
rect 1060 8086 1105 8117
rect 1060 8079 1104 8086
rect 1060 8059 1072 8079
rect 1092 8059 1104 8079
rect 1060 8017 1104 8059
rect 3824 8019 3868 8061
rect 3824 7999 3836 8019
rect 3856 7999 3868 8019
rect 3824 7992 3868 7999
rect 3823 7961 3868 7992
rect 3918 8019 3960 8061
rect 3918 7999 3932 8019
rect 3952 7999 3960 8019
rect 3918 7961 3960 7999
rect 4034 8019 4076 8061
rect 4034 7999 4042 8019
rect 4062 7999 4076 8019
rect 4034 7961 4076 7999
rect 4126 8019 4170 8061
rect 4126 7999 4138 8019
rect 4158 7999 4170 8019
rect 4126 7961 4170 7999
rect 4242 8019 4284 8061
rect 4242 7999 4250 8019
rect 4270 7999 4284 8019
rect 4242 7961 4284 7999
rect 4334 8019 4378 8061
rect 4334 7999 4346 8019
rect 4366 7999 4378 8019
rect 4334 7961 4378 7999
rect 4455 8019 4497 8061
rect 4455 7999 4463 8019
rect 4483 7999 4497 8019
rect 4455 7961 4497 7999
rect 4547 8019 4591 8061
rect 4547 7999 4559 8019
rect 4579 7999 4591 8019
rect 4547 7961 4591 7999
rect 1417 7797 1461 7835
rect 1417 7777 1429 7797
rect 1449 7777 1461 7797
rect 1417 7735 1461 7777
rect 1511 7797 1553 7835
rect 1511 7777 1525 7797
rect 1545 7777 1553 7797
rect 1511 7735 1553 7777
rect 1630 7797 1674 7835
rect 1630 7777 1642 7797
rect 1662 7777 1674 7797
rect 1630 7735 1674 7777
rect 1724 7797 1766 7835
rect 1724 7777 1738 7797
rect 1758 7777 1766 7797
rect 1724 7735 1766 7777
rect 1838 7797 1882 7835
rect 1838 7777 1850 7797
rect 1870 7777 1882 7797
rect 1838 7735 1882 7777
rect 1932 7797 1974 7835
rect 1932 7777 1946 7797
rect 1966 7777 1974 7797
rect 1932 7735 1974 7777
rect 2048 7797 2090 7835
rect 2048 7777 2056 7797
rect 2076 7777 2090 7797
rect 2048 7735 2090 7777
rect 2140 7804 2185 7835
rect 2140 7797 2184 7804
rect 2140 7777 2152 7797
rect 2172 7777 2184 7797
rect 2140 7735 2184 7777
rect 2746 7752 2790 7794
rect 2746 7732 2758 7752
rect 2778 7732 2790 7752
rect 2746 7725 2790 7732
rect 2745 7694 2790 7725
rect 2840 7752 2882 7794
rect 2840 7732 2854 7752
rect 2874 7732 2882 7752
rect 2840 7694 2882 7732
rect 2956 7752 2998 7794
rect 2956 7732 2964 7752
rect 2984 7732 2998 7752
rect 2956 7694 2998 7732
rect 3048 7752 3092 7794
rect 3048 7732 3060 7752
rect 3080 7732 3092 7752
rect 3048 7694 3092 7732
rect 3164 7752 3206 7794
rect 3164 7732 3172 7752
rect 3192 7732 3206 7752
rect 3164 7694 3206 7732
rect 3256 7752 3300 7794
rect 3256 7732 3268 7752
rect 3288 7732 3300 7752
rect 3256 7694 3300 7732
rect 3377 7752 3419 7794
rect 3377 7732 3385 7752
rect 3405 7732 3419 7752
rect 3377 7694 3419 7732
rect 3469 7752 3513 7794
rect 3469 7732 3481 7752
rect 3501 7732 3513 7752
rect 3469 7694 3513 7732
rect 339 7530 383 7568
rect 339 7510 351 7530
rect 371 7510 383 7530
rect 339 7468 383 7510
rect 433 7530 475 7568
rect 433 7510 447 7530
rect 467 7510 475 7530
rect 433 7468 475 7510
rect 552 7530 596 7568
rect 552 7510 564 7530
rect 584 7510 596 7530
rect 552 7468 596 7510
rect 646 7530 688 7568
rect 646 7510 660 7530
rect 680 7510 688 7530
rect 646 7468 688 7510
rect 760 7530 804 7568
rect 760 7510 772 7530
rect 792 7510 804 7530
rect 760 7468 804 7510
rect 854 7530 896 7568
rect 854 7510 868 7530
rect 888 7510 896 7530
rect 854 7468 896 7510
rect 970 7530 1012 7568
rect 970 7510 978 7530
rect 998 7510 1012 7530
rect 970 7468 1012 7510
rect 1062 7537 1107 7568
rect 1062 7530 1106 7537
rect 1062 7510 1074 7530
rect 1094 7510 1106 7530
rect 1062 7468 1106 7510
rect 3826 7470 3870 7512
rect 3826 7450 3838 7470
rect 3858 7450 3870 7470
rect 3826 7443 3870 7450
rect 3825 7412 3870 7443
rect 3920 7470 3962 7512
rect 3920 7450 3934 7470
rect 3954 7450 3962 7470
rect 3920 7412 3962 7450
rect 4036 7470 4078 7512
rect 4036 7450 4044 7470
rect 4064 7450 4078 7470
rect 4036 7412 4078 7450
rect 4128 7470 4172 7512
rect 4128 7450 4140 7470
rect 4160 7450 4172 7470
rect 4128 7412 4172 7450
rect 4244 7470 4286 7512
rect 4244 7450 4252 7470
rect 4272 7450 4286 7470
rect 4244 7412 4286 7450
rect 4336 7470 4380 7512
rect 4336 7450 4348 7470
rect 4368 7450 4380 7470
rect 4336 7412 4380 7450
rect 4457 7470 4499 7512
rect 4457 7450 4465 7470
rect 4485 7450 4499 7470
rect 4457 7412 4499 7450
rect 4549 7470 4593 7512
rect 4549 7450 4561 7470
rect 4581 7450 4593 7470
rect 4549 7412 4593 7450
rect 1277 7286 1321 7324
rect 1277 7266 1289 7286
rect 1309 7266 1321 7286
rect 1277 7224 1321 7266
rect 1371 7286 1413 7324
rect 1371 7266 1385 7286
rect 1405 7266 1413 7286
rect 1371 7224 1413 7266
rect 1490 7286 1534 7324
rect 1490 7266 1502 7286
rect 1522 7266 1534 7286
rect 1490 7224 1534 7266
rect 1584 7286 1626 7324
rect 1584 7266 1598 7286
rect 1618 7266 1626 7286
rect 1584 7224 1626 7266
rect 1698 7286 1742 7324
rect 1698 7266 1710 7286
rect 1730 7266 1742 7286
rect 1698 7224 1742 7266
rect 1792 7286 1834 7324
rect 1792 7266 1806 7286
rect 1826 7266 1834 7286
rect 1792 7224 1834 7266
rect 1908 7286 1950 7324
rect 1908 7266 1916 7286
rect 1936 7266 1950 7286
rect 1908 7224 1950 7266
rect 2000 7293 2045 7324
rect 2000 7286 2044 7293
rect 2000 7266 2012 7286
rect 2032 7266 2044 7286
rect 2000 7224 2044 7266
rect 2887 7160 2931 7202
rect 2887 7140 2899 7160
rect 2919 7140 2931 7160
rect 2887 7133 2931 7140
rect 2886 7102 2931 7133
rect 2981 7160 3023 7202
rect 2981 7140 2995 7160
rect 3015 7140 3023 7160
rect 2981 7102 3023 7140
rect 3097 7160 3139 7202
rect 3097 7140 3105 7160
rect 3125 7140 3139 7160
rect 3097 7102 3139 7140
rect 3189 7160 3233 7202
rect 3189 7140 3201 7160
rect 3221 7140 3233 7160
rect 3189 7102 3233 7140
rect 3305 7160 3347 7202
rect 3305 7140 3313 7160
rect 3333 7140 3347 7160
rect 3305 7102 3347 7140
rect 3397 7160 3441 7202
rect 3397 7140 3409 7160
rect 3429 7140 3441 7160
rect 3397 7102 3441 7140
rect 3518 7160 3560 7202
rect 3518 7140 3526 7160
rect 3546 7140 3560 7160
rect 3518 7102 3560 7140
rect 3610 7160 3654 7202
rect 3610 7140 3622 7160
rect 3642 7140 3654 7160
rect 3610 7102 3654 7140
rect 338 6976 382 7014
rect 338 6956 350 6976
rect 370 6956 382 6976
rect 338 6914 382 6956
rect 432 6976 474 7014
rect 432 6956 446 6976
rect 466 6956 474 6976
rect 432 6914 474 6956
rect 551 6976 595 7014
rect 551 6956 563 6976
rect 583 6956 595 6976
rect 551 6914 595 6956
rect 645 6976 687 7014
rect 645 6956 659 6976
rect 679 6956 687 6976
rect 645 6914 687 6956
rect 759 6976 803 7014
rect 759 6956 771 6976
rect 791 6956 803 6976
rect 759 6914 803 6956
rect 853 6976 895 7014
rect 853 6956 867 6976
rect 887 6956 895 6976
rect 853 6914 895 6956
rect 969 6976 1011 7014
rect 969 6956 977 6976
rect 997 6956 1011 6976
rect 969 6914 1011 6956
rect 1061 6983 1106 7014
rect 1061 6976 1105 6983
rect 1061 6956 1073 6976
rect 1093 6956 1105 6976
rect 1061 6914 1105 6956
rect 3825 6916 3869 6958
rect 3825 6896 3837 6916
rect 3857 6896 3869 6916
rect 3825 6889 3869 6896
rect 3824 6858 3869 6889
rect 3919 6916 3961 6958
rect 3919 6896 3933 6916
rect 3953 6896 3961 6916
rect 3919 6858 3961 6896
rect 4035 6916 4077 6958
rect 4035 6896 4043 6916
rect 4063 6896 4077 6916
rect 4035 6858 4077 6896
rect 4127 6916 4171 6958
rect 4127 6896 4139 6916
rect 4159 6896 4171 6916
rect 4127 6858 4171 6896
rect 4243 6916 4285 6958
rect 4243 6896 4251 6916
rect 4271 6896 4285 6916
rect 4243 6858 4285 6896
rect 4335 6916 4379 6958
rect 4335 6896 4347 6916
rect 4367 6896 4379 6916
rect 4335 6858 4379 6896
rect 4456 6916 4498 6958
rect 4456 6896 4464 6916
rect 4484 6896 4498 6916
rect 4456 6858 4498 6896
rect 4548 6916 4592 6958
rect 4548 6896 4560 6916
rect 4580 6896 4592 6916
rect 4548 6858 4592 6896
rect 1387 6707 1431 6745
rect 1387 6687 1399 6707
rect 1419 6687 1431 6707
rect 1387 6645 1431 6687
rect 1481 6707 1523 6745
rect 1481 6687 1495 6707
rect 1515 6687 1523 6707
rect 1481 6645 1523 6687
rect 1600 6707 1644 6745
rect 1600 6687 1612 6707
rect 1632 6687 1644 6707
rect 1600 6645 1644 6687
rect 1694 6707 1736 6745
rect 1694 6687 1708 6707
rect 1728 6687 1736 6707
rect 1694 6645 1736 6687
rect 1808 6707 1852 6745
rect 1808 6687 1820 6707
rect 1840 6687 1852 6707
rect 1808 6645 1852 6687
rect 1902 6707 1944 6745
rect 1902 6687 1916 6707
rect 1936 6687 1944 6707
rect 1902 6645 1944 6687
rect 2018 6707 2060 6745
rect 2018 6687 2026 6707
rect 2046 6687 2060 6707
rect 2018 6645 2060 6687
rect 2110 6714 2155 6745
rect 2110 6707 2154 6714
rect 2110 6687 2122 6707
rect 2142 6687 2154 6707
rect 2110 6645 2154 6687
rect 2777 6636 2821 6678
rect 2777 6616 2789 6636
rect 2809 6616 2821 6636
rect 2777 6609 2821 6616
rect 2776 6578 2821 6609
rect 2871 6636 2913 6678
rect 2871 6616 2885 6636
rect 2905 6616 2913 6636
rect 2871 6578 2913 6616
rect 2987 6636 3029 6678
rect 2987 6616 2995 6636
rect 3015 6616 3029 6636
rect 2987 6578 3029 6616
rect 3079 6636 3123 6678
rect 3079 6616 3091 6636
rect 3111 6616 3123 6636
rect 3079 6578 3123 6616
rect 3195 6636 3237 6678
rect 3195 6616 3203 6636
rect 3223 6616 3237 6636
rect 3195 6578 3237 6616
rect 3287 6636 3331 6678
rect 3287 6616 3299 6636
rect 3319 6616 3331 6636
rect 3287 6578 3331 6616
rect 3408 6636 3450 6678
rect 3408 6616 3416 6636
rect 3436 6616 3450 6636
rect 3408 6578 3450 6616
rect 3500 6636 3544 6678
rect 3500 6616 3512 6636
rect 3532 6616 3544 6636
rect 3500 6578 3544 6616
rect 339 6427 383 6465
rect 339 6407 351 6427
rect 371 6407 383 6427
rect 339 6365 383 6407
rect 433 6427 475 6465
rect 433 6407 447 6427
rect 467 6407 475 6427
rect 433 6365 475 6407
rect 552 6427 596 6465
rect 552 6407 564 6427
rect 584 6407 596 6427
rect 552 6365 596 6407
rect 646 6427 688 6465
rect 646 6407 660 6427
rect 680 6407 688 6427
rect 646 6365 688 6407
rect 760 6427 804 6465
rect 760 6407 772 6427
rect 792 6407 804 6427
rect 760 6365 804 6407
rect 854 6427 896 6465
rect 854 6407 868 6427
rect 888 6407 896 6427
rect 854 6365 896 6407
rect 970 6427 1012 6465
rect 970 6407 978 6427
rect 998 6407 1012 6427
rect 970 6365 1012 6407
rect 1062 6434 1107 6465
rect 1062 6427 1106 6434
rect 1062 6407 1074 6427
rect 1094 6407 1106 6427
rect 1062 6365 1106 6407
rect 3826 6367 3870 6409
rect 3826 6347 3838 6367
rect 3858 6347 3870 6367
rect 3826 6340 3870 6347
rect 3825 6309 3870 6340
rect 3920 6367 3962 6409
rect 3920 6347 3934 6367
rect 3954 6347 3962 6367
rect 3920 6309 3962 6347
rect 4036 6367 4078 6409
rect 4036 6347 4044 6367
rect 4064 6347 4078 6367
rect 4036 6309 4078 6347
rect 4128 6367 4172 6409
rect 4128 6347 4140 6367
rect 4160 6347 4172 6367
rect 4128 6309 4172 6347
rect 4244 6367 4286 6409
rect 4244 6347 4252 6367
rect 4272 6347 4286 6367
rect 4244 6309 4286 6347
rect 4336 6367 4380 6409
rect 4336 6347 4348 6367
rect 4368 6347 4380 6367
rect 4336 6309 4380 6347
rect 4457 6367 4499 6409
rect 4457 6347 4465 6367
rect 4485 6347 4499 6367
rect 4457 6309 4499 6347
rect 4549 6367 4593 6409
rect 4549 6347 4561 6367
rect 4581 6347 4593 6367
rect 4549 6309 4593 6347
rect 1277 6183 1321 6221
rect 1277 6163 1289 6183
rect 1309 6163 1321 6183
rect 1277 6121 1321 6163
rect 1371 6183 1413 6221
rect 1371 6163 1385 6183
rect 1405 6163 1413 6183
rect 1371 6121 1413 6163
rect 1490 6183 1534 6221
rect 1490 6163 1502 6183
rect 1522 6163 1534 6183
rect 1490 6121 1534 6163
rect 1584 6183 1626 6221
rect 1584 6163 1598 6183
rect 1618 6163 1626 6183
rect 1584 6121 1626 6163
rect 1698 6183 1742 6221
rect 1698 6163 1710 6183
rect 1730 6163 1742 6183
rect 1698 6121 1742 6163
rect 1792 6183 1834 6221
rect 1792 6163 1806 6183
rect 1826 6163 1834 6183
rect 1792 6121 1834 6163
rect 1908 6183 1950 6221
rect 1908 6163 1916 6183
rect 1936 6163 1950 6183
rect 1908 6121 1950 6163
rect 2000 6190 2045 6221
rect 2000 6183 2044 6190
rect 2000 6163 2012 6183
rect 2032 6163 2044 6183
rect 2000 6121 2044 6163
rect 2887 6057 2931 6099
rect 2887 6037 2899 6057
rect 2919 6037 2931 6057
rect 2887 6030 2931 6037
rect 2886 5999 2931 6030
rect 2981 6057 3023 6099
rect 2981 6037 2995 6057
rect 3015 6037 3023 6057
rect 2981 5999 3023 6037
rect 3097 6057 3139 6099
rect 3097 6037 3105 6057
rect 3125 6037 3139 6057
rect 3097 5999 3139 6037
rect 3189 6057 3233 6099
rect 3189 6037 3201 6057
rect 3221 6037 3233 6057
rect 3189 5999 3233 6037
rect 3305 6057 3347 6099
rect 3305 6037 3313 6057
rect 3333 6037 3347 6057
rect 3305 5999 3347 6037
rect 3397 6057 3441 6099
rect 3397 6037 3409 6057
rect 3429 6037 3441 6057
rect 3397 5999 3441 6037
rect 3518 6057 3560 6099
rect 3518 6037 3526 6057
rect 3546 6037 3560 6057
rect 3518 5999 3560 6037
rect 3610 6057 3654 6099
rect 3610 6037 3622 6057
rect 3642 6037 3654 6057
rect 3610 5999 3654 6037
rect 338 5873 382 5911
rect 338 5853 350 5873
rect 370 5853 382 5873
rect 338 5811 382 5853
rect 432 5873 474 5911
rect 432 5853 446 5873
rect 466 5853 474 5873
rect 432 5811 474 5853
rect 551 5873 595 5911
rect 551 5853 563 5873
rect 583 5853 595 5873
rect 551 5811 595 5853
rect 645 5873 687 5911
rect 645 5853 659 5873
rect 679 5853 687 5873
rect 645 5811 687 5853
rect 759 5873 803 5911
rect 759 5853 771 5873
rect 791 5853 803 5873
rect 759 5811 803 5853
rect 853 5873 895 5911
rect 853 5853 867 5873
rect 887 5853 895 5873
rect 853 5811 895 5853
rect 969 5873 1011 5911
rect 969 5853 977 5873
rect 997 5853 1011 5873
rect 969 5811 1011 5853
rect 1061 5880 1106 5911
rect 1061 5873 1105 5880
rect 1061 5853 1073 5873
rect 1093 5853 1105 5873
rect 1061 5811 1105 5853
rect 3825 5813 3869 5855
rect 3825 5793 3837 5813
rect 3857 5793 3869 5813
rect 3825 5786 3869 5793
rect 3824 5755 3869 5786
rect 3919 5813 3961 5855
rect 3919 5793 3933 5813
rect 3953 5793 3961 5813
rect 3919 5755 3961 5793
rect 4035 5813 4077 5855
rect 4035 5793 4043 5813
rect 4063 5793 4077 5813
rect 4035 5755 4077 5793
rect 4127 5813 4171 5855
rect 4127 5793 4139 5813
rect 4159 5793 4171 5813
rect 4127 5755 4171 5793
rect 4243 5813 4285 5855
rect 4243 5793 4251 5813
rect 4271 5793 4285 5813
rect 4243 5755 4285 5793
rect 4335 5813 4379 5855
rect 4335 5793 4347 5813
rect 4367 5793 4379 5813
rect 4335 5755 4379 5793
rect 4456 5813 4498 5855
rect 4456 5793 4464 5813
rect 4484 5793 4498 5813
rect 4456 5755 4498 5793
rect 4548 5813 4592 5855
rect 4548 5793 4560 5813
rect 4580 5793 4592 5813
rect 4548 5755 4592 5793
rect 1418 5591 1462 5629
rect 1418 5571 1430 5591
rect 1450 5571 1462 5591
rect 1418 5529 1462 5571
rect 1512 5591 1554 5629
rect 1512 5571 1526 5591
rect 1546 5571 1554 5591
rect 1512 5529 1554 5571
rect 1631 5591 1675 5629
rect 1631 5571 1643 5591
rect 1663 5571 1675 5591
rect 1631 5529 1675 5571
rect 1725 5591 1767 5629
rect 1725 5571 1739 5591
rect 1759 5571 1767 5591
rect 1725 5529 1767 5571
rect 1839 5591 1883 5629
rect 1839 5571 1851 5591
rect 1871 5571 1883 5591
rect 1839 5529 1883 5571
rect 1933 5591 1975 5629
rect 1933 5571 1947 5591
rect 1967 5571 1975 5591
rect 1933 5529 1975 5571
rect 2049 5591 2091 5629
rect 2049 5571 2057 5591
rect 2077 5571 2091 5591
rect 2049 5529 2091 5571
rect 2141 5598 2186 5629
rect 2141 5591 2185 5598
rect 2141 5571 2153 5591
rect 2173 5571 2185 5591
rect 2141 5529 2185 5571
rect 2747 5546 2791 5588
rect 2747 5526 2759 5546
rect 2779 5526 2791 5546
rect 2747 5519 2791 5526
rect 2746 5488 2791 5519
rect 2841 5546 2883 5588
rect 2841 5526 2855 5546
rect 2875 5526 2883 5546
rect 2841 5488 2883 5526
rect 2957 5546 2999 5588
rect 2957 5526 2965 5546
rect 2985 5526 2999 5546
rect 2957 5488 2999 5526
rect 3049 5546 3093 5588
rect 3049 5526 3061 5546
rect 3081 5526 3093 5546
rect 3049 5488 3093 5526
rect 3165 5546 3207 5588
rect 3165 5526 3173 5546
rect 3193 5526 3207 5546
rect 3165 5488 3207 5526
rect 3257 5546 3301 5588
rect 3257 5526 3269 5546
rect 3289 5526 3301 5546
rect 3257 5488 3301 5526
rect 3378 5546 3420 5588
rect 3378 5526 3386 5546
rect 3406 5526 3420 5546
rect 3378 5488 3420 5526
rect 3470 5546 3514 5588
rect 3470 5526 3482 5546
rect 3502 5526 3514 5546
rect 3470 5488 3514 5526
rect 340 5324 384 5362
rect 340 5304 352 5324
rect 372 5304 384 5324
rect 340 5262 384 5304
rect 434 5324 476 5362
rect 434 5304 448 5324
rect 468 5304 476 5324
rect 434 5262 476 5304
rect 553 5324 597 5362
rect 553 5304 565 5324
rect 585 5304 597 5324
rect 553 5262 597 5304
rect 647 5324 689 5362
rect 647 5304 661 5324
rect 681 5304 689 5324
rect 647 5262 689 5304
rect 761 5324 805 5362
rect 761 5304 773 5324
rect 793 5304 805 5324
rect 761 5262 805 5304
rect 855 5324 897 5362
rect 855 5304 869 5324
rect 889 5304 897 5324
rect 855 5262 897 5304
rect 971 5324 1013 5362
rect 971 5304 979 5324
rect 999 5304 1013 5324
rect 971 5262 1013 5304
rect 1063 5331 1108 5362
rect 1063 5324 1107 5331
rect 1063 5304 1075 5324
rect 1095 5304 1107 5324
rect 1063 5262 1107 5304
rect 3827 5264 3871 5306
rect 3827 5244 3839 5264
rect 3859 5244 3871 5264
rect 3827 5237 3871 5244
rect 3826 5206 3871 5237
rect 3921 5264 3963 5306
rect 3921 5244 3935 5264
rect 3955 5244 3963 5264
rect 3921 5206 3963 5244
rect 4037 5264 4079 5306
rect 4037 5244 4045 5264
rect 4065 5244 4079 5264
rect 4037 5206 4079 5244
rect 4129 5264 4173 5306
rect 4129 5244 4141 5264
rect 4161 5244 4173 5264
rect 4129 5206 4173 5244
rect 4245 5264 4287 5306
rect 4245 5244 4253 5264
rect 4273 5244 4287 5264
rect 4245 5206 4287 5244
rect 4337 5264 4381 5306
rect 4337 5244 4349 5264
rect 4369 5244 4381 5264
rect 4337 5206 4381 5244
rect 4458 5264 4500 5306
rect 4458 5244 4466 5264
rect 4486 5244 4500 5264
rect 4458 5206 4500 5244
rect 4550 5264 4594 5306
rect 4550 5244 4562 5264
rect 4582 5244 4594 5264
rect 4550 5206 4594 5244
rect 1278 5080 1322 5118
rect 1278 5060 1290 5080
rect 1310 5060 1322 5080
rect 1278 5018 1322 5060
rect 1372 5080 1414 5118
rect 1372 5060 1386 5080
rect 1406 5060 1414 5080
rect 1372 5018 1414 5060
rect 1491 5080 1535 5118
rect 1491 5060 1503 5080
rect 1523 5060 1535 5080
rect 1491 5018 1535 5060
rect 1585 5080 1627 5118
rect 1585 5060 1599 5080
rect 1619 5060 1627 5080
rect 1585 5018 1627 5060
rect 1699 5080 1743 5118
rect 1699 5060 1711 5080
rect 1731 5060 1743 5080
rect 1699 5018 1743 5060
rect 1793 5080 1835 5118
rect 1793 5060 1807 5080
rect 1827 5060 1835 5080
rect 1793 5018 1835 5060
rect 1909 5080 1951 5118
rect 1909 5060 1917 5080
rect 1937 5060 1951 5080
rect 1909 5018 1951 5060
rect 2001 5087 2046 5118
rect 2001 5080 2045 5087
rect 2001 5060 2013 5080
rect 2033 5060 2045 5080
rect 2001 5018 2045 5060
rect 2888 4954 2932 4996
rect 2888 4934 2900 4954
rect 2920 4934 2932 4954
rect 2888 4927 2932 4934
rect 2887 4896 2932 4927
rect 2982 4954 3024 4996
rect 2982 4934 2996 4954
rect 3016 4934 3024 4954
rect 2982 4896 3024 4934
rect 3098 4954 3140 4996
rect 3098 4934 3106 4954
rect 3126 4934 3140 4954
rect 3098 4896 3140 4934
rect 3190 4954 3234 4996
rect 3190 4934 3202 4954
rect 3222 4934 3234 4954
rect 3190 4896 3234 4934
rect 3306 4954 3348 4996
rect 3306 4934 3314 4954
rect 3334 4934 3348 4954
rect 3306 4896 3348 4934
rect 3398 4954 3442 4996
rect 3398 4934 3410 4954
rect 3430 4934 3442 4954
rect 3398 4896 3442 4934
rect 3519 4954 3561 4996
rect 3519 4934 3527 4954
rect 3547 4934 3561 4954
rect 3519 4896 3561 4934
rect 3611 4954 3655 4996
rect 3611 4934 3623 4954
rect 3643 4934 3655 4954
rect 3611 4896 3655 4934
rect 339 4770 383 4808
rect 339 4750 351 4770
rect 371 4750 383 4770
rect 339 4708 383 4750
rect 433 4770 475 4808
rect 433 4750 447 4770
rect 467 4750 475 4770
rect 433 4708 475 4750
rect 552 4770 596 4808
rect 552 4750 564 4770
rect 584 4750 596 4770
rect 552 4708 596 4750
rect 646 4770 688 4808
rect 646 4750 660 4770
rect 680 4750 688 4770
rect 646 4708 688 4750
rect 760 4770 804 4808
rect 760 4750 772 4770
rect 792 4750 804 4770
rect 760 4708 804 4750
rect 854 4770 896 4808
rect 854 4750 868 4770
rect 888 4750 896 4770
rect 854 4708 896 4750
rect 970 4770 1012 4808
rect 970 4750 978 4770
rect 998 4750 1012 4770
rect 970 4708 1012 4750
rect 1062 4777 1107 4808
rect 1062 4770 1106 4777
rect 1062 4750 1074 4770
rect 1094 4750 1106 4770
rect 1062 4708 1106 4750
rect 3826 4710 3870 4752
rect 3826 4690 3838 4710
rect 3858 4690 3870 4710
rect 3826 4683 3870 4690
rect 3825 4652 3870 4683
rect 3920 4710 3962 4752
rect 3920 4690 3934 4710
rect 3954 4690 3962 4710
rect 3920 4652 3962 4690
rect 4036 4710 4078 4752
rect 4036 4690 4044 4710
rect 4064 4690 4078 4710
rect 4036 4652 4078 4690
rect 4128 4710 4172 4752
rect 4128 4690 4140 4710
rect 4160 4690 4172 4710
rect 4128 4652 4172 4690
rect 4244 4710 4286 4752
rect 4244 4690 4252 4710
rect 4272 4690 4286 4710
rect 4244 4652 4286 4690
rect 4336 4710 4380 4752
rect 4336 4690 4348 4710
rect 4368 4690 4380 4710
rect 4336 4652 4380 4690
rect 4457 4710 4499 4752
rect 4457 4690 4465 4710
rect 4485 4690 4499 4710
rect 4457 4652 4499 4690
rect 4549 4710 4593 4752
rect 4549 4690 4561 4710
rect 4581 4690 4593 4710
rect 4549 4652 4593 4690
rect 1387 4507 1431 4545
rect 1387 4487 1399 4507
rect 1419 4487 1431 4507
rect 1387 4445 1431 4487
rect 1481 4507 1523 4545
rect 1481 4487 1495 4507
rect 1515 4487 1523 4507
rect 1481 4445 1523 4487
rect 1600 4507 1644 4545
rect 1600 4487 1612 4507
rect 1632 4487 1644 4507
rect 1600 4445 1644 4487
rect 1694 4507 1736 4545
rect 1694 4487 1708 4507
rect 1728 4487 1736 4507
rect 1694 4445 1736 4487
rect 1808 4507 1852 4545
rect 1808 4487 1820 4507
rect 1840 4487 1852 4507
rect 1808 4445 1852 4487
rect 1902 4507 1944 4545
rect 1902 4487 1916 4507
rect 1936 4487 1944 4507
rect 1902 4445 1944 4487
rect 2018 4507 2060 4545
rect 2018 4487 2026 4507
rect 2046 4487 2060 4507
rect 2018 4445 2060 4487
rect 2110 4514 2155 4545
rect 2110 4507 2154 4514
rect 2110 4487 2122 4507
rect 2142 4487 2154 4507
rect 2110 4445 2154 4487
rect 2779 4424 2823 4466
rect 2779 4404 2791 4424
rect 2811 4404 2823 4424
rect 2779 4397 2823 4404
rect 2778 4366 2823 4397
rect 2873 4424 2915 4466
rect 2873 4404 2887 4424
rect 2907 4404 2915 4424
rect 2873 4366 2915 4404
rect 2989 4424 3031 4466
rect 2989 4404 2997 4424
rect 3017 4404 3031 4424
rect 2989 4366 3031 4404
rect 3081 4424 3125 4466
rect 3081 4404 3093 4424
rect 3113 4404 3125 4424
rect 3081 4366 3125 4404
rect 3197 4424 3239 4466
rect 3197 4404 3205 4424
rect 3225 4404 3239 4424
rect 3197 4366 3239 4404
rect 3289 4424 3333 4466
rect 3289 4404 3301 4424
rect 3321 4404 3333 4424
rect 3289 4366 3333 4404
rect 3410 4424 3452 4466
rect 3410 4404 3418 4424
rect 3438 4404 3452 4424
rect 3410 4366 3452 4404
rect 3502 4424 3546 4466
rect 3502 4404 3514 4424
rect 3534 4404 3546 4424
rect 3502 4366 3546 4404
rect 340 4221 384 4259
rect 340 4201 352 4221
rect 372 4201 384 4221
rect 340 4159 384 4201
rect 434 4221 476 4259
rect 434 4201 448 4221
rect 468 4201 476 4221
rect 434 4159 476 4201
rect 553 4221 597 4259
rect 553 4201 565 4221
rect 585 4201 597 4221
rect 553 4159 597 4201
rect 647 4221 689 4259
rect 647 4201 661 4221
rect 681 4201 689 4221
rect 647 4159 689 4201
rect 761 4221 805 4259
rect 761 4201 773 4221
rect 793 4201 805 4221
rect 761 4159 805 4201
rect 855 4221 897 4259
rect 855 4201 869 4221
rect 889 4201 897 4221
rect 855 4159 897 4201
rect 971 4221 1013 4259
rect 971 4201 979 4221
rect 999 4201 1013 4221
rect 971 4159 1013 4201
rect 1063 4228 1108 4259
rect 1063 4221 1107 4228
rect 1063 4201 1075 4221
rect 1095 4201 1107 4221
rect 1063 4159 1107 4201
rect 3827 4161 3871 4203
rect 3827 4141 3839 4161
rect 3859 4141 3871 4161
rect 3827 4134 3871 4141
rect 3826 4103 3871 4134
rect 3921 4161 3963 4203
rect 3921 4141 3935 4161
rect 3955 4141 3963 4161
rect 3921 4103 3963 4141
rect 4037 4161 4079 4203
rect 4037 4141 4045 4161
rect 4065 4141 4079 4161
rect 4037 4103 4079 4141
rect 4129 4161 4173 4203
rect 4129 4141 4141 4161
rect 4161 4141 4173 4161
rect 4129 4103 4173 4141
rect 4245 4161 4287 4203
rect 4245 4141 4253 4161
rect 4273 4141 4287 4161
rect 4245 4103 4287 4141
rect 4337 4161 4381 4203
rect 4337 4141 4349 4161
rect 4369 4141 4381 4161
rect 4337 4103 4381 4141
rect 4458 4161 4500 4203
rect 4458 4141 4466 4161
rect 4486 4141 4500 4161
rect 4458 4103 4500 4141
rect 4550 4161 4594 4203
rect 4550 4141 4562 4161
rect 4582 4141 4594 4161
rect 4550 4103 4594 4141
rect 1278 3977 1322 4015
rect 1278 3957 1290 3977
rect 1310 3957 1322 3977
rect 1278 3915 1322 3957
rect 1372 3977 1414 4015
rect 1372 3957 1386 3977
rect 1406 3957 1414 3977
rect 1372 3915 1414 3957
rect 1491 3977 1535 4015
rect 1491 3957 1503 3977
rect 1523 3957 1535 3977
rect 1491 3915 1535 3957
rect 1585 3977 1627 4015
rect 1585 3957 1599 3977
rect 1619 3957 1627 3977
rect 1585 3915 1627 3957
rect 1699 3977 1743 4015
rect 1699 3957 1711 3977
rect 1731 3957 1743 3977
rect 1699 3915 1743 3957
rect 1793 3977 1835 4015
rect 1793 3957 1807 3977
rect 1827 3957 1835 3977
rect 1793 3915 1835 3957
rect 1909 3977 1951 4015
rect 1909 3957 1917 3977
rect 1937 3957 1951 3977
rect 1909 3915 1951 3957
rect 2001 3984 2046 4015
rect 2001 3977 2045 3984
rect 2001 3957 2013 3977
rect 2033 3957 2045 3977
rect 2001 3915 2045 3957
rect 2888 3851 2932 3893
rect 2888 3831 2900 3851
rect 2920 3831 2932 3851
rect 2888 3824 2932 3831
rect 2887 3793 2932 3824
rect 2982 3851 3024 3893
rect 2982 3831 2996 3851
rect 3016 3831 3024 3851
rect 2982 3793 3024 3831
rect 3098 3851 3140 3893
rect 3098 3831 3106 3851
rect 3126 3831 3140 3851
rect 3098 3793 3140 3831
rect 3190 3851 3234 3893
rect 3190 3831 3202 3851
rect 3222 3831 3234 3851
rect 3190 3793 3234 3831
rect 3306 3851 3348 3893
rect 3306 3831 3314 3851
rect 3334 3831 3348 3851
rect 3306 3793 3348 3831
rect 3398 3851 3442 3893
rect 3398 3831 3410 3851
rect 3430 3831 3442 3851
rect 3398 3793 3442 3831
rect 3519 3851 3561 3893
rect 3519 3831 3527 3851
rect 3547 3831 3561 3851
rect 3519 3793 3561 3831
rect 3611 3851 3655 3893
rect 3611 3831 3623 3851
rect 3643 3831 3655 3851
rect 3611 3793 3655 3831
rect 339 3667 383 3705
rect 339 3647 351 3667
rect 371 3647 383 3667
rect 339 3605 383 3647
rect 433 3667 475 3705
rect 433 3647 447 3667
rect 467 3647 475 3667
rect 433 3605 475 3647
rect 552 3667 596 3705
rect 552 3647 564 3667
rect 584 3647 596 3667
rect 552 3605 596 3647
rect 646 3667 688 3705
rect 646 3647 660 3667
rect 680 3647 688 3667
rect 646 3605 688 3647
rect 760 3667 804 3705
rect 760 3647 772 3667
rect 792 3647 804 3667
rect 760 3605 804 3647
rect 854 3667 896 3705
rect 854 3647 868 3667
rect 888 3647 896 3667
rect 854 3605 896 3647
rect 970 3667 1012 3705
rect 970 3647 978 3667
rect 998 3647 1012 3667
rect 970 3605 1012 3647
rect 1062 3674 1107 3705
rect 1062 3667 1106 3674
rect 1062 3647 1074 3667
rect 1094 3647 1106 3667
rect 1062 3605 1106 3647
rect 3826 3607 3870 3649
rect 3826 3587 3838 3607
rect 3858 3587 3870 3607
rect 3826 3580 3870 3587
rect 3825 3549 3870 3580
rect 3920 3607 3962 3649
rect 3920 3587 3934 3607
rect 3954 3587 3962 3607
rect 3920 3549 3962 3587
rect 4036 3607 4078 3649
rect 4036 3587 4044 3607
rect 4064 3587 4078 3607
rect 4036 3549 4078 3587
rect 4128 3607 4172 3649
rect 4128 3587 4140 3607
rect 4160 3587 4172 3607
rect 4128 3549 4172 3587
rect 4244 3607 4286 3649
rect 4244 3587 4252 3607
rect 4272 3587 4286 3607
rect 4244 3549 4286 3587
rect 4336 3607 4380 3649
rect 4336 3587 4348 3607
rect 4368 3587 4380 3607
rect 4336 3549 4380 3587
rect 4457 3607 4499 3649
rect 4457 3587 4465 3607
rect 4485 3587 4499 3607
rect 4457 3549 4499 3587
rect 4549 3607 4593 3649
rect 4549 3587 4561 3607
rect 4581 3587 4593 3607
rect 4549 3549 4593 3587
rect 1419 3385 1463 3423
rect 1419 3365 1431 3385
rect 1451 3365 1463 3385
rect 1419 3323 1463 3365
rect 1513 3385 1555 3423
rect 1513 3365 1527 3385
rect 1547 3365 1555 3385
rect 1513 3323 1555 3365
rect 1632 3385 1676 3423
rect 1632 3365 1644 3385
rect 1664 3365 1676 3385
rect 1632 3323 1676 3365
rect 1726 3385 1768 3423
rect 1726 3365 1740 3385
rect 1760 3365 1768 3385
rect 1726 3323 1768 3365
rect 1840 3385 1884 3423
rect 1840 3365 1852 3385
rect 1872 3365 1884 3385
rect 1840 3323 1884 3365
rect 1934 3385 1976 3423
rect 1934 3365 1948 3385
rect 1968 3365 1976 3385
rect 1934 3323 1976 3365
rect 2050 3385 2092 3423
rect 2050 3365 2058 3385
rect 2078 3365 2092 3385
rect 2050 3323 2092 3365
rect 2142 3392 2187 3423
rect 2142 3385 2186 3392
rect 2142 3365 2154 3385
rect 2174 3365 2186 3385
rect 2142 3323 2186 3365
rect 2748 3340 2792 3382
rect 2748 3320 2760 3340
rect 2780 3320 2792 3340
rect 2748 3313 2792 3320
rect 2747 3282 2792 3313
rect 2842 3340 2884 3382
rect 2842 3320 2856 3340
rect 2876 3320 2884 3340
rect 2842 3282 2884 3320
rect 2958 3340 3000 3382
rect 2958 3320 2966 3340
rect 2986 3320 3000 3340
rect 2958 3282 3000 3320
rect 3050 3340 3094 3382
rect 3050 3320 3062 3340
rect 3082 3320 3094 3340
rect 3050 3282 3094 3320
rect 3166 3340 3208 3382
rect 3166 3320 3174 3340
rect 3194 3320 3208 3340
rect 3166 3282 3208 3320
rect 3258 3340 3302 3382
rect 3258 3320 3270 3340
rect 3290 3320 3302 3340
rect 3258 3282 3302 3320
rect 3379 3340 3421 3382
rect 3379 3320 3387 3340
rect 3407 3320 3421 3340
rect 3379 3282 3421 3320
rect 3471 3340 3515 3382
rect 3471 3320 3483 3340
rect 3503 3320 3515 3340
rect 3471 3282 3515 3320
rect 341 3118 385 3156
rect 341 3098 353 3118
rect 373 3098 385 3118
rect 341 3056 385 3098
rect 435 3118 477 3156
rect 435 3098 449 3118
rect 469 3098 477 3118
rect 435 3056 477 3098
rect 554 3118 598 3156
rect 554 3098 566 3118
rect 586 3098 598 3118
rect 554 3056 598 3098
rect 648 3118 690 3156
rect 648 3098 662 3118
rect 682 3098 690 3118
rect 648 3056 690 3098
rect 762 3118 806 3156
rect 762 3098 774 3118
rect 794 3098 806 3118
rect 762 3056 806 3098
rect 856 3118 898 3156
rect 856 3098 870 3118
rect 890 3098 898 3118
rect 856 3056 898 3098
rect 972 3118 1014 3156
rect 972 3098 980 3118
rect 1000 3098 1014 3118
rect 972 3056 1014 3098
rect 1064 3125 1109 3156
rect 1064 3118 1108 3125
rect 1064 3098 1076 3118
rect 1096 3098 1108 3118
rect 1064 3056 1108 3098
rect 3828 3058 3872 3100
rect 3828 3038 3840 3058
rect 3860 3038 3872 3058
rect 3828 3031 3872 3038
rect 3827 3000 3872 3031
rect 3922 3058 3964 3100
rect 3922 3038 3936 3058
rect 3956 3038 3964 3058
rect 3922 3000 3964 3038
rect 4038 3058 4080 3100
rect 4038 3038 4046 3058
rect 4066 3038 4080 3058
rect 4038 3000 4080 3038
rect 4130 3058 4174 3100
rect 4130 3038 4142 3058
rect 4162 3038 4174 3058
rect 4130 3000 4174 3038
rect 4246 3058 4288 3100
rect 4246 3038 4254 3058
rect 4274 3038 4288 3058
rect 4246 3000 4288 3038
rect 4338 3058 4382 3100
rect 4338 3038 4350 3058
rect 4370 3038 4382 3058
rect 4338 3000 4382 3038
rect 4459 3058 4501 3100
rect 4459 3038 4467 3058
rect 4487 3038 4501 3058
rect 4459 3000 4501 3038
rect 4551 3058 4595 3100
rect 4551 3038 4563 3058
rect 4583 3038 4595 3058
rect 4551 3000 4595 3038
rect 1279 2874 1323 2912
rect 1279 2854 1291 2874
rect 1311 2854 1323 2874
rect 1279 2812 1323 2854
rect 1373 2874 1415 2912
rect 1373 2854 1387 2874
rect 1407 2854 1415 2874
rect 1373 2812 1415 2854
rect 1492 2874 1536 2912
rect 1492 2854 1504 2874
rect 1524 2854 1536 2874
rect 1492 2812 1536 2854
rect 1586 2874 1628 2912
rect 1586 2854 1600 2874
rect 1620 2854 1628 2874
rect 1586 2812 1628 2854
rect 1700 2874 1744 2912
rect 1700 2854 1712 2874
rect 1732 2854 1744 2874
rect 1700 2812 1744 2854
rect 1794 2874 1836 2912
rect 1794 2854 1808 2874
rect 1828 2854 1836 2874
rect 1794 2812 1836 2854
rect 1910 2874 1952 2912
rect 1910 2854 1918 2874
rect 1938 2854 1952 2874
rect 1910 2812 1952 2854
rect 2002 2881 2047 2912
rect 2002 2874 2046 2881
rect 2002 2854 2014 2874
rect 2034 2854 2046 2874
rect 2002 2812 2046 2854
rect 2889 2748 2933 2790
rect 2889 2728 2901 2748
rect 2921 2728 2933 2748
rect 2889 2721 2933 2728
rect 2888 2690 2933 2721
rect 2983 2748 3025 2790
rect 2983 2728 2997 2748
rect 3017 2728 3025 2748
rect 2983 2690 3025 2728
rect 3099 2748 3141 2790
rect 3099 2728 3107 2748
rect 3127 2728 3141 2748
rect 3099 2690 3141 2728
rect 3191 2748 3235 2790
rect 3191 2728 3203 2748
rect 3223 2728 3235 2748
rect 3191 2690 3235 2728
rect 3307 2748 3349 2790
rect 3307 2728 3315 2748
rect 3335 2728 3349 2748
rect 3307 2690 3349 2728
rect 3399 2748 3443 2790
rect 3399 2728 3411 2748
rect 3431 2728 3443 2748
rect 3399 2690 3443 2728
rect 3520 2748 3562 2790
rect 3520 2728 3528 2748
rect 3548 2728 3562 2748
rect 3520 2690 3562 2728
rect 3612 2748 3656 2790
rect 3612 2728 3624 2748
rect 3644 2728 3656 2748
rect 3612 2690 3656 2728
rect 340 2564 384 2602
rect 340 2544 352 2564
rect 372 2544 384 2564
rect 340 2502 384 2544
rect 434 2564 476 2602
rect 434 2544 448 2564
rect 468 2544 476 2564
rect 434 2502 476 2544
rect 553 2564 597 2602
rect 553 2544 565 2564
rect 585 2544 597 2564
rect 553 2502 597 2544
rect 647 2564 689 2602
rect 647 2544 661 2564
rect 681 2544 689 2564
rect 647 2502 689 2544
rect 761 2564 805 2602
rect 761 2544 773 2564
rect 793 2544 805 2564
rect 761 2502 805 2544
rect 855 2564 897 2602
rect 855 2544 869 2564
rect 889 2544 897 2564
rect 855 2502 897 2544
rect 971 2564 1013 2602
rect 971 2544 979 2564
rect 999 2544 1013 2564
rect 971 2502 1013 2544
rect 1063 2571 1108 2602
rect 1063 2564 1107 2571
rect 1063 2544 1075 2564
rect 1095 2544 1107 2564
rect 1063 2502 1107 2544
rect 3827 2504 3871 2546
rect 3827 2484 3839 2504
rect 3859 2484 3871 2504
rect 3827 2477 3871 2484
rect 3826 2446 3871 2477
rect 3921 2504 3963 2546
rect 3921 2484 3935 2504
rect 3955 2484 3963 2504
rect 3921 2446 3963 2484
rect 4037 2504 4079 2546
rect 4037 2484 4045 2504
rect 4065 2484 4079 2504
rect 4037 2446 4079 2484
rect 4129 2504 4173 2546
rect 4129 2484 4141 2504
rect 4161 2484 4173 2504
rect 4129 2446 4173 2484
rect 4245 2504 4287 2546
rect 4245 2484 4253 2504
rect 4273 2484 4287 2504
rect 4245 2446 4287 2484
rect 4337 2504 4381 2546
rect 4337 2484 4349 2504
rect 4369 2484 4381 2504
rect 4337 2446 4381 2484
rect 4458 2504 4500 2546
rect 4458 2484 4466 2504
rect 4486 2484 4500 2504
rect 4458 2446 4500 2484
rect 4550 2504 4594 2546
rect 4550 2484 4562 2504
rect 4582 2484 4594 2504
rect 4550 2446 4594 2484
rect 1389 2295 1433 2333
rect 1389 2275 1401 2295
rect 1421 2275 1433 2295
rect 1389 2233 1433 2275
rect 1483 2295 1525 2333
rect 1483 2275 1497 2295
rect 1517 2275 1525 2295
rect 1483 2233 1525 2275
rect 1602 2295 1646 2333
rect 1602 2275 1614 2295
rect 1634 2275 1646 2295
rect 1602 2233 1646 2275
rect 1696 2295 1738 2333
rect 1696 2275 1710 2295
rect 1730 2275 1738 2295
rect 1696 2233 1738 2275
rect 1810 2295 1854 2333
rect 1810 2275 1822 2295
rect 1842 2275 1854 2295
rect 1810 2233 1854 2275
rect 1904 2295 1946 2333
rect 1904 2275 1918 2295
rect 1938 2275 1946 2295
rect 1904 2233 1946 2275
rect 2020 2295 2062 2333
rect 2020 2275 2028 2295
rect 2048 2275 2062 2295
rect 2020 2233 2062 2275
rect 2112 2302 2157 2333
rect 2112 2295 2156 2302
rect 2112 2275 2124 2295
rect 2144 2275 2156 2295
rect 2112 2233 2156 2275
rect 2779 2224 2823 2266
rect 2779 2204 2791 2224
rect 2811 2204 2823 2224
rect 2779 2197 2823 2204
rect 2778 2166 2823 2197
rect 2873 2224 2915 2266
rect 2873 2204 2887 2224
rect 2907 2204 2915 2224
rect 2873 2166 2915 2204
rect 2989 2224 3031 2266
rect 2989 2204 2997 2224
rect 3017 2204 3031 2224
rect 2989 2166 3031 2204
rect 3081 2224 3125 2266
rect 3081 2204 3093 2224
rect 3113 2204 3125 2224
rect 3081 2166 3125 2204
rect 3197 2224 3239 2266
rect 3197 2204 3205 2224
rect 3225 2204 3239 2224
rect 3197 2166 3239 2204
rect 3289 2224 3333 2266
rect 3289 2204 3301 2224
rect 3321 2204 3333 2224
rect 3289 2166 3333 2204
rect 3410 2224 3452 2266
rect 3410 2204 3418 2224
rect 3438 2204 3452 2224
rect 3410 2166 3452 2204
rect 3502 2224 3546 2266
rect 3502 2204 3514 2224
rect 3534 2204 3546 2224
rect 3502 2166 3546 2204
rect 341 2015 385 2053
rect 341 1995 353 2015
rect 373 1995 385 2015
rect 341 1953 385 1995
rect 435 2015 477 2053
rect 435 1995 449 2015
rect 469 1995 477 2015
rect 435 1953 477 1995
rect 554 2015 598 2053
rect 554 1995 566 2015
rect 586 1995 598 2015
rect 554 1953 598 1995
rect 648 2015 690 2053
rect 648 1995 662 2015
rect 682 1995 690 2015
rect 648 1953 690 1995
rect 762 2015 806 2053
rect 762 1995 774 2015
rect 794 1995 806 2015
rect 762 1953 806 1995
rect 856 2015 898 2053
rect 856 1995 870 2015
rect 890 1995 898 2015
rect 856 1953 898 1995
rect 972 2015 1014 2053
rect 972 1995 980 2015
rect 1000 1995 1014 2015
rect 972 1953 1014 1995
rect 1064 2022 1109 2053
rect 1064 2015 1108 2022
rect 1064 1995 1076 2015
rect 1096 1995 1108 2015
rect 1064 1953 1108 1995
rect 3828 1955 3872 1997
rect 3828 1935 3840 1955
rect 3860 1935 3872 1955
rect 3828 1928 3872 1935
rect 3827 1897 3872 1928
rect 3922 1955 3964 1997
rect 3922 1935 3936 1955
rect 3956 1935 3964 1955
rect 3922 1897 3964 1935
rect 4038 1955 4080 1997
rect 4038 1935 4046 1955
rect 4066 1935 4080 1955
rect 4038 1897 4080 1935
rect 4130 1955 4174 1997
rect 4130 1935 4142 1955
rect 4162 1935 4174 1955
rect 4130 1897 4174 1935
rect 4246 1955 4288 1997
rect 4246 1935 4254 1955
rect 4274 1935 4288 1955
rect 4246 1897 4288 1935
rect 4338 1955 4382 1997
rect 4338 1935 4350 1955
rect 4370 1935 4382 1955
rect 4338 1897 4382 1935
rect 4459 1955 4501 1997
rect 4459 1935 4467 1955
rect 4487 1935 4501 1955
rect 4459 1897 4501 1935
rect 4551 1955 4595 1997
rect 4551 1935 4563 1955
rect 4583 1935 4595 1955
rect 4551 1897 4595 1935
rect 1279 1771 1323 1809
rect 1279 1751 1291 1771
rect 1311 1751 1323 1771
rect 1279 1709 1323 1751
rect 1373 1771 1415 1809
rect 1373 1751 1387 1771
rect 1407 1751 1415 1771
rect 1373 1709 1415 1751
rect 1492 1771 1536 1809
rect 1492 1751 1504 1771
rect 1524 1751 1536 1771
rect 1492 1709 1536 1751
rect 1586 1771 1628 1809
rect 1586 1751 1600 1771
rect 1620 1751 1628 1771
rect 1586 1709 1628 1751
rect 1700 1771 1744 1809
rect 1700 1751 1712 1771
rect 1732 1751 1744 1771
rect 1700 1709 1744 1751
rect 1794 1771 1836 1809
rect 1794 1751 1808 1771
rect 1828 1751 1836 1771
rect 1794 1709 1836 1751
rect 1910 1771 1952 1809
rect 1910 1751 1918 1771
rect 1938 1751 1952 1771
rect 1910 1709 1952 1751
rect 2002 1778 2047 1809
rect 2002 1771 2046 1778
rect 2002 1751 2014 1771
rect 2034 1751 2046 1771
rect 2002 1709 2046 1751
rect 2889 1645 2933 1687
rect 2889 1625 2901 1645
rect 2921 1625 2933 1645
rect 2889 1618 2933 1625
rect 2888 1587 2933 1618
rect 2983 1645 3025 1687
rect 2983 1625 2997 1645
rect 3017 1625 3025 1645
rect 2983 1587 3025 1625
rect 3099 1645 3141 1687
rect 3099 1625 3107 1645
rect 3127 1625 3141 1645
rect 3099 1587 3141 1625
rect 3191 1645 3235 1687
rect 3191 1625 3203 1645
rect 3223 1625 3235 1645
rect 3191 1587 3235 1625
rect 3307 1645 3349 1687
rect 3307 1625 3315 1645
rect 3335 1625 3349 1645
rect 3307 1587 3349 1625
rect 3399 1645 3443 1687
rect 3399 1625 3411 1645
rect 3431 1625 3443 1645
rect 3399 1587 3443 1625
rect 3520 1645 3562 1687
rect 3520 1625 3528 1645
rect 3548 1625 3562 1645
rect 3520 1587 3562 1625
rect 3612 1645 3656 1687
rect 3612 1625 3624 1645
rect 3644 1625 3656 1645
rect 3612 1587 3656 1625
rect 340 1461 384 1499
rect 340 1441 352 1461
rect 372 1441 384 1461
rect 340 1399 384 1441
rect 434 1461 476 1499
rect 434 1441 448 1461
rect 468 1441 476 1461
rect 434 1399 476 1441
rect 553 1461 597 1499
rect 553 1441 565 1461
rect 585 1441 597 1461
rect 553 1399 597 1441
rect 647 1461 689 1499
rect 647 1441 661 1461
rect 681 1441 689 1461
rect 647 1399 689 1441
rect 761 1461 805 1499
rect 761 1441 773 1461
rect 793 1441 805 1461
rect 761 1399 805 1441
rect 855 1461 897 1499
rect 855 1441 869 1461
rect 889 1441 897 1461
rect 855 1399 897 1441
rect 971 1461 1013 1499
rect 971 1441 979 1461
rect 999 1441 1013 1461
rect 971 1399 1013 1441
rect 1063 1468 1108 1499
rect 1063 1461 1107 1468
rect 1063 1441 1075 1461
rect 1095 1441 1107 1461
rect 1063 1399 1107 1441
rect 3827 1401 3871 1443
rect 3827 1381 3839 1401
rect 3859 1381 3871 1401
rect 3827 1374 3871 1381
rect 3826 1343 3871 1374
rect 3921 1401 3963 1443
rect 3921 1381 3935 1401
rect 3955 1381 3963 1401
rect 3921 1343 3963 1381
rect 4037 1401 4079 1443
rect 4037 1381 4045 1401
rect 4065 1381 4079 1401
rect 4037 1343 4079 1381
rect 4129 1401 4173 1443
rect 4129 1381 4141 1401
rect 4161 1381 4173 1401
rect 4129 1343 4173 1381
rect 4245 1401 4287 1443
rect 4245 1381 4253 1401
rect 4273 1381 4287 1401
rect 4245 1343 4287 1381
rect 4337 1401 4381 1443
rect 4337 1381 4349 1401
rect 4369 1381 4381 1401
rect 4337 1343 4381 1381
rect 4458 1401 4500 1443
rect 4458 1381 4466 1401
rect 4486 1381 4500 1401
rect 4458 1343 4500 1381
rect 4550 1401 4594 1443
rect 4550 1381 4562 1401
rect 4582 1381 4594 1401
rect 4550 1343 4594 1381
rect 1420 1179 1464 1217
rect 1420 1159 1432 1179
rect 1452 1159 1464 1179
rect 1420 1117 1464 1159
rect 1514 1179 1556 1217
rect 1514 1159 1528 1179
rect 1548 1159 1556 1179
rect 1514 1117 1556 1159
rect 1633 1179 1677 1217
rect 1633 1159 1645 1179
rect 1665 1159 1677 1179
rect 1633 1117 1677 1159
rect 1727 1179 1769 1217
rect 1727 1159 1741 1179
rect 1761 1159 1769 1179
rect 1727 1117 1769 1159
rect 1841 1179 1885 1217
rect 1841 1159 1853 1179
rect 1873 1159 1885 1179
rect 1841 1117 1885 1159
rect 1935 1179 1977 1217
rect 1935 1159 1949 1179
rect 1969 1159 1977 1179
rect 1935 1117 1977 1159
rect 2051 1179 2093 1217
rect 2051 1159 2059 1179
rect 2079 1159 2093 1179
rect 2051 1117 2093 1159
rect 2143 1186 2188 1217
rect 2143 1179 2187 1186
rect 2143 1159 2155 1179
rect 2175 1159 2187 1179
rect 2143 1117 2187 1159
rect 2749 1134 2793 1176
rect 2749 1114 2761 1134
rect 2781 1114 2793 1134
rect 2749 1107 2793 1114
rect 2748 1076 2793 1107
rect 2843 1134 2885 1176
rect 2843 1114 2857 1134
rect 2877 1114 2885 1134
rect 2843 1076 2885 1114
rect 2959 1134 3001 1176
rect 2959 1114 2967 1134
rect 2987 1114 3001 1134
rect 2959 1076 3001 1114
rect 3051 1134 3095 1176
rect 3051 1114 3063 1134
rect 3083 1114 3095 1134
rect 3051 1076 3095 1114
rect 3167 1134 3209 1176
rect 3167 1114 3175 1134
rect 3195 1114 3209 1134
rect 3167 1076 3209 1114
rect 3259 1134 3303 1176
rect 3259 1114 3271 1134
rect 3291 1114 3303 1134
rect 3259 1076 3303 1114
rect 3380 1134 3422 1176
rect 3380 1114 3388 1134
rect 3408 1114 3422 1134
rect 3380 1076 3422 1114
rect 3472 1134 3516 1176
rect 3472 1114 3484 1134
rect 3504 1114 3516 1134
rect 3472 1076 3516 1114
rect 342 912 386 950
rect 342 892 354 912
rect 374 892 386 912
rect 342 850 386 892
rect 436 912 478 950
rect 436 892 450 912
rect 470 892 478 912
rect 436 850 478 892
rect 555 912 599 950
rect 555 892 567 912
rect 587 892 599 912
rect 555 850 599 892
rect 649 912 691 950
rect 649 892 663 912
rect 683 892 691 912
rect 649 850 691 892
rect 763 912 807 950
rect 763 892 775 912
rect 795 892 807 912
rect 763 850 807 892
rect 857 912 899 950
rect 857 892 871 912
rect 891 892 899 912
rect 857 850 899 892
rect 973 912 1015 950
rect 973 892 981 912
rect 1001 892 1015 912
rect 973 850 1015 892
rect 1065 919 1110 950
rect 1065 912 1109 919
rect 1065 892 1077 912
rect 1097 892 1109 912
rect 1065 850 1109 892
rect 3829 852 3873 894
rect 3829 832 3841 852
rect 3861 832 3873 852
rect 3829 825 3873 832
rect 3828 794 3873 825
rect 3923 852 3965 894
rect 3923 832 3937 852
rect 3957 832 3965 852
rect 3923 794 3965 832
rect 4039 852 4081 894
rect 4039 832 4047 852
rect 4067 832 4081 852
rect 4039 794 4081 832
rect 4131 852 4175 894
rect 4131 832 4143 852
rect 4163 832 4175 852
rect 4131 794 4175 832
rect 4247 852 4289 894
rect 4247 832 4255 852
rect 4275 832 4289 852
rect 4247 794 4289 832
rect 4339 852 4383 894
rect 4339 832 4351 852
rect 4371 832 4383 852
rect 4339 794 4383 832
rect 4460 852 4502 894
rect 4460 832 4468 852
rect 4488 832 4502 852
rect 4460 794 4502 832
rect 4552 852 4596 894
rect 4552 832 4564 852
rect 4584 832 4596 852
rect 4552 794 4596 832
rect 1280 668 1324 706
rect 1280 648 1292 668
rect 1312 648 1324 668
rect 1280 606 1324 648
rect 1374 668 1416 706
rect 1374 648 1388 668
rect 1408 648 1416 668
rect 1374 606 1416 648
rect 1493 668 1537 706
rect 1493 648 1505 668
rect 1525 648 1537 668
rect 1493 606 1537 648
rect 1587 668 1629 706
rect 1587 648 1601 668
rect 1621 648 1629 668
rect 1587 606 1629 648
rect 1701 668 1745 706
rect 1701 648 1713 668
rect 1733 648 1745 668
rect 1701 606 1745 648
rect 1795 668 1837 706
rect 1795 648 1809 668
rect 1829 648 1837 668
rect 1795 606 1837 648
rect 1911 668 1953 706
rect 1911 648 1919 668
rect 1939 648 1953 668
rect 1911 606 1953 648
rect 2003 675 2048 706
rect 2003 668 2047 675
rect 2003 648 2015 668
rect 2035 648 2047 668
rect 2003 606 2047 648
rect 2890 542 2934 584
rect 2890 522 2902 542
rect 2922 522 2934 542
rect 2890 515 2934 522
rect 2889 484 2934 515
rect 2984 542 3026 584
rect 2984 522 2998 542
rect 3018 522 3026 542
rect 2984 484 3026 522
rect 3100 542 3142 584
rect 3100 522 3108 542
rect 3128 522 3142 542
rect 3100 484 3142 522
rect 3192 542 3236 584
rect 3192 522 3204 542
rect 3224 522 3236 542
rect 3192 484 3236 522
rect 3308 542 3350 584
rect 3308 522 3316 542
rect 3336 522 3350 542
rect 3308 484 3350 522
rect 3400 542 3444 584
rect 3400 522 3412 542
rect 3432 522 3444 542
rect 3400 484 3444 522
rect 3521 542 3563 584
rect 3521 522 3529 542
rect 3549 522 3563 542
rect 3521 484 3563 522
rect 3613 542 3657 584
rect 3613 522 3625 542
rect 3645 522 3657 542
rect 3613 484 3657 522
rect 341 358 385 396
rect 341 338 353 358
rect 373 338 385 358
rect 341 296 385 338
rect 435 358 477 396
rect 435 338 449 358
rect 469 338 477 358
rect 435 296 477 338
rect 554 358 598 396
rect 554 338 566 358
rect 586 338 598 358
rect 554 296 598 338
rect 648 358 690 396
rect 648 338 662 358
rect 682 338 690 358
rect 648 296 690 338
rect 762 358 806 396
rect 762 338 774 358
rect 794 338 806 358
rect 762 296 806 338
rect 856 358 898 396
rect 856 338 870 358
rect 890 338 898 358
rect 856 296 898 338
rect 972 358 1014 396
rect 972 338 980 358
rect 1000 338 1014 358
rect 972 296 1014 338
rect 1064 365 1109 396
rect 1064 358 1108 365
rect 1064 338 1076 358
rect 1096 338 1108 358
rect 1064 296 1108 338
rect 3828 298 3872 340
rect 3828 278 3840 298
rect 3860 278 3872 298
rect 3828 271 3872 278
rect 3827 240 3872 271
rect 3922 298 3964 340
rect 3922 278 3936 298
rect 3956 278 3964 298
rect 3922 240 3964 278
rect 4038 298 4080 340
rect 4038 278 4046 298
rect 4066 278 4080 298
rect 4038 240 4080 278
rect 4130 298 4174 340
rect 4130 278 4142 298
rect 4162 278 4174 298
rect 4130 240 4174 278
rect 4246 298 4288 340
rect 4246 278 4254 298
rect 4274 278 4288 298
rect 4246 240 4288 278
rect 4338 298 4382 340
rect 4338 278 4350 298
rect 4370 278 4382 298
rect 4338 240 4382 278
rect 4459 298 4501 340
rect 4459 278 4467 298
rect 4487 278 4501 298
rect 4459 240 4501 278
rect 4551 298 4595 340
rect 4551 278 4563 298
rect 4583 278 4595 298
rect 4551 240 4595 278
rect 1588 -201 1632 -163
rect 1588 -221 1600 -201
rect 1620 -221 1632 -201
rect 1588 -263 1632 -221
rect 1682 -201 1724 -163
rect 1682 -221 1696 -201
rect 1716 -221 1724 -201
rect 1682 -263 1724 -221
rect 1801 -201 1845 -163
rect 1801 -221 1813 -201
rect 1833 -221 1845 -201
rect 1801 -263 1845 -221
rect 1895 -201 1937 -163
rect 1895 -221 1909 -201
rect 1929 -221 1937 -201
rect 1895 -263 1937 -221
rect 2009 -201 2053 -163
rect 2009 -221 2021 -201
rect 2041 -221 2053 -201
rect 2009 -263 2053 -221
rect 2103 -201 2145 -163
rect 2103 -221 2117 -201
rect 2137 -221 2145 -201
rect 2103 -263 2145 -221
rect 2219 -201 2261 -163
rect 2219 -221 2227 -201
rect 2247 -221 2261 -201
rect 2219 -263 2261 -221
rect 2311 -194 2356 -163
rect 2311 -201 2355 -194
rect 2311 -221 2323 -201
rect 2343 -221 2355 -201
rect 2311 -263 2355 -221
<< ndiffc >>
rect 116 8749 134 8767
rect 3831 8702 3851 8722
rect 3934 8698 3954 8718
rect 4042 8698 4062 8718
rect 4145 8702 4165 8722
rect 4250 8698 4270 8718
rect 4353 8702 4373 8722
rect 4463 8698 4483 8718
rect 4566 8702 4586 8722
rect 118 8650 136 8668
rect 116 8562 134 8580
rect 118 8463 136 8481
rect 344 8464 364 8484
rect 447 8468 467 8488
rect 557 8464 577 8484
rect 660 8468 680 8488
rect 765 8464 785 8484
rect 868 8468 888 8488
rect 976 8468 996 8488
rect 1079 8464 1099 8484
rect 4793 8610 4811 8628
rect 4795 8511 4813 8529
rect 116 8333 134 8351
rect 2892 8392 2912 8412
rect 2995 8388 3015 8408
rect 3103 8388 3123 8408
rect 3206 8392 3226 8412
rect 3311 8388 3331 8408
rect 3414 8392 3434 8412
rect 3524 8388 3544 8408
rect 3627 8392 3647 8412
rect 118 8234 136 8252
rect 4793 8380 4811 8398
rect 1282 8220 1302 8240
rect 1385 8224 1405 8244
rect 1495 8220 1515 8240
rect 1598 8224 1618 8244
rect 1703 8220 1723 8240
rect 1806 8224 1826 8244
rect 1914 8224 1934 8244
rect 2017 8220 2037 8240
rect 4795 8281 4813 8299
rect 116 8103 134 8121
rect 118 8004 136 8022
rect 3830 8148 3850 8168
rect 3933 8144 3953 8164
rect 4041 8144 4061 8164
rect 4144 8148 4164 8168
rect 4249 8144 4269 8164
rect 4352 8148 4372 8168
rect 4462 8144 4482 8164
rect 4565 8148 4585 8168
rect 4793 8151 4811 8169
rect 4795 8052 4813 8070
rect 4793 7964 4811 7982
rect 343 7910 363 7930
rect 446 7914 466 7934
rect 556 7910 576 7930
rect 659 7914 679 7934
rect 764 7910 784 7930
rect 867 7914 887 7934
rect 975 7914 995 7934
rect 1078 7910 1098 7930
rect 2752 7881 2772 7901
rect 2855 7877 2875 7897
rect 2963 7877 2983 7897
rect 3066 7881 3086 7901
rect 3171 7877 3191 7897
rect 3274 7881 3294 7901
rect 3384 7877 3404 7897
rect 3487 7881 3507 7901
rect 4795 7865 4813 7883
rect 117 7646 135 7664
rect 1423 7628 1443 7648
rect 1526 7632 1546 7652
rect 1636 7628 1656 7648
rect 1739 7632 1759 7652
rect 1844 7628 1864 7648
rect 1947 7632 1967 7652
rect 2055 7632 2075 7652
rect 2158 7628 2178 7648
rect 3832 7599 3852 7619
rect 3935 7595 3955 7615
rect 4043 7595 4063 7615
rect 4146 7599 4166 7619
rect 4251 7595 4271 7615
rect 4354 7599 4374 7619
rect 4464 7595 4484 7615
rect 4567 7599 4587 7619
rect 119 7547 137 7565
rect 117 7459 135 7477
rect 119 7360 137 7378
rect 345 7361 365 7381
rect 448 7365 468 7385
rect 558 7361 578 7381
rect 661 7365 681 7385
rect 766 7361 786 7381
rect 869 7365 889 7385
rect 977 7365 997 7385
rect 1080 7361 1100 7381
rect 4794 7507 4812 7525
rect 4796 7408 4814 7426
rect 117 7230 135 7248
rect 2893 7289 2913 7309
rect 2996 7285 3016 7305
rect 3104 7285 3124 7305
rect 3207 7289 3227 7309
rect 3312 7285 3332 7305
rect 3415 7289 3435 7309
rect 3525 7285 3545 7305
rect 3628 7289 3648 7309
rect 119 7131 137 7149
rect 4794 7277 4812 7295
rect 1283 7117 1303 7137
rect 1386 7121 1406 7141
rect 1496 7117 1516 7137
rect 1599 7121 1619 7141
rect 1704 7117 1724 7137
rect 1807 7121 1827 7141
rect 1915 7121 1935 7141
rect 2018 7117 2038 7137
rect 4796 7178 4814 7196
rect 117 7000 135 7018
rect 119 6901 137 6919
rect 3831 7045 3851 7065
rect 3934 7041 3954 7061
rect 4042 7041 4062 7061
rect 4145 7045 4165 7065
rect 4250 7041 4270 7061
rect 4353 7045 4373 7065
rect 4463 7041 4483 7061
rect 4566 7045 4586 7065
rect 4794 7048 4812 7066
rect 4796 6949 4814 6967
rect 4794 6861 4812 6879
rect 344 6807 364 6827
rect 447 6811 467 6831
rect 557 6807 577 6827
rect 660 6811 680 6831
rect 765 6807 785 6827
rect 868 6811 888 6831
rect 976 6811 996 6831
rect 1079 6807 1099 6827
rect 2783 6765 2803 6785
rect 2886 6761 2906 6781
rect 2994 6761 3014 6781
rect 3097 6765 3117 6785
rect 3202 6761 3222 6781
rect 3305 6765 3325 6785
rect 3415 6761 3435 6781
rect 3518 6765 3538 6785
rect 4796 6762 4814 6780
rect 117 6543 135 6561
rect 1393 6538 1413 6558
rect 1496 6542 1516 6562
rect 1606 6538 1626 6558
rect 1709 6542 1729 6562
rect 1814 6538 1834 6558
rect 1917 6542 1937 6562
rect 2025 6542 2045 6562
rect 2128 6538 2148 6558
rect 3832 6496 3852 6516
rect 3935 6492 3955 6512
rect 4043 6492 4063 6512
rect 4146 6496 4166 6516
rect 4251 6492 4271 6512
rect 4354 6496 4374 6516
rect 4464 6492 4484 6512
rect 4567 6496 4587 6516
rect 119 6444 137 6462
rect 117 6356 135 6374
rect 119 6257 137 6275
rect 345 6258 365 6278
rect 448 6262 468 6282
rect 558 6258 578 6278
rect 661 6262 681 6282
rect 766 6258 786 6278
rect 869 6262 889 6282
rect 977 6262 997 6282
rect 1080 6258 1100 6278
rect 4794 6404 4812 6422
rect 4796 6305 4814 6323
rect 117 6127 135 6145
rect 2893 6186 2913 6206
rect 2996 6182 3016 6202
rect 3104 6182 3124 6202
rect 3207 6186 3227 6206
rect 3312 6182 3332 6202
rect 3415 6186 3435 6206
rect 3525 6182 3545 6202
rect 3628 6186 3648 6206
rect 119 6028 137 6046
rect 4794 6174 4812 6192
rect 1283 6014 1303 6034
rect 1386 6018 1406 6038
rect 1496 6014 1516 6034
rect 1599 6018 1619 6038
rect 1704 6014 1724 6034
rect 1807 6018 1827 6038
rect 1915 6018 1935 6038
rect 2018 6014 2038 6034
rect 4796 6075 4814 6093
rect 117 5897 135 5915
rect 119 5798 137 5816
rect 3831 5942 3851 5962
rect 3934 5938 3954 5958
rect 4042 5938 4062 5958
rect 4145 5942 4165 5962
rect 4250 5938 4270 5958
rect 4353 5942 4373 5962
rect 4463 5938 4483 5958
rect 4566 5942 4586 5962
rect 4794 5945 4812 5963
rect 4796 5846 4814 5864
rect 4794 5758 4812 5776
rect 344 5704 364 5724
rect 447 5708 467 5728
rect 557 5704 577 5724
rect 660 5708 680 5728
rect 765 5704 785 5724
rect 868 5708 888 5728
rect 976 5708 996 5728
rect 1079 5704 1099 5724
rect 2753 5675 2773 5695
rect 2856 5671 2876 5691
rect 2964 5671 2984 5691
rect 3067 5675 3087 5695
rect 3172 5671 3192 5691
rect 3275 5675 3295 5695
rect 3385 5671 3405 5691
rect 3488 5675 3508 5695
rect 4796 5659 4814 5677
rect 118 5440 136 5458
rect 1424 5422 1444 5442
rect 1527 5426 1547 5446
rect 1637 5422 1657 5442
rect 1740 5426 1760 5446
rect 1845 5422 1865 5442
rect 1948 5426 1968 5446
rect 2056 5426 2076 5446
rect 2159 5422 2179 5442
rect 3833 5393 3853 5413
rect 3936 5389 3956 5409
rect 4044 5389 4064 5409
rect 4147 5393 4167 5413
rect 4252 5389 4272 5409
rect 4355 5393 4375 5413
rect 4465 5389 4485 5409
rect 4568 5393 4588 5413
rect 120 5341 138 5359
rect 118 5253 136 5271
rect 120 5154 138 5172
rect 346 5155 366 5175
rect 449 5159 469 5179
rect 559 5155 579 5175
rect 662 5159 682 5179
rect 767 5155 787 5175
rect 870 5159 890 5179
rect 978 5159 998 5179
rect 1081 5155 1101 5175
rect 4795 5301 4813 5319
rect 4797 5202 4815 5220
rect 118 5024 136 5042
rect 2894 5083 2914 5103
rect 2997 5079 3017 5099
rect 3105 5079 3125 5099
rect 3208 5083 3228 5103
rect 3313 5079 3333 5099
rect 3416 5083 3436 5103
rect 3526 5079 3546 5099
rect 3629 5083 3649 5103
rect 120 4925 138 4943
rect 4795 5071 4813 5089
rect 1284 4911 1304 4931
rect 1387 4915 1407 4935
rect 1497 4911 1517 4931
rect 1600 4915 1620 4935
rect 1705 4911 1725 4931
rect 1808 4915 1828 4935
rect 1916 4915 1936 4935
rect 2019 4911 2039 4931
rect 4797 4972 4815 4990
rect 118 4794 136 4812
rect 120 4695 138 4713
rect 3832 4839 3852 4859
rect 3935 4835 3955 4855
rect 4043 4835 4063 4855
rect 4146 4839 4166 4859
rect 4251 4835 4271 4855
rect 4354 4839 4374 4859
rect 4464 4835 4484 4855
rect 4567 4839 4587 4859
rect 4795 4842 4813 4860
rect 4797 4743 4815 4761
rect 4795 4655 4813 4673
rect 345 4601 365 4621
rect 448 4605 468 4625
rect 558 4601 578 4621
rect 661 4605 681 4625
rect 766 4601 786 4621
rect 869 4605 889 4625
rect 977 4605 997 4625
rect 1080 4601 1100 4621
rect 2785 4553 2805 4573
rect 2888 4549 2908 4569
rect 2996 4549 3016 4569
rect 3099 4553 3119 4573
rect 3204 4549 3224 4569
rect 3307 4553 3327 4573
rect 3417 4549 3437 4569
rect 3520 4553 3540 4573
rect 4797 4556 4815 4574
rect 118 4337 136 4355
rect 1393 4338 1413 4358
rect 1496 4342 1516 4362
rect 1606 4338 1626 4358
rect 1709 4342 1729 4362
rect 1814 4338 1834 4358
rect 1917 4342 1937 4362
rect 2025 4342 2045 4362
rect 2128 4338 2148 4358
rect 3833 4290 3853 4310
rect 3936 4286 3956 4306
rect 4044 4286 4064 4306
rect 4147 4290 4167 4310
rect 4252 4286 4272 4306
rect 4355 4290 4375 4310
rect 4465 4286 4485 4306
rect 4568 4290 4588 4310
rect 120 4238 138 4256
rect 118 4150 136 4168
rect 120 4051 138 4069
rect 346 4052 366 4072
rect 449 4056 469 4076
rect 559 4052 579 4072
rect 662 4056 682 4076
rect 767 4052 787 4072
rect 870 4056 890 4076
rect 978 4056 998 4076
rect 1081 4052 1101 4072
rect 4795 4198 4813 4216
rect 4797 4099 4815 4117
rect 118 3921 136 3939
rect 2894 3980 2914 4000
rect 2997 3976 3017 3996
rect 3105 3976 3125 3996
rect 3208 3980 3228 4000
rect 3313 3976 3333 3996
rect 3416 3980 3436 4000
rect 3526 3976 3546 3996
rect 3629 3980 3649 4000
rect 120 3822 138 3840
rect 4795 3968 4813 3986
rect 1284 3808 1304 3828
rect 1387 3812 1407 3832
rect 1497 3808 1517 3828
rect 1600 3812 1620 3832
rect 1705 3808 1725 3828
rect 1808 3812 1828 3832
rect 1916 3812 1936 3832
rect 2019 3808 2039 3828
rect 4797 3869 4815 3887
rect 118 3691 136 3709
rect 120 3592 138 3610
rect 3832 3736 3852 3756
rect 3935 3732 3955 3752
rect 4043 3732 4063 3752
rect 4146 3736 4166 3756
rect 4251 3732 4271 3752
rect 4354 3736 4374 3756
rect 4464 3732 4484 3752
rect 4567 3736 4587 3756
rect 4795 3739 4813 3757
rect 4797 3640 4815 3658
rect 4795 3552 4813 3570
rect 345 3498 365 3518
rect 448 3502 468 3522
rect 558 3498 578 3518
rect 661 3502 681 3522
rect 766 3498 786 3518
rect 869 3502 889 3522
rect 977 3502 997 3522
rect 1080 3498 1100 3518
rect 2754 3469 2774 3489
rect 2857 3465 2877 3485
rect 2965 3465 2985 3485
rect 3068 3469 3088 3489
rect 3173 3465 3193 3485
rect 3276 3469 3296 3489
rect 3386 3465 3406 3485
rect 3489 3469 3509 3489
rect 4797 3453 4815 3471
rect 119 3234 137 3252
rect 1425 3216 1445 3236
rect 1528 3220 1548 3240
rect 1638 3216 1658 3236
rect 1741 3220 1761 3240
rect 1846 3216 1866 3236
rect 1949 3220 1969 3240
rect 2057 3220 2077 3240
rect 2160 3216 2180 3236
rect 3834 3187 3854 3207
rect 3937 3183 3957 3203
rect 4045 3183 4065 3203
rect 4148 3187 4168 3207
rect 4253 3183 4273 3203
rect 4356 3187 4376 3207
rect 4466 3183 4486 3203
rect 4569 3187 4589 3207
rect 121 3135 139 3153
rect 119 3047 137 3065
rect 121 2948 139 2966
rect 347 2949 367 2969
rect 450 2953 470 2973
rect 560 2949 580 2969
rect 663 2953 683 2973
rect 768 2949 788 2969
rect 871 2953 891 2973
rect 979 2953 999 2973
rect 1082 2949 1102 2969
rect 4796 3095 4814 3113
rect 4798 2996 4816 3014
rect 119 2818 137 2836
rect 2895 2877 2915 2897
rect 2998 2873 3018 2893
rect 3106 2873 3126 2893
rect 3209 2877 3229 2897
rect 3314 2873 3334 2893
rect 3417 2877 3437 2897
rect 3527 2873 3547 2893
rect 3630 2877 3650 2897
rect 121 2719 139 2737
rect 4796 2865 4814 2883
rect 1285 2705 1305 2725
rect 1388 2709 1408 2729
rect 1498 2705 1518 2725
rect 1601 2709 1621 2729
rect 1706 2705 1726 2725
rect 1809 2709 1829 2729
rect 1917 2709 1937 2729
rect 2020 2705 2040 2725
rect 4798 2766 4816 2784
rect 119 2588 137 2606
rect 121 2489 139 2507
rect 3833 2633 3853 2653
rect 3936 2629 3956 2649
rect 4044 2629 4064 2649
rect 4147 2633 4167 2653
rect 4252 2629 4272 2649
rect 4355 2633 4375 2653
rect 4465 2629 4485 2649
rect 4568 2633 4588 2653
rect 4796 2636 4814 2654
rect 4798 2537 4816 2555
rect 4796 2449 4814 2467
rect 346 2395 366 2415
rect 449 2399 469 2419
rect 559 2395 579 2415
rect 662 2399 682 2419
rect 767 2395 787 2415
rect 870 2399 890 2419
rect 978 2399 998 2419
rect 1081 2395 1101 2415
rect 2785 2353 2805 2373
rect 2888 2349 2908 2369
rect 2996 2349 3016 2369
rect 3099 2353 3119 2373
rect 3204 2349 3224 2369
rect 3307 2353 3327 2373
rect 3417 2349 3437 2369
rect 3520 2353 3540 2373
rect 4798 2350 4816 2368
rect 119 2131 137 2149
rect 1395 2126 1415 2146
rect 1498 2130 1518 2150
rect 1608 2126 1628 2146
rect 1711 2130 1731 2150
rect 1816 2126 1836 2146
rect 1919 2130 1939 2150
rect 2027 2130 2047 2150
rect 2130 2126 2150 2146
rect 3834 2084 3854 2104
rect 3937 2080 3957 2100
rect 4045 2080 4065 2100
rect 4148 2084 4168 2104
rect 4253 2080 4273 2100
rect 4356 2084 4376 2104
rect 4466 2080 4486 2100
rect 4569 2084 4589 2104
rect 121 2032 139 2050
rect 119 1944 137 1962
rect 121 1845 139 1863
rect 347 1846 367 1866
rect 450 1850 470 1870
rect 560 1846 580 1866
rect 663 1850 683 1870
rect 768 1846 788 1866
rect 871 1850 891 1870
rect 979 1850 999 1870
rect 1082 1846 1102 1866
rect 4796 1992 4814 2010
rect 4798 1893 4816 1911
rect 119 1715 137 1733
rect 2895 1774 2915 1794
rect 2998 1770 3018 1790
rect 3106 1770 3126 1790
rect 3209 1774 3229 1794
rect 3314 1770 3334 1790
rect 3417 1774 3437 1794
rect 3527 1770 3547 1790
rect 3630 1774 3650 1794
rect 121 1616 139 1634
rect 4796 1762 4814 1780
rect 1285 1602 1305 1622
rect 1388 1606 1408 1626
rect 1498 1602 1518 1622
rect 1601 1606 1621 1626
rect 1706 1602 1726 1622
rect 1809 1606 1829 1626
rect 1917 1606 1937 1626
rect 2020 1602 2040 1622
rect 4798 1663 4816 1681
rect 119 1485 137 1503
rect 121 1386 139 1404
rect 3833 1530 3853 1550
rect 3936 1526 3956 1546
rect 4044 1526 4064 1546
rect 4147 1530 4167 1550
rect 4252 1526 4272 1546
rect 4355 1530 4375 1550
rect 4465 1526 4485 1546
rect 4568 1530 4588 1550
rect 4796 1533 4814 1551
rect 4798 1434 4816 1452
rect 4796 1346 4814 1364
rect 346 1292 366 1312
rect 449 1296 469 1316
rect 559 1292 579 1312
rect 662 1296 682 1316
rect 767 1292 787 1312
rect 870 1296 890 1316
rect 978 1296 998 1316
rect 1081 1292 1101 1312
rect 2755 1263 2775 1283
rect 2858 1259 2878 1279
rect 2966 1259 2986 1279
rect 3069 1263 3089 1283
rect 3174 1259 3194 1279
rect 3277 1263 3297 1283
rect 3387 1259 3407 1279
rect 3490 1263 3510 1283
rect 4798 1247 4816 1265
rect 120 1028 138 1046
rect 1426 1010 1446 1030
rect 1529 1014 1549 1034
rect 1639 1010 1659 1030
rect 1742 1014 1762 1034
rect 1847 1010 1867 1030
rect 1950 1014 1970 1034
rect 2058 1014 2078 1034
rect 2161 1010 2181 1030
rect 3835 981 3855 1001
rect 3938 977 3958 997
rect 4046 977 4066 997
rect 4149 981 4169 1001
rect 4254 977 4274 997
rect 4357 981 4377 1001
rect 4467 977 4487 997
rect 4570 981 4590 1001
rect 122 929 140 947
rect 120 841 138 859
rect 122 742 140 760
rect 348 743 368 763
rect 451 747 471 767
rect 561 743 581 763
rect 664 747 684 767
rect 769 743 789 763
rect 872 747 892 767
rect 980 747 1000 767
rect 1083 743 1103 763
rect 4797 889 4815 907
rect 4799 790 4817 808
rect 120 612 138 630
rect 2896 671 2916 691
rect 2999 667 3019 687
rect 3107 667 3127 687
rect 3210 671 3230 691
rect 3315 667 3335 687
rect 3418 671 3438 691
rect 3528 667 3548 687
rect 3631 671 3651 691
rect 122 513 140 531
rect 4797 659 4815 677
rect 1286 499 1306 519
rect 1389 503 1409 523
rect 1499 499 1519 519
rect 1602 503 1622 523
rect 1707 499 1727 519
rect 1810 503 1830 523
rect 1918 503 1938 523
rect 2021 499 2041 519
rect 4799 560 4817 578
rect 120 382 138 400
rect 122 283 140 301
rect 3834 427 3854 447
rect 3937 423 3957 443
rect 4045 423 4065 443
rect 4148 427 4168 447
rect 4253 423 4273 443
rect 4356 427 4376 447
rect 4466 423 4486 443
rect 4569 427 4589 447
rect 4797 430 4815 448
rect 4799 331 4817 349
rect 4797 243 4815 261
rect 347 189 367 209
rect 450 193 470 213
rect 560 189 580 209
rect 663 193 683 213
rect 768 189 788 209
rect 871 193 891 213
rect 979 193 999 213
rect 1082 189 1102 209
rect 4799 144 4817 162
rect 1594 -370 1614 -350
rect 1697 -366 1717 -346
rect 1807 -370 1827 -350
rect 1910 -366 1930 -346
rect 2015 -370 2035 -350
rect 2118 -366 2138 -346
rect 2226 -366 2246 -346
rect 2329 -370 2349 -350
<< pdiffc >>
rect 350 8613 370 8633
rect 446 8613 466 8633
rect 563 8613 583 8633
rect 659 8613 679 8633
rect 771 8613 791 8633
rect 867 8613 887 8633
rect 977 8613 997 8633
rect 1073 8613 1093 8633
rect 3837 8553 3857 8573
rect 3933 8553 3953 8573
rect 4043 8553 4063 8573
rect 4139 8553 4159 8573
rect 4251 8553 4271 8573
rect 4347 8553 4367 8573
rect 4464 8553 4484 8573
rect 4560 8553 4580 8573
rect 1288 8369 1308 8389
rect 1384 8369 1404 8389
rect 1501 8369 1521 8389
rect 1597 8369 1617 8389
rect 1709 8369 1729 8389
rect 1805 8369 1825 8389
rect 1915 8369 1935 8389
rect 2011 8369 2031 8389
rect 2898 8243 2918 8263
rect 2994 8243 3014 8263
rect 3104 8243 3124 8263
rect 3200 8243 3220 8263
rect 3312 8243 3332 8263
rect 3408 8243 3428 8263
rect 3525 8243 3545 8263
rect 3621 8243 3641 8263
rect 349 8059 369 8079
rect 445 8059 465 8079
rect 562 8059 582 8079
rect 658 8059 678 8079
rect 770 8059 790 8079
rect 866 8059 886 8079
rect 976 8059 996 8079
rect 1072 8059 1092 8079
rect 3836 7999 3856 8019
rect 3932 7999 3952 8019
rect 4042 7999 4062 8019
rect 4138 7999 4158 8019
rect 4250 7999 4270 8019
rect 4346 7999 4366 8019
rect 4463 7999 4483 8019
rect 4559 7999 4579 8019
rect 1429 7777 1449 7797
rect 1525 7777 1545 7797
rect 1642 7777 1662 7797
rect 1738 7777 1758 7797
rect 1850 7777 1870 7797
rect 1946 7777 1966 7797
rect 2056 7777 2076 7797
rect 2152 7777 2172 7797
rect 2758 7732 2778 7752
rect 2854 7732 2874 7752
rect 2964 7732 2984 7752
rect 3060 7732 3080 7752
rect 3172 7732 3192 7752
rect 3268 7732 3288 7752
rect 3385 7732 3405 7752
rect 3481 7732 3501 7752
rect 351 7510 371 7530
rect 447 7510 467 7530
rect 564 7510 584 7530
rect 660 7510 680 7530
rect 772 7510 792 7530
rect 868 7510 888 7530
rect 978 7510 998 7530
rect 1074 7510 1094 7530
rect 3838 7450 3858 7470
rect 3934 7450 3954 7470
rect 4044 7450 4064 7470
rect 4140 7450 4160 7470
rect 4252 7450 4272 7470
rect 4348 7450 4368 7470
rect 4465 7450 4485 7470
rect 4561 7450 4581 7470
rect 1289 7266 1309 7286
rect 1385 7266 1405 7286
rect 1502 7266 1522 7286
rect 1598 7266 1618 7286
rect 1710 7266 1730 7286
rect 1806 7266 1826 7286
rect 1916 7266 1936 7286
rect 2012 7266 2032 7286
rect 2899 7140 2919 7160
rect 2995 7140 3015 7160
rect 3105 7140 3125 7160
rect 3201 7140 3221 7160
rect 3313 7140 3333 7160
rect 3409 7140 3429 7160
rect 3526 7140 3546 7160
rect 3622 7140 3642 7160
rect 350 6956 370 6976
rect 446 6956 466 6976
rect 563 6956 583 6976
rect 659 6956 679 6976
rect 771 6956 791 6976
rect 867 6956 887 6976
rect 977 6956 997 6976
rect 1073 6956 1093 6976
rect 3837 6896 3857 6916
rect 3933 6896 3953 6916
rect 4043 6896 4063 6916
rect 4139 6896 4159 6916
rect 4251 6896 4271 6916
rect 4347 6896 4367 6916
rect 4464 6896 4484 6916
rect 4560 6896 4580 6916
rect 1399 6687 1419 6707
rect 1495 6687 1515 6707
rect 1612 6687 1632 6707
rect 1708 6687 1728 6707
rect 1820 6687 1840 6707
rect 1916 6687 1936 6707
rect 2026 6687 2046 6707
rect 2122 6687 2142 6707
rect 2789 6616 2809 6636
rect 2885 6616 2905 6636
rect 2995 6616 3015 6636
rect 3091 6616 3111 6636
rect 3203 6616 3223 6636
rect 3299 6616 3319 6636
rect 3416 6616 3436 6636
rect 3512 6616 3532 6636
rect 351 6407 371 6427
rect 447 6407 467 6427
rect 564 6407 584 6427
rect 660 6407 680 6427
rect 772 6407 792 6427
rect 868 6407 888 6427
rect 978 6407 998 6427
rect 1074 6407 1094 6427
rect 3838 6347 3858 6367
rect 3934 6347 3954 6367
rect 4044 6347 4064 6367
rect 4140 6347 4160 6367
rect 4252 6347 4272 6367
rect 4348 6347 4368 6367
rect 4465 6347 4485 6367
rect 4561 6347 4581 6367
rect 1289 6163 1309 6183
rect 1385 6163 1405 6183
rect 1502 6163 1522 6183
rect 1598 6163 1618 6183
rect 1710 6163 1730 6183
rect 1806 6163 1826 6183
rect 1916 6163 1936 6183
rect 2012 6163 2032 6183
rect 2899 6037 2919 6057
rect 2995 6037 3015 6057
rect 3105 6037 3125 6057
rect 3201 6037 3221 6057
rect 3313 6037 3333 6057
rect 3409 6037 3429 6057
rect 3526 6037 3546 6057
rect 3622 6037 3642 6057
rect 350 5853 370 5873
rect 446 5853 466 5873
rect 563 5853 583 5873
rect 659 5853 679 5873
rect 771 5853 791 5873
rect 867 5853 887 5873
rect 977 5853 997 5873
rect 1073 5853 1093 5873
rect 3837 5793 3857 5813
rect 3933 5793 3953 5813
rect 4043 5793 4063 5813
rect 4139 5793 4159 5813
rect 4251 5793 4271 5813
rect 4347 5793 4367 5813
rect 4464 5793 4484 5813
rect 4560 5793 4580 5813
rect 1430 5571 1450 5591
rect 1526 5571 1546 5591
rect 1643 5571 1663 5591
rect 1739 5571 1759 5591
rect 1851 5571 1871 5591
rect 1947 5571 1967 5591
rect 2057 5571 2077 5591
rect 2153 5571 2173 5591
rect 2759 5526 2779 5546
rect 2855 5526 2875 5546
rect 2965 5526 2985 5546
rect 3061 5526 3081 5546
rect 3173 5526 3193 5546
rect 3269 5526 3289 5546
rect 3386 5526 3406 5546
rect 3482 5526 3502 5546
rect 352 5304 372 5324
rect 448 5304 468 5324
rect 565 5304 585 5324
rect 661 5304 681 5324
rect 773 5304 793 5324
rect 869 5304 889 5324
rect 979 5304 999 5324
rect 1075 5304 1095 5324
rect 3839 5244 3859 5264
rect 3935 5244 3955 5264
rect 4045 5244 4065 5264
rect 4141 5244 4161 5264
rect 4253 5244 4273 5264
rect 4349 5244 4369 5264
rect 4466 5244 4486 5264
rect 4562 5244 4582 5264
rect 1290 5060 1310 5080
rect 1386 5060 1406 5080
rect 1503 5060 1523 5080
rect 1599 5060 1619 5080
rect 1711 5060 1731 5080
rect 1807 5060 1827 5080
rect 1917 5060 1937 5080
rect 2013 5060 2033 5080
rect 2900 4934 2920 4954
rect 2996 4934 3016 4954
rect 3106 4934 3126 4954
rect 3202 4934 3222 4954
rect 3314 4934 3334 4954
rect 3410 4934 3430 4954
rect 3527 4934 3547 4954
rect 3623 4934 3643 4954
rect 351 4750 371 4770
rect 447 4750 467 4770
rect 564 4750 584 4770
rect 660 4750 680 4770
rect 772 4750 792 4770
rect 868 4750 888 4770
rect 978 4750 998 4770
rect 1074 4750 1094 4770
rect 3838 4690 3858 4710
rect 3934 4690 3954 4710
rect 4044 4690 4064 4710
rect 4140 4690 4160 4710
rect 4252 4690 4272 4710
rect 4348 4690 4368 4710
rect 4465 4690 4485 4710
rect 4561 4690 4581 4710
rect 1399 4487 1419 4507
rect 1495 4487 1515 4507
rect 1612 4487 1632 4507
rect 1708 4487 1728 4507
rect 1820 4487 1840 4507
rect 1916 4487 1936 4507
rect 2026 4487 2046 4507
rect 2122 4487 2142 4507
rect 2791 4404 2811 4424
rect 2887 4404 2907 4424
rect 2997 4404 3017 4424
rect 3093 4404 3113 4424
rect 3205 4404 3225 4424
rect 3301 4404 3321 4424
rect 3418 4404 3438 4424
rect 3514 4404 3534 4424
rect 352 4201 372 4221
rect 448 4201 468 4221
rect 565 4201 585 4221
rect 661 4201 681 4221
rect 773 4201 793 4221
rect 869 4201 889 4221
rect 979 4201 999 4221
rect 1075 4201 1095 4221
rect 3839 4141 3859 4161
rect 3935 4141 3955 4161
rect 4045 4141 4065 4161
rect 4141 4141 4161 4161
rect 4253 4141 4273 4161
rect 4349 4141 4369 4161
rect 4466 4141 4486 4161
rect 4562 4141 4582 4161
rect 1290 3957 1310 3977
rect 1386 3957 1406 3977
rect 1503 3957 1523 3977
rect 1599 3957 1619 3977
rect 1711 3957 1731 3977
rect 1807 3957 1827 3977
rect 1917 3957 1937 3977
rect 2013 3957 2033 3977
rect 2900 3831 2920 3851
rect 2996 3831 3016 3851
rect 3106 3831 3126 3851
rect 3202 3831 3222 3851
rect 3314 3831 3334 3851
rect 3410 3831 3430 3851
rect 3527 3831 3547 3851
rect 3623 3831 3643 3851
rect 351 3647 371 3667
rect 447 3647 467 3667
rect 564 3647 584 3667
rect 660 3647 680 3667
rect 772 3647 792 3667
rect 868 3647 888 3667
rect 978 3647 998 3667
rect 1074 3647 1094 3667
rect 3838 3587 3858 3607
rect 3934 3587 3954 3607
rect 4044 3587 4064 3607
rect 4140 3587 4160 3607
rect 4252 3587 4272 3607
rect 4348 3587 4368 3607
rect 4465 3587 4485 3607
rect 4561 3587 4581 3607
rect 1431 3365 1451 3385
rect 1527 3365 1547 3385
rect 1644 3365 1664 3385
rect 1740 3365 1760 3385
rect 1852 3365 1872 3385
rect 1948 3365 1968 3385
rect 2058 3365 2078 3385
rect 2154 3365 2174 3385
rect 2760 3320 2780 3340
rect 2856 3320 2876 3340
rect 2966 3320 2986 3340
rect 3062 3320 3082 3340
rect 3174 3320 3194 3340
rect 3270 3320 3290 3340
rect 3387 3320 3407 3340
rect 3483 3320 3503 3340
rect 353 3098 373 3118
rect 449 3098 469 3118
rect 566 3098 586 3118
rect 662 3098 682 3118
rect 774 3098 794 3118
rect 870 3098 890 3118
rect 980 3098 1000 3118
rect 1076 3098 1096 3118
rect 3840 3038 3860 3058
rect 3936 3038 3956 3058
rect 4046 3038 4066 3058
rect 4142 3038 4162 3058
rect 4254 3038 4274 3058
rect 4350 3038 4370 3058
rect 4467 3038 4487 3058
rect 4563 3038 4583 3058
rect 1291 2854 1311 2874
rect 1387 2854 1407 2874
rect 1504 2854 1524 2874
rect 1600 2854 1620 2874
rect 1712 2854 1732 2874
rect 1808 2854 1828 2874
rect 1918 2854 1938 2874
rect 2014 2854 2034 2874
rect 2901 2728 2921 2748
rect 2997 2728 3017 2748
rect 3107 2728 3127 2748
rect 3203 2728 3223 2748
rect 3315 2728 3335 2748
rect 3411 2728 3431 2748
rect 3528 2728 3548 2748
rect 3624 2728 3644 2748
rect 352 2544 372 2564
rect 448 2544 468 2564
rect 565 2544 585 2564
rect 661 2544 681 2564
rect 773 2544 793 2564
rect 869 2544 889 2564
rect 979 2544 999 2564
rect 1075 2544 1095 2564
rect 3839 2484 3859 2504
rect 3935 2484 3955 2504
rect 4045 2484 4065 2504
rect 4141 2484 4161 2504
rect 4253 2484 4273 2504
rect 4349 2484 4369 2504
rect 4466 2484 4486 2504
rect 4562 2484 4582 2504
rect 1401 2275 1421 2295
rect 1497 2275 1517 2295
rect 1614 2275 1634 2295
rect 1710 2275 1730 2295
rect 1822 2275 1842 2295
rect 1918 2275 1938 2295
rect 2028 2275 2048 2295
rect 2124 2275 2144 2295
rect 2791 2204 2811 2224
rect 2887 2204 2907 2224
rect 2997 2204 3017 2224
rect 3093 2204 3113 2224
rect 3205 2204 3225 2224
rect 3301 2204 3321 2224
rect 3418 2204 3438 2224
rect 3514 2204 3534 2224
rect 353 1995 373 2015
rect 449 1995 469 2015
rect 566 1995 586 2015
rect 662 1995 682 2015
rect 774 1995 794 2015
rect 870 1995 890 2015
rect 980 1995 1000 2015
rect 1076 1995 1096 2015
rect 3840 1935 3860 1955
rect 3936 1935 3956 1955
rect 4046 1935 4066 1955
rect 4142 1935 4162 1955
rect 4254 1935 4274 1955
rect 4350 1935 4370 1955
rect 4467 1935 4487 1955
rect 4563 1935 4583 1955
rect 1291 1751 1311 1771
rect 1387 1751 1407 1771
rect 1504 1751 1524 1771
rect 1600 1751 1620 1771
rect 1712 1751 1732 1771
rect 1808 1751 1828 1771
rect 1918 1751 1938 1771
rect 2014 1751 2034 1771
rect 2901 1625 2921 1645
rect 2997 1625 3017 1645
rect 3107 1625 3127 1645
rect 3203 1625 3223 1645
rect 3315 1625 3335 1645
rect 3411 1625 3431 1645
rect 3528 1625 3548 1645
rect 3624 1625 3644 1645
rect 352 1441 372 1461
rect 448 1441 468 1461
rect 565 1441 585 1461
rect 661 1441 681 1461
rect 773 1441 793 1461
rect 869 1441 889 1461
rect 979 1441 999 1461
rect 1075 1441 1095 1461
rect 3839 1381 3859 1401
rect 3935 1381 3955 1401
rect 4045 1381 4065 1401
rect 4141 1381 4161 1401
rect 4253 1381 4273 1401
rect 4349 1381 4369 1401
rect 4466 1381 4486 1401
rect 4562 1381 4582 1401
rect 1432 1159 1452 1179
rect 1528 1159 1548 1179
rect 1645 1159 1665 1179
rect 1741 1159 1761 1179
rect 1853 1159 1873 1179
rect 1949 1159 1969 1179
rect 2059 1159 2079 1179
rect 2155 1159 2175 1179
rect 2761 1114 2781 1134
rect 2857 1114 2877 1134
rect 2967 1114 2987 1134
rect 3063 1114 3083 1134
rect 3175 1114 3195 1134
rect 3271 1114 3291 1134
rect 3388 1114 3408 1134
rect 3484 1114 3504 1134
rect 354 892 374 912
rect 450 892 470 912
rect 567 892 587 912
rect 663 892 683 912
rect 775 892 795 912
rect 871 892 891 912
rect 981 892 1001 912
rect 1077 892 1097 912
rect 3841 832 3861 852
rect 3937 832 3957 852
rect 4047 832 4067 852
rect 4143 832 4163 852
rect 4255 832 4275 852
rect 4351 832 4371 852
rect 4468 832 4488 852
rect 4564 832 4584 852
rect 1292 648 1312 668
rect 1388 648 1408 668
rect 1505 648 1525 668
rect 1601 648 1621 668
rect 1713 648 1733 668
rect 1809 648 1829 668
rect 1919 648 1939 668
rect 2015 648 2035 668
rect 2902 522 2922 542
rect 2998 522 3018 542
rect 3108 522 3128 542
rect 3204 522 3224 542
rect 3316 522 3336 542
rect 3412 522 3432 542
rect 3529 522 3549 542
rect 3625 522 3645 542
rect 353 338 373 358
rect 449 338 469 358
rect 566 338 586 358
rect 662 338 682 358
rect 774 338 794 358
rect 870 338 890 358
rect 980 338 1000 358
rect 1076 338 1096 358
rect 3840 278 3860 298
rect 3936 278 3956 298
rect 4046 278 4066 298
rect 4142 278 4162 298
rect 4254 278 4274 298
rect 4350 278 4370 298
rect 4467 278 4487 298
rect 4563 278 4583 298
rect 1600 -221 1620 -201
rect 1696 -221 1716 -201
rect 1813 -221 1833 -201
rect 1909 -221 1929 -201
rect 2021 -221 2041 -201
rect 2117 -221 2137 -201
rect 2227 -221 2247 -201
rect 2323 -221 2343 -201
<< psubdiff >>
rect 4401 8819 4512 8834
rect 4401 8789 4443 8819
rect 4471 8789 4512 8819
rect 4401 8775 4512 8789
rect 3462 8509 3573 8524
rect 3462 8479 3504 8509
rect 3532 8479 3573 8509
rect 3462 8465 3573 8479
rect 418 8397 529 8411
rect 418 8367 459 8397
rect 487 8367 529 8397
rect 418 8352 529 8367
rect 4400 8265 4511 8280
rect 4400 8235 4442 8265
rect 4470 8235 4511 8265
rect 4400 8221 4511 8235
rect 1356 8153 1467 8167
rect 1356 8123 1397 8153
rect 1425 8123 1467 8153
rect 1356 8108 1467 8123
rect 3322 7998 3433 8013
rect 3322 7968 3364 7998
rect 3392 7968 3433 7998
rect 3322 7954 3433 7968
rect 417 7843 528 7857
rect 417 7813 458 7843
rect 486 7813 528 7843
rect 417 7798 528 7813
rect 4402 7716 4513 7731
rect 4402 7686 4444 7716
rect 4472 7686 4513 7716
rect 4402 7672 4513 7686
rect 1497 7561 1608 7575
rect 1497 7531 1538 7561
rect 1566 7531 1608 7561
rect 1497 7516 1608 7531
rect 3463 7406 3574 7421
rect 3463 7376 3505 7406
rect 3533 7376 3574 7406
rect 3463 7362 3574 7376
rect 419 7294 530 7308
rect 419 7264 460 7294
rect 488 7264 530 7294
rect 419 7249 530 7264
rect 4401 7162 4512 7177
rect 4401 7132 4443 7162
rect 4471 7132 4512 7162
rect 4401 7118 4512 7132
rect 1357 7050 1468 7064
rect 1357 7020 1398 7050
rect 1426 7020 1468 7050
rect 1357 7005 1468 7020
rect 3353 6882 3464 6897
rect 3353 6852 3395 6882
rect 3423 6852 3464 6882
rect 3353 6838 3464 6852
rect 418 6740 529 6754
rect 418 6710 459 6740
rect 487 6710 529 6740
rect 418 6696 529 6710
rect 4402 6613 4513 6627
rect 4402 6583 4444 6613
rect 4472 6583 4513 6613
rect 4402 6569 4513 6583
rect 1467 6471 1578 6485
rect 1467 6441 1508 6471
rect 1536 6441 1578 6471
rect 1467 6426 1578 6441
rect 3463 6303 3574 6318
rect 3463 6273 3505 6303
rect 3533 6273 3574 6303
rect 3463 6259 3574 6273
rect 419 6191 530 6205
rect 419 6161 460 6191
rect 488 6161 530 6191
rect 419 6146 530 6161
rect 4401 6059 4512 6074
rect 4401 6029 4443 6059
rect 4471 6029 4512 6059
rect 4401 6015 4512 6029
rect 1357 5947 1468 5961
rect 1357 5917 1398 5947
rect 1426 5917 1468 5947
rect 1357 5902 1468 5917
rect 3323 5792 3434 5807
rect 3323 5762 3365 5792
rect 3393 5762 3434 5792
rect 3323 5748 3434 5762
rect 418 5637 529 5651
rect 418 5607 459 5637
rect 487 5607 529 5637
rect 418 5592 529 5607
rect 4403 5510 4514 5525
rect 4403 5480 4445 5510
rect 4473 5480 4514 5510
rect 4403 5466 4514 5480
rect 1498 5355 1609 5369
rect 1498 5325 1539 5355
rect 1567 5325 1609 5355
rect 1498 5310 1609 5325
rect 3464 5200 3575 5215
rect 3464 5170 3506 5200
rect 3534 5170 3575 5200
rect 3464 5156 3575 5170
rect 420 5088 531 5102
rect 420 5058 461 5088
rect 489 5058 531 5088
rect 420 5043 531 5058
rect 4402 4956 4513 4971
rect 4402 4926 4444 4956
rect 4472 4926 4513 4956
rect 4402 4912 4513 4926
rect 1358 4844 1469 4858
rect 1358 4814 1399 4844
rect 1427 4814 1469 4844
rect 1358 4799 1469 4814
rect 3355 4670 3466 4685
rect 3355 4640 3397 4670
rect 3425 4640 3466 4670
rect 3355 4626 3466 4640
rect 419 4534 530 4548
rect 419 4504 460 4534
rect 488 4504 530 4534
rect 419 4489 530 4504
rect 4403 4407 4514 4422
rect 4403 4377 4445 4407
rect 4473 4377 4514 4407
rect 4403 4363 4514 4377
rect 1467 4271 1578 4285
rect 1467 4241 1508 4271
rect 1536 4241 1578 4271
rect 1467 4226 1578 4241
rect 3464 4097 3575 4112
rect 3464 4067 3506 4097
rect 3534 4067 3575 4097
rect 3464 4053 3575 4067
rect 420 3985 531 3999
rect 420 3955 461 3985
rect 489 3955 531 3985
rect 420 3940 531 3955
rect 4402 3853 4513 3868
rect 4402 3823 4444 3853
rect 4472 3823 4513 3853
rect 4402 3809 4513 3823
rect 1358 3741 1469 3755
rect 1358 3711 1399 3741
rect 1427 3711 1469 3741
rect 1358 3696 1469 3711
rect 3324 3586 3435 3601
rect 3324 3556 3366 3586
rect 3394 3556 3435 3586
rect 3324 3542 3435 3556
rect 419 3431 530 3445
rect 419 3401 460 3431
rect 488 3401 530 3431
rect 419 3386 530 3401
rect 4404 3304 4515 3319
rect 4404 3274 4446 3304
rect 4474 3274 4515 3304
rect 4404 3260 4515 3274
rect 1499 3149 1610 3163
rect 1499 3119 1540 3149
rect 1568 3119 1610 3149
rect 1499 3104 1610 3119
rect 3465 2994 3576 3009
rect 3465 2964 3507 2994
rect 3535 2964 3576 2994
rect 3465 2950 3576 2964
rect 421 2882 532 2896
rect 421 2852 462 2882
rect 490 2852 532 2882
rect 421 2837 532 2852
rect 4403 2750 4514 2765
rect 4403 2720 4445 2750
rect 4473 2720 4514 2750
rect 4403 2706 4514 2720
rect 1359 2638 1470 2652
rect 1359 2608 1400 2638
rect 1428 2608 1470 2638
rect 1359 2593 1470 2608
rect 3355 2470 3466 2485
rect 3355 2440 3397 2470
rect 3425 2440 3466 2470
rect 3355 2426 3466 2440
rect 420 2328 531 2342
rect 420 2298 461 2328
rect 489 2298 531 2328
rect 420 2284 531 2298
rect 4404 2201 4515 2215
rect 4404 2171 4446 2201
rect 4474 2171 4515 2201
rect 4404 2157 4515 2171
rect 1469 2059 1580 2073
rect 1469 2029 1510 2059
rect 1538 2029 1580 2059
rect 1469 2014 1580 2029
rect 3465 1891 3576 1906
rect 3465 1861 3507 1891
rect 3535 1861 3576 1891
rect 3465 1847 3576 1861
rect 421 1779 532 1793
rect 421 1749 462 1779
rect 490 1749 532 1779
rect 421 1734 532 1749
rect 4403 1647 4514 1662
rect 4403 1617 4445 1647
rect 4473 1617 4514 1647
rect 4403 1603 4514 1617
rect 1359 1535 1470 1549
rect 1359 1505 1400 1535
rect 1428 1505 1470 1535
rect 1359 1490 1470 1505
rect 3325 1380 3436 1395
rect 3325 1350 3367 1380
rect 3395 1350 3436 1380
rect 3325 1336 3436 1350
rect 420 1225 531 1239
rect 420 1195 461 1225
rect 489 1195 531 1225
rect 420 1180 531 1195
rect 4405 1098 4516 1113
rect 4405 1068 4447 1098
rect 4475 1068 4516 1098
rect 4405 1054 4516 1068
rect 1500 943 1611 957
rect 1500 913 1541 943
rect 1569 913 1611 943
rect 1500 898 1611 913
rect 3466 788 3577 803
rect 3466 758 3508 788
rect 3536 758 3577 788
rect 3466 744 3577 758
rect 422 676 533 690
rect 422 646 463 676
rect 491 646 533 676
rect 422 631 533 646
rect 4404 544 4515 559
rect 4404 514 4446 544
rect 4474 514 4515 544
rect 4404 500 4515 514
rect 1360 432 1471 446
rect 1360 402 1401 432
rect 1429 402 1471 432
rect 1360 387 1471 402
rect 421 122 532 136
rect 421 92 462 122
rect 490 116 532 122
rect 490 92 531 116
rect 421 77 531 92
rect 1668 -437 1779 -423
rect 1668 -467 1709 -437
rect 1737 -467 1779 -437
rect 1668 -482 1779 -467
<< nsubdiff >>
rect 419 8744 529 8758
rect 419 8714 462 8744
rect 490 8714 529 8744
rect 419 8699 529 8714
rect 1357 8500 1467 8514
rect 1357 8470 1400 8500
rect 1428 8470 1467 8500
rect 1357 8455 1467 8470
rect 4401 8472 4511 8487
rect 4401 8442 4440 8472
rect 4468 8442 4511 8472
rect 4401 8428 4511 8442
rect 418 8190 528 8204
rect 418 8160 461 8190
rect 489 8160 528 8190
rect 418 8145 528 8160
rect 3462 8162 3572 8177
rect 3462 8132 3501 8162
rect 3529 8132 3572 8162
rect 3462 8118 3572 8132
rect 1498 7908 1608 7922
rect 4400 7918 4510 7933
rect 1498 7878 1541 7908
rect 1569 7878 1608 7908
rect 1498 7863 1608 7878
rect 4400 7888 4439 7918
rect 4467 7888 4510 7918
rect 4400 7874 4510 7888
rect 420 7641 530 7655
rect 420 7611 463 7641
rect 491 7611 530 7641
rect 3322 7651 3432 7666
rect 3322 7621 3361 7651
rect 3389 7621 3432 7651
rect 420 7596 530 7611
rect 3322 7607 3432 7621
rect 1358 7397 1468 7411
rect 1358 7367 1401 7397
rect 1429 7367 1468 7397
rect 1358 7352 1468 7367
rect 4402 7369 4512 7384
rect 4402 7339 4441 7369
rect 4469 7339 4512 7369
rect 4402 7325 4512 7339
rect 419 7087 529 7101
rect 419 7057 462 7087
rect 490 7057 529 7087
rect 419 7042 529 7057
rect 3463 7059 3573 7074
rect 3463 7029 3502 7059
rect 3530 7029 3573 7059
rect 3463 7015 3573 7029
rect 1468 6818 1578 6832
rect 1468 6788 1511 6818
rect 1539 6788 1578 6818
rect 4401 6815 4511 6830
rect 1468 6773 1578 6788
rect 4401 6785 4440 6815
rect 4468 6785 4511 6815
rect 4401 6771 4511 6785
rect 420 6538 530 6552
rect 420 6508 463 6538
rect 491 6508 530 6538
rect 3353 6535 3463 6550
rect 420 6493 530 6508
rect 3353 6505 3392 6535
rect 3420 6505 3463 6535
rect 3353 6491 3463 6505
rect 1358 6294 1468 6308
rect 1358 6264 1401 6294
rect 1429 6264 1468 6294
rect 1358 6249 1468 6264
rect 4402 6266 4512 6281
rect 4402 6236 4441 6266
rect 4469 6236 4512 6266
rect 4402 6222 4512 6236
rect 419 5984 529 5998
rect 419 5954 462 5984
rect 490 5954 529 5984
rect 419 5939 529 5954
rect 3463 5956 3573 5971
rect 3463 5926 3502 5956
rect 3530 5926 3573 5956
rect 3463 5912 3573 5926
rect 1499 5702 1609 5716
rect 4401 5712 4511 5727
rect 1499 5672 1542 5702
rect 1570 5672 1609 5702
rect 1499 5657 1609 5672
rect 4401 5682 4440 5712
rect 4468 5682 4511 5712
rect 4401 5668 4511 5682
rect 421 5435 531 5449
rect 421 5405 464 5435
rect 492 5405 531 5435
rect 3323 5445 3433 5460
rect 3323 5415 3362 5445
rect 3390 5415 3433 5445
rect 421 5390 531 5405
rect 3323 5401 3433 5415
rect 1359 5191 1469 5205
rect 1359 5161 1402 5191
rect 1430 5161 1469 5191
rect 1359 5146 1469 5161
rect 4403 5163 4513 5178
rect 4403 5133 4442 5163
rect 4470 5133 4513 5163
rect 4403 5119 4513 5133
rect 420 4881 530 4895
rect 420 4851 463 4881
rect 491 4851 530 4881
rect 420 4836 530 4851
rect 3464 4853 3574 4868
rect 3464 4823 3503 4853
rect 3531 4823 3574 4853
rect 3464 4809 3574 4823
rect 1468 4618 1578 4632
rect 1468 4588 1511 4618
rect 1539 4588 1578 4618
rect 4402 4609 4512 4624
rect 1468 4573 1578 4588
rect 4402 4579 4441 4609
rect 4469 4579 4512 4609
rect 4402 4565 4512 4579
rect 421 4332 531 4346
rect 421 4302 464 4332
rect 492 4302 531 4332
rect 3355 4323 3465 4338
rect 421 4287 531 4302
rect 3355 4293 3394 4323
rect 3422 4293 3465 4323
rect 3355 4279 3465 4293
rect 1359 4088 1469 4102
rect 1359 4058 1402 4088
rect 1430 4058 1469 4088
rect 1359 4043 1469 4058
rect 4403 4060 4513 4075
rect 4403 4030 4442 4060
rect 4470 4030 4513 4060
rect 4403 4016 4513 4030
rect 420 3778 530 3792
rect 420 3748 463 3778
rect 491 3748 530 3778
rect 420 3733 530 3748
rect 3464 3750 3574 3765
rect 3464 3720 3503 3750
rect 3531 3720 3574 3750
rect 3464 3706 3574 3720
rect 1500 3496 1610 3510
rect 4402 3506 4512 3521
rect 1500 3466 1543 3496
rect 1571 3466 1610 3496
rect 1500 3451 1610 3466
rect 4402 3476 4441 3506
rect 4469 3476 4512 3506
rect 4402 3462 4512 3476
rect 422 3229 532 3243
rect 422 3199 465 3229
rect 493 3199 532 3229
rect 3324 3239 3434 3254
rect 3324 3209 3363 3239
rect 3391 3209 3434 3239
rect 422 3184 532 3199
rect 3324 3195 3434 3209
rect 1360 2985 1470 2999
rect 1360 2955 1403 2985
rect 1431 2955 1470 2985
rect 1360 2940 1470 2955
rect 4404 2957 4514 2972
rect 4404 2927 4443 2957
rect 4471 2927 4514 2957
rect 4404 2913 4514 2927
rect 421 2675 531 2689
rect 421 2645 464 2675
rect 492 2645 531 2675
rect 421 2630 531 2645
rect 3465 2647 3575 2662
rect 3465 2617 3504 2647
rect 3532 2617 3575 2647
rect 3465 2603 3575 2617
rect 1470 2406 1580 2420
rect 1470 2376 1513 2406
rect 1541 2376 1580 2406
rect 4403 2403 4513 2418
rect 1470 2361 1580 2376
rect 4403 2373 4442 2403
rect 4470 2373 4513 2403
rect 4403 2359 4513 2373
rect 422 2126 532 2140
rect 422 2096 465 2126
rect 493 2096 532 2126
rect 3355 2123 3465 2138
rect 422 2081 532 2096
rect 3355 2093 3394 2123
rect 3422 2093 3465 2123
rect 3355 2079 3465 2093
rect 1360 1882 1470 1896
rect 1360 1852 1403 1882
rect 1431 1852 1470 1882
rect 1360 1837 1470 1852
rect 4404 1854 4514 1869
rect 4404 1824 4443 1854
rect 4471 1824 4514 1854
rect 4404 1810 4514 1824
rect 421 1572 531 1586
rect 421 1542 464 1572
rect 492 1542 531 1572
rect 421 1527 531 1542
rect 3465 1544 3575 1559
rect 3465 1514 3504 1544
rect 3532 1514 3575 1544
rect 3465 1500 3575 1514
rect 1501 1290 1611 1304
rect 4403 1300 4513 1315
rect 1501 1260 1544 1290
rect 1572 1260 1611 1290
rect 1501 1245 1611 1260
rect 4403 1270 4442 1300
rect 4470 1270 4513 1300
rect 4403 1256 4513 1270
rect 423 1023 533 1037
rect 423 993 466 1023
rect 494 993 533 1023
rect 3325 1033 3435 1048
rect 3325 1003 3364 1033
rect 3392 1003 3435 1033
rect 423 978 533 993
rect 3325 989 3435 1003
rect 1361 779 1471 793
rect 1361 749 1404 779
rect 1432 749 1471 779
rect 1361 734 1471 749
rect 4405 751 4515 766
rect 4405 721 4444 751
rect 4472 721 4515 751
rect 4405 707 4515 721
rect 422 469 532 483
rect 422 439 465 469
rect 493 439 532 469
rect 422 424 532 439
rect 3466 441 3576 456
rect 3466 411 3505 441
rect 3533 411 3576 441
rect 3466 397 3576 411
rect 4404 197 4514 212
rect 4404 167 4443 197
rect 4471 167 4514 197
rect 4404 153 4514 167
rect 1669 -90 1779 -76
rect 1669 -120 1712 -90
rect 1740 -120 1779 -90
rect 1669 -135 1779 -120
<< psubdiffcont >>
rect 4443 8789 4471 8819
rect 3504 8479 3532 8509
rect 459 8367 487 8397
rect 4442 8235 4470 8265
rect 1397 8123 1425 8153
rect 3364 7968 3392 7998
rect 458 7813 486 7843
rect 4444 7686 4472 7716
rect 1538 7531 1566 7561
rect 3505 7376 3533 7406
rect 460 7264 488 7294
rect 4443 7132 4471 7162
rect 1398 7020 1426 7050
rect 3395 6852 3423 6882
rect 459 6710 487 6740
rect 4444 6583 4472 6613
rect 1508 6441 1536 6471
rect 3505 6273 3533 6303
rect 460 6161 488 6191
rect 4443 6029 4471 6059
rect 1398 5917 1426 5947
rect 3365 5762 3393 5792
rect 459 5607 487 5637
rect 4445 5480 4473 5510
rect 1539 5325 1567 5355
rect 3506 5170 3534 5200
rect 461 5058 489 5088
rect 4444 4926 4472 4956
rect 1399 4814 1427 4844
rect 3397 4640 3425 4670
rect 460 4504 488 4534
rect 4445 4377 4473 4407
rect 1508 4241 1536 4271
rect 3506 4067 3534 4097
rect 461 3955 489 3985
rect 4444 3823 4472 3853
rect 1399 3711 1427 3741
rect 3366 3556 3394 3586
rect 460 3401 488 3431
rect 4446 3274 4474 3304
rect 1540 3119 1568 3149
rect 3507 2964 3535 2994
rect 462 2852 490 2882
rect 4445 2720 4473 2750
rect 1400 2608 1428 2638
rect 3397 2440 3425 2470
rect 461 2298 489 2328
rect 4446 2171 4474 2201
rect 1510 2029 1538 2059
rect 3507 1861 3535 1891
rect 462 1749 490 1779
rect 4445 1617 4473 1647
rect 1400 1505 1428 1535
rect 3367 1350 3395 1380
rect 461 1195 489 1225
rect 4447 1068 4475 1098
rect 1541 913 1569 943
rect 3508 758 3536 788
rect 463 646 491 676
rect 4446 514 4474 544
rect 1401 402 1429 432
rect 462 92 490 122
rect 1709 -467 1737 -437
<< nsubdiffcont >>
rect 462 8714 490 8744
rect 1400 8470 1428 8500
rect 4440 8442 4468 8472
rect 461 8160 489 8190
rect 3501 8132 3529 8162
rect 1541 7878 1569 7908
rect 4439 7888 4467 7918
rect 463 7611 491 7641
rect 3361 7621 3389 7651
rect 1401 7367 1429 7397
rect 4441 7339 4469 7369
rect 462 7057 490 7087
rect 3502 7029 3530 7059
rect 1511 6788 1539 6818
rect 4440 6785 4468 6815
rect 463 6508 491 6538
rect 3392 6505 3420 6535
rect 1401 6264 1429 6294
rect 4441 6236 4469 6266
rect 462 5954 490 5984
rect 3502 5926 3530 5956
rect 1542 5672 1570 5702
rect 4440 5682 4468 5712
rect 464 5405 492 5435
rect 3362 5415 3390 5445
rect 1402 5161 1430 5191
rect 4442 5133 4470 5163
rect 463 4851 491 4881
rect 3503 4823 3531 4853
rect 1511 4588 1539 4618
rect 4441 4579 4469 4609
rect 464 4302 492 4332
rect 3394 4293 3422 4323
rect 1402 4058 1430 4088
rect 4442 4030 4470 4060
rect 463 3748 491 3778
rect 3503 3720 3531 3750
rect 1543 3466 1571 3496
rect 4441 3476 4469 3506
rect 465 3199 493 3229
rect 3363 3209 3391 3239
rect 1403 2955 1431 2985
rect 4443 2927 4471 2957
rect 464 2645 492 2675
rect 3504 2617 3532 2647
rect 1513 2376 1541 2406
rect 4442 2373 4470 2403
rect 465 2096 493 2126
rect 3394 2093 3422 2123
rect 1403 1852 1431 1882
rect 4443 1824 4471 1854
rect 464 1542 492 1572
rect 3504 1514 3532 1544
rect 1544 1260 1572 1290
rect 4442 1270 4470 1300
rect 466 993 494 1023
rect 3364 1003 3392 1033
rect 1404 749 1432 779
rect 4444 721 4472 751
rect 465 439 493 469
rect 3505 411 3533 441
rect 4443 167 4471 197
rect 1712 -120 1740 -90
<< poly >>
rect 3869 8734 3919 8750
rect 4077 8734 4127 8750
rect 4285 8734 4335 8750
rect 4498 8734 4548 8750
rect 382 8671 432 8684
rect 595 8671 645 8684
rect 803 8671 853 8684
rect 1011 8671 1061 8684
rect 3869 8667 3919 8692
rect 3869 8641 3875 8667
rect 3901 8641 3919 8667
rect 3869 8615 3919 8641
rect 4077 8663 4127 8692
rect 4077 8639 4091 8663
rect 4115 8639 4127 8663
rect 4077 8615 4127 8639
rect 4285 8668 4335 8692
rect 4285 8644 4300 8668
rect 4324 8644 4335 8668
rect 4285 8615 4335 8644
rect 4498 8663 4548 8692
rect 4498 8643 4515 8663
rect 4535 8643 4548 8663
rect 4498 8615 4548 8643
rect 382 8543 432 8571
rect 382 8523 395 8543
rect 415 8523 432 8543
rect 382 8494 432 8523
rect 595 8542 645 8571
rect 595 8518 606 8542
rect 630 8518 645 8542
rect 595 8494 645 8518
rect 803 8547 853 8571
rect 803 8523 815 8547
rect 839 8523 853 8547
rect 803 8494 853 8523
rect 1011 8545 1061 8571
rect 1011 8519 1029 8545
rect 1055 8519 1061 8545
rect 1011 8494 1061 8519
rect 3869 8502 3919 8515
rect 4077 8502 4127 8515
rect 4285 8502 4335 8515
rect 4498 8502 4548 8515
rect 382 8436 432 8452
rect 595 8436 645 8452
rect 803 8436 853 8452
rect 1011 8436 1061 8452
rect 1320 8427 1370 8440
rect 1533 8427 1583 8440
rect 1741 8427 1791 8440
rect 1949 8427 1999 8440
rect 2930 8424 2980 8440
rect 3138 8424 3188 8440
rect 3346 8424 3396 8440
rect 3559 8424 3609 8440
rect 2930 8357 2980 8382
rect 2930 8331 2936 8357
rect 2962 8331 2980 8357
rect 1320 8299 1370 8327
rect 1320 8279 1333 8299
rect 1353 8279 1370 8299
rect 1320 8250 1370 8279
rect 1533 8298 1583 8327
rect 1533 8274 1544 8298
rect 1568 8274 1583 8298
rect 1533 8250 1583 8274
rect 1741 8303 1791 8327
rect 1741 8279 1753 8303
rect 1777 8279 1791 8303
rect 1741 8250 1791 8279
rect 1949 8301 1999 8327
rect 2930 8305 2980 8331
rect 3138 8353 3188 8382
rect 3138 8329 3152 8353
rect 3176 8329 3188 8353
rect 3138 8305 3188 8329
rect 3346 8358 3396 8382
rect 3346 8334 3361 8358
rect 3385 8334 3396 8358
rect 3346 8305 3396 8334
rect 3559 8353 3609 8382
rect 3559 8333 3576 8353
rect 3596 8333 3609 8353
rect 3559 8305 3609 8333
rect 1949 8275 1967 8301
rect 1993 8275 1999 8301
rect 1949 8250 1999 8275
rect 1320 8192 1370 8208
rect 1533 8192 1583 8208
rect 1741 8192 1791 8208
rect 1949 8192 1999 8208
rect 2930 8192 2980 8205
rect 3138 8192 3188 8205
rect 3346 8192 3396 8205
rect 3559 8192 3609 8205
rect 3868 8180 3918 8196
rect 4076 8180 4126 8196
rect 4284 8180 4334 8196
rect 4497 8180 4547 8196
rect 381 8117 431 8130
rect 594 8117 644 8130
rect 802 8117 852 8130
rect 1010 8117 1060 8130
rect 3868 8113 3918 8138
rect 3868 8087 3874 8113
rect 3900 8087 3918 8113
rect 3868 8061 3918 8087
rect 4076 8109 4126 8138
rect 4076 8085 4090 8109
rect 4114 8085 4126 8109
rect 4076 8061 4126 8085
rect 4284 8114 4334 8138
rect 4284 8090 4299 8114
rect 4323 8090 4334 8114
rect 4284 8061 4334 8090
rect 4497 8109 4547 8138
rect 4497 8089 4514 8109
rect 4534 8089 4547 8109
rect 4497 8061 4547 8089
rect 381 7989 431 8017
rect 381 7969 394 7989
rect 414 7969 431 7989
rect 381 7940 431 7969
rect 594 7988 644 8017
rect 594 7964 605 7988
rect 629 7964 644 7988
rect 594 7940 644 7964
rect 802 7993 852 8017
rect 802 7969 814 7993
rect 838 7969 852 7993
rect 802 7940 852 7969
rect 1010 7991 1060 8017
rect 1010 7965 1028 7991
rect 1054 7965 1060 7991
rect 1010 7940 1060 7965
rect 3868 7948 3918 7961
rect 4076 7948 4126 7961
rect 4284 7948 4334 7961
rect 4497 7948 4547 7961
rect 2790 7913 2840 7929
rect 2998 7913 3048 7929
rect 3206 7913 3256 7929
rect 3419 7913 3469 7929
rect 381 7882 431 7898
rect 594 7882 644 7898
rect 802 7882 852 7898
rect 1010 7882 1060 7898
rect 1461 7835 1511 7848
rect 1674 7835 1724 7848
rect 1882 7835 1932 7848
rect 2090 7835 2140 7848
rect 2790 7846 2840 7871
rect 2790 7820 2796 7846
rect 2822 7820 2840 7846
rect 2790 7794 2840 7820
rect 2998 7842 3048 7871
rect 2998 7818 3012 7842
rect 3036 7818 3048 7842
rect 2998 7794 3048 7818
rect 3206 7847 3256 7871
rect 3206 7823 3221 7847
rect 3245 7823 3256 7847
rect 3206 7794 3256 7823
rect 3419 7842 3469 7871
rect 3419 7822 3436 7842
rect 3456 7822 3469 7842
rect 3419 7794 3469 7822
rect 1461 7707 1511 7735
rect 1461 7687 1474 7707
rect 1494 7687 1511 7707
rect 1461 7658 1511 7687
rect 1674 7706 1724 7735
rect 1674 7682 1685 7706
rect 1709 7682 1724 7706
rect 1674 7658 1724 7682
rect 1882 7711 1932 7735
rect 1882 7687 1894 7711
rect 1918 7687 1932 7711
rect 1882 7658 1932 7687
rect 2090 7709 2140 7735
rect 2090 7683 2108 7709
rect 2134 7683 2140 7709
rect 2090 7658 2140 7683
rect 2790 7681 2840 7694
rect 2998 7681 3048 7694
rect 3206 7681 3256 7694
rect 3419 7681 3469 7694
rect 3870 7631 3920 7647
rect 4078 7631 4128 7647
rect 4286 7631 4336 7647
rect 4499 7631 4549 7647
rect 1461 7600 1511 7616
rect 1674 7600 1724 7616
rect 1882 7600 1932 7616
rect 2090 7600 2140 7616
rect 383 7568 433 7581
rect 596 7568 646 7581
rect 804 7568 854 7581
rect 1012 7568 1062 7581
rect 3870 7564 3920 7589
rect 3870 7538 3876 7564
rect 3902 7538 3920 7564
rect 3870 7512 3920 7538
rect 4078 7560 4128 7589
rect 4078 7536 4092 7560
rect 4116 7536 4128 7560
rect 4078 7512 4128 7536
rect 4286 7565 4336 7589
rect 4286 7541 4301 7565
rect 4325 7541 4336 7565
rect 4286 7512 4336 7541
rect 4499 7560 4549 7589
rect 4499 7540 4516 7560
rect 4536 7540 4549 7560
rect 4499 7512 4549 7540
rect 383 7440 433 7468
rect 383 7420 396 7440
rect 416 7420 433 7440
rect 383 7391 433 7420
rect 596 7439 646 7468
rect 596 7415 607 7439
rect 631 7415 646 7439
rect 596 7391 646 7415
rect 804 7444 854 7468
rect 804 7420 816 7444
rect 840 7420 854 7444
rect 804 7391 854 7420
rect 1012 7442 1062 7468
rect 1012 7416 1030 7442
rect 1056 7416 1062 7442
rect 1012 7391 1062 7416
rect 3870 7399 3920 7412
rect 4078 7399 4128 7412
rect 4286 7399 4336 7412
rect 4499 7399 4549 7412
rect 383 7333 433 7349
rect 596 7333 646 7349
rect 804 7333 854 7349
rect 1012 7333 1062 7349
rect 1321 7324 1371 7337
rect 1534 7324 1584 7337
rect 1742 7324 1792 7337
rect 1950 7324 2000 7337
rect 2931 7321 2981 7337
rect 3139 7321 3189 7337
rect 3347 7321 3397 7337
rect 3560 7321 3610 7337
rect 2931 7254 2981 7279
rect 2931 7228 2937 7254
rect 2963 7228 2981 7254
rect 1321 7196 1371 7224
rect 1321 7176 1334 7196
rect 1354 7176 1371 7196
rect 1321 7147 1371 7176
rect 1534 7195 1584 7224
rect 1534 7171 1545 7195
rect 1569 7171 1584 7195
rect 1534 7147 1584 7171
rect 1742 7200 1792 7224
rect 1742 7176 1754 7200
rect 1778 7176 1792 7200
rect 1742 7147 1792 7176
rect 1950 7198 2000 7224
rect 2931 7202 2981 7228
rect 3139 7250 3189 7279
rect 3139 7226 3153 7250
rect 3177 7226 3189 7250
rect 3139 7202 3189 7226
rect 3347 7255 3397 7279
rect 3347 7231 3362 7255
rect 3386 7231 3397 7255
rect 3347 7202 3397 7231
rect 3560 7250 3610 7279
rect 3560 7230 3577 7250
rect 3597 7230 3610 7250
rect 3560 7202 3610 7230
rect 1950 7172 1968 7198
rect 1994 7172 2000 7198
rect 1950 7147 2000 7172
rect 1321 7089 1371 7105
rect 1534 7089 1584 7105
rect 1742 7089 1792 7105
rect 1950 7089 2000 7105
rect 2931 7089 2981 7102
rect 3139 7089 3189 7102
rect 3347 7089 3397 7102
rect 3560 7089 3610 7102
rect 3869 7077 3919 7093
rect 4077 7077 4127 7093
rect 4285 7077 4335 7093
rect 4498 7077 4548 7093
rect 382 7014 432 7027
rect 595 7014 645 7027
rect 803 7014 853 7027
rect 1011 7014 1061 7027
rect 3869 7010 3919 7035
rect 3869 6984 3875 7010
rect 3901 6984 3919 7010
rect 3869 6958 3919 6984
rect 4077 7006 4127 7035
rect 4077 6982 4091 7006
rect 4115 6982 4127 7006
rect 4077 6958 4127 6982
rect 4285 7011 4335 7035
rect 4285 6987 4300 7011
rect 4324 6987 4335 7011
rect 4285 6958 4335 6987
rect 4498 7006 4548 7035
rect 4498 6986 4515 7006
rect 4535 6986 4548 7006
rect 4498 6958 4548 6986
rect 382 6886 432 6914
rect 382 6866 395 6886
rect 415 6866 432 6886
rect 382 6837 432 6866
rect 595 6885 645 6914
rect 595 6861 606 6885
rect 630 6861 645 6885
rect 595 6837 645 6861
rect 803 6890 853 6914
rect 803 6866 815 6890
rect 839 6866 853 6890
rect 803 6837 853 6866
rect 1011 6888 1061 6914
rect 1011 6862 1029 6888
rect 1055 6862 1061 6888
rect 1011 6837 1061 6862
rect 3869 6845 3919 6858
rect 4077 6845 4127 6858
rect 4285 6845 4335 6858
rect 4498 6845 4548 6858
rect 382 6779 432 6795
rect 595 6779 645 6795
rect 803 6779 853 6795
rect 1011 6779 1061 6795
rect 2821 6797 2871 6813
rect 3029 6797 3079 6813
rect 3237 6797 3287 6813
rect 3450 6797 3500 6813
rect 1431 6745 1481 6758
rect 1644 6745 1694 6758
rect 1852 6745 1902 6758
rect 2060 6745 2110 6758
rect 2821 6730 2871 6755
rect 2821 6704 2827 6730
rect 2853 6704 2871 6730
rect 2821 6678 2871 6704
rect 3029 6726 3079 6755
rect 3029 6702 3043 6726
rect 3067 6702 3079 6726
rect 3029 6678 3079 6702
rect 3237 6731 3287 6755
rect 3237 6707 3252 6731
rect 3276 6707 3287 6731
rect 3237 6678 3287 6707
rect 3450 6726 3500 6755
rect 3450 6706 3467 6726
rect 3487 6706 3500 6726
rect 3450 6678 3500 6706
rect 1431 6617 1481 6645
rect 1431 6597 1444 6617
rect 1464 6597 1481 6617
rect 1431 6568 1481 6597
rect 1644 6616 1694 6645
rect 1644 6592 1655 6616
rect 1679 6592 1694 6616
rect 1644 6568 1694 6592
rect 1852 6621 1902 6645
rect 1852 6597 1864 6621
rect 1888 6597 1902 6621
rect 1852 6568 1902 6597
rect 2060 6619 2110 6645
rect 2060 6593 2078 6619
rect 2104 6593 2110 6619
rect 2060 6568 2110 6593
rect 2821 6565 2871 6578
rect 3029 6565 3079 6578
rect 3237 6565 3287 6578
rect 3450 6565 3500 6578
rect 1431 6510 1481 6526
rect 1644 6510 1694 6526
rect 1852 6510 1902 6526
rect 2060 6510 2110 6526
rect 3870 6528 3920 6544
rect 4078 6528 4128 6544
rect 4286 6528 4336 6544
rect 4499 6528 4549 6544
rect 383 6465 433 6478
rect 596 6465 646 6478
rect 804 6465 854 6478
rect 1012 6465 1062 6478
rect 3870 6461 3920 6486
rect 3870 6435 3876 6461
rect 3902 6435 3920 6461
rect 3870 6409 3920 6435
rect 4078 6457 4128 6486
rect 4078 6433 4092 6457
rect 4116 6433 4128 6457
rect 4078 6409 4128 6433
rect 4286 6462 4336 6486
rect 4286 6438 4301 6462
rect 4325 6438 4336 6462
rect 4286 6409 4336 6438
rect 4499 6457 4549 6486
rect 4499 6437 4516 6457
rect 4536 6437 4549 6457
rect 4499 6409 4549 6437
rect 383 6337 433 6365
rect 383 6317 396 6337
rect 416 6317 433 6337
rect 383 6288 433 6317
rect 596 6336 646 6365
rect 596 6312 607 6336
rect 631 6312 646 6336
rect 596 6288 646 6312
rect 804 6341 854 6365
rect 804 6317 816 6341
rect 840 6317 854 6341
rect 804 6288 854 6317
rect 1012 6339 1062 6365
rect 1012 6313 1030 6339
rect 1056 6313 1062 6339
rect 1012 6288 1062 6313
rect 3870 6296 3920 6309
rect 4078 6296 4128 6309
rect 4286 6296 4336 6309
rect 4499 6296 4549 6309
rect 383 6230 433 6246
rect 596 6230 646 6246
rect 804 6230 854 6246
rect 1012 6230 1062 6246
rect 1321 6221 1371 6234
rect 1534 6221 1584 6234
rect 1742 6221 1792 6234
rect 1950 6221 2000 6234
rect 2931 6218 2981 6234
rect 3139 6218 3189 6234
rect 3347 6218 3397 6234
rect 3560 6218 3610 6234
rect 2931 6151 2981 6176
rect 2931 6125 2937 6151
rect 2963 6125 2981 6151
rect 1321 6093 1371 6121
rect 1321 6073 1334 6093
rect 1354 6073 1371 6093
rect 1321 6044 1371 6073
rect 1534 6092 1584 6121
rect 1534 6068 1545 6092
rect 1569 6068 1584 6092
rect 1534 6044 1584 6068
rect 1742 6097 1792 6121
rect 1742 6073 1754 6097
rect 1778 6073 1792 6097
rect 1742 6044 1792 6073
rect 1950 6095 2000 6121
rect 2931 6099 2981 6125
rect 3139 6147 3189 6176
rect 3139 6123 3153 6147
rect 3177 6123 3189 6147
rect 3139 6099 3189 6123
rect 3347 6152 3397 6176
rect 3347 6128 3362 6152
rect 3386 6128 3397 6152
rect 3347 6099 3397 6128
rect 3560 6147 3610 6176
rect 3560 6127 3577 6147
rect 3597 6127 3610 6147
rect 3560 6099 3610 6127
rect 1950 6069 1968 6095
rect 1994 6069 2000 6095
rect 1950 6044 2000 6069
rect 1321 5986 1371 6002
rect 1534 5986 1584 6002
rect 1742 5986 1792 6002
rect 1950 5986 2000 6002
rect 2931 5986 2981 5999
rect 3139 5986 3189 5999
rect 3347 5986 3397 5999
rect 3560 5986 3610 5999
rect 3869 5974 3919 5990
rect 4077 5974 4127 5990
rect 4285 5974 4335 5990
rect 4498 5974 4548 5990
rect 382 5911 432 5924
rect 595 5911 645 5924
rect 803 5911 853 5924
rect 1011 5911 1061 5924
rect 3869 5907 3919 5932
rect 3869 5881 3875 5907
rect 3901 5881 3919 5907
rect 3869 5855 3919 5881
rect 4077 5903 4127 5932
rect 4077 5879 4091 5903
rect 4115 5879 4127 5903
rect 4077 5855 4127 5879
rect 4285 5908 4335 5932
rect 4285 5884 4300 5908
rect 4324 5884 4335 5908
rect 4285 5855 4335 5884
rect 4498 5903 4548 5932
rect 4498 5883 4515 5903
rect 4535 5883 4548 5903
rect 4498 5855 4548 5883
rect 382 5783 432 5811
rect 382 5763 395 5783
rect 415 5763 432 5783
rect 382 5734 432 5763
rect 595 5782 645 5811
rect 595 5758 606 5782
rect 630 5758 645 5782
rect 595 5734 645 5758
rect 803 5787 853 5811
rect 803 5763 815 5787
rect 839 5763 853 5787
rect 803 5734 853 5763
rect 1011 5785 1061 5811
rect 1011 5759 1029 5785
rect 1055 5759 1061 5785
rect 1011 5734 1061 5759
rect 3869 5742 3919 5755
rect 4077 5742 4127 5755
rect 4285 5742 4335 5755
rect 4498 5742 4548 5755
rect 2791 5707 2841 5723
rect 2999 5707 3049 5723
rect 3207 5707 3257 5723
rect 3420 5707 3470 5723
rect 382 5676 432 5692
rect 595 5676 645 5692
rect 803 5676 853 5692
rect 1011 5676 1061 5692
rect 1462 5629 1512 5642
rect 1675 5629 1725 5642
rect 1883 5629 1933 5642
rect 2091 5629 2141 5642
rect 2791 5640 2841 5665
rect 2791 5614 2797 5640
rect 2823 5614 2841 5640
rect 2791 5588 2841 5614
rect 2999 5636 3049 5665
rect 2999 5612 3013 5636
rect 3037 5612 3049 5636
rect 2999 5588 3049 5612
rect 3207 5641 3257 5665
rect 3207 5617 3222 5641
rect 3246 5617 3257 5641
rect 3207 5588 3257 5617
rect 3420 5636 3470 5665
rect 3420 5616 3437 5636
rect 3457 5616 3470 5636
rect 3420 5588 3470 5616
rect 1462 5501 1512 5529
rect 1462 5481 1475 5501
rect 1495 5481 1512 5501
rect 1462 5452 1512 5481
rect 1675 5500 1725 5529
rect 1675 5476 1686 5500
rect 1710 5476 1725 5500
rect 1675 5452 1725 5476
rect 1883 5505 1933 5529
rect 1883 5481 1895 5505
rect 1919 5481 1933 5505
rect 1883 5452 1933 5481
rect 2091 5503 2141 5529
rect 2091 5477 2109 5503
rect 2135 5477 2141 5503
rect 2091 5452 2141 5477
rect 2791 5475 2841 5488
rect 2999 5475 3049 5488
rect 3207 5475 3257 5488
rect 3420 5475 3470 5488
rect 3871 5425 3921 5441
rect 4079 5425 4129 5441
rect 4287 5425 4337 5441
rect 4500 5425 4550 5441
rect 1462 5394 1512 5410
rect 1675 5394 1725 5410
rect 1883 5394 1933 5410
rect 2091 5394 2141 5410
rect 384 5362 434 5375
rect 597 5362 647 5375
rect 805 5362 855 5375
rect 1013 5362 1063 5375
rect 3871 5358 3921 5383
rect 3871 5332 3877 5358
rect 3903 5332 3921 5358
rect 3871 5306 3921 5332
rect 4079 5354 4129 5383
rect 4079 5330 4093 5354
rect 4117 5330 4129 5354
rect 4079 5306 4129 5330
rect 4287 5359 4337 5383
rect 4287 5335 4302 5359
rect 4326 5335 4337 5359
rect 4287 5306 4337 5335
rect 4500 5354 4550 5383
rect 4500 5334 4517 5354
rect 4537 5334 4550 5354
rect 4500 5306 4550 5334
rect 384 5234 434 5262
rect 384 5214 397 5234
rect 417 5214 434 5234
rect 384 5185 434 5214
rect 597 5233 647 5262
rect 597 5209 608 5233
rect 632 5209 647 5233
rect 597 5185 647 5209
rect 805 5238 855 5262
rect 805 5214 817 5238
rect 841 5214 855 5238
rect 805 5185 855 5214
rect 1013 5236 1063 5262
rect 1013 5210 1031 5236
rect 1057 5210 1063 5236
rect 1013 5185 1063 5210
rect 3871 5193 3921 5206
rect 4079 5193 4129 5206
rect 4287 5193 4337 5206
rect 4500 5193 4550 5206
rect 384 5127 434 5143
rect 597 5127 647 5143
rect 805 5127 855 5143
rect 1013 5127 1063 5143
rect 1322 5118 1372 5131
rect 1535 5118 1585 5131
rect 1743 5118 1793 5131
rect 1951 5118 2001 5131
rect 2932 5115 2982 5131
rect 3140 5115 3190 5131
rect 3348 5115 3398 5131
rect 3561 5115 3611 5131
rect 2932 5048 2982 5073
rect 2932 5022 2938 5048
rect 2964 5022 2982 5048
rect 1322 4990 1372 5018
rect 1322 4970 1335 4990
rect 1355 4970 1372 4990
rect 1322 4941 1372 4970
rect 1535 4989 1585 5018
rect 1535 4965 1546 4989
rect 1570 4965 1585 4989
rect 1535 4941 1585 4965
rect 1743 4994 1793 5018
rect 1743 4970 1755 4994
rect 1779 4970 1793 4994
rect 1743 4941 1793 4970
rect 1951 4992 2001 5018
rect 2932 4996 2982 5022
rect 3140 5044 3190 5073
rect 3140 5020 3154 5044
rect 3178 5020 3190 5044
rect 3140 4996 3190 5020
rect 3348 5049 3398 5073
rect 3348 5025 3363 5049
rect 3387 5025 3398 5049
rect 3348 4996 3398 5025
rect 3561 5044 3611 5073
rect 3561 5024 3578 5044
rect 3598 5024 3611 5044
rect 3561 4996 3611 5024
rect 1951 4966 1969 4992
rect 1995 4966 2001 4992
rect 1951 4941 2001 4966
rect 1322 4883 1372 4899
rect 1535 4883 1585 4899
rect 1743 4883 1793 4899
rect 1951 4883 2001 4899
rect 2932 4883 2982 4896
rect 3140 4883 3190 4896
rect 3348 4883 3398 4896
rect 3561 4883 3611 4896
rect 3870 4871 3920 4887
rect 4078 4871 4128 4887
rect 4286 4871 4336 4887
rect 4499 4871 4549 4887
rect 383 4808 433 4821
rect 596 4808 646 4821
rect 804 4808 854 4821
rect 1012 4808 1062 4821
rect 3870 4804 3920 4829
rect 3870 4778 3876 4804
rect 3902 4778 3920 4804
rect 3870 4752 3920 4778
rect 4078 4800 4128 4829
rect 4078 4776 4092 4800
rect 4116 4776 4128 4800
rect 4078 4752 4128 4776
rect 4286 4805 4336 4829
rect 4286 4781 4301 4805
rect 4325 4781 4336 4805
rect 4286 4752 4336 4781
rect 4499 4800 4549 4829
rect 4499 4780 4516 4800
rect 4536 4780 4549 4800
rect 4499 4752 4549 4780
rect 383 4680 433 4708
rect 383 4660 396 4680
rect 416 4660 433 4680
rect 383 4631 433 4660
rect 596 4679 646 4708
rect 596 4655 607 4679
rect 631 4655 646 4679
rect 596 4631 646 4655
rect 804 4684 854 4708
rect 804 4660 816 4684
rect 840 4660 854 4684
rect 804 4631 854 4660
rect 1012 4682 1062 4708
rect 1012 4656 1030 4682
rect 1056 4656 1062 4682
rect 1012 4631 1062 4656
rect 3870 4639 3920 4652
rect 4078 4639 4128 4652
rect 4286 4639 4336 4652
rect 4499 4639 4549 4652
rect 383 4573 433 4589
rect 596 4573 646 4589
rect 804 4573 854 4589
rect 1012 4573 1062 4589
rect 2823 4585 2873 4601
rect 3031 4585 3081 4601
rect 3239 4585 3289 4601
rect 3452 4585 3502 4601
rect 1431 4545 1481 4558
rect 1644 4545 1694 4558
rect 1852 4545 1902 4558
rect 2060 4545 2110 4558
rect 2823 4518 2873 4543
rect 2823 4492 2829 4518
rect 2855 4492 2873 4518
rect 2823 4466 2873 4492
rect 3031 4514 3081 4543
rect 3031 4490 3045 4514
rect 3069 4490 3081 4514
rect 3031 4466 3081 4490
rect 3239 4519 3289 4543
rect 3239 4495 3254 4519
rect 3278 4495 3289 4519
rect 3239 4466 3289 4495
rect 3452 4514 3502 4543
rect 3452 4494 3469 4514
rect 3489 4494 3502 4514
rect 3452 4466 3502 4494
rect 1431 4417 1481 4445
rect 1431 4397 1444 4417
rect 1464 4397 1481 4417
rect 1431 4368 1481 4397
rect 1644 4416 1694 4445
rect 1644 4392 1655 4416
rect 1679 4392 1694 4416
rect 1644 4368 1694 4392
rect 1852 4421 1902 4445
rect 1852 4397 1864 4421
rect 1888 4397 1902 4421
rect 1852 4368 1902 4397
rect 2060 4419 2110 4445
rect 2060 4393 2078 4419
rect 2104 4393 2110 4419
rect 2060 4368 2110 4393
rect 2823 4353 2873 4366
rect 3031 4353 3081 4366
rect 3239 4353 3289 4366
rect 3452 4353 3502 4366
rect 1431 4310 1481 4326
rect 1644 4310 1694 4326
rect 1852 4310 1902 4326
rect 2060 4310 2110 4326
rect 3871 4322 3921 4338
rect 4079 4322 4129 4338
rect 4287 4322 4337 4338
rect 4500 4322 4550 4338
rect 384 4259 434 4272
rect 597 4259 647 4272
rect 805 4259 855 4272
rect 1013 4259 1063 4272
rect 3871 4255 3921 4280
rect 3871 4229 3877 4255
rect 3903 4229 3921 4255
rect 3871 4203 3921 4229
rect 4079 4251 4129 4280
rect 4079 4227 4093 4251
rect 4117 4227 4129 4251
rect 4079 4203 4129 4227
rect 4287 4256 4337 4280
rect 4287 4232 4302 4256
rect 4326 4232 4337 4256
rect 4287 4203 4337 4232
rect 4500 4251 4550 4280
rect 4500 4231 4517 4251
rect 4537 4231 4550 4251
rect 4500 4203 4550 4231
rect 384 4131 434 4159
rect 384 4111 397 4131
rect 417 4111 434 4131
rect 384 4082 434 4111
rect 597 4130 647 4159
rect 597 4106 608 4130
rect 632 4106 647 4130
rect 597 4082 647 4106
rect 805 4135 855 4159
rect 805 4111 817 4135
rect 841 4111 855 4135
rect 805 4082 855 4111
rect 1013 4133 1063 4159
rect 1013 4107 1031 4133
rect 1057 4107 1063 4133
rect 1013 4082 1063 4107
rect 3871 4090 3921 4103
rect 4079 4090 4129 4103
rect 4287 4090 4337 4103
rect 4500 4090 4550 4103
rect 384 4024 434 4040
rect 597 4024 647 4040
rect 805 4024 855 4040
rect 1013 4024 1063 4040
rect 1322 4015 1372 4028
rect 1535 4015 1585 4028
rect 1743 4015 1793 4028
rect 1951 4015 2001 4028
rect 2932 4012 2982 4028
rect 3140 4012 3190 4028
rect 3348 4012 3398 4028
rect 3561 4012 3611 4028
rect 2932 3945 2982 3970
rect 2932 3919 2938 3945
rect 2964 3919 2982 3945
rect 1322 3887 1372 3915
rect 1322 3867 1335 3887
rect 1355 3867 1372 3887
rect 1322 3838 1372 3867
rect 1535 3886 1585 3915
rect 1535 3862 1546 3886
rect 1570 3862 1585 3886
rect 1535 3838 1585 3862
rect 1743 3891 1793 3915
rect 1743 3867 1755 3891
rect 1779 3867 1793 3891
rect 1743 3838 1793 3867
rect 1951 3889 2001 3915
rect 2932 3893 2982 3919
rect 3140 3941 3190 3970
rect 3140 3917 3154 3941
rect 3178 3917 3190 3941
rect 3140 3893 3190 3917
rect 3348 3946 3398 3970
rect 3348 3922 3363 3946
rect 3387 3922 3398 3946
rect 3348 3893 3398 3922
rect 3561 3941 3611 3970
rect 3561 3921 3578 3941
rect 3598 3921 3611 3941
rect 3561 3893 3611 3921
rect 1951 3863 1969 3889
rect 1995 3863 2001 3889
rect 1951 3838 2001 3863
rect 1322 3780 1372 3796
rect 1535 3780 1585 3796
rect 1743 3780 1793 3796
rect 1951 3780 2001 3796
rect 2932 3780 2982 3793
rect 3140 3780 3190 3793
rect 3348 3780 3398 3793
rect 3561 3780 3611 3793
rect 3870 3768 3920 3784
rect 4078 3768 4128 3784
rect 4286 3768 4336 3784
rect 4499 3768 4549 3784
rect 383 3705 433 3718
rect 596 3705 646 3718
rect 804 3705 854 3718
rect 1012 3705 1062 3718
rect 3870 3701 3920 3726
rect 3870 3675 3876 3701
rect 3902 3675 3920 3701
rect 3870 3649 3920 3675
rect 4078 3697 4128 3726
rect 4078 3673 4092 3697
rect 4116 3673 4128 3697
rect 4078 3649 4128 3673
rect 4286 3702 4336 3726
rect 4286 3678 4301 3702
rect 4325 3678 4336 3702
rect 4286 3649 4336 3678
rect 4499 3697 4549 3726
rect 4499 3677 4516 3697
rect 4536 3677 4549 3697
rect 4499 3649 4549 3677
rect 383 3577 433 3605
rect 383 3557 396 3577
rect 416 3557 433 3577
rect 383 3528 433 3557
rect 596 3576 646 3605
rect 596 3552 607 3576
rect 631 3552 646 3576
rect 596 3528 646 3552
rect 804 3581 854 3605
rect 804 3557 816 3581
rect 840 3557 854 3581
rect 804 3528 854 3557
rect 1012 3579 1062 3605
rect 1012 3553 1030 3579
rect 1056 3553 1062 3579
rect 1012 3528 1062 3553
rect 3870 3536 3920 3549
rect 4078 3536 4128 3549
rect 4286 3536 4336 3549
rect 4499 3536 4549 3549
rect 2792 3501 2842 3517
rect 3000 3501 3050 3517
rect 3208 3501 3258 3517
rect 3421 3501 3471 3517
rect 383 3470 433 3486
rect 596 3470 646 3486
rect 804 3470 854 3486
rect 1012 3470 1062 3486
rect 1463 3423 1513 3436
rect 1676 3423 1726 3436
rect 1884 3423 1934 3436
rect 2092 3423 2142 3436
rect 2792 3434 2842 3459
rect 2792 3408 2798 3434
rect 2824 3408 2842 3434
rect 2792 3382 2842 3408
rect 3000 3430 3050 3459
rect 3000 3406 3014 3430
rect 3038 3406 3050 3430
rect 3000 3382 3050 3406
rect 3208 3435 3258 3459
rect 3208 3411 3223 3435
rect 3247 3411 3258 3435
rect 3208 3382 3258 3411
rect 3421 3430 3471 3459
rect 3421 3410 3438 3430
rect 3458 3410 3471 3430
rect 3421 3382 3471 3410
rect 1463 3295 1513 3323
rect 1463 3275 1476 3295
rect 1496 3275 1513 3295
rect 1463 3246 1513 3275
rect 1676 3294 1726 3323
rect 1676 3270 1687 3294
rect 1711 3270 1726 3294
rect 1676 3246 1726 3270
rect 1884 3299 1934 3323
rect 1884 3275 1896 3299
rect 1920 3275 1934 3299
rect 1884 3246 1934 3275
rect 2092 3297 2142 3323
rect 2092 3271 2110 3297
rect 2136 3271 2142 3297
rect 2092 3246 2142 3271
rect 2792 3269 2842 3282
rect 3000 3269 3050 3282
rect 3208 3269 3258 3282
rect 3421 3269 3471 3282
rect 3872 3219 3922 3235
rect 4080 3219 4130 3235
rect 4288 3219 4338 3235
rect 4501 3219 4551 3235
rect 1463 3188 1513 3204
rect 1676 3188 1726 3204
rect 1884 3188 1934 3204
rect 2092 3188 2142 3204
rect 385 3156 435 3169
rect 598 3156 648 3169
rect 806 3156 856 3169
rect 1014 3156 1064 3169
rect 3872 3152 3922 3177
rect 3872 3126 3878 3152
rect 3904 3126 3922 3152
rect 3872 3100 3922 3126
rect 4080 3148 4130 3177
rect 4080 3124 4094 3148
rect 4118 3124 4130 3148
rect 4080 3100 4130 3124
rect 4288 3153 4338 3177
rect 4288 3129 4303 3153
rect 4327 3129 4338 3153
rect 4288 3100 4338 3129
rect 4501 3148 4551 3177
rect 4501 3128 4518 3148
rect 4538 3128 4551 3148
rect 4501 3100 4551 3128
rect 385 3028 435 3056
rect 385 3008 398 3028
rect 418 3008 435 3028
rect 385 2979 435 3008
rect 598 3027 648 3056
rect 598 3003 609 3027
rect 633 3003 648 3027
rect 598 2979 648 3003
rect 806 3032 856 3056
rect 806 3008 818 3032
rect 842 3008 856 3032
rect 806 2979 856 3008
rect 1014 3030 1064 3056
rect 1014 3004 1032 3030
rect 1058 3004 1064 3030
rect 1014 2979 1064 3004
rect 3872 2987 3922 3000
rect 4080 2987 4130 3000
rect 4288 2987 4338 3000
rect 4501 2987 4551 3000
rect 385 2921 435 2937
rect 598 2921 648 2937
rect 806 2921 856 2937
rect 1014 2921 1064 2937
rect 1323 2912 1373 2925
rect 1536 2912 1586 2925
rect 1744 2912 1794 2925
rect 1952 2912 2002 2925
rect 2933 2909 2983 2925
rect 3141 2909 3191 2925
rect 3349 2909 3399 2925
rect 3562 2909 3612 2925
rect 2933 2842 2983 2867
rect 2933 2816 2939 2842
rect 2965 2816 2983 2842
rect 1323 2784 1373 2812
rect 1323 2764 1336 2784
rect 1356 2764 1373 2784
rect 1323 2735 1373 2764
rect 1536 2783 1586 2812
rect 1536 2759 1547 2783
rect 1571 2759 1586 2783
rect 1536 2735 1586 2759
rect 1744 2788 1794 2812
rect 1744 2764 1756 2788
rect 1780 2764 1794 2788
rect 1744 2735 1794 2764
rect 1952 2786 2002 2812
rect 2933 2790 2983 2816
rect 3141 2838 3191 2867
rect 3141 2814 3155 2838
rect 3179 2814 3191 2838
rect 3141 2790 3191 2814
rect 3349 2843 3399 2867
rect 3349 2819 3364 2843
rect 3388 2819 3399 2843
rect 3349 2790 3399 2819
rect 3562 2838 3612 2867
rect 3562 2818 3579 2838
rect 3599 2818 3612 2838
rect 3562 2790 3612 2818
rect 1952 2760 1970 2786
rect 1996 2760 2002 2786
rect 1952 2735 2002 2760
rect 1323 2677 1373 2693
rect 1536 2677 1586 2693
rect 1744 2677 1794 2693
rect 1952 2677 2002 2693
rect 2933 2677 2983 2690
rect 3141 2677 3191 2690
rect 3349 2677 3399 2690
rect 3562 2677 3612 2690
rect 3871 2665 3921 2681
rect 4079 2665 4129 2681
rect 4287 2665 4337 2681
rect 4500 2665 4550 2681
rect 384 2602 434 2615
rect 597 2602 647 2615
rect 805 2602 855 2615
rect 1013 2602 1063 2615
rect 3871 2598 3921 2623
rect 3871 2572 3877 2598
rect 3903 2572 3921 2598
rect 3871 2546 3921 2572
rect 4079 2594 4129 2623
rect 4079 2570 4093 2594
rect 4117 2570 4129 2594
rect 4079 2546 4129 2570
rect 4287 2599 4337 2623
rect 4287 2575 4302 2599
rect 4326 2575 4337 2599
rect 4287 2546 4337 2575
rect 4500 2594 4550 2623
rect 4500 2574 4517 2594
rect 4537 2574 4550 2594
rect 4500 2546 4550 2574
rect 384 2474 434 2502
rect 384 2454 397 2474
rect 417 2454 434 2474
rect 384 2425 434 2454
rect 597 2473 647 2502
rect 597 2449 608 2473
rect 632 2449 647 2473
rect 597 2425 647 2449
rect 805 2478 855 2502
rect 805 2454 817 2478
rect 841 2454 855 2478
rect 805 2425 855 2454
rect 1013 2476 1063 2502
rect 1013 2450 1031 2476
rect 1057 2450 1063 2476
rect 1013 2425 1063 2450
rect 3871 2433 3921 2446
rect 4079 2433 4129 2446
rect 4287 2433 4337 2446
rect 4500 2433 4550 2446
rect 384 2367 434 2383
rect 597 2367 647 2383
rect 805 2367 855 2383
rect 1013 2367 1063 2383
rect 2823 2385 2873 2401
rect 3031 2385 3081 2401
rect 3239 2385 3289 2401
rect 3452 2385 3502 2401
rect 1433 2333 1483 2346
rect 1646 2333 1696 2346
rect 1854 2333 1904 2346
rect 2062 2333 2112 2346
rect 2823 2318 2873 2343
rect 2823 2292 2829 2318
rect 2855 2292 2873 2318
rect 2823 2266 2873 2292
rect 3031 2314 3081 2343
rect 3031 2290 3045 2314
rect 3069 2290 3081 2314
rect 3031 2266 3081 2290
rect 3239 2319 3289 2343
rect 3239 2295 3254 2319
rect 3278 2295 3289 2319
rect 3239 2266 3289 2295
rect 3452 2314 3502 2343
rect 3452 2294 3469 2314
rect 3489 2294 3502 2314
rect 3452 2266 3502 2294
rect 1433 2205 1483 2233
rect 1433 2185 1446 2205
rect 1466 2185 1483 2205
rect 1433 2156 1483 2185
rect 1646 2204 1696 2233
rect 1646 2180 1657 2204
rect 1681 2180 1696 2204
rect 1646 2156 1696 2180
rect 1854 2209 1904 2233
rect 1854 2185 1866 2209
rect 1890 2185 1904 2209
rect 1854 2156 1904 2185
rect 2062 2207 2112 2233
rect 2062 2181 2080 2207
rect 2106 2181 2112 2207
rect 2062 2156 2112 2181
rect 2823 2153 2873 2166
rect 3031 2153 3081 2166
rect 3239 2153 3289 2166
rect 3452 2153 3502 2166
rect 1433 2098 1483 2114
rect 1646 2098 1696 2114
rect 1854 2098 1904 2114
rect 2062 2098 2112 2114
rect 3872 2116 3922 2132
rect 4080 2116 4130 2132
rect 4288 2116 4338 2132
rect 4501 2116 4551 2132
rect 385 2053 435 2066
rect 598 2053 648 2066
rect 806 2053 856 2066
rect 1014 2053 1064 2066
rect 3872 2049 3922 2074
rect 3872 2023 3878 2049
rect 3904 2023 3922 2049
rect 3872 1997 3922 2023
rect 4080 2045 4130 2074
rect 4080 2021 4094 2045
rect 4118 2021 4130 2045
rect 4080 1997 4130 2021
rect 4288 2050 4338 2074
rect 4288 2026 4303 2050
rect 4327 2026 4338 2050
rect 4288 1997 4338 2026
rect 4501 2045 4551 2074
rect 4501 2025 4518 2045
rect 4538 2025 4551 2045
rect 4501 1997 4551 2025
rect 385 1925 435 1953
rect 385 1905 398 1925
rect 418 1905 435 1925
rect 385 1876 435 1905
rect 598 1924 648 1953
rect 598 1900 609 1924
rect 633 1900 648 1924
rect 598 1876 648 1900
rect 806 1929 856 1953
rect 806 1905 818 1929
rect 842 1905 856 1929
rect 806 1876 856 1905
rect 1014 1927 1064 1953
rect 1014 1901 1032 1927
rect 1058 1901 1064 1927
rect 1014 1876 1064 1901
rect 3872 1884 3922 1897
rect 4080 1884 4130 1897
rect 4288 1884 4338 1897
rect 4501 1884 4551 1897
rect 385 1818 435 1834
rect 598 1818 648 1834
rect 806 1818 856 1834
rect 1014 1818 1064 1834
rect 1323 1809 1373 1822
rect 1536 1809 1586 1822
rect 1744 1809 1794 1822
rect 1952 1809 2002 1822
rect 2933 1806 2983 1822
rect 3141 1806 3191 1822
rect 3349 1806 3399 1822
rect 3562 1806 3612 1822
rect 2933 1739 2983 1764
rect 2933 1713 2939 1739
rect 2965 1713 2983 1739
rect 1323 1681 1373 1709
rect 1323 1661 1336 1681
rect 1356 1661 1373 1681
rect 1323 1632 1373 1661
rect 1536 1680 1586 1709
rect 1536 1656 1547 1680
rect 1571 1656 1586 1680
rect 1536 1632 1586 1656
rect 1744 1685 1794 1709
rect 1744 1661 1756 1685
rect 1780 1661 1794 1685
rect 1744 1632 1794 1661
rect 1952 1683 2002 1709
rect 2933 1687 2983 1713
rect 3141 1735 3191 1764
rect 3141 1711 3155 1735
rect 3179 1711 3191 1735
rect 3141 1687 3191 1711
rect 3349 1740 3399 1764
rect 3349 1716 3364 1740
rect 3388 1716 3399 1740
rect 3349 1687 3399 1716
rect 3562 1735 3612 1764
rect 3562 1715 3579 1735
rect 3599 1715 3612 1735
rect 3562 1687 3612 1715
rect 1952 1657 1970 1683
rect 1996 1657 2002 1683
rect 1952 1632 2002 1657
rect 1323 1574 1373 1590
rect 1536 1574 1586 1590
rect 1744 1574 1794 1590
rect 1952 1574 2002 1590
rect 2933 1574 2983 1587
rect 3141 1574 3191 1587
rect 3349 1574 3399 1587
rect 3562 1574 3612 1587
rect 3871 1562 3921 1578
rect 4079 1562 4129 1578
rect 4287 1562 4337 1578
rect 4500 1562 4550 1578
rect 384 1499 434 1512
rect 597 1499 647 1512
rect 805 1499 855 1512
rect 1013 1499 1063 1512
rect 3871 1495 3921 1520
rect 3871 1469 3877 1495
rect 3903 1469 3921 1495
rect 3871 1443 3921 1469
rect 4079 1491 4129 1520
rect 4079 1467 4093 1491
rect 4117 1467 4129 1491
rect 4079 1443 4129 1467
rect 4287 1496 4337 1520
rect 4287 1472 4302 1496
rect 4326 1472 4337 1496
rect 4287 1443 4337 1472
rect 4500 1491 4550 1520
rect 4500 1471 4517 1491
rect 4537 1471 4550 1491
rect 4500 1443 4550 1471
rect 384 1371 434 1399
rect 384 1351 397 1371
rect 417 1351 434 1371
rect 384 1322 434 1351
rect 597 1370 647 1399
rect 597 1346 608 1370
rect 632 1346 647 1370
rect 597 1322 647 1346
rect 805 1375 855 1399
rect 805 1351 817 1375
rect 841 1351 855 1375
rect 805 1322 855 1351
rect 1013 1373 1063 1399
rect 1013 1347 1031 1373
rect 1057 1347 1063 1373
rect 1013 1322 1063 1347
rect 3871 1330 3921 1343
rect 4079 1330 4129 1343
rect 4287 1330 4337 1343
rect 4500 1330 4550 1343
rect 2793 1295 2843 1311
rect 3001 1295 3051 1311
rect 3209 1295 3259 1311
rect 3422 1295 3472 1311
rect 384 1264 434 1280
rect 597 1264 647 1280
rect 805 1264 855 1280
rect 1013 1264 1063 1280
rect 1464 1217 1514 1230
rect 1677 1217 1727 1230
rect 1885 1217 1935 1230
rect 2093 1217 2143 1230
rect 2793 1228 2843 1253
rect 2793 1202 2799 1228
rect 2825 1202 2843 1228
rect 2793 1176 2843 1202
rect 3001 1224 3051 1253
rect 3001 1200 3015 1224
rect 3039 1200 3051 1224
rect 3001 1176 3051 1200
rect 3209 1229 3259 1253
rect 3209 1205 3224 1229
rect 3248 1205 3259 1229
rect 3209 1176 3259 1205
rect 3422 1224 3472 1253
rect 3422 1204 3439 1224
rect 3459 1204 3472 1224
rect 3422 1176 3472 1204
rect 1464 1089 1514 1117
rect 1464 1069 1477 1089
rect 1497 1069 1514 1089
rect 1464 1040 1514 1069
rect 1677 1088 1727 1117
rect 1677 1064 1688 1088
rect 1712 1064 1727 1088
rect 1677 1040 1727 1064
rect 1885 1093 1935 1117
rect 1885 1069 1897 1093
rect 1921 1069 1935 1093
rect 1885 1040 1935 1069
rect 2093 1091 2143 1117
rect 2093 1065 2111 1091
rect 2137 1065 2143 1091
rect 2093 1040 2143 1065
rect 2793 1063 2843 1076
rect 3001 1063 3051 1076
rect 3209 1063 3259 1076
rect 3422 1063 3472 1076
rect 3873 1013 3923 1029
rect 4081 1013 4131 1029
rect 4289 1013 4339 1029
rect 4502 1013 4552 1029
rect 1464 982 1514 998
rect 1677 982 1727 998
rect 1885 982 1935 998
rect 2093 982 2143 998
rect 386 950 436 963
rect 599 950 649 963
rect 807 950 857 963
rect 1015 950 1065 963
rect 3873 946 3923 971
rect 3873 920 3879 946
rect 3905 920 3923 946
rect 3873 894 3923 920
rect 4081 942 4131 971
rect 4081 918 4095 942
rect 4119 918 4131 942
rect 4081 894 4131 918
rect 4289 947 4339 971
rect 4289 923 4304 947
rect 4328 923 4339 947
rect 4289 894 4339 923
rect 4502 942 4552 971
rect 4502 922 4519 942
rect 4539 922 4552 942
rect 4502 894 4552 922
rect 386 822 436 850
rect 386 802 399 822
rect 419 802 436 822
rect 386 773 436 802
rect 599 821 649 850
rect 599 797 610 821
rect 634 797 649 821
rect 599 773 649 797
rect 807 826 857 850
rect 807 802 819 826
rect 843 802 857 826
rect 807 773 857 802
rect 1015 824 1065 850
rect 1015 798 1033 824
rect 1059 798 1065 824
rect 1015 773 1065 798
rect 3873 781 3923 794
rect 4081 781 4131 794
rect 4289 781 4339 794
rect 4502 781 4552 794
rect 386 715 436 731
rect 599 715 649 731
rect 807 715 857 731
rect 1015 715 1065 731
rect 1324 706 1374 719
rect 1537 706 1587 719
rect 1745 706 1795 719
rect 1953 706 2003 719
rect 2934 703 2984 719
rect 3142 703 3192 719
rect 3350 703 3400 719
rect 3563 703 3613 719
rect 2934 636 2984 661
rect 2934 610 2940 636
rect 2966 610 2984 636
rect 1324 578 1374 606
rect 1324 558 1337 578
rect 1357 558 1374 578
rect 1324 529 1374 558
rect 1537 577 1587 606
rect 1537 553 1548 577
rect 1572 553 1587 577
rect 1537 529 1587 553
rect 1745 582 1795 606
rect 1745 558 1757 582
rect 1781 558 1795 582
rect 1745 529 1795 558
rect 1953 580 2003 606
rect 2934 584 2984 610
rect 3142 632 3192 661
rect 3142 608 3156 632
rect 3180 608 3192 632
rect 3142 584 3192 608
rect 3350 637 3400 661
rect 3350 613 3365 637
rect 3389 613 3400 637
rect 3350 584 3400 613
rect 3563 632 3613 661
rect 3563 612 3580 632
rect 3600 612 3613 632
rect 3563 584 3613 612
rect 1953 554 1971 580
rect 1997 554 2003 580
rect 1953 529 2003 554
rect 1324 471 1374 487
rect 1537 471 1587 487
rect 1745 471 1795 487
rect 1953 471 2003 487
rect 2934 471 2984 484
rect 3142 471 3192 484
rect 3350 471 3400 484
rect 3563 471 3613 484
rect 3872 459 3922 475
rect 4080 459 4130 475
rect 4288 459 4338 475
rect 4501 459 4551 475
rect 385 396 435 409
rect 598 396 648 409
rect 806 396 856 409
rect 1014 396 1064 409
rect 3872 392 3922 417
rect 3872 366 3878 392
rect 3904 366 3922 392
rect 3872 340 3922 366
rect 4080 388 4130 417
rect 4080 364 4094 388
rect 4118 364 4130 388
rect 4080 340 4130 364
rect 4288 393 4338 417
rect 4288 369 4303 393
rect 4327 369 4338 393
rect 4288 340 4338 369
rect 4501 388 4551 417
rect 4501 368 4518 388
rect 4538 368 4551 388
rect 4501 340 4551 368
rect 385 268 435 296
rect 385 248 398 268
rect 418 248 435 268
rect 385 219 435 248
rect 598 267 648 296
rect 598 243 609 267
rect 633 243 648 267
rect 598 219 648 243
rect 806 272 856 296
rect 806 248 818 272
rect 842 248 856 272
rect 806 219 856 248
rect 1014 270 1064 296
rect 1014 244 1032 270
rect 1058 244 1064 270
rect 1014 219 1064 244
rect 3872 227 3922 240
rect 4080 227 4130 240
rect 4288 227 4338 240
rect 4501 227 4551 240
rect 385 161 435 177
rect 598 161 648 177
rect 806 161 856 177
rect 1014 161 1064 177
rect 1632 -163 1682 -150
rect 1845 -163 1895 -150
rect 2053 -163 2103 -150
rect 2261 -163 2311 -150
rect 1632 -291 1682 -263
rect 1632 -311 1645 -291
rect 1665 -311 1682 -291
rect 1632 -340 1682 -311
rect 1845 -292 1895 -263
rect 1845 -316 1856 -292
rect 1880 -316 1895 -292
rect 1845 -340 1895 -316
rect 2053 -287 2103 -263
rect 2053 -311 2065 -287
rect 2089 -311 2103 -287
rect 2053 -340 2103 -311
rect 2261 -289 2311 -263
rect 2261 -315 2279 -289
rect 2305 -315 2311 -289
rect 2261 -340 2311 -315
rect 1632 -398 1682 -382
rect 1845 -398 1895 -382
rect 2053 -398 2103 -382
rect 2261 -398 2311 -382
<< polycont >>
rect 3875 8641 3901 8667
rect 4091 8639 4115 8663
rect 4300 8644 4324 8668
rect 4515 8643 4535 8663
rect 395 8523 415 8543
rect 606 8518 630 8542
rect 815 8523 839 8547
rect 1029 8519 1055 8545
rect 2936 8331 2962 8357
rect 1333 8279 1353 8299
rect 1544 8274 1568 8298
rect 1753 8279 1777 8303
rect 3152 8329 3176 8353
rect 3361 8334 3385 8358
rect 3576 8333 3596 8353
rect 1967 8275 1993 8301
rect 3874 8087 3900 8113
rect 4090 8085 4114 8109
rect 4299 8090 4323 8114
rect 4514 8089 4534 8109
rect 394 7969 414 7989
rect 605 7964 629 7988
rect 814 7969 838 7993
rect 1028 7965 1054 7991
rect 2796 7820 2822 7846
rect 3012 7818 3036 7842
rect 3221 7823 3245 7847
rect 3436 7822 3456 7842
rect 1474 7687 1494 7707
rect 1685 7682 1709 7706
rect 1894 7687 1918 7711
rect 2108 7683 2134 7709
rect 3876 7538 3902 7564
rect 4092 7536 4116 7560
rect 4301 7541 4325 7565
rect 4516 7540 4536 7560
rect 396 7420 416 7440
rect 607 7415 631 7439
rect 816 7420 840 7444
rect 1030 7416 1056 7442
rect 2937 7228 2963 7254
rect 1334 7176 1354 7196
rect 1545 7171 1569 7195
rect 1754 7176 1778 7200
rect 3153 7226 3177 7250
rect 3362 7231 3386 7255
rect 3577 7230 3597 7250
rect 1968 7172 1994 7198
rect 3875 6984 3901 7010
rect 4091 6982 4115 7006
rect 4300 6987 4324 7011
rect 4515 6986 4535 7006
rect 395 6866 415 6886
rect 606 6861 630 6885
rect 815 6866 839 6890
rect 1029 6862 1055 6888
rect 2827 6704 2853 6730
rect 3043 6702 3067 6726
rect 3252 6707 3276 6731
rect 3467 6706 3487 6726
rect 1444 6597 1464 6617
rect 1655 6592 1679 6616
rect 1864 6597 1888 6621
rect 2078 6593 2104 6619
rect 3876 6435 3902 6461
rect 4092 6433 4116 6457
rect 4301 6438 4325 6462
rect 4516 6437 4536 6457
rect 396 6317 416 6337
rect 607 6312 631 6336
rect 816 6317 840 6341
rect 1030 6313 1056 6339
rect 2937 6125 2963 6151
rect 1334 6073 1354 6093
rect 1545 6068 1569 6092
rect 1754 6073 1778 6097
rect 3153 6123 3177 6147
rect 3362 6128 3386 6152
rect 3577 6127 3597 6147
rect 1968 6069 1994 6095
rect 3875 5881 3901 5907
rect 4091 5879 4115 5903
rect 4300 5884 4324 5908
rect 4515 5883 4535 5903
rect 395 5763 415 5783
rect 606 5758 630 5782
rect 815 5763 839 5787
rect 1029 5759 1055 5785
rect 2797 5614 2823 5640
rect 3013 5612 3037 5636
rect 3222 5617 3246 5641
rect 3437 5616 3457 5636
rect 1475 5481 1495 5501
rect 1686 5476 1710 5500
rect 1895 5481 1919 5505
rect 2109 5477 2135 5503
rect 3877 5332 3903 5358
rect 4093 5330 4117 5354
rect 4302 5335 4326 5359
rect 4517 5334 4537 5354
rect 397 5214 417 5234
rect 608 5209 632 5233
rect 817 5214 841 5238
rect 1031 5210 1057 5236
rect 2938 5022 2964 5048
rect 1335 4970 1355 4990
rect 1546 4965 1570 4989
rect 1755 4970 1779 4994
rect 3154 5020 3178 5044
rect 3363 5025 3387 5049
rect 3578 5024 3598 5044
rect 1969 4966 1995 4992
rect 3876 4778 3902 4804
rect 4092 4776 4116 4800
rect 4301 4781 4325 4805
rect 4516 4780 4536 4800
rect 396 4660 416 4680
rect 607 4655 631 4679
rect 816 4660 840 4684
rect 1030 4656 1056 4682
rect 2829 4492 2855 4518
rect 3045 4490 3069 4514
rect 3254 4495 3278 4519
rect 3469 4494 3489 4514
rect 1444 4397 1464 4417
rect 1655 4392 1679 4416
rect 1864 4397 1888 4421
rect 2078 4393 2104 4419
rect 3877 4229 3903 4255
rect 4093 4227 4117 4251
rect 4302 4232 4326 4256
rect 4517 4231 4537 4251
rect 397 4111 417 4131
rect 608 4106 632 4130
rect 817 4111 841 4135
rect 1031 4107 1057 4133
rect 2938 3919 2964 3945
rect 1335 3867 1355 3887
rect 1546 3862 1570 3886
rect 1755 3867 1779 3891
rect 3154 3917 3178 3941
rect 3363 3922 3387 3946
rect 3578 3921 3598 3941
rect 1969 3863 1995 3889
rect 3876 3675 3902 3701
rect 4092 3673 4116 3697
rect 4301 3678 4325 3702
rect 4516 3677 4536 3697
rect 396 3557 416 3577
rect 607 3552 631 3576
rect 816 3557 840 3581
rect 1030 3553 1056 3579
rect 2798 3408 2824 3434
rect 3014 3406 3038 3430
rect 3223 3411 3247 3435
rect 3438 3410 3458 3430
rect 1476 3275 1496 3295
rect 1687 3270 1711 3294
rect 1896 3275 1920 3299
rect 2110 3271 2136 3297
rect 3878 3126 3904 3152
rect 4094 3124 4118 3148
rect 4303 3129 4327 3153
rect 4518 3128 4538 3148
rect 398 3008 418 3028
rect 609 3003 633 3027
rect 818 3008 842 3032
rect 1032 3004 1058 3030
rect 2939 2816 2965 2842
rect 1336 2764 1356 2784
rect 1547 2759 1571 2783
rect 1756 2764 1780 2788
rect 3155 2814 3179 2838
rect 3364 2819 3388 2843
rect 3579 2818 3599 2838
rect 1970 2760 1996 2786
rect 3877 2572 3903 2598
rect 4093 2570 4117 2594
rect 4302 2575 4326 2599
rect 4517 2574 4537 2594
rect 397 2454 417 2474
rect 608 2449 632 2473
rect 817 2454 841 2478
rect 1031 2450 1057 2476
rect 2829 2292 2855 2318
rect 3045 2290 3069 2314
rect 3254 2295 3278 2319
rect 3469 2294 3489 2314
rect 1446 2185 1466 2205
rect 1657 2180 1681 2204
rect 1866 2185 1890 2209
rect 2080 2181 2106 2207
rect 3878 2023 3904 2049
rect 4094 2021 4118 2045
rect 4303 2026 4327 2050
rect 4518 2025 4538 2045
rect 398 1905 418 1925
rect 609 1900 633 1924
rect 818 1905 842 1929
rect 1032 1901 1058 1927
rect 2939 1713 2965 1739
rect 1336 1661 1356 1681
rect 1547 1656 1571 1680
rect 1756 1661 1780 1685
rect 3155 1711 3179 1735
rect 3364 1716 3388 1740
rect 3579 1715 3599 1735
rect 1970 1657 1996 1683
rect 3877 1469 3903 1495
rect 4093 1467 4117 1491
rect 4302 1472 4326 1496
rect 4517 1471 4537 1491
rect 397 1351 417 1371
rect 608 1346 632 1370
rect 817 1351 841 1375
rect 1031 1347 1057 1373
rect 2799 1202 2825 1228
rect 3015 1200 3039 1224
rect 3224 1205 3248 1229
rect 3439 1204 3459 1224
rect 1477 1069 1497 1089
rect 1688 1064 1712 1088
rect 1897 1069 1921 1093
rect 2111 1065 2137 1091
rect 3879 920 3905 946
rect 4095 918 4119 942
rect 4304 923 4328 947
rect 4519 922 4539 942
rect 399 802 419 822
rect 610 797 634 821
rect 819 802 843 826
rect 1033 798 1059 824
rect 2940 610 2966 636
rect 1337 558 1357 578
rect 1548 553 1572 577
rect 1757 558 1781 582
rect 3156 608 3180 632
rect 3365 613 3389 637
rect 3580 612 3600 632
rect 1971 554 1997 580
rect 3878 366 3904 392
rect 4094 364 4118 388
rect 4303 369 4327 393
rect 4518 368 4538 388
rect 398 248 418 268
rect 609 243 633 267
rect 818 248 842 272
rect 1032 244 1058 270
rect 1645 -311 1665 -291
rect 1856 -316 1880 -292
rect 2065 -311 2089 -287
rect 2279 -315 2305 -289
<< ndiffres >>
rect 95 8767 152 8786
rect 95 8764 116 8767
rect 1 8749 116 8764
rect 134 8749 152 8767
rect 1 8726 152 8749
rect 1 8690 43 8726
rect 0 8689 100 8690
rect 0 8668 156 8689
rect 0 8650 118 8668
rect 136 8650 156 8668
rect 0 8646 156 8650
rect 95 8630 156 8646
rect 95 8580 152 8599
rect 95 8577 116 8580
rect 1 8562 116 8577
rect 134 8562 152 8580
rect 4773 8632 4834 8648
rect 4773 8628 4929 8632
rect 1 8539 152 8562
rect 1 8503 43 8539
rect 0 8502 100 8503
rect 0 8481 156 8502
rect 0 8463 118 8481
rect 136 8463 156 8481
rect 0 8459 156 8463
rect 95 8443 156 8459
rect 4773 8610 4793 8628
rect 4811 8610 4929 8628
rect 4773 8589 4929 8610
rect 4829 8588 4929 8589
rect 4886 8552 4928 8588
rect 4777 8529 4928 8552
rect 4777 8511 4795 8529
rect 4813 8514 4928 8529
rect 4813 8511 4834 8514
rect 4777 8492 4834 8511
rect 95 8351 152 8370
rect 95 8348 116 8351
rect 1 8333 116 8348
rect 134 8333 152 8351
rect 1 8310 152 8333
rect 4773 8402 4834 8418
rect 4773 8398 4929 8402
rect 1 8274 43 8310
rect 0 8273 100 8274
rect 0 8252 156 8273
rect 0 8234 118 8252
rect 136 8234 156 8252
rect 4773 8380 4793 8398
rect 4811 8380 4929 8398
rect 4773 8359 4929 8380
rect 4829 8358 4929 8359
rect 4886 8322 4928 8358
rect 0 8230 156 8234
rect 95 8214 156 8230
rect 4777 8299 4928 8322
rect 4777 8281 4795 8299
rect 4813 8284 4928 8299
rect 4813 8281 4834 8284
rect 4777 8262 4834 8281
rect 95 8121 152 8140
rect 95 8118 116 8121
rect 1 8103 116 8118
rect 134 8103 152 8121
rect 1 8080 152 8103
rect 1 8044 43 8080
rect 0 8043 100 8044
rect 0 8022 156 8043
rect 0 8004 118 8022
rect 136 8004 156 8022
rect 4773 8173 4834 8189
rect 4773 8169 4929 8173
rect 4773 8151 4793 8169
rect 4811 8151 4929 8169
rect 4773 8130 4929 8151
rect 4829 8129 4929 8130
rect 4886 8093 4928 8129
rect 4777 8070 4928 8093
rect 0 8000 156 8004
rect 95 7984 156 8000
rect 4777 8052 4795 8070
rect 4813 8055 4928 8070
rect 4813 8052 4834 8055
rect 4777 8033 4834 8052
rect 4773 7986 4834 8002
rect 4773 7982 4929 7986
rect 4773 7964 4793 7982
rect 4811 7964 4929 7982
rect 4773 7943 4929 7964
rect 4829 7942 4929 7943
rect 4886 7906 4928 7942
rect 4777 7883 4928 7906
rect 4777 7865 4795 7883
rect 4813 7868 4928 7883
rect 4813 7865 4834 7868
rect 4777 7846 4834 7865
rect 96 7664 153 7683
rect 96 7661 117 7664
rect 2 7646 117 7661
rect 135 7646 153 7664
rect 2 7623 153 7646
rect 2 7587 44 7623
rect 1 7586 101 7587
rect 1 7565 157 7586
rect 1 7547 119 7565
rect 137 7547 157 7565
rect 1 7543 157 7547
rect 96 7527 157 7543
rect 96 7477 153 7496
rect 96 7474 117 7477
rect 2 7459 117 7474
rect 135 7459 153 7477
rect 4774 7529 4835 7545
rect 4774 7525 4930 7529
rect 2 7436 153 7459
rect 2 7400 44 7436
rect 1 7399 101 7400
rect 1 7378 157 7399
rect 1 7360 119 7378
rect 137 7360 157 7378
rect 1 7356 157 7360
rect 96 7340 157 7356
rect 4774 7507 4794 7525
rect 4812 7507 4930 7525
rect 4774 7486 4930 7507
rect 4830 7485 4930 7486
rect 4887 7449 4929 7485
rect 4778 7426 4929 7449
rect 4778 7408 4796 7426
rect 4814 7411 4929 7426
rect 4814 7408 4835 7411
rect 4778 7389 4835 7408
rect 96 7248 153 7267
rect 96 7245 117 7248
rect 2 7230 117 7245
rect 135 7230 153 7248
rect 2 7207 153 7230
rect 4774 7299 4835 7315
rect 4774 7295 4930 7299
rect 2 7171 44 7207
rect 1 7170 101 7171
rect 1 7149 157 7170
rect 1 7131 119 7149
rect 137 7131 157 7149
rect 4774 7277 4794 7295
rect 4812 7277 4930 7295
rect 4774 7256 4930 7277
rect 4830 7255 4930 7256
rect 4887 7219 4929 7255
rect 1 7127 157 7131
rect 96 7111 157 7127
rect 4778 7196 4929 7219
rect 4778 7178 4796 7196
rect 4814 7181 4929 7196
rect 4814 7178 4835 7181
rect 4778 7159 4835 7178
rect 96 7018 153 7037
rect 96 7015 117 7018
rect 2 7000 117 7015
rect 135 7000 153 7018
rect 2 6977 153 7000
rect 2 6941 44 6977
rect 1 6940 101 6941
rect 1 6919 157 6940
rect 1 6901 119 6919
rect 137 6901 157 6919
rect 4774 7070 4835 7086
rect 4774 7066 4930 7070
rect 4774 7048 4794 7066
rect 4812 7048 4930 7066
rect 4774 7027 4930 7048
rect 4830 7026 4930 7027
rect 4887 6990 4929 7026
rect 4778 6967 4929 6990
rect 1 6897 157 6901
rect 96 6881 157 6897
rect 4778 6949 4796 6967
rect 4814 6952 4929 6967
rect 4814 6949 4835 6952
rect 4778 6930 4835 6949
rect 4774 6883 4835 6899
rect 4774 6879 4930 6883
rect 4774 6861 4794 6879
rect 4812 6861 4930 6879
rect 4774 6840 4930 6861
rect 4830 6839 4930 6840
rect 4887 6803 4929 6839
rect 4778 6780 4929 6803
rect 4778 6762 4796 6780
rect 4814 6765 4929 6780
rect 4814 6762 4835 6765
rect 4778 6743 4835 6762
rect 96 6561 153 6580
rect 96 6558 117 6561
rect 2 6543 117 6558
rect 135 6543 153 6561
rect 2 6520 153 6543
rect 2 6484 44 6520
rect 1 6483 101 6484
rect 1 6462 157 6483
rect 1 6444 119 6462
rect 137 6444 157 6462
rect 1 6440 157 6444
rect 96 6424 157 6440
rect 96 6374 153 6393
rect 96 6371 117 6374
rect 2 6356 117 6371
rect 135 6356 153 6374
rect 4774 6426 4835 6442
rect 4774 6422 4930 6426
rect 2 6333 153 6356
rect 2 6297 44 6333
rect 1 6296 101 6297
rect 1 6275 157 6296
rect 1 6257 119 6275
rect 137 6257 157 6275
rect 1 6253 157 6257
rect 96 6237 157 6253
rect 4774 6404 4794 6422
rect 4812 6404 4930 6422
rect 4774 6383 4930 6404
rect 4830 6382 4930 6383
rect 4887 6346 4929 6382
rect 4778 6323 4929 6346
rect 4778 6305 4796 6323
rect 4814 6308 4929 6323
rect 4814 6305 4835 6308
rect 4778 6286 4835 6305
rect 96 6145 153 6164
rect 96 6142 117 6145
rect 2 6127 117 6142
rect 135 6127 153 6145
rect 2 6104 153 6127
rect 4774 6196 4835 6212
rect 4774 6192 4930 6196
rect 2 6068 44 6104
rect 1 6067 101 6068
rect 1 6046 157 6067
rect 1 6028 119 6046
rect 137 6028 157 6046
rect 4774 6174 4794 6192
rect 4812 6174 4930 6192
rect 4774 6153 4930 6174
rect 4830 6152 4930 6153
rect 4887 6116 4929 6152
rect 1 6024 157 6028
rect 96 6008 157 6024
rect 4778 6093 4929 6116
rect 4778 6075 4796 6093
rect 4814 6078 4929 6093
rect 4814 6075 4835 6078
rect 4778 6056 4835 6075
rect 96 5915 153 5934
rect 96 5912 117 5915
rect 2 5897 117 5912
rect 135 5897 153 5915
rect 2 5874 153 5897
rect 2 5838 44 5874
rect 1 5837 101 5838
rect 1 5816 157 5837
rect 1 5798 119 5816
rect 137 5798 157 5816
rect 4774 5967 4835 5983
rect 4774 5963 4930 5967
rect 4774 5945 4794 5963
rect 4812 5945 4930 5963
rect 4774 5924 4930 5945
rect 4830 5923 4930 5924
rect 4887 5887 4929 5923
rect 4778 5864 4929 5887
rect 1 5794 157 5798
rect 96 5778 157 5794
rect 4778 5846 4796 5864
rect 4814 5849 4929 5864
rect 4814 5846 4835 5849
rect 4778 5827 4835 5846
rect 4774 5780 4835 5796
rect 4774 5776 4930 5780
rect 4774 5758 4794 5776
rect 4812 5758 4930 5776
rect 4774 5737 4930 5758
rect 4830 5736 4930 5737
rect 4887 5700 4929 5736
rect 4778 5677 4929 5700
rect 4778 5659 4796 5677
rect 4814 5662 4929 5677
rect 4814 5659 4835 5662
rect 4778 5640 4835 5659
rect 97 5458 154 5477
rect 97 5455 118 5458
rect 3 5440 118 5455
rect 136 5440 154 5458
rect 3 5417 154 5440
rect 3 5381 45 5417
rect 2 5380 102 5381
rect 2 5359 158 5380
rect 2 5341 120 5359
rect 138 5341 158 5359
rect 2 5337 158 5341
rect 97 5321 158 5337
rect 97 5271 154 5290
rect 97 5268 118 5271
rect 3 5253 118 5268
rect 136 5253 154 5271
rect 4775 5323 4836 5339
rect 4775 5319 4931 5323
rect 3 5230 154 5253
rect 3 5194 45 5230
rect 2 5193 102 5194
rect 2 5172 158 5193
rect 2 5154 120 5172
rect 138 5154 158 5172
rect 2 5150 158 5154
rect 97 5134 158 5150
rect 4775 5301 4795 5319
rect 4813 5301 4931 5319
rect 4775 5280 4931 5301
rect 4831 5279 4931 5280
rect 4888 5243 4930 5279
rect 4779 5220 4930 5243
rect 4779 5202 4797 5220
rect 4815 5205 4930 5220
rect 4815 5202 4836 5205
rect 4779 5183 4836 5202
rect 97 5042 154 5061
rect 97 5039 118 5042
rect 3 5024 118 5039
rect 136 5024 154 5042
rect 3 5001 154 5024
rect 4775 5093 4836 5109
rect 4775 5089 4931 5093
rect 3 4965 45 5001
rect 2 4964 102 4965
rect 2 4943 158 4964
rect 2 4925 120 4943
rect 138 4925 158 4943
rect 4775 5071 4795 5089
rect 4813 5071 4931 5089
rect 4775 5050 4931 5071
rect 4831 5049 4931 5050
rect 4888 5013 4930 5049
rect 2 4921 158 4925
rect 97 4905 158 4921
rect 4779 4990 4930 5013
rect 4779 4972 4797 4990
rect 4815 4975 4930 4990
rect 4815 4972 4836 4975
rect 4779 4953 4836 4972
rect 97 4812 154 4831
rect 97 4809 118 4812
rect 3 4794 118 4809
rect 136 4794 154 4812
rect 3 4771 154 4794
rect 3 4735 45 4771
rect 2 4734 102 4735
rect 2 4713 158 4734
rect 2 4695 120 4713
rect 138 4695 158 4713
rect 4775 4864 4836 4880
rect 4775 4860 4931 4864
rect 4775 4842 4795 4860
rect 4813 4842 4931 4860
rect 4775 4821 4931 4842
rect 4831 4820 4931 4821
rect 4888 4784 4930 4820
rect 4779 4761 4930 4784
rect 2 4691 158 4695
rect 97 4675 158 4691
rect 4779 4743 4797 4761
rect 4815 4746 4930 4761
rect 4815 4743 4836 4746
rect 4779 4724 4836 4743
rect 4775 4677 4836 4693
rect 4775 4673 4931 4677
rect 4775 4655 4795 4673
rect 4813 4655 4931 4673
rect 4775 4634 4931 4655
rect 4831 4633 4931 4634
rect 4888 4597 4930 4633
rect 4779 4574 4930 4597
rect 4779 4556 4797 4574
rect 4815 4559 4930 4574
rect 4815 4556 4836 4559
rect 4779 4537 4836 4556
rect 97 4355 154 4374
rect 97 4352 118 4355
rect 3 4337 118 4352
rect 136 4337 154 4355
rect 3 4314 154 4337
rect 3 4278 45 4314
rect 2 4277 102 4278
rect 2 4256 158 4277
rect 2 4238 120 4256
rect 138 4238 158 4256
rect 2 4234 158 4238
rect 97 4218 158 4234
rect 97 4168 154 4187
rect 97 4165 118 4168
rect 3 4150 118 4165
rect 136 4150 154 4168
rect 4775 4220 4836 4236
rect 4775 4216 4931 4220
rect 3 4127 154 4150
rect 3 4091 45 4127
rect 2 4090 102 4091
rect 2 4069 158 4090
rect 2 4051 120 4069
rect 138 4051 158 4069
rect 2 4047 158 4051
rect 97 4031 158 4047
rect 4775 4198 4795 4216
rect 4813 4198 4931 4216
rect 4775 4177 4931 4198
rect 4831 4176 4931 4177
rect 4888 4140 4930 4176
rect 4779 4117 4930 4140
rect 4779 4099 4797 4117
rect 4815 4102 4930 4117
rect 4815 4099 4836 4102
rect 4779 4080 4836 4099
rect 97 3939 154 3958
rect 97 3936 118 3939
rect 3 3921 118 3936
rect 136 3921 154 3939
rect 3 3898 154 3921
rect 4775 3990 4836 4006
rect 4775 3986 4931 3990
rect 3 3862 45 3898
rect 2 3861 102 3862
rect 2 3840 158 3861
rect 2 3822 120 3840
rect 138 3822 158 3840
rect 4775 3968 4795 3986
rect 4813 3968 4931 3986
rect 4775 3947 4931 3968
rect 4831 3946 4931 3947
rect 4888 3910 4930 3946
rect 2 3818 158 3822
rect 97 3802 158 3818
rect 4779 3887 4930 3910
rect 4779 3869 4797 3887
rect 4815 3872 4930 3887
rect 4815 3869 4836 3872
rect 4779 3850 4836 3869
rect 97 3709 154 3728
rect 97 3706 118 3709
rect 3 3691 118 3706
rect 136 3691 154 3709
rect 3 3668 154 3691
rect 3 3632 45 3668
rect 2 3631 102 3632
rect 2 3610 158 3631
rect 2 3592 120 3610
rect 138 3592 158 3610
rect 4775 3761 4836 3777
rect 4775 3757 4931 3761
rect 4775 3739 4795 3757
rect 4813 3739 4931 3757
rect 4775 3718 4931 3739
rect 4831 3717 4931 3718
rect 4888 3681 4930 3717
rect 4779 3658 4930 3681
rect 2 3588 158 3592
rect 97 3572 158 3588
rect 4779 3640 4797 3658
rect 4815 3643 4930 3658
rect 4815 3640 4836 3643
rect 4779 3621 4836 3640
rect 4775 3574 4836 3590
rect 4775 3570 4931 3574
rect 4775 3552 4795 3570
rect 4813 3552 4931 3570
rect 4775 3531 4931 3552
rect 4831 3530 4931 3531
rect 4888 3494 4930 3530
rect 4779 3471 4930 3494
rect 4779 3453 4797 3471
rect 4815 3456 4930 3471
rect 4815 3453 4836 3456
rect 4779 3434 4836 3453
rect 98 3252 155 3271
rect 98 3249 119 3252
rect 4 3234 119 3249
rect 137 3234 155 3252
rect 4 3211 155 3234
rect 4 3175 46 3211
rect 3 3174 103 3175
rect 3 3153 159 3174
rect 3 3135 121 3153
rect 139 3135 159 3153
rect 3 3131 159 3135
rect 98 3115 159 3131
rect 98 3065 155 3084
rect 98 3062 119 3065
rect 4 3047 119 3062
rect 137 3047 155 3065
rect 4776 3117 4837 3133
rect 4776 3113 4932 3117
rect 4 3024 155 3047
rect 4 2988 46 3024
rect 3 2987 103 2988
rect 3 2966 159 2987
rect 3 2948 121 2966
rect 139 2948 159 2966
rect 3 2944 159 2948
rect 98 2928 159 2944
rect 4776 3095 4796 3113
rect 4814 3095 4932 3113
rect 4776 3074 4932 3095
rect 4832 3073 4932 3074
rect 4889 3037 4931 3073
rect 4780 3014 4931 3037
rect 4780 2996 4798 3014
rect 4816 2999 4931 3014
rect 4816 2996 4837 2999
rect 4780 2977 4837 2996
rect 98 2836 155 2855
rect 98 2833 119 2836
rect 4 2818 119 2833
rect 137 2818 155 2836
rect 4 2795 155 2818
rect 4776 2887 4837 2903
rect 4776 2883 4932 2887
rect 4 2759 46 2795
rect 3 2758 103 2759
rect 3 2737 159 2758
rect 3 2719 121 2737
rect 139 2719 159 2737
rect 4776 2865 4796 2883
rect 4814 2865 4932 2883
rect 4776 2844 4932 2865
rect 4832 2843 4932 2844
rect 4889 2807 4931 2843
rect 3 2715 159 2719
rect 98 2699 159 2715
rect 4780 2784 4931 2807
rect 4780 2766 4798 2784
rect 4816 2769 4931 2784
rect 4816 2766 4837 2769
rect 4780 2747 4837 2766
rect 98 2606 155 2625
rect 98 2603 119 2606
rect 4 2588 119 2603
rect 137 2588 155 2606
rect 4 2565 155 2588
rect 4 2529 46 2565
rect 3 2528 103 2529
rect 3 2507 159 2528
rect 3 2489 121 2507
rect 139 2489 159 2507
rect 4776 2658 4837 2674
rect 4776 2654 4932 2658
rect 4776 2636 4796 2654
rect 4814 2636 4932 2654
rect 4776 2615 4932 2636
rect 4832 2614 4932 2615
rect 4889 2578 4931 2614
rect 4780 2555 4931 2578
rect 3 2485 159 2489
rect 98 2469 159 2485
rect 4780 2537 4798 2555
rect 4816 2540 4931 2555
rect 4816 2537 4837 2540
rect 4780 2518 4837 2537
rect 4776 2471 4837 2487
rect 4776 2467 4932 2471
rect 4776 2449 4796 2467
rect 4814 2449 4932 2467
rect 4776 2428 4932 2449
rect 4832 2427 4932 2428
rect 4889 2391 4931 2427
rect 4780 2368 4931 2391
rect 4780 2350 4798 2368
rect 4816 2353 4931 2368
rect 4816 2350 4837 2353
rect 4780 2331 4837 2350
rect 98 2149 155 2168
rect 98 2146 119 2149
rect 4 2131 119 2146
rect 137 2131 155 2149
rect 4 2108 155 2131
rect 4 2072 46 2108
rect 3 2071 103 2072
rect 3 2050 159 2071
rect 3 2032 121 2050
rect 139 2032 159 2050
rect 3 2028 159 2032
rect 98 2012 159 2028
rect 98 1962 155 1981
rect 98 1959 119 1962
rect 4 1944 119 1959
rect 137 1944 155 1962
rect 4776 2014 4837 2030
rect 4776 2010 4932 2014
rect 4 1921 155 1944
rect 4 1885 46 1921
rect 3 1884 103 1885
rect 3 1863 159 1884
rect 3 1845 121 1863
rect 139 1845 159 1863
rect 3 1841 159 1845
rect 98 1825 159 1841
rect 4776 1992 4796 2010
rect 4814 1992 4932 2010
rect 4776 1971 4932 1992
rect 4832 1970 4932 1971
rect 4889 1934 4931 1970
rect 4780 1911 4931 1934
rect 4780 1893 4798 1911
rect 4816 1896 4931 1911
rect 4816 1893 4837 1896
rect 4780 1874 4837 1893
rect 98 1733 155 1752
rect 98 1730 119 1733
rect 4 1715 119 1730
rect 137 1715 155 1733
rect 4 1692 155 1715
rect 4776 1784 4837 1800
rect 4776 1780 4932 1784
rect 4 1656 46 1692
rect 3 1655 103 1656
rect 3 1634 159 1655
rect 3 1616 121 1634
rect 139 1616 159 1634
rect 4776 1762 4796 1780
rect 4814 1762 4932 1780
rect 4776 1741 4932 1762
rect 4832 1740 4932 1741
rect 4889 1704 4931 1740
rect 3 1612 159 1616
rect 98 1596 159 1612
rect 4780 1681 4931 1704
rect 4780 1663 4798 1681
rect 4816 1666 4931 1681
rect 4816 1663 4837 1666
rect 4780 1644 4837 1663
rect 98 1503 155 1522
rect 98 1500 119 1503
rect 4 1485 119 1500
rect 137 1485 155 1503
rect 4 1462 155 1485
rect 4 1426 46 1462
rect 3 1425 103 1426
rect 3 1404 159 1425
rect 3 1386 121 1404
rect 139 1386 159 1404
rect 4776 1555 4837 1571
rect 4776 1551 4932 1555
rect 4776 1533 4796 1551
rect 4814 1533 4932 1551
rect 4776 1512 4932 1533
rect 4832 1511 4932 1512
rect 4889 1475 4931 1511
rect 4780 1452 4931 1475
rect 3 1382 159 1386
rect 98 1366 159 1382
rect 4780 1434 4798 1452
rect 4816 1437 4931 1452
rect 4816 1434 4837 1437
rect 4780 1415 4837 1434
rect 4776 1368 4837 1384
rect 4776 1364 4932 1368
rect 4776 1346 4796 1364
rect 4814 1346 4932 1364
rect 4776 1325 4932 1346
rect 4832 1324 4932 1325
rect 4889 1288 4931 1324
rect 4780 1265 4931 1288
rect 4780 1247 4798 1265
rect 4816 1250 4931 1265
rect 4816 1247 4837 1250
rect 4780 1228 4837 1247
rect 99 1046 156 1065
rect 99 1043 120 1046
rect 5 1028 120 1043
rect 138 1028 156 1046
rect 5 1005 156 1028
rect 5 969 47 1005
rect 4 968 104 969
rect 4 947 160 968
rect 4 929 122 947
rect 140 929 160 947
rect 4 925 160 929
rect 99 909 160 925
rect 99 859 156 878
rect 99 856 120 859
rect 5 841 120 856
rect 138 841 156 859
rect 4777 911 4838 927
rect 4777 907 4933 911
rect 5 818 156 841
rect 5 782 47 818
rect 4 781 104 782
rect 4 760 160 781
rect 4 742 122 760
rect 140 742 160 760
rect 4 738 160 742
rect 99 722 160 738
rect 4777 889 4797 907
rect 4815 889 4933 907
rect 4777 868 4933 889
rect 4833 867 4933 868
rect 4890 831 4932 867
rect 4781 808 4932 831
rect 4781 790 4799 808
rect 4817 793 4932 808
rect 4817 790 4838 793
rect 4781 771 4838 790
rect 99 630 156 649
rect 99 627 120 630
rect 5 612 120 627
rect 138 612 156 630
rect 5 589 156 612
rect 4777 681 4838 697
rect 4777 677 4933 681
rect 5 553 47 589
rect 4 552 104 553
rect 4 531 160 552
rect 4 513 122 531
rect 140 513 160 531
rect 4777 659 4797 677
rect 4815 659 4933 677
rect 4777 638 4933 659
rect 4833 637 4933 638
rect 4890 601 4932 637
rect 4 509 160 513
rect 99 493 160 509
rect 4781 578 4932 601
rect 4781 560 4799 578
rect 4817 563 4932 578
rect 4817 560 4838 563
rect 4781 541 4838 560
rect 99 400 156 419
rect 99 397 120 400
rect 5 382 120 397
rect 138 382 156 400
rect 5 359 156 382
rect 5 323 47 359
rect 4 322 104 323
rect 4 301 160 322
rect 4 283 122 301
rect 140 283 160 301
rect 4777 452 4838 468
rect 4777 448 4933 452
rect 4777 430 4797 448
rect 4815 430 4933 448
rect 4777 409 4933 430
rect 4833 408 4933 409
rect 4890 372 4932 408
rect 4781 349 4932 372
rect 4 279 160 283
rect 99 263 160 279
rect 4781 331 4799 349
rect 4817 334 4932 349
rect 4817 331 4838 334
rect 4781 312 4838 331
rect 4777 265 4838 281
rect 4777 261 4933 265
rect 4777 243 4797 261
rect 4815 243 4933 261
rect 4777 222 4933 243
rect 4833 221 4933 222
rect 4890 185 4932 221
rect 4781 162 4932 185
rect 4781 144 4799 162
rect 4817 147 4932 162
rect 4817 144 4838 147
rect 4781 125 4838 144
<< locali >>
rect 4137 8909 4175 8911
rect 4137 8876 4823 8909
rect 105 8769 144 8826
rect 3729 8788 3897 8789
rect 4137 8788 4175 8876
rect 4436 8858 4483 8876
rect 4400 8819 4512 8858
rect 4783 8852 4823 8876
rect 4400 8818 4443 8819
rect 105 8767 153 8769
rect 105 8749 116 8767
rect 134 8749 153 8767
rect 3729 8765 4175 8788
rect 4401 8817 4443 8818
rect 4401 8797 4408 8817
rect 4427 8797 4443 8817
rect 4401 8789 4443 8797
rect 4471 8817 4512 8819
rect 4471 8797 4485 8817
rect 4504 8797 4512 8817
rect 4784 8808 4823 8852
rect 4471 8789 4512 8797
rect 4401 8783 4512 8789
rect 3729 8762 4173 8765
rect 3729 8760 3897 8762
rect 105 8740 153 8749
rect 106 8739 153 8740
rect 419 8744 529 8758
rect 419 8741 462 8744
rect 419 8736 423 8741
rect 341 8714 423 8736
rect 452 8714 462 8741
rect 490 8717 497 8744
rect 526 8736 529 8744
rect 526 8717 591 8736
rect 490 8714 591 8717
rect 341 8712 591 8714
rect 109 8676 146 8677
rect 105 8673 146 8676
rect 105 8668 147 8673
rect 105 8650 118 8668
rect 136 8650 147 8668
rect 105 8636 147 8650
rect 185 8636 232 8640
rect 105 8630 232 8636
rect 105 8601 193 8630
rect 222 8601 232 8630
rect 341 8633 378 8712
rect 419 8699 529 8712
rect 493 8643 524 8644
rect 341 8613 350 8633
rect 370 8613 378 8633
rect 341 8603 378 8613
rect 437 8633 524 8643
rect 437 8613 446 8633
rect 466 8613 524 8633
rect 437 8604 524 8613
rect 437 8603 474 8604
rect 105 8597 232 8601
rect 105 8580 144 8597
rect 185 8596 232 8597
rect 105 8562 116 8580
rect 134 8562 144 8580
rect 105 8553 144 8562
rect 106 8552 143 8553
rect 493 8551 524 8604
rect 554 8633 591 8712
rect 762 8709 1155 8729
rect 1175 8709 1178 8729
rect 762 8704 1178 8709
rect 762 8703 1103 8704
rect 706 8643 737 8644
rect 554 8613 563 8633
rect 583 8613 591 8633
rect 554 8603 591 8613
rect 650 8636 737 8643
rect 650 8633 711 8636
rect 650 8613 659 8633
rect 679 8616 711 8633
rect 732 8616 737 8636
rect 679 8613 737 8616
rect 650 8606 737 8613
rect 762 8633 799 8703
rect 1065 8702 1102 8703
rect 914 8643 950 8644
rect 762 8613 771 8633
rect 791 8613 799 8633
rect 650 8604 706 8606
rect 650 8603 687 8604
rect 762 8603 799 8613
rect 858 8633 1006 8643
rect 1106 8640 1202 8642
rect 858 8613 867 8633
rect 887 8613 977 8633
rect 997 8613 1006 8633
rect 858 8604 1006 8613
rect 1064 8633 1202 8640
rect 1064 8613 1073 8633
rect 1093 8613 1202 8633
rect 1064 8604 1202 8613
rect 858 8603 895 8604
rect 914 8552 950 8604
rect 969 8603 1006 8604
rect 1065 8603 1102 8604
rect 385 8550 426 8551
rect 277 8543 426 8550
rect 277 8523 395 8543
rect 415 8523 426 8543
rect 277 8515 426 8523
rect 493 8547 852 8551
rect 493 8542 815 8547
rect 493 8518 606 8542
rect 630 8523 815 8542
rect 839 8523 852 8547
rect 630 8518 852 8523
rect 493 8515 852 8518
rect 914 8515 949 8552
rect 1017 8549 1117 8552
rect 1017 8545 1084 8549
rect 1017 8519 1029 8545
rect 1055 8523 1084 8545
rect 1110 8523 1117 8549
rect 1055 8519 1117 8523
rect 1017 8515 1117 8519
rect 493 8494 524 8515
rect 914 8494 950 8515
rect 336 8493 373 8494
rect 110 8490 144 8491
rect 109 8481 146 8490
rect 109 8463 118 8481
rect 136 8463 146 8481
rect 109 8453 146 8463
rect 335 8484 373 8493
rect 335 8464 344 8484
rect 364 8464 373 8484
rect 335 8456 373 8464
rect 439 8488 524 8494
rect 549 8493 586 8494
rect 439 8468 447 8488
rect 467 8468 524 8488
rect 439 8460 524 8468
rect 548 8484 586 8493
rect 548 8464 557 8484
rect 577 8464 586 8484
rect 439 8459 475 8460
rect 548 8456 586 8464
rect 652 8488 737 8494
rect 757 8493 794 8494
rect 652 8468 660 8488
rect 680 8487 737 8488
rect 680 8468 709 8487
rect 652 8467 709 8468
rect 730 8467 737 8487
rect 652 8460 737 8467
rect 756 8484 794 8493
rect 756 8464 765 8484
rect 785 8464 794 8484
rect 652 8459 688 8460
rect 756 8456 794 8464
rect 860 8488 1004 8494
rect 860 8468 868 8488
rect 888 8487 976 8488
rect 888 8468 919 8487
rect 860 8467 919 8468
rect 944 8468 976 8487
rect 996 8468 1004 8488
rect 944 8467 1004 8468
rect 860 8460 1004 8467
rect 860 8459 896 8460
rect 968 8459 1004 8460
rect 1070 8493 1107 8494
rect 1070 8492 1108 8493
rect 1070 8484 1134 8492
rect 1070 8464 1079 8484
rect 1099 8470 1134 8484
rect 1154 8470 1157 8490
rect 1099 8465 1157 8470
rect 1099 8464 1134 8465
rect 110 8425 144 8453
rect 336 8427 373 8456
rect 337 8425 373 8427
rect 549 8425 586 8456
rect 110 8424 282 8425
rect 110 8392 296 8424
rect 337 8403 586 8425
rect 757 8424 794 8456
rect 1070 8452 1134 8464
rect 1174 8426 1201 8604
rect 3729 8582 3756 8760
rect 3796 8722 3860 8734
rect 4136 8730 4173 8762
rect 4344 8761 4593 8783
rect 4344 8730 4381 8761
rect 4557 8759 4593 8761
rect 4557 8730 4594 8759
rect 3796 8721 3831 8722
rect 3773 8716 3831 8721
rect 3773 8696 3776 8716
rect 3796 8702 3831 8716
rect 3851 8702 3860 8722
rect 3796 8694 3860 8702
rect 3822 8693 3860 8694
rect 3823 8692 3860 8693
rect 3926 8726 3962 8727
rect 4034 8726 4070 8727
rect 3926 8721 4070 8726
rect 3926 8718 3988 8721
rect 3926 8698 3934 8718
rect 3954 8701 3988 8718
rect 4011 8718 4070 8721
rect 4011 8701 4042 8718
rect 3954 8698 4042 8701
rect 4062 8698 4070 8718
rect 3926 8692 4070 8698
rect 4136 8722 4174 8730
rect 4242 8726 4278 8727
rect 4136 8702 4145 8722
rect 4165 8702 4174 8722
rect 4136 8693 4174 8702
rect 4193 8719 4278 8726
rect 4193 8699 4200 8719
rect 4221 8718 4278 8719
rect 4221 8699 4250 8718
rect 4193 8698 4250 8699
rect 4270 8698 4278 8718
rect 4136 8692 4173 8693
rect 4193 8692 4278 8698
rect 4344 8722 4382 8730
rect 4455 8726 4491 8727
rect 4344 8702 4353 8722
rect 4373 8702 4382 8722
rect 4344 8693 4382 8702
rect 4406 8718 4491 8726
rect 4406 8698 4463 8718
rect 4483 8698 4491 8718
rect 4344 8692 4381 8693
rect 4406 8692 4491 8698
rect 4557 8722 4595 8730
rect 4557 8702 4566 8722
rect 4586 8702 4595 8722
rect 4557 8693 4595 8702
rect 4557 8692 4594 8693
rect 3980 8671 4016 8692
rect 4406 8671 4437 8692
rect 3813 8667 3913 8671
rect 3813 8663 3875 8667
rect 3813 8637 3820 8663
rect 3846 8641 3875 8663
rect 3901 8641 3913 8667
rect 3846 8637 3913 8641
rect 3813 8634 3913 8637
rect 3981 8634 4016 8671
rect 4078 8668 4437 8671
rect 4078 8663 4300 8668
rect 4078 8639 4091 8663
rect 4115 8644 4300 8663
rect 4324 8644 4437 8668
rect 4115 8639 4437 8644
rect 4078 8635 4437 8639
rect 4504 8663 4653 8671
rect 4504 8643 4515 8663
rect 4535 8643 4653 8663
rect 4504 8636 4653 8643
rect 4504 8635 4545 8636
rect 3828 8582 3865 8583
rect 3924 8582 3961 8583
rect 3980 8582 4016 8634
rect 4035 8582 4072 8583
rect 3728 8573 3866 8582
rect 3728 8553 3837 8573
rect 3857 8553 3866 8573
rect 3728 8546 3866 8553
rect 3924 8573 4072 8582
rect 3924 8553 3933 8573
rect 3953 8553 4043 8573
rect 4063 8553 4072 8573
rect 3728 8544 3824 8546
rect 3924 8543 4072 8553
rect 4131 8573 4168 8583
rect 4243 8582 4280 8583
rect 4224 8580 4280 8582
rect 4131 8553 4139 8573
rect 4159 8553 4168 8573
rect 3980 8542 4016 8543
rect 1357 8500 1467 8514
rect 1357 8497 1400 8500
rect 1357 8492 1361 8497
rect 1033 8424 1201 8426
rect 757 8418 1201 8424
rect 110 8360 144 8392
rect 106 8351 144 8360
rect 106 8333 116 8351
rect 134 8333 144 8351
rect 106 8327 144 8333
rect 262 8329 296 8392
rect 418 8397 529 8403
rect 418 8389 459 8397
rect 418 8369 426 8389
rect 445 8369 459 8389
rect 418 8367 459 8369
rect 487 8389 529 8397
rect 487 8369 503 8389
rect 522 8369 529 8389
rect 487 8367 529 8369
rect 418 8352 529 8367
rect 756 8398 1201 8418
rect 756 8329 794 8398
rect 1033 8397 1201 8398
rect 1279 8470 1361 8492
rect 1390 8470 1400 8497
rect 1428 8473 1435 8500
rect 1464 8492 1467 8500
rect 3462 8509 3573 8524
rect 3462 8507 3504 8509
rect 1464 8473 1529 8492
rect 1428 8470 1529 8473
rect 1279 8468 1529 8470
rect 1279 8389 1316 8468
rect 1357 8455 1467 8468
rect 1431 8399 1462 8400
rect 1279 8369 1288 8389
rect 1308 8369 1316 8389
rect 1279 8359 1316 8369
rect 1375 8389 1462 8399
rect 1375 8369 1384 8389
rect 1404 8369 1462 8389
rect 1375 8360 1462 8369
rect 1375 8359 1412 8360
rect 106 8323 143 8327
rect 262 8318 794 8329
rect 261 8302 794 8318
rect 1431 8307 1462 8360
rect 1492 8389 1529 8468
rect 1700 8465 2093 8485
rect 2113 8465 2116 8485
rect 3195 8480 3236 8489
rect 1700 8460 2116 8465
rect 2790 8478 2958 8479
rect 3195 8478 3204 8480
rect 1700 8459 2041 8460
rect 1644 8399 1675 8400
rect 1492 8369 1501 8389
rect 1521 8369 1529 8389
rect 1492 8359 1529 8369
rect 1588 8392 1675 8399
rect 1588 8389 1649 8392
rect 1588 8369 1597 8389
rect 1617 8372 1649 8389
rect 1670 8372 1675 8392
rect 1617 8369 1675 8372
rect 1588 8362 1675 8369
rect 1700 8389 1737 8459
rect 2003 8458 2040 8459
rect 2790 8458 3204 8478
rect 3230 8458 3236 8480
rect 3462 8487 3469 8507
rect 3488 8487 3504 8507
rect 3462 8479 3504 8487
rect 3532 8507 3573 8509
rect 3532 8487 3546 8507
rect 3565 8487 3573 8507
rect 3532 8479 3573 8487
rect 3828 8483 3865 8484
rect 4131 8483 4168 8553
rect 4193 8573 4280 8580
rect 4193 8570 4251 8573
rect 4193 8550 4198 8570
rect 4219 8553 4251 8570
rect 4271 8553 4280 8573
rect 4219 8550 4280 8553
rect 4193 8543 4280 8550
rect 4339 8573 4376 8583
rect 4339 8553 4347 8573
rect 4367 8553 4376 8573
rect 4193 8542 4224 8543
rect 3827 8482 4168 8483
rect 3462 8473 3573 8479
rect 3752 8477 4168 8482
rect 2790 8452 3236 8458
rect 2790 8450 2958 8452
rect 1852 8399 1888 8400
rect 1700 8369 1709 8389
rect 1729 8369 1737 8389
rect 1588 8360 1644 8362
rect 1588 8359 1625 8360
rect 1700 8359 1737 8369
rect 1796 8389 1944 8399
rect 2044 8396 2140 8398
rect 1796 8369 1805 8389
rect 1825 8369 1915 8389
rect 1935 8369 1944 8389
rect 1796 8360 1944 8369
rect 2002 8389 2140 8396
rect 2002 8369 2011 8389
rect 2031 8369 2140 8389
rect 2002 8360 2140 8369
rect 1796 8359 1833 8360
rect 1852 8308 1888 8360
rect 1907 8359 1944 8360
rect 2003 8359 2040 8360
rect 1323 8306 1364 8307
rect 261 8301 775 8302
rect 1215 8299 1364 8306
rect 1215 8279 1333 8299
rect 1353 8279 1364 8299
rect 1215 8271 1364 8279
rect 1431 8303 1790 8307
rect 1431 8298 1753 8303
rect 1431 8274 1544 8298
rect 1568 8279 1753 8298
rect 1777 8279 1790 8303
rect 1568 8274 1790 8279
rect 1431 8271 1790 8274
rect 1852 8271 1887 8308
rect 1955 8305 2055 8308
rect 1955 8301 2022 8305
rect 1955 8275 1967 8301
rect 1993 8279 2022 8301
rect 2048 8279 2055 8305
rect 1993 8275 2055 8279
rect 1955 8271 2055 8275
rect 109 8260 146 8261
rect 107 8252 147 8260
rect 107 8234 118 8252
rect 136 8234 147 8252
rect 1431 8250 1462 8271
rect 1852 8250 1888 8271
rect 1274 8249 1311 8250
rect 107 8186 147 8234
rect 1273 8240 1311 8249
rect 1273 8220 1282 8240
rect 1302 8220 1311 8240
rect 1273 8212 1311 8220
rect 1377 8244 1462 8250
rect 1487 8249 1524 8250
rect 1377 8224 1385 8244
rect 1405 8224 1462 8244
rect 1377 8216 1462 8224
rect 1486 8240 1524 8249
rect 1486 8220 1495 8240
rect 1515 8220 1524 8240
rect 1377 8215 1413 8216
rect 1486 8212 1524 8220
rect 1590 8244 1675 8250
rect 1695 8249 1732 8250
rect 1590 8224 1598 8244
rect 1618 8243 1675 8244
rect 1618 8224 1647 8243
rect 1590 8223 1647 8224
rect 1668 8223 1675 8243
rect 1590 8216 1675 8223
rect 1694 8240 1732 8249
rect 1694 8220 1703 8240
rect 1723 8220 1732 8240
rect 1590 8215 1626 8216
rect 1694 8212 1732 8220
rect 1798 8244 1942 8250
rect 1798 8224 1806 8244
rect 1826 8227 1862 8244
rect 1882 8227 1914 8244
rect 1826 8224 1914 8227
rect 1934 8224 1942 8244
rect 1798 8216 1942 8224
rect 1798 8215 1834 8216
rect 1906 8215 1942 8216
rect 2008 8249 2045 8250
rect 2008 8248 2046 8249
rect 2008 8240 2072 8248
rect 2008 8220 2017 8240
rect 2037 8226 2072 8240
rect 2092 8226 2095 8246
rect 2037 8221 2095 8226
rect 2037 8220 2072 8221
rect 418 8190 528 8204
rect 418 8187 461 8190
rect 107 8179 232 8186
rect 418 8182 422 8187
rect 107 8160 199 8179
rect 224 8160 232 8179
rect 107 8150 232 8160
rect 340 8160 422 8182
rect 451 8160 461 8187
rect 489 8163 496 8190
rect 525 8182 528 8190
rect 1274 8183 1311 8212
rect 525 8163 590 8182
rect 1275 8181 1311 8183
rect 1487 8181 1524 8212
rect 1695 8185 1732 8212
rect 2008 8208 2072 8220
rect 489 8160 590 8163
rect 340 8158 590 8160
rect 107 8130 147 8150
rect 106 8121 147 8130
rect 106 8103 116 8121
rect 134 8103 147 8121
rect 106 8094 147 8103
rect 106 8093 143 8094
rect 340 8079 377 8158
rect 418 8145 528 8158
rect 492 8089 523 8090
rect 340 8059 349 8079
rect 369 8059 377 8079
rect 340 8049 377 8059
rect 436 8079 523 8089
rect 436 8059 445 8079
rect 465 8059 523 8079
rect 436 8050 523 8059
rect 436 8049 473 8050
rect 109 8027 146 8031
rect 106 8022 146 8027
rect 106 8004 118 8022
rect 136 8004 146 8022
rect 106 7824 146 8004
rect 492 7997 523 8050
rect 553 8079 590 8158
rect 761 8155 1154 8175
rect 1174 8155 1177 8175
rect 1275 8159 1524 8181
rect 1693 8180 1734 8185
rect 2112 8182 2139 8360
rect 2790 8272 2817 8450
rect 3195 8447 3236 8452
rect 3405 8451 3654 8473
rect 3752 8457 3755 8477
rect 3775 8457 4168 8477
rect 4339 8474 4376 8553
rect 4406 8582 4437 8635
rect 4783 8628 4823 8808
rect 4783 8610 4793 8628
rect 4811 8610 4823 8628
rect 4783 8605 4823 8610
rect 4783 8601 4820 8605
rect 4456 8582 4493 8583
rect 4406 8573 4493 8582
rect 4406 8553 4464 8573
rect 4484 8553 4493 8573
rect 4406 8543 4493 8553
rect 4552 8573 4589 8583
rect 4552 8553 4560 8573
rect 4580 8553 4589 8573
rect 4406 8542 4437 8543
rect 4401 8474 4511 8487
rect 4552 8474 4589 8553
rect 4786 8538 4823 8539
rect 4782 8529 4823 8538
rect 4782 8511 4795 8529
rect 4813 8511 4823 8529
rect 4782 8502 4823 8511
rect 4782 8482 4822 8502
rect 4339 8472 4589 8474
rect 4339 8469 4440 8472
rect 2857 8412 2921 8424
rect 3197 8420 3234 8447
rect 3405 8420 3442 8451
rect 3618 8449 3654 8451
rect 4339 8450 4404 8469
rect 3618 8420 3655 8449
rect 4401 8442 4404 8450
rect 4433 8442 4440 8469
rect 4468 8445 4478 8472
rect 4507 8450 4589 8472
rect 4697 8472 4822 8482
rect 4697 8453 4705 8472
rect 4730 8453 4822 8472
rect 4507 8445 4511 8450
rect 4697 8446 4822 8453
rect 4468 8442 4511 8445
rect 4401 8428 4511 8442
rect 2857 8411 2892 8412
rect 2834 8406 2892 8411
rect 2834 8386 2837 8406
rect 2857 8392 2892 8406
rect 2912 8392 2921 8412
rect 2857 8384 2921 8392
rect 2883 8383 2921 8384
rect 2884 8382 2921 8383
rect 2987 8416 3023 8417
rect 3095 8416 3131 8417
rect 2987 8408 3131 8416
rect 2987 8388 2995 8408
rect 3015 8388 3103 8408
rect 3123 8388 3131 8408
rect 2987 8382 3131 8388
rect 3197 8412 3235 8420
rect 3303 8416 3339 8417
rect 3197 8392 3206 8412
rect 3226 8392 3235 8412
rect 3197 8383 3235 8392
rect 3254 8409 3339 8416
rect 3254 8389 3261 8409
rect 3282 8408 3339 8409
rect 3282 8389 3311 8408
rect 3254 8388 3311 8389
rect 3331 8388 3339 8408
rect 3197 8382 3234 8383
rect 3254 8382 3339 8388
rect 3405 8412 3443 8420
rect 3516 8416 3552 8417
rect 3405 8392 3414 8412
rect 3434 8392 3443 8412
rect 3405 8383 3443 8392
rect 3467 8408 3552 8416
rect 3467 8388 3524 8408
rect 3544 8388 3552 8408
rect 3405 8382 3442 8383
rect 3467 8382 3552 8388
rect 3618 8412 3656 8420
rect 3618 8392 3627 8412
rect 3647 8392 3656 8412
rect 3618 8383 3656 8392
rect 4782 8398 4822 8446
rect 3618 8382 3655 8383
rect 3041 8361 3077 8382
rect 3467 8361 3498 8382
rect 4782 8380 4793 8398
rect 4811 8380 4822 8398
rect 4782 8372 4822 8380
rect 4783 8371 4820 8372
rect 2874 8357 2974 8361
rect 2874 8353 2936 8357
rect 2874 8327 2881 8353
rect 2907 8331 2936 8353
rect 2962 8331 2974 8357
rect 2907 8327 2974 8331
rect 2874 8324 2974 8327
rect 3042 8324 3077 8361
rect 3139 8358 3498 8361
rect 3139 8353 3361 8358
rect 3139 8329 3152 8353
rect 3176 8334 3361 8353
rect 3385 8334 3498 8358
rect 3176 8329 3498 8334
rect 3139 8325 3498 8329
rect 3565 8353 3714 8361
rect 3565 8333 3576 8353
rect 3596 8333 3714 8353
rect 3565 8326 3714 8333
rect 4154 8330 4668 8331
rect 3565 8325 3606 8326
rect 3041 8289 3077 8324
rect 2889 8272 2926 8273
rect 2985 8272 3022 8273
rect 3041 8272 3048 8289
rect 2789 8263 2927 8272
rect 2789 8243 2898 8263
rect 2918 8243 2927 8263
rect 2789 8236 2927 8243
rect 2985 8263 3048 8272
rect 2985 8243 2994 8263
rect 3014 8248 3048 8263
rect 3069 8272 3077 8289
rect 3096 8272 3133 8273
rect 3069 8263 3133 8272
rect 3069 8248 3104 8263
rect 3014 8243 3104 8248
rect 3124 8243 3133 8263
rect 2789 8234 2885 8236
rect 2985 8233 3133 8243
rect 3192 8263 3229 8273
rect 3304 8272 3341 8273
rect 3285 8270 3341 8272
rect 3192 8243 3200 8263
rect 3220 8243 3229 8263
rect 3041 8232 3077 8233
rect 1971 8180 2139 8182
rect 1693 8174 2139 8180
rect 761 8150 1177 8155
rect 1356 8153 1467 8159
rect 761 8149 1102 8150
rect 705 8089 736 8090
rect 553 8059 562 8079
rect 582 8059 590 8079
rect 553 8049 590 8059
rect 649 8082 736 8089
rect 649 8079 710 8082
rect 649 8059 658 8079
rect 678 8062 710 8079
rect 731 8062 736 8082
rect 678 8059 736 8062
rect 649 8052 736 8059
rect 761 8079 798 8149
rect 1064 8148 1101 8149
rect 1356 8145 1397 8153
rect 1356 8125 1364 8145
rect 1383 8125 1397 8145
rect 1356 8123 1397 8125
rect 1425 8145 1467 8153
rect 1425 8125 1441 8145
rect 1460 8125 1467 8145
rect 1693 8152 1699 8174
rect 1725 8154 2139 8174
rect 2889 8173 2926 8174
rect 3192 8173 3229 8243
rect 3254 8263 3341 8270
rect 3254 8260 3312 8263
rect 3254 8240 3259 8260
rect 3280 8243 3312 8260
rect 3332 8243 3341 8263
rect 3280 8240 3341 8243
rect 3254 8233 3341 8240
rect 3400 8263 3437 8273
rect 3400 8243 3408 8263
rect 3428 8243 3437 8263
rect 3254 8232 3285 8233
rect 2888 8172 3229 8173
rect 1725 8152 1734 8154
rect 1971 8153 2139 8154
rect 2813 8171 3229 8172
rect 2813 8167 3189 8171
rect 1693 8143 1734 8152
rect 2813 8147 2816 8167
rect 2836 8154 3189 8167
rect 3221 8154 3229 8171
rect 2836 8147 3229 8154
rect 3400 8164 3437 8243
rect 3467 8272 3498 8325
rect 4135 8314 4668 8330
rect 4135 8303 4667 8314
rect 4786 8305 4823 8309
rect 3517 8272 3554 8273
rect 3467 8263 3554 8272
rect 3467 8243 3525 8263
rect 3545 8243 3554 8263
rect 3467 8233 3554 8243
rect 3613 8263 3650 8273
rect 3613 8243 3621 8263
rect 3641 8243 3650 8263
rect 3467 8232 3498 8233
rect 3462 8164 3572 8177
rect 3613 8164 3650 8243
rect 3400 8162 3650 8164
rect 3400 8159 3501 8162
rect 3400 8140 3465 8159
rect 1425 8123 1467 8125
rect 1356 8108 1467 8123
rect 3462 8132 3465 8140
rect 3494 8132 3501 8159
rect 3529 8135 3539 8162
rect 3568 8140 3650 8162
rect 3728 8234 3896 8235
rect 4135 8234 4173 8303
rect 3728 8214 4173 8234
rect 4400 8265 4511 8280
rect 4400 8263 4442 8265
rect 4400 8243 4407 8263
rect 4426 8243 4442 8263
rect 4400 8235 4442 8243
rect 4470 8263 4511 8265
rect 4470 8243 4484 8263
rect 4503 8243 4511 8263
rect 4470 8235 4511 8243
rect 4400 8229 4511 8235
rect 4633 8240 4667 8303
rect 4785 8299 4823 8305
rect 4785 8281 4795 8299
rect 4813 8281 4823 8299
rect 4785 8272 4823 8281
rect 4785 8240 4819 8272
rect 3728 8208 4172 8214
rect 3728 8206 3896 8208
rect 3568 8135 3572 8140
rect 3529 8132 3572 8135
rect 3462 8118 3572 8132
rect 913 8089 949 8090
rect 761 8059 770 8079
rect 790 8059 798 8079
rect 649 8050 705 8052
rect 649 8049 686 8050
rect 761 8049 798 8059
rect 857 8079 1005 8089
rect 1105 8086 1201 8088
rect 857 8059 866 8079
rect 886 8059 976 8079
rect 996 8059 1005 8079
rect 857 8050 1005 8059
rect 1063 8079 1201 8086
rect 1063 8059 1072 8079
rect 1092 8059 1201 8079
rect 1063 8050 1201 8059
rect 857 8049 894 8050
rect 913 7998 949 8050
rect 968 8049 1005 8050
rect 1064 8049 1101 8050
rect 384 7996 425 7997
rect 276 7989 425 7996
rect 276 7969 394 7989
rect 414 7969 425 7989
rect 276 7961 425 7969
rect 492 7993 851 7997
rect 492 7988 814 7993
rect 492 7964 605 7988
rect 629 7969 814 7988
rect 838 7969 851 7993
rect 629 7964 851 7969
rect 492 7961 851 7964
rect 913 7961 948 7998
rect 1016 7995 1116 7998
rect 1016 7991 1083 7995
rect 1016 7965 1028 7991
rect 1054 7969 1083 7991
rect 1109 7969 1116 7995
rect 1054 7965 1116 7969
rect 1016 7961 1116 7965
rect 492 7940 523 7961
rect 913 7940 949 7961
rect 335 7939 372 7940
rect 334 7930 372 7939
rect 334 7910 343 7930
rect 363 7910 372 7930
rect 334 7902 372 7910
rect 438 7934 523 7940
rect 548 7939 585 7940
rect 438 7914 446 7934
rect 466 7914 523 7934
rect 438 7906 523 7914
rect 547 7930 585 7939
rect 547 7910 556 7930
rect 576 7910 585 7930
rect 438 7905 474 7906
rect 547 7902 585 7910
rect 651 7934 736 7940
rect 756 7939 793 7940
rect 651 7914 659 7934
rect 679 7933 736 7934
rect 679 7914 708 7933
rect 651 7913 708 7914
rect 729 7913 736 7933
rect 651 7906 736 7913
rect 755 7930 793 7939
rect 755 7910 764 7930
rect 784 7910 793 7930
rect 651 7905 687 7906
rect 755 7902 793 7910
rect 859 7934 1003 7940
rect 859 7914 867 7934
rect 887 7931 975 7934
rect 887 7914 918 7931
rect 859 7911 918 7914
rect 941 7914 975 7931
rect 995 7914 1003 7934
rect 941 7911 1003 7914
rect 859 7906 1003 7911
rect 859 7905 895 7906
rect 967 7905 1003 7906
rect 1069 7939 1106 7940
rect 1069 7938 1107 7939
rect 1069 7930 1133 7938
rect 1069 7910 1078 7930
rect 1098 7916 1133 7930
rect 1153 7916 1156 7936
rect 1098 7911 1156 7916
rect 1098 7910 1133 7911
rect 335 7873 372 7902
rect 336 7871 372 7873
rect 548 7871 585 7902
rect 336 7849 585 7871
rect 756 7870 793 7902
rect 1069 7898 1133 7910
rect 1173 7872 1200 8050
rect 3728 8028 3755 8206
rect 3795 8168 3859 8180
rect 4135 8176 4172 8208
rect 4343 8207 4592 8229
rect 4633 8208 4819 8240
rect 4647 8207 4819 8208
rect 4343 8176 4380 8207
rect 4556 8205 4592 8207
rect 4556 8176 4593 8205
rect 4785 8179 4819 8207
rect 3795 8167 3830 8168
rect 3772 8162 3830 8167
rect 3772 8142 3775 8162
rect 3795 8148 3830 8162
rect 3850 8148 3859 8168
rect 3795 8140 3859 8148
rect 3821 8139 3859 8140
rect 3822 8138 3859 8139
rect 3925 8172 3961 8173
rect 4033 8172 4069 8173
rect 3925 8165 4069 8172
rect 3925 8164 3985 8165
rect 3925 8144 3933 8164
rect 3953 8145 3985 8164
rect 4010 8164 4069 8165
rect 4010 8145 4041 8164
rect 3953 8144 4041 8145
rect 4061 8144 4069 8164
rect 3925 8138 4069 8144
rect 4135 8168 4173 8176
rect 4241 8172 4277 8173
rect 4135 8148 4144 8168
rect 4164 8148 4173 8168
rect 4135 8139 4173 8148
rect 4192 8165 4277 8172
rect 4192 8145 4199 8165
rect 4220 8164 4277 8165
rect 4220 8145 4249 8164
rect 4192 8144 4249 8145
rect 4269 8144 4277 8164
rect 4135 8138 4172 8139
rect 4192 8138 4277 8144
rect 4343 8168 4381 8176
rect 4454 8172 4490 8173
rect 4343 8148 4352 8168
rect 4372 8148 4381 8168
rect 4343 8139 4381 8148
rect 4405 8164 4490 8172
rect 4405 8144 4462 8164
rect 4482 8144 4490 8164
rect 4343 8138 4380 8139
rect 4405 8138 4490 8144
rect 4556 8168 4594 8176
rect 4556 8148 4565 8168
rect 4585 8148 4594 8168
rect 4556 8139 4594 8148
rect 4783 8169 4820 8179
rect 4783 8151 4793 8169
rect 4811 8151 4820 8169
rect 4783 8142 4820 8151
rect 4785 8141 4819 8142
rect 4556 8138 4593 8139
rect 3979 8117 4015 8138
rect 4405 8117 4436 8138
rect 3812 8113 3912 8117
rect 3812 8109 3874 8113
rect 3812 8083 3819 8109
rect 3845 8087 3874 8109
rect 3900 8087 3912 8113
rect 3845 8083 3912 8087
rect 3812 8080 3912 8083
rect 3980 8080 4015 8117
rect 4077 8114 4436 8117
rect 4077 8109 4299 8114
rect 4077 8085 4090 8109
rect 4114 8090 4299 8109
rect 4323 8090 4436 8114
rect 4114 8085 4436 8090
rect 4077 8081 4436 8085
rect 4503 8109 4652 8117
rect 4503 8089 4514 8109
rect 4534 8089 4652 8109
rect 4503 8082 4652 8089
rect 4503 8081 4544 8082
rect 3827 8028 3864 8029
rect 3923 8028 3960 8029
rect 3979 8028 4015 8080
rect 4034 8028 4071 8029
rect 3727 8019 3865 8028
rect 3322 7998 3433 8013
rect 3322 7996 3364 7998
rect 2992 7975 3097 7977
rect 2648 7967 2818 7968
rect 2992 7967 3041 7975
rect 2648 7948 3041 7967
rect 3072 7948 3097 7975
rect 3322 7976 3329 7996
rect 3348 7976 3364 7996
rect 3322 7968 3364 7976
rect 3392 7996 3433 7998
rect 3392 7976 3406 7996
rect 3425 7976 3433 7996
rect 3727 7999 3836 8019
rect 3856 7999 3865 8019
rect 3727 7992 3865 7999
rect 3923 8019 4071 8028
rect 3923 7999 3932 8019
rect 3952 7999 4042 8019
rect 4062 7999 4071 8019
rect 3727 7990 3823 7992
rect 3923 7989 4071 7999
rect 4130 8019 4167 8029
rect 4242 8028 4279 8029
rect 4223 8026 4279 8028
rect 4130 7999 4138 8019
rect 4158 7999 4167 8019
rect 3979 7988 4015 7989
rect 3392 7968 3433 7976
rect 3322 7962 3433 7968
rect 2648 7941 3097 7948
rect 2648 7939 2818 7941
rect 1498 7908 1608 7922
rect 1498 7905 1541 7908
rect 1498 7900 1502 7905
rect 1032 7870 1200 7872
rect 756 7867 1200 7870
rect 417 7843 528 7849
rect 417 7835 458 7843
rect 106 7780 145 7824
rect 417 7815 425 7835
rect 444 7815 458 7835
rect 417 7813 458 7815
rect 486 7835 528 7843
rect 486 7815 502 7835
rect 521 7815 528 7835
rect 486 7813 528 7815
rect 417 7798 528 7813
rect 754 7844 1200 7867
rect 106 7756 146 7780
rect 446 7756 493 7758
rect 754 7756 792 7844
rect 1032 7843 1200 7844
rect 1420 7878 1502 7900
rect 1531 7878 1541 7905
rect 1569 7881 1576 7908
rect 1605 7900 1608 7908
rect 1605 7881 1670 7900
rect 1569 7878 1670 7881
rect 1420 7876 1670 7878
rect 1420 7797 1457 7876
rect 1498 7863 1608 7876
rect 1572 7807 1603 7808
rect 1420 7777 1429 7797
rect 1449 7777 1457 7797
rect 1420 7767 1457 7777
rect 1516 7797 1603 7807
rect 1516 7777 1525 7797
rect 1545 7777 1603 7797
rect 1516 7768 1603 7777
rect 1516 7767 1553 7768
rect 106 7723 792 7756
rect 106 7666 145 7723
rect 754 7721 792 7723
rect 1572 7715 1603 7768
rect 1633 7797 1670 7876
rect 1841 7889 2234 7893
rect 1841 7872 1860 7889
rect 1880 7873 2234 7889
rect 2254 7873 2257 7893
rect 1880 7872 2257 7873
rect 1841 7868 2257 7872
rect 1841 7867 2182 7868
rect 1785 7807 1816 7808
rect 1633 7777 1642 7797
rect 1662 7777 1670 7797
rect 1633 7767 1670 7777
rect 1729 7800 1816 7807
rect 1729 7797 1790 7800
rect 1729 7777 1738 7797
rect 1758 7780 1790 7797
rect 1811 7780 1816 7800
rect 1758 7777 1816 7780
rect 1729 7770 1816 7777
rect 1841 7797 1878 7867
rect 2144 7866 2181 7867
rect 1993 7807 2029 7808
rect 1841 7777 1850 7797
rect 1870 7777 1878 7797
rect 1729 7768 1785 7770
rect 1729 7767 1766 7768
rect 1841 7767 1878 7777
rect 1937 7797 2085 7807
rect 2185 7804 2281 7806
rect 1937 7777 1946 7797
rect 1966 7777 2056 7797
rect 2076 7777 2085 7797
rect 1937 7768 2085 7777
rect 2143 7797 2281 7804
rect 2143 7777 2152 7797
rect 2172 7777 2281 7797
rect 2143 7768 2281 7777
rect 1937 7767 1974 7768
rect 1993 7716 2029 7768
rect 2048 7767 2085 7768
rect 2144 7767 2181 7768
rect 1464 7714 1505 7715
rect 1356 7707 1505 7714
rect 1356 7687 1474 7707
rect 1494 7687 1505 7707
rect 1356 7679 1505 7687
rect 1572 7711 1931 7715
rect 1572 7706 1894 7711
rect 1572 7682 1685 7706
rect 1709 7687 1894 7706
rect 1918 7687 1931 7711
rect 1709 7682 1931 7687
rect 1572 7679 1931 7682
rect 1993 7679 2028 7716
rect 2096 7713 2196 7716
rect 2096 7709 2163 7713
rect 2096 7683 2108 7709
rect 2134 7687 2163 7709
rect 2189 7687 2196 7713
rect 2134 7683 2196 7687
rect 2096 7679 2196 7683
rect 106 7664 154 7666
rect 106 7646 117 7664
rect 135 7646 154 7664
rect 1572 7658 1603 7679
rect 1993 7658 2029 7679
rect 1415 7657 1452 7658
rect 106 7637 154 7646
rect 107 7636 154 7637
rect 420 7641 530 7655
rect 420 7638 463 7641
rect 420 7633 424 7638
rect 342 7611 424 7633
rect 453 7611 463 7638
rect 491 7614 498 7641
rect 527 7633 530 7641
rect 1414 7648 1452 7657
rect 527 7614 592 7633
rect 1414 7628 1423 7648
rect 1443 7628 1452 7648
rect 491 7611 592 7614
rect 342 7609 592 7611
rect 110 7573 147 7574
rect 106 7570 147 7573
rect 106 7565 148 7570
rect 106 7547 119 7565
rect 137 7547 148 7565
rect 106 7533 148 7547
rect 186 7533 233 7537
rect 106 7527 233 7533
rect 106 7498 194 7527
rect 223 7498 233 7527
rect 342 7530 379 7609
rect 420 7596 530 7609
rect 494 7540 525 7541
rect 342 7510 351 7530
rect 371 7510 379 7530
rect 342 7500 379 7510
rect 438 7530 525 7540
rect 438 7510 447 7530
rect 467 7510 525 7530
rect 438 7501 525 7510
rect 438 7500 475 7501
rect 106 7494 233 7498
rect 106 7477 145 7494
rect 186 7493 233 7494
rect 106 7459 117 7477
rect 135 7459 145 7477
rect 106 7450 145 7459
rect 107 7449 144 7450
rect 494 7448 525 7501
rect 555 7530 592 7609
rect 763 7606 1156 7626
rect 1176 7606 1179 7626
rect 1414 7620 1452 7628
rect 1518 7652 1603 7658
rect 1628 7657 1665 7658
rect 1518 7632 1526 7652
rect 1546 7632 1603 7652
rect 1518 7624 1603 7632
rect 1627 7648 1665 7657
rect 1627 7628 1636 7648
rect 1656 7628 1665 7648
rect 1518 7623 1554 7624
rect 1627 7620 1665 7628
rect 1731 7652 1816 7658
rect 1836 7657 1873 7658
rect 1731 7632 1739 7652
rect 1759 7651 1816 7652
rect 1759 7632 1788 7651
rect 1731 7631 1788 7632
rect 1809 7631 1816 7651
rect 1731 7624 1816 7631
rect 1835 7648 1873 7657
rect 1835 7628 1844 7648
rect 1864 7628 1873 7648
rect 1731 7623 1767 7624
rect 1835 7620 1873 7628
rect 1939 7652 2083 7658
rect 1939 7632 1947 7652
rect 1967 7650 2055 7652
rect 1967 7632 1996 7650
rect 1939 7629 1996 7632
rect 2023 7632 2055 7650
rect 2075 7632 2083 7652
rect 2023 7629 2083 7632
rect 1939 7624 2083 7629
rect 1939 7623 1975 7624
rect 2047 7623 2083 7624
rect 2149 7657 2186 7658
rect 2149 7656 2187 7657
rect 2149 7648 2213 7656
rect 2149 7628 2158 7648
rect 2178 7634 2213 7648
rect 2233 7634 2236 7654
rect 2178 7629 2236 7634
rect 2178 7628 2213 7629
rect 763 7601 1179 7606
rect 763 7600 1104 7601
rect 707 7540 738 7541
rect 555 7510 564 7530
rect 584 7510 592 7530
rect 555 7500 592 7510
rect 651 7533 738 7540
rect 651 7530 712 7533
rect 651 7510 660 7530
rect 680 7513 712 7530
rect 733 7513 738 7533
rect 680 7510 738 7513
rect 651 7503 738 7510
rect 763 7530 800 7600
rect 1066 7599 1103 7600
rect 1415 7591 1452 7620
rect 1416 7589 1452 7591
rect 1628 7589 1665 7620
rect 1416 7567 1665 7589
rect 1836 7588 1873 7620
rect 2149 7616 2213 7628
rect 2253 7590 2280 7768
rect 2648 7761 2677 7939
rect 2717 7901 2781 7913
rect 3057 7909 3094 7941
rect 3265 7940 3514 7962
rect 3265 7909 3302 7940
rect 3478 7938 3514 7940
rect 3478 7909 3515 7938
rect 3827 7929 3864 7930
rect 4130 7929 4167 7999
rect 4192 8019 4279 8026
rect 4192 8016 4250 8019
rect 4192 7996 4197 8016
rect 4218 7999 4250 8016
rect 4270 7999 4279 8019
rect 4218 7996 4279 7999
rect 4192 7989 4279 7996
rect 4338 8019 4375 8029
rect 4338 7999 4346 8019
rect 4366 7999 4375 8019
rect 4192 7988 4223 7989
rect 3826 7928 4167 7929
rect 3751 7923 4167 7928
rect 2717 7900 2752 7901
rect 2694 7895 2752 7900
rect 2694 7875 2697 7895
rect 2717 7881 2752 7895
rect 2772 7881 2781 7901
rect 2717 7873 2781 7881
rect 2743 7872 2781 7873
rect 2744 7871 2781 7872
rect 2847 7905 2883 7906
rect 2955 7905 2991 7906
rect 2847 7897 2991 7905
rect 2847 7877 2855 7897
rect 2875 7877 2963 7897
rect 2983 7877 2991 7897
rect 2847 7871 2991 7877
rect 3057 7901 3095 7909
rect 3163 7905 3199 7906
rect 3057 7881 3066 7901
rect 3086 7881 3095 7901
rect 3057 7872 3095 7881
rect 3114 7898 3199 7905
rect 3114 7878 3121 7898
rect 3142 7897 3199 7898
rect 3142 7878 3171 7897
rect 3114 7877 3171 7878
rect 3191 7877 3199 7897
rect 3057 7871 3094 7872
rect 3114 7871 3199 7877
rect 3265 7901 3303 7909
rect 3376 7905 3412 7906
rect 3265 7881 3274 7901
rect 3294 7881 3303 7901
rect 3265 7872 3303 7881
rect 3327 7897 3412 7905
rect 3327 7877 3384 7897
rect 3404 7877 3412 7897
rect 3265 7871 3302 7872
rect 3327 7871 3412 7877
rect 3478 7901 3516 7909
rect 3751 7903 3754 7923
rect 3774 7903 4167 7923
rect 4338 7920 4375 7999
rect 4405 8028 4436 8081
rect 4786 8079 4823 8080
rect 4785 8070 4824 8079
rect 4785 8052 4795 8070
rect 4813 8052 4824 8070
rect 4697 8035 4744 8036
rect 4785 8035 4824 8052
rect 4697 8031 4824 8035
rect 4455 8028 4492 8029
rect 4405 8019 4492 8028
rect 4405 7999 4463 8019
rect 4483 7999 4492 8019
rect 4405 7989 4492 7999
rect 4551 8019 4588 8029
rect 4551 7999 4559 8019
rect 4579 7999 4588 8019
rect 4405 7988 4436 7989
rect 4400 7920 4510 7933
rect 4551 7920 4588 7999
rect 4697 8002 4707 8031
rect 4736 8002 4824 8031
rect 4697 7996 4824 8002
rect 4697 7992 4744 7996
rect 4782 7982 4824 7996
rect 4782 7964 4793 7982
rect 4811 7964 4824 7982
rect 4782 7959 4824 7964
rect 4783 7956 4824 7959
rect 4783 7955 4820 7956
rect 4338 7918 4588 7920
rect 4338 7915 4439 7918
rect 3478 7881 3487 7901
rect 3507 7881 3516 7901
rect 4338 7896 4403 7915
rect 3478 7872 3516 7881
rect 4400 7888 4403 7896
rect 4432 7888 4439 7915
rect 4467 7891 4477 7918
rect 4506 7896 4588 7918
rect 4506 7891 4510 7896
rect 4467 7888 4510 7891
rect 4400 7874 4510 7888
rect 4776 7892 4823 7893
rect 4776 7883 4824 7892
rect 3478 7871 3515 7872
rect 2901 7850 2937 7871
rect 3327 7850 3358 7871
rect 4776 7865 4795 7883
rect 4813 7865 4824 7883
rect 4776 7863 4824 7865
rect 2734 7846 2834 7850
rect 2734 7842 2796 7846
rect 2734 7816 2741 7842
rect 2767 7820 2796 7842
rect 2822 7820 2834 7846
rect 2767 7816 2834 7820
rect 2734 7813 2834 7816
rect 2902 7813 2937 7850
rect 2999 7847 3358 7850
rect 2999 7842 3221 7847
rect 2999 7818 3012 7842
rect 3036 7823 3221 7842
rect 3245 7823 3358 7847
rect 3036 7818 3358 7823
rect 2999 7814 3358 7818
rect 3425 7842 3574 7850
rect 3425 7822 3436 7842
rect 3456 7822 3574 7842
rect 3425 7815 3574 7822
rect 3425 7814 3466 7815
rect 2901 7774 2937 7813
rect 2749 7761 2786 7762
rect 2845 7761 2882 7762
rect 2901 7761 2908 7774
rect 2648 7752 2787 7761
rect 2648 7732 2758 7752
rect 2778 7732 2787 7752
rect 2648 7725 2787 7732
rect 2845 7752 2908 7761
rect 2845 7732 2854 7752
rect 2874 7736 2908 7752
rect 2931 7761 2937 7774
rect 2956 7761 2993 7762
rect 2931 7752 2993 7761
rect 2931 7736 2964 7752
rect 2874 7732 2964 7736
rect 2984 7732 2993 7752
rect 2648 7723 2745 7725
rect 2648 7722 2677 7723
rect 2845 7722 2993 7732
rect 3052 7752 3089 7762
rect 3164 7761 3201 7762
rect 3145 7759 3201 7761
rect 3052 7732 3060 7752
rect 3080 7732 3089 7752
rect 2901 7721 2937 7722
rect 2749 7662 2786 7663
rect 3052 7662 3089 7732
rect 3114 7752 3201 7759
rect 3114 7749 3172 7752
rect 3114 7729 3119 7749
rect 3140 7732 3172 7749
rect 3192 7732 3201 7752
rect 3140 7729 3201 7732
rect 3114 7722 3201 7729
rect 3260 7752 3297 7762
rect 3260 7732 3268 7752
rect 3288 7732 3297 7752
rect 3114 7721 3145 7722
rect 2748 7661 3089 7662
rect 2673 7657 3089 7661
rect 2673 7656 3050 7657
rect 2673 7636 2676 7656
rect 2696 7640 3050 7656
rect 3070 7640 3089 7657
rect 2696 7636 3089 7640
rect 3260 7653 3297 7732
rect 3327 7761 3358 7814
rect 4138 7806 4176 7808
rect 4785 7806 4824 7863
rect 4138 7773 4824 7806
rect 3377 7761 3414 7762
rect 3327 7752 3414 7761
rect 3327 7732 3385 7752
rect 3405 7732 3414 7752
rect 3327 7722 3414 7732
rect 3473 7752 3510 7762
rect 3473 7732 3481 7752
rect 3501 7732 3510 7752
rect 3327 7721 3358 7722
rect 3322 7653 3432 7666
rect 3473 7653 3510 7732
rect 3260 7651 3510 7653
rect 3260 7648 3361 7651
rect 3260 7629 3325 7648
rect 3322 7621 3325 7629
rect 3354 7621 3361 7648
rect 3389 7624 3399 7651
rect 3428 7629 3510 7651
rect 3730 7685 3898 7686
rect 4138 7685 4176 7773
rect 4437 7771 4484 7773
rect 4784 7749 4824 7773
rect 3730 7662 4176 7685
rect 4402 7716 4513 7731
rect 4402 7714 4444 7716
rect 4402 7694 4409 7714
rect 4428 7694 4444 7714
rect 4402 7686 4444 7694
rect 4472 7714 4513 7716
rect 4472 7694 4486 7714
rect 4505 7694 4513 7714
rect 4785 7705 4824 7749
rect 4472 7686 4513 7694
rect 4402 7680 4513 7686
rect 3730 7659 4174 7662
rect 3730 7657 3898 7659
rect 3428 7624 3432 7629
rect 3389 7621 3432 7624
rect 3322 7607 3432 7621
rect 2112 7588 2280 7590
rect 1833 7581 2280 7588
rect 1497 7561 1608 7567
rect 1497 7553 1538 7561
rect 915 7540 951 7541
rect 763 7510 772 7530
rect 792 7510 800 7530
rect 651 7501 707 7503
rect 651 7500 688 7501
rect 763 7500 800 7510
rect 859 7530 1007 7540
rect 1107 7537 1203 7539
rect 859 7510 868 7530
rect 888 7510 978 7530
rect 998 7510 1007 7530
rect 859 7501 1007 7510
rect 1065 7530 1203 7537
rect 1065 7510 1074 7530
rect 1094 7510 1203 7530
rect 1497 7533 1505 7553
rect 1524 7533 1538 7553
rect 1497 7531 1538 7533
rect 1566 7553 1608 7561
rect 1566 7533 1582 7553
rect 1601 7533 1608 7553
rect 1833 7554 1858 7581
rect 1889 7562 2280 7581
rect 1889 7554 1938 7562
rect 2112 7561 2280 7562
rect 1833 7552 1938 7554
rect 1566 7531 1608 7533
rect 1497 7516 1608 7531
rect 1065 7501 1203 7510
rect 859 7500 896 7501
rect 915 7449 951 7501
rect 970 7500 1007 7501
rect 1066 7500 1103 7501
rect 386 7447 427 7448
rect 278 7440 427 7447
rect 278 7420 396 7440
rect 416 7420 427 7440
rect 278 7412 427 7420
rect 494 7444 853 7448
rect 494 7439 816 7444
rect 494 7415 607 7439
rect 631 7420 816 7439
rect 840 7420 853 7444
rect 631 7415 853 7420
rect 494 7412 853 7415
rect 915 7412 950 7449
rect 1018 7446 1118 7449
rect 1018 7442 1085 7446
rect 1018 7416 1030 7442
rect 1056 7420 1085 7442
rect 1111 7420 1118 7446
rect 1056 7416 1118 7420
rect 1018 7412 1118 7416
rect 494 7391 525 7412
rect 915 7391 951 7412
rect 337 7390 374 7391
rect 111 7387 145 7388
rect 110 7378 147 7387
rect 110 7360 119 7378
rect 137 7360 147 7378
rect 110 7350 147 7360
rect 336 7381 374 7390
rect 336 7361 345 7381
rect 365 7361 374 7381
rect 336 7353 374 7361
rect 440 7385 525 7391
rect 550 7390 587 7391
rect 440 7365 448 7385
rect 468 7365 525 7385
rect 440 7357 525 7365
rect 549 7381 587 7390
rect 549 7361 558 7381
rect 578 7361 587 7381
rect 440 7356 476 7357
rect 549 7353 587 7361
rect 653 7385 738 7391
rect 758 7390 795 7391
rect 653 7365 661 7385
rect 681 7384 738 7385
rect 681 7365 710 7384
rect 653 7364 710 7365
rect 731 7364 738 7384
rect 653 7357 738 7364
rect 757 7381 795 7390
rect 757 7361 766 7381
rect 786 7361 795 7381
rect 653 7356 689 7357
rect 757 7353 795 7361
rect 861 7385 1005 7391
rect 861 7365 869 7385
rect 889 7384 977 7385
rect 889 7365 920 7384
rect 861 7364 920 7365
rect 945 7365 977 7384
rect 997 7365 1005 7385
rect 945 7364 1005 7365
rect 861 7357 1005 7364
rect 861 7356 897 7357
rect 969 7356 1005 7357
rect 1071 7390 1108 7391
rect 1071 7389 1109 7390
rect 1071 7381 1135 7389
rect 1071 7361 1080 7381
rect 1100 7367 1135 7381
rect 1155 7367 1158 7387
rect 1100 7362 1158 7367
rect 1100 7361 1135 7362
rect 111 7322 145 7350
rect 337 7324 374 7353
rect 338 7322 374 7324
rect 550 7322 587 7353
rect 111 7321 283 7322
rect 111 7289 297 7321
rect 338 7300 587 7322
rect 758 7321 795 7353
rect 1071 7349 1135 7361
rect 1175 7323 1202 7501
rect 3730 7479 3757 7657
rect 3797 7619 3861 7631
rect 4137 7627 4174 7659
rect 4345 7658 4594 7680
rect 4345 7627 4382 7658
rect 4558 7656 4594 7658
rect 4558 7627 4595 7656
rect 3797 7618 3832 7619
rect 3774 7613 3832 7618
rect 3774 7593 3777 7613
rect 3797 7599 3832 7613
rect 3852 7599 3861 7619
rect 3797 7591 3861 7599
rect 3823 7590 3861 7591
rect 3824 7589 3861 7590
rect 3927 7623 3963 7624
rect 4035 7623 4071 7624
rect 3927 7618 4071 7623
rect 3927 7615 3989 7618
rect 3927 7595 3935 7615
rect 3955 7598 3989 7615
rect 4012 7615 4071 7618
rect 4012 7598 4043 7615
rect 3955 7595 4043 7598
rect 4063 7595 4071 7615
rect 3927 7589 4071 7595
rect 4137 7619 4175 7627
rect 4243 7623 4279 7624
rect 4137 7599 4146 7619
rect 4166 7599 4175 7619
rect 4137 7590 4175 7599
rect 4194 7616 4279 7623
rect 4194 7596 4201 7616
rect 4222 7615 4279 7616
rect 4222 7596 4251 7615
rect 4194 7595 4251 7596
rect 4271 7595 4279 7615
rect 4137 7589 4174 7590
rect 4194 7589 4279 7595
rect 4345 7619 4383 7627
rect 4456 7623 4492 7624
rect 4345 7599 4354 7619
rect 4374 7599 4383 7619
rect 4345 7590 4383 7599
rect 4407 7615 4492 7623
rect 4407 7595 4464 7615
rect 4484 7595 4492 7615
rect 4345 7589 4382 7590
rect 4407 7589 4492 7595
rect 4558 7619 4596 7627
rect 4558 7599 4567 7619
rect 4587 7599 4596 7619
rect 4558 7590 4596 7599
rect 4558 7589 4595 7590
rect 3981 7568 4017 7589
rect 4407 7568 4438 7589
rect 3814 7564 3914 7568
rect 3814 7560 3876 7564
rect 3814 7534 3821 7560
rect 3847 7538 3876 7560
rect 3902 7538 3914 7564
rect 3847 7534 3914 7538
rect 3814 7531 3914 7534
rect 3982 7531 4017 7568
rect 4079 7565 4438 7568
rect 4079 7560 4301 7565
rect 4079 7536 4092 7560
rect 4116 7541 4301 7560
rect 4325 7541 4438 7565
rect 4116 7536 4438 7541
rect 4079 7532 4438 7536
rect 4505 7560 4654 7568
rect 4505 7540 4516 7560
rect 4536 7540 4654 7560
rect 4505 7533 4654 7540
rect 4505 7532 4546 7533
rect 3829 7479 3866 7480
rect 3925 7479 3962 7480
rect 3981 7479 4017 7531
rect 4036 7479 4073 7480
rect 3729 7470 3867 7479
rect 3729 7450 3838 7470
rect 3858 7450 3867 7470
rect 3729 7443 3867 7450
rect 3925 7470 4073 7479
rect 3925 7450 3934 7470
rect 3954 7450 4044 7470
rect 4064 7450 4073 7470
rect 3729 7441 3825 7443
rect 3925 7440 4073 7450
rect 4132 7470 4169 7480
rect 4244 7479 4281 7480
rect 4225 7477 4281 7479
rect 4132 7450 4140 7470
rect 4160 7450 4169 7470
rect 3981 7439 4017 7440
rect 1358 7397 1468 7411
rect 1358 7394 1401 7397
rect 1358 7389 1362 7394
rect 1034 7321 1202 7323
rect 758 7315 1202 7321
rect 111 7257 145 7289
rect 107 7248 145 7257
rect 107 7230 117 7248
rect 135 7230 145 7248
rect 107 7224 145 7230
rect 263 7226 297 7289
rect 419 7294 530 7300
rect 419 7286 460 7294
rect 419 7266 427 7286
rect 446 7266 460 7286
rect 419 7264 460 7266
rect 488 7286 530 7294
rect 488 7266 504 7286
rect 523 7266 530 7286
rect 488 7264 530 7266
rect 419 7249 530 7264
rect 757 7295 1202 7315
rect 757 7226 795 7295
rect 1034 7294 1202 7295
rect 1280 7367 1362 7389
rect 1391 7367 1401 7394
rect 1429 7370 1436 7397
rect 1465 7389 1468 7397
rect 3463 7406 3574 7421
rect 3463 7404 3505 7406
rect 1465 7370 1530 7389
rect 1429 7367 1530 7370
rect 1280 7365 1530 7367
rect 1280 7286 1317 7365
rect 1358 7352 1468 7365
rect 1432 7296 1463 7297
rect 1280 7266 1289 7286
rect 1309 7266 1317 7286
rect 1280 7256 1317 7266
rect 1376 7286 1463 7296
rect 1376 7266 1385 7286
rect 1405 7266 1463 7286
rect 1376 7257 1463 7266
rect 1376 7256 1413 7257
rect 107 7220 144 7224
rect 263 7215 795 7226
rect 262 7199 795 7215
rect 1432 7204 1463 7257
rect 1493 7286 1530 7365
rect 1701 7375 2094 7382
rect 1701 7358 1709 7375
rect 1741 7362 2094 7375
rect 2114 7362 2117 7382
rect 3196 7377 3237 7386
rect 1741 7358 2117 7362
rect 1701 7357 2117 7358
rect 2791 7375 2959 7376
rect 3196 7375 3205 7377
rect 1701 7356 2042 7357
rect 1645 7296 1676 7297
rect 1493 7266 1502 7286
rect 1522 7266 1530 7286
rect 1493 7256 1530 7266
rect 1589 7289 1676 7296
rect 1589 7286 1650 7289
rect 1589 7266 1598 7286
rect 1618 7269 1650 7286
rect 1671 7269 1676 7289
rect 1618 7266 1676 7269
rect 1589 7259 1676 7266
rect 1701 7286 1738 7356
rect 2004 7355 2041 7356
rect 2791 7355 3205 7375
rect 3231 7355 3237 7377
rect 3463 7384 3470 7404
rect 3489 7384 3505 7404
rect 3463 7376 3505 7384
rect 3533 7404 3574 7406
rect 3533 7384 3547 7404
rect 3566 7384 3574 7404
rect 3533 7376 3574 7384
rect 3829 7380 3866 7381
rect 4132 7380 4169 7450
rect 4194 7470 4281 7477
rect 4194 7467 4252 7470
rect 4194 7447 4199 7467
rect 4220 7450 4252 7467
rect 4272 7450 4281 7470
rect 4220 7447 4281 7450
rect 4194 7440 4281 7447
rect 4340 7470 4377 7480
rect 4340 7450 4348 7470
rect 4368 7450 4377 7470
rect 4194 7439 4225 7440
rect 3828 7379 4169 7380
rect 3463 7370 3574 7376
rect 3753 7374 4169 7379
rect 2791 7349 3237 7355
rect 2791 7347 2959 7349
rect 1853 7296 1889 7297
rect 1701 7266 1710 7286
rect 1730 7266 1738 7286
rect 1589 7257 1645 7259
rect 1589 7256 1626 7257
rect 1701 7256 1738 7266
rect 1797 7286 1945 7296
rect 2045 7293 2141 7295
rect 1797 7266 1806 7286
rect 1826 7281 1916 7286
rect 1826 7266 1861 7281
rect 1797 7257 1861 7266
rect 1797 7256 1834 7257
rect 1853 7240 1861 7257
rect 1882 7266 1916 7281
rect 1936 7266 1945 7286
rect 1882 7257 1945 7266
rect 2003 7286 2141 7293
rect 2003 7266 2012 7286
rect 2032 7266 2141 7286
rect 2003 7257 2141 7266
rect 1882 7240 1889 7257
rect 1908 7256 1945 7257
rect 2004 7256 2041 7257
rect 1853 7205 1889 7240
rect 1324 7203 1365 7204
rect 262 7198 776 7199
rect 1216 7196 1365 7203
rect 1216 7176 1334 7196
rect 1354 7176 1365 7196
rect 1216 7168 1365 7176
rect 1432 7200 1791 7204
rect 1432 7195 1754 7200
rect 1432 7171 1545 7195
rect 1569 7176 1754 7195
rect 1778 7176 1791 7200
rect 1569 7171 1791 7176
rect 1432 7168 1791 7171
rect 1853 7168 1888 7205
rect 1956 7202 2056 7205
rect 1956 7198 2023 7202
rect 1956 7172 1968 7198
rect 1994 7176 2023 7198
rect 2049 7176 2056 7202
rect 1994 7172 2056 7176
rect 1956 7168 2056 7172
rect 110 7157 147 7158
rect 108 7149 148 7157
rect 108 7131 119 7149
rect 137 7131 148 7149
rect 1432 7147 1463 7168
rect 1853 7147 1889 7168
rect 1275 7146 1312 7147
rect 108 7083 148 7131
rect 1274 7137 1312 7146
rect 1274 7117 1283 7137
rect 1303 7117 1312 7137
rect 1274 7109 1312 7117
rect 1378 7141 1463 7147
rect 1488 7146 1525 7147
rect 1378 7121 1386 7141
rect 1406 7121 1463 7141
rect 1378 7113 1463 7121
rect 1487 7137 1525 7146
rect 1487 7117 1496 7137
rect 1516 7117 1525 7137
rect 1378 7112 1414 7113
rect 1487 7109 1525 7117
rect 1591 7141 1676 7147
rect 1696 7146 1733 7147
rect 1591 7121 1599 7141
rect 1619 7140 1676 7141
rect 1619 7121 1648 7140
rect 1591 7120 1648 7121
rect 1669 7120 1676 7140
rect 1591 7113 1676 7120
rect 1695 7137 1733 7146
rect 1695 7117 1704 7137
rect 1724 7117 1733 7137
rect 1591 7112 1627 7113
rect 1695 7109 1733 7117
rect 1799 7141 1943 7147
rect 1799 7121 1807 7141
rect 1827 7121 1915 7141
rect 1935 7121 1943 7141
rect 1799 7113 1943 7121
rect 1799 7112 1835 7113
rect 1907 7112 1943 7113
rect 2009 7146 2046 7147
rect 2009 7145 2047 7146
rect 2009 7137 2073 7145
rect 2009 7117 2018 7137
rect 2038 7123 2073 7137
rect 2093 7123 2096 7143
rect 2038 7118 2096 7123
rect 2038 7117 2073 7118
rect 419 7087 529 7101
rect 419 7084 462 7087
rect 108 7076 233 7083
rect 419 7079 423 7084
rect 108 7057 200 7076
rect 225 7057 233 7076
rect 108 7047 233 7057
rect 341 7057 423 7079
rect 452 7057 462 7084
rect 490 7060 497 7087
rect 526 7079 529 7087
rect 1275 7080 1312 7109
rect 526 7060 591 7079
rect 1276 7078 1312 7080
rect 1488 7078 1525 7109
rect 1696 7082 1733 7109
rect 2009 7105 2073 7117
rect 490 7057 591 7060
rect 341 7055 591 7057
rect 108 7027 148 7047
rect 107 7018 148 7027
rect 107 7000 117 7018
rect 135 7000 148 7018
rect 107 6991 148 7000
rect 107 6990 144 6991
rect 341 6976 378 7055
rect 419 7042 529 7055
rect 493 6986 524 6987
rect 341 6956 350 6976
rect 370 6956 378 6976
rect 341 6946 378 6956
rect 437 6976 524 6986
rect 437 6956 446 6976
rect 466 6956 524 6976
rect 437 6947 524 6956
rect 437 6946 474 6947
rect 110 6924 147 6928
rect 107 6919 147 6924
rect 107 6901 119 6919
rect 137 6901 147 6919
rect 107 6721 147 6901
rect 493 6894 524 6947
rect 554 6976 591 7055
rect 762 7052 1155 7072
rect 1175 7052 1178 7072
rect 1276 7056 1525 7078
rect 1694 7077 1735 7082
rect 2113 7079 2140 7257
rect 2791 7169 2818 7347
rect 3196 7344 3237 7349
rect 3406 7348 3655 7370
rect 3753 7354 3756 7374
rect 3776 7354 4169 7374
rect 4340 7371 4377 7450
rect 4407 7479 4438 7532
rect 4784 7525 4824 7705
rect 4784 7507 4794 7525
rect 4812 7507 4824 7525
rect 4784 7502 4824 7507
rect 4784 7498 4821 7502
rect 4457 7479 4494 7480
rect 4407 7470 4494 7479
rect 4407 7450 4465 7470
rect 4485 7450 4494 7470
rect 4407 7440 4494 7450
rect 4553 7470 4590 7480
rect 4553 7450 4561 7470
rect 4581 7450 4590 7470
rect 4407 7439 4438 7440
rect 4402 7371 4512 7384
rect 4553 7371 4590 7450
rect 4787 7435 4824 7436
rect 4783 7426 4824 7435
rect 4783 7408 4796 7426
rect 4814 7408 4824 7426
rect 4783 7399 4824 7408
rect 4783 7379 4823 7399
rect 4340 7369 4590 7371
rect 4340 7366 4441 7369
rect 2858 7309 2922 7321
rect 3198 7317 3235 7344
rect 3406 7317 3443 7348
rect 3619 7346 3655 7348
rect 4340 7347 4405 7366
rect 3619 7317 3656 7346
rect 4402 7339 4405 7347
rect 4434 7339 4441 7366
rect 4469 7342 4479 7369
rect 4508 7347 4590 7369
rect 4698 7369 4823 7379
rect 4698 7350 4706 7369
rect 4731 7350 4823 7369
rect 4508 7342 4512 7347
rect 4698 7343 4823 7350
rect 4469 7339 4512 7342
rect 4402 7325 4512 7339
rect 2858 7308 2893 7309
rect 2835 7303 2893 7308
rect 2835 7283 2838 7303
rect 2858 7289 2893 7303
rect 2913 7289 2922 7309
rect 2858 7281 2922 7289
rect 2884 7280 2922 7281
rect 2885 7279 2922 7280
rect 2988 7313 3024 7314
rect 3096 7313 3132 7314
rect 2988 7305 3132 7313
rect 2988 7285 2996 7305
rect 3016 7302 3104 7305
rect 3016 7285 3048 7302
rect 3068 7285 3104 7302
rect 3124 7285 3132 7305
rect 2988 7279 3132 7285
rect 3198 7309 3236 7317
rect 3304 7313 3340 7314
rect 3198 7289 3207 7309
rect 3227 7289 3236 7309
rect 3198 7280 3236 7289
rect 3255 7306 3340 7313
rect 3255 7286 3262 7306
rect 3283 7305 3340 7306
rect 3283 7286 3312 7305
rect 3255 7285 3312 7286
rect 3332 7285 3340 7305
rect 3198 7279 3235 7280
rect 3255 7279 3340 7285
rect 3406 7309 3444 7317
rect 3517 7313 3553 7314
rect 3406 7289 3415 7309
rect 3435 7289 3444 7309
rect 3406 7280 3444 7289
rect 3468 7305 3553 7313
rect 3468 7285 3525 7305
rect 3545 7285 3553 7305
rect 3406 7279 3443 7280
rect 3468 7279 3553 7285
rect 3619 7309 3657 7317
rect 3619 7289 3628 7309
rect 3648 7289 3657 7309
rect 3619 7280 3657 7289
rect 4783 7295 4823 7343
rect 3619 7279 3656 7280
rect 3042 7258 3078 7279
rect 3468 7258 3499 7279
rect 4783 7277 4794 7295
rect 4812 7277 4823 7295
rect 4783 7269 4823 7277
rect 4784 7268 4821 7269
rect 2875 7254 2975 7258
rect 2875 7250 2937 7254
rect 2875 7224 2882 7250
rect 2908 7228 2937 7250
rect 2963 7228 2975 7254
rect 2908 7224 2975 7228
rect 2875 7221 2975 7224
rect 3043 7221 3078 7258
rect 3140 7255 3499 7258
rect 3140 7250 3362 7255
rect 3140 7226 3153 7250
rect 3177 7231 3362 7250
rect 3386 7231 3499 7255
rect 3177 7226 3499 7231
rect 3140 7222 3499 7226
rect 3566 7250 3715 7258
rect 3566 7230 3577 7250
rect 3597 7230 3715 7250
rect 3566 7223 3715 7230
rect 4155 7227 4669 7228
rect 3566 7222 3607 7223
rect 2890 7169 2927 7170
rect 2986 7169 3023 7170
rect 3042 7169 3078 7221
rect 3097 7169 3134 7170
rect 2790 7160 2928 7169
rect 2790 7140 2899 7160
rect 2919 7140 2928 7160
rect 2790 7133 2928 7140
rect 2986 7160 3134 7169
rect 2986 7140 2995 7160
rect 3015 7140 3105 7160
rect 3125 7140 3134 7160
rect 2790 7131 2886 7133
rect 2986 7130 3134 7140
rect 3193 7160 3230 7170
rect 3305 7169 3342 7170
rect 3286 7167 3342 7169
rect 3193 7140 3201 7160
rect 3221 7140 3230 7160
rect 3042 7129 3078 7130
rect 1972 7077 2140 7079
rect 1694 7071 2140 7077
rect 762 7047 1178 7052
rect 1357 7050 1468 7056
rect 762 7046 1103 7047
rect 706 6986 737 6987
rect 554 6956 563 6976
rect 583 6956 591 6976
rect 554 6946 591 6956
rect 650 6979 737 6986
rect 650 6976 711 6979
rect 650 6956 659 6976
rect 679 6959 711 6976
rect 732 6959 737 6979
rect 679 6956 737 6959
rect 650 6949 737 6956
rect 762 6976 799 7046
rect 1065 7045 1102 7046
rect 1357 7042 1398 7050
rect 1357 7022 1365 7042
rect 1384 7022 1398 7042
rect 1357 7020 1398 7022
rect 1426 7042 1468 7050
rect 1426 7022 1442 7042
rect 1461 7022 1468 7042
rect 1694 7049 1700 7071
rect 1726 7051 2140 7071
rect 2890 7070 2927 7071
rect 3193 7070 3230 7140
rect 3255 7160 3342 7167
rect 3255 7157 3313 7160
rect 3255 7137 3260 7157
rect 3281 7140 3313 7157
rect 3333 7140 3342 7160
rect 3281 7137 3342 7140
rect 3255 7130 3342 7137
rect 3401 7160 3438 7170
rect 3401 7140 3409 7160
rect 3429 7140 3438 7160
rect 3255 7129 3286 7130
rect 2889 7069 3230 7070
rect 1726 7049 1735 7051
rect 1972 7050 2140 7051
rect 2814 7064 3230 7069
rect 1694 7040 1735 7049
rect 2814 7044 2817 7064
rect 2837 7044 3230 7064
rect 3401 7061 3438 7140
rect 3468 7169 3499 7222
rect 4136 7211 4669 7227
rect 4136 7200 4668 7211
rect 4787 7202 4824 7206
rect 3518 7169 3555 7170
rect 3468 7160 3555 7169
rect 3468 7140 3526 7160
rect 3546 7140 3555 7160
rect 3468 7130 3555 7140
rect 3614 7160 3651 7170
rect 3614 7140 3622 7160
rect 3642 7140 3651 7160
rect 3468 7129 3499 7130
rect 3463 7061 3573 7074
rect 3614 7061 3651 7140
rect 3401 7059 3651 7061
rect 3401 7056 3502 7059
rect 3401 7037 3466 7056
rect 1426 7020 1468 7022
rect 1357 7005 1468 7020
rect 3463 7029 3466 7037
rect 3495 7029 3502 7056
rect 3530 7032 3540 7059
rect 3569 7037 3651 7059
rect 3729 7131 3897 7132
rect 4136 7131 4174 7200
rect 3729 7111 4174 7131
rect 4401 7162 4512 7177
rect 4401 7160 4443 7162
rect 4401 7140 4408 7160
rect 4427 7140 4443 7160
rect 4401 7132 4443 7140
rect 4471 7160 4512 7162
rect 4471 7140 4485 7160
rect 4504 7140 4512 7160
rect 4471 7132 4512 7140
rect 4401 7126 4512 7132
rect 4634 7137 4668 7200
rect 4786 7196 4824 7202
rect 4786 7178 4796 7196
rect 4814 7178 4824 7196
rect 4786 7169 4824 7178
rect 4786 7137 4820 7169
rect 3729 7105 4173 7111
rect 3729 7103 3897 7105
rect 3569 7032 3573 7037
rect 3530 7029 3573 7032
rect 3463 7015 3573 7029
rect 914 6986 950 6987
rect 762 6956 771 6976
rect 791 6956 799 6976
rect 650 6947 706 6949
rect 650 6946 687 6947
rect 762 6946 799 6956
rect 858 6976 1006 6986
rect 1106 6983 1202 6985
rect 858 6956 867 6976
rect 887 6956 977 6976
rect 997 6956 1006 6976
rect 858 6947 1006 6956
rect 1064 6976 1202 6983
rect 1064 6956 1073 6976
rect 1093 6956 1202 6976
rect 1064 6947 1202 6956
rect 858 6946 895 6947
rect 914 6895 950 6947
rect 969 6946 1006 6947
rect 1065 6946 1102 6947
rect 385 6893 426 6894
rect 277 6886 426 6893
rect 277 6866 395 6886
rect 415 6866 426 6886
rect 277 6858 426 6866
rect 493 6890 852 6894
rect 493 6885 815 6890
rect 493 6861 606 6885
rect 630 6866 815 6885
rect 839 6866 852 6890
rect 630 6861 852 6866
rect 493 6858 852 6861
rect 914 6858 949 6895
rect 1017 6892 1117 6895
rect 1017 6888 1084 6892
rect 1017 6862 1029 6888
rect 1055 6866 1084 6888
rect 1110 6866 1117 6892
rect 1055 6862 1117 6866
rect 1017 6858 1117 6862
rect 493 6837 524 6858
rect 914 6837 950 6858
rect 336 6836 373 6837
rect 335 6827 373 6836
rect 335 6807 344 6827
rect 364 6807 373 6827
rect 335 6799 373 6807
rect 439 6831 524 6837
rect 549 6836 586 6837
rect 439 6811 447 6831
rect 467 6811 524 6831
rect 439 6803 524 6811
rect 548 6827 586 6836
rect 548 6807 557 6827
rect 577 6807 586 6827
rect 439 6802 475 6803
rect 548 6799 586 6807
rect 652 6831 737 6837
rect 757 6836 794 6837
rect 652 6811 660 6831
rect 680 6830 737 6831
rect 680 6811 709 6830
rect 652 6810 709 6811
rect 730 6810 737 6830
rect 652 6803 737 6810
rect 756 6827 794 6836
rect 756 6807 765 6827
rect 785 6807 794 6827
rect 652 6802 688 6803
rect 756 6799 794 6807
rect 860 6831 1004 6837
rect 860 6811 868 6831
rect 888 6828 976 6831
rect 888 6811 919 6828
rect 860 6808 919 6811
rect 942 6811 976 6828
rect 996 6811 1004 6831
rect 942 6808 1004 6811
rect 860 6803 1004 6808
rect 860 6802 896 6803
rect 968 6802 1004 6803
rect 1070 6836 1107 6837
rect 1070 6835 1108 6836
rect 1070 6827 1134 6835
rect 1070 6807 1079 6827
rect 1099 6813 1134 6827
rect 1154 6813 1157 6833
rect 1099 6808 1157 6813
rect 1099 6807 1134 6808
rect 336 6770 373 6799
rect 337 6768 373 6770
rect 549 6768 586 6799
rect 337 6746 586 6768
rect 757 6767 794 6799
rect 1070 6795 1134 6807
rect 1174 6769 1201 6947
rect 3729 6925 3756 7103
rect 3796 7065 3860 7077
rect 4136 7073 4173 7105
rect 4344 7104 4593 7126
rect 4634 7105 4820 7137
rect 4648 7104 4820 7105
rect 4344 7073 4381 7104
rect 4557 7102 4593 7104
rect 4557 7073 4594 7102
rect 4786 7076 4820 7104
rect 3796 7064 3831 7065
rect 3773 7059 3831 7064
rect 3773 7039 3776 7059
rect 3796 7045 3831 7059
rect 3851 7045 3860 7065
rect 3796 7037 3860 7045
rect 3822 7036 3860 7037
rect 3823 7035 3860 7036
rect 3926 7069 3962 7070
rect 4034 7069 4070 7070
rect 3926 7062 4070 7069
rect 3926 7061 3986 7062
rect 3926 7041 3934 7061
rect 3954 7042 3986 7061
rect 4011 7061 4070 7062
rect 4011 7042 4042 7061
rect 3954 7041 4042 7042
rect 4062 7041 4070 7061
rect 3926 7035 4070 7041
rect 4136 7065 4174 7073
rect 4242 7069 4278 7070
rect 4136 7045 4145 7065
rect 4165 7045 4174 7065
rect 4136 7036 4174 7045
rect 4193 7062 4278 7069
rect 4193 7042 4200 7062
rect 4221 7061 4278 7062
rect 4221 7042 4250 7061
rect 4193 7041 4250 7042
rect 4270 7041 4278 7061
rect 4136 7035 4173 7036
rect 4193 7035 4278 7041
rect 4344 7065 4382 7073
rect 4455 7069 4491 7070
rect 4344 7045 4353 7065
rect 4373 7045 4382 7065
rect 4344 7036 4382 7045
rect 4406 7061 4491 7069
rect 4406 7041 4463 7061
rect 4483 7041 4491 7061
rect 4344 7035 4381 7036
rect 4406 7035 4491 7041
rect 4557 7065 4595 7073
rect 4557 7045 4566 7065
rect 4586 7045 4595 7065
rect 4557 7036 4595 7045
rect 4784 7066 4821 7076
rect 4784 7048 4794 7066
rect 4812 7048 4821 7066
rect 4784 7039 4821 7048
rect 4786 7038 4820 7039
rect 4557 7035 4594 7036
rect 3980 7014 4016 7035
rect 4406 7014 4437 7035
rect 3813 7010 3913 7014
rect 3813 7006 3875 7010
rect 3813 6980 3820 7006
rect 3846 6984 3875 7006
rect 3901 6984 3913 7010
rect 3846 6980 3913 6984
rect 3813 6977 3913 6980
rect 3981 6977 4016 7014
rect 4078 7011 4437 7014
rect 4078 7006 4300 7011
rect 4078 6982 4091 7006
rect 4115 6987 4300 7006
rect 4324 6987 4437 7011
rect 4115 6982 4437 6987
rect 4078 6978 4437 6982
rect 4504 7006 4653 7014
rect 4504 6986 4515 7006
rect 4535 6986 4653 7006
rect 4504 6979 4653 6986
rect 4504 6978 4545 6979
rect 3828 6925 3865 6926
rect 3924 6925 3961 6926
rect 3980 6925 4016 6977
rect 4035 6925 4072 6926
rect 3728 6916 3866 6925
rect 3353 6882 3464 6897
rect 3728 6896 3837 6916
rect 3857 6896 3866 6916
rect 3728 6889 3866 6896
rect 3924 6916 4072 6925
rect 3924 6896 3933 6916
rect 3953 6896 4043 6916
rect 4063 6896 4072 6916
rect 3728 6887 3824 6889
rect 3924 6886 4072 6896
rect 4131 6916 4168 6926
rect 4243 6925 4280 6926
rect 4224 6923 4280 6925
rect 4131 6896 4139 6916
rect 4159 6896 4168 6916
rect 3980 6885 4016 6886
rect 3353 6880 3395 6882
rect 2690 6861 2760 6870
rect 2690 6852 2707 6861
rect 2681 6832 2707 6852
rect 2755 6852 2760 6861
rect 3353 6860 3360 6880
rect 3379 6860 3395 6880
rect 3353 6852 3395 6860
rect 3423 6880 3464 6882
rect 3423 6860 3437 6880
rect 3456 6860 3464 6880
rect 3423 6852 3464 6860
rect 2755 6851 2849 6852
rect 2755 6832 3125 6851
rect 3353 6846 3464 6852
rect 1468 6818 1578 6832
rect 1468 6815 1511 6818
rect 1468 6810 1472 6815
rect 1033 6767 1201 6769
rect 757 6764 1201 6767
rect 418 6740 529 6746
rect 418 6732 459 6740
rect 107 6677 146 6721
rect 418 6712 426 6732
rect 445 6712 459 6732
rect 418 6710 459 6712
rect 487 6732 529 6740
rect 487 6712 503 6732
rect 522 6712 529 6732
rect 487 6710 529 6712
rect 418 6696 529 6710
rect 755 6741 1201 6764
rect 107 6653 147 6677
rect 447 6653 494 6655
rect 755 6653 793 6741
rect 1033 6740 1201 6741
rect 1390 6788 1472 6810
rect 1501 6788 1511 6815
rect 1539 6791 1546 6818
rect 1575 6810 1578 6818
rect 2681 6825 3125 6832
rect 2681 6823 2849 6825
rect 2681 6815 2760 6823
rect 1575 6791 1640 6810
rect 1539 6788 1640 6791
rect 1390 6786 1640 6788
rect 1390 6707 1427 6786
rect 1468 6773 1578 6786
rect 1542 6717 1573 6718
rect 1390 6687 1399 6707
rect 1419 6687 1427 6707
rect 1390 6677 1427 6687
rect 1486 6707 1573 6717
rect 1486 6687 1495 6707
rect 1515 6687 1573 6707
rect 1486 6678 1573 6687
rect 1486 6677 1523 6678
rect 107 6620 793 6653
rect 1542 6625 1573 6678
rect 1603 6707 1640 6786
rect 1811 6783 2204 6803
rect 2224 6783 2227 6803
rect 1811 6778 2227 6783
rect 1811 6777 2152 6778
rect 1755 6717 1786 6718
rect 1603 6687 1612 6707
rect 1632 6687 1640 6707
rect 1603 6677 1640 6687
rect 1699 6710 1786 6717
rect 1699 6707 1760 6710
rect 1699 6687 1708 6707
rect 1728 6690 1760 6707
rect 1781 6690 1786 6710
rect 1728 6687 1786 6690
rect 1699 6680 1786 6687
rect 1811 6707 1848 6777
rect 2114 6776 2151 6777
rect 1963 6717 1999 6718
rect 1811 6687 1820 6707
rect 1840 6687 1848 6707
rect 1699 6678 1755 6680
rect 1699 6677 1736 6678
rect 1811 6677 1848 6687
rect 1907 6707 2055 6717
rect 2155 6714 2251 6716
rect 1907 6687 1916 6707
rect 1936 6687 2026 6707
rect 2046 6687 2055 6707
rect 1907 6678 2055 6687
rect 2113 6707 2251 6714
rect 2113 6687 2122 6707
rect 2142 6687 2251 6707
rect 2113 6678 2251 6687
rect 1907 6677 1944 6678
rect 1963 6626 1999 6678
rect 2018 6677 2055 6678
rect 2114 6677 2151 6678
rect 1434 6624 1475 6625
rect 106 6563 145 6620
rect 755 6618 793 6620
rect 1326 6617 1475 6624
rect 1326 6597 1444 6617
rect 1464 6597 1475 6617
rect 1326 6589 1475 6597
rect 1542 6621 1901 6625
rect 1542 6616 1864 6621
rect 1542 6592 1655 6616
rect 1679 6597 1864 6616
rect 1888 6597 1901 6621
rect 1679 6592 1901 6597
rect 1542 6589 1901 6592
rect 1963 6589 1998 6626
rect 2066 6623 2166 6626
rect 2066 6619 2133 6623
rect 2066 6593 2078 6619
rect 2104 6597 2133 6619
rect 2159 6597 2166 6623
rect 2104 6593 2166 6597
rect 2066 6589 2166 6593
rect 1542 6568 1573 6589
rect 1963 6568 1999 6589
rect 1385 6567 1422 6568
rect 106 6561 154 6563
rect 106 6543 117 6561
rect 135 6543 154 6561
rect 1384 6558 1422 6567
rect 106 6534 154 6543
rect 107 6533 154 6534
rect 420 6538 530 6552
rect 420 6535 463 6538
rect 420 6530 424 6535
rect 342 6508 424 6530
rect 453 6508 463 6535
rect 491 6511 498 6538
rect 527 6530 530 6538
rect 1384 6538 1393 6558
rect 1413 6538 1422 6558
rect 1384 6530 1422 6538
rect 1488 6562 1573 6568
rect 1598 6567 1635 6568
rect 1488 6542 1496 6562
rect 1516 6542 1573 6562
rect 1488 6534 1573 6542
rect 1597 6558 1635 6567
rect 1597 6538 1606 6558
rect 1626 6538 1635 6558
rect 1488 6533 1524 6534
rect 1597 6530 1635 6538
rect 1701 6562 1786 6568
rect 1806 6567 1843 6568
rect 1701 6542 1709 6562
rect 1729 6561 1786 6562
rect 1729 6542 1758 6561
rect 1701 6541 1758 6542
rect 1779 6541 1786 6561
rect 1701 6534 1786 6541
rect 1805 6558 1843 6567
rect 1805 6538 1814 6558
rect 1834 6538 1843 6558
rect 1701 6533 1737 6534
rect 1805 6530 1843 6538
rect 1909 6562 2053 6568
rect 1909 6542 1917 6562
rect 1937 6560 2025 6562
rect 1937 6542 1966 6560
rect 1909 6541 1966 6542
rect 1995 6542 2025 6560
rect 2045 6542 2053 6562
rect 1995 6541 2053 6542
rect 1909 6534 2053 6541
rect 1909 6533 1945 6534
rect 2017 6533 2053 6534
rect 2119 6567 2156 6568
rect 2119 6566 2157 6567
rect 2119 6558 2183 6566
rect 2119 6538 2128 6558
rect 2148 6544 2183 6558
rect 2203 6544 2206 6564
rect 2148 6539 2206 6544
rect 2148 6538 2183 6539
rect 527 6511 592 6530
rect 491 6508 592 6511
rect 342 6506 592 6508
rect 110 6470 147 6471
rect 106 6467 147 6470
rect 106 6462 148 6467
rect 106 6444 119 6462
rect 137 6444 148 6462
rect 106 6430 148 6444
rect 186 6430 233 6434
rect 106 6424 233 6430
rect 106 6395 194 6424
rect 223 6395 233 6424
rect 342 6427 379 6506
rect 420 6493 530 6506
rect 494 6437 525 6438
rect 342 6407 351 6427
rect 371 6407 379 6427
rect 342 6397 379 6407
rect 438 6427 525 6437
rect 438 6407 447 6427
rect 467 6407 525 6427
rect 438 6398 525 6407
rect 438 6397 475 6398
rect 106 6391 233 6395
rect 106 6374 145 6391
rect 186 6390 233 6391
rect 106 6356 117 6374
rect 135 6356 145 6374
rect 106 6347 145 6356
rect 107 6346 144 6347
rect 494 6345 525 6398
rect 555 6427 592 6506
rect 763 6503 1156 6523
rect 1176 6503 1179 6523
rect 763 6498 1179 6503
rect 1385 6501 1422 6530
rect 1386 6499 1422 6501
rect 1598 6499 1635 6530
rect 763 6497 1104 6498
rect 707 6437 738 6438
rect 555 6407 564 6427
rect 584 6407 592 6427
rect 555 6397 592 6407
rect 651 6430 738 6437
rect 651 6427 712 6430
rect 651 6407 660 6427
rect 680 6410 712 6427
rect 733 6410 738 6430
rect 680 6407 738 6410
rect 651 6400 738 6407
rect 763 6427 800 6497
rect 1066 6496 1103 6497
rect 1386 6477 1635 6499
rect 1806 6498 1843 6530
rect 2119 6526 2183 6538
rect 2223 6502 2250 6678
rect 2681 6645 2708 6815
rect 2748 6785 2812 6797
rect 3088 6793 3125 6825
rect 3296 6824 3545 6846
rect 3828 6826 3865 6827
rect 4131 6826 4168 6896
rect 4193 6916 4280 6923
rect 4193 6913 4251 6916
rect 4193 6893 4198 6913
rect 4219 6896 4251 6913
rect 4271 6896 4280 6916
rect 4219 6893 4280 6896
rect 4193 6886 4280 6893
rect 4339 6916 4376 6926
rect 4339 6896 4347 6916
rect 4367 6896 4376 6916
rect 4193 6885 4224 6886
rect 3827 6825 4168 6826
rect 3296 6793 3333 6824
rect 3509 6822 3545 6824
rect 3509 6793 3546 6822
rect 3752 6820 4168 6825
rect 3752 6800 3755 6820
rect 3775 6800 4168 6820
rect 4339 6817 4376 6896
rect 4406 6925 4437 6978
rect 4787 6976 4824 6977
rect 4786 6967 4825 6976
rect 4786 6949 4796 6967
rect 4814 6949 4825 6967
rect 4698 6932 4745 6933
rect 4786 6932 4825 6949
rect 4698 6928 4825 6932
rect 4456 6925 4493 6926
rect 4406 6916 4493 6925
rect 4406 6896 4464 6916
rect 4484 6896 4493 6916
rect 4406 6886 4493 6896
rect 4552 6916 4589 6926
rect 4552 6896 4560 6916
rect 4580 6896 4589 6916
rect 4406 6885 4437 6886
rect 4401 6817 4511 6830
rect 4552 6817 4589 6896
rect 4698 6899 4708 6928
rect 4737 6899 4825 6928
rect 4698 6893 4825 6899
rect 4698 6889 4745 6893
rect 4783 6879 4825 6893
rect 4783 6861 4794 6879
rect 4812 6861 4825 6879
rect 4783 6856 4825 6861
rect 4784 6853 4825 6856
rect 4784 6852 4821 6853
rect 4339 6815 4589 6817
rect 4339 6812 4440 6815
rect 4339 6793 4404 6812
rect 2748 6784 2783 6785
rect 2725 6779 2783 6784
rect 2725 6759 2728 6779
rect 2748 6765 2783 6779
rect 2803 6765 2812 6785
rect 2748 6757 2812 6765
rect 2774 6756 2812 6757
rect 2775 6755 2812 6756
rect 2878 6789 2914 6790
rect 2986 6789 3022 6790
rect 2878 6781 3022 6789
rect 2878 6761 2886 6781
rect 2906 6761 2994 6781
rect 3014 6761 3022 6781
rect 2878 6755 3022 6761
rect 3088 6785 3126 6793
rect 3194 6789 3230 6790
rect 3088 6765 3097 6785
rect 3117 6765 3126 6785
rect 3088 6756 3126 6765
rect 3145 6782 3230 6789
rect 3145 6762 3152 6782
rect 3173 6781 3230 6782
rect 3173 6762 3202 6781
rect 3145 6761 3202 6762
rect 3222 6761 3230 6781
rect 3088 6755 3125 6756
rect 3145 6755 3230 6761
rect 3296 6785 3334 6793
rect 3407 6789 3443 6790
rect 3296 6765 3305 6785
rect 3325 6765 3334 6785
rect 3296 6756 3334 6765
rect 3358 6781 3443 6789
rect 3358 6761 3415 6781
rect 3435 6761 3443 6781
rect 3296 6755 3333 6756
rect 3358 6755 3443 6761
rect 3509 6785 3547 6793
rect 3509 6765 3518 6785
rect 3538 6765 3547 6785
rect 4401 6785 4404 6793
rect 4433 6785 4440 6812
rect 4468 6788 4478 6815
rect 4507 6793 4589 6815
rect 4507 6788 4511 6793
rect 4468 6785 4511 6788
rect 4401 6771 4511 6785
rect 4777 6789 4824 6790
rect 4777 6780 4825 6789
rect 3509 6756 3547 6765
rect 4777 6762 4796 6780
rect 4814 6762 4825 6780
rect 4777 6760 4825 6762
rect 3509 6755 3546 6756
rect 2932 6734 2968 6755
rect 3358 6734 3389 6755
rect 2765 6730 2865 6734
rect 2765 6726 2827 6730
rect 2765 6700 2772 6726
rect 2798 6704 2827 6726
rect 2853 6704 2865 6730
rect 2798 6700 2865 6704
rect 2765 6697 2865 6700
rect 2933 6697 2968 6734
rect 3030 6731 3389 6734
rect 3030 6726 3252 6731
rect 3030 6702 3043 6726
rect 3067 6707 3252 6726
rect 3276 6707 3389 6731
rect 3067 6702 3389 6707
rect 3030 6698 3389 6702
rect 3456 6726 3605 6734
rect 3456 6706 3467 6726
rect 3487 6706 3605 6726
rect 3456 6699 3605 6706
rect 4138 6703 4176 6705
rect 4786 6703 4825 6760
rect 3456 6698 3497 6699
rect 2932 6657 2968 6697
rect 2780 6645 2817 6646
rect 2876 6645 2913 6646
rect 2932 6645 2937 6657
rect 2680 6636 2818 6645
rect 2680 6616 2789 6636
rect 2809 6616 2818 6636
rect 2680 6609 2818 6616
rect 2876 6636 2937 6645
rect 2876 6616 2885 6636
rect 2905 6625 2937 6636
rect 2964 6645 2968 6657
rect 2987 6645 3024 6646
rect 2964 6636 3024 6645
rect 2964 6625 2995 6636
rect 2905 6616 2995 6625
rect 3015 6616 3024 6636
rect 2680 6607 2776 6609
rect 2876 6606 3024 6616
rect 3083 6636 3120 6646
rect 3195 6645 3232 6646
rect 3176 6643 3232 6645
rect 3083 6616 3091 6636
rect 3111 6616 3120 6636
rect 2932 6605 2968 6606
rect 2780 6546 2817 6547
rect 3083 6546 3120 6616
rect 3145 6636 3232 6643
rect 3145 6633 3203 6636
rect 3145 6613 3150 6633
rect 3171 6616 3203 6633
rect 3223 6616 3232 6636
rect 3171 6613 3232 6616
rect 3145 6606 3232 6613
rect 3291 6636 3328 6646
rect 3291 6616 3299 6636
rect 3319 6616 3328 6636
rect 3145 6605 3176 6606
rect 2779 6545 3120 6546
rect 2704 6540 3120 6545
rect 2704 6522 2707 6540
rect 2727 6538 3120 6540
rect 2727 6522 3097 6538
rect 2745 6520 3097 6522
rect 3088 6518 3097 6520
rect 3118 6518 3120 6538
rect 3088 6506 3120 6518
rect 3291 6537 3328 6616
rect 3358 6645 3389 6698
rect 4138 6670 4824 6703
rect 3408 6645 3445 6646
rect 3358 6636 3445 6645
rect 3358 6616 3416 6636
rect 3436 6616 3445 6636
rect 3358 6606 3445 6616
rect 3504 6636 3541 6646
rect 3504 6616 3512 6636
rect 3532 6616 3541 6636
rect 3358 6605 3389 6606
rect 3353 6537 3463 6550
rect 3504 6537 3541 6616
rect 3291 6535 3541 6537
rect 3291 6532 3392 6535
rect 3291 6513 3356 6532
rect 2131 6500 2250 6502
rect 2082 6498 2250 6500
rect 1467 6471 1578 6477
rect 1806 6472 2250 6498
rect 3353 6505 3356 6513
rect 3385 6505 3392 6532
rect 3420 6508 3430 6535
rect 3459 6513 3541 6535
rect 3730 6582 3898 6583
rect 4138 6582 4176 6670
rect 4437 6668 4484 6670
rect 4784 6646 4824 6670
rect 3730 6559 4176 6582
rect 4402 6613 4513 6627
rect 4402 6611 4444 6613
rect 4402 6591 4409 6611
rect 4428 6591 4444 6611
rect 4402 6583 4444 6591
rect 4472 6611 4513 6613
rect 4472 6591 4486 6611
rect 4505 6591 4513 6611
rect 4785 6602 4824 6646
rect 4472 6583 4513 6591
rect 4402 6577 4513 6583
rect 3730 6556 4174 6559
rect 3730 6554 3898 6556
rect 3459 6508 3463 6513
rect 3420 6505 3463 6508
rect 3353 6491 3463 6505
rect 2082 6471 2250 6472
rect 1467 6463 1508 6471
rect 1467 6443 1475 6463
rect 1494 6443 1508 6463
rect 1467 6441 1508 6443
rect 1536 6463 1578 6471
rect 2131 6470 2239 6471
rect 1536 6443 1552 6463
rect 1571 6443 1578 6463
rect 1536 6441 1578 6443
rect 915 6437 951 6438
rect 763 6407 772 6427
rect 792 6407 800 6427
rect 651 6398 707 6400
rect 651 6397 688 6398
rect 763 6397 800 6407
rect 859 6427 1007 6437
rect 1107 6434 1203 6436
rect 859 6407 868 6427
rect 888 6407 978 6427
rect 998 6407 1007 6427
rect 859 6398 1007 6407
rect 1065 6427 1203 6434
rect 1065 6407 1074 6427
rect 1094 6407 1203 6427
rect 1467 6426 1578 6441
rect 2169 6469 2239 6470
rect 1065 6398 1203 6407
rect 859 6397 896 6398
rect 915 6346 951 6398
rect 970 6397 1007 6398
rect 1066 6397 1103 6398
rect 386 6344 427 6345
rect 278 6337 427 6344
rect 278 6317 396 6337
rect 416 6317 427 6337
rect 278 6309 427 6317
rect 494 6341 853 6345
rect 494 6336 816 6341
rect 494 6312 607 6336
rect 631 6317 816 6336
rect 840 6317 853 6341
rect 631 6312 853 6317
rect 494 6309 853 6312
rect 915 6309 950 6346
rect 1018 6343 1118 6346
rect 1018 6339 1085 6343
rect 1018 6313 1030 6339
rect 1056 6317 1085 6339
rect 1111 6317 1118 6343
rect 1056 6313 1118 6317
rect 1018 6309 1118 6313
rect 494 6288 525 6309
rect 915 6288 951 6309
rect 337 6287 374 6288
rect 111 6284 145 6285
rect 110 6275 147 6284
rect 110 6257 119 6275
rect 137 6257 147 6275
rect 110 6247 147 6257
rect 336 6278 374 6287
rect 336 6258 345 6278
rect 365 6258 374 6278
rect 336 6250 374 6258
rect 440 6282 525 6288
rect 550 6287 587 6288
rect 440 6262 448 6282
rect 468 6262 525 6282
rect 440 6254 525 6262
rect 549 6278 587 6287
rect 549 6258 558 6278
rect 578 6258 587 6278
rect 440 6253 476 6254
rect 549 6250 587 6258
rect 653 6282 738 6288
rect 758 6287 795 6288
rect 653 6262 661 6282
rect 681 6281 738 6282
rect 681 6262 710 6281
rect 653 6261 710 6262
rect 731 6261 738 6281
rect 653 6254 738 6261
rect 757 6278 795 6287
rect 757 6258 766 6278
rect 786 6258 795 6278
rect 653 6253 689 6254
rect 757 6250 795 6258
rect 861 6282 1005 6288
rect 861 6262 869 6282
rect 889 6281 977 6282
rect 889 6262 920 6281
rect 861 6261 920 6262
rect 945 6262 977 6281
rect 997 6262 1005 6282
rect 945 6261 1005 6262
rect 861 6254 1005 6261
rect 861 6253 897 6254
rect 969 6253 1005 6254
rect 1071 6287 1108 6288
rect 1071 6286 1109 6287
rect 1071 6278 1135 6286
rect 1071 6258 1080 6278
rect 1100 6264 1135 6278
rect 1155 6264 1158 6284
rect 1100 6259 1158 6264
rect 1100 6258 1135 6259
rect 111 6219 145 6247
rect 337 6221 374 6250
rect 338 6219 374 6221
rect 550 6219 587 6250
rect 111 6218 283 6219
rect 111 6186 297 6218
rect 338 6197 587 6219
rect 758 6218 795 6250
rect 1071 6246 1135 6258
rect 1175 6220 1202 6398
rect 2169 6362 2230 6469
rect 3730 6376 3757 6554
rect 3797 6516 3861 6528
rect 4137 6524 4174 6556
rect 4345 6555 4594 6577
rect 4345 6524 4382 6555
rect 4558 6553 4594 6555
rect 4558 6524 4595 6553
rect 3797 6515 3832 6516
rect 3774 6510 3832 6515
rect 3774 6490 3777 6510
rect 3797 6496 3832 6510
rect 3852 6496 3861 6516
rect 3797 6488 3861 6496
rect 3823 6487 3861 6488
rect 3824 6486 3861 6487
rect 3927 6520 3963 6521
rect 4035 6520 4071 6521
rect 3927 6515 4071 6520
rect 3927 6512 3989 6515
rect 3927 6492 3935 6512
rect 3955 6495 3989 6512
rect 4012 6512 4071 6515
rect 4012 6495 4043 6512
rect 3955 6492 4043 6495
rect 4063 6492 4071 6512
rect 3927 6486 4071 6492
rect 4137 6516 4175 6524
rect 4243 6520 4279 6521
rect 4137 6496 4146 6516
rect 4166 6496 4175 6516
rect 4137 6487 4175 6496
rect 4194 6513 4279 6520
rect 4194 6493 4201 6513
rect 4222 6512 4279 6513
rect 4222 6493 4251 6512
rect 4194 6492 4251 6493
rect 4271 6492 4279 6512
rect 4137 6486 4174 6487
rect 4194 6486 4279 6492
rect 4345 6516 4383 6524
rect 4456 6520 4492 6521
rect 4345 6496 4354 6516
rect 4374 6496 4383 6516
rect 4345 6487 4383 6496
rect 4407 6512 4492 6520
rect 4407 6492 4464 6512
rect 4484 6492 4492 6512
rect 4345 6486 4382 6487
rect 4407 6486 4492 6492
rect 4558 6516 4596 6524
rect 4558 6496 4567 6516
rect 4587 6496 4596 6516
rect 4558 6487 4596 6496
rect 4558 6486 4595 6487
rect 3981 6465 4017 6486
rect 4407 6465 4438 6486
rect 3814 6461 3914 6465
rect 3814 6457 3876 6461
rect 3814 6431 3821 6457
rect 3847 6435 3876 6457
rect 3902 6435 3914 6461
rect 3847 6431 3914 6435
rect 3814 6428 3914 6431
rect 3982 6428 4017 6465
rect 4079 6462 4438 6465
rect 4079 6457 4301 6462
rect 4079 6433 4092 6457
rect 4116 6438 4301 6457
rect 4325 6438 4438 6462
rect 4116 6433 4438 6438
rect 4079 6429 4438 6433
rect 4505 6457 4654 6465
rect 4505 6437 4516 6457
rect 4536 6437 4654 6457
rect 4505 6430 4654 6437
rect 4505 6429 4546 6430
rect 3829 6376 3866 6377
rect 3925 6376 3962 6377
rect 3981 6376 4017 6428
rect 4036 6376 4073 6377
rect 3729 6367 3867 6376
rect 2169 6351 2239 6362
rect 2169 6342 2176 6351
rect 2171 6322 2176 6342
rect 2224 6322 2239 6351
rect 3729 6347 3838 6367
rect 3858 6347 3867 6367
rect 3729 6340 3867 6347
rect 3925 6367 4073 6376
rect 3925 6347 3934 6367
rect 3954 6347 4044 6367
rect 4064 6347 4073 6367
rect 3729 6338 3825 6340
rect 3925 6337 4073 6347
rect 4132 6367 4169 6377
rect 4244 6376 4281 6377
rect 4225 6374 4281 6376
rect 4132 6347 4140 6367
rect 4160 6347 4169 6367
rect 3981 6336 4017 6337
rect 2171 6313 2239 6322
rect 1358 6294 1468 6308
rect 1358 6291 1401 6294
rect 1358 6286 1362 6291
rect 1034 6218 1202 6220
rect 758 6212 1202 6218
rect 111 6154 145 6186
rect 107 6145 145 6154
rect 107 6127 117 6145
rect 135 6127 145 6145
rect 107 6121 145 6127
rect 263 6123 297 6186
rect 419 6191 530 6197
rect 419 6183 460 6191
rect 419 6163 427 6183
rect 446 6163 460 6183
rect 419 6161 460 6163
rect 488 6183 530 6191
rect 488 6163 504 6183
rect 523 6163 530 6183
rect 488 6161 530 6163
rect 419 6146 530 6161
rect 757 6192 1202 6212
rect 757 6123 795 6192
rect 1034 6191 1202 6192
rect 1280 6264 1362 6286
rect 1391 6264 1401 6291
rect 1429 6267 1436 6294
rect 1465 6286 1468 6294
rect 3463 6303 3574 6318
rect 3463 6301 3505 6303
rect 1465 6267 1530 6286
rect 1429 6264 1530 6267
rect 1280 6262 1530 6264
rect 1280 6183 1317 6262
rect 1358 6249 1468 6262
rect 1432 6193 1463 6194
rect 1280 6163 1289 6183
rect 1309 6163 1317 6183
rect 1280 6153 1317 6163
rect 1376 6183 1463 6193
rect 1376 6163 1385 6183
rect 1405 6163 1463 6183
rect 1376 6154 1463 6163
rect 1376 6153 1413 6154
rect 107 6117 144 6121
rect 263 6112 795 6123
rect 262 6096 795 6112
rect 1432 6101 1463 6154
rect 1493 6183 1530 6262
rect 1701 6259 2094 6279
rect 2114 6259 2117 6279
rect 3196 6274 3237 6283
rect 1701 6254 2117 6259
rect 2791 6272 2959 6273
rect 3196 6272 3205 6274
rect 1701 6253 2042 6254
rect 1645 6193 1676 6194
rect 1493 6163 1502 6183
rect 1522 6163 1530 6183
rect 1493 6153 1530 6163
rect 1589 6186 1676 6193
rect 1589 6183 1650 6186
rect 1589 6163 1598 6183
rect 1618 6166 1650 6183
rect 1671 6166 1676 6186
rect 1618 6163 1676 6166
rect 1589 6156 1676 6163
rect 1701 6183 1738 6253
rect 2004 6252 2041 6253
rect 2791 6252 3205 6272
rect 3231 6252 3237 6274
rect 3463 6281 3470 6301
rect 3489 6281 3505 6301
rect 3463 6273 3505 6281
rect 3533 6301 3574 6303
rect 3533 6281 3547 6301
rect 3566 6281 3574 6301
rect 3533 6273 3574 6281
rect 3829 6277 3866 6278
rect 4132 6277 4169 6347
rect 4194 6367 4281 6374
rect 4194 6364 4252 6367
rect 4194 6344 4199 6364
rect 4220 6347 4252 6364
rect 4272 6347 4281 6367
rect 4220 6344 4281 6347
rect 4194 6337 4281 6344
rect 4340 6367 4377 6377
rect 4340 6347 4348 6367
rect 4368 6347 4377 6367
rect 4194 6336 4225 6337
rect 3828 6276 4169 6277
rect 3463 6267 3574 6273
rect 3753 6271 4169 6276
rect 2791 6246 3237 6252
rect 2791 6244 2959 6246
rect 1853 6193 1889 6194
rect 1701 6163 1710 6183
rect 1730 6163 1738 6183
rect 1589 6154 1645 6156
rect 1589 6153 1626 6154
rect 1701 6153 1738 6163
rect 1797 6183 1945 6193
rect 2045 6190 2141 6192
rect 1797 6163 1806 6183
rect 1826 6163 1916 6183
rect 1936 6163 1945 6183
rect 1797 6154 1945 6163
rect 2003 6183 2141 6190
rect 2003 6163 2012 6183
rect 2032 6163 2141 6183
rect 2003 6154 2141 6163
rect 1797 6153 1834 6154
rect 1853 6102 1889 6154
rect 1908 6153 1945 6154
rect 2004 6153 2041 6154
rect 1324 6100 1365 6101
rect 262 6095 776 6096
rect 1216 6093 1365 6100
rect 1216 6073 1334 6093
rect 1354 6073 1365 6093
rect 1216 6065 1365 6073
rect 1432 6097 1791 6101
rect 1432 6092 1754 6097
rect 1432 6068 1545 6092
rect 1569 6073 1754 6092
rect 1778 6073 1791 6097
rect 1569 6068 1791 6073
rect 1432 6065 1791 6068
rect 1853 6065 1888 6102
rect 1956 6099 2056 6102
rect 1956 6095 2023 6099
rect 1956 6069 1968 6095
rect 1994 6073 2023 6095
rect 2049 6073 2056 6099
rect 1994 6069 2056 6073
rect 1956 6065 2056 6069
rect 110 6054 147 6055
rect 108 6046 148 6054
rect 108 6028 119 6046
rect 137 6028 148 6046
rect 1432 6044 1463 6065
rect 1853 6044 1889 6065
rect 1275 6043 1312 6044
rect 108 5980 148 6028
rect 1274 6034 1312 6043
rect 1274 6014 1283 6034
rect 1303 6014 1312 6034
rect 1274 6006 1312 6014
rect 1378 6038 1463 6044
rect 1488 6043 1525 6044
rect 1378 6018 1386 6038
rect 1406 6018 1463 6038
rect 1378 6010 1463 6018
rect 1487 6034 1525 6043
rect 1487 6014 1496 6034
rect 1516 6014 1525 6034
rect 1378 6009 1414 6010
rect 1487 6006 1525 6014
rect 1591 6038 1676 6044
rect 1696 6043 1733 6044
rect 1591 6018 1599 6038
rect 1619 6037 1676 6038
rect 1619 6018 1648 6037
rect 1591 6017 1648 6018
rect 1669 6017 1676 6037
rect 1591 6010 1676 6017
rect 1695 6034 1733 6043
rect 1695 6014 1704 6034
rect 1724 6014 1733 6034
rect 1591 6009 1627 6010
rect 1695 6006 1733 6014
rect 1799 6038 1943 6044
rect 1799 6018 1807 6038
rect 1827 6021 1863 6038
rect 1883 6021 1915 6038
rect 1827 6018 1915 6021
rect 1935 6018 1943 6038
rect 1799 6010 1943 6018
rect 1799 6009 1835 6010
rect 1907 6009 1943 6010
rect 2009 6043 2046 6044
rect 2009 6042 2047 6043
rect 2009 6034 2073 6042
rect 2009 6014 2018 6034
rect 2038 6020 2073 6034
rect 2093 6020 2096 6040
rect 2038 6015 2096 6020
rect 2038 6014 2073 6015
rect 419 5984 529 5998
rect 419 5981 462 5984
rect 108 5973 233 5980
rect 419 5976 423 5981
rect 108 5954 200 5973
rect 225 5954 233 5973
rect 108 5944 233 5954
rect 341 5954 423 5976
rect 452 5954 462 5981
rect 490 5957 497 5984
rect 526 5976 529 5984
rect 1275 5977 1312 6006
rect 526 5957 591 5976
rect 1276 5975 1312 5977
rect 1488 5975 1525 6006
rect 1696 5979 1733 6006
rect 2009 6002 2073 6014
rect 490 5954 591 5957
rect 341 5952 591 5954
rect 108 5924 148 5944
rect 107 5915 148 5924
rect 107 5897 117 5915
rect 135 5897 148 5915
rect 107 5888 148 5897
rect 107 5887 144 5888
rect 341 5873 378 5952
rect 419 5939 529 5952
rect 493 5883 524 5884
rect 341 5853 350 5873
rect 370 5853 378 5873
rect 341 5843 378 5853
rect 437 5873 524 5883
rect 437 5853 446 5873
rect 466 5853 524 5873
rect 437 5844 524 5853
rect 437 5843 474 5844
rect 110 5821 147 5825
rect 107 5816 147 5821
rect 107 5798 119 5816
rect 137 5798 147 5816
rect 107 5618 147 5798
rect 493 5791 524 5844
rect 554 5873 591 5952
rect 762 5949 1155 5969
rect 1175 5949 1178 5969
rect 1276 5953 1525 5975
rect 1694 5974 1735 5979
rect 2113 5976 2140 6154
rect 2791 6066 2818 6244
rect 3196 6241 3237 6246
rect 3406 6245 3655 6267
rect 3753 6251 3756 6271
rect 3776 6251 4169 6271
rect 4340 6268 4377 6347
rect 4407 6376 4438 6429
rect 4784 6422 4824 6602
rect 4784 6404 4794 6422
rect 4812 6404 4824 6422
rect 4784 6399 4824 6404
rect 4784 6395 4821 6399
rect 4457 6376 4494 6377
rect 4407 6367 4494 6376
rect 4407 6347 4465 6367
rect 4485 6347 4494 6367
rect 4407 6337 4494 6347
rect 4553 6367 4590 6377
rect 4553 6347 4561 6367
rect 4581 6347 4590 6367
rect 4407 6336 4438 6337
rect 4402 6268 4512 6281
rect 4553 6268 4590 6347
rect 4787 6332 4824 6333
rect 4783 6323 4824 6332
rect 4783 6305 4796 6323
rect 4814 6305 4824 6323
rect 4783 6296 4824 6305
rect 4783 6276 4823 6296
rect 4340 6266 4590 6268
rect 4340 6263 4441 6266
rect 2858 6206 2922 6218
rect 3198 6214 3235 6241
rect 3406 6214 3443 6245
rect 3619 6243 3655 6245
rect 4340 6244 4405 6263
rect 3619 6214 3656 6243
rect 4402 6236 4405 6244
rect 4434 6236 4441 6263
rect 4469 6239 4479 6266
rect 4508 6244 4590 6266
rect 4698 6266 4823 6276
rect 4698 6247 4706 6266
rect 4731 6247 4823 6266
rect 4508 6239 4512 6244
rect 4698 6240 4823 6247
rect 4469 6236 4512 6239
rect 4402 6222 4512 6236
rect 2858 6205 2893 6206
rect 2835 6200 2893 6205
rect 2835 6180 2838 6200
rect 2858 6186 2893 6200
rect 2913 6186 2922 6206
rect 2858 6178 2922 6186
rect 2884 6177 2922 6178
rect 2885 6176 2922 6177
rect 2988 6210 3024 6211
rect 3096 6210 3132 6211
rect 2988 6202 3132 6210
rect 2988 6182 2996 6202
rect 3016 6182 3104 6202
rect 3124 6182 3132 6202
rect 2988 6176 3132 6182
rect 3198 6206 3236 6214
rect 3304 6210 3340 6211
rect 3198 6186 3207 6206
rect 3227 6186 3236 6206
rect 3198 6177 3236 6186
rect 3255 6203 3340 6210
rect 3255 6183 3262 6203
rect 3283 6202 3340 6203
rect 3283 6183 3312 6202
rect 3255 6182 3312 6183
rect 3332 6182 3340 6202
rect 3198 6176 3235 6177
rect 3255 6176 3340 6182
rect 3406 6206 3444 6214
rect 3517 6210 3553 6211
rect 3406 6186 3415 6206
rect 3435 6186 3444 6206
rect 3406 6177 3444 6186
rect 3468 6202 3553 6210
rect 3468 6182 3525 6202
rect 3545 6182 3553 6202
rect 3406 6176 3443 6177
rect 3468 6176 3553 6182
rect 3619 6206 3657 6214
rect 3619 6186 3628 6206
rect 3648 6186 3657 6206
rect 3619 6177 3657 6186
rect 4783 6192 4823 6240
rect 3619 6176 3656 6177
rect 3042 6155 3078 6176
rect 3468 6155 3499 6176
rect 4783 6174 4794 6192
rect 4812 6174 4823 6192
rect 4783 6166 4823 6174
rect 4784 6165 4821 6166
rect 2875 6151 2975 6155
rect 2875 6147 2937 6151
rect 2875 6121 2882 6147
rect 2908 6125 2937 6147
rect 2963 6125 2975 6151
rect 2908 6121 2975 6125
rect 2875 6118 2975 6121
rect 3043 6118 3078 6155
rect 3140 6152 3499 6155
rect 3140 6147 3362 6152
rect 3140 6123 3153 6147
rect 3177 6128 3362 6147
rect 3386 6128 3499 6152
rect 3177 6123 3499 6128
rect 3140 6119 3499 6123
rect 3566 6147 3715 6155
rect 3566 6127 3577 6147
rect 3597 6127 3715 6147
rect 3566 6120 3715 6127
rect 4155 6124 4669 6125
rect 3566 6119 3607 6120
rect 3042 6083 3078 6118
rect 2890 6066 2927 6067
rect 2986 6066 3023 6067
rect 3042 6066 3049 6083
rect 2790 6057 2928 6066
rect 2790 6037 2899 6057
rect 2919 6037 2928 6057
rect 2790 6030 2928 6037
rect 2986 6057 3049 6066
rect 2986 6037 2995 6057
rect 3015 6042 3049 6057
rect 3070 6066 3078 6083
rect 3097 6066 3134 6067
rect 3070 6057 3134 6066
rect 3070 6042 3105 6057
rect 3015 6037 3105 6042
rect 3125 6037 3134 6057
rect 2790 6028 2886 6030
rect 2986 6027 3134 6037
rect 3193 6057 3230 6067
rect 3305 6066 3342 6067
rect 3286 6064 3342 6066
rect 3193 6037 3201 6057
rect 3221 6037 3230 6057
rect 3042 6026 3078 6027
rect 1972 5974 2140 5976
rect 1694 5968 2140 5974
rect 762 5944 1178 5949
rect 1357 5947 1468 5953
rect 762 5943 1103 5944
rect 706 5883 737 5884
rect 554 5853 563 5873
rect 583 5853 591 5873
rect 554 5843 591 5853
rect 650 5876 737 5883
rect 650 5873 711 5876
rect 650 5853 659 5873
rect 679 5856 711 5873
rect 732 5856 737 5876
rect 679 5853 737 5856
rect 650 5846 737 5853
rect 762 5873 799 5943
rect 1065 5942 1102 5943
rect 1357 5939 1398 5947
rect 1357 5919 1365 5939
rect 1384 5919 1398 5939
rect 1357 5917 1398 5919
rect 1426 5939 1468 5947
rect 1426 5919 1442 5939
rect 1461 5919 1468 5939
rect 1694 5946 1700 5968
rect 1726 5948 2140 5968
rect 2890 5967 2927 5968
rect 3193 5967 3230 6037
rect 3255 6057 3342 6064
rect 3255 6054 3313 6057
rect 3255 6034 3260 6054
rect 3281 6037 3313 6054
rect 3333 6037 3342 6057
rect 3281 6034 3342 6037
rect 3255 6027 3342 6034
rect 3401 6057 3438 6067
rect 3401 6037 3409 6057
rect 3429 6037 3438 6057
rect 3255 6026 3286 6027
rect 2889 5966 3230 5967
rect 1726 5946 1735 5948
rect 1972 5947 2140 5948
rect 2814 5965 3230 5966
rect 2814 5961 3190 5965
rect 1694 5937 1735 5946
rect 2814 5941 2817 5961
rect 2837 5948 3190 5961
rect 3222 5948 3230 5965
rect 2837 5941 3230 5948
rect 3401 5958 3438 6037
rect 3468 6066 3499 6119
rect 4136 6108 4669 6124
rect 4136 6097 4668 6108
rect 4787 6099 4824 6103
rect 3518 6066 3555 6067
rect 3468 6057 3555 6066
rect 3468 6037 3526 6057
rect 3546 6037 3555 6057
rect 3468 6027 3555 6037
rect 3614 6057 3651 6067
rect 3614 6037 3622 6057
rect 3642 6037 3651 6057
rect 3468 6026 3499 6027
rect 3463 5958 3573 5971
rect 3614 5958 3651 6037
rect 3401 5956 3651 5958
rect 3401 5953 3502 5956
rect 3401 5934 3466 5953
rect 1426 5917 1468 5919
rect 1357 5902 1468 5917
rect 3463 5926 3466 5934
rect 3495 5926 3502 5953
rect 3530 5929 3540 5956
rect 3569 5934 3651 5956
rect 3729 6028 3897 6029
rect 4136 6028 4174 6097
rect 3729 6008 4174 6028
rect 4401 6059 4512 6074
rect 4401 6057 4443 6059
rect 4401 6037 4408 6057
rect 4427 6037 4443 6057
rect 4401 6029 4443 6037
rect 4471 6057 4512 6059
rect 4471 6037 4485 6057
rect 4504 6037 4512 6057
rect 4471 6029 4512 6037
rect 4401 6023 4512 6029
rect 4634 6034 4668 6097
rect 4786 6093 4824 6099
rect 4786 6075 4796 6093
rect 4814 6075 4824 6093
rect 4786 6066 4824 6075
rect 4786 6034 4820 6066
rect 3729 6002 4173 6008
rect 3729 6000 3897 6002
rect 3569 5929 3573 5934
rect 3530 5926 3573 5929
rect 3463 5912 3573 5926
rect 914 5883 950 5884
rect 762 5853 771 5873
rect 791 5853 799 5873
rect 650 5844 706 5846
rect 650 5843 687 5844
rect 762 5843 799 5853
rect 858 5873 1006 5883
rect 1106 5880 1202 5882
rect 858 5853 867 5873
rect 887 5853 977 5873
rect 997 5853 1006 5873
rect 858 5844 1006 5853
rect 1064 5873 1202 5880
rect 1064 5853 1073 5873
rect 1093 5853 1202 5873
rect 1064 5844 1202 5853
rect 858 5843 895 5844
rect 914 5792 950 5844
rect 969 5843 1006 5844
rect 1065 5843 1102 5844
rect 385 5790 426 5791
rect 277 5783 426 5790
rect 277 5763 395 5783
rect 415 5763 426 5783
rect 277 5755 426 5763
rect 493 5787 852 5791
rect 493 5782 815 5787
rect 493 5758 606 5782
rect 630 5763 815 5782
rect 839 5763 852 5787
rect 630 5758 852 5763
rect 493 5755 852 5758
rect 914 5755 949 5792
rect 1017 5789 1117 5792
rect 1017 5785 1084 5789
rect 1017 5759 1029 5785
rect 1055 5763 1084 5785
rect 1110 5763 1117 5789
rect 1055 5759 1117 5763
rect 1017 5755 1117 5759
rect 493 5734 524 5755
rect 914 5734 950 5755
rect 336 5733 373 5734
rect 335 5724 373 5733
rect 335 5704 344 5724
rect 364 5704 373 5724
rect 335 5696 373 5704
rect 439 5728 524 5734
rect 549 5733 586 5734
rect 439 5708 447 5728
rect 467 5708 524 5728
rect 439 5700 524 5708
rect 548 5724 586 5733
rect 548 5704 557 5724
rect 577 5704 586 5724
rect 439 5699 475 5700
rect 548 5696 586 5704
rect 652 5728 737 5734
rect 757 5733 794 5734
rect 652 5708 660 5728
rect 680 5727 737 5728
rect 680 5708 709 5727
rect 652 5707 709 5708
rect 730 5707 737 5727
rect 652 5700 737 5707
rect 756 5724 794 5733
rect 756 5704 765 5724
rect 785 5704 794 5724
rect 652 5699 688 5700
rect 756 5696 794 5704
rect 860 5728 1004 5734
rect 860 5708 868 5728
rect 888 5725 976 5728
rect 888 5708 919 5725
rect 860 5705 919 5708
rect 942 5708 976 5725
rect 996 5708 1004 5728
rect 942 5705 1004 5708
rect 860 5700 1004 5705
rect 860 5699 896 5700
rect 968 5699 1004 5700
rect 1070 5733 1107 5734
rect 1070 5732 1108 5733
rect 1070 5724 1134 5732
rect 1070 5704 1079 5724
rect 1099 5710 1134 5724
rect 1154 5710 1157 5730
rect 1099 5705 1157 5710
rect 1099 5704 1134 5705
rect 336 5667 373 5696
rect 337 5665 373 5667
rect 549 5665 586 5696
rect 337 5643 586 5665
rect 757 5664 794 5696
rect 1070 5692 1134 5704
rect 1174 5666 1201 5844
rect 3729 5822 3756 6000
rect 3796 5962 3860 5974
rect 4136 5970 4173 6002
rect 4344 6001 4593 6023
rect 4634 6002 4820 6034
rect 4648 6001 4820 6002
rect 4344 5970 4381 6001
rect 4557 5999 4593 6001
rect 4557 5970 4594 5999
rect 4786 5973 4820 6001
rect 3796 5961 3831 5962
rect 3773 5956 3831 5961
rect 3773 5936 3776 5956
rect 3796 5942 3831 5956
rect 3851 5942 3860 5962
rect 3796 5934 3860 5942
rect 3822 5933 3860 5934
rect 3823 5932 3860 5933
rect 3926 5966 3962 5967
rect 4034 5966 4070 5967
rect 3926 5959 4070 5966
rect 3926 5958 3986 5959
rect 3926 5938 3934 5958
rect 3954 5939 3986 5958
rect 4011 5958 4070 5959
rect 4011 5939 4042 5958
rect 3954 5938 4042 5939
rect 4062 5938 4070 5958
rect 3926 5932 4070 5938
rect 4136 5962 4174 5970
rect 4242 5966 4278 5967
rect 4136 5942 4145 5962
rect 4165 5942 4174 5962
rect 4136 5933 4174 5942
rect 4193 5959 4278 5966
rect 4193 5939 4200 5959
rect 4221 5958 4278 5959
rect 4221 5939 4250 5958
rect 4193 5938 4250 5939
rect 4270 5938 4278 5958
rect 4136 5932 4173 5933
rect 4193 5932 4278 5938
rect 4344 5962 4382 5970
rect 4455 5966 4491 5967
rect 4344 5942 4353 5962
rect 4373 5942 4382 5962
rect 4344 5933 4382 5942
rect 4406 5958 4491 5966
rect 4406 5938 4463 5958
rect 4483 5938 4491 5958
rect 4344 5932 4381 5933
rect 4406 5932 4491 5938
rect 4557 5962 4595 5970
rect 4557 5942 4566 5962
rect 4586 5942 4595 5962
rect 4557 5933 4595 5942
rect 4784 5963 4821 5973
rect 4784 5945 4794 5963
rect 4812 5945 4821 5963
rect 4784 5936 4821 5945
rect 4786 5935 4820 5936
rect 4557 5932 4594 5933
rect 3980 5911 4016 5932
rect 4406 5911 4437 5932
rect 3813 5907 3913 5911
rect 3813 5903 3875 5907
rect 3813 5877 3820 5903
rect 3846 5881 3875 5903
rect 3901 5881 3913 5907
rect 3846 5877 3913 5881
rect 3813 5874 3913 5877
rect 3981 5874 4016 5911
rect 4078 5908 4437 5911
rect 4078 5903 4300 5908
rect 4078 5879 4091 5903
rect 4115 5884 4300 5903
rect 4324 5884 4437 5908
rect 4115 5879 4437 5884
rect 4078 5875 4437 5879
rect 4504 5903 4653 5911
rect 4504 5883 4515 5903
rect 4535 5883 4653 5903
rect 4504 5876 4653 5883
rect 4504 5875 4545 5876
rect 3828 5822 3865 5823
rect 3924 5822 3961 5823
rect 3980 5822 4016 5874
rect 4035 5822 4072 5823
rect 3728 5813 3866 5822
rect 3323 5792 3434 5807
rect 3323 5790 3365 5792
rect 2993 5769 3098 5771
rect 2651 5761 2819 5762
rect 2993 5761 3042 5769
rect 2651 5742 3042 5761
rect 3073 5742 3098 5769
rect 3323 5770 3330 5790
rect 3349 5770 3365 5790
rect 3323 5762 3365 5770
rect 3393 5790 3434 5792
rect 3393 5770 3407 5790
rect 3426 5770 3434 5790
rect 3728 5793 3837 5813
rect 3857 5793 3866 5813
rect 3728 5786 3866 5793
rect 3924 5813 4072 5822
rect 3924 5793 3933 5813
rect 3953 5793 4043 5813
rect 4063 5793 4072 5813
rect 3728 5784 3824 5786
rect 3924 5783 4072 5793
rect 4131 5813 4168 5823
rect 4243 5822 4280 5823
rect 4224 5820 4280 5822
rect 4131 5793 4139 5813
rect 4159 5793 4168 5813
rect 3980 5782 4016 5783
rect 3393 5762 3434 5770
rect 3323 5756 3434 5762
rect 2651 5735 3098 5742
rect 2651 5733 2819 5735
rect 1499 5702 1609 5716
rect 1499 5699 1542 5702
rect 1499 5694 1503 5699
rect 1033 5664 1201 5666
rect 757 5661 1201 5664
rect 418 5637 529 5643
rect 418 5629 459 5637
rect 107 5574 146 5618
rect 418 5609 426 5629
rect 445 5609 459 5629
rect 418 5607 459 5609
rect 487 5629 529 5637
rect 487 5609 503 5629
rect 522 5609 529 5629
rect 487 5607 529 5609
rect 418 5592 529 5607
rect 755 5638 1201 5661
rect 107 5550 147 5574
rect 447 5550 494 5552
rect 755 5550 793 5638
rect 1033 5637 1201 5638
rect 1421 5672 1503 5694
rect 1532 5672 1542 5699
rect 1570 5675 1577 5702
rect 1606 5694 1609 5702
rect 1606 5675 1671 5694
rect 1570 5672 1671 5675
rect 1421 5670 1671 5672
rect 1421 5591 1458 5670
rect 1499 5657 1609 5670
rect 1573 5601 1604 5602
rect 1421 5571 1430 5591
rect 1450 5571 1458 5591
rect 1421 5561 1458 5571
rect 1517 5591 1604 5601
rect 1517 5571 1526 5591
rect 1546 5571 1604 5591
rect 1517 5562 1604 5571
rect 1517 5561 1554 5562
rect 107 5517 793 5550
rect 107 5460 146 5517
rect 755 5515 793 5517
rect 1573 5509 1604 5562
rect 1634 5591 1671 5670
rect 1842 5683 2235 5687
rect 1842 5666 1861 5683
rect 1881 5667 2235 5683
rect 2255 5667 2258 5687
rect 1881 5666 2258 5667
rect 1842 5662 2258 5666
rect 1842 5661 2183 5662
rect 1786 5601 1817 5602
rect 1634 5571 1643 5591
rect 1663 5571 1671 5591
rect 1634 5561 1671 5571
rect 1730 5594 1817 5601
rect 1730 5591 1791 5594
rect 1730 5571 1739 5591
rect 1759 5574 1791 5591
rect 1812 5574 1817 5594
rect 1759 5571 1817 5574
rect 1730 5564 1817 5571
rect 1842 5591 1879 5661
rect 2145 5660 2182 5661
rect 1994 5601 2030 5602
rect 1842 5571 1851 5591
rect 1871 5571 1879 5591
rect 1730 5562 1786 5564
rect 1730 5561 1767 5562
rect 1842 5561 1879 5571
rect 1938 5591 2086 5601
rect 2254 5600 2283 5601
rect 2186 5598 2283 5600
rect 1938 5571 1947 5591
rect 1967 5587 2057 5591
rect 1967 5571 2000 5587
rect 1938 5562 2000 5571
rect 1938 5561 1975 5562
rect 1994 5549 2000 5562
rect 2023 5571 2057 5587
rect 2077 5571 2086 5591
rect 2023 5562 2086 5571
rect 2144 5591 2283 5598
rect 2144 5571 2153 5591
rect 2173 5571 2283 5591
rect 2144 5562 2283 5571
rect 2023 5549 2030 5562
rect 2049 5561 2086 5562
rect 2145 5561 2182 5562
rect 1994 5510 2030 5549
rect 1465 5508 1506 5509
rect 1357 5501 1506 5508
rect 1357 5481 1475 5501
rect 1495 5481 1506 5501
rect 1357 5473 1506 5481
rect 1573 5505 1932 5509
rect 1573 5500 1895 5505
rect 1573 5476 1686 5500
rect 1710 5481 1895 5500
rect 1919 5481 1932 5505
rect 1710 5476 1932 5481
rect 1573 5473 1932 5476
rect 1994 5473 2029 5510
rect 2097 5507 2197 5510
rect 2097 5503 2164 5507
rect 2097 5477 2109 5503
rect 2135 5481 2164 5503
rect 2190 5481 2197 5507
rect 2135 5477 2197 5481
rect 2097 5473 2197 5477
rect 107 5458 155 5460
rect 107 5440 118 5458
rect 136 5440 155 5458
rect 1573 5452 1604 5473
rect 1994 5452 2030 5473
rect 1416 5451 1453 5452
rect 107 5431 155 5440
rect 108 5430 155 5431
rect 421 5435 531 5449
rect 421 5432 464 5435
rect 421 5427 425 5432
rect 343 5405 425 5427
rect 454 5405 464 5432
rect 492 5408 499 5435
rect 528 5427 531 5435
rect 1415 5442 1453 5451
rect 528 5408 593 5427
rect 1415 5422 1424 5442
rect 1444 5422 1453 5442
rect 492 5405 593 5408
rect 343 5403 593 5405
rect 111 5367 148 5368
rect 107 5364 148 5367
rect 107 5359 149 5364
rect 107 5341 120 5359
rect 138 5341 149 5359
rect 107 5327 149 5341
rect 187 5327 234 5331
rect 107 5321 234 5327
rect 107 5292 195 5321
rect 224 5292 234 5321
rect 343 5324 380 5403
rect 421 5390 531 5403
rect 495 5334 526 5335
rect 343 5304 352 5324
rect 372 5304 380 5324
rect 343 5294 380 5304
rect 439 5324 526 5334
rect 439 5304 448 5324
rect 468 5304 526 5324
rect 439 5295 526 5304
rect 439 5294 476 5295
rect 107 5288 234 5292
rect 107 5271 146 5288
rect 187 5287 234 5288
rect 107 5253 118 5271
rect 136 5253 146 5271
rect 107 5244 146 5253
rect 108 5243 145 5244
rect 495 5242 526 5295
rect 556 5324 593 5403
rect 764 5400 1157 5420
rect 1177 5400 1180 5420
rect 1415 5414 1453 5422
rect 1519 5446 1604 5452
rect 1629 5451 1666 5452
rect 1519 5426 1527 5446
rect 1547 5426 1604 5446
rect 1519 5418 1604 5426
rect 1628 5442 1666 5451
rect 1628 5422 1637 5442
rect 1657 5422 1666 5442
rect 1519 5417 1555 5418
rect 1628 5414 1666 5422
rect 1732 5446 1817 5452
rect 1837 5451 1874 5452
rect 1732 5426 1740 5446
rect 1760 5445 1817 5446
rect 1760 5426 1789 5445
rect 1732 5425 1789 5426
rect 1810 5425 1817 5445
rect 1732 5418 1817 5425
rect 1836 5442 1874 5451
rect 1836 5422 1845 5442
rect 1865 5422 1874 5442
rect 1732 5417 1768 5418
rect 1836 5414 1874 5422
rect 1940 5446 2084 5452
rect 1940 5426 1948 5446
rect 1968 5426 2056 5446
rect 2076 5426 2084 5446
rect 1940 5418 2084 5426
rect 1940 5417 1976 5418
rect 2048 5417 2084 5418
rect 2150 5451 2187 5452
rect 2150 5450 2188 5451
rect 2150 5442 2214 5450
rect 2150 5422 2159 5442
rect 2179 5428 2214 5442
rect 2234 5428 2237 5448
rect 2179 5423 2237 5428
rect 2179 5422 2214 5423
rect 764 5395 1180 5400
rect 764 5394 1105 5395
rect 708 5334 739 5335
rect 556 5304 565 5324
rect 585 5304 593 5324
rect 556 5294 593 5304
rect 652 5327 739 5334
rect 652 5324 713 5327
rect 652 5304 661 5324
rect 681 5307 713 5324
rect 734 5307 739 5327
rect 681 5304 739 5307
rect 652 5297 739 5304
rect 764 5324 801 5394
rect 1067 5393 1104 5394
rect 1416 5385 1453 5414
rect 1417 5383 1453 5385
rect 1629 5383 1666 5414
rect 1417 5361 1666 5383
rect 1837 5382 1874 5414
rect 2150 5410 2214 5422
rect 2254 5384 2283 5562
rect 2651 5555 2678 5733
rect 2718 5695 2782 5707
rect 3058 5703 3095 5735
rect 3266 5734 3515 5756
rect 3266 5703 3303 5734
rect 3479 5732 3515 5734
rect 3479 5703 3516 5732
rect 3828 5723 3865 5724
rect 4131 5723 4168 5793
rect 4193 5813 4280 5820
rect 4193 5810 4251 5813
rect 4193 5790 4198 5810
rect 4219 5793 4251 5810
rect 4271 5793 4280 5813
rect 4219 5790 4280 5793
rect 4193 5783 4280 5790
rect 4339 5813 4376 5823
rect 4339 5793 4347 5813
rect 4367 5793 4376 5813
rect 4193 5782 4224 5783
rect 3827 5722 4168 5723
rect 3752 5717 4168 5722
rect 2718 5694 2753 5695
rect 2695 5689 2753 5694
rect 2695 5669 2698 5689
rect 2718 5675 2753 5689
rect 2773 5675 2782 5695
rect 2718 5667 2782 5675
rect 2744 5666 2782 5667
rect 2745 5665 2782 5666
rect 2848 5699 2884 5700
rect 2956 5699 2992 5700
rect 2848 5694 2992 5699
rect 2848 5691 2908 5694
rect 2848 5671 2856 5691
rect 2876 5673 2908 5691
rect 2935 5691 2992 5694
rect 2935 5673 2964 5691
rect 2876 5671 2964 5673
rect 2984 5671 2992 5691
rect 2848 5665 2992 5671
rect 3058 5695 3096 5703
rect 3164 5699 3200 5700
rect 3058 5675 3067 5695
rect 3087 5675 3096 5695
rect 3058 5666 3096 5675
rect 3115 5692 3200 5699
rect 3115 5672 3122 5692
rect 3143 5691 3200 5692
rect 3143 5672 3172 5691
rect 3115 5671 3172 5672
rect 3192 5671 3200 5691
rect 3058 5665 3095 5666
rect 3115 5665 3200 5671
rect 3266 5695 3304 5703
rect 3377 5699 3413 5700
rect 3266 5675 3275 5695
rect 3295 5675 3304 5695
rect 3266 5666 3304 5675
rect 3328 5691 3413 5699
rect 3328 5671 3385 5691
rect 3405 5671 3413 5691
rect 3266 5665 3303 5666
rect 3328 5665 3413 5671
rect 3479 5695 3517 5703
rect 3752 5697 3755 5717
rect 3775 5697 4168 5717
rect 4339 5714 4376 5793
rect 4406 5822 4437 5875
rect 4787 5873 4824 5874
rect 4786 5864 4825 5873
rect 4786 5846 4796 5864
rect 4814 5846 4825 5864
rect 4698 5829 4745 5830
rect 4786 5829 4825 5846
rect 4698 5825 4825 5829
rect 4456 5822 4493 5823
rect 4406 5813 4493 5822
rect 4406 5793 4464 5813
rect 4484 5793 4493 5813
rect 4406 5783 4493 5793
rect 4552 5813 4589 5823
rect 4552 5793 4560 5813
rect 4580 5793 4589 5813
rect 4406 5782 4437 5783
rect 4401 5714 4511 5727
rect 4552 5714 4589 5793
rect 4698 5796 4708 5825
rect 4737 5796 4825 5825
rect 4698 5790 4825 5796
rect 4698 5786 4745 5790
rect 4783 5776 4825 5790
rect 4783 5758 4794 5776
rect 4812 5758 4825 5776
rect 4783 5753 4825 5758
rect 4784 5750 4825 5753
rect 4784 5749 4821 5750
rect 4339 5712 4589 5714
rect 4339 5709 4440 5712
rect 3479 5675 3488 5695
rect 3508 5675 3517 5695
rect 4339 5690 4404 5709
rect 3479 5666 3517 5675
rect 4401 5682 4404 5690
rect 4433 5682 4440 5709
rect 4468 5685 4478 5712
rect 4507 5690 4589 5712
rect 4507 5685 4511 5690
rect 4468 5682 4511 5685
rect 4401 5668 4511 5682
rect 4777 5686 4824 5687
rect 4777 5677 4825 5686
rect 3479 5665 3516 5666
rect 2902 5644 2938 5665
rect 3328 5644 3359 5665
rect 4777 5659 4796 5677
rect 4814 5659 4825 5677
rect 4777 5657 4825 5659
rect 2735 5640 2835 5644
rect 2735 5636 2797 5640
rect 2735 5610 2742 5636
rect 2768 5614 2797 5636
rect 2823 5614 2835 5640
rect 2768 5610 2835 5614
rect 2735 5607 2835 5610
rect 2903 5607 2938 5644
rect 3000 5641 3359 5644
rect 3000 5636 3222 5641
rect 3000 5612 3013 5636
rect 3037 5617 3222 5636
rect 3246 5617 3359 5641
rect 3037 5612 3359 5617
rect 3000 5608 3359 5612
rect 3426 5636 3575 5644
rect 3426 5616 3437 5636
rect 3457 5616 3575 5636
rect 3426 5609 3575 5616
rect 3426 5608 3467 5609
rect 2750 5555 2787 5556
rect 2846 5555 2883 5556
rect 2902 5555 2938 5607
rect 2957 5555 2994 5556
rect 2650 5546 2788 5555
rect 2650 5526 2759 5546
rect 2779 5526 2788 5546
rect 2650 5519 2788 5526
rect 2846 5546 2994 5555
rect 2846 5526 2855 5546
rect 2875 5526 2965 5546
rect 2985 5526 2994 5546
rect 2650 5517 2746 5519
rect 2846 5516 2994 5526
rect 3053 5546 3090 5556
rect 3165 5555 3202 5556
rect 3146 5553 3202 5555
rect 3053 5526 3061 5546
rect 3081 5526 3090 5546
rect 2902 5515 2938 5516
rect 2750 5456 2787 5457
rect 3053 5456 3090 5526
rect 3115 5546 3202 5553
rect 3115 5543 3173 5546
rect 3115 5523 3120 5543
rect 3141 5526 3173 5543
rect 3193 5526 3202 5546
rect 3141 5523 3202 5526
rect 3115 5516 3202 5523
rect 3261 5546 3298 5556
rect 3261 5526 3269 5546
rect 3289 5526 3298 5546
rect 3115 5515 3146 5516
rect 2749 5455 3090 5456
rect 2674 5451 3090 5455
rect 2674 5450 3051 5451
rect 2674 5430 2677 5450
rect 2697 5434 3051 5450
rect 3071 5434 3090 5451
rect 2697 5430 3090 5434
rect 3261 5447 3298 5526
rect 3328 5555 3359 5608
rect 4139 5600 4177 5602
rect 4786 5600 4825 5657
rect 4139 5567 4825 5600
rect 3378 5555 3415 5556
rect 3328 5546 3415 5555
rect 3328 5526 3386 5546
rect 3406 5526 3415 5546
rect 3328 5516 3415 5526
rect 3474 5546 3511 5556
rect 3474 5526 3482 5546
rect 3502 5526 3511 5546
rect 3328 5515 3359 5516
rect 3323 5447 3433 5460
rect 3474 5447 3511 5526
rect 3261 5445 3511 5447
rect 3261 5442 3362 5445
rect 3261 5423 3326 5442
rect 3323 5415 3326 5423
rect 3355 5415 3362 5442
rect 3390 5418 3400 5445
rect 3429 5423 3511 5445
rect 3731 5479 3899 5480
rect 4139 5479 4177 5567
rect 4438 5565 4485 5567
rect 4785 5543 4825 5567
rect 3731 5456 4177 5479
rect 4403 5510 4514 5525
rect 4403 5508 4445 5510
rect 4403 5488 4410 5508
rect 4429 5488 4445 5508
rect 4403 5480 4445 5488
rect 4473 5508 4514 5510
rect 4473 5488 4487 5508
rect 4506 5488 4514 5508
rect 4786 5499 4825 5543
rect 4473 5480 4514 5488
rect 4403 5474 4514 5480
rect 3731 5453 4175 5456
rect 3731 5451 3899 5453
rect 3429 5418 3433 5423
rect 3390 5415 3433 5418
rect 3323 5401 3433 5415
rect 2113 5382 2283 5384
rect 1834 5375 2283 5382
rect 1498 5355 1609 5361
rect 1498 5347 1539 5355
rect 916 5334 952 5335
rect 764 5304 773 5324
rect 793 5304 801 5324
rect 652 5295 708 5297
rect 652 5294 689 5295
rect 764 5294 801 5304
rect 860 5324 1008 5334
rect 1108 5331 1204 5333
rect 860 5304 869 5324
rect 889 5304 979 5324
rect 999 5304 1008 5324
rect 860 5295 1008 5304
rect 1066 5324 1204 5331
rect 1066 5304 1075 5324
rect 1095 5304 1204 5324
rect 1498 5327 1506 5347
rect 1525 5327 1539 5347
rect 1498 5325 1539 5327
rect 1567 5347 1609 5355
rect 1567 5327 1583 5347
rect 1602 5327 1609 5347
rect 1834 5348 1859 5375
rect 1890 5356 2283 5375
rect 1890 5348 1939 5356
rect 2113 5355 2283 5356
rect 1834 5346 1939 5348
rect 1567 5325 1609 5327
rect 1498 5310 1609 5325
rect 1066 5295 1204 5304
rect 860 5294 897 5295
rect 916 5243 952 5295
rect 971 5294 1008 5295
rect 1067 5294 1104 5295
rect 387 5241 428 5242
rect 279 5234 428 5241
rect 279 5214 397 5234
rect 417 5214 428 5234
rect 279 5206 428 5214
rect 495 5238 854 5242
rect 495 5233 817 5238
rect 495 5209 608 5233
rect 632 5214 817 5233
rect 841 5214 854 5238
rect 632 5209 854 5214
rect 495 5206 854 5209
rect 916 5206 951 5243
rect 1019 5240 1119 5243
rect 1019 5236 1086 5240
rect 1019 5210 1031 5236
rect 1057 5214 1086 5236
rect 1112 5214 1119 5240
rect 1057 5210 1119 5214
rect 1019 5206 1119 5210
rect 495 5185 526 5206
rect 916 5185 952 5206
rect 338 5184 375 5185
rect 112 5181 146 5182
rect 111 5172 148 5181
rect 111 5154 120 5172
rect 138 5154 148 5172
rect 111 5144 148 5154
rect 337 5175 375 5184
rect 337 5155 346 5175
rect 366 5155 375 5175
rect 337 5147 375 5155
rect 441 5179 526 5185
rect 551 5184 588 5185
rect 441 5159 449 5179
rect 469 5159 526 5179
rect 441 5151 526 5159
rect 550 5175 588 5184
rect 550 5155 559 5175
rect 579 5155 588 5175
rect 441 5150 477 5151
rect 550 5147 588 5155
rect 654 5179 739 5185
rect 759 5184 796 5185
rect 654 5159 662 5179
rect 682 5178 739 5179
rect 682 5159 711 5178
rect 654 5158 711 5159
rect 732 5158 739 5178
rect 654 5151 739 5158
rect 758 5175 796 5184
rect 758 5155 767 5175
rect 787 5155 796 5175
rect 654 5150 690 5151
rect 758 5147 796 5155
rect 862 5179 1006 5185
rect 862 5159 870 5179
rect 890 5178 978 5179
rect 890 5159 921 5178
rect 862 5158 921 5159
rect 946 5159 978 5178
rect 998 5159 1006 5179
rect 946 5158 1006 5159
rect 862 5151 1006 5158
rect 862 5150 898 5151
rect 970 5150 1006 5151
rect 1072 5184 1109 5185
rect 1072 5183 1110 5184
rect 1072 5175 1136 5183
rect 1072 5155 1081 5175
rect 1101 5161 1136 5175
rect 1156 5161 1159 5181
rect 1101 5156 1159 5161
rect 1101 5155 1136 5156
rect 112 5116 146 5144
rect 338 5118 375 5147
rect 339 5116 375 5118
rect 551 5116 588 5147
rect 112 5115 284 5116
rect 112 5083 298 5115
rect 339 5094 588 5116
rect 759 5115 796 5147
rect 1072 5143 1136 5155
rect 1176 5117 1203 5295
rect 3731 5273 3758 5451
rect 3798 5413 3862 5425
rect 4138 5421 4175 5453
rect 4346 5452 4595 5474
rect 4346 5421 4383 5452
rect 4559 5450 4595 5452
rect 4559 5421 4596 5450
rect 3798 5412 3833 5413
rect 3775 5407 3833 5412
rect 3775 5387 3778 5407
rect 3798 5393 3833 5407
rect 3853 5393 3862 5413
rect 3798 5385 3862 5393
rect 3824 5384 3862 5385
rect 3825 5383 3862 5384
rect 3928 5417 3964 5418
rect 4036 5417 4072 5418
rect 3928 5412 4072 5417
rect 3928 5409 3990 5412
rect 3928 5389 3936 5409
rect 3956 5392 3990 5409
rect 4013 5409 4072 5412
rect 4013 5392 4044 5409
rect 3956 5389 4044 5392
rect 4064 5389 4072 5409
rect 3928 5383 4072 5389
rect 4138 5413 4176 5421
rect 4244 5417 4280 5418
rect 4138 5393 4147 5413
rect 4167 5393 4176 5413
rect 4138 5384 4176 5393
rect 4195 5410 4280 5417
rect 4195 5390 4202 5410
rect 4223 5409 4280 5410
rect 4223 5390 4252 5409
rect 4195 5389 4252 5390
rect 4272 5389 4280 5409
rect 4138 5383 4175 5384
rect 4195 5383 4280 5389
rect 4346 5413 4384 5421
rect 4457 5417 4493 5418
rect 4346 5393 4355 5413
rect 4375 5393 4384 5413
rect 4346 5384 4384 5393
rect 4408 5409 4493 5417
rect 4408 5389 4465 5409
rect 4485 5389 4493 5409
rect 4346 5383 4383 5384
rect 4408 5383 4493 5389
rect 4559 5413 4597 5421
rect 4559 5393 4568 5413
rect 4588 5393 4597 5413
rect 4559 5384 4597 5393
rect 4559 5383 4596 5384
rect 3982 5362 4018 5383
rect 4408 5362 4439 5383
rect 3815 5358 3915 5362
rect 3815 5354 3877 5358
rect 3815 5328 3822 5354
rect 3848 5332 3877 5354
rect 3903 5332 3915 5358
rect 3848 5328 3915 5332
rect 3815 5325 3915 5328
rect 3983 5325 4018 5362
rect 4080 5359 4439 5362
rect 4080 5354 4302 5359
rect 4080 5330 4093 5354
rect 4117 5335 4302 5354
rect 4326 5335 4439 5359
rect 4117 5330 4439 5335
rect 4080 5326 4439 5330
rect 4506 5354 4655 5362
rect 4506 5334 4517 5354
rect 4537 5334 4655 5354
rect 4506 5327 4655 5334
rect 4506 5326 4547 5327
rect 3830 5273 3867 5274
rect 3926 5273 3963 5274
rect 3982 5273 4018 5325
rect 4037 5273 4074 5274
rect 3730 5264 3868 5273
rect 3730 5244 3839 5264
rect 3859 5244 3868 5264
rect 3730 5237 3868 5244
rect 3926 5264 4074 5273
rect 3926 5244 3935 5264
rect 3955 5244 4045 5264
rect 4065 5244 4074 5264
rect 3730 5235 3826 5237
rect 3926 5234 4074 5244
rect 4133 5264 4170 5274
rect 4245 5273 4282 5274
rect 4226 5271 4282 5273
rect 4133 5244 4141 5264
rect 4161 5244 4170 5264
rect 3982 5233 4018 5234
rect 1359 5191 1469 5205
rect 1359 5188 1402 5191
rect 1359 5183 1363 5188
rect 1035 5115 1203 5117
rect 759 5109 1203 5115
rect 112 5051 146 5083
rect 108 5042 146 5051
rect 108 5024 118 5042
rect 136 5024 146 5042
rect 108 5018 146 5024
rect 264 5020 298 5083
rect 420 5088 531 5094
rect 420 5080 461 5088
rect 420 5060 428 5080
rect 447 5060 461 5080
rect 420 5058 461 5060
rect 489 5080 531 5088
rect 489 5060 505 5080
rect 524 5060 531 5080
rect 489 5058 531 5060
rect 420 5043 531 5058
rect 758 5089 1203 5109
rect 758 5020 796 5089
rect 1035 5088 1203 5089
rect 1281 5161 1363 5183
rect 1392 5161 1402 5188
rect 1430 5164 1437 5191
rect 1466 5183 1469 5191
rect 3464 5200 3575 5215
rect 3464 5198 3506 5200
rect 1466 5164 1531 5183
rect 1430 5161 1531 5164
rect 1281 5159 1531 5161
rect 1281 5080 1318 5159
rect 1359 5146 1469 5159
rect 1433 5090 1464 5091
rect 1281 5060 1290 5080
rect 1310 5060 1318 5080
rect 1281 5050 1318 5060
rect 1377 5080 1464 5090
rect 1377 5060 1386 5080
rect 1406 5060 1464 5080
rect 1377 5051 1464 5060
rect 1377 5050 1414 5051
rect 108 5014 145 5018
rect 264 5009 796 5020
rect 263 4993 796 5009
rect 1433 4998 1464 5051
rect 1494 5080 1531 5159
rect 1702 5169 2095 5176
rect 1702 5152 1710 5169
rect 1742 5156 2095 5169
rect 2115 5156 2118 5176
rect 3197 5171 3238 5180
rect 1742 5152 2118 5156
rect 1702 5151 2118 5152
rect 2792 5169 2960 5170
rect 3197 5169 3206 5171
rect 1702 5150 2043 5151
rect 1646 5090 1677 5091
rect 1494 5060 1503 5080
rect 1523 5060 1531 5080
rect 1494 5050 1531 5060
rect 1590 5083 1677 5090
rect 1590 5080 1651 5083
rect 1590 5060 1599 5080
rect 1619 5063 1651 5080
rect 1672 5063 1677 5083
rect 1619 5060 1677 5063
rect 1590 5053 1677 5060
rect 1702 5080 1739 5150
rect 2005 5149 2042 5150
rect 2792 5149 3206 5169
rect 3232 5149 3238 5171
rect 3464 5178 3471 5198
rect 3490 5178 3506 5198
rect 3464 5170 3506 5178
rect 3534 5198 3575 5200
rect 3534 5178 3548 5198
rect 3567 5178 3575 5198
rect 3534 5170 3575 5178
rect 3830 5174 3867 5175
rect 4133 5174 4170 5244
rect 4195 5264 4282 5271
rect 4195 5261 4253 5264
rect 4195 5241 4200 5261
rect 4221 5244 4253 5261
rect 4273 5244 4282 5264
rect 4221 5241 4282 5244
rect 4195 5234 4282 5241
rect 4341 5264 4378 5274
rect 4341 5244 4349 5264
rect 4369 5244 4378 5264
rect 4195 5233 4226 5234
rect 3829 5173 4170 5174
rect 3464 5164 3575 5170
rect 3754 5168 4170 5173
rect 2792 5143 3238 5149
rect 2792 5141 2960 5143
rect 1854 5090 1890 5091
rect 1702 5060 1711 5080
rect 1731 5060 1739 5080
rect 1590 5051 1646 5053
rect 1590 5050 1627 5051
rect 1702 5050 1739 5060
rect 1798 5080 1946 5090
rect 2046 5087 2142 5089
rect 1798 5060 1807 5080
rect 1827 5075 1917 5080
rect 1827 5060 1862 5075
rect 1798 5051 1862 5060
rect 1798 5050 1835 5051
rect 1854 5034 1862 5051
rect 1883 5060 1917 5075
rect 1937 5060 1946 5080
rect 1883 5051 1946 5060
rect 2004 5080 2142 5087
rect 2004 5060 2013 5080
rect 2033 5060 2142 5080
rect 2004 5051 2142 5060
rect 1883 5034 1890 5051
rect 1909 5050 1946 5051
rect 2005 5050 2042 5051
rect 1854 4999 1890 5034
rect 1325 4997 1366 4998
rect 263 4992 777 4993
rect 1217 4990 1366 4997
rect 1217 4970 1335 4990
rect 1355 4970 1366 4990
rect 1217 4962 1366 4970
rect 1433 4994 1792 4998
rect 1433 4989 1755 4994
rect 1433 4965 1546 4989
rect 1570 4970 1755 4989
rect 1779 4970 1792 4994
rect 1570 4965 1792 4970
rect 1433 4962 1792 4965
rect 1854 4962 1889 4999
rect 1957 4996 2057 4999
rect 1957 4992 2024 4996
rect 1957 4966 1969 4992
rect 1995 4970 2024 4992
rect 2050 4970 2057 4996
rect 1995 4966 2057 4970
rect 1957 4962 2057 4966
rect 111 4951 148 4952
rect 109 4943 149 4951
rect 109 4925 120 4943
rect 138 4925 149 4943
rect 1433 4941 1464 4962
rect 1854 4941 1890 4962
rect 1276 4940 1313 4941
rect 109 4877 149 4925
rect 1275 4931 1313 4940
rect 1275 4911 1284 4931
rect 1304 4911 1313 4931
rect 1275 4903 1313 4911
rect 1379 4935 1464 4941
rect 1489 4940 1526 4941
rect 1379 4915 1387 4935
rect 1407 4915 1464 4935
rect 1379 4907 1464 4915
rect 1488 4931 1526 4940
rect 1488 4911 1497 4931
rect 1517 4911 1526 4931
rect 1379 4906 1415 4907
rect 1488 4903 1526 4911
rect 1592 4935 1677 4941
rect 1697 4940 1734 4941
rect 1592 4915 1600 4935
rect 1620 4934 1677 4935
rect 1620 4915 1649 4934
rect 1592 4914 1649 4915
rect 1670 4914 1677 4934
rect 1592 4907 1677 4914
rect 1696 4931 1734 4940
rect 1696 4911 1705 4931
rect 1725 4911 1734 4931
rect 1592 4906 1628 4907
rect 1696 4903 1734 4911
rect 1800 4935 1944 4941
rect 1800 4915 1808 4935
rect 1828 4915 1916 4935
rect 1936 4915 1944 4935
rect 1800 4907 1944 4915
rect 1800 4906 1836 4907
rect 1908 4906 1944 4907
rect 2010 4940 2047 4941
rect 2010 4939 2048 4940
rect 2010 4931 2074 4939
rect 2010 4911 2019 4931
rect 2039 4917 2074 4931
rect 2094 4917 2097 4937
rect 2039 4912 2097 4917
rect 2039 4911 2074 4912
rect 420 4881 530 4895
rect 420 4878 463 4881
rect 109 4870 234 4877
rect 420 4873 424 4878
rect 109 4851 201 4870
rect 226 4851 234 4870
rect 109 4841 234 4851
rect 342 4851 424 4873
rect 453 4851 463 4878
rect 491 4854 498 4881
rect 527 4873 530 4881
rect 1276 4874 1313 4903
rect 527 4854 592 4873
rect 1277 4872 1313 4874
rect 1489 4872 1526 4903
rect 1697 4876 1734 4903
rect 2010 4899 2074 4911
rect 491 4851 592 4854
rect 342 4849 592 4851
rect 109 4821 149 4841
rect 108 4812 149 4821
rect 108 4794 118 4812
rect 136 4794 149 4812
rect 108 4785 149 4794
rect 108 4784 145 4785
rect 342 4770 379 4849
rect 420 4836 530 4849
rect 494 4780 525 4781
rect 342 4750 351 4770
rect 371 4750 379 4770
rect 342 4740 379 4750
rect 438 4770 525 4780
rect 438 4750 447 4770
rect 467 4750 525 4770
rect 438 4741 525 4750
rect 438 4740 475 4741
rect 111 4718 148 4722
rect 108 4713 148 4718
rect 108 4695 120 4713
rect 138 4695 148 4713
rect 108 4515 148 4695
rect 494 4688 525 4741
rect 555 4770 592 4849
rect 763 4846 1156 4866
rect 1176 4846 1179 4866
rect 1277 4850 1526 4872
rect 1695 4871 1736 4876
rect 2114 4873 2141 5051
rect 2792 4963 2819 5141
rect 3197 5138 3238 5143
rect 3407 5142 3656 5164
rect 3754 5148 3757 5168
rect 3777 5148 4170 5168
rect 4341 5165 4378 5244
rect 4408 5273 4439 5326
rect 4785 5319 4825 5499
rect 4785 5301 4795 5319
rect 4813 5301 4825 5319
rect 4785 5296 4825 5301
rect 4785 5292 4822 5296
rect 4458 5273 4495 5274
rect 4408 5264 4495 5273
rect 4408 5244 4466 5264
rect 4486 5244 4495 5264
rect 4408 5234 4495 5244
rect 4554 5264 4591 5274
rect 4554 5244 4562 5264
rect 4582 5244 4591 5264
rect 4408 5233 4439 5234
rect 4403 5165 4513 5178
rect 4554 5165 4591 5244
rect 4788 5229 4825 5230
rect 4784 5220 4825 5229
rect 4784 5202 4797 5220
rect 4815 5202 4825 5220
rect 4784 5193 4825 5202
rect 4784 5173 4824 5193
rect 4341 5163 4591 5165
rect 4341 5160 4442 5163
rect 2859 5103 2923 5115
rect 3199 5111 3236 5138
rect 3407 5111 3444 5142
rect 3620 5140 3656 5142
rect 4341 5141 4406 5160
rect 3620 5111 3657 5140
rect 4403 5133 4406 5141
rect 4435 5133 4442 5160
rect 4470 5136 4480 5163
rect 4509 5141 4591 5163
rect 4699 5163 4824 5173
rect 4699 5144 4707 5163
rect 4732 5144 4824 5163
rect 4509 5136 4513 5141
rect 4699 5137 4824 5144
rect 4470 5133 4513 5136
rect 4403 5119 4513 5133
rect 2859 5102 2894 5103
rect 2836 5097 2894 5102
rect 2836 5077 2839 5097
rect 2859 5083 2894 5097
rect 2914 5083 2923 5103
rect 2859 5075 2923 5083
rect 2885 5074 2923 5075
rect 2886 5073 2923 5074
rect 2989 5107 3025 5108
rect 3097 5107 3133 5108
rect 2989 5099 3133 5107
rect 2989 5079 2997 5099
rect 3017 5096 3105 5099
rect 3017 5079 3049 5096
rect 3069 5079 3105 5096
rect 3125 5079 3133 5099
rect 2989 5073 3133 5079
rect 3199 5103 3237 5111
rect 3305 5107 3341 5108
rect 3199 5083 3208 5103
rect 3228 5083 3237 5103
rect 3199 5074 3237 5083
rect 3256 5100 3341 5107
rect 3256 5080 3263 5100
rect 3284 5099 3341 5100
rect 3284 5080 3313 5099
rect 3256 5079 3313 5080
rect 3333 5079 3341 5099
rect 3199 5073 3236 5074
rect 3256 5073 3341 5079
rect 3407 5103 3445 5111
rect 3518 5107 3554 5108
rect 3407 5083 3416 5103
rect 3436 5083 3445 5103
rect 3407 5074 3445 5083
rect 3469 5099 3554 5107
rect 3469 5079 3526 5099
rect 3546 5079 3554 5099
rect 3407 5073 3444 5074
rect 3469 5073 3554 5079
rect 3620 5103 3658 5111
rect 3620 5083 3629 5103
rect 3649 5083 3658 5103
rect 3620 5074 3658 5083
rect 4784 5089 4824 5137
rect 3620 5073 3657 5074
rect 3043 5052 3079 5073
rect 3469 5052 3500 5073
rect 4784 5071 4795 5089
rect 4813 5071 4824 5089
rect 4784 5063 4824 5071
rect 4785 5062 4822 5063
rect 2876 5048 2976 5052
rect 2876 5044 2938 5048
rect 2876 5018 2883 5044
rect 2909 5022 2938 5044
rect 2964 5022 2976 5048
rect 2909 5018 2976 5022
rect 2876 5015 2976 5018
rect 3044 5015 3079 5052
rect 3141 5049 3500 5052
rect 3141 5044 3363 5049
rect 3141 5020 3154 5044
rect 3178 5025 3363 5044
rect 3387 5025 3500 5049
rect 3178 5020 3500 5025
rect 3141 5016 3500 5020
rect 3567 5044 3716 5052
rect 3567 5024 3578 5044
rect 3598 5024 3716 5044
rect 3567 5017 3716 5024
rect 4156 5021 4670 5022
rect 3567 5016 3608 5017
rect 2891 4963 2928 4964
rect 2987 4963 3024 4964
rect 3043 4963 3079 5015
rect 3098 4963 3135 4964
rect 2791 4954 2929 4963
rect 2791 4934 2900 4954
rect 2920 4934 2929 4954
rect 2791 4927 2929 4934
rect 2987 4954 3135 4963
rect 2987 4934 2996 4954
rect 3016 4934 3106 4954
rect 3126 4934 3135 4954
rect 2791 4925 2887 4927
rect 2987 4924 3135 4934
rect 3194 4954 3231 4964
rect 3306 4963 3343 4964
rect 3287 4961 3343 4963
rect 3194 4934 3202 4954
rect 3222 4934 3231 4954
rect 3043 4923 3079 4924
rect 1973 4871 2141 4873
rect 1695 4865 2141 4871
rect 763 4841 1179 4846
rect 1358 4844 1469 4850
rect 763 4840 1104 4841
rect 707 4780 738 4781
rect 555 4750 564 4770
rect 584 4750 592 4770
rect 555 4740 592 4750
rect 651 4773 738 4780
rect 651 4770 712 4773
rect 651 4750 660 4770
rect 680 4753 712 4770
rect 733 4753 738 4773
rect 680 4750 738 4753
rect 651 4743 738 4750
rect 763 4770 800 4840
rect 1066 4839 1103 4840
rect 1358 4836 1399 4844
rect 1358 4816 1366 4836
rect 1385 4816 1399 4836
rect 1358 4814 1399 4816
rect 1427 4836 1469 4844
rect 1427 4816 1443 4836
rect 1462 4816 1469 4836
rect 1695 4843 1701 4865
rect 1727 4845 2141 4865
rect 2891 4864 2928 4865
rect 3194 4864 3231 4934
rect 3256 4954 3343 4961
rect 3256 4951 3314 4954
rect 3256 4931 3261 4951
rect 3282 4934 3314 4951
rect 3334 4934 3343 4954
rect 3282 4931 3343 4934
rect 3256 4924 3343 4931
rect 3402 4954 3439 4964
rect 3402 4934 3410 4954
rect 3430 4934 3439 4954
rect 3256 4923 3287 4924
rect 2890 4863 3231 4864
rect 1727 4843 1736 4845
rect 1973 4844 2141 4845
rect 2815 4858 3231 4863
rect 1695 4834 1736 4843
rect 2815 4838 2818 4858
rect 2838 4838 3231 4858
rect 3402 4855 3439 4934
rect 3469 4963 3500 5016
rect 4137 5005 4670 5021
rect 4137 4994 4669 5005
rect 4788 4996 4825 5000
rect 3519 4963 3556 4964
rect 3469 4954 3556 4963
rect 3469 4934 3527 4954
rect 3547 4934 3556 4954
rect 3469 4924 3556 4934
rect 3615 4954 3652 4964
rect 3615 4934 3623 4954
rect 3643 4934 3652 4954
rect 3469 4923 3500 4924
rect 3464 4855 3574 4868
rect 3615 4855 3652 4934
rect 3402 4853 3652 4855
rect 3402 4850 3503 4853
rect 3402 4831 3467 4850
rect 3464 4823 3467 4831
rect 3496 4823 3503 4850
rect 3531 4826 3541 4853
rect 3570 4831 3652 4853
rect 3730 4925 3898 4926
rect 4137 4925 4175 4994
rect 3730 4905 4175 4925
rect 4402 4956 4513 4971
rect 4402 4954 4444 4956
rect 4402 4934 4409 4954
rect 4428 4934 4444 4954
rect 4402 4926 4444 4934
rect 4472 4954 4513 4956
rect 4472 4934 4486 4954
rect 4505 4934 4513 4954
rect 4472 4926 4513 4934
rect 4402 4920 4513 4926
rect 4635 4931 4669 4994
rect 4787 4990 4825 4996
rect 4787 4972 4797 4990
rect 4815 4972 4825 4990
rect 4787 4963 4825 4972
rect 4787 4931 4821 4963
rect 3730 4899 4174 4905
rect 3730 4897 3898 4899
rect 3570 4826 3574 4831
rect 3531 4823 3574 4826
rect 1427 4814 1469 4816
rect 1358 4799 1469 4814
rect 2554 4805 2602 4819
rect 3464 4809 3574 4823
rect 915 4780 951 4781
rect 763 4750 772 4770
rect 792 4750 800 4770
rect 651 4741 707 4743
rect 651 4740 688 4741
rect 763 4740 800 4750
rect 859 4770 1007 4780
rect 1107 4777 1203 4779
rect 859 4750 868 4770
rect 888 4750 978 4770
rect 998 4750 1007 4770
rect 859 4741 1007 4750
rect 1065 4770 1203 4777
rect 1065 4750 1074 4770
rect 1094 4750 1203 4770
rect 1065 4741 1203 4750
rect 2554 4765 2567 4805
rect 2594 4765 2602 4805
rect 2554 4747 2602 4765
rect 859 4740 896 4741
rect 915 4689 951 4741
rect 970 4740 1007 4741
rect 1066 4740 1103 4741
rect 386 4687 427 4688
rect 278 4680 427 4687
rect 278 4660 396 4680
rect 416 4660 427 4680
rect 278 4652 427 4660
rect 494 4684 853 4688
rect 494 4679 816 4684
rect 494 4655 607 4679
rect 631 4660 816 4679
rect 840 4660 853 4684
rect 631 4655 853 4660
rect 494 4652 853 4655
rect 915 4652 950 4689
rect 1018 4686 1118 4689
rect 1018 4682 1085 4686
rect 1018 4656 1030 4682
rect 1056 4660 1085 4682
rect 1111 4660 1118 4686
rect 1056 4656 1118 4660
rect 1018 4652 1118 4656
rect 494 4631 525 4652
rect 915 4631 951 4652
rect 337 4630 374 4631
rect 336 4621 374 4630
rect 336 4601 345 4621
rect 365 4601 374 4621
rect 336 4593 374 4601
rect 440 4625 525 4631
rect 550 4630 587 4631
rect 440 4605 448 4625
rect 468 4605 525 4625
rect 440 4597 525 4605
rect 549 4621 587 4630
rect 549 4601 558 4621
rect 578 4601 587 4621
rect 440 4596 476 4597
rect 549 4593 587 4601
rect 653 4625 738 4631
rect 758 4630 795 4631
rect 653 4605 661 4625
rect 681 4624 738 4625
rect 681 4605 710 4624
rect 653 4604 710 4605
rect 731 4604 738 4624
rect 653 4597 738 4604
rect 757 4621 795 4630
rect 757 4601 766 4621
rect 786 4601 795 4621
rect 653 4596 689 4597
rect 757 4593 795 4601
rect 861 4625 1005 4631
rect 861 4605 869 4625
rect 889 4622 977 4625
rect 889 4605 920 4622
rect 861 4602 920 4605
rect 943 4605 977 4622
rect 997 4605 1005 4625
rect 943 4602 1005 4605
rect 861 4597 1005 4602
rect 861 4596 897 4597
rect 969 4596 1005 4597
rect 1071 4630 1108 4631
rect 1071 4629 1109 4630
rect 1071 4621 1135 4629
rect 1071 4601 1080 4621
rect 1100 4607 1135 4621
rect 1155 4607 1158 4627
rect 1100 4602 1158 4607
rect 1100 4601 1135 4602
rect 337 4564 374 4593
rect 338 4562 374 4564
rect 550 4562 587 4593
rect 338 4540 587 4562
rect 758 4561 795 4593
rect 1071 4589 1135 4601
rect 1175 4563 1202 4741
rect 2549 4640 2602 4747
rect 3730 4719 3757 4897
rect 3797 4859 3861 4871
rect 4137 4867 4174 4899
rect 4345 4898 4594 4920
rect 4635 4899 4821 4931
rect 4649 4898 4821 4899
rect 4345 4867 4382 4898
rect 4558 4896 4594 4898
rect 4558 4867 4595 4896
rect 4787 4870 4821 4898
rect 3797 4858 3832 4859
rect 3774 4853 3832 4858
rect 3774 4833 3777 4853
rect 3797 4839 3832 4853
rect 3852 4839 3861 4859
rect 3797 4831 3861 4839
rect 3823 4830 3861 4831
rect 3824 4829 3861 4830
rect 3927 4863 3963 4864
rect 4035 4863 4071 4864
rect 3927 4856 4071 4863
rect 3927 4855 3987 4856
rect 3927 4835 3935 4855
rect 3955 4836 3987 4855
rect 4012 4855 4071 4856
rect 4012 4836 4043 4855
rect 3955 4835 4043 4836
rect 4063 4835 4071 4855
rect 3927 4829 4071 4835
rect 4137 4859 4175 4867
rect 4243 4863 4279 4864
rect 4137 4839 4146 4859
rect 4166 4839 4175 4859
rect 4137 4830 4175 4839
rect 4194 4856 4279 4863
rect 4194 4836 4201 4856
rect 4222 4855 4279 4856
rect 4222 4836 4251 4855
rect 4194 4835 4251 4836
rect 4271 4835 4279 4855
rect 4137 4829 4174 4830
rect 4194 4829 4279 4835
rect 4345 4859 4383 4867
rect 4456 4863 4492 4864
rect 4345 4839 4354 4859
rect 4374 4839 4383 4859
rect 4345 4830 4383 4839
rect 4407 4855 4492 4863
rect 4407 4835 4464 4855
rect 4484 4835 4492 4855
rect 4345 4829 4382 4830
rect 4407 4829 4492 4835
rect 4558 4859 4596 4867
rect 4558 4839 4567 4859
rect 4587 4839 4596 4859
rect 4558 4830 4596 4839
rect 4785 4860 4822 4870
rect 4785 4842 4795 4860
rect 4813 4842 4822 4860
rect 4785 4833 4822 4842
rect 4787 4832 4821 4833
rect 4558 4829 4595 4830
rect 3981 4808 4017 4829
rect 4407 4808 4438 4829
rect 3814 4804 3914 4808
rect 3814 4800 3876 4804
rect 3814 4774 3821 4800
rect 3847 4778 3876 4800
rect 3902 4778 3914 4804
rect 3847 4774 3914 4778
rect 3814 4771 3914 4774
rect 3982 4771 4017 4808
rect 4079 4805 4438 4808
rect 4079 4800 4301 4805
rect 4079 4776 4092 4800
rect 4116 4781 4301 4800
rect 4325 4781 4438 4805
rect 4116 4776 4438 4781
rect 4079 4772 4438 4776
rect 4505 4800 4654 4808
rect 4505 4780 4516 4800
rect 4536 4780 4654 4800
rect 4505 4773 4654 4780
rect 4505 4772 4546 4773
rect 3829 4719 3866 4720
rect 3925 4719 3962 4720
rect 3981 4719 4017 4771
rect 4036 4719 4073 4720
rect 3729 4710 3867 4719
rect 3729 4690 3838 4710
rect 3858 4690 3867 4710
rect 3355 4670 3466 4685
rect 3729 4683 3867 4690
rect 3925 4710 4073 4719
rect 3925 4690 3934 4710
rect 3954 4690 4044 4710
rect 4064 4690 4073 4710
rect 3729 4681 3825 4683
rect 3925 4680 4073 4690
rect 4132 4710 4169 4720
rect 4244 4719 4281 4720
rect 4225 4717 4281 4719
rect 4132 4690 4140 4710
rect 4160 4690 4169 4710
rect 3981 4679 4017 4680
rect 3355 4668 3397 4670
rect 3355 4648 3362 4668
rect 3381 4648 3397 4668
rect 3355 4640 3397 4648
rect 3425 4668 3466 4670
rect 3425 4648 3439 4668
rect 3458 4648 3466 4668
rect 3425 4640 3466 4648
rect 2549 4639 2851 4640
rect 1468 4618 1578 4632
rect 1468 4615 1511 4618
rect 1468 4610 1472 4615
rect 1034 4561 1202 4563
rect 758 4558 1202 4561
rect 419 4534 530 4540
rect 419 4526 460 4534
rect 108 4471 147 4515
rect 419 4506 427 4526
rect 446 4506 460 4526
rect 419 4504 460 4506
rect 488 4526 530 4534
rect 488 4506 504 4526
rect 523 4506 530 4526
rect 488 4505 530 4506
rect 756 4535 1202 4558
rect 488 4504 531 4505
rect 419 4485 531 4504
rect 108 4447 148 4471
rect 448 4447 495 4448
rect 756 4447 794 4535
rect 1034 4534 1202 4535
rect 1390 4588 1472 4610
rect 1501 4588 1511 4615
rect 1539 4591 1546 4618
rect 1575 4610 1578 4618
rect 2549 4613 3127 4639
rect 3355 4634 3466 4640
rect 2549 4611 2851 4613
rect 2549 4610 2735 4611
rect 1575 4591 1640 4610
rect 1539 4588 1640 4591
rect 1390 4586 1640 4588
rect 1390 4507 1427 4586
rect 1468 4573 1578 4586
rect 1542 4517 1573 4518
rect 1390 4487 1399 4507
rect 1419 4487 1427 4507
rect 1390 4477 1427 4487
rect 1486 4507 1573 4517
rect 1486 4487 1495 4507
rect 1515 4487 1573 4507
rect 1486 4478 1573 4487
rect 1486 4477 1523 4478
rect 108 4437 794 4447
rect 104 4414 794 4437
rect 1542 4425 1573 4478
rect 1603 4507 1640 4586
rect 1811 4583 2204 4603
rect 2224 4583 2227 4603
rect 2549 4602 2602 4610
rect 1811 4578 2227 4583
rect 1811 4577 2152 4578
rect 1755 4517 1786 4518
rect 1603 4487 1612 4507
rect 1632 4487 1640 4507
rect 1603 4477 1640 4487
rect 1699 4510 1786 4517
rect 1699 4507 1760 4510
rect 1699 4487 1708 4507
rect 1728 4490 1760 4507
rect 1781 4490 1786 4510
rect 1728 4487 1786 4490
rect 1699 4480 1786 4487
rect 1811 4507 1848 4577
rect 2114 4576 2151 4577
rect 1963 4517 1999 4518
rect 1811 4487 1820 4507
rect 1840 4487 1848 4507
rect 1699 4478 1755 4480
rect 1699 4477 1736 4478
rect 1811 4477 1848 4487
rect 1907 4507 2055 4517
rect 2155 4514 2251 4516
rect 1907 4487 1916 4507
rect 1936 4487 2026 4507
rect 2046 4487 2055 4507
rect 1907 4478 2055 4487
rect 2113 4507 2251 4514
rect 2113 4487 2122 4507
rect 2142 4487 2251 4507
rect 2113 4478 2251 4487
rect 1907 4477 1944 4478
rect 1963 4426 1999 4478
rect 2018 4477 2055 4478
rect 2114 4477 2151 4478
rect 1434 4424 1475 4425
rect 104 4395 146 4414
rect 756 4412 794 4414
rect 1326 4417 1475 4424
rect 107 4357 146 4395
rect 1326 4397 1444 4417
rect 1464 4397 1475 4417
rect 1326 4389 1475 4397
rect 1542 4421 1901 4425
rect 1542 4416 1864 4421
rect 1542 4392 1655 4416
rect 1679 4397 1864 4416
rect 1888 4397 1901 4421
rect 1679 4392 1901 4397
rect 1542 4389 1901 4392
rect 1963 4389 1998 4426
rect 2066 4423 2166 4426
rect 2066 4419 2133 4423
rect 2066 4393 2078 4419
rect 2104 4397 2133 4419
rect 2159 4397 2166 4423
rect 2104 4393 2166 4397
rect 2066 4389 2166 4393
rect 1542 4368 1573 4389
rect 1963 4368 1999 4389
rect 1385 4367 1422 4368
rect 1384 4358 1422 4367
rect 107 4355 155 4357
rect 107 4337 118 4355
rect 136 4337 155 4355
rect 107 4328 155 4337
rect 108 4327 155 4328
rect 421 4332 531 4346
rect 421 4329 464 4332
rect 421 4324 425 4329
rect 343 4302 425 4324
rect 454 4302 464 4329
rect 492 4305 499 4332
rect 528 4324 531 4332
rect 1384 4338 1393 4358
rect 1413 4338 1422 4358
rect 1384 4330 1422 4338
rect 1488 4362 1573 4368
rect 1598 4367 1635 4368
rect 1488 4342 1496 4362
rect 1516 4342 1573 4362
rect 1488 4334 1573 4342
rect 1597 4358 1635 4367
rect 1597 4338 1606 4358
rect 1626 4338 1635 4358
rect 1488 4333 1524 4334
rect 1597 4330 1635 4338
rect 1701 4362 1786 4368
rect 1806 4367 1843 4368
rect 1701 4342 1709 4362
rect 1729 4361 1786 4362
rect 1729 4342 1758 4361
rect 1701 4341 1758 4342
rect 1779 4341 1786 4361
rect 1701 4334 1786 4341
rect 1805 4358 1843 4367
rect 1805 4338 1814 4358
rect 1834 4338 1843 4358
rect 1701 4333 1737 4334
rect 1805 4330 1843 4338
rect 1909 4364 2053 4368
rect 1909 4362 1966 4364
rect 1909 4342 1917 4362
rect 1937 4342 1966 4362
rect 1909 4340 1966 4342
rect 1992 4362 2053 4364
rect 1992 4342 2025 4362
rect 2045 4342 2053 4362
rect 1992 4340 2053 4342
rect 1909 4334 2053 4340
rect 1909 4333 1945 4334
rect 2017 4333 2053 4334
rect 2119 4367 2156 4368
rect 2119 4366 2157 4367
rect 2119 4358 2183 4366
rect 2119 4338 2128 4358
rect 2148 4344 2183 4358
rect 2203 4344 2206 4364
rect 2148 4339 2206 4344
rect 2148 4338 2183 4339
rect 528 4305 593 4324
rect 492 4302 593 4305
rect 343 4300 593 4302
rect 111 4264 148 4265
rect 107 4261 148 4264
rect 107 4256 149 4261
rect 107 4238 120 4256
rect 138 4238 149 4256
rect 107 4224 149 4238
rect 187 4224 234 4228
rect 107 4218 234 4224
rect 107 4189 195 4218
rect 224 4189 234 4218
rect 343 4221 380 4300
rect 421 4287 531 4300
rect 495 4231 526 4232
rect 343 4201 352 4221
rect 372 4201 380 4221
rect 343 4191 380 4201
rect 439 4221 526 4231
rect 439 4201 448 4221
rect 468 4201 526 4221
rect 439 4192 526 4201
rect 439 4191 476 4192
rect 107 4185 234 4189
rect 107 4168 146 4185
rect 187 4184 234 4185
rect 107 4150 118 4168
rect 136 4150 146 4168
rect 107 4141 146 4150
rect 108 4140 145 4141
rect 495 4139 526 4192
rect 556 4221 593 4300
rect 764 4297 1157 4317
rect 1177 4297 1180 4317
rect 1385 4301 1422 4330
rect 764 4292 1180 4297
rect 1386 4299 1422 4301
rect 1598 4299 1635 4330
rect 764 4291 1105 4292
rect 708 4231 739 4232
rect 556 4201 565 4221
rect 585 4201 593 4221
rect 556 4191 593 4201
rect 652 4224 739 4231
rect 652 4221 713 4224
rect 652 4201 661 4221
rect 681 4204 713 4221
rect 734 4204 739 4224
rect 681 4201 739 4204
rect 652 4194 739 4201
rect 764 4221 801 4291
rect 1067 4290 1104 4291
rect 1386 4277 1635 4299
rect 1806 4298 1843 4330
rect 2119 4326 2183 4338
rect 2223 4301 2250 4478
rect 2683 4433 2710 4610
rect 2750 4573 2814 4585
rect 3090 4581 3127 4613
rect 3298 4612 3547 4634
rect 3829 4620 3866 4621
rect 4132 4620 4169 4690
rect 4194 4710 4281 4717
rect 4194 4707 4252 4710
rect 4194 4687 4199 4707
rect 4220 4690 4252 4707
rect 4272 4690 4281 4710
rect 4220 4687 4281 4690
rect 4194 4680 4281 4687
rect 4340 4710 4377 4720
rect 4340 4690 4348 4710
rect 4368 4690 4377 4710
rect 4194 4679 4225 4680
rect 3828 4619 4169 4620
rect 3298 4581 3335 4612
rect 3511 4610 3547 4612
rect 3753 4614 4169 4619
rect 3511 4581 3548 4610
rect 3753 4594 3756 4614
rect 3776 4594 4169 4614
rect 4340 4611 4377 4690
rect 4407 4719 4438 4772
rect 4788 4770 4825 4771
rect 4787 4761 4826 4770
rect 4787 4743 4797 4761
rect 4815 4743 4826 4761
rect 4699 4726 4746 4727
rect 4787 4726 4826 4743
rect 4699 4722 4826 4726
rect 4457 4719 4494 4720
rect 4407 4710 4494 4719
rect 4407 4690 4465 4710
rect 4485 4690 4494 4710
rect 4407 4680 4494 4690
rect 4553 4710 4590 4720
rect 4553 4690 4561 4710
rect 4581 4690 4590 4710
rect 4407 4679 4438 4680
rect 4402 4611 4512 4624
rect 4553 4611 4590 4690
rect 4699 4693 4709 4722
rect 4738 4693 4826 4722
rect 4699 4687 4826 4693
rect 4699 4683 4746 4687
rect 4784 4673 4826 4687
rect 4784 4655 4795 4673
rect 4813 4655 4826 4673
rect 4784 4650 4826 4655
rect 4785 4647 4826 4650
rect 4785 4646 4822 4647
rect 4340 4609 4590 4611
rect 4340 4606 4441 4609
rect 4340 4587 4405 4606
rect 2750 4572 2785 4573
rect 2727 4567 2785 4572
rect 2727 4547 2730 4567
rect 2750 4553 2785 4567
rect 2805 4553 2814 4573
rect 2750 4545 2814 4553
rect 2776 4544 2814 4545
rect 2777 4543 2814 4544
rect 2880 4577 2916 4578
rect 2988 4577 3024 4578
rect 2880 4570 3024 4577
rect 2880 4569 2937 4570
rect 2880 4549 2888 4569
rect 2908 4550 2937 4569
rect 2962 4569 3024 4570
rect 2962 4550 2996 4569
rect 2908 4549 2996 4550
rect 3016 4549 3024 4569
rect 2880 4543 3024 4549
rect 3090 4573 3128 4581
rect 3196 4577 3232 4578
rect 3090 4553 3099 4573
rect 3119 4553 3128 4573
rect 3090 4544 3128 4553
rect 3147 4570 3232 4577
rect 3147 4550 3154 4570
rect 3175 4569 3232 4570
rect 3175 4550 3204 4569
rect 3147 4549 3204 4550
rect 3224 4549 3232 4569
rect 3090 4543 3127 4544
rect 3147 4543 3232 4549
rect 3298 4573 3336 4581
rect 3409 4577 3445 4578
rect 3298 4553 3307 4573
rect 3327 4553 3336 4573
rect 3298 4544 3336 4553
rect 3360 4569 3445 4577
rect 3360 4549 3417 4569
rect 3437 4549 3445 4569
rect 3298 4543 3335 4544
rect 3360 4543 3445 4549
rect 3511 4573 3549 4581
rect 3511 4553 3520 4573
rect 3540 4553 3549 4573
rect 4402 4579 4405 4587
rect 4434 4579 4441 4606
rect 4469 4582 4479 4609
rect 4508 4587 4590 4609
rect 4508 4582 4512 4587
rect 4469 4579 4512 4582
rect 4402 4565 4512 4579
rect 4778 4583 4825 4584
rect 4778 4574 4826 4583
rect 4778 4556 4797 4574
rect 4815 4556 4826 4574
rect 4778 4554 4826 4556
rect 3511 4544 3549 4553
rect 3511 4543 3548 4544
rect 2934 4522 2970 4543
rect 3360 4522 3391 4543
rect 2767 4518 2867 4522
rect 2767 4514 2829 4518
rect 2767 4488 2774 4514
rect 2800 4492 2829 4514
rect 2855 4492 2867 4518
rect 2800 4488 2867 4492
rect 2767 4485 2867 4488
rect 2935 4485 2970 4522
rect 3032 4519 3391 4522
rect 3032 4514 3254 4519
rect 3032 4490 3045 4514
rect 3069 4495 3254 4514
rect 3278 4495 3391 4519
rect 3069 4490 3391 4495
rect 3032 4486 3391 4490
rect 3458 4514 3607 4522
rect 3458 4494 3469 4514
rect 3489 4494 3607 4514
rect 4787 4516 4826 4554
rect 3458 4487 3607 4494
rect 4139 4497 4177 4499
rect 4787 4497 4829 4516
rect 3458 4486 3499 4487
rect 2934 4481 2970 4485
rect 2934 4452 2971 4481
rect 2782 4433 2819 4434
rect 2878 4433 2915 4434
rect 2934 4433 2970 4452
rect 2989 4433 3026 4434
rect 2682 4424 2820 4433
rect 2682 4404 2791 4424
rect 2811 4404 2820 4424
rect 2682 4397 2820 4404
rect 2878 4424 3026 4433
rect 2878 4404 2887 4424
rect 2907 4404 2997 4424
rect 3017 4404 3026 4424
rect 2682 4395 2778 4397
rect 2878 4394 3026 4404
rect 3085 4424 3122 4434
rect 3197 4433 3234 4434
rect 3178 4431 3234 4433
rect 3085 4404 3093 4424
rect 3113 4404 3122 4424
rect 2934 4393 2970 4394
rect 2782 4334 2819 4335
rect 3085 4334 3122 4404
rect 3147 4424 3234 4431
rect 3147 4421 3205 4424
rect 3147 4401 3152 4421
rect 3173 4404 3205 4421
rect 3225 4404 3234 4424
rect 3173 4401 3234 4404
rect 3147 4394 3234 4401
rect 3293 4424 3330 4434
rect 3293 4404 3301 4424
rect 3321 4404 3330 4424
rect 3147 4393 3178 4394
rect 2781 4333 3122 4334
rect 2706 4328 3122 4333
rect 2331 4301 2384 4309
rect 2706 4308 2709 4328
rect 2729 4308 3122 4328
rect 3293 4325 3330 4404
rect 3360 4433 3391 4486
rect 4139 4474 4829 4497
rect 4139 4464 4825 4474
rect 3410 4433 3447 4434
rect 3360 4424 3447 4433
rect 3360 4404 3418 4424
rect 3438 4404 3447 4424
rect 3360 4394 3447 4404
rect 3506 4424 3543 4434
rect 3506 4404 3514 4424
rect 3534 4404 3543 4424
rect 3360 4393 3391 4394
rect 3355 4325 3465 4338
rect 3506 4325 3543 4404
rect 3293 4323 3543 4325
rect 3293 4320 3394 4323
rect 3293 4301 3358 4320
rect 2198 4300 2384 4301
rect 2082 4298 2384 4300
rect 1467 4271 1578 4277
rect 1806 4272 2384 4298
rect 3355 4293 3358 4301
rect 3387 4293 3394 4320
rect 3422 4296 3432 4323
rect 3461 4301 3543 4323
rect 3731 4376 3899 4377
rect 4139 4376 4177 4464
rect 4438 4463 4485 4464
rect 4785 4440 4825 4464
rect 4402 4407 4514 4426
rect 4402 4406 4445 4407
rect 3731 4353 4177 4376
rect 4403 4405 4445 4406
rect 4403 4385 4410 4405
rect 4429 4385 4445 4405
rect 4403 4377 4445 4385
rect 4473 4405 4514 4407
rect 4473 4385 4487 4405
rect 4506 4385 4514 4405
rect 4786 4396 4825 4440
rect 4473 4377 4514 4385
rect 4403 4371 4514 4377
rect 3731 4350 4175 4353
rect 3731 4348 3899 4350
rect 3461 4296 3465 4301
rect 3422 4293 3465 4296
rect 3355 4279 3465 4293
rect 2082 4271 2384 4272
rect 1467 4263 1508 4271
rect 1467 4243 1475 4263
rect 1494 4243 1508 4263
rect 1467 4241 1508 4243
rect 1536 4263 1578 4271
rect 1536 4243 1552 4263
rect 1571 4243 1578 4263
rect 1536 4241 1578 4243
rect 916 4231 952 4232
rect 764 4201 773 4221
rect 793 4201 801 4221
rect 652 4192 708 4194
rect 652 4191 689 4192
rect 764 4191 801 4201
rect 860 4221 1008 4231
rect 1108 4228 1204 4230
rect 860 4201 869 4221
rect 889 4201 979 4221
rect 999 4201 1008 4221
rect 860 4192 1008 4201
rect 1066 4221 1204 4228
rect 1467 4226 1578 4241
rect 1066 4201 1075 4221
rect 1095 4201 1204 4221
rect 1066 4192 1204 4201
rect 860 4191 897 4192
rect 916 4140 952 4192
rect 971 4191 1008 4192
rect 1067 4191 1104 4192
rect 387 4138 428 4139
rect 279 4131 428 4138
rect 279 4111 397 4131
rect 417 4111 428 4131
rect 279 4103 428 4111
rect 495 4135 854 4139
rect 495 4130 817 4135
rect 495 4106 608 4130
rect 632 4111 817 4130
rect 841 4111 854 4135
rect 632 4106 854 4111
rect 495 4103 854 4106
rect 916 4103 951 4140
rect 1019 4137 1119 4140
rect 1019 4133 1086 4137
rect 1019 4107 1031 4133
rect 1057 4111 1086 4133
rect 1112 4111 1119 4137
rect 1057 4107 1119 4111
rect 1019 4103 1119 4107
rect 495 4082 526 4103
rect 916 4082 952 4103
rect 338 4081 375 4082
rect 112 4078 146 4079
rect 111 4069 148 4078
rect 111 4051 120 4069
rect 138 4051 148 4069
rect 111 4041 148 4051
rect 337 4072 375 4081
rect 337 4052 346 4072
rect 366 4052 375 4072
rect 337 4044 375 4052
rect 441 4076 526 4082
rect 551 4081 588 4082
rect 441 4056 449 4076
rect 469 4056 526 4076
rect 441 4048 526 4056
rect 550 4072 588 4081
rect 550 4052 559 4072
rect 579 4052 588 4072
rect 441 4047 477 4048
rect 550 4044 588 4052
rect 654 4076 739 4082
rect 759 4081 796 4082
rect 654 4056 662 4076
rect 682 4075 739 4076
rect 682 4056 711 4075
rect 654 4055 711 4056
rect 732 4055 739 4075
rect 654 4048 739 4055
rect 758 4072 796 4081
rect 758 4052 767 4072
rect 787 4052 796 4072
rect 654 4047 690 4048
rect 758 4044 796 4052
rect 862 4076 1006 4082
rect 862 4056 870 4076
rect 890 4075 978 4076
rect 890 4056 921 4075
rect 862 4055 921 4056
rect 946 4056 978 4075
rect 998 4056 1006 4076
rect 946 4055 1006 4056
rect 862 4048 1006 4055
rect 862 4047 898 4048
rect 970 4047 1006 4048
rect 1072 4081 1109 4082
rect 1072 4080 1110 4081
rect 1072 4072 1136 4080
rect 1072 4052 1081 4072
rect 1101 4058 1136 4072
rect 1156 4058 1159 4078
rect 1101 4053 1159 4058
rect 1101 4052 1136 4053
rect 112 4013 146 4041
rect 338 4015 375 4044
rect 339 4013 375 4015
rect 551 4013 588 4044
rect 112 4012 284 4013
rect 112 3980 298 4012
rect 339 3991 588 4013
rect 759 4012 796 4044
rect 1072 4040 1136 4052
rect 1176 4014 1203 4192
rect 2331 4164 2384 4271
rect 3731 4170 3758 4348
rect 3798 4310 3862 4322
rect 4138 4318 4175 4350
rect 4346 4349 4595 4371
rect 4346 4318 4383 4349
rect 4559 4347 4595 4349
rect 4559 4318 4596 4347
rect 3798 4309 3833 4310
rect 3775 4304 3833 4309
rect 3775 4284 3778 4304
rect 3798 4290 3833 4304
rect 3853 4290 3862 4310
rect 3798 4282 3862 4290
rect 3824 4281 3862 4282
rect 3825 4280 3862 4281
rect 3928 4314 3964 4315
rect 4036 4314 4072 4315
rect 3928 4309 4072 4314
rect 3928 4306 3990 4309
rect 3928 4286 3936 4306
rect 3956 4289 3990 4306
rect 4013 4306 4072 4309
rect 4013 4289 4044 4306
rect 3956 4286 4044 4289
rect 4064 4286 4072 4306
rect 3928 4280 4072 4286
rect 4138 4310 4176 4318
rect 4244 4314 4280 4315
rect 4138 4290 4147 4310
rect 4167 4290 4176 4310
rect 4138 4281 4176 4290
rect 4195 4307 4280 4314
rect 4195 4287 4202 4307
rect 4223 4306 4280 4307
rect 4223 4287 4252 4306
rect 4195 4286 4252 4287
rect 4272 4286 4280 4306
rect 4138 4280 4175 4281
rect 4195 4280 4280 4286
rect 4346 4310 4384 4318
rect 4457 4314 4493 4315
rect 4346 4290 4355 4310
rect 4375 4290 4384 4310
rect 4346 4281 4384 4290
rect 4408 4306 4493 4314
rect 4408 4286 4465 4306
rect 4485 4286 4493 4306
rect 4346 4280 4383 4281
rect 4408 4280 4493 4286
rect 4559 4310 4597 4318
rect 4559 4290 4568 4310
rect 4588 4290 4597 4310
rect 4559 4281 4597 4290
rect 4559 4280 4596 4281
rect 3982 4259 4018 4280
rect 4408 4259 4439 4280
rect 3815 4255 3915 4259
rect 3815 4251 3877 4255
rect 3815 4225 3822 4251
rect 3848 4229 3877 4251
rect 3903 4229 3915 4255
rect 3848 4225 3915 4229
rect 3815 4222 3915 4225
rect 3983 4222 4018 4259
rect 4080 4256 4439 4259
rect 4080 4251 4302 4256
rect 4080 4227 4093 4251
rect 4117 4232 4302 4251
rect 4326 4232 4439 4256
rect 4117 4227 4439 4232
rect 4080 4223 4439 4227
rect 4506 4251 4655 4259
rect 4506 4231 4517 4251
rect 4537 4231 4655 4251
rect 4506 4224 4655 4231
rect 4506 4223 4547 4224
rect 3830 4170 3867 4171
rect 3926 4170 3963 4171
rect 3982 4170 4018 4222
rect 4037 4170 4074 4171
rect 2331 4146 2379 4164
rect 2331 4106 2339 4146
rect 2366 4106 2379 4146
rect 3730 4161 3868 4170
rect 3730 4141 3839 4161
rect 3859 4141 3868 4161
rect 3730 4134 3868 4141
rect 3926 4161 4074 4170
rect 3926 4141 3935 4161
rect 3955 4141 4045 4161
rect 4065 4141 4074 4161
rect 3730 4132 3826 4134
rect 3926 4131 4074 4141
rect 4133 4161 4170 4171
rect 4245 4170 4282 4171
rect 4226 4168 4282 4170
rect 4133 4141 4141 4161
rect 4161 4141 4170 4161
rect 3982 4130 4018 4131
rect 1359 4088 1469 4102
rect 2331 4092 2379 4106
rect 3464 4097 3575 4112
rect 3464 4095 3506 4097
rect 1359 4085 1402 4088
rect 1359 4080 1363 4085
rect 1035 4012 1203 4014
rect 759 4006 1203 4012
rect 112 3948 146 3980
rect 108 3939 146 3948
rect 108 3921 118 3939
rect 136 3921 146 3939
rect 108 3915 146 3921
rect 264 3917 298 3980
rect 420 3985 531 3991
rect 420 3977 461 3985
rect 420 3957 428 3977
rect 447 3957 461 3977
rect 420 3955 461 3957
rect 489 3977 531 3985
rect 489 3957 505 3977
rect 524 3957 531 3977
rect 489 3955 531 3957
rect 420 3940 531 3955
rect 758 3986 1203 4006
rect 758 3917 796 3986
rect 1035 3985 1203 3986
rect 1281 4058 1363 4080
rect 1392 4058 1402 4085
rect 1430 4061 1437 4088
rect 1466 4080 1469 4088
rect 1466 4061 1531 4080
rect 1430 4058 1531 4061
rect 1281 4056 1531 4058
rect 1281 3977 1318 4056
rect 1359 4043 1469 4056
rect 1433 3987 1464 3988
rect 1281 3957 1290 3977
rect 1310 3957 1318 3977
rect 1281 3947 1318 3957
rect 1377 3977 1464 3987
rect 1377 3957 1386 3977
rect 1406 3957 1464 3977
rect 1377 3948 1464 3957
rect 1377 3947 1414 3948
rect 108 3911 145 3915
rect 264 3906 796 3917
rect 263 3890 796 3906
rect 1433 3895 1464 3948
rect 1494 3977 1531 4056
rect 1702 4053 2095 4073
rect 2115 4053 2118 4073
rect 3197 4068 3238 4077
rect 1702 4048 2118 4053
rect 2792 4066 2960 4067
rect 3197 4066 3206 4068
rect 1702 4047 2043 4048
rect 1646 3987 1677 3988
rect 1494 3957 1503 3977
rect 1523 3957 1531 3977
rect 1494 3947 1531 3957
rect 1590 3980 1677 3987
rect 1590 3977 1651 3980
rect 1590 3957 1599 3977
rect 1619 3960 1651 3977
rect 1672 3960 1677 3980
rect 1619 3957 1677 3960
rect 1590 3950 1677 3957
rect 1702 3977 1739 4047
rect 2005 4046 2042 4047
rect 2792 4046 3206 4066
rect 3232 4046 3238 4068
rect 3464 4075 3471 4095
rect 3490 4075 3506 4095
rect 3464 4067 3506 4075
rect 3534 4095 3575 4097
rect 3534 4075 3548 4095
rect 3567 4075 3575 4095
rect 3534 4067 3575 4075
rect 3830 4071 3867 4072
rect 4133 4071 4170 4141
rect 4195 4161 4282 4168
rect 4195 4158 4253 4161
rect 4195 4138 4200 4158
rect 4221 4141 4253 4158
rect 4273 4141 4282 4161
rect 4221 4138 4282 4141
rect 4195 4131 4282 4138
rect 4341 4161 4378 4171
rect 4341 4141 4349 4161
rect 4369 4141 4378 4161
rect 4195 4130 4226 4131
rect 3829 4070 4170 4071
rect 3464 4061 3575 4067
rect 3754 4065 4170 4070
rect 2792 4040 3238 4046
rect 2792 4038 2960 4040
rect 1854 3987 1890 3988
rect 1702 3957 1711 3977
rect 1731 3957 1739 3977
rect 1590 3948 1646 3950
rect 1590 3947 1627 3948
rect 1702 3947 1739 3957
rect 1798 3977 1946 3987
rect 2046 3984 2142 3986
rect 1798 3957 1807 3977
rect 1827 3957 1917 3977
rect 1937 3957 1946 3977
rect 1798 3948 1946 3957
rect 2004 3977 2142 3984
rect 2004 3957 2013 3977
rect 2033 3957 2142 3977
rect 2004 3948 2142 3957
rect 1798 3947 1835 3948
rect 1854 3896 1890 3948
rect 1909 3947 1946 3948
rect 2005 3947 2042 3948
rect 1325 3894 1366 3895
rect 263 3889 777 3890
rect 1217 3887 1366 3894
rect 1217 3867 1335 3887
rect 1355 3867 1366 3887
rect 1217 3859 1366 3867
rect 1433 3891 1792 3895
rect 1433 3886 1755 3891
rect 1433 3862 1546 3886
rect 1570 3867 1755 3886
rect 1779 3867 1792 3891
rect 1570 3862 1792 3867
rect 1433 3859 1792 3862
rect 1854 3859 1889 3896
rect 1957 3893 2057 3896
rect 1957 3889 2024 3893
rect 1957 3863 1969 3889
rect 1995 3867 2024 3889
rect 2050 3867 2057 3893
rect 1995 3863 2057 3867
rect 1957 3859 2057 3863
rect 111 3848 148 3849
rect 109 3840 149 3848
rect 109 3822 120 3840
rect 138 3822 149 3840
rect 1433 3838 1464 3859
rect 1854 3838 1890 3859
rect 1276 3837 1313 3838
rect 109 3774 149 3822
rect 1275 3828 1313 3837
rect 1275 3808 1284 3828
rect 1304 3808 1313 3828
rect 1275 3800 1313 3808
rect 1379 3832 1464 3838
rect 1489 3837 1526 3838
rect 1379 3812 1387 3832
rect 1407 3812 1464 3832
rect 1379 3804 1464 3812
rect 1488 3828 1526 3837
rect 1488 3808 1497 3828
rect 1517 3808 1526 3828
rect 1379 3803 1415 3804
rect 1488 3800 1526 3808
rect 1592 3832 1677 3838
rect 1697 3837 1734 3838
rect 1592 3812 1600 3832
rect 1620 3831 1677 3832
rect 1620 3812 1649 3831
rect 1592 3811 1649 3812
rect 1670 3811 1677 3831
rect 1592 3804 1677 3811
rect 1696 3828 1734 3837
rect 1696 3808 1705 3828
rect 1725 3808 1734 3828
rect 1592 3803 1628 3804
rect 1696 3800 1734 3808
rect 1800 3832 1944 3838
rect 1800 3812 1808 3832
rect 1828 3815 1864 3832
rect 1884 3815 1916 3832
rect 1828 3812 1916 3815
rect 1936 3812 1944 3832
rect 1800 3804 1944 3812
rect 1800 3803 1836 3804
rect 1908 3803 1944 3804
rect 2010 3837 2047 3838
rect 2010 3836 2048 3837
rect 2010 3828 2074 3836
rect 2010 3808 2019 3828
rect 2039 3814 2074 3828
rect 2094 3814 2097 3834
rect 2039 3809 2097 3814
rect 2039 3808 2074 3809
rect 420 3778 530 3792
rect 420 3775 463 3778
rect 109 3767 234 3774
rect 420 3770 424 3775
rect 109 3748 201 3767
rect 226 3748 234 3767
rect 109 3738 234 3748
rect 342 3748 424 3770
rect 453 3748 463 3775
rect 491 3751 498 3778
rect 527 3770 530 3778
rect 1276 3771 1313 3800
rect 527 3751 592 3770
rect 1277 3769 1313 3771
rect 1489 3769 1526 3800
rect 1697 3773 1734 3800
rect 2010 3796 2074 3808
rect 491 3748 592 3751
rect 342 3746 592 3748
rect 109 3718 149 3738
rect 108 3709 149 3718
rect 108 3691 118 3709
rect 136 3691 149 3709
rect 108 3682 149 3691
rect 108 3681 145 3682
rect 342 3667 379 3746
rect 420 3733 530 3746
rect 494 3677 525 3678
rect 342 3647 351 3667
rect 371 3647 379 3667
rect 342 3637 379 3647
rect 438 3667 525 3677
rect 438 3647 447 3667
rect 467 3647 525 3667
rect 438 3638 525 3647
rect 438 3637 475 3638
rect 111 3615 148 3619
rect 108 3610 148 3615
rect 108 3592 120 3610
rect 138 3592 148 3610
rect 108 3412 148 3592
rect 494 3585 525 3638
rect 555 3667 592 3746
rect 763 3743 1156 3763
rect 1176 3743 1179 3763
rect 1277 3747 1526 3769
rect 1695 3768 1736 3773
rect 2114 3770 2141 3948
rect 2792 3860 2819 4038
rect 3197 4035 3238 4040
rect 3407 4039 3656 4061
rect 3754 4045 3757 4065
rect 3777 4045 4170 4065
rect 4341 4062 4378 4141
rect 4408 4170 4439 4223
rect 4785 4216 4825 4396
rect 4785 4198 4795 4216
rect 4813 4198 4825 4216
rect 4785 4193 4825 4198
rect 4785 4189 4822 4193
rect 4458 4170 4495 4171
rect 4408 4161 4495 4170
rect 4408 4141 4466 4161
rect 4486 4141 4495 4161
rect 4408 4131 4495 4141
rect 4554 4161 4591 4171
rect 4554 4141 4562 4161
rect 4582 4141 4591 4161
rect 4408 4130 4439 4131
rect 4403 4062 4513 4075
rect 4554 4062 4591 4141
rect 4788 4126 4825 4127
rect 4784 4117 4825 4126
rect 4784 4099 4797 4117
rect 4815 4099 4825 4117
rect 4784 4090 4825 4099
rect 4784 4070 4824 4090
rect 4341 4060 4591 4062
rect 4341 4057 4442 4060
rect 2859 4000 2923 4012
rect 3199 4008 3236 4035
rect 3407 4008 3444 4039
rect 3620 4037 3656 4039
rect 4341 4038 4406 4057
rect 3620 4008 3657 4037
rect 4403 4030 4406 4038
rect 4435 4030 4442 4057
rect 4470 4033 4480 4060
rect 4509 4038 4591 4060
rect 4699 4060 4824 4070
rect 4699 4041 4707 4060
rect 4732 4041 4824 4060
rect 4509 4033 4513 4038
rect 4699 4034 4824 4041
rect 4470 4030 4513 4033
rect 4403 4016 4513 4030
rect 2859 3999 2894 4000
rect 2836 3994 2894 3999
rect 2836 3974 2839 3994
rect 2859 3980 2894 3994
rect 2914 3980 2923 4000
rect 2859 3972 2923 3980
rect 2885 3971 2923 3972
rect 2886 3970 2923 3971
rect 2989 4004 3025 4005
rect 3097 4004 3133 4005
rect 2989 3996 3133 4004
rect 2989 3976 2997 3996
rect 3017 3976 3105 3996
rect 3125 3976 3133 3996
rect 2989 3970 3133 3976
rect 3199 4000 3237 4008
rect 3305 4004 3341 4005
rect 3199 3980 3208 4000
rect 3228 3980 3237 4000
rect 3199 3971 3237 3980
rect 3256 3997 3341 4004
rect 3256 3977 3263 3997
rect 3284 3996 3341 3997
rect 3284 3977 3313 3996
rect 3256 3976 3313 3977
rect 3333 3976 3341 3996
rect 3199 3970 3236 3971
rect 3256 3970 3341 3976
rect 3407 4000 3445 4008
rect 3518 4004 3554 4005
rect 3407 3980 3416 4000
rect 3436 3980 3445 4000
rect 3407 3971 3445 3980
rect 3469 3996 3554 4004
rect 3469 3976 3526 3996
rect 3546 3976 3554 3996
rect 3407 3970 3444 3971
rect 3469 3970 3554 3976
rect 3620 4000 3658 4008
rect 3620 3980 3629 4000
rect 3649 3980 3658 4000
rect 3620 3971 3658 3980
rect 4784 3986 4824 4034
rect 3620 3970 3657 3971
rect 3043 3949 3079 3970
rect 3469 3949 3500 3970
rect 4784 3968 4795 3986
rect 4813 3968 4824 3986
rect 4784 3960 4824 3968
rect 4785 3959 4822 3960
rect 2876 3945 2976 3949
rect 2876 3941 2938 3945
rect 2876 3915 2883 3941
rect 2909 3919 2938 3941
rect 2964 3919 2976 3945
rect 2909 3915 2976 3919
rect 2876 3912 2976 3915
rect 3044 3912 3079 3949
rect 3141 3946 3500 3949
rect 3141 3941 3363 3946
rect 3141 3917 3154 3941
rect 3178 3922 3363 3941
rect 3387 3922 3500 3946
rect 3178 3917 3500 3922
rect 3141 3913 3500 3917
rect 3567 3941 3716 3949
rect 3567 3921 3578 3941
rect 3598 3921 3716 3941
rect 3567 3914 3716 3921
rect 4156 3918 4670 3919
rect 3567 3913 3608 3914
rect 3043 3877 3079 3912
rect 2891 3860 2928 3861
rect 2987 3860 3024 3861
rect 3043 3860 3050 3877
rect 2791 3851 2929 3860
rect 2791 3831 2900 3851
rect 2920 3831 2929 3851
rect 2791 3824 2929 3831
rect 2987 3851 3050 3860
rect 2987 3831 2996 3851
rect 3016 3836 3050 3851
rect 3071 3860 3079 3877
rect 3098 3860 3135 3861
rect 3071 3851 3135 3860
rect 3071 3836 3106 3851
rect 3016 3831 3106 3836
rect 3126 3831 3135 3851
rect 2791 3822 2887 3824
rect 2987 3821 3135 3831
rect 3194 3851 3231 3861
rect 3306 3860 3343 3861
rect 3287 3858 3343 3860
rect 3194 3831 3202 3851
rect 3222 3831 3231 3851
rect 3043 3820 3079 3821
rect 1973 3768 2141 3770
rect 1695 3762 2141 3768
rect 763 3738 1179 3743
rect 1358 3741 1469 3747
rect 763 3737 1104 3738
rect 707 3677 738 3678
rect 555 3647 564 3667
rect 584 3647 592 3667
rect 555 3637 592 3647
rect 651 3670 738 3677
rect 651 3667 712 3670
rect 651 3647 660 3667
rect 680 3650 712 3667
rect 733 3650 738 3670
rect 680 3647 738 3650
rect 651 3640 738 3647
rect 763 3667 800 3737
rect 1066 3736 1103 3737
rect 1358 3733 1399 3741
rect 1358 3713 1366 3733
rect 1385 3713 1399 3733
rect 1358 3711 1399 3713
rect 1427 3733 1469 3741
rect 1427 3713 1443 3733
rect 1462 3713 1469 3733
rect 1695 3740 1701 3762
rect 1727 3742 2141 3762
rect 2891 3761 2928 3762
rect 3194 3761 3231 3831
rect 3256 3851 3343 3858
rect 3256 3848 3314 3851
rect 3256 3828 3261 3848
rect 3282 3831 3314 3848
rect 3334 3831 3343 3851
rect 3282 3828 3343 3831
rect 3256 3821 3343 3828
rect 3402 3851 3439 3861
rect 3402 3831 3410 3851
rect 3430 3831 3439 3851
rect 3256 3820 3287 3821
rect 2890 3760 3231 3761
rect 1727 3740 1736 3742
rect 1973 3741 2141 3742
rect 2815 3759 3231 3760
rect 2815 3755 3191 3759
rect 1695 3731 1736 3740
rect 2815 3735 2818 3755
rect 2838 3742 3191 3755
rect 3223 3742 3231 3759
rect 2838 3735 3231 3742
rect 3402 3752 3439 3831
rect 3469 3860 3500 3913
rect 4137 3902 4670 3918
rect 4137 3891 4669 3902
rect 4788 3893 4825 3897
rect 3519 3860 3556 3861
rect 3469 3851 3556 3860
rect 3469 3831 3527 3851
rect 3547 3831 3556 3851
rect 3469 3821 3556 3831
rect 3615 3851 3652 3861
rect 3615 3831 3623 3851
rect 3643 3831 3652 3851
rect 3469 3820 3500 3821
rect 3464 3752 3574 3765
rect 3615 3752 3652 3831
rect 3402 3750 3652 3752
rect 3402 3747 3503 3750
rect 3402 3728 3467 3747
rect 1427 3711 1469 3713
rect 1358 3696 1469 3711
rect 3464 3720 3467 3728
rect 3496 3720 3503 3747
rect 3531 3723 3541 3750
rect 3570 3728 3652 3750
rect 3730 3822 3898 3823
rect 4137 3822 4175 3891
rect 3730 3802 4175 3822
rect 4402 3853 4513 3868
rect 4402 3851 4444 3853
rect 4402 3831 4409 3851
rect 4428 3831 4444 3851
rect 4402 3823 4444 3831
rect 4472 3851 4513 3853
rect 4472 3831 4486 3851
rect 4505 3831 4513 3851
rect 4472 3823 4513 3831
rect 4402 3817 4513 3823
rect 4635 3828 4669 3891
rect 4787 3887 4825 3893
rect 4787 3869 4797 3887
rect 4815 3869 4825 3887
rect 4787 3860 4825 3869
rect 4787 3828 4821 3860
rect 3730 3796 4174 3802
rect 3730 3794 3898 3796
rect 3570 3723 3574 3728
rect 3531 3720 3574 3723
rect 3464 3706 3574 3720
rect 915 3677 951 3678
rect 763 3647 772 3667
rect 792 3647 800 3667
rect 651 3638 707 3640
rect 651 3637 688 3638
rect 763 3637 800 3647
rect 859 3667 1007 3677
rect 1107 3674 1203 3676
rect 859 3647 868 3667
rect 888 3647 978 3667
rect 998 3647 1007 3667
rect 859 3638 1007 3647
rect 1065 3667 1203 3674
rect 1065 3647 1074 3667
rect 1094 3647 1203 3667
rect 1065 3638 1203 3647
rect 859 3637 896 3638
rect 915 3586 951 3638
rect 970 3637 1007 3638
rect 1066 3637 1103 3638
rect 386 3584 427 3585
rect 278 3577 427 3584
rect 278 3557 396 3577
rect 416 3557 427 3577
rect 278 3549 427 3557
rect 494 3581 853 3585
rect 494 3576 816 3581
rect 494 3552 607 3576
rect 631 3557 816 3576
rect 840 3557 853 3581
rect 631 3552 853 3557
rect 494 3549 853 3552
rect 915 3549 950 3586
rect 1018 3583 1118 3586
rect 1018 3579 1085 3583
rect 1018 3553 1030 3579
rect 1056 3557 1085 3579
rect 1111 3557 1118 3583
rect 1056 3553 1118 3557
rect 1018 3549 1118 3553
rect 494 3528 525 3549
rect 915 3528 951 3549
rect 337 3527 374 3528
rect 336 3518 374 3527
rect 336 3498 345 3518
rect 365 3498 374 3518
rect 336 3490 374 3498
rect 440 3522 525 3528
rect 550 3527 587 3528
rect 440 3502 448 3522
rect 468 3502 525 3522
rect 440 3494 525 3502
rect 549 3518 587 3527
rect 549 3498 558 3518
rect 578 3498 587 3518
rect 440 3493 476 3494
rect 549 3490 587 3498
rect 653 3522 738 3528
rect 758 3527 795 3528
rect 653 3502 661 3522
rect 681 3521 738 3522
rect 681 3502 710 3521
rect 653 3501 710 3502
rect 731 3501 738 3521
rect 653 3494 738 3501
rect 757 3518 795 3527
rect 757 3498 766 3518
rect 786 3498 795 3518
rect 653 3493 689 3494
rect 757 3490 795 3498
rect 861 3522 1005 3528
rect 861 3502 869 3522
rect 889 3519 977 3522
rect 889 3502 920 3519
rect 861 3499 920 3502
rect 943 3502 977 3519
rect 997 3502 1005 3522
rect 943 3499 1005 3502
rect 861 3494 1005 3499
rect 861 3493 897 3494
rect 969 3493 1005 3494
rect 1071 3527 1108 3528
rect 1071 3526 1109 3527
rect 1071 3518 1135 3526
rect 1071 3498 1080 3518
rect 1100 3504 1135 3518
rect 1155 3504 1158 3524
rect 1100 3499 1158 3504
rect 1100 3498 1135 3499
rect 337 3461 374 3490
rect 338 3459 374 3461
rect 550 3459 587 3490
rect 338 3437 587 3459
rect 758 3458 795 3490
rect 1071 3486 1135 3498
rect 1175 3460 1202 3638
rect 3730 3616 3757 3794
rect 3797 3756 3861 3768
rect 4137 3764 4174 3796
rect 4345 3795 4594 3817
rect 4635 3796 4821 3828
rect 4649 3795 4821 3796
rect 4345 3764 4382 3795
rect 4558 3793 4594 3795
rect 4558 3764 4595 3793
rect 4787 3767 4821 3795
rect 3797 3755 3832 3756
rect 3774 3750 3832 3755
rect 3774 3730 3777 3750
rect 3797 3736 3832 3750
rect 3852 3736 3861 3756
rect 3797 3728 3861 3736
rect 3823 3727 3861 3728
rect 3824 3726 3861 3727
rect 3927 3760 3963 3761
rect 4035 3760 4071 3761
rect 3927 3753 4071 3760
rect 3927 3752 3987 3753
rect 3927 3732 3935 3752
rect 3955 3733 3987 3752
rect 4012 3752 4071 3753
rect 4012 3733 4043 3752
rect 3955 3732 4043 3733
rect 4063 3732 4071 3752
rect 3927 3726 4071 3732
rect 4137 3756 4175 3764
rect 4243 3760 4279 3761
rect 4137 3736 4146 3756
rect 4166 3736 4175 3756
rect 4137 3727 4175 3736
rect 4194 3753 4279 3760
rect 4194 3733 4201 3753
rect 4222 3752 4279 3753
rect 4222 3733 4251 3752
rect 4194 3732 4251 3733
rect 4271 3732 4279 3752
rect 4137 3726 4174 3727
rect 4194 3726 4279 3732
rect 4345 3756 4383 3764
rect 4456 3760 4492 3761
rect 4345 3736 4354 3756
rect 4374 3736 4383 3756
rect 4345 3727 4383 3736
rect 4407 3752 4492 3760
rect 4407 3732 4464 3752
rect 4484 3732 4492 3752
rect 4345 3726 4382 3727
rect 4407 3726 4492 3732
rect 4558 3756 4596 3764
rect 4558 3736 4567 3756
rect 4587 3736 4596 3756
rect 4558 3727 4596 3736
rect 4785 3757 4822 3767
rect 4785 3739 4795 3757
rect 4813 3739 4822 3757
rect 4785 3730 4822 3739
rect 4787 3729 4821 3730
rect 4558 3726 4595 3727
rect 3981 3705 4017 3726
rect 4407 3705 4438 3726
rect 3814 3701 3914 3705
rect 3814 3697 3876 3701
rect 3814 3671 3821 3697
rect 3847 3675 3876 3697
rect 3902 3675 3914 3701
rect 3847 3671 3914 3675
rect 3814 3668 3914 3671
rect 3982 3668 4017 3705
rect 4079 3702 4438 3705
rect 4079 3697 4301 3702
rect 4079 3673 4092 3697
rect 4116 3678 4301 3697
rect 4325 3678 4438 3702
rect 4116 3673 4438 3678
rect 4079 3669 4438 3673
rect 4505 3697 4654 3705
rect 4505 3677 4516 3697
rect 4536 3677 4654 3697
rect 4505 3670 4654 3677
rect 4505 3669 4546 3670
rect 3829 3616 3866 3617
rect 3925 3616 3962 3617
rect 3981 3616 4017 3668
rect 4036 3616 4073 3617
rect 3729 3607 3867 3616
rect 3324 3586 3435 3601
rect 3324 3584 3366 3586
rect 2994 3563 3099 3565
rect 2650 3555 2820 3556
rect 2994 3555 3043 3563
rect 2650 3536 3043 3555
rect 3074 3536 3099 3563
rect 3324 3564 3331 3584
rect 3350 3564 3366 3584
rect 3324 3556 3366 3564
rect 3394 3584 3435 3586
rect 3394 3564 3408 3584
rect 3427 3564 3435 3584
rect 3729 3587 3838 3607
rect 3858 3587 3867 3607
rect 3729 3580 3867 3587
rect 3925 3607 4073 3616
rect 3925 3587 3934 3607
rect 3954 3587 4044 3607
rect 4064 3587 4073 3607
rect 3729 3578 3825 3580
rect 3925 3577 4073 3587
rect 4132 3607 4169 3617
rect 4244 3616 4281 3617
rect 4225 3614 4281 3616
rect 4132 3587 4140 3607
rect 4160 3587 4169 3607
rect 3981 3576 4017 3577
rect 3394 3556 3435 3564
rect 3324 3550 3435 3556
rect 2650 3529 3099 3536
rect 2650 3527 2820 3529
rect 1500 3496 1610 3510
rect 1500 3493 1543 3496
rect 1500 3488 1504 3493
rect 1034 3458 1202 3460
rect 758 3455 1202 3458
rect 419 3431 530 3437
rect 419 3423 460 3431
rect 108 3368 147 3412
rect 419 3403 427 3423
rect 446 3403 460 3423
rect 419 3401 460 3403
rect 488 3423 530 3431
rect 488 3403 504 3423
rect 523 3403 530 3423
rect 488 3401 530 3403
rect 419 3386 530 3401
rect 756 3432 1202 3455
rect 108 3344 148 3368
rect 448 3344 495 3346
rect 756 3344 794 3432
rect 1034 3431 1202 3432
rect 1422 3466 1504 3488
rect 1533 3466 1543 3493
rect 1571 3469 1578 3496
rect 1607 3488 1610 3496
rect 1607 3469 1672 3488
rect 1571 3466 1672 3469
rect 1422 3464 1672 3466
rect 1422 3385 1459 3464
rect 1500 3451 1610 3464
rect 1574 3395 1605 3396
rect 1422 3365 1431 3385
rect 1451 3365 1459 3385
rect 1422 3355 1459 3365
rect 1518 3385 1605 3395
rect 1518 3365 1527 3385
rect 1547 3365 1605 3385
rect 1518 3356 1605 3365
rect 1518 3355 1555 3356
rect 108 3311 794 3344
rect 108 3254 147 3311
rect 756 3309 794 3311
rect 1574 3303 1605 3356
rect 1635 3385 1672 3464
rect 1843 3477 2236 3481
rect 1843 3460 1862 3477
rect 1882 3461 2236 3477
rect 2256 3461 2259 3481
rect 1882 3460 2259 3461
rect 1843 3456 2259 3460
rect 1843 3455 2184 3456
rect 1787 3395 1818 3396
rect 1635 3365 1644 3385
rect 1664 3365 1672 3385
rect 1635 3355 1672 3365
rect 1731 3388 1818 3395
rect 1731 3385 1792 3388
rect 1731 3365 1740 3385
rect 1760 3368 1792 3385
rect 1813 3368 1818 3388
rect 1760 3365 1818 3368
rect 1731 3358 1818 3365
rect 1843 3385 1880 3455
rect 2146 3454 2183 3455
rect 1995 3395 2031 3396
rect 1843 3365 1852 3385
rect 1872 3365 1880 3385
rect 1731 3356 1787 3358
rect 1731 3355 1768 3356
rect 1843 3355 1880 3365
rect 1939 3385 2087 3395
rect 2187 3392 2283 3394
rect 1939 3365 1948 3385
rect 1968 3365 2058 3385
rect 2078 3365 2087 3385
rect 1939 3356 2087 3365
rect 2145 3385 2283 3392
rect 2145 3365 2154 3385
rect 2174 3365 2283 3385
rect 2145 3356 2283 3365
rect 1939 3355 1976 3356
rect 1995 3304 2031 3356
rect 2050 3355 2087 3356
rect 2146 3355 2183 3356
rect 1466 3302 1507 3303
rect 1358 3295 1507 3302
rect 1358 3275 1476 3295
rect 1496 3275 1507 3295
rect 1358 3267 1507 3275
rect 1574 3299 1933 3303
rect 1574 3294 1896 3299
rect 1574 3270 1687 3294
rect 1711 3275 1896 3294
rect 1920 3275 1933 3299
rect 1711 3270 1933 3275
rect 1574 3267 1933 3270
rect 1995 3267 2030 3304
rect 2098 3301 2198 3304
rect 2098 3297 2165 3301
rect 2098 3271 2110 3297
rect 2136 3275 2165 3297
rect 2191 3275 2198 3301
rect 2136 3271 2198 3275
rect 2098 3267 2198 3271
rect 108 3252 156 3254
rect 108 3234 119 3252
rect 137 3234 156 3252
rect 1574 3246 1605 3267
rect 1995 3246 2031 3267
rect 1417 3245 1454 3246
rect 108 3225 156 3234
rect 109 3224 156 3225
rect 422 3229 532 3243
rect 422 3226 465 3229
rect 422 3221 426 3226
rect 344 3199 426 3221
rect 455 3199 465 3226
rect 493 3202 500 3229
rect 529 3221 532 3229
rect 1416 3236 1454 3245
rect 529 3202 594 3221
rect 1416 3216 1425 3236
rect 1445 3216 1454 3236
rect 493 3199 594 3202
rect 344 3197 594 3199
rect 112 3161 149 3162
rect 108 3158 149 3161
rect 108 3153 150 3158
rect 108 3135 121 3153
rect 139 3135 150 3153
rect 108 3121 150 3135
rect 188 3121 235 3125
rect 108 3115 235 3121
rect 108 3086 196 3115
rect 225 3086 235 3115
rect 344 3118 381 3197
rect 422 3184 532 3197
rect 496 3128 527 3129
rect 344 3098 353 3118
rect 373 3098 381 3118
rect 344 3088 381 3098
rect 440 3118 527 3128
rect 440 3098 449 3118
rect 469 3098 527 3118
rect 440 3089 527 3098
rect 440 3088 477 3089
rect 108 3082 235 3086
rect 108 3065 147 3082
rect 188 3081 235 3082
rect 108 3047 119 3065
rect 137 3047 147 3065
rect 108 3038 147 3047
rect 109 3037 146 3038
rect 496 3036 527 3089
rect 557 3118 594 3197
rect 765 3194 1158 3214
rect 1178 3194 1181 3214
rect 1416 3208 1454 3216
rect 1520 3240 1605 3246
rect 1630 3245 1667 3246
rect 1520 3220 1528 3240
rect 1548 3220 1605 3240
rect 1520 3212 1605 3220
rect 1629 3236 1667 3245
rect 1629 3216 1638 3236
rect 1658 3216 1667 3236
rect 1520 3211 1556 3212
rect 1629 3208 1667 3216
rect 1733 3240 1818 3246
rect 1838 3245 1875 3246
rect 1733 3220 1741 3240
rect 1761 3239 1818 3240
rect 1761 3220 1790 3239
rect 1733 3219 1790 3220
rect 1811 3219 1818 3239
rect 1733 3212 1818 3219
rect 1837 3236 1875 3245
rect 1837 3216 1846 3236
rect 1866 3216 1875 3236
rect 1733 3211 1769 3212
rect 1837 3208 1875 3216
rect 1941 3240 2085 3246
rect 1941 3220 1949 3240
rect 1969 3238 2057 3240
rect 1969 3220 1998 3238
rect 1941 3217 1998 3220
rect 2025 3220 2057 3238
rect 2077 3220 2085 3240
rect 2025 3217 2085 3220
rect 1941 3212 2085 3217
rect 1941 3211 1977 3212
rect 2049 3211 2085 3212
rect 2151 3245 2188 3246
rect 2151 3244 2189 3245
rect 2151 3236 2215 3244
rect 2151 3216 2160 3236
rect 2180 3222 2215 3236
rect 2235 3222 2238 3242
rect 2180 3217 2238 3222
rect 2180 3216 2215 3217
rect 765 3189 1181 3194
rect 765 3188 1106 3189
rect 709 3128 740 3129
rect 557 3098 566 3118
rect 586 3098 594 3118
rect 557 3088 594 3098
rect 653 3121 740 3128
rect 653 3118 714 3121
rect 653 3098 662 3118
rect 682 3101 714 3118
rect 735 3101 740 3121
rect 682 3098 740 3101
rect 653 3091 740 3098
rect 765 3118 802 3188
rect 1068 3187 1105 3188
rect 1417 3179 1454 3208
rect 1418 3177 1454 3179
rect 1630 3177 1667 3208
rect 1418 3155 1667 3177
rect 1838 3176 1875 3208
rect 2151 3204 2215 3216
rect 2255 3178 2282 3356
rect 2650 3349 2679 3527
rect 2719 3489 2783 3501
rect 3059 3497 3096 3529
rect 3267 3528 3516 3550
rect 3267 3497 3304 3528
rect 3480 3526 3516 3528
rect 3480 3497 3517 3526
rect 3829 3517 3866 3518
rect 4132 3517 4169 3587
rect 4194 3607 4281 3614
rect 4194 3604 4252 3607
rect 4194 3584 4199 3604
rect 4220 3587 4252 3604
rect 4272 3587 4281 3607
rect 4220 3584 4281 3587
rect 4194 3577 4281 3584
rect 4340 3607 4377 3617
rect 4340 3587 4348 3607
rect 4368 3587 4377 3607
rect 4194 3576 4225 3577
rect 3828 3516 4169 3517
rect 3753 3511 4169 3516
rect 2719 3488 2754 3489
rect 2696 3483 2754 3488
rect 2696 3463 2699 3483
rect 2719 3469 2754 3483
rect 2774 3469 2783 3489
rect 2719 3461 2783 3469
rect 2745 3460 2783 3461
rect 2746 3459 2783 3460
rect 2849 3493 2885 3494
rect 2957 3493 2993 3494
rect 2849 3485 2993 3493
rect 2849 3465 2857 3485
rect 2877 3465 2965 3485
rect 2985 3465 2993 3485
rect 2849 3459 2993 3465
rect 3059 3489 3097 3497
rect 3165 3493 3201 3494
rect 3059 3469 3068 3489
rect 3088 3469 3097 3489
rect 3059 3460 3097 3469
rect 3116 3486 3201 3493
rect 3116 3466 3123 3486
rect 3144 3485 3201 3486
rect 3144 3466 3173 3485
rect 3116 3465 3173 3466
rect 3193 3465 3201 3485
rect 3059 3459 3096 3460
rect 3116 3459 3201 3465
rect 3267 3489 3305 3497
rect 3378 3493 3414 3494
rect 3267 3469 3276 3489
rect 3296 3469 3305 3489
rect 3267 3460 3305 3469
rect 3329 3485 3414 3493
rect 3329 3465 3386 3485
rect 3406 3465 3414 3485
rect 3267 3459 3304 3460
rect 3329 3459 3414 3465
rect 3480 3489 3518 3497
rect 3753 3491 3756 3511
rect 3776 3491 4169 3511
rect 4340 3508 4377 3587
rect 4407 3616 4438 3669
rect 4788 3667 4825 3668
rect 4787 3658 4826 3667
rect 4787 3640 4797 3658
rect 4815 3640 4826 3658
rect 4699 3623 4746 3624
rect 4787 3623 4826 3640
rect 4699 3619 4826 3623
rect 4457 3616 4494 3617
rect 4407 3607 4494 3616
rect 4407 3587 4465 3607
rect 4485 3587 4494 3607
rect 4407 3577 4494 3587
rect 4553 3607 4590 3617
rect 4553 3587 4561 3607
rect 4581 3587 4590 3607
rect 4407 3576 4438 3577
rect 4402 3508 4512 3521
rect 4553 3508 4590 3587
rect 4699 3590 4709 3619
rect 4738 3590 4826 3619
rect 4699 3584 4826 3590
rect 4699 3580 4746 3584
rect 4784 3570 4826 3584
rect 4784 3552 4795 3570
rect 4813 3552 4826 3570
rect 4784 3547 4826 3552
rect 4785 3544 4826 3547
rect 4785 3543 4822 3544
rect 4340 3506 4590 3508
rect 4340 3503 4441 3506
rect 3480 3469 3489 3489
rect 3509 3469 3518 3489
rect 4340 3484 4405 3503
rect 3480 3460 3518 3469
rect 4402 3476 4405 3484
rect 4434 3476 4441 3503
rect 4469 3479 4479 3506
rect 4508 3484 4590 3506
rect 4508 3479 4512 3484
rect 4469 3476 4512 3479
rect 4402 3462 4512 3476
rect 4778 3480 4825 3481
rect 4778 3471 4826 3480
rect 3480 3459 3517 3460
rect 2903 3438 2939 3459
rect 3329 3438 3360 3459
rect 4778 3453 4797 3471
rect 4815 3453 4826 3471
rect 4778 3451 4826 3453
rect 2736 3434 2836 3438
rect 2736 3430 2798 3434
rect 2736 3404 2743 3430
rect 2769 3408 2798 3430
rect 2824 3408 2836 3434
rect 2769 3404 2836 3408
rect 2736 3401 2836 3404
rect 2904 3401 2939 3438
rect 3001 3435 3360 3438
rect 3001 3430 3223 3435
rect 3001 3406 3014 3430
rect 3038 3411 3223 3430
rect 3247 3411 3360 3435
rect 3038 3406 3360 3411
rect 3001 3402 3360 3406
rect 3427 3430 3576 3438
rect 3427 3410 3438 3430
rect 3458 3410 3576 3430
rect 3427 3403 3576 3410
rect 3427 3402 3468 3403
rect 2903 3362 2939 3401
rect 2751 3349 2788 3350
rect 2847 3349 2884 3350
rect 2903 3349 2910 3362
rect 2650 3340 2789 3349
rect 2650 3320 2760 3340
rect 2780 3320 2789 3340
rect 2650 3313 2789 3320
rect 2847 3340 2910 3349
rect 2847 3320 2856 3340
rect 2876 3324 2910 3340
rect 2933 3349 2939 3362
rect 2958 3349 2995 3350
rect 2933 3340 2995 3349
rect 2933 3324 2966 3340
rect 2876 3320 2966 3324
rect 2986 3320 2995 3340
rect 2650 3311 2747 3313
rect 2650 3310 2679 3311
rect 2847 3310 2995 3320
rect 3054 3340 3091 3350
rect 3166 3349 3203 3350
rect 3147 3347 3203 3349
rect 3054 3320 3062 3340
rect 3082 3320 3091 3340
rect 2903 3309 2939 3310
rect 2751 3250 2788 3251
rect 3054 3250 3091 3320
rect 3116 3340 3203 3347
rect 3116 3337 3174 3340
rect 3116 3317 3121 3337
rect 3142 3320 3174 3337
rect 3194 3320 3203 3340
rect 3142 3317 3203 3320
rect 3116 3310 3203 3317
rect 3262 3340 3299 3350
rect 3262 3320 3270 3340
rect 3290 3320 3299 3340
rect 3116 3309 3147 3310
rect 2750 3249 3091 3250
rect 2675 3245 3091 3249
rect 2675 3244 3052 3245
rect 2675 3224 2678 3244
rect 2698 3228 3052 3244
rect 3072 3228 3091 3245
rect 2698 3224 3091 3228
rect 3262 3241 3299 3320
rect 3329 3349 3360 3402
rect 4140 3394 4178 3396
rect 4787 3394 4826 3451
rect 4140 3361 4826 3394
rect 3379 3349 3416 3350
rect 3329 3340 3416 3349
rect 3329 3320 3387 3340
rect 3407 3320 3416 3340
rect 3329 3310 3416 3320
rect 3475 3340 3512 3350
rect 3475 3320 3483 3340
rect 3503 3320 3512 3340
rect 3329 3309 3360 3310
rect 3324 3241 3434 3254
rect 3475 3241 3512 3320
rect 3262 3239 3512 3241
rect 3262 3236 3363 3239
rect 3262 3217 3327 3236
rect 3324 3209 3327 3217
rect 3356 3209 3363 3236
rect 3391 3212 3401 3239
rect 3430 3217 3512 3239
rect 3732 3273 3900 3274
rect 4140 3273 4178 3361
rect 4439 3359 4486 3361
rect 4786 3337 4826 3361
rect 3732 3250 4178 3273
rect 4404 3304 4515 3319
rect 4404 3302 4446 3304
rect 4404 3282 4411 3302
rect 4430 3282 4446 3302
rect 4404 3274 4446 3282
rect 4474 3302 4515 3304
rect 4474 3282 4488 3302
rect 4507 3282 4515 3302
rect 4787 3293 4826 3337
rect 4474 3274 4515 3282
rect 4404 3268 4515 3274
rect 3732 3247 4176 3250
rect 3732 3245 3900 3247
rect 3430 3212 3434 3217
rect 3391 3209 3434 3212
rect 3324 3195 3434 3209
rect 2114 3176 2282 3178
rect 1835 3169 2282 3176
rect 1499 3149 1610 3155
rect 1499 3141 1540 3149
rect 917 3128 953 3129
rect 765 3098 774 3118
rect 794 3098 802 3118
rect 653 3089 709 3091
rect 653 3088 690 3089
rect 765 3088 802 3098
rect 861 3118 1009 3128
rect 1109 3125 1205 3127
rect 861 3098 870 3118
rect 890 3098 980 3118
rect 1000 3098 1009 3118
rect 861 3089 1009 3098
rect 1067 3118 1205 3125
rect 1067 3098 1076 3118
rect 1096 3098 1205 3118
rect 1499 3121 1507 3141
rect 1526 3121 1540 3141
rect 1499 3119 1540 3121
rect 1568 3141 1610 3149
rect 1568 3121 1584 3141
rect 1603 3121 1610 3141
rect 1835 3142 1860 3169
rect 1891 3150 2282 3169
rect 1891 3142 1940 3150
rect 2114 3149 2282 3150
rect 1835 3140 1940 3142
rect 1568 3119 1610 3121
rect 1499 3104 1610 3119
rect 1067 3089 1205 3098
rect 861 3088 898 3089
rect 917 3037 953 3089
rect 972 3088 1009 3089
rect 1068 3088 1105 3089
rect 388 3035 429 3036
rect 280 3028 429 3035
rect 280 3008 398 3028
rect 418 3008 429 3028
rect 280 3000 429 3008
rect 496 3032 855 3036
rect 496 3027 818 3032
rect 496 3003 609 3027
rect 633 3008 818 3027
rect 842 3008 855 3032
rect 633 3003 855 3008
rect 496 3000 855 3003
rect 917 3000 952 3037
rect 1020 3034 1120 3037
rect 1020 3030 1087 3034
rect 1020 3004 1032 3030
rect 1058 3008 1087 3030
rect 1113 3008 1120 3034
rect 1058 3004 1120 3008
rect 1020 3000 1120 3004
rect 496 2979 527 3000
rect 917 2979 953 3000
rect 339 2978 376 2979
rect 113 2975 147 2976
rect 112 2966 149 2975
rect 112 2948 121 2966
rect 139 2948 149 2966
rect 112 2938 149 2948
rect 338 2969 376 2978
rect 338 2949 347 2969
rect 367 2949 376 2969
rect 338 2941 376 2949
rect 442 2973 527 2979
rect 552 2978 589 2979
rect 442 2953 450 2973
rect 470 2953 527 2973
rect 442 2945 527 2953
rect 551 2969 589 2978
rect 551 2949 560 2969
rect 580 2949 589 2969
rect 442 2944 478 2945
rect 551 2941 589 2949
rect 655 2973 740 2979
rect 760 2978 797 2979
rect 655 2953 663 2973
rect 683 2972 740 2973
rect 683 2953 712 2972
rect 655 2952 712 2953
rect 733 2952 740 2972
rect 655 2945 740 2952
rect 759 2969 797 2978
rect 759 2949 768 2969
rect 788 2949 797 2969
rect 655 2944 691 2945
rect 759 2941 797 2949
rect 863 2973 1007 2979
rect 863 2953 871 2973
rect 891 2972 979 2973
rect 891 2953 922 2972
rect 863 2952 922 2953
rect 947 2953 979 2972
rect 999 2953 1007 2973
rect 947 2952 1007 2953
rect 863 2945 1007 2952
rect 863 2944 899 2945
rect 971 2944 1007 2945
rect 1073 2978 1110 2979
rect 1073 2977 1111 2978
rect 1073 2969 1137 2977
rect 1073 2949 1082 2969
rect 1102 2955 1137 2969
rect 1157 2955 1160 2975
rect 1102 2950 1160 2955
rect 1102 2949 1137 2950
rect 113 2910 147 2938
rect 339 2912 376 2941
rect 340 2910 376 2912
rect 552 2910 589 2941
rect 113 2909 285 2910
rect 113 2877 299 2909
rect 340 2888 589 2910
rect 760 2909 797 2941
rect 1073 2937 1137 2949
rect 1177 2911 1204 3089
rect 3732 3067 3759 3245
rect 3799 3207 3863 3219
rect 4139 3215 4176 3247
rect 4347 3246 4596 3268
rect 4347 3215 4384 3246
rect 4560 3244 4596 3246
rect 4560 3215 4597 3244
rect 3799 3206 3834 3207
rect 3776 3201 3834 3206
rect 3776 3181 3779 3201
rect 3799 3187 3834 3201
rect 3854 3187 3863 3207
rect 3799 3179 3863 3187
rect 3825 3178 3863 3179
rect 3826 3177 3863 3178
rect 3929 3211 3965 3212
rect 4037 3211 4073 3212
rect 3929 3206 4073 3211
rect 3929 3203 3991 3206
rect 3929 3183 3937 3203
rect 3957 3186 3991 3203
rect 4014 3203 4073 3206
rect 4014 3186 4045 3203
rect 3957 3183 4045 3186
rect 4065 3183 4073 3203
rect 3929 3177 4073 3183
rect 4139 3207 4177 3215
rect 4245 3211 4281 3212
rect 4139 3187 4148 3207
rect 4168 3187 4177 3207
rect 4139 3178 4177 3187
rect 4196 3204 4281 3211
rect 4196 3184 4203 3204
rect 4224 3203 4281 3204
rect 4224 3184 4253 3203
rect 4196 3183 4253 3184
rect 4273 3183 4281 3203
rect 4139 3177 4176 3178
rect 4196 3177 4281 3183
rect 4347 3207 4385 3215
rect 4458 3211 4494 3212
rect 4347 3187 4356 3207
rect 4376 3187 4385 3207
rect 4347 3178 4385 3187
rect 4409 3203 4494 3211
rect 4409 3183 4466 3203
rect 4486 3183 4494 3203
rect 4347 3177 4384 3178
rect 4409 3177 4494 3183
rect 4560 3207 4598 3215
rect 4560 3187 4569 3207
rect 4589 3187 4598 3207
rect 4560 3178 4598 3187
rect 4560 3177 4597 3178
rect 3983 3156 4019 3177
rect 4409 3156 4440 3177
rect 3816 3152 3916 3156
rect 3816 3148 3878 3152
rect 3816 3122 3823 3148
rect 3849 3126 3878 3148
rect 3904 3126 3916 3152
rect 3849 3122 3916 3126
rect 3816 3119 3916 3122
rect 3984 3119 4019 3156
rect 4081 3153 4440 3156
rect 4081 3148 4303 3153
rect 4081 3124 4094 3148
rect 4118 3129 4303 3148
rect 4327 3129 4440 3153
rect 4118 3124 4440 3129
rect 4081 3120 4440 3124
rect 4507 3148 4656 3156
rect 4507 3128 4518 3148
rect 4538 3128 4656 3148
rect 4507 3121 4656 3128
rect 4507 3120 4548 3121
rect 3831 3067 3868 3068
rect 3927 3067 3964 3068
rect 3983 3067 4019 3119
rect 4038 3067 4075 3068
rect 3731 3058 3869 3067
rect 3731 3038 3840 3058
rect 3860 3038 3869 3058
rect 3731 3031 3869 3038
rect 3927 3058 4075 3067
rect 3927 3038 3936 3058
rect 3956 3038 4046 3058
rect 4066 3038 4075 3058
rect 3731 3029 3827 3031
rect 3927 3028 4075 3038
rect 4134 3058 4171 3068
rect 4246 3067 4283 3068
rect 4227 3065 4283 3067
rect 4134 3038 4142 3058
rect 4162 3038 4171 3058
rect 3983 3027 4019 3028
rect 1360 2985 1470 2999
rect 1360 2982 1403 2985
rect 1360 2977 1364 2982
rect 1036 2909 1204 2911
rect 760 2903 1204 2909
rect 113 2845 147 2877
rect 109 2836 147 2845
rect 109 2818 119 2836
rect 137 2818 147 2836
rect 109 2812 147 2818
rect 265 2814 299 2877
rect 421 2882 532 2888
rect 421 2874 462 2882
rect 421 2854 429 2874
rect 448 2854 462 2874
rect 421 2852 462 2854
rect 490 2874 532 2882
rect 490 2854 506 2874
rect 525 2854 532 2874
rect 490 2852 532 2854
rect 421 2837 532 2852
rect 759 2883 1204 2903
rect 759 2814 797 2883
rect 1036 2882 1204 2883
rect 1282 2955 1364 2977
rect 1393 2955 1403 2982
rect 1431 2958 1438 2985
rect 1467 2977 1470 2985
rect 3465 2994 3576 3009
rect 3465 2992 3507 2994
rect 1467 2958 1532 2977
rect 1431 2955 1532 2958
rect 1282 2953 1532 2955
rect 1282 2874 1319 2953
rect 1360 2940 1470 2953
rect 1434 2884 1465 2885
rect 1282 2854 1291 2874
rect 1311 2854 1319 2874
rect 1282 2844 1319 2854
rect 1378 2874 1465 2884
rect 1378 2854 1387 2874
rect 1407 2854 1465 2874
rect 1378 2845 1465 2854
rect 1378 2844 1415 2845
rect 109 2808 146 2812
rect 265 2803 797 2814
rect 264 2787 797 2803
rect 1434 2792 1465 2845
rect 1495 2874 1532 2953
rect 1703 2963 2096 2970
rect 1703 2946 1711 2963
rect 1743 2950 2096 2963
rect 2116 2950 2119 2970
rect 3198 2965 3239 2974
rect 1743 2946 2119 2950
rect 1703 2945 2119 2946
rect 2793 2963 2961 2964
rect 3198 2963 3207 2965
rect 1703 2944 2044 2945
rect 1647 2884 1678 2885
rect 1495 2854 1504 2874
rect 1524 2854 1532 2874
rect 1495 2844 1532 2854
rect 1591 2877 1678 2884
rect 1591 2874 1652 2877
rect 1591 2854 1600 2874
rect 1620 2857 1652 2874
rect 1673 2857 1678 2877
rect 1620 2854 1678 2857
rect 1591 2847 1678 2854
rect 1703 2874 1740 2944
rect 2006 2943 2043 2944
rect 2793 2943 3207 2963
rect 3233 2943 3239 2965
rect 3465 2972 3472 2992
rect 3491 2972 3507 2992
rect 3465 2964 3507 2972
rect 3535 2992 3576 2994
rect 3535 2972 3549 2992
rect 3568 2972 3576 2992
rect 3535 2964 3576 2972
rect 3831 2968 3868 2969
rect 4134 2968 4171 3038
rect 4196 3058 4283 3065
rect 4196 3055 4254 3058
rect 4196 3035 4201 3055
rect 4222 3038 4254 3055
rect 4274 3038 4283 3058
rect 4222 3035 4283 3038
rect 4196 3028 4283 3035
rect 4342 3058 4379 3068
rect 4342 3038 4350 3058
rect 4370 3038 4379 3058
rect 4196 3027 4227 3028
rect 3830 2967 4171 2968
rect 3465 2958 3576 2964
rect 3755 2962 4171 2967
rect 2793 2937 3239 2943
rect 2793 2935 2961 2937
rect 1855 2884 1891 2885
rect 1703 2854 1712 2874
rect 1732 2854 1740 2874
rect 1591 2845 1647 2847
rect 1591 2844 1628 2845
rect 1703 2844 1740 2854
rect 1799 2874 1947 2884
rect 2047 2881 2143 2883
rect 1799 2854 1808 2874
rect 1828 2869 1918 2874
rect 1828 2854 1863 2869
rect 1799 2845 1863 2854
rect 1799 2844 1836 2845
rect 1855 2828 1863 2845
rect 1884 2854 1918 2869
rect 1938 2854 1947 2874
rect 1884 2845 1947 2854
rect 2005 2874 2143 2881
rect 2005 2854 2014 2874
rect 2034 2854 2143 2874
rect 2005 2845 2143 2854
rect 1884 2828 1891 2845
rect 1910 2844 1947 2845
rect 2006 2844 2043 2845
rect 1855 2793 1891 2828
rect 1326 2791 1367 2792
rect 264 2786 778 2787
rect 1218 2784 1367 2791
rect 1218 2764 1336 2784
rect 1356 2764 1367 2784
rect 1218 2756 1367 2764
rect 1434 2788 1793 2792
rect 1434 2783 1756 2788
rect 1434 2759 1547 2783
rect 1571 2764 1756 2783
rect 1780 2764 1793 2788
rect 1571 2759 1793 2764
rect 1434 2756 1793 2759
rect 1855 2756 1890 2793
rect 1958 2790 2058 2793
rect 1958 2786 2025 2790
rect 1958 2760 1970 2786
rect 1996 2764 2025 2786
rect 2051 2764 2058 2790
rect 1996 2760 2058 2764
rect 1958 2756 2058 2760
rect 112 2745 149 2746
rect 110 2737 150 2745
rect 110 2719 121 2737
rect 139 2719 150 2737
rect 1434 2735 1465 2756
rect 1855 2735 1891 2756
rect 1277 2734 1314 2735
rect 110 2671 150 2719
rect 1276 2725 1314 2734
rect 1276 2705 1285 2725
rect 1305 2705 1314 2725
rect 1276 2697 1314 2705
rect 1380 2729 1465 2735
rect 1490 2734 1527 2735
rect 1380 2709 1388 2729
rect 1408 2709 1465 2729
rect 1380 2701 1465 2709
rect 1489 2725 1527 2734
rect 1489 2705 1498 2725
rect 1518 2705 1527 2725
rect 1380 2700 1416 2701
rect 1489 2697 1527 2705
rect 1593 2729 1678 2735
rect 1698 2734 1735 2735
rect 1593 2709 1601 2729
rect 1621 2728 1678 2729
rect 1621 2709 1650 2728
rect 1593 2708 1650 2709
rect 1671 2708 1678 2728
rect 1593 2701 1678 2708
rect 1697 2725 1735 2734
rect 1697 2705 1706 2725
rect 1726 2705 1735 2725
rect 1593 2700 1629 2701
rect 1697 2697 1735 2705
rect 1801 2729 1945 2735
rect 1801 2709 1809 2729
rect 1829 2709 1917 2729
rect 1937 2709 1945 2729
rect 1801 2701 1945 2709
rect 1801 2700 1837 2701
rect 1909 2700 1945 2701
rect 2011 2734 2048 2735
rect 2011 2733 2049 2734
rect 2011 2725 2075 2733
rect 2011 2705 2020 2725
rect 2040 2711 2075 2725
rect 2095 2711 2098 2731
rect 2040 2706 2098 2711
rect 2040 2705 2075 2706
rect 421 2675 531 2689
rect 421 2672 464 2675
rect 110 2664 235 2671
rect 421 2667 425 2672
rect 110 2645 202 2664
rect 227 2645 235 2664
rect 110 2635 235 2645
rect 343 2645 425 2667
rect 454 2645 464 2672
rect 492 2648 499 2675
rect 528 2667 531 2675
rect 1277 2668 1314 2697
rect 528 2648 593 2667
rect 1278 2666 1314 2668
rect 1490 2666 1527 2697
rect 1698 2670 1735 2697
rect 2011 2693 2075 2705
rect 492 2645 593 2648
rect 343 2643 593 2645
rect 110 2615 150 2635
rect 109 2606 150 2615
rect 109 2588 119 2606
rect 137 2588 150 2606
rect 109 2579 150 2588
rect 109 2578 146 2579
rect 343 2564 380 2643
rect 421 2630 531 2643
rect 495 2574 526 2575
rect 343 2544 352 2564
rect 372 2544 380 2564
rect 343 2534 380 2544
rect 439 2564 526 2574
rect 439 2544 448 2564
rect 468 2544 526 2564
rect 439 2535 526 2544
rect 439 2534 476 2535
rect 112 2512 149 2516
rect 109 2507 149 2512
rect 109 2489 121 2507
rect 139 2489 149 2507
rect 109 2309 149 2489
rect 495 2482 526 2535
rect 556 2564 593 2643
rect 764 2640 1157 2660
rect 1177 2640 1180 2660
rect 1278 2644 1527 2666
rect 1696 2665 1737 2670
rect 2115 2667 2142 2845
rect 2793 2757 2820 2935
rect 3198 2932 3239 2937
rect 3408 2936 3657 2958
rect 3755 2942 3758 2962
rect 3778 2942 4171 2962
rect 4342 2959 4379 3038
rect 4409 3067 4440 3120
rect 4786 3113 4826 3293
rect 4786 3095 4796 3113
rect 4814 3095 4826 3113
rect 4786 3090 4826 3095
rect 4786 3086 4823 3090
rect 4459 3067 4496 3068
rect 4409 3058 4496 3067
rect 4409 3038 4467 3058
rect 4487 3038 4496 3058
rect 4409 3028 4496 3038
rect 4555 3058 4592 3068
rect 4555 3038 4563 3058
rect 4583 3038 4592 3058
rect 4409 3027 4440 3028
rect 4404 2959 4514 2972
rect 4555 2959 4592 3038
rect 4789 3023 4826 3024
rect 4785 3014 4826 3023
rect 4785 2996 4798 3014
rect 4816 2996 4826 3014
rect 4785 2987 4826 2996
rect 4785 2967 4825 2987
rect 4342 2957 4592 2959
rect 4342 2954 4443 2957
rect 2860 2897 2924 2909
rect 3200 2905 3237 2932
rect 3408 2905 3445 2936
rect 3621 2934 3657 2936
rect 4342 2935 4407 2954
rect 3621 2905 3658 2934
rect 4404 2927 4407 2935
rect 4436 2927 4443 2954
rect 4471 2930 4481 2957
rect 4510 2935 4592 2957
rect 4700 2957 4825 2967
rect 4700 2938 4708 2957
rect 4733 2938 4825 2957
rect 4510 2930 4514 2935
rect 4700 2931 4825 2938
rect 4471 2927 4514 2930
rect 4404 2913 4514 2927
rect 2860 2896 2895 2897
rect 2837 2891 2895 2896
rect 2837 2871 2840 2891
rect 2860 2877 2895 2891
rect 2915 2877 2924 2897
rect 2860 2869 2924 2877
rect 2886 2868 2924 2869
rect 2887 2867 2924 2868
rect 2990 2901 3026 2902
rect 3098 2901 3134 2902
rect 2990 2893 3134 2901
rect 2990 2873 2998 2893
rect 3018 2890 3106 2893
rect 3018 2873 3050 2890
rect 3070 2873 3106 2890
rect 3126 2873 3134 2893
rect 2990 2867 3134 2873
rect 3200 2897 3238 2905
rect 3306 2901 3342 2902
rect 3200 2877 3209 2897
rect 3229 2877 3238 2897
rect 3200 2868 3238 2877
rect 3257 2894 3342 2901
rect 3257 2874 3264 2894
rect 3285 2893 3342 2894
rect 3285 2874 3314 2893
rect 3257 2873 3314 2874
rect 3334 2873 3342 2893
rect 3200 2867 3237 2868
rect 3257 2867 3342 2873
rect 3408 2897 3446 2905
rect 3519 2901 3555 2902
rect 3408 2877 3417 2897
rect 3437 2877 3446 2897
rect 3408 2868 3446 2877
rect 3470 2893 3555 2901
rect 3470 2873 3527 2893
rect 3547 2873 3555 2893
rect 3408 2867 3445 2868
rect 3470 2867 3555 2873
rect 3621 2897 3659 2905
rect 3621 2877 3630 2897
rect 3650 2877 3659 2897
rect 3621 2868 3659 2877
rect 4785 2883 4825 2931
rect 3621 2867 3658 2868
rect 3044 2846 3080 2867
rect 3470 2846 3501 2867
rect 4785 2865 4796 2883
rect 4814 2865 4825 2883
rect 4785 2857 4825 2865
rect 4786 2856 4823 2857
rect 2877 2842 2977 2846
rect 2877 2838 2939 2842
rect 2877 2812 2884 2838
rect 2910 2816 2939 2838
rect 2965 2816 2977 2842
rect 2910 2812 2977 2816
rect 2877 2809 2977 2812
rect 3045 2809 3080 2846
rect 3142 2843 3501 2846
rect 3142 2838 3364 2843
rect 3142 2814 3155 2838
rect 3179 2819 3364 2838
rect 3388 2819 3501 2843
rect 3179 2814 3501 2819
rect 3142 2810 3501 2814
rect 3568 2838 3717 2846
rect 3568 2818 3579 2838
rect 3599 2818 3717 2838
rect 3568 2811 3717 2818
rect 4157 2815 4671 2816
rect 3568 2810 3609 2811
rect 2892 2757 2929 2758
rect 2988 2757 3025 2758
rect 3044 2757 3080 2809
rect 3099 2757 3136 2758
rect 2792 2748 2930 2757
rect 2792 2728 2901 2748
rect 2921 2728 2930 2748
rect 2792 2721 2930 2728
rect 2988 2748 3136 2757
rect 2988 2728 2997 2748
rect 3017 2728 3107 2748
rect 3127 2728 3136 2748
rect 2792 2719 2888 2721
rect 2988 2718 3136 2728
rect 3195 2748 3232 2758
rect 3307 2757 3344 2758
rect 3288 2755 3344 2757
rect 3195 2728 3203 2748
rect 3223 2728 3232 2748
rect 3044 2717 3080 2718
rect 1974 2665 2142 2667
rect 1696 2659 2142 2665
rect 764 2635 1180 2640
rect 1359 2638 1470 2644
rect 764 2634 1105 2635
rect 708 2574 739 2575
rect 556 2544 565 2564
rect 585 2544 593 2564
rect 556 2534 593 2544
rect 652 2567 739 2574
rect 652 2564 713 2567
rect 652 2544 661 2564
rect 681 2547 713 2564
rect 734 2547 739 2567
rect 681 2544 739 2547
rect 652 2537 739 2544
rect 764 2564 801 2634
rect 1067 2633 1104 2634
rect 1359 2630 1400 2638
rect 1359 2610 1367 2630
rect 1386 2610 1400 2630
rect 1359 2608 1400 2610
rect 1428 2630 1470 2638
rect 1428 2610 1444 2630
rect 1463 2610 1470 2630
rect 1696 2637 1702 2659
rect 1728 2639 2142 2659
rect 2892 2658 2929 2659
rect 3195 2658 3232 2728
rect 3257 2748 3344 2755
rect 3257 2745 3315 2748
rect 3257 2725 3262 2745
rect 3283 2728 3315 2745
rect 3335 2728 3344 2748
rect 3283 2725 3344 2728
rect 3257 2718 3344 2725
rect 3403 2748 3440 2758
rect 3403 2728 3411 2748
rect 3431 2728 3440 2748
rect 3257 2717 3288 2718
rect 2891 2657 3232 2658
rect 1728 2637 1737 2639
rect 1974 2638 2142 2639
rect 2816 2652 3232 2657
rect 1696 2628 1737 2637
rect 2816 2632 2819 2652
rect 2839 2632 3232 2652
rect 3403 2649 3440 2728
rect 3470 2757 3501 2810
rect 4138 2799 4671 2815
rect 4138 2788 4670 2799
rect 4789 2790 4826 2794
rect 3520 2757 3557 2758
rect 3470 2748 3557 2757
rect 3470 2728 3528 2748
rect 3548 2728 3557 2748
rect 3470 2718 3557 2728
rect 3616 2748 3653 2758
rect 3616 2728 3624 2748
rect 3644 2728 3653 2748
rect 3470 2717 3501 2718
rect 3465 2649 3575 2662
rect 3616 2649 3653 2728
rect 3403 2647 3653 2649
rect 3403 2644 3504 2647
rect 3403 2625 3468 2644
rect 1428 2608 1470 2610
rect 1359 2593 1470 2608
rect 3465 2617 3468 2625
rect 3497 2617 3504 2644
rect 3532 2620 3542 2647
rect 3571 2625 3653 2647
rect 3731 2719 3899 2720
rect 4138 2719 4176 2788
rect 3731 2699 4176 2719
rect 4403 2750 4514 2765
rect 4403 2748 4445 2750
rect 4403 2728 4410 2748
rect 4429 2728 4445 2748
rect 4403 2720 4445 2728
rect 4473 2748 4514 2750
rect 4473 2728 4487 2748
rect 4506 2728 4514 2748
rect 4473 2720 4514 2728
rect 4403 2714 4514 2720
rect 4636 2725 4670 2788
rect 4788 2784 4826 2790
rect 4788 2766 4798 2784
rect 4816 2766 4826 2784
rect 4788 2757 4826 2766
rect 4788 2725 4822 2757
rect 3731 2693 4175 2699
rect 3731 2691 3899 2693
rect 3571 2620 3575 2625
rect 3532 2617 3575 2620
rect 3465 2603 3575 2617
rect 2694 2589 2762 2598
rect 916 2574 952 2575
rect 764 2544 773 2564
rect 793 2544 801 2564
rect 652 2535 708 2537
rect 652 2534 689 2535
rect 764 2534 801 2544
rect 860 2564 1008 2574
rect 1108 2571 1204 2573
rect 860 2544 869 2564
rect 889 2544 979 2564
rect 999 2544 1008 2564
rect 860 2535 1008 2544
rect 1066 2564 1204 2571
rect 1066 2544 1075 2564
rect 1095 2544 1204 2564
rect 2694 2560 2709 2589
rect 2757 2569 2762 2589
rect 2757 2560 2764 2569
rect 2694 2549 2764 2560
rect 1066 2535 1204 2544
rect 860 2534 897 2535
rect 916 2483 952 2535
rect 971 2534 1008 2535
rect 1067 2534 1104 2535
rect 387 2481 428 2482
rect 279 2474 428 2481
rect 279 2454 397 2474
rect 417 2454 428 2474
rect 279 2446 428 2454
rect 495 2478 854 2482
rect 495 2473 817 2478
rect 495 2449 608 2473
rect 632 2454 817 2473
rect 841 2454 854 2478
rect 632 2449 854 2454
rect 495 2446 854 2449
rect 916 2446 951 2483
rect 1019 2480 1119 2483
rect 1019 2476 1086 2480
rect 1019 2450 1031 2476
rect 1057 2454 1086 2476
rect 1112 2454 1119 2480
rect 1057 2450 1119 2454
rect 1019 2446 1119 2450
rect 495 2425 526 2446
rect 916 2425 952 2446
rect 338 2424 375 2425
rect 337 2415 375 2424
rect 337 2395 346 2415
rect 366 2395 375 2415
rect 337 2387 375 2395
rect 441 2419 526 2425
rect 551 2424 588 2425
rect 441 2399 449 2419
rect 469 2399 526 2419
rect 441 2391 526 2399
rect 550 2415 588 2424
rect 550 2395 559 2415
rect 579 2395 588 2415
rect 441 2390 477 2391
rect 550 2387 588 2395
rect 654 2419 739 2425
rect 759 2424 796 2425
rect 654 2399 662 2419
rect 682 2418 739 2419
rect 682 2399 711 2418
rect 654 2398 711 2399
rect 732 2398 739 2418
rect 654 2391 739 2398
rect 758 2415 796 2424
rect 758 2395 767 2415
rect 787 2395 796 2415
rect 654 2390 690 2391
rect 758 2387 796 2395
rect 862 2419 1006 2425
rect 862 2399 870 2419
rect 890 2416 978 2419
rect 890 2399 921 2416
rect 862 2396 921 2399
rect 944 2399 978 2416
rect 998 2399 1006 2419
rect 944 2396 1006 2399
rect 862 2391 1006 2396
rect 862 2390 898 2391
rect 970 2390 1006 2391
rect 1072 2424 1109 2425
rect 1072 2423 1110 2424
rect 1072 2415 1136 2423
rect 1072 2395 1081 2415
rect 1101 2401 1136 2415
rect 1156 2401 1159 2421
rect 1101 2396 1159 2401
rect 1101 2395 1136 2396
rect 338 2358 375 2387
rect 339 2356 375 2358
rect 551 2356 588 2387
rect 339 2334 588 2356
rect 759 2355 796 2387
rect 1072 2383 1136 2395
rect 1176 2357 1203 2535
rect 2703 2442 2764 2549
rect 3731 2513 3758 2691
rect 3798 2653 3862 2665
rect 4138 2661 4175 2693
rect 4346 2692 4595 2714
rect 4636 2693 4822 2725
rect 4650 2692 4822 2693
rect 4346 2661 4383 2692
rect 4559 2690 4595 2692
rect 4559 2661 4596 2690
rect 4788 2664 4822 2692
rect 3798 2652 3833 2653
rect 3775 2647 3833 2652
rect 3775 2627 3778 2647
rect 3798 2633 3833 2647
rect 3853 2633 3862 2653
rect 3798 2625 3862 2633
rect 3824 2624 3862 2625
rect 3825 2623 3862 2624
rect 3928 2657 3964 2658
rect 4036 2657 4072 2658
rect 3928 2650 4072 2657
rect 3928 2649 3988 2650
rect 3928 2629 3936 2649
rect 3956 2630 3988 2649
rect 4013 2649 4072 2650
rect 4013 2630 4044 2649
rect 3956 2629 4044 2630
rect 4064 2629 4072 2649
rect 3928 2623 4072 2629
rect 4138 2653 4176 2661
rect 4244 2657 4280 2658
rect 4138 2633 4147 2653
rect 4167 2633 4176 2653
rect 4138 2624 4176 2633
rect 4195 2650 4280 2657
rect 4195 2630 4202 2650
rect 4223 2649 4280 2650
rect 4223 2630 4252 2649
rect 4195 2629 4252 2630
rect 4272 2629 4280 2649
rect 4138 2623 4175 2624
rect 4195 2623 4280 2629
rect 4346 2653 4384 2661
rect 4457 2657 4493 2658
rect 4346 2633 4355 2653
rect 4375 2633 4384 2653
rect 4346 2624 4384 2633
rect 4408 2649 4493 2657
rect 4408 2629 4465 2649
rect 4485 2629 4493 2649
rect 4346 2623 4383 2624
rect 4408 2623 4493 2629
rect 4559 2653 4597 2661
rect 4559 2633 4568 2653
rect 4588 2633 4597 2653
rect 4559 2624 4597 2633
rect 4786 2654 4823 2664
rect 4786 2636 4796 2654
rect 4814 2636 4823 2654
rect 4786 2627 4823 2636
rect 4788 2626 4822 2627
rect 4559 2623 4596 2624
rect 3982 2602 4018 2623
rect 4408 2602 4439 2623
rect 3815 2598 3915 2602
rect 3815 2594 3877 2598
rect 3815 2568 3822 2594
rect 3848 2572 3877 2594
rect 3903 2572 3915 2598
rect 3848 2568 3915 2572
rect 3815 2565 3915 2568
rect 3983 2565 4018 2602
rect 4080 2599 4439 2602
rect 4080 2594 4302 2599
rect 4080 2570 4093 2594
rect 4117 2575 4302 2594
rect 4326 2575 4439 2599
rect 4117 2570 4439 2575
rect 4080 2566 4439 2570
rect 4506 2594 4655 2602
rect 4506 2574 4517 2594
rect 4537 2574 4655 2594
rect 4506 2567 4655 2574
rect 4506 2566 4547 2567
rect 3830 2513 3867 2514
rect 3926 2513 3963 2514
rect 3982 2513 4018 2565
rect 4037 2513 4074 2514
rect 3730 2504 3868 2513
rect 2694 2441 2764 2442
rect 3355 2470 3466 2485
rect 3730 2484 3839 2504
rect 3859 2484 3868 2504
rect 3730 2477 3868 2484
rect 3926 2504 4074 2513
rect 3926 2484 3935 2504
rect 3955 2484 4045 2504
rect 4065 2484 4074 2504
rect 3730 2475 3826 2477
rect 3926 2474 4074 2484
rect 4133 2504 4170 2514
rect 4245 2513 4282 2514
rect 4226 2511 4282 2513
rect 4133 2484 4141 2504
rect 4161 2484 4170 2504
rect 3982 2473 4018 2474
rect 3355 2468 3397 2470
rect 3355 2448 3362 2468
rect 3381 2448 3397 2468
rect 2694 2440 2802 2441
rect 3355 2440 3397 2448
rect 3425 2468 3466 2470
rect 3425 2448 3439 2468
rect 3458 2448 3466 2468
rect 3425 2440 3466 2448
rect 2683 2439 2851 2440
rect 1470 2406 1580 2420
rect 1470 2403 1513 2406
rect 1470 2398 1474 2403
rect 1035 2355 1203 2357
rect 759 2352 1203 2355
rect 420 2328 531 2334
rect 420 2320 461 2328
rect 109 2265 148 2309
rect 420 2300 428 2320
rect 447 2300 461 2320
rect 420 2298 461 2300
rect 489 2320 531 2328
rect 489 2300 505 2320
rect 524 2300 531 2320
rect 489 2298 531 2300
rect 420 2284 531 2298
rect 757 2329 1203 2352
rect 109 2241 149 2265
rect 449 2241 496 2243
rect 757 2241 795 2329
rect 1035 2328 1203 2329
rect 1392 2376 1474 2398
rect 1503 2376 1513 2403
rect 1541 2379 1548 2406
rect 1577 2398 1580 2406
rect 2683 2413 3127 2439
rect 3355 2434 3466 2440
rect 2683 2411 2851 2413
rect 2683 2409 2802 2411
rect 1577 2379 1642 2398
rect 1541 2376 1642 2379
rect 1392 2374 1642 2376
rect 1392 2295 1429 2374
rect 1470 2361 1580 2374
rect 1544 2305 1575 2306
rect 1392 2275 1401 2295
rect 1421 2275 1429 2295
rect 1392 2265 1429 2275
rect 1488 2295 1575 2305
rect 1488 2275 1497 2295
rect 1517 2275 1575 2295
rect 1488 2266 1575 2275
rect 1488 2265 1525 2266
rect 109 2208 795 2241
rect 1544 2213 1575 2266
rect 1605 2295 1642 2374
rect 1813 2393 1845 2405
rect 1813 2373 1815 2393
rect 1836 2391 1845 2393
rect 1836 2389 2188 2391
rect 1836 2373 2206 2389
rect 1813 2371 2206 2373
rect 2226 2371 2229 2389
rect 1813 2366 2229 2371
rect 1813 2365 2154 2366
rect 1757 2305 1788 2306
rect 1605 2275 1614 2295
rect 1634 2275 1642 2295
rect 1605 2265 1642 2275
rect 1701 2298 1788 2305
rect 1701 2295 1762 2298
rect 1701 2275 1710 2295
rect 1730 2278 1762 2295
rect 1783 2278 1788 2298
rect 1730 2275 1788 2278
rect 1701 2268 1788 2275
rect 1813 2295 1850 2365
rect 2116 2364 2153 2365
rect 1965 2305 2001 2306
rect 1813 2275 1822 2295
rect 1842 2275 1850 2295
rect 1701 2266 1757 2268
rect 1701 2265 1738 2266
rect 1813 2265 1850 2275
rect 1909 2295 2057 2305
rect 2157 2302 2253 2304
rect 1909 2275 1918 2295
rect 1938 2286 2028 2295
rect 1938 2275 1969 2286
rect 1909 2266 1969 2275
rect 1909 2265 1946 2266
rect 1965 2254 1969 2266
rect 1996 2275 2028 2286
rect 2048 2275 2057 2295
rect 1996 2266 2057 2275
rect 2115 2295 2253 2302
rect 2115 2275 2124 2295
rect 2144 2275 2253 2295
rect 2115 2266 2253 2275
rect 1996 2254 2001 2266
rect 2020 2265 2057 2266
rect 2116 2265 2153 2266
rect 1965 2214 2001 2254
rect 1436 2212 1477 2213
rect 108 2151 147 2208
rect 757 2206 795 2208
rect 1328 2205 1477 2212
rect 1328 2185 1446 2205
rect 1466 2185 1477 2205
rect 1328 2177 1477 2185
rect 1544 2209 1903 2213
rect 1544 2204 1866 2209
rect 1544 2180 1657 2204
rect 1681 2185 1866 2204
rect 1890 2185 1903 2209
rect 1681 2180 1903 2185
rect 1544 2177 1903 2180
rect 1965 2177 2000 2214
rect 2068 2211 2168 2214
rect 2068 2207 2135 2211
rect 2068 2181 2080 2207
rect 2106 2185 2135 2207
rect 2161 2185 2168 2211
rect 2106 2181 2168 2185
rect 2068 2177 2168 2181
rect 1544 2156 1575 2177
rect 1965 2156 2001 2177
rect 1387 2155 1424 2156
rect 108 2149 156 2151
rect 108 2131 119 2149
rect 137 2131 156 2149
rect 1386 2146 1424 2155
rect 108 2122 156 2131
rect 109 2121 156 2122
rect 422 2126 532 2140
rect 422 2123 465 2126
rect 422 2118 426 2123
rect 344 2096 426 2118
rect 455 2096 465 2123
rect 493 2099 500 2126
rect 529 2118 532 2126
rect 1386 2126 1395 2146
rect 1415 2126 1424 2146
rect 1386 2118 1424 2126
rect 1490 2150 1575 2156
rect 1600 2155 1637 2156
rect 1490 2130 1498 2150
rect 1518 2130 1575 2150
rect 1490 2122 1575 2130
rect 1599 2146 1637 2155
rect 1599 2126 1608 2146
rect 1628 2126 1637 2146
rect 1490 2121 1526 2122
rect 1599 2118 1637 2126
rect 1703 2150 1788 2156
rect 1808 2155 1845 2156
rect 1703 2130 1711 2150
rect 1731 2149 1788 2150
rect 1731 2130 1760 2149
rect 1703 2129 1760 2130
rect 1781 2129 1788 2149
rect 1703 2122 1788 2129
rect 1807 2146 1845 2155
rect 1807 2126 1816 2146
rect 1836 2126 1845 2146
rect 1703 2121 1739 2122
rect 1807 2118 1845 2126
rect 1911 2150 2055 2156
rect 1911 2130 1919 2150
rect 1939 2130 2027 2150
rect 2047 2130 2055 2150
rect 1911 2122 2055 2130
rect 1911 2121 1947 2122
rect 2019 2121 2055 2122
rect 2121 2155 2158 2156
rect 2121 2154 2159 2155
rect 2121 2146 2185 2154
rect 2121 2126 2130 2146
rect 2150 2132 2185 2146
rect 2205 2132 2208 2152
rect 2150 2127 2208 2132
rect 2150 2126 2185 2127
rect 529 2099 594 2118
rect 493 2096 594 2099
rect 344 2094 594 2096
rect 112 2058 149 2059
rect 108 2055 149 2058
rect 108 2050 150 2055
rect 108 2032 121 2050
rect 139 2032 150 2050
rect 108 2018 150 2032
rect 188 2018 235 2022
rect 108 2012 235 2018
rect 108 1983 196 2012
rect 225 1983 235 2012
rect 344 2015 381 2094
rect 422 2081 532 2094
rect 496 2025 527 2026
rect 344 1995 353 2015
rect 373 1995 381 2015
rect 344 1985 381 1995
rect 440 2015 527 2025
rect 440 1995 449 2015
rect 469 1995 527 2015
rect 440 1986 527 1995
rect 440 1985 477 1986
rect 108 1979 235 1983
rect 108 1962 147 1979
rect 188 1978 235 1979
rect 108 1944 119 1962
rect 137 1944 147 1962
rect 108 1935 147 1944
rect 109 1934 146 1935
rect 496 1933 527 1986
rect 557 2015 594 2094
rect 765 2091 1158 2111
rect 1178 2091 1181 2111
rect 765 2086 1181 2091
rect 1387 2089 1424 2118
rect 1388 2087 1424 2089
rect 1600 2087 1637 2118
rect 765 2085 1106 2086
rect 709 2025 740 2026
rect 557 1995 566 2015
rect 586 1995 594 2015
rect 557 1985 594 1995
rect 653 2018 740 2025
rect 653 2015 714 2018
rect 653 1995 662 2015
rect 682 1998 714 2015
rect 735 1998 740 2018
rect 682 1995 740 1998
rect 653 1988 740 1995
rect 765 2015 802 2085
rect 1068 2084 1105 2085
rect 1388 2065 1637 2087
rect 1808 2086 1845 2118
rect 2121 2114 2185 2126
rect 2225 2096 2252 2266
rect 2683 2233 2710 2409
rect 2750 2373 2814 2385
rect 3090 2381 3127 2413
rect 3298 2412 3547 2434
rect 3830 2414 3867 2415
rect 4133 2414 4170 2484
rect 4195 2504 4282 2511
rect 4195 2501 4253 2504
rect 4195 2481 4200 2501
rect 4221 2484 4253 2501
rect 4273 2484 4282 2504
rect 4221 2481 4282 2484
rect 4195 2474 4282 2481
rect 4341 2504 4378 2514
rect 4341 2484 4349 2504
rect 4369 2484 4378 2504
rect 4195 2473 4226 2474
rect 3829 2413 4170 2414
rect 3298 2381 3335 2412
rect 3511 2410 3547 2412
rect 3511 2381 3548 2410
rect 3754 2408 4170 2413
rect 3754 2388 3757 2408
rect 3777 2388 4170 2408
rect 4341 2405 4378 2484
rect 4408 2513 4439 2566
rect 4789 2564 4826 2565
rect 4788 2555 4827 2564
rect 4788 2537 4798 2555
rect 4816 2537 4827 2555
rect 4700 2520 4747 2521
rect 4788 2520 4827 2537
rect 4700 2516 4827 2520
rect 4458 2513 4495 2514
rect 4408 2504 4495 2513
rect 4408 2484 4466 2504
rect 4486 2484 4495 2504
rect 4408 2474 4495 2484
rect 4554 2504 4591 2514
rect 4554 2484 4562 2504
rect 4582 2484 4591 2504
rect 4408 2473 4439 2474
rect 4403 2405 4513 2418
rect 4554 2405 4591 2484
rect 4700 2487 4710 2516
rect 4739 2487 4827 2516
rect 4700 2481 4827 2487
rect 4700 2477 4747 2481
rect 4785 2467 4827 2481
rect 4785 2449 4796 2467
rect 4814 2449 4827 2467
rect 4785 2444 4827 2449
rect 4786 2441 4827 2444
rect 4786 2440 4823 2441
rect 4341 2403 4591 2405
rect 4341 2400 4442 2403
rect 4341 2381 4406 2400
rect 2750 2372 2785 2373
rect 2727 2367 2785 2372
rect 2727 2347 2730 2367
rect 2750 2353 2785 2367
rect 2805 2353 2814 2373
rect 2750 2345 2814 2353
rect 2776 2344 2814 2345
rect 2777 2343 2814 2344
rect 2880 2377 2916 2378
rect 2988 2377 3024 2378
rect 2880 2370 3024 2377
rect 2880 2369 2938 2370
rect 2880 2349 2888 2369
rect 2908 2351 2938 2369
rect 2967 2369 3024 2370
rect 2967 2351 2996 2369
rect 2908 2349 2996 2351
rect 3016 2349 3024 2369
rect 2880 2343 3024 2349
rect 3090 2373 3128 2381
rect 3196 2377 3232 2378
rect 3090 2353 3099 2373
rect 3119 2353 3128 2373
rect 3090 2344 3128 2353
rect 3147 2370 3232 2377
rect 3147 2350 3154 2370
rect 3175 2369 3232 2370
rect 3175 2350 3204 2369
rect 3147 2349 3204 2350
rect 3224 2349 3232 2369
rect 3090 2343 3127 2344
rect 3147 2343 3232 2349
rect 3298 2373 3336 2381
rect 3409 2377 3445 2378
rect 3298 2353 3307 2373
rect 3327 2353 3336 2373
rect 3298 2344 3336 2353
rect 3360 2369 3445 2377
rect 3360 2349 3417 2369
rect 3437 2349 3445 2369
rect 3298 2343 3335 2344
rect 3360 2343 3445 2349
rect 3511 2373 3549 2381
rect 3511 2353 3520 2373
rect 3540 2353 3549 2373
rect 4403 2373 4406 2381
rect 4435 2373 4442 2400
rect 4470 2376 4480 2403
rect 4509 2381 4591 2403
rect 4509 2376 4513 2381
rect 4470 2373 4513 2376
rect 4403 2359 4513 2373
rect 4779 2377 4826 2378
rect 4779 2368 4827 2377
rect 3511 2344 3549 2353
rect 4779 2350 4798 2368
rect 4816 2350 4827 2368
rect 4779 2348 4827 2350
rect 3511 2343 3548 2344
rect 2934 2322 2970 2343
rect 3360 2322 3391 2343
rect 2767 2318 2867 2322
rect 2767 2314 2829 2318
rect 2767 2288 2774 2314
rect 2800 2292 2829 2314
rect 2855 2292 2867 2318
rect 2800 2288 2867 2292
rect 2767 2285 2867 2288
rect 2935 2285 2970 2322
rect 3032 2319 3391 2322
rect 3032 2314 3254 2319
rect 3032 2290 3045 2314
rect 3069 2295 3254 2314
rect 3278 2295 3391 2319
rect 3069 2290 3391 2295
rect 3032 2286 3391 2290
rect 3458 2314 3607 2322
rect 3458 2294 3469 2314
rect 3489 2294 3607 2314
rect 3458 2287 3607 2294
rect 4140 2291 4178 2293
rect 4788 2291 4827 2348
rect 3458 2286 3499 2287
rect 2782 2233 2819 2234
rect 2878 2233 2915 2234
rect 2934 2233 2970 2285
rect 2989 2233 3026 2234
rect 2682 2224 2820 2233
rect 2682 2204 2791 2224
rect 2811 2204 2820 2224
rect 2682 2197 2820 2204
rect 2878 2224 3026 2233
rect 2878 2204 2887 2224
rect 2907 2204 2997 2224
rect 3017 2204 3026 2224
rect 2682 2195 2778 2197
rect 2878 2194 3026 2204
rect 3085 2224 3122 2234
rect 3197 2233 3234 2234
rect 3178 2231 3234 2233
rect 3085 2204 3093 2224
rect 3113 2204 3122 2224
rect 2934 2193 2970 2194
rect 2782 2134 2819 2135
rect 3085 2134 3122 2204
rect 3147 2224 3234 2231
rect 3147 2221 3205 2224
rect 3147 2201 3152 2221
rect 3173 2204 3205 2221
rect 3225 2204 3234 2224
rect 3173 2201 3234 2204
rect 3147 2194 3234 2201
rect 3293 2224 3330 2234
rect 3293 2204 3301 2224
rect 3321 2204 3330 2224
rect 3147 2193 3178 2194
rect 2781 2133 3122 2134
rect 2706 2128 3122 2133
rect 2706 2108 2709 2128
rect 2729 2108 3122 2128
rect 3293 2125 3330 2204
rect 3360 2233 3391 2286
rect 4140 2258 4826 2291
rect 3410 2233 3447 2234
rect 3360 2224 3447 2233
rect 3360 2204 3418 2224
rect 3438 2204 3447 2224
rect 3360 2194 3447 2204
rect 3506 2224 3543 2234
rect 3506 2204 3514 2224
rect 3534 2204 3543 2224
rect 3360 2193 3391 2194
rect 3355 2125 3465 2138
rect 3506 2125 3543 2204
rect 3293 2123 3543 2125
rect 3293 2120 3394 2123
rect 3293 2101 3358 2120
rect 2173 2088 2252 2096
rect 2084 2086 2252 2088
rect 1808 2079 2252 2086
rect 3355 2093 3358 2101
rect 3387 2093 3394 2120
rect 3422 2096 3432 2123
rect 3461 2101 3543 2123
rect 3732 2170 3900 2171
rect 4140 2170 4178 2258
rect 4439 2256 4486 2258
rect 4786 2234 4826 2258
rect 3732 2147 4178 2170
rect 4404 2201 4515 2215
rect 4404 2199 4446 2201
rect 4404 2179 4411 2199
rect 4430 2179 4446 2199
rect 4404 2171 4446 2179
rect 4474 2199 4515 2201
rect 4474 2179 4488 2199
rect 4507 2179 4515 2199
rect 4787 2190 4826 2234
rect 4474 2171 4515 2179
rect 4404 2165 4515 2171
rect 3732 2144 4176 2147
rect 3732 2142 3900 2144
rect 3461 2096 3465 2101
rect 3422 2093 3465 2096
rect 3355 2079 3465 2093
rect 1469 2059 1580 2065
rect 1808 2060 2178 2079
rect 2084 2059 2178 2060
rect 1469 2051 1510 2059
rect 1469 2031 1477 2051
rect 1496 2031 1510 2051
rect 1469 2029 1510 2031
rect 1538 2051 1580 2059
rect 1538 2031 1554 2051
rect 1573 2031 1580 2051
rect 2173 2050 2178 2059
rect 2226 2059 2252 2079
rect 2226 2050 2243 2059
rect 2173 2041 2243 2050
rect 1538 2029 1580 2031
rect 917 2025 953 2026
rect 765 1995 774 2015
rect 794 1995 802 2015
rect 653 1986 709 1988
rect 653 1985 690 1986
rect 765 1985 802 1995
rect 861 2015 1009 2025
rect 1109 2022 1205 2024
rect 861 1995 870 2015
rect 890 1995 980 2015
rect 1000 1995 1009 2015
rect 861 1986 1009 1995
rect 1067 2015 1205 2022
rect 1067 1995 1076 2015
rect 1096 1995 1205 2015
rect 1469 2014 1580 2029
rect 1067 1986 1205 1995
rect 861 1985 898 1986
rect 917 1934 953 1986
rect 972 1985 1009 1986
rect 1068 1985 1105 1986
rect 388 1932 429 1933
rect 280 1925 429 1932
rect 280 1905 398 1925
rect 418 1905 429 1925
rect 280 1897 429 1905
rect 496 1929 855 1933
rect 496 1924 818 1929
rect 496 1900 609 1924
rect 633 1905 818 1924
rect 842 1905 855 1929
rect 633 1900 855 1905
rect 496 1897 855 1900
rect 917 1897 952 1934
rect 1020 1931 1120 1934
rect 1020 1927 1087 1931
rect 1020 1901 1032 1927
rect 1058 1905 1087 1927
rect 1113 1905 1120 1931
rect 1058 1901 1120 1905
rect 1020 1897 1120 1901
rect 496 1876 527 1897
rect 917 1876 953 1897
rect 339 1875 376 1876
rect 113 1872 147 1873
rect 112 1863 149 1872
rect 112 1845 121 1863
rect 139 1845 149 1863
rect 112 1835 149 1845
rect 338 1866 376 1875
rect 338 1846 347 1866
rect 367 1846 376 1866
rect 338 1838 376 1846
rect 442 1870 527 1876
rect 552 1875 589 1876
rect 442 1850 450 1870
rect 470 1850 527 1870
rect 442 1842 527 1850
rect 551 1866 589 1875
rect 551 1846 560 1866
rect 580 1846 589 1866
rect 442 1841 478 1842
rect 551 1838 589 1846
rect 655 1870 740 1876
rect 760 1875 797 1876
rect 655 1850 663 1870
rect 683 1869 740 1870
rect 683 1850 712 1869
rect 655 1849 712 1850
rect 733 1849 740 1869
rect 655 1842 740 1849
rect 759 1866 797 1875
rect 759 1846 768 1866
rect 788 1846 797 1866
rect 655 1841 691 1842
rect 759 1838 797 1846
rect 863 1870 1007 1876
rect 863 1850 871 1870
rect 891 1869 979 1870
rect 891 1850 922 1869
rect 863 1849 922 1850
rect 947 1850 979 1869
rect 999 1850 1007 1870
rect 947 1849 1007 1850
rect 863 1842 1007 1849
rect 863 1841 899 1842
rect 971 1841 1007 1842
rect 1073 1875 1110 1876
rect 1073 1874 1111 1875
rect 1073 1866 1137 1874
rect 1073 1846 1082 1866
rect 1102 1852 1137 1866
rect 1157 1852 1160 1872
rect 1102 1847 1160 1852
rect 1102 1846 1137 1847
rect 113 1807 147 1835
rect 339 1809 376 1838
rect 340 1807 376 1809
rect 552 1807 589 1838
rect 113 1806 285 1807
rect 113 1774 299 1806
rect 340 1785 589 1807
rect 760 1806 797 1838
rect 1073 1834 1137 1846
rect 1177 1808 1204 1986
rect 3732 1964 3759 2142
rect 3799 2104 3863 2116
rect 4139 2112 4176 2144
rect 4347 2143 4596 2165
rect 4347 2112 4384 2143
rect 4560 2141 4596 2143
rect 4560 2112 4597 2141
rect 3799 2103 3834 2104
rect 3776 2098 3834 2103
rect 3776 2078 3779 2098
rect 3799 2084 3834 2098
rect 3854 2084 3863 2104
rect 3799 2076 3863 2084
rect 3825 2075 3863 2076
rect 3826 2074 3863 2075
rect 3929 2108 3965 2109
rect 4037 2108 4073 2109
rect 3929 2103 4073 2108
rect 3929 2100 3991 2103
rect 3929 2080 3937 2100
rect 3957 2083 3991 2100
rect 4014 2100 4073 2103
rect 4014 2083 4045 2100
rect 3957 2080 4045 2083
rect 4065 2080 4073 2100
rect 3929 2074 4073 2080
rect 4139 2104 4177 2112
rect 4245 2108 4281 2109
rect 4139 2084 4148 2104
rect 4168 2084 4177 2104
rect 4139 2075 4177 2084
rect 4196 2101 4281 2108
rect 4196 2081 4203 2101
rect 4224 2100 4281 2101
rect 4224 2081 4253 2100
rect 4196 2080 4253 2081
rect 4273 2080 4281 2100
rect 4139 2074 4176 2075
rect 4196 2074 4281 2080
rect 4347 2104 4385 2112
rect 4458 2108 4494 2109
rect 4347 2084 4356 2104
rect 4376 2084 4385 2104
rect 4347 2075 4385 2084
rect 4409 2100 4494 2108
rect 4409 2080 4466 2100
rect 4486 2080 4494 2100
rect 4347 2074 4384 2075
rect 4409 2074 4494 2080
rect 4560 2104 4598 2112
rect 4560 2084 4569 2104
rect 4589 2084 4598 2104
rect 4560 2075 4598 2084
rect 4560 2074 4597 2075
rect 3983 2053 4019 2074
rect 4409 2053 4440 2074
rect 3816 2049 3916 2053
rect 3816 2045 3878 2049
rect 3816 2019 3823 2045
rect 3849 2023 3878 2045
rect 3904 2023 3916 2049
rect 3849 2019 3916 2023
rect 3816 2016 3916 2019
rect 3984 2016 4019 2053
rect 4081 2050 4440 2053
rect 4081 2045 4303 2050
rect 4081 2021 4094 2045
rect 4118 2026 4303 2045
rect 4327 2026 4440 2050
rect 4118 2021 4440 2026
rect 4081 2017 4440 2021
rect 4507 2045 4656 2053
rect 4507 2025 4518 2045
rect 4538 2025 4656 2045
rect 4507 2018 4656 2025
rect 4507 2017 4548 2018
rect 3831 1964 3868 1965
rect 3927 1964 3964 1965
rect 3983 1964 4019 2016
rect 4038 1964 4075 1965
rect 3731 1955 3869 1964
rect 3731 1935 3840 1955
rect 3860 1935 3869 1955
rect 3731 1928 3869 1935
rect 3927 1955 4075 1964
rect 3927 1935 3936 1955
rect 3956 1935 4046 1955
rect 4066 1935 4075 1955
rect 3731 1926 3827 1928
rect 3927 1925 4075 1935
rect 4134 1955 4171 1965
rect 4246 1964 4283 1965
rect 4227 1962 4283 1964
rect 4134 1935 4142 1955
rect 4162 1935 4171 1955
rect 3983 1924 4019 1925
rect 1360 1882 1470 1896
rect 1360 1879 1403 1882
rect 1360 1874 1364 1879
rect 1036 1806 1204 1808
rect 760 1800 1204 1806
rect 113 1742 147 1774
rect 109 1733 147 1742
rect 109 1715 119 1733
rect 137 1715 147 1733
rect 109 1709 147 1715
rect 265 1711 299 1774
rect 421 1779 532 1785
rect 421 1771 462 1779
rect 421 1751 429 1771
rect 448 1751 462 1771
rect 421 1749 462 1751
rect 490 1771 532 1779
rect 490 1751 506 1771
rect 525 1751 532 1771
rect 490 1749 532 1751
rect 421 1734 532 1749
rect 759 1780 1204 1800
rect 759 1711 797 1780
rect 1036 1779 1204 1780
rect 1282 1852 1364 1874
rect 1393 1852 1403 1879
rect 1431 1855 1438 1882
rect 1467 1874 1470 1882
rect 3465 1891 3576 1906
rect 3465 1889 3507 1891
rect 1467 1855 1532 1874
rect 1431 1852 1532 1855
rect 1282 1850 1532 1852
rect 1282 1771 1319 1850
rect 1360 1837 1470 1850
rect 1434 1781 1465 1782
rect 1282 1751 1291 1771
rect 1311 1751 1319 1771
rect 1282 1741 1319 1751
rect 1378 1771 1465 1781
rect 1378 1751 1387 1771
rect 1407 1751 1465 1771
rect 1378 1742 1465 1751
rect 1378 1741 1415 1742
rect 109 1705 146 1709
rect 265 1700 797 1711
rect 264 1684 797 1700
rect 1434 1689 1465 1742
rect 1495 1771 1532 1850
rect 1703 1847 2096 1867
rect 2116 1847 2119 1867
rect 3198 1862 3239 1871
rect 1703 1842 2119 1847
rect 2793 1860 2961 1861
rect 3198 1860 3207 1862
rect 1703 1841 2044 1842
rect 1647 1781 1678 1782
rect 1495 1751 1504 1771
rect 1524 1751 1532 1771
rect 1495 1741 1532 1751
rect 1591 1774 1678 1781
rect 1591 1771 1652 1774
rect 1591 1751 1600 1771
rect 1620 1754 1652 1771
rect 1673 1754 1678 1774
rect 1620 1751 1678 1754
rect 1591 1744 1678 1751
rect 1703 1771 1740 1841
rect 2006 1840 2043 1841
rect 2793 1840 3207 1860
rect 3233 1840 3239 1862
rect 3465 1869 3472 1889
rect 3491 1869 3507 1889
rect 3465 1861 3507 1869
rect 3535 1889 3576 1891
rect 3535 1869 3549 1889
rect 3568 1869 3576 1889
rect 3535 1861 3576 1869
rect 3831 1865 3868 1866
rect 4134 1865 4171 1935
rect 4196 1955 4283 1962
rect 4196 1952 4254 1955
rect 4196 1932 4201 1952
rect 4222 1935 4254 1952
rect 4274 1935 4283 1955
rect 4222 1932 4283 1935
rect 4196 1925 4283 1932
rect 4342 1955 4379 1965
rect 4342 1935 4350 1955
rect 4370 1935 4379 1955
rect 4196 1924 4227 1925
rect 3830 1864 4171 1865
rect 3465 1855 3576 1861
rect 3755 1859 4171 1864
rect 2793 1834 3239 1840
rect 2793 1832 2961 1834
rect 1855 1781 1891 1782
rect 1703 1751 1712 1771
rect 1732 1751 1740 1771
rect 1591 1742 1647 1744
rect 1591 1741 1628 1742
rect 1703 1741 1740 1751
rect 1799 1771 1947 1781
rect 2047 1778 2143 1780
rect 1799 1751 1808 1771
rect 1828 1751 1918 1771
rect 1938 1751 1947 1771
rect 1799 1742 1947 1751
rect 2005 1771 2143 1778
rect 2005 1751 2014 1771
rect 2034 1751 2143 1771
rect 2005 1742 2143 1751
rect 1799 1741 1836 1742
rect 1855 1690 1891 1742
rect 1910 1741 1947 1742
rect 2006 1741 2043 1742
rect 1326 1688 1367 1689
rect 264 1683 778 1684
rect 1218 1681 1367 1688
rect 1218 1661 1336 1681
rect 1356 1661 1367 1681
rect 1218 1653 1367 1661
rect 1434 1685 1793 1689
rect 1434 1680 1756 1685
rect 1434 1656 1547 1680
rect 1571 1661 1756 1680
rect 1780 1661 1793 1685
rect 1571 1656 1793 1661
rect 1434 1653 1793 1656
rect 1855 1653 1890 1690
rect 1958 1687 2058 1690
rect 1958 1683 2025 1687
rect 1958 1657 1970 1683
rect 1996 1661 2025 1683
rect 2051 1661 2058 1687
rect 1996 1657 2058 1661
rect 1958 1653 2058 1657
rect 112 1642 149 1643
rect 110 1634 150 1642
rect 110 1616 121 1634
rect 139 1616 150 1634
rect 1434 1632 1465 1653
rect 1855 1632 1891 1653
rect 1277 1631 1314 1632
rect 110 1568 150 1616
rect 1276 1622 1314 1631
rect 1276 1602 1285 1622
rect 1305 1602 1314 1622
rect 1276 1594 1314 1602
rect 1380 1626 1465 1632
rect 1490 1631 1527 1632
rect 1380 1606 1388 1626
rect 1408 1606 1465 1626
rect 1380 1598 1465 1606
rect 1489 1622 1527 1631
rect 1489 1602 1498 1622
rect 1518 1602 1527 1622
rect 1380 1597 1416 1598
rect 1489 1594 1527 1602
rect 1593 1626 1678 1632
rect 1698 1631 1735 1632
rect 1593 1606 1601 1626
rect 1621 1625 1678 1626
rect 1621 1606 1650 1625
rect 1593 1605 1650 1606
rect 1671 1605 1678 1625
rect 1593 1598 1678 1605
rect 1697 1622 1735 1631
rect 1697 1602 1706 1622
rect 1726 1602 1735 1622
rect 1593 1597 1629 1598
rect 1697 1594 1735 1602
rect 1801 1626 1945 1632
rect 1801 1606 1809 1626
rect 1829 1609 1865 1626
rect 1885 1609 1917 1626
rect 1829 1606 1917 1609
rect 1937 1606 1945 1626
rect 1801 1598 1945 1606
rect 1801 1597 1837 1598
rect 1909 1597 1945 1598
rect 2011 1631 2048 1632
rect 2011 1630 2049 1631
rect 2011 1622 2075 1630
rect 2011 1602 2020 1622
rect 2040 1608 2075 1622
rect 2095 1608 2098 1628
rect 2040 1603 2098 1608
rect 2040 1602 2075 1603
rect 421 1572 531 1586
rect 421 1569 464 1572
rect 110 1561 235 1568
rect 421 1564 425 1569
rect 110 1542 202 1561
rect 227 1542 235 1561
rect 110 1532 235 1542
rect 343 1542 425 1564
rect 454 1542 464 1569
rect 492 1545 499 1572
rect 528 1564 531 1572
rect 1277 1565 1314 1594
rect 528 1545 593 1564
rect 1278 1563 1314 1565
rect 1490 1563 1527 1594
rect 1698 1567 1735 1594
rect 2011 1590 2075 1602
rect 492 1542 593 1545
rect 343 1540 593 1542
rect 110 1512 150 1532
rect 109 1503 150 1512
rect 109 1485 119 1503
rect 137 1485 150 1503
rect 109 1476 150 1485
rect 109 1475 146 1476
rect 343 1461 380 1540
rect 421 1527 531 1540
rect 495 1471 526 1472
rect 343 1441 352 1461
rect 372 1441 380 1461
rect 343 1431 380 1441
rect 439 1461 526 1471
rect 439 1441 448 1461
rect 468 1441 526 1461
rect 439 1432 526 1441
rect 439 1431 476 1432
rect 112 1409 149 1413
rect 109 1404 149 1409
rect 109 1386 121 1404
rect 139 1386 149 1404
rect 109 1206 149 1386
rect 495 1379 526 1432
rect 556 1461 593 1540
rect 764 1537 1157 1557
rect 1177 1537 1180 1557
rect 1278 1541 1527 1563
rect 1696 1562 1737 1567
rect 2115 1564 2142 1742
rect 2793 1654 2820 1832
rect 3198 1829 3239 1834
rect 3408 1833 3657 1855
rect 3755 1839 3758 1859
rect 3778 1839 4171 1859
rect 4342 1856 4379 1935
rect 4409 1964 4440 2017
rect 4786 2010 4826 2190
rect 4786 1992 4796 2010
rect 4814 1992 4826 2010
rect 4786 1987 4826 1992
rect 4786 1983 4823 1987
rect 4459 1964 4496 1965
rect 4409 1955 4496 1964
rect 4409 1935 4467 1955
rect 4487 1935 4496 1955
rect 4409 1925 4496 1935
rect 4555 1955 4592 1965
rect 4555 1935 4563 1955
rect 4583 1935 4592 1955
rect 4409 1924 4440 1925
rect 4404 1856 4514 1869
rect 4555 1856 4592 1935
rect 4789 1920 4826 1921
rect 4785 1911 4826 1920
rect 4785 1893 4798 1911
rect 4816 1893 4826 1911
rect 4785 1884 4826 1893
rect 4785 1864 4825 1884
rect 4342 1854 4592 1856
rect 4342 1851 4443 1854
rect 2860 1794 2924 1806
rect 3200 1802 3237 1829
rect 3408 1802 3445 1833
rect 3621 1831 3657 1833
rect 4342 1832 4407 1851
rect 3621 1802 3658 1831
rect 4404 1824 4407 1832
rect 4436 1824 4443 1851
rect 4471 1827 4481 1854
rect 4510 1832 4592 1854
rect 4700 1854 4825 1864
rect 4700 1835 4708 1854
rect 4733 1835 4825 1854
rect 4510 1827 4514 1832
rect 4700 1828 4825 1835
rect 4471 1824 4514 1827
rect 4404 1810 4514 1824
rect 2860 1793 2895 1794
rect 2837 1788 2895 1793
rect 2837 1768 2840 1788
rect 2860 1774 2895 1788
rect 2915 1774 2924 1794
rect 2860 1766 2924 1774
rect 2886 1765 2924 1766
rect 2887 1764 2924 1765
rect 2990 1798 3026 1799
rect 3098 1798 3134 1799
rect 2990 1790 3134 1798
rect 2990 1770 2998 1790
rect 3018 1770 3106 1790
rect 3126 1770 3134 1790
rect 2990 1764 3134 1770
rect 3200 1794 3238 1802
rect 3306 1798 3342 1799
rect 3200 1774 3209 1794
rect 3229 1774 3238 1794
rect 3200 1765 3238 1774
rect 3257 1791 3342 1798
rect 3257 1771 3264 1791
rect 3285 1790 3342 1791
rect 3285 1771 3314 1790
rect 3257 1770 3314 1771
rect 3334 1770 3342 1790
rect 3200 1764 3237 1765
rect 3257 1764 3342 1770
rect 3408 1794 3446 1802
rect 3519 1798 3555 1799
rect 3408 1774 3417 1794
rect 3437 1774 3446 1794
rect 3408 1765 3446 1774
rect 3470 1790 3555 1798
rect 3470 1770 3527 1790
rect 3547 1770 3555 1790
rect 3408 1764 3445 1765
rect 3470 1764 3555 1770
rect 3621 1794 3659 1802
rect 3621 1774 3630 1794
rect 3650 1774 3659 1794
rect 3621 1765 3659 1774
rect 4785 1780 4825 1828
rect 3621 1764 3658 1765
rect 3044 1743 3080 1764
rect 3470 1743 3501 1764
rect 4785 1762 4796 1780
rect 4814 1762 4825 1780
rect 4785 1754 4825 1762
rect 4786 1753 4823 1754
rect 2877 1739 2977 1743
rect 2877 1735 2939 1739
rect 2877 1709 2884 1735
rect 2910 1713 2939 1735
rect 2965 1713 2977 1739
rect 2910 1709 2977 1713
rect 2877 1706 2977 1709
rect 3045 1706 3080 1743
rect 3142 1740 3501 1743
rect 3142 1735 3364 1740
rect 3142 1711 3155 1735
rect 3179 1716 3364 1735
rect 3388 1716 3501 1740
rect 3179 1711 3501 1716
rect 3142 1707 3501 1711
rect 3568 1735 3717 1743
rect 3568 1715 3579 1735
rect 3599 1715 3717 1735
rect 3568 1708 3717 1715
rect 4157 1712 4671 1713
rect 3568 1707 3609 1708
rect 3044 1671 3080 1706
rect 2892 1654 2929 1655
rect 2988 1654 3025 1655
rect 3044 1654 3051 1671
rect 2792 1645 2930 1654
rect 2792 1625 2901 1645
rect 2921 1625 2930 1645
rect 2792 1618 2930 1625
rect 2988 1645 3051 1654
rect 2988 1625 2997 1645
rect 3017 1630 3051 1645
rect 3072 1654 3080 1671
rect 3099 1654 3136 1655
rect 3072 1645 3136 1654
rect 3072 1630 3107 1645
rect 3017 1625 3107 1630
rect 3127 1625 3136 1645
rect 2792 1616 2888 1618
rect 2988 1615 3136 1625
rect 3195 1645 3232 1655
rect 3307 1654 3344 1655
rect 3288 1652 3344 1654
rect 3195 1625 3203 1645
rect 3223 1625 3232 1645
rect 3044 1614 3080 1615
rect 1974 1562 2142 1564
rect 1696 1556 2142 1562
rect 764 1532 1180 1537
rect 1359 1535 1470 1541
rect 764 1531 1105 1532
rect 708 1471 739 1472
rect 556 1441 565 1461
rect 585 1441 593 1461
rect 556 1431 593 1441
rect 652 1464 739 1471
rect 652 1461 713 1464
rect 652 1441 661 1461
rect 681 1444 713 1461
rect 734 1444 739 1464
rect 681 1441 739 1444
rect 652 1434 739 1441
rect 764 1461 801 1531
rect 1067 1530 1104 1531
rect 1359 1527 1400 1535
rect 1359 1507 1367 1527
rect 1386 1507 1400 1527
rect 1359 1505 1400 1507
rect 1428 1527 1470 1535
rect 1428 1507 1444 1527
rect 1463 1507 1470 1527
rect 1696 1534 1702 1556
rect 1728 1536 2142 1556
rect 2892 1555 2929 1556
rect 3195 1555 3232 1625
rect 3257 1645 3344 1652
rect 3257 1642 3315 1645
rect 3257 1622 3262 1642
rect 3283 1625 3315 1642
rect 3335 1625 3344 1645
rect 3283 1622 3344 1625
rect 3257 1615 3344 1622
rect 3403 1645 3440 1655
rect 3403 1625 3411 1645
rect 3431 1625 3440 1645
rect 3257 1614 3288 1615
rect 2891 1554 3232 1555
rect 1728 1534 1737 1536
rect 1974 1535 2142 1536
rect 2816 1553 3232 1554
rect 2816 1549 3192 1553
rect 1696 1525 1737 1534
rect 2816 1529 2819 1549
rect 2839 1536 3192 1549
rect 3224 1536 3232 1553
rect 2839 1529 3232 1536
rect 3403 1546 3440 1625
rect 3470 1654 3501 1707
rect 4138 1696 4671 1712
rect 4138 1685 4670 1696
rect 4789 1687 4826 1691
rect 3520 1654 3557 1655
rect 3470 1645 3557 1654
rect 3470 1625 3528 1645
rect 3548 1625 3557 1645
rect 3470 1615 3557 1625
rect 3616 1645 3653 1655
rect 3616 1625 3624 1645
rect 3644 1625 3653 1645
rect 3470 1614 3501 1615
rect 3465 1546 3575 1559
rect 3616 1546 3653 1625
rect 3403 1544 3653 1546
rect 3403 1541 3504 1544
rect 3403 1522 3468 1541
rect 1428 1505 1470 1507
rect 1359 1490 1470 1505
rect 3465 1514 3468 1522
rect 3497 1514 3504 1541
rect 3532 1517 3542 1544
rect 3571 1522 3653 1544
rect 3731 1616 3899 1617
rect 4138 1616 4176 1685
rect 3731 1596 4176 1616
rect 4403 1647 4514 1662
rect 4403 1645 4445 1647
rect 4403 1625 4410 1645
rect 4429 1625 4445 1645
rect 4403 1617 4445 1625
rect 4473 1645 4514 1647
rect 4473 1625 4487 1645
rect 4506 1625 4514 1645
rect 4473 1617 4514 1625
rect 4403 1611 4514 1617
rect 4636 1622 4670 1685
rect 4788 1681 4826 1687
rect 4788 1663 4798 1681
rect 4816 1663 4826 1681
rect 4788 1654 4826 1663
rect 4788 1622 4822 1654
rect 3731 1590 4175 1596
rect 3731 1588 3899 1590
rect 3571 1517 3575 1522
rect 3532 1514 3575 1517
rect 3465 1500 3575 1514
rect 916 1471 952 1472
rect 764 1441 773 1461
rect 793 1441 801 1461
rect 652 1432 708 1434
rect 652 1431 689 1432
rect 764 1431 801 1441
rect 860 1461 1008 1471
rect 1108 1468 1204 1470
rect 860 1441 869 1461
rect 889 1441 979 1461
rect 999 1441 1008 1461
rect 860 1432 1008 1441
rect 1066 1461 1204 1468
rect 1066 1441 1075 1461
rect 1095 1441 1204 1461
rect 1066 1432 1204 1441
rect 860 1431 897 1432
rect 916 1380 952 1432
rect 971 1431 1008 1432
rect 1067 1431 1104 1432
rect 387 1378 428 1379
rect 279 1371 428 1378
rect 279 1351 397 1371
rect 417 1351 428 1371
rect 279 1343 428 1351
rect 495 1375 854 1379
rect 495 1370 817 1375
rect 495 1346 608 1370
rect 632 1351 817 1370
rect 841 1351 854 1375
rect 632 1346 854 1351
rect 495 1343 854 1346
rect 916 1343 951 1380
rect 1019 1377 1119 1380
rect 1019 1373 1086 1377
rect 1019 1347 1031 1373
rect 1057 1351 1086 1373
rect 1112 1351 1119 1377
rect 1057 1347 1119 1351
rect 1019 1343 1119 1347
rect 495 1322 526 1343
rect 916 1322 952 1343
rect 338 1321 375 1322
rect 337 1312 375 1321
rect 337 1292 346 1312
rect 366 1292 375 1312
rect 337 1284 375 1292
rect 441 1316 526 1322
rect 551 1321 588 1322
rect 441 1296 449 1316
rect 469 1296 526 1316
rect 441 1288 526 1296
rect 550 1312 588 1321
rect 550 1292 559 1312
rect 579 1292 588 1312
rect 441 1287 477 1288
rect 550 1284 588 1292
rect 654 1316 739 1322
rect 759 1321 796 1322
rect 654 1296 662 1316
rect 682 1315 739 1316
rect 682 1296 711 1315
rect 654 1295 711 1296
rect 732 1295 739 1315
rect 654 1288 739 1295
rect 758 1312 796 1321
rect 758 1292 767 1312
rect 787 1292 796 1312
rect 654 1287 690 1288
rect 758 1284 796 1292
rect 862 1316 1006 1322
rect 862 1296 870 1316
rect 890 1313 978 1316
rect 890 1296 921 1313
rect 862 1293 921 1296
rect 944 1296 978 1313
rect 998 1296 1006 1316
rect 944 1293 1006 1296
rect 862 1288 1006 1293
rect 862 1287 898 1288
rect 970 1287 1006 1288
rect 1072 1321 1109 1322
rect 1072 1320 1110 1321
rect 1072 1312 1136 1320
rect 1072 1292 1081 1312
rect 1101 1298 1136 1312
rect 1156 1298 1159 1318
rect 1101 1293 1159 1298
rect 1101 1292 1136 1293
rect 338 1255 375 1284
rect 339 1253 375 1255
rect 551 1253 588 1284
rect 339 1231 588 1253
rect 759 1252 796 1284
rect 1072 1280 1136 1292
rect 1176 1254 1203 1432
rect 3731 1410 3758 1588
rect 3798 1550 3862 1562
rect 4138 1558 4175 1590
rect 4346 1589 4595 1611
rect 4636 1590 4822 1622
rect 4650 1589 4822 1590
rect 4346 1558 4383 1589
rect 4559 1587 4595 1589
rect 4559 1558 4596 1587
rect 4788 1561 4822 1589
rect 3798 1549 3833 1550
rect 3775 1544 3833 1549
rect 3775 1524 3778 1544
rect 3798 1530 3833 1544
rect 3853 1530 3862 1550
rect 3798 1522 3862 1530
rect 3824 1521 3862 1522
rect 3825 1520 3862 1521
rect 3928 1554 3964 1555
rect 4036 1554 4072 1555
rect 3928 1547 4072 1554
rect 3928 1546 3988 1547
rect 3928 1526 3936 1546
rect 3956 1527 3988 1546
rect 4013 1546 4072 1547
rect 4013 1527 4044 1546
rect 3956 1526 4044 1527
rect 4064 1526 4072 1546
rect 3928 1520 4072 1526
rect 4138 1550 4176 1558
rect 4244 1554 4280 1555
rect 4138 1530 4147 1550
rect 4167 1530 4176 1550
rect 4138 1521 4176 1530
rect 4195 1547 4280 1554
rect 4195 1527 4202 1547
rect 4223 1546 4280 1547
rect 4223 1527 4252 1546
rect 4195 1526 4252 1527
rect 4272 1526 4280 1546
rect 4138 1520 4175 1521
rect 4195 1520 4280 1526
rect 4346 1550 4384 1558
rect 4457 1554 4493 1555
rect 4346 1530 4355 1550
rect 4375 1530 4384 1550
rect 4346 1521 4384 1530
rect 4408 1546 4493 1554
rect 4408 1526 4465 1546
rect 4485 1526 4493 1546
rect 4346 1520 4383 1521
rect 4408 1520 4493 1526
rect 4559 1550 4597 1558
rect 4559 1530 4568 1550
rect 4588 1530 4597 1550
rect 4559 1521 4597 1530
rect 4786 1551 4823 1561
rect 4786 1533 4796 1551
rect 4814 1533 4823 1551
rect 4786 1524 4823 1533
rect 4788 1523 4822 1524
rect 4559 1520 4596 1521
rect 3982 1499 4018 1520
rect 4408 1499 4439 1520
rect 3815 1495 3915 1499
rect 3815 1491 3877 1495
rect 3815 1465 3822 1491
rect 3848 1469 3877 1491
rect 3903 1469 3915 1495
rect 3848 1465 3915 1469
rect 3815 1462 3915 1465
rect 3983 1462 4018 1499
rect 4080 1496 4439 1499
rect 4080 1491 4302 1496
rect 4080 1467 4093 1491
rect 4117 1472 4302 1491
rect 4326 1472 4439 1496
rect 4117 1467 4439 1472
rect 4080 1463 4439 1467
rect 4506 1491 4655 1499
rect 4506 1471 4517 1491
rect 4537 1471 4655 1491
rect 4506 1464 4655 1471
rect 4506 1463 4547 1464
rect 3830 1410 3867 1411
rect 3926 1410 3963 1411
rect 3982 1410 4018 1462
rect 4037 1410 4074 1411
rect 3730 1401 3868 1410
rect 3325 1380 3436 1395
rect 3325 1378 3367 1380
rect 2995 1357 3100 1359
rect 2653 1349 2821 1350
rect 2995 1349 3044 1357
rect 2653 1330 3044 1349
rect 3075 1330 3100 1357
rect 3325 1358 3332 1378
rect 3351 1358 3367 1378
rect 3325 1350 3367 1358
rect 3395 1378 3436 1380
rect 3395 1358 3409 1378
rect 3428 1358 3436 1378
rect 3730 1381 3839 1401
rect 3859 1381 3868 1401
rect 3730 1374 3868 1381
rect 3926 1401 4074 1410
rect 3926 1381 3935 1401
rect 3955 1381 4045 1401
rect 4065 1381 4074 1401
rect 3730 1372 3826 1374
rect 3926 1371 4074 1381
rect 4133 1401 4170 1411
rect 4245 1410 4282 1411
rect 4226 1408 4282 1410
rect 4133 1381 4141 1401
rect 4161 1381 4170 1401
rect 3982 1370 4018 1371
rect 3395 1350 3436 1358
rect 3325 1344 3436 1350
rect 2653 1323 3100 1330
rect 2653 1321 2821 1323
rect 1501 1290 1611 1304
rect 1501 1287 1544 1290
rect 1501 1282 1505 1287
rect 1035 1252 1203 1254
rect 759 1249 1203 1252
rect 420 1225 531 1231
rect 420 1217 461 1225
rect 109 1162 148 1206
rect 420 1197 428 1217
rect 447 1197 461 1217
rect 420 1195 461 1197
rect 489 1217 531 1225
rect 489 1197 505 1217
rect 524 1197 531 1217
rect 489 1195 531 1197
rect 420 1180 531 1195
rect 757 1226 1203 1249
rect 109 1138 149 1162
rect 449 1138 496 1140
rect 757 1138 795 1226
rect 1035 1225 1203 1226
rect 1423 1260 1505 1282
rect 1534 1260 1544 1287
rect 1572 1263 1579 1290
rect 1608 1282 1611 1290
rect 1608 1263 1673 1282
rect 1572 1260 1673 1263
rect 1423 1258 1673 1260
rect 1423 1179 1460 1258
rect 1501 1245 1611 1258
rect 1575 1189 1606 1190
rect 1423 1159 1432 1179
rect 1452 1159 1460 1179
rect 1423 1149 1460 1159
rect 1519 1179 1606 1189
rect 1519 1159 1528 1179
rect 1548 1159 1606 1179
rect 1519 1150 1606 1159
rect 1519 1149 1556 1150
rect 109 1105 795 1138
rect 109 1048 148 1105
rect 757 1103 795 1105
rect 1575 1097 1606 1150
rect 1636 1179 1673 1258
rect 1844 1271 2237 1275
rect 1844 1254 1863 1271
rect 1883 1255 2237 1271
rect 2257 1255 2260 1275
rect 1883 1254 2260 1255
rect 1844 1250 2260 1254
rect 1844 1249 2185 1250
rect 1788 1189 1819 1190
rect 1636 1159 1645 1179
rect 1665 1159 1673 1179
rect 1636 1149 1673 1159
rect 1732 1182 1819 1189
rect 1732 1179 1793 1182
rect 1732 1159 1741 1179
rect 1761 1162 1793 1179
rect 1814 1162 1819 1182
rect 1761 1159 1819 1162
rect 1732 1152 1819 1159
rect 1844 1179 1881 1249
rect 2147 1248 2184 1249
rect 1996 1189 2032 1190
rect 1844 1159 1853 1179
rect 1873 1159 1881 1179
rect 1732 1150 1788 1152
rect 1732 1149 1769 1150
rect 1844 1149 1881 1159
rect 1940 1179 2088 1189
rect 2256 1188 2285 1189
rect 2188 1186 2285 1188
rect 1940 1159 1949 1179
rect 1969 1175 2059 1179
rect 1969 1159 2002 1175
rect 1940 1150 2002 1159
rect 1940 1149 1977 1150
rect 1996 1137 2002 1150
rect 2025 1159 2059 1175
rect 2079 1159 2088 1179
rect 2025 1150 2088 1159
rect 2146 1179 2285 1186
rect 2146 1159 2155 1179
rect 2175 1159 2285 1179
rect 2146 1150 2285 1159
rect 2025 1137 2032 1150
rect 2051 1149 2088 1150
rect 2147 1149 2184 1150
rect 1996 1098 2032 1137
rect 1467 1096 1508 1097
rect 1359 1089 1508 1096
rect 1359 1069 1477 1089
rect 1497 1069 1508 1089
rect 1359 1061 1508 1069
rect 1575 1093 1934 1097
rect 1575 1088 1897 1093
rect 1575 1064 1688 1088
rect 1712 1069 1897 1088
rect 1921 1069 1934 1093
rect 1712 1064 1934 1069
rect 1575 1061 1934 1064
rect 1996 1061 2031 1098
rect 2099 1095 2199 1098
rect 2099 1091 2166 1095
rect 2099 1065 2111 1091
rect 2137 1069 2166 1091
rect 2192 1069 2199 1095
rect 2137 1065 2199 1069
rect 2099 1061 2199 1065
rect 109 1046 157 1048
rect 109 1028 120 1046
rect 138 1028 157 1046
rect 1575 1040 1606 1061
rect 1996 1040 2032 1061
rect 1418 1039 1455 1040
rect 109 1019 157 1028
rect 110 1018 157 1019
rect 423 1023 533 1037
rect 423 1020 466 1023
rect 423 1015 427 1020
rect 345 993 427 1015
rect 456 993 466 1020
rect 494 996 501 1023
rect 530 1015 533 1023
rect 1417 1030 1455 1039
rect 530 996 595 1015
rect 1417 1010 1426 1030
rect 1446 1010 1455 1030
rect 494 993 595 996
rect 345 991 595 993
rect 113 955 150 956
rect 109 952 150 955
rect 109 947 151 952
rect 109 929 122 947
rect 140 929 151 947
rect 109 915 151 929
rect 189 915 236 919
rect 109 909 236 915
rect 109 880 197 909
rect 226 880 236 909
rect 345 912 382 991
rect 423 978 533 991
rect 497 922 528 923
rect 345 892 354 912
rect 374 892 382 912
rect 345 882 382 892
rect 441 912 528 922
rect 441 892 450 912
rect 470 892 528 912
rect 441 883 528 892
rect 441 882 478 883
rect 109 876 236 880
rect 109 859 148 876
rect 189 875 236 876
rect 109 841 120 859
rect 138 841 148 859
rect 109 832 148 841
rect 110 831 147 832
rect 497 830 528 883
rect 558 912 595 991
rect 766 988 1159 1008
rect 1179 988 1182 1008
rect 1417 1002 1455 1010
rect 1521 1034 1606 1040
rect 1631 1039 1668 1040
rect 1521 1014 1529 1034
rect 1549 1014 1606 1034
rect 1521 1006 1606 1014
rect 1630 1030 1668 1039
rect 1630 1010 1639 1030
rect 1659 1010 1668 1030
rect 1521 1005 1557 1006
rect 1630 1002 1668 1010
rect 1734 1034 1819 1040
rect 1839 1039 1876 1040
rect 1734 1014 1742 1034
rect 1762 1033 1819 1034
rect 1762 1014 1791 1033
rect 1734 1013 1791 1014
rect 1812 1013 1819 1033
rect 1734 1006 1819 1013
rect 1838 1030 1876 1039
rect 1838 1010 1847 1030
rect 1867 1010 1876 1030
rect 1734 1005 1770 1006
rect 1838 1002 1876 1010
rect 1942 1034 2086 1040
rect 1942 1014 1950 1034
rect 1970 1014 2058 1034
rect 2078 1014 2086 1034
rect 1942 1006 2086 1014
rect 1942 1005 1978 1006
rect 2050 1005 2086 1006
rect 2152 1039 2189 1040
rect 2152 1038 2190 1039
rect 2152 1030 2216 1038
rect 2152 1010 2161 1030
rect 2181 1016 2216 1030
rect 2236 1016 2239 1036
rect 2181 1011 2239 1016
rect 2181 1010 2216 1011
rect 766 983 1182 988
rect 766 982 1107 983
rect 710 922 741 923
rect 558 892 567 912
rect 587 892 595 912
rect 558 882 595 892
rect 654 915 741 922
rect 654 912 715 915
rect 654 892 663 912
rect 683 895 715 912
rect 736 895 741 915
rect 683 892 741 895
rect 654 885 741 892
rect 766 912 803 982
rect 1069 981 1106 982
rect 1418 973 1455 1002
rect 1419 971 1455 973
rect 1631 971 1668 1002
rect 1419 949 1668 971
rect 1839 970 1876 1002
rect 2152 998 2216 1010
rect 2256 972 2285 1150
rect 2653 1143 2680 1321
rect 2720 1283 2784 1295
rect 3060 1291 3097 1323
rect 3268 1322 3517 1344
rect 3268 1291 3305 1322
rect 3481 1320 3517 1322
rect 3481 1291 3518 1320
rect 3830 1311 3867 1312
rect 4133 1311 4170 1381
rect 4195 1401 4282 1408
rect 4195 1398 4253 1401
rect 4195 1378 4200 1398
rect 4221 1381 4253 1398
rect 4273 1381 4282 1401
rect 4221 1378 4282 1381
rect 4195 1371 4282 1378
rect 4341 1401 4378 1411
rect 4341 1381 4349 1401
rect 4369 1381 4378 1401
rect 4195 1370 4226 1371
rect 3829 1310 4170 1311
rect 3754 1305 4170 1310
rect 2720 1282 2755 1283
rect 2697 1277 2755 1282
rect 2697 1257 2700 1277
rect 2720 1263 2755 1277
rect 2775 1263 2784 1283
rect 2720 1255 2784 1263
rect 2746 1254 2784 1255
rect 2747 1253 2784 1254
rect 2850 1287 2886 1288
rect 2958 1287 2994 1288
rect 2850 1282 2994 1287
rect 2850 1279 2910 1282
rect 2850 1259 2858 1279
rect 2878 1261 2910 1279
rect 2937 1279 2994 1282
rect 2937 1261 2966 1279
rect 2878 1259 2966 1261
rect 2986 1259 2994 1279
rect 2850 1253 2994 1259
rect 3060 1283 3098 1291
rect 3166 1287 3202 1288
rect 3060 1263 3069 1283
rect 3089 1263 3098 1283
rect 3060 1254 3098 1263
rect 3117 1280 3202 1287
rect 3117 1260 3124 1280
rect 3145 1279 3202 1280
rect 3145 1260 3174 1279
rect 3117 1259 3174 1260
rect 3194 1259 3202 1279
rect 3060 1253 3097 1254
rect 3117 1253 3202 1259
rect 3268 1283 3306 1291
rect 3379 1287 3415 1288
rect 3268 1263 3277 1283
rect 3297 1263 3306 1283
rect 3268 1254 3306 1263
rect 3330 1279 3415 1287
rect 3330 1259 3387 1279
rect 3407 1259 3415 1279
rect 3268 1253 3305 1254
rect 3330 1253 3415 1259
rect 3481 1283 3519 1291
rect 3754 1285 3757 1305
rect 3777 1285 4170 1305
rect 4341 1302 4378 1381
rect 4408 1410 4439 1463
rect 4789 1461 4826 1462
rect 4788 1452 4827 1461
rect 4788 1434 4798 1452
rect 4816 1434 4827 1452
rect 4700 1417 4747 1418
rect 4788 1417 4827 1434
rect 4700 1413 4827 1417
rect 4458 1410 4495 1411
rect 4408 1401 4495 1410
rect 4408 1381 4466 1401
rect 4486 1381 4495 1401
rect 4408 1371 4495 1381
rect 4554 1401 4591 1411
rect 4554 1381 4562 1401
rect 4582 1381 4591 1401
rect 4408 1370 4439 1371
rect 4403 1302 4513 1315
rect 4554 1302 4591 1381
rect 4700 1384 4710 1413
rect 4739 1384 4827 1413
rect 4700 1378 4827 1384
rect 4700 1374 4747 1378
rect 4785 1364 4827 1378
rect 4785 1346 4796 1364
rect 4814 1346 4827 1364
rect 4785 1341 4827 1346
rect 4786 1338 4827 1341
rect 4786 1337 4823 1338
rect 4341 1300 4591 1302
rect 4341 1297 4442 1300
rect 3481 1263 3490 1283
rect 3510 1263 3519 1283
rect 4341 1278 4406 1297
rect 3481 1254 3519 1263
rect 4403 1270 4406 1278
rect 4435 1270 4442 1297
rect 4470 1273 4480 1300
rect 4509 1278 4591 1300
rect 4509 1273 4513 1278
rect 4470 1270 4513 1273
rect 4403 1256 4513 1270
rect 4779 1274 4826 1275
rect 4779 1265 4827 1274
rect 3481 1253 3518 1254
rect 2904 1232 2940 1253
rect 3330 1232 3361 1253
rect 4779 1247 4798 1265
rect 4816 1247 4827 1265
rect 4779 1245 4827 1247
rect 2737 1228 2837 1232
rect 2737 1224 2799 1228
rect 2737 1198 2744 1224
rect 2770 1202 2799 1224
rect 2825 1202 2837 1228
rect 2770 1198 2837 1202
rect 2737 1195 2837 1198
rect 2905 1195 2940 1232
rect 3002 1229 3361 1232
rect 3002 1224 3224 1229
rect 3002 1200 3015 1224
rect 3039 1205 3224 1224
rect 3248 1205 3361 1229
rect 3039 1200 3361 1205
rect 3002 1196 3361 1200
rect 3428 1224 3577 1232
rect 3428 1204 3439 1224
rect 3459 1204 3577 1224
rect 3428 1197 3577 1204
rect 3428 1196 3469 1197
rect 2752 1143 2789 1144
rect 2848 1143 2885 1144
rect 2904 1143 2940 1195
rect 2959 1143 2996 1144
rect 2652 1134 2790 1143
rect 2652 1114 2761 1134
rect 2781 1114 2790 1134
rect 2652 1107 2790 1114
rect 2848 1134 2996 1143
rect 2848 1114 2857 1134
rect 2877 1114 2967 1134
rect 2987 1114 2996 1134
rect 2652 1105 2748 1107
rect 2848 1104 2996 1114
rect 3055 1134 3092 1144
rect 3167 1143 3204 1144
rect 3148 1141 3204 1143
rect 3055 1114 3063 1134
rect 3083 1114 3092 1134
rect 2904 1103 2940 1104
rect 2752 1044 2789 1045
rect 3055 1044 3092 1114
rect 3117 1134 3204 1141
rect 3117 1131 3175 1134
rect 3117 1111 3122 1131
rect 3143 1114 3175 1131
rect 3195 1114 3204 1134
rect 3143 1111 3204 1114
rect 3117 1104 3204 1111
rect 3263 1134 3300 1144
rect 3263 1114 3271 1134
rect 3291 1114 3300 1134
rect 3117 1103 3148 1104
rect 2751 1043 3092 1044
rect 2676 1039 3092 1043
rect 2676 1038 3053 1039
rect 2676 1018 2679 1038
rect 2699 1022 3053 1038
rect 3073 1022 3092 1039
rect 2699 1018 3092 1022
rect 3263 1035 3300 1114
rect 3330 1143 3361 1196
rect 4141 1188 4179 1190
rect 4788 1188 4827 1245
rect 4141 1155 4827 1188
rect 3380 1143 3417 1144
rect 3330 1134 3417 1143
rect 3330 1114 3388 1134
rect 3408 1114 3417 1134
rect 3330 1104 3417 1114
rect 3476 1134 3513 1144
rect 3476 1114 3484 1134
rect 3504 1114 3513 1134
rect 3330 1103 3361 1104
rect 3325 1035 3435 1048
rect 3476 1035 3513 1114
rect 3263 1033 3513 1035
rect 3263 1030 3364 1033
rect 3263 1011 3328 1030
rect 3325 1003 3328 1011
rect 3357 1003 3364 1030
rect 3392 1006 3402 1033
rect 3431 1011 3513 1033
rect 3733 1067 3901 1068
rect 4141 1067 4179 1155
rect 4440 1153 4487 1155
rect 4787 1131 4827 1155
rect 3733 1044 4179 1067
rect 4405 1098 4516 1113
rect 4405 1096 4447 1098
rect 4405 1076 4412 1096
rect 4431 1076 4447 1096
rect 4405 1068 4447 1076
rect 4475 1096 4516 1098
rect 4475 1076 4489 1096
rect 4508 1076 4516 1096
rect 4788 1087 4827 1131
rect 4475 1068 4516 1076
rect 4405 1062 4516 1068
rect 3733 1041 4177 1044
rect 3733 1039 3901 1041
rect 3431 1006 3435 1011
rect 3392 1003 3435 1006
rect 3325 989 3435 1003
rect 2115 970 2285 972
rect 1836 963 2285 970
rect 1500 943 1611 949
rect 1500 935 1541 943
rect 918 922 954 923
rect 766 892 775 912
rect 795 892 803 912
rect 654 883 710 885
rect 654 882 691 883
rect 766 882 803 892
rect 862 912 1010 922
rect 1110 919 1206 921
rect 862 892 871 912
rect 891 892 981 912
rect 1001 892 1010 912
rect 862 883 1010 892
rect 1068 912 1206 919
rect 1068 892 1077 912
rect 1097 892 1206 912
rect 1500 915 1508 935
rect 1527 915 1541 935
rect 1500 913 1541 915
rect 1569 935 1611 943
rect 1569 915 1585 935
rect 1604 915 1611 935
rect 1836 936 1861 963
rect 1892 944 2285 963
rect 1892 936 1941 944
rect 2115 943 2285 944
rect 1836 934 1941 936
rect 1569 913 1611 915
rect 1500 898 1611 913
rect 1068 883 1206 892
rect 862 882 899 883
rect 918 831 954 883
rect 973 882 1010 883
rect 1069 882 1106 883
rect 389 829 430 830
rect 281 822 430 829
rect 281 802 399 822
rect 419 802 430 822
rect 281 794 430 802
rect 497 826 856 830
rect 497 821 819 826
rect 497 797 610 821
rect 634 802 819 821
rect 843 802 856 826
rect 634 797 856 802
rect 497 794 856 797
rect 918 794 953 831
rect 1021 828 1121 831
rect 1021 824 1088 828
rect 1021 798 1033 824
rect 1059 802 1088 824
rect 1114 802 1121 828
rect 1059 798 1121 802
rect 1021 794 1121 798
rect 497 773 528 794
rect 918 773 954 794
rect 340 772 377 773
rect 114 769 148 770
rect 113 760 150 769
rect 113 742 122 760
rect 140 742 150 760
rect 113 732 150 742
rect 339 763 377 772
rect 339 743 348 763
rect 368 743 377 763
rect 339 735 377 743
rect 443 767 528 773
rect 553 772 590 773
rect 443 747 451 767
rect 471 747 528 767
rect 443 739 528 747
rect 552 763 590 772
rect 552 743 561 763
rect 581 743 590 763
rect 443 738 479 739
rect 552 735 590 743
rect 656 767 741 773
rect 761 772 798 773
rect 656 747 664 767
rect 684 766 741 767
rect 684 747 713 766
rect 656 746 713 747
rect 734 746 741 766
rect 656 739 741 746
rect 760 763 798 772
rect 760 743 769 763
rect 789 743 798 763
rect 656 738 692 739
rect 760 735 798 743
rect 864 767 1008 773
rect 864 747 872 767
rect 892 766 980 767
rect 892 747 923 766
rect 864 746 923 747
rect 948 747 980 766
rect 1000 747 1008 767
rect 948 746 1008 747
rect 864 739 1008 746
rect 864 738 900 739
rect 972 738 1008 739
rect 1074 772 1111 773
rect 1074 771 1112 772
rect 1074 763 1138 771
rect 1074 743 1083 763
rect 1103 749 1138 763
rect 1158 749 1161 769
rect 1103 744 1161 749
rect 1103 743 1138 744
rect 114 704 148 732
rect 340 706 377 735
rect 341 704 377 706
rect 553 704 590 735
rect 114 703 286 704
rect 114 671 300 703
rect 341 682 590 704
rect 761 703 798 735
rect 1074 731 1138 743
rect 1178 705 1205 883
rect 3733 861 3760 1039
rect 3800 1001 3864 1013
rect 4140 1009 4177 1041
rect 4348 1040 4597 1062
rect 4348 1009 4385 1040
rect 4561 1038 4597 1040
rect 4561 1009 4598 1038
rect 3800 1000 3835 1001
rect 3777 995 3835 1000
rect 3777 975 3780 995
rect 3800 981 3835 995
rect 3855 981 3864 1001
rect 3800 973 3864 981
rect 3826 972 3864 973
rect 3827 971 3864 972
rect 3930 1005 3966 1006
rect 4038 1005 4074 1006
rect 3930 1000 4074 1005
rect 3930 997 3992 1000
rect 3930 977 3938 997
rect 3958 980 3992 997
rect 4015 997 4074 1000
rect 4015 980 4046 997
rect 3958 977 4046 980
rect 4066 977 4074 997
rect 3930 971 4074 977
rect 4140 1001 4178 1009
rect 4246 1005 4282 1006
rect 4140 981 4149 1001
rect 4169 981 4178 1001
rect 4140 972 4178 981
rect 4197 998 4282 1005
rect 4197 978 4204 998
rect 4225 997 4282 998
rect 4225 978 4254 997
rect 4197 977 4254 978
rect 4274 977 4282 997
rect 4140 971 4177 972
rect 4197 971 4282 977
rect 4348 1001 4386 1009
rect 4459 1005 4495 1006
rect 4348 981 4357 1001
rect 4377 981 4386 1001
rect 4348 972 4386 981
rect 4410 997 4495 1005
rect 4410 977 4467 997
rect 4487 977 4495 997
rect 4348 971 4385 972
rect 4410 971 4495 977
rect 4561 1001 4599 1009
rect 4561 981 4570 1001
rect 4590 981 4599 1001
rect 4561 972 4599 981
rect 4561 971 4598 972
rect 3984 950 4020 971
rect 4410 950 4441 971
rect 3817 946 3917 950
rect 3817 942 3879 946
rect 3817 916 3824 942
rect 3850 920 3879 942
rect 3905 920 3917 946
rect 3850 916 3917 920
rect 3817 913 3917 916
rect 3985 913 4020 950
rect 4082 947 4441 950
rect 4082 942 4304 947
rect 4082 918 4095 942
rect 4119 923 4304 942
rect 4328 923 4441 947
rect 4119 918 4441 923
rect 4082 914 4441 918
rect 4508 942 4657 950
rect 4508 922 4519 942
rect 4539 922 4657 942
rect 4508 915 4657 922
rect 4508 914 4549 915
rect 3832 861 3869 862
rect 3928 861 3965 862
rect 3984 861 4020 913
rect 4039 861 4076 862
rect 3732 852 3870 861
rect 3732 832 3841 852
rect 3861 832 3870 852
rect 3732 825 3870 832
rect 3928 852 4076 861
rect 3928 832 3937 852
rect 3957 832 4047 852
rect 4067 832 4076 852
rect 3732 823 3828 825
rect 3928 822 4076 832
rect 4135 852 4172 862
rect 4247 861 4284 862
rect 4228 859 4284 861
rect 4135 832 4143 852
rect 4163 832 4172 852
rect 3984 821 4020 822
rect 1361 779 1471 793
rect 1361 776 1404 779
rect 1361 771 1365 776
rect 1037 703 1205 705
rect 761 697 1205 703
rect 114 639 148 671
rect 110 630 148 639
rect 110 612 120 630
rect 138 612 148 630
rect 110 606 148 612
rect 266 608 300 671
rect 422 676 533 682
rect 422 668 463 676
rect 422 648 430 668
rect 449 648 463 668
rect 422 646 463 648
rect 491 668 533 676
rect 491 648 507 668
rect 526 648 533 668
rect 491 646 533 648
rect 422 631 533 646
rect 760 677 1205 697
rect 760 608 798 677
rect 1037 676 1205 677
rect 1283 749 1365 771
rect 1394 749 1404 776
rect 1432 752 1439 779
rect 1468 771 1471 779
rect 3466 788 3577 803
rect 3466 786 3508 788
rect 1468 752 1533 771
rect 1432 749 1533 752
rect 1283 747 1533 749
rect 1283 668 1320 747
rect 1361 734 1471 747
rect 1435 678 1466 679
rect 1283 648 1292 668
rect 1312 648 1320 668
rect 1283 638 1320 648
rect 1379 668 1466 678
rect 1379 648 1388 668
rect 1408 648 1466 668
rect 1379 639 1466 648
rect 1379 638 1416 639
rect 110 602 147 606
rect 266 597 798 608
rect 265 581 798 597
rect 1435 586 1466 639
rect 1496 668 1533 747
rect 1704 757 2097 764
rect 1704 740 1712 757
rect 1744 744 2097 757
rect 2117 744 2120 764
rect 3199 759 3240 768
rect 1744 740 2120 744
rect 1704 739 2120 740
rect 2794 757 2962 758
rect 3199 757 3208 759
rect 1704 738 2045 739
rect 1648 678 1679 679
rect 1496 648 1505 668
rect 1525 648 1533 668
rect 1496 638 1533 648
rect 1592 671 1679 678
rect 1592 668 1653 671
rect 1592 648 1601 668
rect 1621 651 1653 668
rect 1674 651 1679 671
rect 1621 648 1679 651
rect 1592 641 1679 648
rect 1704 668 1741 738
rect 2007 737 2044 738
rect 2794 737 3208 757
rect 3234 737 3240 759
rect 3466 766 3473 786
rect 3492 766 3508 786
rect 3466 758 3508 766
rect 3536 786 3577 788
rect 3536 766 3550 786
rect 3569 766 3577 786
rect 3536 758 3577 766
rect 3832 762 3869 763
rect 4135 762 4172 832
rect 4197 852 4284 859
rect 4197 849 4255 852
rect 4197 829 4202 849
rect 4223 832 4255 849
rect 4275 832 4284 852
rect 4223 829 4284 832
rect 4197 822 4284 829
rect 4343 852 4380 862
rect 4343 832 4351 852
rect 4371 832 4380 852
rect 4197 821 4228 822
rect 3831 761 4172 762
rect 3466 752 3577 758
rect 3756 756 4172 761
rect 2794 731 3240 737
rect 2794 729 2962 731
rect 1856 678 1892 679
rect 1704 648 1713 668
rect 1733 648 1741 668
rect 1592 639 1648 641
rect 1592 638 1629 639
rect 1704 638 1741 648
rect 1800 668 1948 678
rect 2048 675 2144 677
rect 1800 648 1809 668
rect 1829 663 1919 668
rect 1829 648 1864 663
rect 1800 639 1864 648
rect 1800 638 1837 639
rect 1856 622 1864 639
rect 1885 648 1919 663
rect 1939 648 1948 668
rect 1885 639 1948 648
rect 2006 668 2144 675
rect 2006 648 2015 668
rect 2035 648 2144 668
rect 2006 639 2144 648
rect 1885 622 1892 639
rect 1911 638 1948 639
rect 2007 638 2044 639
rect 1856 587 1892 622
rect 1327 585 1368 586
rect 265 580 779 581
rect 1219 578 1368 585
rect 1219 558 1337 578
rect 1357 558 1368 578
rect 1219 550 1368 558
rect 1435 582 1794 586
rect 1435 577 1757 582
rect 1435 553 1548 577
rect 1572 558 1757 577
rect 1781 558 1794 582
rect 1572 553 1794 558
rect 1435 550 1794 553
rect 1856 550 1891 587
rect 1959 584 2059 587
rect 1959 580 2026 584
rect 1959 554 1971 580
rect 1997 558 2026 580
rect 2052 558 2059 584
rect 1997 554 2059 558
rect 1959 550 2059 554
rect 113 539 150 540
rect 111 531 151 539
rect 111 513 122 531
rect 140 513 151 531
rect 1435 529 1466 550
rect 1856 529 1892 550
rect 1278 528 1315 529
rect 111 465 151 513
rect 1277 519 1315 528
rect 1277 499 1286 519
rect 1306 499 1315 519
rect 1277 491 1315 499
rect 1381 523 1466 529
rect 1491 528 1528 529
rect 1381 503 1389 523
rect 1409 503 1466 523
rect 1381 495 1466 503
rect 1490 519 1528 528
rect 1490 499 1499 519
rect 1519 499 1528 519
rect 1381 494 1417 495
rect 1490 491 1528 499
rect 1594 523 1679 529
rect 1699 528 1736 529
rect 1594 503 1602 523
rect 1622 522 1679 523
rect 1622 503 1651 522
rect 1594 502 1651 503
rect 1672 502 1679 522
rect 1594 495 1679 502
rect 1698 519 1736 528
rect 1698 499 1707 519
rect 1727 499 1736 519
rect 1594 494 1630 495
rect 1698 491 1736 499
rect 1802 523 1946 529
rect 1802 503 1810 523
rect 1830 503 1918 523
rect 1938 503 1946 523
rect 1802 495 1946 503
rect 1802 494 1838 495
rect 1910 494 1946 495
rect 2012 528 2049 529
rect 2012 527 2050 528
rect 2012 519 2076 527
rect 2012 499 2021 519
rect 2041 505 2076 519
rect 2096 505 2099 525
rect 2041 500 2099 505
rect 2041 499 2076 500
rect 422 469 532 483
rect 422 466 465 469
rect 111 458 236 465
rect 422 461 426 466
rect 111 439 203 458
rect 228 439 236 458
rect 111 429 236 439
rect 344 439 426 461
rect 455 439 465 466
rect 493 442 500 469
rect 529 461 532 469
rect 1278 462 1315 491
rect 529 442 594 461
rect 1279 460 1315 462
rect 1491 460 1528 491
rect 1699 464 1736 491
rect 2012 487 2076 499
rect 493 439 594 442
rect 344 437 594 439
rect 111 409 151 429
rect 110 400 151 409
rect 110 382 120 400
rect 138 382 151 400
rect 110 373 151 382
rect 110 372 147 373
rect 344 358 381 437
rect 422 424 532 437
rect 496 368 527 369
rect 344 338 353 358
rect 373 338 381 358
rect 344 328 381 338
rect 440 358 527 368
rect 440 338 449 358
rect 469 338 527 358
rect 440 329 527 338
rect 440 328 477 329
rect 113 306 150 310
rect 110 301 150 306
rect 110 283 122 301
rect 140 283 150 301
rect 110 103 150 283
rect 496 276 527 329
rect 557 358 594 437
rect 765 434 1158 454
rect 1178 434 1181 454
rect 1279 438 1528 460
rect 1697 459 1738 464
rect 2116 461 2143 639
rect 2794 551 2821 729
rect 3199 726 3240 731
rect 3409 730 3658 752
rect 3756 736 3759 756
rect 3779 736 4172 756
rect 4343 753 4380 832
rect 4410 861 4441 914
rect 4787 907 4827 1087
rect 4787 889 4797 907
rect 4815 889 4827 907
rect 4787 884 4827 889
rect 4787 880 4824 884
rect 4460 861 4497 862
rect 4410 852 4497 861
rect 4410 832 4468 852
rect 4488 832 4497 852
rect 4410 822 4497 832
rect 4556 852 4593 862
rect 4556 832 4564 852
rect 4584 832 4593 852
rect 4410 821 4441 822
rect 4405 753 4515 766
rect 4556 753 4593 832
rect 4790 817 4827 818
rect 4786 808 4827 817
rect 4786 790 4799 808
rect 4817 790 4827 808
rect 4786 781 4827 790
rect 4786 761 4826 781
rect 4343 751 4593 753
rect 4343 748 4444 751
rect 2861 691 2925 703
rect 3201 699 3238 726
rect 3409 699 3446 730
rect 3622 728 3658 730
rect 4343 729 4408 748
rect 3622 699 3659 728
rect 4405 721 4408 729
rect 4437 721 4444 748
rect 4472 724 4482 751
rect 4511 729 4593 751
rect 4701 751 4826 761
rect 4701 732 4709 751
rect 4734 732 4826 751
rect 4511 724 4515 729
rect 4701 725 4826 732
rect 4472 721 4515 724
rect 4405 707 4515 721
rect 2861 690 2896 691
rect 2838 685 2896 690
rect 2838 665 2841 685
rect 2861 671 2896 685
rect 2916 671 2925 691
rect 2861 663 2925 671
rect 2887 662 2925 663
rect 2888 661 2925 662
rect 2991 695 3027 696
rect 3099 695 3135 696
rect 2991 687 3135 695
rect 2991 667 2999 687
rect 3019 684 3107 687
rect 3019 667 3051 684
rect 3071 667 3107 684
rect 3127 667 3135 687
rect 2991 661 3135 667
rect 3201 691 3239 699
rect 3307 695 3343 696
rect 3201 671 3210 691
rect 3230 671 3239 691
rect 3201 662 3239 671
rect 3258 688 3343 695
rect 3258 668 3265 688
rect 3286 687 3343 688
rect 3286 668 3315 687
rect 3258 667 3315 668
rect 3335 667 3343 687
rect 3201 661 3238 662
rect 3258 661 3343 667
rect 3409 691 3447 699
rect 3520 695 3556 696
rect 3409 671 3418 691
rect 3438 671 3447 691
rect 3409 662 3447 671
rect 3471 687 3556 695
rect 3471 667 3528 687
rect 3548 667 3556 687
rect 3409 661 3446 662
rect 3471 661 3556 667
rect 3622 691 3660 699
rect 3622 671 3631 691
rect 3651 671 3660 691
rect 3622 662 3660 671
rect 4786 677 4826 725
rect 3622 661 3659 662
rect 3045 640 3081 661
rect 3471 640 3502 661
rect 4786 659 4797 677
rect 4815 659 4826 677
rect 4786 651 4826 659
rect 4787 650 4824 651
rect 2878 636 2978 640
rect 2878 632 2940 636
rect 2878 606 2885 632
rect 2911 610 2940 632
rect 2966 610 2978 636
rect 2911 606 2978 610
rect 2878 603 2978 606
rect 3046 603 3081 640
rect 3143 637 3502 640
rect 3143 632 3365 637
rect 3143 608 3156 632
rect 3180 613 3365 632
rect 3389 613 3502 637
rect 3180 608 3502 613
rect 3143 604 3502 608
rect 3569 632 3718 640
rect 3569 612 3580 632
rect 3600 612 3718 632
rect 3569 605 3718 612
rect 4158 609 4672 610
rect 3569 604 3610 605
rect 2893 551 2930 552
rect 2989 551 3026 552
rect 3045 551 3081 603
rect 3100 551 3137 552
rect 2793 542 2931 551
rect 2793 522 2902 542
rect 2922 522 2931 542
rect 2793 515 2931 522
rect 2989 542 3137 551
rect 2989 522 2998 542
rect 3018 522 3108 542
rect 3128 522 3137 542
rect 2793 513 2889 515
rect 2989 512 3137 522
rect 3196 542 3233 552
rect 3308 551 3345 552
rect 3289 549 3345 551
rect 3196 522 3204 542
rect 3224 522 3233 542
rect 3045 511 3081 512
rect 1975 459 2143 461
rect 1697 453 2143 459
rect 765 429 1181 434
rect 1360 432 1471 438
rect 765 428 1106 429
rect 709 368 740 369
rect 557 338 566 358
rect 586 338 594 358
rect 557 328 594 338
rect 653 361 740 368
rect 653 358 714 361
rect 653 338 662 358
rect 682 341 714 358
rect 735 341 740 361
rect 682 338 740 341
rect 653 331 740 338
rect 765 358 802 428
rect 1068 427 1105 428
rect 1360 424 1401 432
rect 1360 404 1368 424
rect 1387 404 1401 424
rect 1360 402 1401 404
rect 1429 424 1471 432
rect 1429 404 1445 424
rect 1464 404 1471 424
rect 1697 431 1703 453
rect 1729 433 2143 453
rect 2893 452 2930 453
rect 3196 452 3233 522
rect 3258 542 3345 549
rect 3258 539 3316 542
rect 3258 519 3263 539
rect 3284 522 3316 539
rect 3336 522 3345 542
rect 3284 519 3345 522
rect 3258 512 3345 519
rect 3404 542 3441 552
rect 3404 522 3412 542
rect 3432 522 3441 542
rect 3258 511 3289 512
rect 2892 451 3233 452
rect 1729 431 1738 433
rect 1975 432 2143 433
rect 2817 446 3233 451
rect 1697 422 1738 431
rect 2817 426 2820 446
rect 2840 426 3233 446
rect 3404 443 3441 522
rect 3471 551 3502 604
rect 4139 593 4672 609
rect 4139 582 4671 593
rect 4790 584 4827 588
rect 3521 551 3558 552
rect 3471 542 3558 551
rect 3471 522 3529 542
rect 3549 522 3558 542
rect 3471 512 3558 522
rect 3617 542 3654 552
rect 3617 522 3625 542
rect 3645 522 3654 542
rect 3471 511 3502 512
rect 3466 443 3576 456
rect 3617 443 3654 522
rect 3404 441 3654 443
rect 3404 438 3505 441
rect 3404 419 3469 438
rect 1429 402 1471 404
rect 1360 387 1471 402
rect 3466 411 3469 419
rect 3498 411 3505 438
rect 3533 414 3543 441
rect 3572 419 3654 441
rect 3732 513 3900 514
rect 4139 513 4177 582
rect 3732 493 4177 513
rect 4404 544 4515 559
rect 4404 542 4446 544
rect 4404 522 4411 542
rect 4430 522 4446 542
rect 4404 514 4446 522
rect 4474 542 4515 544
rect 4474 522 4488 542
rect 4507 522 4515 542
rect 4474 514 4515 522
rect 4404 508 4515 514
rect 4637 519 4671 582
rect 4789 578 4827 584
rect 4789 560 4799 578
rect 4817 560 4827 578
rect 4789 551 4827 560
rect 4789 519 4823 551
rect 3732 487 4176 493
rect 3732 485 3900 487
rect 3572 414 3576 419
rect 3533 411 3576 414
rect 3466 397 3576 411
rect 917 368 953 369
rect 765 338 774 358
rect 794 338 802 358
rect 653 329 709 331
rect 653 328 690 329
rect 765 328 802 338
rect 861 358 1009 368
rect 1109 365 1205 367
rect 861 338 870 358
rect 890 338 980 358
rect 1000 338 1009 358
rect 861 329 1009 338
rect 1067 358 1205 365
rect 1067 338 1076 358
rect 1096 338 1205 358
rect 1067 329 1205 338
rect 861 328 898 329
rect 917 277 953 329
rect 972 328 1009 329
rect 1068 328 1105 329
rect 388 275 429 276
rect 280 268 429 275
rect 280 248 398 268
rect 418 248 429 268
rect 280 240 429 248
rect 496 272 855 276
rect 496 267 818 272
rect 496 243 609 267
rect 633 248 818 267
rect 842 248 855 272
rect 633 243 855 248
rect 496 240 855 243
rect 917 240 952 277
rect 1020 274 1120 277
rect 1020 270 1087 274
rect 1020 244 1032 270
rect 1058 248 1087 270
rect 1113 248 1120 274
rect 1058 244 1120 248
rect 1020 240 1120 244
rect 496 219 527 240
rect 917 219 953 240
rect 339 218 376 219
rect 338 209 376 218
rect 338 189 347 209
rect 367 189 376 209
rect 338 181 376 189
rect 442 213 527 219
rect 552 218 589 219
rect 442 193 450 213
rect 470 193 527 213
rect 442 185 527 193
rect 551 209 589 218
rect 551 189 560 209
rect 580 189 589 209
rect 442 184 478 185
rect 551 181 589 189
rect 655 213 740 219
rect 760 218 797 219
rect 655 193 663 213
rect 683 212 740 213
rect 683 193 712 212
rect 655 192 712 193
rect 733 192 740 212
rect 655 185 740 192
rect 759 209 797 218
rect 759 189 768 209
rect 788 189 797 209
rect 655 184 691 185
rect 759 181 797 189
rect 863 213 1007 219
rect 863 193 871 213
rect 891 210 979 213
rect 891 193 922 210
rect 863 190 922 193
rect 945 193 979 210
rect 999 193 1007 213
rect 945 190 1007 193
rect 863 185 1007 190
rect 863 184 899 185
rect 971 184 1007 185
rect 1073 218 1110 219
rect 1073 217 1111 218
rect 1073 209 1137 217
rect 1073 189 1082 209
rect 1102 195 1137 209
rect 1157 195 1160 215
rect 1102 190 1160 195
rect 1102 189 1137 190
rect 339 152 376 181
rect 340 150 376 152
rect 552 150 589 181
rect 340 128 589 150
rect 760 149 797 181
rect 1073 177 1137 189
rect 1177 151 1204 329
rect 3732 307 3759 485
rect 3799 447 3863 459
rect 4139 455 4176 487
rect 4347 486 4596 508
rect 4637 487 4823 519
rect 4651 486 4823 487
rect 4347 455 4384 486
rect 4560 484 4596 486
rect 4560 455 4597 484
rect 4789 458 4823 486
rect 3799 446 3834 447
rect 3776 441 3834 446
rect 3776 421 3779 441
rect 3799 427 3834 441
rect 3854 427 3863 447
rect 3799 419 3863 427
rect 3825 418 3863 419
rect 3826 417 3863 418
rect 3929 451 3965 452
rect 4037 451 4073 452
rect 3929 444 4073 451
rect 3929 443 3989 444
rect 3929 423 3937 443
rect 3957 424 3989 443
rect 4014 443 4073 444
rect 4014 424 4045 443
rect 3957 423 4045 424
rect 4065 423 4073 443
rect 3929 417 4073 423
rect 4139 447 4177 455
rect 4245 451 4281 452
rect 4139 427 4148 447
rect 4168 427 4177 447
rect 4139 418 4177 427
rect 4196 444 4281 451
rect 4196 424 4203 444
rect 4224 443 4281 444
rect 4224 424 4253 443
rect 4196 423 4253 424
rect 4273 423 4281 443
rect 4139 417 4176 418
rect 4196 417 4281 423
rect 4347 447 4385 455
rect 4458 451 4494 452
rect 4347 427 4356 447
rect 4376 427 4385 447
rect 4347 418 4385 427
rect 4409 443 4494 451
rect 4409 423 4466 443
rect 4486 423 4494 443
rect 4347 417 4384 418
rect 4409 417 4494 423
rect 4560 447 4598 455
rect 4560 427 4569 447
rect 4589 427 4598 447
rect 4560 418 4598 427
rect 4787 448 4824 458
rect 4787 430 4797 448
rect 4815 430 4824 448
rect 4787 421 4824 430
rect 4789 420 4823 421
rect 4560 417 4597 418
rect 3983 396 4019 417
rect 4409 396 4440 417
rect 3816 392 3916 396
rect 3816 388 3878 392
rect 3816 362 3823 388
rect 3849 366 3878 388
rect 3904 366 3916 392
rect 3849 362 3916 366
rect 3816 359 3916 362
rect 3984 359 4019 396
rect 4081 393 4440 396
rect 4081 388 4303 393
rect 4081 364 4094 388
rect 4118 369 4303 388
rect 4327 369 4440 393
rect 4118 364 4440 369
rect 4081 360 4440 364
rect 4507 388 4656 396
rect 4507 368 4518 388
rect 4538 368 4656 388
rect 4507 361 4656 368
rect 4507 360 4548 361
rect 3831 307 3868 308
rect 3927 307 3964 308
rect 3983 307 4019 359
rect 4038 307 4075 308
rect 3731 298 3869 307
rect 3731 278 3840 298
rect 3860 278 3869 298
rect 3731 271 3869 278
rect 3927 298 4075 307
rect 3927 278 3936 298
rect 3956 278 4046 298
rect 4066 278 4075 298
rect 3731 269 3827 271
rect 3927 268 4075 278
rect 4134 298 4171 308
rect 4246 307 4283 308
rect 4227 305 4283 307
rect 4134 278 4142 298
rect 4162 278 4171 298
rect 3983 267 4019 268
rect 3831 208 3868 209
rect 4134 208 4171 278
rect 4196 298 4283 305
rect 4196 295 4254 298
rect 4196 275 4201 295
rect 4222 278 4254 295
rect 4274 278 4283 298
rect 4222 275 4283 278
rect 4196 268 4283 275
rect 4342 298 4379 308
rect 4342 278 4350 298
rect 4370 278 4379 298
rect 4196 267 4227 268
rect 3830 207 4171 208
rect 3755 202 4171 207
rect 3755 182 3758 202
rect 3778 182 4171 202
rect 4342 199 4379 278
rect 4409 307 4440 360
rect 4790 358 4827 359
rect 4789 349 4828 358
rect 4789 331 4799 349
rect 4817 331 4828 349
rect 4701 314 4748 315
rect 4789 314 4828 331
rect 4701 310 4828 314
rect 4459 307 4496 308
rect 4409 298 4496 307
rect 4409 278 4467 298
rect 4487 278 4496 298
rect 4409 268 4496 278
rect 4555 298 4592 308
rect 4555 278 4563 298
rect 4583 278 4592 298
rect 4409 267 4440 268
rect 4404 199 4514 212
rect 4555 199 4592 278
rect 4701 281 4711 310
rect 4740 281 4828 310
rect 4701 275 4828 281
rect 4701 271 4748 275
rect 4786 261 4828 275
rect 4786 243 4797 261
rect 4815 243 4828 261
rect 4786 238 4828 243
rect 4787 235 4828 238
rect 4787 234 4824 235
rect 4342 197 4592 199
rect 4342 194 4443 197
rect 4342 175 4407 194
rect 4404 167 4407 175
rect 4436 167 4443 194
rect 4471 170 4481 197
rect 4510 175 4592 197
rect 4510 170 4514 175
rect 4471 167 4514 170
rect 4404 153 4514 167
rect 4780 171 4827 172
rect 4780 162 4828 171
rect 1036 149 1204 151
rect 760 146 1204 149
rect 421 122 532 128
rect 421 114 462 122
rect 110 59 149 103
rect 421 94 429 114
rect 448 94 462 114
rect 421 92 462 94
rect 490 116 532 122
rect 758 123 1204 146
rect 4780 144 4799 162
rect 4817 144 4828 162
rect 4780 142 4828 144
rect 4789 123 4828 142
rect 490 114 531 116
rect 490 94 506 114
rect 525 94 531 114
rect 490 92 531 94
rect 421 77 531 92
rect 110 35 150 59
rect 758 49 796 123
rect 1036 122 1204 123
rect 718 35 797 49
rect 110 34 400 35
rect 566 34 797 35
rect 110 32 797 34
rect 110 11 757 32
rect 786 11 797 32
rect 110 2 797 11
rect 4787 36 4831 123
rect 4787 15 4792 36
rect 4821 15 4831 36
rect 4787 2 4831 15
rect 718 -8 797 2
rect 1669 -90 1779 -76
rect 1669 -93 1712 -90
rect 1669 -98 1673 -93
rect 1591 -120 1673 -98
rect 1702 -120 1712 -93
rect 1740 -117 1747 -90
rect 1776 -98 1779 -90
rect 1776 -117 1841 -98
rect 1740 -120 1841 -117
rect 1591 -122 1841 -120
rect 1591 -201 1628 -122
rect 1669 -135 1779 -122
rect 1743 -191 1774 -190
rect 1591 -221 1600 -201
rect 1620 -221 1628 -201
rect 1591 -231 1628 -221
rect 1687 -201 1774 -191
rect 1687 -221 1696 -201
rect 1716 -221 1774 -201
rect 1687 -230 1774 -221
rect 1687 -231 1724 -230
rect 1743 -283 1774 -230
rect 1804 -201 1841 -122
rect 2012 -125 2405 -105
rect 2425 -125 2428 -105
rect 2012 -130 2428 -125
rect 2012 -131 2353 -130
rect 1956 -191 1987 -190
rect 1804 -221 1813 -201
rect 1833 -221 1841 -201
rect 1804 -231 1841 -221
rect 1900 -198 1987 -191
rect 1900 -201 1961 -198
rect 1900 -221 1909 -201
rect 1929 -218 1961 -201
rect 1982 -218 1987 -198
rect 1929 -221 1987 -218
rect 1900 -228 1987 -221
rect 2012 -201 2049 -131
rect 2315 -132 2352 -131
rect 2164 -191 2200 -190
rect 2012 -221 2021 -201
rect 2041 -221 2049 -201
rect 1900 -230 1956 -228
rect 1900 -231 1937 -230
rect 2012 -231 2049 -221
rect 2108 -201 2256 -191
rect 2356 -194 2452 -192
rect 2108 -221 2117 -201
rect 2137 -221 2227 -201
rect 2247 -221 2256 -201
rect 2108 -230 2256 -221
rect 2314 -201 2452 -194
rect 2314 -221 2323 -201
rect 2343 -221 2452 -201
rect 2314 -230 2452 -221
rect 2108 -231 2145 -230
rect 2164 -282 2200 -230
rect 2219 -231 2256 -230
rect 2315 -231 2352 -230
rect 1635 -284 1676 -283
rect 1527 -291 1676 -284
rect 1527 -311 1645 -291
rect 1665 -311 1676 -291
rect 1527 -319 1676 -311
rect 1743 -287 2102 -283
rect 1743 -292 2065 -287
rect 1743 -316 1856 -292
rect 1880 -311 2065 -292
rect 2089 -311 2102 -287
rect 1880 -316 2102 -311
rect 1743 -319 2102 -316
rect 2164 -319 2199 -282
rect 2267 -285 2367 -282
rect 2267 -289 2334 -285
rect 2267 -315 2279 -289
rect 2305 -311 2334 -289
rect 2360 -311 2367 -285
rect 2305 -315 2367 -311
rect 2267 -319 2367 -315
rect 1743 -340 1774 -319
rect 2164 -340 2200 -319
rect 1586 -341 1623 -340
rect 1585 -350 1623 -341
rect 1585 -370 1594 -350
rect 1614 -370 1623 -350
rect 1585 -378 1623 -370
rect 1689 -346 1774 -340
rect 1799 -341 1836 -340
rect 1689 -366 1697 -346
rect 1717 -366 1774 -346
rect 1689 -374 1774 -366
rect 1798 -350 1836 -341
rect 1798 -370 1807 -350
rect 1827 -370 1836 -350
rect 1689 -375 1725 -374
rect 1798 -378 1836 -370
rect 1902 -346 1987 -340
rect 2007 -341 2044 -340
rect 1902 -366 1910 -346
rect 1930 -347 1987 -346
rect 1930 -366 1959 -347
rect 1902 -367 1959 -366
rect 1980 -367 1987 -347
rect 1902 -374 1987 -367
rect 2006 -350 2044 -341
rect 2006 -370 2015 -350
rect 2035 -370 2044 -350
rect 1902 -375 1938 -374
rect 2006 -378 2044 -370
rect 2110 -346 2254 -340
rect 2110 -366 2118 -346
rect 2138 -348 2226 -346
rect 2138 -366 2165 -348
rect 2110 -368 2165 -366
rect 2199 -366 2226 -348
rect 2246 -366 2254 -346
rect 2199 -368 2254 -366
rect 2110 -374 2254 -368
rect 2110 -375 2146 -374
rect 2218 -375 2254 -374
rect 2320 -341 2357 -340
rect 2320 -342 2358 -341
rect 2320 -350 2384 -342
rect 2320 -370 2329 -350
rect 2349 -364 2384 -350
rect 2404 -364 2407 -344
rect 2349 -369 2407 -364
rect 2349 -370 2384 -369
rect 1586 -407 1623 -378
rect 1587 -409 1623 -407
rect 1799 -409 1836 -378
rect 1587 -431 1836 -409
rect 2007 -410 2044 -378
rect 2320 -382 2384 -370
rect 2424 -399 2451 -230
rect 2397 -405 2525 -399
rect 2397 -408 2486 -405
rect 2283 -410 2486 -408
rect 2007 -426 2486 -410
rect 2513 -426 2525 -405
rect 1668 -437 1779 -431
rect 2007 -436 2525 -426
rect 2283 -437 2525 -436
rect 1668 -445 1709 -437
rect 1668 -465 1676 -445
rect 1695 -465 1709 -445
rect 1668 -467 1709 -465
rect 1737 -445 1779 -437
rect 2397 -439 2525 -437
rect 1737 -465 1753 -445
rect 1772 -465 1779 -445
rect 1737 -467 1779 -465
rect 1668 -482 1779 -467
<< viali >>
rect 4408 8797 4427 8817
rect 4485 8797 4504 8817
rect 423 8714 452 8741
rect 497 8717 526 8744
rect 193 8601 222 8630
rect 1155 8709 1175 8729
rect 711 8616 732 8636
rect 1084 8523 1110 8549
rect 709 8467 730 8487
rect 919 8467 944 8487
rect 1134 8470 1154 8490
rect 3776 8696 3796 8716
rect 3988 8701 4011 8721
rect 4200 8699 4221 8719
rect 3820 8637 3846 8663
rect 426 8369 445 8389
rect 503 8369 522 8389
rect 1361 8470 1390 8497
rect 1435 8473 1464 8500
rect 2093 8465 2113 8485
rect 1649 8372 1670 8392
rect 3204 8458 3230 8480
rect 3469 8487 3488 8507
rect 3546 8487 3565 8507
rect 4198 8550 4219 8570
rect 2022 8279 2048 8305
rect 1647 8223 1668 8243
rect 1862 8227 1882 8244
rect 2072 8226 2092 8246
rect 199 8160 224 8179
rect 422 8160 451 8187
rect 496 8163 525 8190
rect 1154 8155 1174 8175
rect 3755 8457 3775 8477
rect 4404 8442 4433 8469
rect 4478 8445 4507 8472
rect 4705 8453 4730 8472
rect 2837 8386 2857 8406
rect 3261 8389 3282 8409
rect 2881 8327 2907 8353
rect 3048 8248 3069 8289
rect 710 8062 731 8082
rect 1364 8125 1383 8145
rect 1441 8125 1460 8145
rect 1699 8152 1725 8174
rect 3259 8240 3280 8260
rect 2816 8147 2836 8167
rect 3189 8154 3221 8171
rect 3465 8132 3494 8159
rect 3539 8135 3568 8162
rect 4407 8243 4426 8263
rect 4484 8243 4503 8263
rect 1083 7969 1109 7995
rect 708 7913 729 7933
rect 918 7911 941 7931
rect 1133 7916 1153 7936
rect 3775 8142 3795 8162
rect 3985 8145 4010 8165
rect 4199 8145 4220 8165
rect 3819 8083 3845 8109
rect 3041 7948 3072 7975
rect 3329 7976 3348 7996
rect 3406 7976 3425 7996
rect 425 7815 444 7835
rect 502 7815 521 7835
rect 1502 7878 1531 7905
rect 1576 7881 1605 7908
rect 1860 7872 1880 7889
rect 2234 7873 2254 7893
rect 1790 7780 1811 7800
rect 2163 7687 2189 7713
rect 424 7611 453 7638
rect 498 7614 527 7641
rect 194 7498 223 7527
rect 1156 7606 1176 7626
rect 1788 7631 1809 7651
rect 1996 7629 2023 7650
rect 2213 7634 2233 7654
rect 712 7513 733 7533
rect 4197 7996 4218 8016
rect 2697 7875 2717 7895
rect 3121 7878 3142 7898
rect 3754 7903 3774 7923
rect 4707 8002 4736 8031
rect 4403 7888 4432 7915
rect 4477 7891 4506 7918
rect 2741 7816 2767 7842
rect 2908 7736 2931 7774
rect 3119 7729 3140 7749
rect 2676 7636 2696 7656
rect 3050 7640 3070 7657
rect 3325 7621 3354 7648
rect 3399 7624 3428 7651
rect 4409 7694 4428 7714
rect 4486 7694 4505 7714
rect 1505 7533 1524 7553
rect 1582 7533 1601 7553
rect 1858 7554 1889 7581
rect 1085 7420 1111 7446
rect 710 7364 731 7384
rect 920 7364 945 7384
rect 1135 7367 1155 7387
rect 3777 7593 3797 7613
rect 3989 7598 4012 7618
rect 4201 7596 4222 7616
rect 3821 7534 3847 7560
rect 427 7266 446 7286
rect 504 7266 523 7286
rect 1362 7367 1391 7394
rect 1436 7370 1465 7397
rect 1709 7358 1741 7375
rect 2094 7362 2114 7382
rect 1650 7269 1671 7289
rect 3205 7355 3231 7377
rect 3470 7384 3489 7404
rect 3547 7384 3566 7404
rect 4199 7447 4220 7467
rect 1861 7240 1882 7281
rect 2023 7176 2049 7202
rect 1648 7120 1669 7140
rect 2073 7123 2093 7143
rect 200 7057 225 7076
rect 423 7057 452 7084
rect 497 7060 526 7087
rect 1155 7052 1175 7072
rect 3756 7354 3776 7374
rect 4405 7339 4434 7366
rect 4479 7342 4508 7369
rect 4706 7350 4731 7369
rect 2838 7283 2858 7303
rect 3048 7285 3068 7302
rect 3262 7286 3283 7306
rect 2882 7224 2908 7250
rect 711 6959 732 6979
rect 1365 7022 1384 7042
rect 1442 7022 1461 7042
rect 1700 7049 1726 7071
rect 3260 7137 3281 7157
rect 2817 7044 2837 7064
rect 3466 7029 3495 7056
rect 3540 7032 3569 7059
rect 4408 7140 4427 7160
rect 4485 7140 4504 7160
rect 1084 6866 1110 6892
rect 709 6810 730 6830
rect 919 6808 942 6828
rect 1134 6813 1154 6833
rect 3776 7039 3796 7059
rect 3986 7042 4011 7062
rect 4200 7042 4221 7062
rect 3820 6980 3846 7006
rect 2707 6832 2755 6861
rect 3360 6860 3379 6880
rect 3437 6860 3456 6880
rect 426 6712 445 6732
rect 503 6712 522 6732
rect 1472 6788 1501 6815
rect 1546 6791 1575 6818
rect 2204 6783 2224 6803
rect 1760 6690 1781 6710
rect 2133 6597 2159 6623
rect 424 6508 453 6535
rect 498 6511 527 6538
rect 1758 6541 1779 6561
rect 1966 6541 1995 6560
rect 2183 6544 2203 6564
rect 194 6395 223 6424
rect 1156 6503 1176 6523
rect 712 6410 733 6430
rect 4198 6893 4219 6913
rect 3755 6800 3775 6820
rect 4708 6899 4737 6928
rect 2728 6759 2748 6779
rect 3152 6762 3173 6782
rect 4404 6785 4433 6812
rect 4478 6788 4507 6815
rect 2772 6700 2798 6726
rect 2937 6625 2964 6657
rect 3150 6613 3171 6633
rect 2707 6522 2727 6540
rect 3097 6518 3118 6538
rect 3356 6505 3385 6532
rect 3430 6508 3459 6535
rect 4409 6591 4428 6611
rect 4486 6591 4505 6611
rect 1475 6443 1494 6463
rect 1552 6443 1571 6463
rect 1085 6317 1111 6343
rect 710 6261 731 6281
rect 920 6261 945 6281
rect 1135 6264 1155 6284
rect 3777 6490 3797 6510
rect 3989 6495 4012 6515
rect 4201 6493 4222 6513
rect 3821 6431 3847 6457
rect 2176 6322 2224 6351
rect 427 6163 446 6183
rect 504 6163 523 6183
rect 1362 6264 1391 6291
rect 1436 6267 1465 6294
rect 2094 6259 2114 6279
rect 1650 6166 1671 6186
rect 3205 6252 3231 6274
rect 3470 6281 3489 6301
rect 3547 6281 3566 6301
rect 4199 6344 4220 6364
rect 2023 6073 2049 6099
rect 1648 6017 1669 6037
rect 1863 6021 1883 6038
rect 2073 6020 2093 6040
rect 200 5954 225 5973
rect 423 5954 452 5981
rect 497 5957 526 5984
rect 1155 5949 1175 5969
rect 3756 6251 3776 6271
rect 4405 6236 4434 6263
rect 4479 6239 4508 6266
rect 4706 6247 4731 6266
rect 2838 6180 2858 6200
rect 3262 6183 3283 6203
rect 2882 6121 2908 6147
rect 3049 6042 3070 6083
rect 711 5856 732 5876
rect 1365 5919 1384 5939
rect 1442 5919 1461 5939
rect 1700 5946 1726 5968
rect 3260 6034 3281 6054
rect 2817 5941 2837 5961
rect 3190 5948 3222 5965
rect 3466 5926 3495 5953
rect 3540 5929 3569 5956
rect 4408 6037 4427 6057
rect 4485 6037 4504 6057
rect 1084 5763 1110 5789
rect 709 5707 730 5727
rect 919 5705 942 5725
rect 1134 5710 1154 5730
rect 3776 5936 3796 5956
rect 3986 5939 4011 5959
rect 4200 5939 4221 5959
rect 3820 5877 3846 5903
rect 3042 5742 3073 5769
rect 3330 5770 3349 5790
rect 3407 5770 3426 5790
rect 426 5609 445 5629
rect 503 5609 522 5629
rect 1503 5672 1532 5699
rect 1577 5675 1606 5702
rect 1861 5666 1881 5683
rect 2235 5667 2255 5687
rect 1791 5574 1812 5594
rect 2000 5549 2023 5587
rect 2164 5481 2190 5507
rect 425 5405 454 5432
rect 499 5408 528 5435
rect 195 5292 224 5321
rect 1157 5400 1177 5420
rect 1789 5425 1810 5445
rect 2214 5428 2234 5448
rect 713 5307 734 5327
rect 4198 5790 4219 5810
rect 2698 5669 2718 5689
rect 2908 5673 2935 5694
rect 3122 5672 3143 5692
rect 3755 5697 3775 5717
rect 4708 5796 4737 5825
rect 4404 5682 4433 5709
rect 4478 5685 4507 5712
rect 2742 5610 2768 5636
rect 3120 5523 3141 5543
rect 2677 5430 2697 5450
rect 3051 5434 3071 5451
rect 3326 5415 3355 5442
rect 3400 5418 3429 5445
rect 4410 5488 4429 5508
rect 4487 5488 4506 5508
rect 1506 5327 1525 5347
rect 1583 5327 1602 5347
rect 1859 5348 1890 5375
rect 1086 5214 1112 5240
rect 711 5158 732 5178
rect 921 5158 946 5178
rect 1136 5161 1156 5181
rect 3778 5387 3798 5407
rect 3990 5392 4013 5412
rect 4202 5390 4223 5410
rect 3822 5328 3848 5354
rect 428 5060 447 5080
rect 505 5060 524 5080
rect 1363 5161 1392 5188
rect 1437 5164 1466 5191
rect 1710 5152 1742 5169
rect 2095 5156 2115 5176
rect 1651 5063 1672 5083
rect 3206 5149 3232 5171
rect 3471 5178 3490 5198
rect 3548 5178 3567 5198
rect 4200 5241 4221 5261
rect 1862 5034 1883 5075
rect 2024 4970 2050 4996
rect 1649 4914 1670 4934
rect 2074 4917 2094 4937
rect 201 4851 226 4870
rect 424 4851 453 4878
rect 498 4854 527 4881
rect 1156 4846 1176 4866
rect 3757 5148 3777 5168
rect 4406 5133 4435 5160
rect 4480 5136 4509 5163
rect 4707 5144 4732 5163
rect 2839 5077 2859 5097
rect 3049 5079 3069 5096
rect 3263 5080 3284 5100
rect 2883 5018 2909 5044
rect 712 4753 733 4773
rect 1366 4816 1385 4836
rect 1443 4816 1462 4836
rect 1701 4843 1727 4865
rect 3261 4931 3282 4951
rect 2818 4838 2838 4858
rect 3467 4823 3496 4850
rect 3541 4826 3570 4853
rect 4409 4934 4428 4954
rect 4486 4934 4505 4954
rect 2567 4765 2594 4805
rect 1085 4660 1111 4686
rect 710 4604 731 4624
rect 920 4602 943 4622
rect 1135 4607 1155 4627
rect 3777 4833 3797 4853
rect 3987 4836 4012 4856
rect 4201 4836 4222 4856
rect 3821 4774 3847 4800
rect 3362 4648 3381 4668
rect 3439 4648 3458 4668
rect 427 4506 446 4526
rect 504 4506 523 4526
rect 1472 4588 1501 4615
rect 1546 4591 1575 4618
rect 2204 4583 2224 4603
rect 1760 4490 1781 4510
rect 2133 4397 2159 4423
rect 425 4302 454 4329
rect 499 4305 528 4332
rect 1758 4341 1779 4361
rect 1966 4340 1992 4364
rect 2183 4344 2203 4364
rect 195 4189 224 4218
rect 1157 4297 1177 4317
rect 713 4204 734 4224
rect 4199 4687 4220 4707
rect 3756 4594 3776 4614
rect 4709 4693 4738 4722
rect 2730 4547 2750 4567
rect 2937 4550 2962 4570
rect 3154 4550 3175 4570
rect 4405 4579 4434 4606
rect 4479 4582 4508 4609
rect 2774 4488 2800 4514
rect 3152 4401 3173 4421
rect 2709 4308 2729 4328
rect 3358 4293 3387 4320
rect 3432 4296 3461 4323
rect 4410 4385 4429 4405
rect 4487 4385 4506 4405
rect 1475 4243 1494 4263
rect 1552 4243 1571 4263
rect 1086 4111 1112 4137
rect 711 4055 732 4075
rect 921 4055 946 4075
rect 1136 4058 1156 4078
rect 3778 4284 3798 4304
rect 3990 4289 4013 4309
rect 4202 4287 4223 4307
rect 3822 4225 3848 4251
rect 2339 4106 2366 4146
rect 428 3957 447 3977
rect 505 3957 524 3977
rect 1363 4058 1392 4085
rect 1437 4061 1466 4088
rect 2095 4053 2115 4073
rect 1651 3960 1672 3980
rect 3206 4046 3232 4068
rect 3471 4075 3490 4095
rect 3548 4075 3567 4095
rect 4200 4138 4221 4158
rect 2024 3867 2050 3893
rect 1649 3811 1670 3831
rect 1864 3815 1884 3832
rect 2074 3814 2094 3834
rect 201 3748 226 3767
rect 424 3748 453 3775
rect 498 3751 527 3778
rect 1156 3743 1176 3763
rect 3757 4045 3777 4065
rect 4406 4030 4435 4057
rect 4480 4033 4509 4060
rect 4707 4041 4732 4060
rect 2839 3974 2859 3994
rect 3263 3977 3284 3997
rect 2883 3915 2909 3941
rect 3050 3836 3071 3877
rect 712 3650 733 3670
rect 1366 3713 1385 3733
rect 1443 3713 1462 3733
rect 1701 3740 1727 3762
rect 3261 3828 3282 3848
rect 2818 3735 2838 3755
rect 3191 3742 3223 3759
rect 3467 3720 3496 3747
rect 3541 3723 3570 3750
rect 4409 3831 4428 3851
rect 4486 3831 4505 3851
rect 1085 3557 1111 3583
rect 710 3501 731 3521
rect 920 3499 943 3519
rect 1135 3504 1155 3524
rect 3777 3730 3797 3750
rect 3987 3733 4012 3753
rect 4201 3733 4222 3753
rect 3821 3671 3847 3697
rect 3043 3536 3074 3563
rect 3331 3564 3350 3584
rect 3408 3564 3427 3584
rect 427 3403 446 3423
rect 504 3403 523 3423
rect 1504 3466 1533 3493
rect 1578 3469 1607 3496
rect 1862 3460 1882 3477
rect 2236 3461 2256 3481
rect 1792 3368 1813 3388
rect 2165 3275 2191 3301
rect 426 3199 455 3226
rect 500 3202 529 3229
rect 196 3086 225 3115
rect 1158 3194 1178 3214
rect 1790 3219 1811 3239
rect 1998 3217 2025 3238
rect 2215 3222 2235 3242
rect 714 3101 735 3121
rect 4199 3584 4220 3604
rect 2699 3463 2719 3483
rect 3123 3466 3144 3486
rect 3756 3491 3776 3511
rect 4709 3590 4738 3619
rect 4405 3476 4434 3503
rect 4479 3479 4508 3506
rect 2743 3404 2769 3430
rect 2910 3324 2933 3362
rect 3121 3317 3142 3337
rect 2678 3224 2698 3244
rect 3052 3228 3072 3245
rect 3327 3209 3356 3236
rect 3401 3212 3430 3239
rect 4411 3282 4430 3302
rect 4488 3282 4507 3302
rect 1507 3121 1526 3141
rect 1584 3121 1603 3141
rect 1860 3142 1891 3169
rect 1087 3008 1113 3034
rect 712 2952 733 2972
rect 922 2952 947 2972
rect 1137 2955 1157 2975
rect 3779 3181 3799 3201
rect 3991 3186 4014 3206
rect 4203 3184 4224 3204
rect 3823 3122 3849 3148
rect 429 2854 448 2874
rect 506 2854 525 2874
rect 1364 2955 1393 2982
rect 1438 2958 1467 2985
rect 1711 2946 1743 2963
rect 2096 2950 2116 2970
rect 1652 2857 1673 2877
rect 3207 2943 3233 2965
rect 3472 2972 3491 2992
rect 3549 2972 3568 2992
rect 4201 3035 4222 3055
rect 1863 2828 1884 2869
rect 2025 2764 2051 2790
rect 1650 2708 1671 2728
rect 2075 2711 2095 2731
rect 202 2645 227 2664
rect 425 2645 454 2672
rect 499 2648 528 2675
rect 1157 2640 1177 2660
rect 3758 2942 3778 2962
rect 4407 2927 4436 2954
rect 4481 2930 4510 2957
rect 4708 2938 4733 2957
rect 2840 2871 2860 2891
rect 3050 2873 3070 2890
rect 3264 2874 3285 2894
rect 2884 2812 2910 2838
rect 713 2547 734 2567
rect 1367 2610 1386 2630
rect 1444 2610 1463 2630
rect 1702 2637 1728 2659
rect 3262 2725 3283 2745
rect 2819 2632 2839 2652
rect 3468 2617 3497 2644
rect 3542 2620 3571 2647
rect 4410 2728 4429 2748
rect 4487 2728 4506 2748
rect 2709 2560 2757 2589
rect 1086 2454 1112 2480
rect 711 2398 732 2418
rect 921 2396 944 2416
rect 1136 2401 1156 2421
rect 3778 2627 3798 2647
rect 3988 2630 4013 2650
rect 4202 2630 4223 2650
rect 3822 2568 3848 2594
rect 3362 2448 3381 2468
rect 3439 2448 3458 2468
rect 428 2300 447 2320
rect 505 2300 524 2320
rect 1474 2376 1503 2403
rect 1548 2379 1577 2406
rect 1815 2373 1836 2393
rect 2206 2371 2226 2389
rect 1762 2278 1783 2298
rect 1969 2254 1996 2286
rect 2135 2185 2161 2211
rect 426 2096 455 2123
rect 500 2099 529 2126
rect 1760 2129 1781 2149
rect 2185 2132 2205 2152
rect 196 1983 225 2012
rect 1158 2091 1178 2111
rect 714 1998 735 2018
rect 4200 2481 4221 2501
rect 3757 2388 3777 2408
rect 4710 2487 4739 2516
rect 2730 2347 2750 2367
rect 2938 2351 2967 2370
rect 3154 2350 3175 2370
rect 4406 2373 4435 2400
rect 4480 2376 4509 2403
rect 2774 2288 2800 2314
rect 3152 2201 3173 2221
rect 2709 2108 2729 2128
rect 3358 2093 3387 2120
rect 3432 2096 3461 2123
rect 4411 2179 4430 2199
rect 4488 2179 4507 2199
rect 1477 2031 1496 2051
rect 1554 2031 1573 2051
rect 2178 2050 2226 2079
rect 1087 1905 1113 1931
rect 712 1849 733 1869
rect 922 1849 947 1869
rect 1137 1852 1157 1872
rect 3779 2078 3799 2098
rect 3991 2083 4014 2103
rect 4203 2081 4224 2101
rect 3823 2019 3849 2045
rect 429 1751 448 1771
rect 506 1751 525 1771
rect 1364 1852 1393 1879
rect 1438 1855 1467 1882
rect 2096 1847 2116 1867
rect 1652 1754 1673 1774
rect 3207 1840 3233 1862
rect 3472 1869 3491 1889
rect 3549 1869 3568 1889
rect 4201 1932 4222 1952
rect 2025 1661 2051 1687
rect 1650 1605 1671 1625
rect 1865 1609 1885 1626
rect 2075 1608 2095 1628
rect 202 1542 227 1561
rect 425 1542 454 1569
rect 499 1545 528 1572
rect 1157 1537 1177 1557
rect 3758 1839 3778 1859
rect 4407 1824 4436 1851
rect 4481 1827 4510 1854
rect 4708 1835 4733 1854
rect 2840 1768 2860 1788
rect 3264 1771 3285 1791
rect 2884 1709 2910 1735
rect 3051 1630 3072 1671
rect 713 1444 734 1464
rect 1367 1507 1386 1527
rect 1444 1507 1463 1527
rect 1702 1534 1728 1556
rect 3262 1622 3283 1642
rect 2819 1529 2839 1549
rect 3192 1536 3224 1553
rect 3468 1514 3497 1541
rect 3542 1517 3571 1544
rect 4410 1625 4429 1645
rect 4487 1625 4506 1645
rect 1086 1351 1112 1377
rect 711 1295 732 1315
rect 921 1293 944 1313
rect 1136 1298 1156 1318
rect 3778 1524 3798 1544
rect 3988 1527 4013 1547
rect 4202 1527 4223 1547
rect 3822 1465 3848 1491
rect 3044 1330 3075 1357
rect 3332 1358 3351 1378
rect 3409 1358 3428 1378
rect 428 1197 447 1217
rect 505 1197 524 1217
rect 1505 1260 1534 1287
rect 1579 1263 1608 1290
rect 1863 1254 1883 1271
rect 2237 1255 2257 1275
rect 1793 1162 1814 1182
rect 2002 1137 2025 1175
rect 2166 1069 2192 1095
rect 427 993 456 1020
rect 501 996 530 1023
rect 197 880 226 909
rect 1159 988 1179 1008
rect 1791 1013 1812 1033
rect 2216 1016 2236 1036
rect 715 895 736 915
rect 4200 1378 4221 1398
rect 2700 1257 2720 1277
rect 2910 1261 2937 1282
rect 3124 1260 3145 1280
rect 3757 1285 3777 1305
rect 4710 1384 4739 1413
rect 4406 1270 4435 1297
rect 4480 1273 4509 1300
rect 2744 1198 2770 1224
rect 3122 1111 3143 1131
rect 2679 1018 2699 1038
rect 3053 1022 3073 1039
rect 3328 1003 3357 1030
rect 3402 1006 3431 1033
rect 4412 1076 4431 1096
rect 4489 1076 4508 1096
rect 1508 915 1527 935
rect 1585 915 1604 935
rect 1861 936 1892 963
rect 1088 802 1114 828
rect 713 746 734 766
rect 923 746 948 766
rect 1138 749 1158 769
rect 3780 975 3800 995
rect 3992 980 4015 1000
rect 4204 978 4225 998
rect 3824 916 3850 942
rect 430 648 449 668
rect 507 648 526 668
rect 1365 749 1394 776
rect 1439 752 1468 779
rect 1712 740 1744 757
rect 2097 744 2117 764
rect 1653 651 1674 671
rect 3208 737 3234 759
rect 3473 766 3492 786
rect 3550 766 3569 786
rect 4202 829 4223 849
rect 1864 622 1885 663
rect 2026 558 2052 584
rect 1651 502 1672 522
rect 2076 505 2096 525
rect 203 439 228 458
rect 426 439 455 466
rect 500 442 529 469
rect 1158 434 1178 454
rect 3759 736 3779 756
rect 4408 721 4437 748
rect 4482 724 4511 751
rect 4709 732 4734 751
rect 2841 665 2861 685
rect 3051 667 3071 684
rect 3265 668 3286 688
rect 2885 606 2911 632
rect 714 341 735 361
rect 1368 404 1387 424
rect 1445 404 1464 424
rect 1703 431 1729 453
rect 3263 519 3284 539
rect 2820 426 2840 446
rect 3469 411 3498 438
rect 3543 414 3572 441
rect 4411 522 4430 542
rect 4488 522 4507 542
rect 1087 248 1113 274
rect 712 192 733 212
rect 922 190 945 210
rect 1137 195 1157 215
rect 3779 421 3799 441
rect 3989 424 4014 444
rect 4203 424 4224 444
rect 3823 362 3849 388
rect 4201 275 4222 295
rect 3758 182 3778 202
rect 4711 281 4740 310
rect 4407 167 4436 194
rect 4481 170 4510 197
rect 429 94 448 114
rect 506 94 525 114
rect 757 11 786 32
rect 4792 15 4821 36
rect 1673 -120 1702 -93
rect 1747 -117 1776 -90
rect 2405 -125 2425 -105
rect 1961 -218 1982 -198
rect 2334 -311 2360 -285
rect 1959 -367 1980 -347
rect 2165 -368 2199 -348
rect 2384 -364 2404 -344
rect 2486 -426 2513 -405
rect 1676 -465 1695 -445
rect 1753 -465 1772 -445
<< metal1 >>
rect 3719 8835 4021 8837
rect 1150 8812 1185 8814
rect 186 8809 1185 8812
rect 185 8785 1185 8809
rect 185 8630 233 8785
rect 419 8744 529 8758
rect 419 8741 497 8744
rect 419 8714 423 8741
rect 452 8717 497 8741
rect 526 8717 529 8744
rect 1150 8734 1185 8785
rect 452 8714 529 8717
rect 419 8699 529 8714
rect 1148 8729 1185 8734
rect 1148 8709 1155 8729
rect 1175 8709 1185 8729
rect 1148 8702 1185 8709
rect 3658 8806 4021 8835
rect 3658 8804 3719 8806
rect 1148 8701 1183 8702
rect 185 8601 193 8630
rect 222 8601 233 8630
rect 185 8596 233 8601
rect 704 8636 736 8643
rect 704 8616 711 8636
rect 732 8616 736 8636
rect 704 8551 736 8616
rect 1074 8551 1114 8552
rect 704 8549 1116 8551
rect 704 8523 1084 8549
rect 1110 8523 1116 8549
rect 704 8515 1116 8523
rect 704 8487 736 8515
rect 1149 8495 1183 8701
rect 3200 8584 3237 8586
rect 3658 8584 3691 8804
rect 3979 8725 4021 8806
rect 4401 8817 4512 8834
rect 4401 8797 4408 8817
rect 4427 8797 4485 8817
rect 4504 8797 4512 8817
rect 4401 8775 4512 8797
rect 3768 8723 3803 8724
rect 2087 8568 2121 8569
rect 1218 8533 2122 8568
rect 3200 8555 3691 8584
rect 704 8467 709 8487
rect 730 8467 736 8487
rect 704 8460 736 8467
rect 911 8487 950 8493
rect 911 8467 919 8487
rect 944 8467 950 8487
rect 911 8460 950 8467
rect 1127 8490 1183 8495
rect 1127 8470 1134 8490
rect 1154 8470 1183 8490
rect 1127 8463 1183 8470
rect 1127 8462 1162 8463
rect 919 8414 950 8460
rect 418 8389 529 8411
rect 418 8369 426 8389
rect 445 8369 503 8389
rect 522 8369 529 8389
rect 918 8397 950 8414
rect 1219 8397 1256 8533
rect 1357 8500 1467 8514
rect 1357 8497 1435 8500
rect 1357 8470 1361 8497
rect 1390 8473 1435 8497
rect 1464 8473 1467 8500
rect 2087 8490 2121 8533
rect 1390 8470 1467 8473
rect 1357 8455 1467 8470
rect 2086 8485 2121 8490
rect 3200 8489 3237 8555
rect 3658 8554 3691 8555
rect 3747 8716 3803 8723
rect 3747 8696 3776 8716
rect 3796 8696 3803 8716
rect 3747 8691 3803 8696
rect 3977 8721 4021 8725
rect 3977 8701 3988 8721
rect 4011 8701 4021 8721
rect 3977 8694 4021 8701
rect 4194 8719 4226 8726
rect 4194 8699 4200 8719
rect 4221 8699 4226 8719
rect 3977 8692 4020 8694
rect 2086 8465 2093 8485
rect 2113 8465 2121 8485
rect 2086 8457 2121 8465
rect 918 8384 1256 8397
rect 418 8352 529 8369
rect 919 8365 1256 8384
rect 1198 8364 1256 8365
rect 1642 8392 1674 8399
rect 1642 8372 1649 8392
rect 1670 8372 1674 8392
rect 1642 8307 1674 8372
rect 2012 8307 2052 8308
rect 1642 8305 2054 8307
rect 1642 8279 2022 8305
rect 2048 8279 2054 8305
rect 1642 8271 2054 8279
rect 188 8232 1184 8258
rect 1642 8243 1674 8271
rect 190 8179 232 8232
rect 190 8160 199 8179
rect 224 8160 232 8179
rect 190 8150 232 8160
rect 418 8190 528 8204
rect 418 8187 496 8190
rect 418 8160 422 8187
rect 451 8163 496 8187
rect 525 8163 528 8190
rect 1148 8180 1182 8232
rect 1642 8223 1647 8243
rect 1668 8223 1674 8243
rect 1642 8216 1674 8223
rect 1852 8244 1890 8254
rect 2087 8251 2121 8457
rect 3195 8480 3237 8489
rect 3195 8458 3204 8480
rect 3230 8458 3237 8480
rect 3462 8507 3573 8524
rect 3462 8487 3469 8507
rect 3488 8487 3546 8507
rect 3565 8487 3573 8507
rect 3462 8465 3573 8487
rect 3747 8485 3781 8691
rect 4194 8671 4226 8699
rect 3814 8663 4226 8671
rect 3814 8637 3820 8663
rect 3846 8637 4226 8663
rect 3814 8635 4226 8637
rect 3816 8634 3856 8635
rect 4194 8570 4226 8635
rect 4194 8550 4198 8570
rect 4219 8550 4226 8570
rect 4194 8543 4226 8550
rect 3747 8477 3782 8485
rect 3195 8448 3237 8458
rect 3747 8457 3755 8477
rect 3775 8457 3782 8477
rect 3747 8452 3782 8457
rect 4401 8472 4511 8487
rect 4401 8469 4478 8472
rect 3195 8447 3236 8448
rect 2829 8413 2864 8414
rect 1852 8227 1862 8244
rect 1882 8227 1890 8244
rect 1693 8184 1734 8185
rect 451 8160 528 8163
rect 418 8145 528 8160
rect 1147 8175 1182 8180
rect 1147 8155 1154 8175
rect 1174 8155 1182 8175
rect 1692 8174 1734 8184
rect 1147 8147 1182 8155
rect 703 8082 735 8089
rect 703 8062 710 8082
rect 731 8062 735 8082
rect 703 7997 735 8062
rect 1073 7997 1113 7998
rect 703 7995 1115 7997
rect 703 7969 1083 7995
rect 1109 7969 1115 7995
rect 703 7961 1115 7969
rect 703 7933 735 7961
rect 1148 7941 1182 8147
rect 1356 8145 1467 8167
rect 1356 8125 1364 8145
rect 1383 8125 1441 8145
rect 1460 8125 1467 8145
rect 1356 8108 1467 8125
rect 1692 8152 1699 8174
rect 1725 8152 1734 8174
rect 1692 8143 1734 8152
rect 909 7938 952 7940
rect 703 7913 708 7933
rect 729 7913 735 7933
rect 703 7906 735 7913
rect 908 7931 952 7938
rect 908 7911 918 7931
rect 941 7911 952 7931
rect 908 7907 952 7911
rect 1126 7936 1182 7941
rect 1126 7916 1133 7936
rect 1153 7916 1182 7936
rect 1126 7909 1182 7916
rect 1238 8077 1271 8078
rect 1692 8077 1729 8143
rect 1238 8048 1729 8077
rect 1126 7908 1161 7909
rect 417 7835 528 7857
rect 417 7815 425 7835
rect 444 7815 502 7835
rect 521 7815 528 7835
rect 417 7798 528 7815
rect 908 7826 950 7907
rect 1238 7828 1271 8048
rect 1692 8046 1729 8048
rect 1498 7908 1608 7922
rect 1498 7905 1576 7908
rect 1498 7878 1502 7905
rect 1531 7881 1576 7905
rect 1605 7881 1608 7908
rect 1531 7878 1608 7881
rect 1498 7863 1608 7878
rect 1852 7889 1890 8227
rect 2065 8246 2121 8251
rect 2065 8226 2072 8246
rect 2092 8226 2121 8246
rect 2065 8219 2121 8226
rect 2808 8406 2864 8413
rect 2808 8386 2837 8406
rect 2857 8386 2864 8406
rect 2808 8381 2864 8386
rect 3255 8409 3287 8416
rect 3255 8389 3261 8409
rect 3282 8389 3287 8409
rect 3747 8400 3781 8452
rect 4401 8442 4404 8469
rect 4433 8445 4478 8469
rect 4507 8445 4511 8472
rect 4433 8442 4511 8445
rect 4401 8428 4511 8442
rect 4697 8472 4739 8482
rect 4697 8453 4705 8472
rect 4730 8453 4739 8472
rect 4697 8400 4739 8453
rect 2065 8218 2100 8219
rect 2808 8175 2842 8381
rect 3255 8361 3287 8389
rect 3745 8374 4741 8400
rect 2875 8353 3287 8361
rect 2875 8327 2881 8353
rect 2907 8327 3287 8353
rect 2875 8325 3287 8327
rect 2877 8324 2917 8325
rect 3037 8289 3076 8304
rect 3037 8248 3048 8289
rect 3069 8248 3076 8289
rect 2807 8167 2843 8175
rect 2807 8147 2816 8167
rect 2836 8147 2843 8167
rect 2807 8146 2843 8147
rect 2807 8135 2841 8146
rect 3037 7975 3076 8248
rect 3255 8260 3287 8325
rect 3255 8240 3259 8260
rect 3280 8240 3287 8260
rect 3255 8233 3287 8240
rect 3673 8267 3731 8268
rect 3673 8248 4010 8267
rect 4400 8263 4511 8280
rect 3673 8235 4011 8248
rect 3177 8171 3230 8174
rect 3177 8154 3189 8171
rect 3221 8154 3230 8171
rect 3177 8146 3230 8154
rect 3176 8099 3230 8146
rect 3462 8162 3572 8177
rect 3462 8159 3539 8162
rect 3462 8132 3465 8159
rect 3494 8135 3539 8159
rect 3568 8135 3572 8162
rect 3494 8132 3572 8135
rect 3462 8118 3572 8132
rect 3673 8099 3710 8235
rect 3979 8218 4011 8235
rect 4400 8243 4407 8263
rect 4426 8243 4484 8263
rect 4503 8243 4511 8263
rect 4400 8221 4511 8243
rect 3979 8172 4010 8218
rect 3767 8169 3802 8170
rect 3746 8162 3802 8169
rect 3746 8142 3775 8162
rect 3795 8142 3802 8162
rect 3746 8137 3802 8142
rect 3979 8165 4018 8172
rect 3979 8145 3985 8165
rect 4010 8145 4018 8165
rect 3979 8139 4018 8145
rect 4193 8165 4225 8172
rect 4193 8145 4199 8165
rect 4220 8145 4225 8165
rect 3176 8064 3711 8099
rect 3176 8060 3229 8064
rect 3037 7948 3041 7975
rect 3072 7948 3076 7975
rect 3322 7996 3433 8013
rect 3322 7976 3329 7996
rect 3348 7976 3406 7996
rect 3425 7976 3433 7996
rect 3322 7954 3433 7976
rect 3037 7941 3076 7948
rect 3746 7931 3780 8137
rect 4193 8117 4225 8145
rect 3813 8109 4225 8117
rect 3813 8083 3819 8109
rect 3845 8083 4225 8109
rect 3813 8081 4225 8083
rect 3815 8080 3855 8081
rect 4193 8016 4225 8081
rect 4193 7996 4197 8016
rect 4218 7996 4225 8016
rect 4193 7989 4225 7996
rect 4696 8031 4744 8036
rect 4696 8002 4707 8031
rect 4736 8002 4744 8031
rect 3746 7930 3781 7931
rect 3744 7923 3781 7930
rect 2689 7902 2724 7903
rect 2230 7898 2262 7899
rect 1852 7872 1860 7889
rect 1880 7872 1890 7889
rect 1852 7866 1890 7872
rect 2227 7893 2262 7898
rect 2227 7873 2234 7893
rect 2254 7873 2262 7893
rect 2227 7865 2262 7873
rect 1210 7826 1271 7828
rect 908 7797 1271 7826
rect 1783 7800 1815 7807
rect 908 7795 1210 7797
rect 1783 7780 1790 7800
rect 1811 7780 1815 7800
rect 1783 7715 1815 7780
rect 2153 7715 2193 7716
rect 1783 7713 2195 7715
rect 1151 7709 1186 7711
rect 187 7706 1186 7709
rect 186 7682 1186 7706
rect 186 7527 234 7682
rect 420 7641 530 7655
rect 420 7638 498 7641
rect 420 7611 424 7638
rect 453 7614 498 7638
rect 527 7614 530 7641
rect 1151 7631 1186 7682
rect 453 7611 530 7614
rect 420 7596 530 7611
rect 1149 7626 1186 7631
rect 1149 7606 1156 7626
rect 1176 7606 1186 7626
rect 1783 7687 2163 7713
rect 2189 7687 2195 7713
rect 1783 7679 2195 7687
rect 1783 7651 1815 7679
rect 1783 7631 1788 7651
rect 1809 7631 1815 7651
rect 1783 7624 1815 7631
rect 1989 7650 2031 7661
rect 2228 7659 2262 7865
rect 2666 7895 2724 7902
rect 2666 7875 2697 7895
rect 2717 7875 2724 7895
rect 2666 7870 2724 7875
rect 3115 7898 3147 7905
rect 3115 7878 3121 7898
rect 3142 7878 3147 7898
rect 2666 7722 2702 7870
rect 3115 7850 3147 7878
rect 2735 7842 3147 7850
rect 2735 7816 2741 7842
rect 2767 7816 3147 7842
rect 3744 7903 3754 7923
rect 3774 7903 3781 7923
rect 3744 7898 3781 7903
rect 4400 7918 4510 7933
rect 4400 7915 4477 7918
rect 3744 7847 3779 7898
rect 4400 7888 4403 7915
rect 4432 7891 4477 7915
rect 4506 7891 4510 7918
rect 4432 7888 4510 7891
rect 4400 7874 4510 7888
rect 4696 7847 4744 8002
rect 3744 7823 4744 7847
rect 3744 7820 4743 7823
rect 3744 7818 3779 7820
rect 2735 7814 3147 7816
rect 2737 7813 2777 7814
rect 1989 7629 1996 7650
rect 2023 7629 2031 7650
rect 1149 7599 1186 7606
rect 1149 7598 1184 7599
rect 186 7498 194 7527
rect 223 7498 234 7527
rect 186 7493 234 7498
rect 705 7533 737 7540
rect 705 7513 712 7533
rect 733 7513 737 7533
rect 705 7448 737 7513
rect 1075 7448 1115 7449
rect 705 7446 1117 7448
rect 705 7420 1085 7446
rect 1111 7420 1117 7446
rect 705 7412 1117 7420
rect 705 7384 737 7412
rect 1150 7392 1184 7598
rect 1854 7581 1893 7588
rect 1497 7553 1608 7575
rect 1497 7533 1505 7553
rect 1524 7533 1582 7553
rect 1601 7533 1608 7553
rect 1497 7516 1608 7533
rect 1854 7554 1858 7581
rect 1889 7554 1893 7581
rect 1701 7465 1754 7469
rect 1219 7430 1754 7465
rect 705 7364 710 7384
rect 731 7364 737 7384
rect 705 7357 737 7364
rect 912 7384 951 7390
rect 912 7364 920 7384
rect 945 7364 951 7384
rect 912 7357 951 7364
rect 1128 7387 1184 7392
rect 1128 7367 1135 7387
rect 1155 7367 1184 7387
rect 1128 7360 1184 7367
rect 1128 7359 1163 7360
rect 920 7311 951 7357
rect 419 7286 530 7308
rect 419 7266 427 7286
rect 446 7266 504 7286
rect 523 7266 530 7286
rect 919 7294 951 7311
rect 1220 7294 1257 7430
rect 1358 7397 1468 7411
rect 1358 7394 1436 7397
rect 1358 7367 1362 7394
rect 1391 7370 1436 7394
rect 1465 7370 1468 7397
rect 1391 7367 1468 7370
rect 1358 7352 1468 7367
rect 1700 7383 1754 7430
rect 1700 7375 1753 7383
rect 1700 7358 1709 7375
rect 1741 7358 1753 7375
rect 1700 7355 1753 7358
rect 919 7281 1257 7294
rect 419 7249 530 7266
rect 920 7262 1257 7281
rect 1199 7261 1257 7262
rect 1643 7289 1675 7296
rect 1643 7269 1650 7289
rect 1671 7269 1675 7289
rect 1643 7204 1675 7269
rect 1854 7281 1893 7554
rect 1989 7458 2031 7629
rect 2206 7654 2262 7659
rect 2206 7634 2213 7654
rect 2233 7634 2262 7654
rect 2206 7627 2262 7634
rect 2669 7664 2702 7722
rect 2899 7774 2937 7784
rect 2899 7736 2908 7774
rect 2931 7736 2937 7774
rect 2669 7656 2703 7664
rect 2669 7636 2676 7656
rect 2696 7636 2703 7656
rect 2669 7631 2703 7636
rect 2669 7630 2700 7631
rect 2206 7626 2241 7627
rect 2899 7600 2937 7736
rect 3115 7749 3147 7814
rect 3115 7729 3119 7749
rect 3140 7729 3147 7749
rect 3720 7732 4022 7734
rect 3115 7722 3147 7729
rect 3659 7703 4022 7732
rect 3659 7701 3720 7703
rect 3040 7657 3078 7663
rect 3040 7640 3050 7657
rect 3070 7640 3078 7657
rect 1989 7424 2233 7458
rect 2899 7446 2943 7600
rect 2736 7444 2943 7446
rect 2196 7416 2233 7424
rect 2089 7383 2123 7394
rect 2087 7382 2123 7383
rect 2087 7362 2094 7382
rect 2114 7362 2123 7382
rect 2087 7354 2123 7362
rect 1854 7240 1861 7281
rect 1882 7240 1893 7281
rect 1854 7225 1893 7240
rect 2013 7204 2053 7205
rect 1643 7202 2055 7204
rect 1643 7176 2023 7202
rect 2049 7176 2055 7202
rect 1643 7168 2055 7176
rect 189 7129 1185 7155
rect 1643 7140 1675 7168
rect 2088 7148 2122 7354
rect 191 7076 233 7129
rect 191 7057 200 7076
rect 225 7057 233 7076
rect 191 7047 233 7057
rect 419 7087 529 7101
rect 419 7084 497 7087
rect 419 7057 423 7084
rect 452 7060 497 7084
rect 526 7060 529 7087
rect 1149 7077 1183 7129
rect 1643 7120 1648 7140
rect 1669 7120 1675 7140
rect 1643 7113 1675 7120
rect 2066 7143 2122 7148
rect 2066 7123 2073 7143
rect 2093 7123 2122 7143
rect 2066 7116 2122 7123
rect 2066 7115 2101 7116
rect 1694 7081 1735 7082
rect 452 7057 529 7060
rect 419 7042 529 7057
rect 1148 7072 1183 7077
rect 1148 7052 1155 7072
rect 1175 7052 1183 7072
rect 1693 7071 1735 7081
rect 1148 7044 1183 7052
rect 704 6979 736 6986
rect 704 6959 711 6979
rect 732 6959 736 6979
rect 704 6894 736 6959
rect 1074 6894 1114 6895
rect 704 6892 1116 6894
rect 704 6866 1084 6892
rect 1110 6866 1116 6892
rect 704 6858 1116 6866
rect 704 6830 736 6858
rect 1149 6838 1183 7044
rect 1357 7042 1468 7064
rect 1357 7022 1365 7042
rect 1384 7022 1442 7042
rect 1461 7022 1468 7042
rect 1357 7005 1468 7022
rect 1693 7049 1700 7071
rect 1726 7049 1735 7071
rect 1693 7040 1735 7049
rect 910 6835 953 6837
rect 704 6810 709 6830
rect 730 6810 736 6830
rect 704 6803 736 6810
rect 909 6828 953 6835
rect 909 6808 919 6828
rect 942 6808 953 6828
rect 909 6804 953 6808
rect 1127 6833 1183 6838
rect 1127 6813 1134 6833
rect 1154 6813 1183 6833
rect 1127 6806 1183 6813
rect 1239 6974 1272 6975
rect 1693 6974 1730 7040
rect 1239 6945 1730 6974
rect 1127 6805 1162 6806
rect 418 6732 529 6754
rect 418 6712 426 6732
rect 445 6712 503 6732
rect 522 6712 529 6732
rect 418 6696 529 6712
rect 909 6723 951 6804
rect 1239 6725 1272 6945
rect 1693 6943 1730 6945
rect 1468 6818 1578 6832
rect 1468 6815 1546 6818
rect 1468 6788 1472 6815
rect 1501 6791 1546 6815
rect 1575 6791 1578 6818
rect 1501 6788 1578 6791
rect 1468 6773 1578 6788
rect 2196 6803 2234 7416
rect 2712 7411 2943 7444
rect 2712 6870 2762 7411
rect 2899 7407 2943 7411
rect 2830 7310 2865 7311
rect 2809 7303 2865 7310
rect 2809 7283 2838 7303
rect 2858 7283 2865 7303
rect 2809 7278 2865 7283
rect 3040 7302 3078 7640
rect 3322 7651 3432 7666
rect 3322 7648 3399 7651
rect 3322 7621 3325 7648
rect 3354 7624 3399 7648
rect 3428 7624 3432 7651
rect 3354 7621 3432 7624
rect 3322 7607 3432 7621
rect 3201 7481 3238 7483
rect 3659 7481 3692 7701
rect 3980 7622 4022 7703
rect 4402 7714 4513 7731
rect 4402 7694 4409 7714
rect 4428 7694 4486 7714
rect 4505 7694 4513 7714
rect 4402 7672 4513 7694
rect 3769 7620 3804 7621
rect 3201 7452 3692 7481
rect 3201 7386 3238 7452
rect 3659 7451 3692 7452
rect 3748 7613 3804 7620
rect 3748 7593 3777 7613
rect 3797 7593 3804 7613
rect 3748 7588 3804 7593
rect 3978 7618 4022 7622
rect 3978 7598 3989 7618
rect 4012 7598 4022 7618
rect 3978 7591 4022 7598
rect 4195 7616 4227 7623
rect 4195 7596 4201 7616
rect 4222 7596 4227 7616
rect 3978 7589 4021 7591
rect 3196 7377 3238 7386
rect 3196 7355 3205 7377
rect 3231 7355 3238 7377
rect 3463 7404 3574 7421
rect 3463 7384 3470 7404
rect 3489 7384 3547 7404
rect 3566 7384 3574 7404
rect 3463 7362 3574 7384
rect 3748 7382 3782 7588
rect 4195 7568 4227 7596
rect 3815 7560 4227 7568
rect 3815 7534 3821 7560
rect 3847 7534 4227 7560
rect 3815 7532 4227 7534
rect 3817 7531 3857 7532
rect 4195 7467 4227 7532
rect 4195 7447 4199 7467
rect 4220 7447 4227 7467
rect 4195 7440 4227 7447
rect 3748 7374 3783 7382
rect 3196 7345 3238 7355
rect 3748 7354 3756 7374
rect 3776 7354 3783 7374
rect 3748 7349 3783 7354
rect 4402 7369 4512 7384
rect 4402 7366 4479 7369
rect 3196 7344 3237 7345
rect 3040 7285 3048 7302
rect 3068 7285 3078 7302
rect 2809 7072 2843 7278
rect 3040 7275 3078 7285
rect 3256 7306 3288 7313
rect 3256 7286 3262 7306
rect 3283 7286 3288 7306
rect 3748 7297 3782 7349
rect 4402 7339 4405 7366
rect 4434 7342 4479 7366
rect 4508 7342 4512 7369
rect 4434 7339 4512 7342
rect 4402 7325 4512 7339
rect 4698 7369 4740 7379
rect 4698 7350 4706 7369
rect 4731 7350 4740 7369
rect 4698 7297 4740 7350
rect 3256 7258 3288 7286
rect 3746 7271 4742 7297
rect 2876 7250 3288 7258
rect 2876 7224 2882 7250
rect 2908 7224 3288 7250
rect 2876 7222 3288 7224
rect 2878 7221 2918 7222
rect 3256 7157 3288 7222
rect 3256 7137 3260 7157
rect 3281 7137 3288 7157
rect 3256 7130 3288 7137
rect 3674 7164 3732 7165
rect 3674 7145 4011 7164
rect 4401 7160 4512 7177
rect 3674 7132 4012 7145
rect 2809 7064 2844 7072
rect 2809 7044 2817 7064
rect 2837 7044 2844 7064
rect 2809 7039 2844 7044
rect 3463 7059 3573 7074
rect 3463 7056 3540 7059
rect 2809 6996 2843 7039
rect 3463 7029 3466 7056
rect 3495 7032 3540 7056
rect 3569 7032 3573 7059
rect 3495 7029 3573 7032
rect 3463 7015 3573 7029
rect 3674 6996 3711 7132
rect 3980 7115 4012 7132
rect 4401 7140 4408 7160
rect 4427 7140 4485 7160
rect 4504 7140 4512 7160
rect 4401 7118 4512 7140
rect 3980 7069 4011 7115
rect 3768 7066 3803 7067
rect 3747 7059 3803 7066
rect 3747 7039 3776 7059
rect 3796 7039 3803 7059
rect 3747 7034 3803 7039
rect 3980 7062 4019 7069
rect 3980 7042 3986 7062
rect 4011 7042 4019 7062
rect 3980 7036 4019 7042
rect 4194 7062 4226 7069
rect 4194 7042 4200 7062
rect 4221 7042 4226 7062
rect 2808 6961 3712 6996
rect 2809 6960 2843 6961
rect 2690 6861 2762 6870
rect 2690 6832 2707 6861
rect 2755 6832 2762 6861
rect 3353 6880 3464 6897
rect 3353 6860 3360 6880
rect 3379 6860 3437 6880
rect 3456 6860 3464 6880
rect 3353 6838 3464 6860
rect 2690 6825 2762 6832
rect 3747 6828 3781 7034
rect 4194 7014 4226 7042
rect 3814 7006 4226 7014
rect 3814 6980 3820 7006
rect 3846 6980 4226 7006
rect 3814 6978 4226 6980
rect 3816 6977 3856 6978
rect 4194 6913 4226 6978
rect 4194 6893 4198 6913
rect 4219 6893 4226 6913
rect 4194 6886 4226 6893
rect 4697 6928 4745 6933
rect 4697 6899 4708 6928
rect 4737 6899 4745 6928
rect 3747 6827 3782 6828
rect 2690 6815 2760 6825
rect 3745 6820 3782 6827
rect 2196 6783 2204 6803
rect 2224 6783 2234 6803
rect 3745 6800 3755 6820
rect 3775 6800 3782 6820
rect 3745 6795 3782 6800
rect 4401 6815 4511 6830
rect 4401 6812 4478 6815
rect 2720 6786 2755 6787
rect 2196 6776 2234 6783
rect 2699 6779 2755 6786
rect 2197 6775 2232 6776
rect 1211 6723 1272 6725
rect 909 6694 1272 6723
rect 1753 6710 1785 6717
rect 909 6692 1211 6694
rect 1753 6690 1760 6710
rect 1781 6690 1785 6710
rect 1753 6625 1785 6690
rect 2123 6625 2163 6626
rect 1753 6623 2165 6625
rect 1151 6606 1186 6608
rect 187 6603 1186 6606
rect 186 6579 1186 6603
rect 186 6424 234 6579
rect 420 6538 530 6552
rect 420 6535 498 6538
rect 420 6508 424 6535
rect 453 6511 498 6535
rect 527 6511 530 6538
rect 1151 6528 1186 6579
rect 1753 6597 2133 6623
rect 2159 6597 2165 6623
rect 1753 6589 2165 6597
rect 1753 6561 1785 6589
rect 1753 6541 1758 6561
rect 1779 6541 1785 6561
rect 1753 6534 1785 6541
rect 1959 6560 2004 6572
rect 2198 6569 2232 6775
rect 1959 6541 1966 6560
rect 1995 6541 2004 6560
rect 453 6508 530 6511
rect 420 6493 530 6508
rect 1149 6523 1186 6528
rect 1149 6503 1156 6523
rect 1176 6503 1186 6523
rect 1149 6496 1186 6503
rect 1149 6495 1184 6496
rect 186 6395 194 6424
rect 223 6395 234 6424
rect 186 6390 234 6395
rect 705 6430 737 6437
rect 705 6410 712 6430
rect 733 6410 737 6430
rect 705 6345 737 6410
rect 1075 6345 1115 6346
rect 705 6343 1117 6345
rect 705 6317 1085 6343
rect 1111 6317 1117 6343
rect 705 6309 1117 6317
rect 705 6281 737 6309
rect 1150 6289 1184 6495
rect 1467 6463 1578 6485
rect 1467 6443 1475 6463
rect 1494 6443 1552 6463
rect 1571 6443 1578 6463
rect 1467 6426 1578 6443
rect 1959 6458 2004 6541
rect 2176 6564 2232 6569
rect 2176 6544 2183 6564
rect 2203 6544 2232 6564
rect 2699 6759 2728 6779
rect 2748 6759 2755 6779
rect 2699 6754 2755 6759
rect 3146 6782 3178 6789
rect 3146 6762 3152 6782
rect 3173 6762 3178 6782
rect 2699 6548 2733 6754
rect 3146 6734 3178 6762
rect 2766 6726 3178 6734
rect 2766 6700 2772 6726
rect 2798 6700 3178 6726
rect 3745 6744 3780 6795
rect 4401 6785 4404 6812
rect 4433 6788 4478 6812
rect 4507 6788 4511 6815
rect 4433 6785 4511 6788
rect 4401 6771 4511 6785
rect 4697 6744 4745 6899
rect 3745 6720 4745 6744
rect 3745 6717 4744 6720
rect 3745 6715 3780 6717
rect 2766 6698 3178 6700
rect 2768 6697 2808 6698
rect 2934 6657 2969 6675
rect 2934 6625 2937 6657
rect 2964 6625 2969 6657
rect 2699 6547 2734 6548
rect 2176 6537 2232 6544
rect 2697 6540 2735 6547
rect 2176 6536 2211 6537
rect 2697 6536 2707 6540
rect 2691 6522 2707 6536
rect 2727 6536 2735 6540
rect 2727 6522 2741 6536
rect 2691 6515 2741 6522
rect 2324 6458 2374 6460
rect 1959 6424 2374 6458
rect 2088 6362 2122 6363
rect 1219 6327 2123 6362
rect 2171 6351 2239 6362
rect 2171 6330 2176 6351
rect 705 6261 710 6281
rect 731 6261 737 6281
rect 705 6254 737 6261
rect 912 6281 951 6287
rect 912 6261 920 6281
rect 945 6261 951 6281
rect 912 6254 951 6261
rect 1128 6284 1184 6289
rect 1128 6264 1135 6284
rect 1155 6264 1184 6284
rect 1128 6257 1184 6264
rect 1128 6256 1163 6257
rect 920 6208 951 6254
rect 419 6183 530 6205
rect 419 6163 427 6183
rect 446 6163 504 6183
rect 523 6163 530 6183
rect 919 6191 951 6208
rect 1220 6191 1257 6327
rect 1358 6294 1468 6308
rect 1358 6291 1436 6294
rect 1358 6264 1362 6291
rect 1391 6267 1436 6291
rect 1465 6267 1468 6294
rect 2088 6284 2122 6327
rect 1391 6264 1468 6267
rect 1358 6249 1468 6264
rect 2087 6279 2122 6284
rect 2087 6259 2094 6279
rect 2114 6259 2122 6279
rect 2087 6251 2122 6259
rect 919 6178 1257 6191
rect 419 6146 530 6163
rect 920 6159 1257 6178
rect 1199 6158 1257 6159
rect 1643 6186 1675 6193
rect 1643 6166 1650 6186
rect 1671 6166 1675 6186
rect 1643 6101 1675 6166
rect 2013 6101 2053 6102
rect 1643 6099 2055 6101
rect 1643 6073 2023 6099
rect 2049 6073 2055 6099
rect 1643 6065 2055 6073
rect 189 6026 1185 6052
rect 1643 6037 1675 6065
rect 191 5973 233 6026
rect 191 5954 200 5973
rect 225 5954 233 5973
rect 191 5944 233 5954
rect 419 5984 529 5998
rect 419 5981 497 5984
rect 419 5954 423 5981
rect 452 5957 497 5981
rect 526 5957 529 5984
rect 1149 5974 1183 6026
rect 1643 6017 1648 6037
rect 1669 6017 1675 6037
rect 1643 6010 1675 6017
rect 1853 6038 1891 6048
rect 2088 6045 2122 6251
rect 1853 6021 1863 6038
rect 1883 6021 1891 6038
rect 1694 5978 1735 5979
rect 452 5954 529 5957
rect 419 5939 529 5954
rect 1148 5969 1183 5974
rect 1148 5949 1155 5969
rect 1175 5949 1183 5969
rect 1693 5968 1735 5978
rect 1148 5941 1183 5949
rect 704 5876 736 5883
rect 704 5856 711 5876
rect 732 5856 736 5876
rect 704 5791 736 5856
rect 1074 5791 1114 5792
rect 704 5789 1116 5791
rect 704 5763 1084 5789
rect 1110 5763 1116 5789
rect 704 5755 1116 5763
rect 704 5727 736 5755
rect 1149 5735 1183 5941
rect 1357 5939 1468 5961
rect 1357 5919 1365 5939
rect 1384 5919 1442 5939
rect 1461 5919 1468 5939
rect 1357 5902 1468 5919
rect 1693 5946 1700 5968
rect 1726 5946 1735 5968
rect 1693 5937 1735 5946
rect 910 5732 953 5734
rect 704 5707 709 5727
rect 730 5707 736 5727
rect 704 5700 736 5707
rect 909 5725 953 5732
rect 909 5705 919 5725
rect 942 5705 953 5725
rect 909 5701 953 5705
rect 1127 5730 1183 5735
rect 1127 5710 1134 5730
rect 1154 5710 1183 5730
rect 1127 5703 1183 5710
rect 1239 5871 1272 5872
rect 1693 5871 1730 5937
rect 1239 5842 1730 5871
rect 1127 5702 1162 5703
rect 418 5629 529 5651
rect 418 5609 426 5629
rect 445 5609 503 5629
rect 522 5609 529 5629
rect 418 5592 529 5609
rect 909 5620 951 5701
rect 1239 5622 1272 5842
rect 1693 5840 1730 5842
rect 1499 5702 1609 5716
rect 1499 5699 1577 5702
rect 1499 5672 1503 5699
rect 1532 5675 1577 5699
rect 1606 5675 1609 5702
rect 1532 5672 1609 5675
rect 1499 5657 1609 5672
rect 1853 5683 1891 6021
rect 2066 6040 2122 6045
rect 2066 6020 2073 6040
rect 2093 6020 2122 6040
rect 2066 6013 2122 6020
rect 2169 6322 2176 6330
rect 2224 6322 2239 6351
rect 2169 6313 2239 6322
rect 2066 6012 2101 6013
rect 1988 5912 2032 5916
rect 2169 5912 2219 6313
rect 2324 6296 2374 6424
rect 2557 6437 2667 6439
rect 2934 6437 2969 6625
rect 3146 6633 3178 6698
rect 3146 6613 3150 6633
rect 3171 6613 3178 6633
rect 3720 6629 4022 6631
rect 3146 6606 3178 6613
rect 3659 6600 4022 6629
rect 3659 6598 3720 6600
rect 2557 6407 2969 6437
rect 2557 6382 2601 6407
rect 2640 6404 2969 6407
rect 3088 6538 3122 6544
rect 3088 6518 3097 6538
rect 3118 6518 3122 6538
rect 1988 5879 2219 5912
rect 1988 5877 2195 5879
rect 1988 5723 2032 5877
rect 1853 5666 1861 5683
rect 1881 5666 1891 5683
rect 1853 5660 1891 5666
rect 1211 5620 1272 5622
rect 909 5591 1272 5620
rect 1784 5594 1816 5601
rect 909 5589 1211 5591
rect 1784 5574 1791 5594
rect 1812 5574 1816 5594
rect 1784 5509 1816 5574
rect 1994 5587 2032 5723
rect 2231 5692 2262 5693
rect 2228 5687 2262 5692
rect 2228 5667 2235 5687
rect 2255 5667 2262 5687
rect 2228 5659 2262 5667
rect 1994 5549 2000 5587
rect 2023 5549 2032 5587
rect 1994 5539 2032 5549
rect 2229 5601 2262 5659
rect 2154 5509 2194 5510
rect 1784 5507 2196 5509
rect 1152 5503 1187 5505
rect 188 5500 1187 5503
rect 187 5476 1187 5500
rect 187 5321 235 5476
rect 421 5435 531 5449
rect 421 5432 499 5435
rect 421 5405 425 5432
rect 454 5408 499 5432
rect 528 5408 531 5435
rect 1152 5425 1187 5476
rect 454 5405 531 5408
rect 421 5390 531 5405
rect 1150 5420 1187 5425
rect 1150 5400 1157 5420
rect 1177 5400 1187 5420
rect 1784 5481 2164 5507
rect 2190 5481 2196 5507
rect 1784 5473 2196 5481
rect 1784 5445 1816 5473
rect 2229 5453 2265 5601
rect 1784 5425 1789 5445
rect 1810 5425 1816 5445
rect 1784 5418 1816 5425
rect 2207 5448 2265 5453
rect 2207 5428 2214 5448
rect 2234 5428 2265 5448
rect 2207 5421 2265 5428
rect 2207 5420 2242 5421
rect 1150 5393 1187 5400
rect 1150 5392 1185 5393
rect 187 5292 195 5321
rect 224 5292 235 5321
rect 187 5287 235 5292
rect 706 5327 738 5334
rect 706 5307 713 5327
rect 734 5307 738 5327
rect 706 5242 738 5307
rect 1076 5242 1116 5243
rect 706 5240 1118 5242
rect 706 5214 1086 5240
rect 1112 5214 1118 5240
rect 706 5206 1118 5214
rect 706 5178 738 5206
rect 1151 5186 1185 5392
rect 1855 5375 1894 5382
rect 1498 5347 1609 5369
rect 1498 5327 1506 5347
rect 1525 5327 1583 5347
rect 1602 5327 1609 5347
rect 1498 5310 1609 5327
rect 1855 5348 1859 5375
rect 1890 5348 1894 5375
rect 1702 5259 1755 5263
rect 1220 5224 1755 5259
rect 706 5158 711 5178
rect 732 5158 738 5178
rect 706 5151 738 5158
rect 913 5178 952 5184
rect 913 5158 921 5178
rect 946 5158 952 5178
rect 913 5151 952 5158
rect 1129 5181 1185 5186
rect 1129 5161 1136 5181
rect 1156 5161 1185 5181
rect 1129 5154 1185 5161
rect 1129 5153 1164 5154
rect 921 5105 952 5151
rect 420 5080 531 5102
rect 420 5060 428 5080
rect 447 5060 505 5080
rect 524 5060 531 5080
rect 920 5088 952 5105
rect 1221 5088 1258 5224
rect 1359 5191 1469 5205
rect 1359 5188 1437 5191
rect 1359 5161 1363 5188
rect 1392 5164 1437 5188
rect 1466 5164 1469 5191
rect 1392 5161 1469 5164
rect 1359 5146 1469 5161
rect 1701 5177 1755 5224
rect 1701 5169 1754 5177
rect 1701 5152 1710 5169
rect 1742 5152 1754 5169
rect 1701 5149 1754 5152
rect 920 5075 1258 5088
rect 420 5043 531 5060
rect 921 5056 1258 5075
rect 1200 5055 1258 5056
rect 1644 5083 1676 5090
rect 1644 5063 1651 5083
rect 1672 5063 1676 5083
rect 1644 4998 1676 5063
rect 1855 5075 1894 5348
rect 2090 5177 2124 5188
rect 2088 5176 2124 5177
rect 2088 5156 2095 5176
rect 2115 5156 2124 5176
rect 2088 5148 2124 5156
rect 1855 5034 1862 5075
rect 1883 5034 1894 5075
rect 1855 5019 1894 5034
rect 2014 4998 2054 4999
rect 1644 4996 2056 4998
rect 1644 4970 2024 4996
rect 2050 4970 2056 4996
rect 1644 4962 2056 4970
rect 190 4923 1186 4949
rect 1644 4934 1676 4962
rect 2089 4942 2123 5148
rect 192 4870 234 4923
rect 192 4851 201 4870
rect 226 4851 234 4870
rect 192 4841 234 4851
rect 420 4881 530 4895
rect 420 4878 498 4881
rect 420 4851 424 4878
rect 453 4854 498 4878
rect 527 4854 530 4881
rect 1150 4871 1184 4923
rect 1644 4914 1649 4934
rect 1670 4914 1676 4934
rect 1644 4907 1676 4914
rect 2067 4937 2123 4942
rect 2067 4917 2074 4937
rect 2094 4917 2123 4937
rect 2067 4910 2123 4917
rect 2067 4909 2102 4910
rect 1695 4875 1736 4876
rect 453 4851 530 4854
rect 420 4836 530 4851
rect 1149 4866 1184 4871
rect 1149 4846 1156 4866
rect 1176 4846 1184 4866
rect 1694 4865 1736 4875
rect 1149 4838 1184 4846
rect 705 4773 737 4780
rect 705 4753 712 4773
rect 733 4753 737 4773
rect 705 4688 737 4753
rect 1075 4688 1115 4689
rect 705 4686 1117 4688
rect 705 4660 1085 4686
rect 1111 4660 1117 4686
rect 705 4652 1117 4660
rect 705 4624 737 4652
rect 1150 4632 1184 4838
rect 1358 4836 1469 4858
rect 1358 4816 1366 4836
rect 1385 4816 1443 4836
rect 1462 4816 1469 4836
rect 1358 4799 1469 4816
rect 1694 4843 1701 4865
rect 1727 4843 1736 4865
rect 1694 4834 1736 4843
rect 911 4629 954 4631
rect 705 4604 710 4624
rect 731 4604 737 4624
rect 705 4597 737 4604
rect 910 4622 954 4629
rect 910 4602 920 4622
rect 943 4602 954 4622
rect 910 4598 954 4602
rect 1128 4627 1184 4632
rect 1128 4607 1135 4627
rect 1155 4607 1184 4627
rect 1128 4600 1184 4607
rect 1240 4768 1273 4769
rect 1694 4768 1731 4834
rect 2326 4811 2372 6296
rect 1240 4739 1731 4768
rect 1128 4599 1163 4600
rect 419 4526 530 4548
rect 419 4506 427 4526
rect 446 4506 504 4526
rect 523 4506 530 4526
rect 419 4489 530 4506
rect 910 4517 952 4598
rect 1240 4519 1273 4739
rect 1694 4737 1731 4739
rect 2324 4787 2372 4811
rect 2554 4805 2601 6382
rect 3088 6339 3122 6518
rect 3353 6535 3463 6550
rect 3353 6532 3430 6535
rect 3353 6505 3356 6532
rect 3385 6508 3430 6532
rect 3459 6508 3463 6535
rect 3385 6505 3463 6508
rect 3353 6491 3463 6505
rect 2697 6314 3122 6339
rect 3201 6378 3238 6380
rect 3659 6378 3692 6598
rect 3980 6519 4022 6600
rect 4402 6611 4513 6627
rect 4402 6591 4409 6611
rect 4428 6591 4486 6611
rect 4505 6591 4513 6611
rect 4402 6569 4513 6591
rect 3769 6517 3804 6518
rect 3201 6349 3692 6378
rect 2697 6298 3121 6314
rect 2697 5907 2735 6298
rect 3201 6283 3238 6349
rect 3659 6348 3692 6349
rect 3748 6510 3804 6517
rect 3748 6490 3777 6510
rect 3797 6490 3804 6510
rect 3748 6485 3804 6490
rect 3978 6515 4022 6519
rect 3978 6495 3989 6515
rect 4012 6495 4022 6515
rect 3978 6488 4022 6495
rect 4195 6513 4227 6520
rect 4195 6493 4201 6513
rect 4222 6493 4227 6513
rect 3978 6486 4021 6488
rect 3196 6274 3238 6283
rect 3196 6252 3205 6274
rect 3231 6252 3238 6274
rect 3463 6301 3574 6318
rect 3463 6281 3470 6301
rect 3489 6281 3547 6301
rect 3566 6281 3574 6301
rect 3463 6259 3574 6281
rect 3748 6279 3782 6485
rect 4195 6465 4227 6493
rect 3815 6457 4227 6465
rect 3815 6431 3821 6457
rect 3847 6431 4227 6457
rect 3815 6429 4227 6431
rect 3817 6428 3857 6429
rect 4195 6364 4227 6429
rect 4195 6344 4199 6364
rect 4220 6344 4227 6364
rect 4195 6337 4227 6344
rect 3748 6271 3783 6279
rect 3196 6242 3238 6252
rect 3748 6251 3756 6271
rect 3776 6251 3783 6271
rect 3748 6246 3783 6251
rect 4402 6266 4512 6281
rect 4402 6263 4479 6266
rect 3196 6241 3237 6242
rect 2830 6207 2865 6208
rect 2809 6200 2865 6207
rect 2809 6180 2838 6200
rect 2858 6180 2865 6200
rect 2809 6175 2865 6180
rect 3256 6203 3288 6210
rect 3256 6183 3262 6203
rect 3283 6183 3288 6203
rect 3748 6194 3782 6246
rect 4402 6236 4405 6263
rect 4434 6239 4479 6263
rect 4508 6239 4512 6266
rect 4434 6236 4512 6239
rect 4402 6222 4512 6236
rect 4698 6266 4740 6276
rect 4698 6247 4706 6266
rect 4731 6247 4740 6266
rect 4698 6194 4740 6247
rect 2809 5969 2843 6175
rect 3256 6155 3288 6183
rect 3746 6168 4742 6194
rect 2876 6147 3288 6155
rect 2876 6121 2882 6147
rect 2908 6121 3288 6147
rect 2876 6119 3288 6121
rect 2878 6118 2918 6119
rect 3038 6083 3077 6098
rect 3038 6042 3049 6083
rect 3070 6042 3077 6083
rect 2808 5961 2844 5969
rect 2808 5941 2817 5961
rect 2837 5941 2844 5961
rect 2808 5940 2844 5941
rect 2808 5929 2842 5940
rect 2698 5899 2735 5907
rect 2698 5865 2942 5899
rect 2690 5696 2725 5697
rect 2669 5689 2725 5696
rect 2669 5669 2698 5689
rect 2718 5669 2725 5689
rect 2669 5664 2725 5669
rect 2900 5694 2942 5865
rect 3038 5769 3077 6042
rect 3256 6054 3288 6119
rect 3256 6034 3260 6054
rect 3281 6034 3288 6054
rect 3256 6027 3288 6034
rect 3674 6061 3732 6062
rect 3674 6042 4011 6061
rect 4401 6057 4512 6074
rect 3674 6029 4012 6042
rect 3178 5965 3231 5968
rect 3178 5948 3190 5965
rect 3222 5948 3231 5965
rect 3178 5940 3231 5948
rect 3177 5893 3231 5940
rect 3463 5956 3573 5971
rect 3463 5953 3540 5956
rect 3463 5926 3466 5953
rect 3495 5929 3540 5953
rect 3569 5929 3573 5956
rect 3495 5926 3573 5929
rect 3463 5912 3573 5926
rect 3674 5893 3711 6029
rect 3980 6012 4012 6029
rect 4401 6037 4408 6057
rect 4427 6037 4485 6057
rect 4504 6037 4512 6057
rect 4401 6015 4512 6037
rect 3980 5966 4011 6012
rect 3768 5963 3803 5964
rect 3747 5956 3803 5963
rect 3747 5936 3776 5956
rect 3796 5936 3803 5956
rect 3747 5931 3803 5936
rect 3980 5959 4019 5966
rect 3980 5939 3986 5959
rect 4011 5939 4019 5959
rect 3980 5933 4019 5939
rect 4194 5959 4226 5966
rect 4194 5939 4200 5959
rect 4221 5939 4226 5959
rect 3177 5858 3712 5893
rect 3177 5854 3230 5858
rect 3038 5742 3042 5769
rect 3073 5742 3077 5769
rect 3323 5790 3434 5807
rect 3323 5770 3330 5790
rect 3349 5770 3407 5790
rect 3426 5770 3434 5790
rect 3323 5748 3434 5770
rect 3038 5735 3077 5742
rect 3747 5725 3781 5931
rect 4194 5911 4226 5939
rect 3814 5903 4226 5911
rect 3814 5877 3820 5903
rect 3846 5877 4226 5903
rect 3814 5875 4226 5877
rect 3816 5874 3856 5875
rect 4194 5810 4226 5875
rect 4194 5790 4198 5810
rect 4219 5790 4226 5810
rect 4194 5783 4226 5790
rect 4697 5825 4745 5830
rect 4697 5796 4708 5825
rect 4737 5796 4745 5825
rect 3747 5724 3782 5725
rect 3745 5717 3782 5724
rect 2900 5673 2908 5694
rect 2935 5673 2942 5694
rect 2669 5458 2703 5664
rect 2900 5662 2942 5673
rect 3116 5692 3148 5699
rect 3116 5672 3122 5692
rect 3143 5672 3148 5692
rect 3116 5644 3148 5672
rect 2736 5636 3148 5644
rect 2736 5610 2742 5636
rect 2768 5610 3148 5636
rect 3745 5697 3755 5717
rect 3775 5697 3782 5717
rect 3745 5692 3782 5697
rect 4401 5712 4511 5727
rect 4401 5709 4478 5712
rect 3745 5641 3780 5692
rect 4401 5682 4404 5709
rect 4433 5685 4478 5709
rect 4507 5685 4511 5712
rect 4433 5682 4511 5685
rect 4401 5668 4511 5682
rect 4697 5641 4745 5796
rect 3745 5617 4745 5641
rect 3745 5614 4744 5617
rect 3745 5612 3780 5614
rect 2736 5608 3148 5610
rect 2738 5607 2778 5608
rect 3116 5543 3148 5608
rect 3116 5523 3120 5543
rect 3141 5523 3148 5543
rect 3721 5526 4023 5528
rect 3116 5516 3148 5523
rect 3660 5497 4023 5526
rect 3660 5495 3721 5497
rect 2669 5450 2704 5458
rect 2669 5430 2677 5450
rect 2697 5430 2704 5450
rect 2669 5425 2704 5430
rect 3041 5451 3079 5457
rect 3041 5434 3051 5451
rect 3071 5434 3079 5451
rect 2669 5424 2701 5425
rect 2831 5104 2866 5105
rect 1468 4618 1578 4632
rect 1468 4615 1546 4618
rect 1468 4588 1472 4615
rect 1501 4591 1546 4615
rect 1575 4591 1578 4618
rect 2324 4609 2371 4787
rect 2554 4765 2567 4805
rect 2594 4765 2601 4805
rect 2810 5097 2866 5104
rect 2810 5077 2839 5097
rect 2859 5077 2866 5097
rect 2810 5072 2866 5077
rect 3041 5096 3079 5434
rect 3323 5445 3433 5460
rect 3323 5442 3400 5445
rect 3323 5415 3326 5442
rect 3355 5418 3400 5442
rect 3429 5418 3433 5445
rect 3355 5415 3433 5418
rect 3323 5401 3433 5415
rect 3202 5275 3239 5277
rect 3660 5275 3693 5495
rect 3981 5416 4023 5497
rect 4403 5508 4514 5525
rect 4403 5488 4410 5508
rect 4429 5488 4487 5508
rect 4506 5488 4514 5508
rect 4403 5466 4514 5488
rect 3770 5414 3805 5415
rect 3202 5246 3693 5275
rect 3202 5180 3239 5246
rect 3660 5245 3693 5246
rect 3749 5407 3805 5414
rect 3749 5387 3778 5407
rect 3798 5387 3805 5407
rect 3749 5382 3805 5387
rect 3979 5412 4023 5416
rect 3979 5392 3990 5412
rect 4013 5392 4023 5412
rect 3979 5385 4023 5392
rect 4196 5410 4228 5417
rect 4196 5390 4202 5410
rect 4223 5390 4228 5410
rect 3979 5383 4022 5385
rect 3197 5171 3239 5180
rect 3197 5149 3206 5171
rect 3232 5149 3239 5171
rect 3464 5198 3575 5215
rect 3464 5178 3471 5198
rect 3490 5178 3548 5198
rect 3567 5178 3575 5198
rect 3464 5156 3575 5178
rect 3749 5176 3783 5382
rect 4196 5362 4228 5390
rect 3816 5354 4228 5362
rect 3816 5328 3822 5354
rect 3848 5328 4228 5354
rect 3816 5326 4228 5328
rect 3818 5325 3858 5326
rect 4196 5261 4228 5326
rect 4196 5241 4200 5261
rect 4221 5241 4228 5261
rect 4196 5234 4228 5241
rect 3749 5168 3784 5176
rect 3197 5139 3239 5149
rect 3749 5148 3757 5168
rect 3777 5148 3784 5168
rect 3749 5143 3784 5148
rect 4403 5163 4513 5178
rect 4403 5160 4480 5163
rect 3197 5138 3238 5139
rect 3041 5079 3049 5096
rect 3069 5079 3079 5096
rect 2810 4866 2844 5072
rect 3041 5069 3079 5079
rect 3257 5100 3289 5107
rect 3257 5080 3263 5100
rect 3284 5080 3289 5100
rect 3749 5091 3783 5143
rect 4403 5133 4406 5160
rect 4435 5136 4480 5160
rect 4509 5136 4513 5163
rect 4435 5133 4513 5136
rect 4403 5119 4513 5133
rect 4699 5163 4741 5173
rect 4699 5144 4707 5163
rect 4732 5144 4741 5163
rect 4699 5091 4741 5144
rect 3257 5052 3289 5080
rect 3747 5065 4743 5091
rect 2877 5044 3289 5052
rect 2877 5018 2883 5044
rect 2909 5018 3289 5044
rect 2877 5016 3289 5018
rect 2879 5015 2919 5016
rect 3257 4951 3289 5016
rect 3257 4931 3261 4951
rect 3282 4931 3289 4951
rect 3257 4924 3289 4931
rect 3675 4958 3733 4959
rect 3675 4939 4012 4958
rect 4402 4954 4513 4971
rect 3675 4926 4013 4939
rect 2810 4858 2845 4866
rect 2810 4838 2818 4858
rect 2838 4838 2845 4858
rect 2810 4833 2845 4838
rect 3464 4853 3574 4868
rect 3464 4850 3541 4853
rect 2810 4790 2844 4833
rect 3464 4823 3467 4850
rect 3496 4826 3541 4850
rect 3570 4826 3574 4853
rect 3496 4823 3574 4826
rect 3464 4809 3574 4823
rect 3675 4790 3712 4926
rect 3981 4909 4013 4926
rect 4402 4934 4409 4954
rect 4428 4934 4486 4954
rect 4505 4934 4513 4954
rect 4402 4912 4513 4934
rect 3981 4863 4012 4909
rect 3769 4860 3804 4861
rect 3748 4853 3804 4860
rect 3748 4833 3777 4853
rect 3797 4833 3804 4853
rect 3748 4828 3804 4833
rect 3981 4856 4020 4863
rect 3981 4836 3987 4856
rect 4012 4836 4020 4856
rect 3981 4830 4020 4836
rect 4195 4856 4227 4863
rect 4195 4836 4201 4856
rect 4222 4836 4227 4856
rect 2554 4747 2601 4765
rect 2809 4755 3713 4790
rect 2810 4754 2844 4755
rect 2471 4688 2523 4693
rect 2926 4688 2971 4690
rect 2471 4673 2971 4688
rect 2471 4620 2485 4673
rect 2516 4649 2971 4673
rect 2516 4648 2541 4649
rect 2516 4620 2523 4648
rect 1501 4588 1578 4591
rect 1468 4573 1578 4588
rect 2193 4603 2374 4609
rect 2193 4583 2204 4603
rect 2224 4583 2374 4603
rect 2471 4596 2523 4620
rect 2193 4577 2374 4583
rect 2197 4575 2232 4577
rect 1212 4517 1273 4519
rect 910 4488 1273 4517
rect 1753 4510 1785 4517
rect 1753 4490 1760 4510
rect 1781 4490 1785 4510
rect 910 4486 1212 4488
rect 1753 4425 1785 4490
rect 2123 4425 2163 4426
rect 1753 4423 2165 4425
rect 1152 4400 1187 4402
rect 188 4397 1187 4400
rect 187 4373 1187 4397
rect 187 4218 235 4373
rect 421 4332 531 4346
rect 421 4329 499 4332
rect 421 4302 425 4329
rect 454 4305 499 4329
rect 528 4305 531 4332
rect 1152 4322 1187 4373
rect 1753 4397 2133 4423
rect 2159 4397 2165 4423
rect 1753 4389 2165 4397
rect 1753 4361 1785 4389
rect 2198 4369 2232 4575
rect 2722 4574 2757 4575
rect 1753 4341 1758 4361
rect 1779 4341 1785 4361
rect 1753 4334 1785 4341
rect 1955 4364 2000 4369
rect 1955 4340 1966 4364
rect 1992 4340 2000 4364
rect 1955 4329 2000 4340
rect 2176 4364 2232 4369
rect 2176 4344 2183 4364
rect 2203 4344 2232 4364
rect 2176 4337 2232 4344
rect 2701 4567 2757 4574
rect 2701 4547 2730 4567
rect 2750 4547 2757 4567
rect 2701 4542 2757 4547
rect 2926 4570 2971 4649
rect 3355 4668 3466 4685
rect 3355 4648 3362 4668
rect 3381 4648 3439 4668
rect 3458 4648 3466 4668
rect 3355 4626 3466 4648
rect 3748 4622 3782 4828
rect 4195 4808 4227 4836
rect 3815 4800 4227 4808
rect 3815 4774 3821 4800
rect 3847 4774 4227 4800
rect 3815 4772 4227 4774
rect 3817 4771 3857 4772
rect 4195 4707 4227 4772
rect 4195 4687 4199 4707
rect 4220 4687 4227 4707
rect 4195 4680 4227 4687
rect 4698 4722 4746 4727
rect 4698 4693 4709 4722
rect 4738 4693 4746 4722
rect 3748 4621 3783 4622
rect 3746 4614 3783 4621
rect 3746 4594 3756 4614
rect 3776 4594 3783 4614
rect 3746 4589 3783 4594
rect 4402 4609 4512 4624
rect 4402 4606 4479 4609
rect 2926 4550 2937 4570
rect 2962 4550 2971 4570
rect 2926 4546 2971 4550
rect 3148 4570 3180 4577
rect 3148 4550 3154 4570
rect 3175 4550 3180 4570
rect 2176 4336 2211 4337
rect 2701 4336 2735 4542
rect 3148 4522 3180 4550
rect 2768 4514 3180 4522
rect 2768 4488 2774 4514
rect 2800 4488 3180 4514
rect 3746 4538 3781 4589
rect 4402 4579 4405 4606
rect 4434 4582 4479 4606
rect 4508 4582 4512 4609
rect 4434 4579 4512 4582
rect 4402 4565 4512 4579
rect 4698 4538 4746 4693
rect 3746 4514 4746 4538
rect 3746 4511 4745 4514
rect 3746 4509 3781 4511
rect 2768 4486 3180 4488
rect 2770 4485 2810 4486
rect 3148 4421 3180 4486
rect 3721 4423 4023 4425
rect 3148 4401 3152 4421
rect 3173 4401 3180 4421
rect 3148 4394 3180 4401
rect 3660 4394 4023 4423
rect 3660 4392 3721 4394
rect 2701 4334 2736 4336
rect 454 4302 531 4305
rect 421 4287 531 4302
rect 1150 4317 1187 4322
rect 1150 4297 1157 4317
rect 1177 4297 1187 4317
rect 1150 4290 1187 4297
rect 1956 4295 1994 4329
rect 2559 4328 2740 4334
rect 2559 4308 2709 4328
rect 2729 4308 2740 4328
rect 2559 4302 2740 4308
rect 3355 4323 3465 4338
rect 3355 4320 3432 4323
rect 2392 4295 2442 4299
rect 1150 4289 1185 4290
rect 187 4189 195 4218
rect 224 4189 235 4218
rect 187 4184 235 4189
rect 706 4224 738 4231
rect 706 4204 713 4224
rect 734 4204 738 4224
rect 706 4139 738 4204
rect 1076 4139 1116 4140
rect 706 4137 1118 4139
rect 706 4111 1086 4137
rect 1112 4111 1118 4137
rect 706 4103 1118 4111
rect 706 4075 738 4103
rect 1151 4083 1185 4289
rect 1956 4285 2442 4295
rect 1467 4263 1578 4285
rect 1467 4243 1475 4263
rect 1494 4243 1552 4263
rect 1571 4243 1578 4263
rect 1956 4253 2405 4285
rect 1467 4226 1578 4243
rect 2392 4232 2405 4253
rect 2436 4232 2442 4285
rect 2392 4215 2442 4232
rect 2089 4156 2123 4157
rect 1220 4121 2124 4156
rect 2332 4146 2379 4164
rect 706 4055 711 4075
rect 732 4055 738 4075
rect 706 4048 738 4055
rect 913 4075 952 4081
rect 913 4055 921 4075
rect 946 4055 952 4075
rect 913 4048 952 4055
rect 1129 4078 1185 4083
rect 1129 4058 1136 4078
rect 1156 4058 1185 4078
rect 1129 4051 1185 4058
rect 1129 4050 1164 4051
rect 921 4002 952 4048
rect 420 3977 531 3999
rect 420 3957 428 3977
rect 447 3957 505 3977
rect 524 3957 531 3977
rect 920 3985 952 4002
rect 1221 3985 1258 4121
rect 1359 4088 1469 4102
rect 1359 4085 1437 4088
rect 1359 4058 1363 4085
rect 1392 4061 1437 4085
rect 1466 4061 1469 4088
rect 2089 4078 2123 4121
rect 1392 4058 1469 4061
rect 1359 4043 1469 4058
rect 2088 4073 2123 4078
rect 2088 4053 2095 4073
rect 2115 4053 2123 4073
rect 2088 4045 2123 4053
rect 920 3972 1258 3985
rect 420 3940 531 3957
rect 921 3953 1258 3972
rect 1200 3952 1258 3953
rect 1644 3980 1676 3987
rect 1644 3960 1651 3980
rect 1672 3960 1676 3980
rect 1644 3895 1676 3960
rect 2014 3895 2054 3896
rect 1644 3893 2056 3895
rect 1644 3867 2024 3893
rect 2050 3867 2056 3893
rect 1644 3859 2056 3867
rect 190 3820 1186 3846
rect 1644 3831 1676 3859
rect 192 3767 234 3820
rect 192 3748 201 3767
rect 226 3748 234 3767
rect 192 3738 234 3748
rect 420 3778 530 3792
rect 420 3775 498 3778
rect 420 3748 424 3775
rect 453 3751 498 3775
rect 527 3751 530 3778
rect 1150 3768 1184 3820
rect 1644 3811 1649 3831
rect 1670 3811 1676 3831
rect 1644 3804 1676 3811
rect 1854 3832 1892 3842
rect 2089 3839 2123 4045
rect 1854 3815 1864 3832
rect 1884 3815 1892 3832
rect 1695 3772 1736 3773
rect 453 3748 530 3751
rect 420 3733 530 3748
rect 1149 3763 1184 3768
rect 1149 3743 1156 3763
rect 1176 3743 1184 3763
rect 1694 3762 1736 3772
rect 1149 3735 1184 3743
rect 705 3670 737 3677
rect 705 3650 712 3670
rect 733 3650 737 3670
rect 705 3585 737 3650
rect 1075 3585 1115 3586
rect 705 3583 1117 3585
rect 705 3557 1085 3583
rect 1111 3557 1117 3583
rect 705 3549 1117 3557
rect 705 3521 737 3549
rect 1150 3529 1184 3735
rect 1358 3733 1469 3755
rect 1358 3713 1366 3733
rect 1385 3713 1443 3733
rect 1462 3713 1469 3733
rect 1358 3696 1469 3713
rect 1694 3740 1701 3762
rect 1727 3740 1736 3762
rect 1694 3731 1736 3740
rect 911 3526 954 3528
rect 705 3501 710 3521
rect 731 3501 737 3521
rect 705 3494 737 3501
rect 910 3519 954 3526
rect 910 3499 920 3519
rect 943 3499 954 3519
rect 910 3495 954 3499
rect 1128 3524 1184 3529
rect 1128 3504 1135 3524
rect 1155 3504 1184 3524
rect 1128 3497 1184 3504
rect 1240 3665 1273 3666
rect 1694 3665 1731 3731
rect 1240 3636 1731 3665
rect 1128 3496 1163 3497
rect 419 3423 530 3445
rect 419 3403 427 3423
rect 446 3403 504 3423
rect 523 3403 530 3423
rect 419 3386 530 3403
rect 910 3414 952 3495
rect 1240 3416 1273 3636
rect 1694 3634 1731 3636
rect 1500 3496 1610 3510
rect 1500 3493 1578 3496
rect 1500 3466 1504 3493
rect 1533 3469 1578 3493
rect 1607 3469 1610 3496
rect 1533 3466 1610 3469
rect 1500 3451 1610 3466
rect 1854 3477 1892 3815
rect 2067 3834 2123 3839
rect 2067 3814 2074 3834
rect 2094 3814 2123 3834
rect 2067 3807 2123 3814
rect 2332 4106 2339 4146
rect 2366 4106 2379 4146
rect 2562 4124 2609 4302
rect 3355 4293 3358 4320
rect 3387 4296 3432 4320
rect 3461 4296 3465 4323
rect 3387 4293 3465 4296
rect 3355 4279 3465 4293
rect 2067 3806 2102 3807
rect 2232 3486 2264 3487
rect 1854 3460 1862 3477
rect 1882 3460 1892 3477
rect 1854 3454 1892 3460
rect 2229 3481 2264 3486
rect 2229 3461 2236 3481
rect 2256 3461 2264 3481
rect 2229 3453 2264 3461
rect 1212 3414 1273 3416
rect 910 3385 1273 3414
rect 1785 3388 1817 3395
rect 910 3383 1212 3385
rect 1785 3368 1792 3388
rect 1813 3368 1817 3388
rect 1785 3303 1817 3368
rect 2155 3303 2195 3304
rect 1785 3301 2197 3303
rect 1153 3297 1188 3299
rect 189 3294 1188 3297
rect 188 3270 1188 3294
rect 188 3115 236 3270
rect 422 3229 532 3243
rect 422 3226 500 3229
rect 422 3199 426 3226
rect 455 3202 500 3226
rect 529 3202 532 3229
rect 1153 3219 1188 3270
rect 455 3199 532 3202
rect 422 3184 532 3199
rect 1151 3214 1188 3219
rect 1151 3194 1158 3214
rect 1178 3194 1188 3214
rect 1785 3275 2165 3301
rect 2191 3275 2197 3301
rect 1785 3267 2197 3275
rect 1785 3239 1817 3267
rect 1785 3219 1790 3239
rect 1811 3219 1817 3239
rect 1785 3212 1817 3219
rect 1991 3238 2033 3249
rect 2230 3247 2264 3453
rect 1991 3217 1998 3238
rect 2025 3217 2033 3238
rect 1151 3187 1188 3194
rect 1151 3186 1186 3187
rect 188 3086 196 3115
rect 225 3086 236 3115
rect 188 3081 236 3086
rect 707 3121 739 3128
rect 707 3101 714 3121
rect 735 3101 739 3121
rect 707 3036 739 3101
rect 1077 3036 1117 3037
rect 707 3034 1119 3036
rect 707 3008 1087 3034
rect 1113 3008 1119 3034
rect 707 3000 1119 3008
rect 707 2972 739 3000
rect 1152 2980 1186 3186
rect 1856 3169 1895 3176
rect 1499 3141 1610 3163
rect 1499 3121 1507 3141
rect 1526 3121 1584 3141
rect 1603 3121 1610 3141
rect 1499 3104 1610 3121
rect 1856 3142 1860 3169
rect 1891 3142 1895 3169
rect 1703 3053 1756 3057
rect 1221 3018 1756 3053
rect 707 2952 712 2972
rect 733 2952 739 2972
rect 707 2945 739 2952
rect 914 2972 953 2978
rect 914 2952 922 2972
rect 947 2952 953 2972
rect 914 2945 953 2952
rect 1130 2975 1186 2980
rect 1130 2955 1137 2975
rect 1157 2955 1186 2975
rect 1130 2948 1186 2955
rect 1130 2947 1165 2948
rect 922 2899 953 2945
rect 421 2874 532 2896
rect 421 2854 429 2874
rect 448 2854 506 2874
rect 525 2854 532 2874
rect 921 2882 953 2899
rect 1222 2882 1259 3018
rect 1360 2985 1470 2999
rect 1360 2982 1438 2985
rect 1360 2955 1364 2982
rect 1393 2958 1438 2982
rect 1467 2958 1470 2985
rect 1393 2955 1470 2958
rect 1360 2940 1470 2955
rect 1702 2971 1756 3018
rect 1702 2963 1755 2971
rect 1702 2946 1711 2963
rect 1743 2946 1755 2963
rect 1702 2943 1755 2946
rect 921 2869 1259 2882
rect 421 2837 532 2854
rect 922 2850 1259 2869
rect 1201 2849 1259 2850
rect 1645 2877 1677 2884
rect 1645 2857 1652 2877
rect 1673 2857 1677 2877
rect 1645 2792 1677 2857
rect 1856 2869 1895 3142
rect 1991 3046 2033 3217
rect 2208 3242 2264 3247
rect 2208 3222 2215 3242
rect 2235 3222 2264 3242
rect 2208 3215 2264 3222
rect 2208 3214 2243 3215
rect 1991 3012 2235 3046
rect 2198 3004 2235 3012
rect 2091 2971 2125 2982
rect 2089 2970 2125 2971
rect 2089 2950 2096 2970
rect 2116 2950 2125 2970
rect 2089 2942 2125 2950
rect 1856 2828 1863 2869
rect 1884 2828 1895 2869
rect 1856 2813 1895 2828
rect 2015 2792 2055 2793
rect 1645 2790 2057 2792
rect 1645 2764 2025 2790
rect 2051 2764 2057 2790
rect 1645 2756 2057 2764
rect 191 2717 1187 2743
rect 1645 2728 1677 2756
rect 2090 2736 2124 2942
rect 193 2664 235 2717
rect 193 2645 202 2664
rect 227 2645 235 2664
rect 193 2635 235 2645
rect 421 2675 531 2689
rect 421 2672 499 2675
rect 421 2645 425 2672
rect 454 2648 499 2672
rect 528 2648 531 2675
rect 1151 2665 1185 2717
rect 1645 2708 1650 2728
rect 1671 2708 1677 2728
rect 1645 2701 1677 2708
rect 2068 2731 2124 2736
rect 2068 2711 2075 2731
rect 2095 2711 2124 2731
rect 2068 2704 2124 2711
rect 2068 2703 2103 2704
rect 1696 2669 1737 2670
rect 454 2645 531 2648
rect 421 2630 531 2645
rect 1150 2660 1185 2665
rect 1150 2640 1157 2660
rect 1177 2640 1185 2660
rect 1695 2659 1737 2669
rect 1150 2632 1185 2640
rect 706 2567 738 2574
rect 706 2547 713 2567
rect 734 2547 738 2567
rect 706 2482 738 2547
rect 1076 2482 1116 2483
rect 706 2480 1118 2482
rect 706 2454 1086 2480
rect 1112 2454 1118 2480
rect 706 2446 1118 2454
rect 706 2418 738 2446
rect 1151 2426 1185 2632
rect 1359 2630 1470 2652
rect 1359 2610 1367 2630
rect 1386 2610 1444 2630
rect 1463 2610 1470 2630
rect 1359 2593 1470 2610
rect 1695 2637 1702 2659
rect 1728 2637 1737 2659
rect 1695 2628 1737 2637
rect 912 2423 955 2425
rect 706 2398 711 2418
rect 732 2398 738 2418
rect 706 2391 738 2398
rect 911 2416 955 2423
rect 911 2396 921 2416
rect 944 2396 955 2416
rect 911 2392 955 2396
rect 1129 2421 1185 2426
rect 1129 2401 1136 2421
rect 1156 2401 1185 2421
rect 1129 2394 1185 2401
rect 1241 2562 1274 2563
rect 1695 2562 1732 2628
rect 2198 2613 2236 3004
rect 1812 2597 2236 2613
rect 1241 2533 1732 2562
rect 1129 2393 1164 2394
rect 420 2320 531 2342
rect 420 2300 428 2320
rect 447 2300 505 2320
rect 524 2300 531 2320
rect 420 2284 531 2300
rect 911 2311 953 2392
rect 1241 2313 1274 2533
rect 1695 2531 1732 2533
rect 1811 2572 2236 2597
rect 1470 2406 1580 2420
rect 1470 2403 1548 2406
rect 1470 2376 1474 2403
rect 1503 2379 1548 2403
rect 1577 2379 1580 2406
rect 1503 2376 1580 2379
rect 1470 2361 1580 2376
rect 1811 2393 1845 2572
rect 2332 2529 2379 4106
rect 2561 4100 2609 4124
rect 3202 4172 3239 4174
rect 3660 4172 3693 4392
rect 3981 4313 4023 4394
rect 4403 4405 4514 4422
rect 4403 4385 4410 4405
rect 4429 4385 4487 4405
rect 4506 4385 4514 4405
rect 4403 4363 4514 4385
rect 3770 4311 3805 4312
rect 3202 4143 3693 4172
rect 2561 2615 2607 4100
rect 3202 4077 3239 4143
rect 3660 4142 3693 4143
rect 3749 4304 3805 4311
rect 3749 4284 3778 4304
rect 3798 4284 3805 4304
rect 3749 4279 3805 4284
rect 3979 4309 4023 4313
rect 3979 4289 3990 4309
rect 4013 4289 4023 4309
rect 3979 4282 4023 4289
rect 4196 4307 4228 4314
rect 4196 4287 4202 4307
rect 4223 4287 4228 4307
rect 3979 4280 4022 4282
rect 3197 4068 3239 4077
rect 3197 4046 3206 4068
rect 3232 4046 3239 4068
rect 3464 4095 3575 4112
rect 3464 4075 3471 4095
rect 3490 4075 3548 4095
rect 3567 4075 3575 4095
rect 3464 4053 3575 4075
rect 3749 4073 3783 4279
rect 4196 4259 4228 4287
rect 3816 4251 4228 4259
rect 3816 4225 3822 4251
rect 3848 4225 4228 4251
rect 3816 4223 4228 4225
rect 3818 4222 3858 4223
rect 4196 4158 4228 4223
rect 4196 4138 4200 4158
rect 4221 4138 4228 4158
rect 4196 4131 4228 4138
rect 3749 4065 3784 4073
rect 3197 4036 3239 4046
rect 3749 4045 3757 4065
rect 3777 4045 3784 4065
rect 3749 4040 3784 4045
rect 4403 4060 4513 4075
rect 4403 4057 4480 4060
rect 3197 4035 3238 4036
rect 2831 4001 2866 4002
rect 2810 3994 2866 4001
rect 2810 3974 2839 3994
rect 2859 3974 2866 3994
rect 2810 3969 2866 3974
rect 3257 3997 3289 4004
rect 3257 3977 3263 3997
rect 3284 3977 3289 3997
rect 3749 3988 3783 4040
rect 4403 4030 4406 4057
rect 4435 4033 4480 4057
rect 4509 4033 4513 4060
rect 4435 4030 4513 4033
rect 4403 4016 4513 4030
rect 4699 4060 4741 4070
rect 4699 4041 4707 4060
rect 4732 4041 4741 4060
rect 4699 3988 4741 4041
rect 2810 3763 2844 3969
rect 3257 3949 3289 3977
rect 3747 3962 4743 3988
rect 2877 3941 3289 3949
rect 2877 3915 2883 3941
rect 2909 3915 3289 3941
rect 2877 3913 3289 3915
rect 2879 3912 2919 3913
rect 3039 3877 3078 3892
rect 3039 3836 3050 3877
rect 3071 3836 3078 3877
rect 2809 3755 2845 3763
rect 2809 3735 2818 3755
rect 2838 3735 2845 3755
rect 2809 3734 2845 3735
rect 2809 3723 2843 3734
rect 3039 3563 3078 3836
rect 3257 3848 3289 3913
rect 3257 3828 3261 3848
rect 3282 3828 3289 3848
rect 3257 3821 3289 3828
rect 3675 3855 3733 3856
rect 3675 3836 4012 3855
rect 4402 3851 4513 3868
rect 3675 3823 4013 3836
rect 3179 3759 3232 3762
rect 3179 3742 3191 3759
rect 3223 3742 3232 3759
rect 3179 3734 3232 3742
rect 3178 3687 3232 3734
rect 3464 3750 3574 3765
rect 3464 3747 3541 3750
rect 3464 3720 3467 3747
rect 3496 3723 3541 3747
rect 3570 3723 3574 3750
rect 3496 3720 3574 3723
rect 3464 3706 3574 3720
rect 3675 3687 3712 3823
rect 3981 3806 4013 3823
rect 4402 3831 4409 3851
rect 4428 3831 4486 3851
rect 4505 3831 4513 3851
rect 4402 3809 4513 3831
rect 3981 3760 4012 3806
rect 3769 3757 3804 3758
rect 3748 3750 3804 3757
rect 3748 3730 3777 3750
rect 3797 3730 3804 3750
rect 3748 3725 3804 3730
rect 3981 3753 4020 3760
rect 3981 3733 3987 3753
rect 4012 3733 4020 3753
rect 3981 3727 4020 3733
rect 4195 3753 4227 3760
rect 4195 3733 4201 3753
rect 4222 3733 4227 3753
rect 3178 3652 3713 3687
rect 3178 3648 3231 3652
rect 3039 3536 3043 3563
rect 3074 3536 3078 3563
rect 3324 3584 3435 3601
rect 3324 3564 3331 3584
rect 3350 3564 3408 3584
rect 3427 3564 3435 3584
rect 3324 3542 3435 3564
rect 3039 3529 3078 3536
rect 3748 3519 3782 3725
rect 4195 3705 4227 3733
rect 3815 3697 4227 3705
rect 3815 3671 3821 3697
rect 3847 3671 4227 3697
rect 3815 3669 4227 3671
rect 3817 3668 3857 3669
rect 4195 3604 4227 3669
rect 4195 3584 4199 3604
rect 4220 3584 4227 3604
rect 4195 3577 4227 3584
rect 4698 3619 4746 3624
rect 4698 3590 4709 3619
rect 4738 3590 4746 3619
rect 3748 3518 3783 3519
rect 3746 3511 3783 3518
rect 2691 3490 2726 3491
rect 2668 3483 2726 3490
rect 2668 3463 2699 3483
rect 2719 3463 2726 3483
rect 2668 3458 2726 3463
rect 3117 3486 3149 3493
rect 3117 3466 3123 3486
rect 3144 3466 3149 3486
rect 2668 3310 2704 3458
rect 3117 3438 3149 3466
rect 2737 3430 3149 3438
rect 2737 3404 2743 3430
rect 2769 3404 3149 3430
rect 3746 3491 3756 3511
rect 3776 3491 3783 3511
rect 3746 3486 3783 3491
rect 4402 3506 4512 3521
rect 4402 3503 4479 3506
rect 3746 3435 3781 3486
rect 4402 3476 4405 3503
rect 4434 3479 4479 3503
rect 4508 3479 4512 3506
rect 4434 3476 4512 3479
rect 4402 3462 4512 3476
rect 4698 3435 4746 3590
rect 3746 3411 4746 3435
rect 3746 3408 4745 3411
rect 3746 3406 3781 3408
rect 2737 3402 3149 3404
rect 2739 3401 2779 3402
rect 2671 3252 2704 3310
rect 2901 3362 2939 3372
rect 2901 3324 2910 3362
rect 2933 3324 2939 3362
rect 2671 3244 2705 3252
rect 2671 3224 2678 3244
rect 2698 3224 2705 3244
rect 2671 3219 2705 3224
rect 2671 3218 2702 3219
rect 2901 3188 2939 3324
rect 3117 3337 3149 3402
rect 3117 3317 3121 3337
rect 3142 3317 3149 3337
rect 3722 3320 4024 3322
rect 3117 3310 3149 3317
rect 3661 3291 4024 3320
rect 3661 3289 3722 3291
rect 3042 3245 3080 3251
rect 3042 3228 3052 3245
rect 3072 3228 3080 3245
rect 2901 3034 2945 3188
rect 2738 3032 2945 3034
rect 2714 2999 2945 3032
rect 1811 2373 1815 2393
rect 1836 2373 1845 2393
rect 1811 2367 1845 2373
rect 1964 2504 2293 2507
rect 2332 2504 2376 2529
rect 1964 2474 2376 2504
rect 1213 2311 1274 2313
rect 911 2282 1274 2311
rect 1755 2298 1787 2305
rect 911 2280 1213 2282
rect 1755 2278 1762 2298
rect 1783 2278 1787 2298
rect 1755 2213 1787 2278
rect 1964 2286 1999 2474
rect 2266 2472 2376 2474
rect 2559 2487 2609 2615
rect 2714 2598 2764 2999
rect 2901 2995 2945 2999
rect 2832 2898 2867 2899
rect 2694 2589 2764 2598
rect 2694 2560 2709 2589
rect 2757 2581 2764 2589
rect 2811 2891 2867 2898
rect 2811 2871 2840 2891
rect 2860 2871 2867 2891
rect 2811 2866 2867 2871
rect 3042 2890 3080 3228
rect 3324 3239 3434 3254
rect 3324 3236 3401 3239
rect 3324 3209 3327 3236
rect 3356 3212 3401 3236
rect 3430 3212 3434 3239
rect 3356 3209 3434 3212
rect 3324 3195 3434 3209
rect 3203 3069 3240 3071
rect 3661 3069 3694 3289
rect 3982 3210 4024 3291
rect 4404 3302 4515 3319
rect 4404 3282 4411 3302
rect 4430 3282 4488 3302
rect 4507 3282 4515 3302
rect 4404 3260 4515 3282
rect 3771 3208 3806 3209
rect 3203 3040 3694 3069
rect 3203 2974 3240 3040
rect 3661 3039 3694 3040
rect 3750 3201 3806 3208
rect 3750 3181 3779 3201
rect 3799 3181 3806 3201
rect 3750 3176 3806 3181
rect 3980 3206 4024 3210
rect 3980 3186 3991 3206
rect 4014 3186 4024 3206
rect 3980 3179 4024 3186
rect 4197 3204 4229 3211
rect 4197 3184 4203 3204
rect 4224 3184 4229 3204
rect 3980 3177 4023 3179
rect 3198 2965 3240 2974
rect 3198 2943 3207 2965
rect 3233 2943 3240 2965
rect 3465 2992 3576 3009
rect 3465 2972 3472 2992
rect 3491 2972 3549 2992
rect 3568 2972 3576 2992
rect 3465 2950 3576 2972
rect 3750 2970 3784 3176
rect 4197 3156 4229 3184
rect 3817 3148 4229 3156
rect 3817 3122 3823 3148
rect 3849 3122 4229 3148
rect 3817 3120 4229 3122
rect 3819 3119 3859 3120
rect 4197 3055 4229 3120
rect 4197 3035 4201 3055
rect 4222 3035 4229 3055
rect 4197 3028 4229 3035
rect 3750 2962 3785 2970
rect 3198 2933 3240 2943
rect 3750 2942 3758 2962
rect 3778 2942 3785 2962
rect 3750 2937 3785 2942
rect 4404 2957 4514 2972
rect 4404 2954 4481 2957
rect 3198 2932 3239 2933
rect 3042 2873 3050 2890
rect 3070 2873 3080 2890
rect 2811 2660 2845 2866
rect 3042 2863 3080 2873
rect 3258 2894 3290 2901
rect 3258 2874 3264 2894
rect 3285 2874 3290 2894
rect 3750 2885 3784 2937
rect 4404 2927 4407 2954
rect 4436 2930 4481 2954
rect 4510 2930 4514 2957
rect 4436 2927 4514 2930
rect 4404 2913 4514 2927
rect 4700 2957 4742 2967
rect 4700 2938 4708 2957
rect 4733 2938 4742 2957
rect 4700 2885 4742 2938
rect 3258 2846 3290 2874
rect 3748 2859 4744 2885
rect 2878 2838 3290 2846
rect 2878 2812 2884 2838
rect 2910 2812 3290 2838
rect 2878 2810 3290 2812
rect 2880 2809 2920 2810
rect 3258 2745 3290 2810
rect 3258 2725 3262 2745
rect 3283 2725 3290 2745
rect 3258 2718 3290 2725
rect 3676 2752 3734 2753
rect 3676 2733 4013 2752
rect 4403 2748 4514 2765
rect 3676 2720 4014 2733
rect 2811 2652 2846 2660
rect 2811 2632 2819 2652
rect 2839 2632 2846 2652
rect 2811 2627 2846 2632
rect 3465 2647 3575 2662
rect 3465 2644 3542 2647
rect 2811 2584 2845 2627
rect 3465 2617 3468 2644
rect 3497 2620 3542 2644
rect 3571 2620 3575 2647
rect 3497 2617 3575 2620
rect 3465 2603 3575 2617
rect 3676 2584 3713 2720
rect 3982 2703 4014 2720
rect 4403 2728 4410 2748
rect 4429 2728 4487 2748
rect 4506 2728 4514 2748
rect 4403 2706 4514 2728
rect 3982 2657 4013 2703
rect 3770 2654 3805 2655
rect 3749 2647 3805 2654
rect 3749 2627 3778 2647
rect 3798 2627 3805 2647
rect 3749 2622 3805 2627
rect 3982 2650 4021 2657
rect 3982 2630 3988 2650
rect 4013 2630 4021 2650
rect 3982 2624 4021 2630
rect 4196 2650 4228 2657
rect 4196 2630 4202 2650
rect 4223 2630 4228 2650
rect 2757 2560 2762 2581
rect 2694 2549 2762 2560
rect 2810 2549 3714 2584
rect 2811 2548 2845 2549
rect 2559 2453 2974 2487
rect 2559 2451 2609 2453
rect 2192 2389 2242 2396
rect 2192 2375 2206 2389
rect 2198 2371 2206 2375
rect 2226 2375 2242 2389
rect 2226 2371 2236 2375
rect 2722 2374 2757 2375
rect 2198 2364 2236 2371
rect 2701 2367 2757 2374
rect 2199 2363 2234 2364
rect 1964 2254 1969 2286
rect 1996 2254 1999 2286
rect 1964 2236 1999 2254
rect 2125 2213 2165 2214
rect 1755 2211 2167 2213
rect 1153 2194 1188 2196
rect 189 2191 1188 2194
rect 188 2167 1188 2191
rect 188 2012 236 2167
rect 422 2126 532 2140
rect 422 2123 500 2126
rect 422 2096 426 2123
rect 455 2099 500 2123
rect 529 2099 532 2126
rect 1153 2116 1188 2167
rect 1755 2185 2135 2211
rect 2161 2185 2167 2211
rect 1755 2177 2167 2185
rect 1755 2149 1787 2177
rect 2200 2157 2234 2363
rect 1755 2129 1760 2149
rect 1781 2129 1787 2149
rect 1755 2122 1787 2129
rect 2178 2152 2234 2157
rect 2178 2132 2185 2152
rect 2205 2132 2234 2152
rect 2701 2347 2730 2367
rect 2750 2347 2757 2367
rect 2701 2342 2757 2347
rect 2929 2370 2974 2453
rect 3355 2468 3466 2485
rect 3355 2448 3362 2468
rect 3381 2448 3439 2468
rect 3458 2448 3466 2468
rect 3355 2426 3466 2448
rect 3749 2416 3783 2622
rect 4196 2602 4228 2630
rect 3816 2594 4228 2602
rect 3816 2568 3822 2594
rect 3848 2568 4228 2594
rect 3816 2566 4228 2568
rect 3818 2565 3858 2566
rect 4196 2501 4228 2566
rect 4196 2481 4200 2501
rect 4221 2481 4228 2501
rect 4196 2474 4228 2481
rect 4699 2516 4747 2521
rect 4699 2487 4710 2516
rect 4739 2487 4747 2516
rect 3749 2415 3784 2416
rect 3747 2408 3784 2415
rect 3747 2388 3757 2408
rect 3777 2388 3784 2408
rect 3747 2383 3784 2388
rect 4403 2403 4513 2418
rect 4403 2400 4480 2403
rect 2929 2351 2938 2370
rect 2967 2351 2974 2370
rect 2701 2136 2735 2342
rect 2929 2339 2974 2351
rect 3148 2370 3180 2377
rect 3148 2350 3154 2370
rect 3175 2350 3180 2370
rect 3148 2322 3180 2350
rect 2768 2314 3180 2322
rect 2768 2288 2774 2314
rect 2800 2288 3180 2314
rect 3747 2332 3782 2383
rect 4403 2373 4406 2400
rect 4435 2376 4480 2400
rect 4509 2376 4513 2403
rect 4435 2373 4513 2376
rect 4403 2359 4513 2373
rect 4699 2332 4747 2487
rect 3747 2308 4747 2332
rect 3747 2305 4746 2308
rect 3747 2303 3782 2305
rect 2768 2286 3180 2288
rect 2770 2285 2810 2286
rect 3148 2221 3180 2286
rect 3148 2201 3152 2221
rect 3173 2201 3180 2221
rect 3722 2217 4024 2219
rect 3148 2194 3180 2201
rect 3661 2188 4024 2217
rect 3661 2186 3722 2188
rect 2701 2135 2736 2136
rect 2178 2125 2234 2132
rect 2699 2128 2737 2135
rect 2178 2124 2213 2125
rect 455 2096 532 2099
rect 422 2081 532 2096
rect 1151 2111 1188 2116
rect 1151 2091 1158 2111
rect 1178 2091 1188 2111
rect 2699 2108 2709 2128
rect 2729 2108 2737 2128
rect 1151 2084 1188 2091
rect 2173 2086 2243 2096
rect 1151 2083 1186 2084
rect 188 1983 196 2012
rect 225 1983 236 2012
rect 188 1978 236 1983
rect 707 2018 739 2025
rect 707 1998 714 2018
rect 735 1998 739 2018
rect 707 1933 739 1998
rect 1077 1933 1117 1934
rect 707 1931 1119 1933
rect 707 1905 1087 1931
rect 1113 1905 1119 1931
rect 707 1897 1119 1905
rect 707 1869 739 1897
rect 1152 1877 1186 2083
rect 2171 2079 2243 2086
rect 1469 2051 1580 2073
rect 1469 2031 1477 2051
rect 1496 2031 1554 2051
rect 1573 2031 1580 2051
rect 1469 2014 1580 2031
rect 2171 2050 2178 2079
rect 2226 2050 2243 2079
rect 2171 2041 2243 2050
rect 2090 1950 2124 1951
rect 1221 1915 2125 1950
rect 707 1849 712 1869
rect 733 1849 739 1869
rect 707 1842 739 1849
rect 914 1869 953 1875
rect 914 1849 922 1869
rect 947 1849 953 1869
rect 914 1842 953 1849
rect 1130 1872 1186 1877
rect 1130 1852 1137 1872
rect 1157 1852 1186 1872
rect 1130 1845 1186 1852
rect 1130 1844 1165 1845
rect 922 1796 953 1842
rect 421 1771 532 1793
rect 421 1751 429 1771
rect 448 1751 506 1771
rect 525 1751 532 1771
rect 921 1779 953 1796
rect 1222 1779 1259 1915
rect 1360 1882 1470 1896
rect 1360 1879 1438 1882
rect 1360 1852 1364 1879
rect 1393 1855 1438 1879
rect 1467 1855 1470 1882
rect 2090 1872 2124 1915
rect 1393 1852 1470 1855
rect 1360 1837 1470 1852
rect 2089 1867 2124 1872
rect 2089 1847 2096 1867
rect 2116 1847 2124 1867
rect 2089 1839 2124 1847
rect 921 1766 1259 1779
rect 421 1734 532 1751
rect 922 1747 1259 1766
rect 1201 1746 1259 1747
rect 1645 1774 1677 1781
rect 1645 1754 1652 1774
rect 1673 1754 1677 1774
rect 1645 1689 1677 1754
rect 2015 1689 2055 1690
rect 1645 1687 2057 1689
rect 1645 1661 2025 1687
rect 2051 1661 2057 1687
rect 1645 1653 2057 1661
rect 191 1614 1187 1640
rect 1645 1625 1677 1653
rect 193 1561 235 1614
rect 193 1542 202 1561
rect 227 1542 235 1561
rect 193 1532 235 1542
rect 421 1572 531 1586
rect 421 1569 499 1572
rect 421 1542 425 1569
rect 454 1545 499 1569
rect 528 1545 531 1572
rect 1151 1562 1185 1614
rect 1645 1605 1650 1625
rect 1671 1605 1677 1625
rect 1645 1598 1677 1605
rect 1855 1626 1893 1636
rect 2090 1633 2124 1839
rect 1855 1609 1865 1626
rect 1885 1609 1893 1626
rect 1696 1566 1737 1567
rect 454 1542 531 1545
rect 421 1527 531 1542
rect 1150 1557 1185 1562
rect 1150 1537 1157 1557
rect 1177 1537 1185 1557
rect 1695 1556 1737 1566
rect 1150 1529 1185 1537
rect 706 1464 738 1471
rect 706 1444 713 1464
rect 734 1444 738 1464
rect 706 1379 738 1444
rect 1076 1379 1116 1380
rect 706 1377 1118 1379
rect 706 1351 1086 1377
rect 1112 1351 1118 1377
rect 706 1343 1118 1351
rect 706 1315 738 1343
rect 1151 1323 1185 1529
rect 1359 1527 1470 1549
rect 1359 1507 1367 1527
rect 1386 1507 1444 1527
rect 1463 1507 1470 1527
rect 1359 1490 1470 1507
rect 1695 1534 1702 1556
rect 1728 1534 1737 1556
rect 1695 1525 1737 1534
rect 912 1320 955 1322
rect 706 1295 711 1315
rect 732 1295 738 1315
rect 706 1288 738 1295
rect 911 1313 955 1320
rect 911 1293 921 1313
rect 944 1293 955 1313
rect 911 1289 955 1293
rect 1129 1318 1185 1323
rect 1129 1298 1136 1318
rect 1156 1298 1185 1318
rect 1129 1291 1185 1298
rect 1241 1459 1274 1460
rect 1695 1459 1732 1525
rect 1241 1430 1732 1459
rect 1129 1290 1164 1291
rect 420 1217 531 1239
rect 420 1197 428 1217
rect 447 1197 505 1217
rect 524 1197 531 1217
rect 420 1180 531 1197
rect 911 1208 953 1289
rect 1241 1210 1274 1430
rect 1695 1428 1732 1430
rect 1501 1290 1611 1304
rect 1501 1287 1579 1290
rect 1501 1260 1505 1287
rect 1534 1263 1579 1287
rect 1608 1263 1611 1290
rect 1534 1260 1611 1263
rect 1501 1245 1611 1260
rect 1855 1271 1893 1609
rect 2068 1628 2124 1633
rect 2068 1608 2075 1628
rect 2095 1608 2124 1628
rect 2068 1601 2124 1608
rect 2068 1600 2103 1601
rect 1990 1500 2034 1504
rect 2171 1500 2221 2041
rect 1990 1467 2221 1500
rect 2699 1495 2737 2108
rect 3355 2123 3465 2138
rect 3355 2120 3432 2123
rect 3355 2093 3358 2120
rect 3387 2096 3432 2120
rect 3461 2096 3465 2123
rect 3387 2093 3465 2096
rect 3355 2079 3465 2093
rect 3203 1966 3240 1968
rect 3661 1966 3694 2186
rect 3982 2107 4024 2188
rect 4404 2199 4515 2215
rect 4404 2179 4411 2199
rect 4430 2179 4488 2199
rect 4507 2179 4515 2199
rect 4404 2157 4515 2179
rect 3771 2105 3806 2106
rect 3203 1937 3694 1966
rect 3203 1871 3240 1937
rect 3661 1936 3694 1937
rect 3750 2098 3806 2105
rect 3750 2078 3779 2098
rect 3799 2078 3806 2098
rect 3750 2073 3806 2078
rect 3980 2103 4024 2107
rect 3980 2083 3991 2103
rect 4014 2083 4024 2103
rect 3980 2076 4024 2083
rect 4197 2101 4229 2108
rect 4197 2081 4203 2101
rect 4224 2081 4229 2101
rect 3980 2074 4023 2076
rect 3198 1862 3240 1871
rect 3198 1840 3207 1862
rect 3233 1840 3240 1862
rect 3465 1889 3576 1906
rect 3465 1869 3472 1889
rect 3491 1869 3549 1889
rect 3568 1869 3576 1889
rect 3465 1847 3576 1869
rect 3750 1867 3784 2073
rect 4197 2053 4229 2081
rect 3817 2045 4229 2053
rect 3817 2019 3823 2045
rect 3849 2019 4229 2045
rect 3817 2017 4229 2019
rect 3819 2016 3859 2017
rect 4197 1952 4229 2017
rect 4197 1932 4201 1952
rect 4222 1932 4229 1952
rect 4197 1925 4229 1932
rect 3750 1859 3785 1867
rect 3198 1830 3240 1840
rect 3750 1839 3758 1859
rect 3778 1839 3785 1859
rect 3750 1834 3785 1839
rect 4404 1854 4514 1869
rect 4404 1851 4481 1854
rect 3198 1829 3239 1830
rect 2832 1795 2867 1796
rect 2811 1788 2867 1795
rect 2811 1768 2840 1788
rect 2860 1768 2867 1788
rect 2811 1763 2867 1768
rect 3258 1791 3290 1798
rect 3258 1771 3264 1791
rect 3285 1771 3290 1791
rect 3750 1782 3784 1834
rect 4404 1824 4407 1851
rect 4436 1827 4481 1851
rect 4510 1827 4514 1854
rect 4436 1824 4514 1827
rect 4404 1810 4514 1824
rect 4700 1854 4742 1864
rect 4700 1835 4708 1854
rect 4733 1835 4742 1854
rect 4700 1782 4742 1835
rect 2811 1557 2845 1763
rect 3258 1743 3290 1771
rect 3748 1756 4744 1782
rect 2878 1735 3290 1743
rect 2878 1709 2884 1735
rect 2910 1709 3290 1735
rect 2878 1707 3290 1709
rect 2880 1706 2920 1707
rect 3040 1671 3079 1686
rect 3040 1630 3051 1671
rect 3072 1630 3079 1671
rect 2810 1549 2846 1557
rect 2810 1529 2819 1549
rect 2839 1529 2846 1549
rect 2810 1528 2846 1529
rect 2810 1517 2844 1528
rect 2700 1487 2737 1495
rect 1990 1465 2197 1467
rect 1990 1311 2034 1465
rect 2700 1453 2944 1487
rect 1855 1254 1863 1271
rect 1883 1254 1893 1271
rect 1855 1248 1893 1254
rect 1213 1208 1274 1210
rect 911 1179 1274 1208
rect 1786 1182 1818 1189
rect 911 1177 1213 1179
rect 1786 1162 1793 1182
rect 1814 1162 1818 1182
rect 1786 1097 1818 1162
rect 1996 1175 2034 1311
rect 2692 1284 2727 1285
rect 2233 1280 2264 1281
rect 2230 1275 2264 1280
rect 2230 1255 2237 1275
rect 2257 1255 2264 1275
rect 2230 1247 2264 1255
rect 1996 1137 2002 1175
rect 2025 1137 2034 1175
rect 1996 1127 2034 1137
rect 2231 1189 2264 1247
rect 2671 1277 2727 1284
rect 2671 1257 2700 1277
rect 2720 1257 2727 1277
rect 2671 1252 2727 1257
rect 2902 1282 2944 1453
rect 3040 1357 3079 1630
rect 3258 1642 3290 1707
rect 3258 1622 3262 1642
rect 3283 1622 3290 1642
rect 3258 1615 3290 1622
rect 3676 1649 3734 1650
rect 3676 1630 4013 1649
rect 4403 1645 4514 1662
rect 3676 1617 4014 1630
rect 3180 1553 3233 1556
rect 3180 1536 3192 1553
rect 3224 1536 3233 1553
rect 3180 1528 3233 1536
rect 3179 1481 3233 1528
rect 3465 1544 3575 1559
rect 3465 1541 3542 1544
rect 3465 1514 3468 1541
rect 3497 1517 3542 1541
rect 3571 1517 3575 1544
rect 3497 1514 3575 1517
rect 3465 1500 3575 1514
rect 3676 1481 3713 1617
rect 3982 1600 4014 1617
rect 4403 1625 4410 1645
rect 4429 1625 4487 1645
rect 4506 1625 4514 1645
rect 4403 1603 4514 1625
rect 3982 1554 4013 1600
rect 3770 1551 3805 1552
rect 3749 1544 3805 1551
rect 3749 1524 3778 1544
rect 3798 1524 3805 1544
rect 3749 1519 3805 1524
rect 3982 1547 4021 1554
rect 3982 1527 3988 1547
rect 4013 1527 4021 1547
rect 3982 1521 4021 1527
rect 4196 1547 4228 1554
rect 4196 1527 4202 1547
rect 4223 1527 4228 1547
rect 3179 1446 3714 1481
rect 3179 1442 3232 1446
rect 3040 1330 3044 1357
rect 3075 1330 3079 1357
rect 3325 1378 3436 1395
rect 3325 1358 3332 1378
rect 3351 1358 3409 1378
rect 3428 1358 3436 1378
rect 3325 1336 3436 1358
rect 3040 1323 3079 1330
rect 3749 1313 3783 1519
rect 4196 1499 4228 1527
rect 3816 1491 4228 1499
rect 3816 1465 3822 1491
rect 3848 1465 4228 1491
rect 3816 1463 4228 1465
rect 3818 1462 3858 1463
rect 4196 1398 4228 1463
rect 4196 1378 4200 1398
rect 4221 1378 4228 1398
rect 4196 1371 4228 1378
rect 4699 1413 4747 1418
rect 4699 1384 4710 1413
rect 4739 1384 4747 1413
rect 3749 1312 3784 1313
rect 3747 1305 3784 1312
rect 2902 1261 2910 1282
rect 2937 1261 2944 1282
rect 2156 1097 2196 1098
rect 1786 1095 2198 1097
rect 1154 1091 1189 1093
rect 190 1088 1189 1091
rect 189 1064 1189 1088
rect 189 909 237 1064
rect 423 1023 533 1037
rect 423 1020 501 1023
rect 423 993 427 1020
rect 456 996 501 1020
rect 530 996 533 1023
rect 1154 1013 1189 1064
rect 456 993 533 996
rect 423 978 533 993
rect 1152 1008 1189 1013
rect 1152 988 1159 1008
rect 1179 988 1189 1008
rect 1786 1069 2166 1095
rect 2192 1069 2198 1095
rect 1786 1061 2198 1069
rect 1786 1033 1818 1061
rect 2231 1041 2267 1189
rect 1786 1013 1791 1033
rect 1812 1013 1818 1033
rect 1786 1006 1818 1013
rect 2209 1036 2267 1041
rect 2209 1016 2216 1036
rect 2236 1016 2267 1036
rect 2209 1009 2267 1016
rect 2671 1046 2705 1252
rect 2902 1250 2944 1261
rect 3118 1280 3150 1287
rect 3118 1260 3124 1280
rect 3145 1260 3150 1280
rect 3118 1232 3150 1260
rect 2738 1224 3150 1232
rect 2738 1198 2744 1224
rect 2770 1198 3150 1224
rect 3747 1285 3757 1305
rect 3777 1285 3784 1305
rect 3747 1280 3784 1285
rect 4403 1300 4513 1315
rect 4403 1297 4480 1300
rect 3747 1229 3782 1280
rect 4403 1270 4406 1297
rect 4435 1273 4480 1297
rect 4509 1273 4513 1300
rect 4435 1270 4513 1273
rect 4403 1256 4513 1270
rect 4699 1229 4747 1384
rect 3747 1205 4747 1229
rect 3747 1202 4746 1205
rect 3747 1200 3782 1202
rect 2738 1196 3150 1198
rect 2740 1195 2780 1196
rect 3118 1131 3150 1196
rect 3118 1111 3122 1131
rect 3143 1111 3150 1131
rect 3723 1114 4025 1116
rect 3118 1104 3150 1111
rect 3662 1085 4025 1114
rect 3662 1083 3723 1085
rect 2671 1038 2706 1046
rect 2671 1018 2679 1038
rect 2699 1018 2706 1038
rect 2671 1013 2706 1018
rect 3043 1039 3081 1045
rect 3043 1022 3053 1039
rect 3073 1022 3081 1039
rect 2671 1012 2703 1013
rect 2209 1008 2244 1009
rect 1152 981 1189 988
rect 1152 980 1187 981
rect 189 880 197 909
rect 226 880 237 909
rect 189 875 237 880
rect 708 915 740 922
rect 708 895 715 915
rect 736 895 740 915
rect 708 830 740 895
rect 1078 830 1118 831
rect 708 828 1120 830
rect 708 802 1088 828
rect 1114 802 1120 828
rect 708 794 1120 802
rect 708 766 740 794
rect 1153 774 1187 980
rect 1857 963 1896 970
rect 1500 935 1611 957
rect 1500 915 1508 935
rect 1527 915 1585 935
rect 1604 915 1611 935
rect 1500 898 1611 915
rect 1857 936 1861 963
rect 1892 936 1896 963
rect 1704 847 1757 851
rect 1222 812 1757 847
rect 708 746 713 766
rect 734 746 740 766
rect 708 739 740 746
rect 915 766 954 772
rect 915 746 923 766
rect 948 746 954 766
rect 915 739 954 746
rect 1131 769 1187 774
rect 1131 749 1138 769
rect 1158 749 1187 769
rect 1131 742 1187 749
rect 1131 741 1166 742
rect 923 693 954 739
rect 422 668 533 690
rect 422 648 430 668
rect 449 648 507 668
rect 526 648 533 668
rect 922 676 954 693
rect 1223 676 1260 812
rect 1361 779 1471 793
rect 1361 776 1439 779
rect 1361 749 1365 776
rect 1394 752 1439 776
rect 1468 752 1471 779
rect 1394 749 1471 752
rect 1361 734 1471 749
rect 1703 765 1757 812
rect 1703 757 1756 765
rect 1703 740 1712 757
rect 1744 740 1756 757
rect 1703 737 1756 740
rect 922 663 1260 676
rect 422 631 533 648
rect 923 644 1260 663
rect 1202 643 1260 644
rect 1646 671 1678 678
rect 1646 651 1653 671
rect 1674 651 1678 671
rect 1646 586 1678 651
rect 1857 663 1896 936
rect 2092 765 2126 776
rect 2090 764 2126 765
rect 2090 744 2097 764
rect 2117 744 2126 764
rect 2090 736 2126 744
rect 1857 622 1864 663
rect 1885 622 1896 663
rect 1857 607 1896 622
rect 2016 586 2056 587
rect 1646 584 2058 586
rect 1646 558 2026 584
rect 2052 558 2058 584
rect 1646 550 2058 558
rect 192 511 1188 537
rect 1646 522 1678 550
rect 2091 530 2125 736
rect 2833 692 2868 693
rect 194 458 236 511
rect 194 439 203 458
rect 228 439 236 458
rect 194 429 236 439
rect 422 469 532 483
rect 422 466 500 469
rect 422 439 426 466
rect 455 442 500 466
rect 529 442 532 469
rect 1152 459 1186 511
rect 1646 502 1651 522
rect 1672 502 1678 522
rect 1646 495 1678 502
rect 2069 525 2125 530
rect 2069 505 2076 525
rect 2096 505 2125 525
rect 2069 498 2125 505
rect 2812 685 2868 692
rect 2812 665 2841 685
rect 2861 665 2868 685
rect 2812 660 2868 665
rect 3043 684 3081 1022
rect 3325 1033 3435 1048
rect 3325 1030 3402 1033
rect 3325 1003 3328 1030
rect 3357 1006 3402 1030
rect 3431 1006 3435 1033
rect 3357 1003 3435 1006
rect 3325 989 3435 1003
rect 3204 863 3241 865
rect 3662 863 3695 1083
rect 3983 1004 4025 1085
rect 4405 1096 4516 1113
rect 4405 1076 4412 1096
rect 4431 1076 4489 1096
rect 4508 1076 4516 1096
rect 4405 1054 4516 1076
rect 3772 1002 3807 1003
rect 3204 834 3695 863
rect 3204 768 3241 834
rect 3662 833 3695 834
rect 3751 995 3807 1002
rect 3751 975 3780 995
rect 3800 975 3807 995
rect 3751 970 3807 975
rect 3981 1000 4025 1004
rect 3981 980 3992 1000
rect 4015 980 4025 1000
rect 3981 973 4025 980
rect 4198 998 4230 1005
rect 4198 978 4204 998
rect 4225 978 4230 998
rect 3981 971 4024 973
rect 3199 759 3241 768
rect 3199 737 3208 759
rect 3234 737 3241 759
rect 3466 786 3577 803
rect 3466 766 3473 786
rect 3492 766 3550 786
rect 3569 766 3577 786
rect 3466 744 3577 766
rect 3751 764 3785 970
rect 4198 950 4230 978
rect 3818 942 4230 950
rect 3818 916 3824 942
rect 3850 916 4230 942
rect 3818 914 4230 916
rect 3820 913 3860 914
rect 4198 849 4230 914
rect 4198 829 4202 849
rect 4223 829 4230 849
rect 4198 822 4230 829
rect 3751 756 3786 764
rect 3199 727 3241 737
rect 3751 736 3759 756
rect 3779 736 3786 756
rect 3751 731 3786 736
rect 4405 751 4515 766
rect 4405 748 4482 751
rect 3199 726 3240 727
rect 3043 667 3051 684
rect 3071 667 3081 684
rect 2069 497 2104 498
rect 1697 463 1738 464
rect 455 439 532 442
rect 422 424 532 439
rect 1151 454 1186 459
rect 1151 434 1158 454
rect 1178 434 1186 454
rect 1696 453 1738 463
rect 1151 426 1186 434
rect 707 361 739 368
rect 707 341 714 361
rect 735 341 739 361
rect 707 276 739 341
rect 1077 276 1117 277
rect 707 274 1119 276
rect 707 248 1087 274
rect 1113 248 1119 274
rect 707 240 1119 248
rect 707 212 739 240
rect 1152 220 1186 426
rect 1360 424 1471 446
rect 1360 404 1368 424
rect 1387 404 1445 424
rect 1464 404 1471 424
rect 1360 387 1471 404
rect 1696 431 1703 453
rect 1729 431 1738 453
rect 1696 422 1738 431
rect 2812 454 2846 660
rect 3043 657 3081 667
rect 3259 688 3291 695
rect 3259 668 3265 688
rect 3286 668 3291 688
rect 3751 679 3785 731
rect 4405 721 4408 748
rect 4437 724 4482 748
rect 4511 724 4515 751
rect 4437 721 4515 724
rect 4405 707 4515 721
rect 4701 751 4743 761
rect 4701 732 4709 751
rect 4734 732 4743 751
rect 4701 679 4743 732
rect 3259 640 3291 668
rect 3749 653 4745 679
rect 2879 632 3291 640
rect 2879 606 2885 632
rect 2911 606 3291 632
rect 2879 604 3291 606
rect 2881 603 2921 604
rect 3259 539 3291 604
rect 3259 519 3263 539
rect 3284 519 3291 539
rect 3259 512 3291 519
rect 3677 546 3735 547
rect 3677 527 4014 546
rect 4404 542 4515 559
rect 3677 514 4015 527
rect 2812 446 2847 454
rect 2812 426 2820 446
rect 2840 426 2847 446
rect 913 217 956 219
rect 707 192 712 212
rect 733 192 739 212
rect 707 185 739 192
rect 912 210 956 217
rect 912 190 922 210
rect 945 190 956 210
rect 912 186 956 190
rect 1130 215 1186 220
rect 1130 195 1137 215
rect 1157 195 1186 215
rect 1130 188 1186 195
rect 1242 356 1275 357
rect 1696 356 1733 422
rect 2812 421 2847 426
rect 3466 441 3576 456
rect 3466 438 3543 441
rect 2812 378 2846 421
rect 3466 411 3469 438
rect 3498 414 3543 438
rect 3572 414 3576 441
rect 3498 411 3576 414
rect 3466 397 3576 411
rect 3677 378 3714 514
rect 3983 497 4015 514
rect 4404 522 4411 542
rect 4430 522 4488 542
rect 4507 522 4515 542
rect 4404 500 4515 522
rect 3983 451 4014 497
rect 3771 448 3806 449
rect 3750 441 3806 448
rect 3750 421 3779 441
rect 3799 421 3806 441
rect 3750 416 3806 421
rect 3983 444 4022 451
rect 3983 424 3989 444
rect 4014 424 4022 444
rect 3983 418 4022 424
rect 4197 444 4229 451
rect 4197 424 4203 444
rect 4224 424 4229 444
rect 1242 327 1733 356
rect 2811 343 3715 378
rect 2812 342 2846 343
rect 1130 187 1165 188
rect 421 116 532 136
rect 421 114 531 116
rect 421 94 429 114
rect 448 94 506 114
rect 525 94 531 114
rect 421 77 531 94
rect 912 105 954 186
rect 1242 107 1275 327
rect 1696 325 1733 327
rect 3750 210 3784 416
rect 4197 396 4229 424
rect 3817 388 4229 396
rect 3817 362 3823 388
rect 3849 362 4229 388
rect 3817 360 4229 362
rect 3819 359 3859 360
rect 4197 295 4229 360
rect 4197 275 4201 295
rect 4222 275 4229 295
rect 4197 268 4229 275
rect 4700 310 4748 315
rect 4700 281 4711 310
rect 4740 281 4748 310
rect 3750 209 3785 210
rect 1214 105 1275 107
rect 912 76 1275 105
rect 3748 202 3785 209
rect 3748 182 3758 202
rect 3778 182 3785 202
rect 3748 177 3785 182
rect 4404 197 4514 212
rect 4404 194 4481 197
rect 3748 126 3783 177
rect 4404 167 4407 194
rect 4436 170 4481 194
rect 4510 170 4514 197
rect 4436 167 4514 170
rect 4404 153 4514 167
rect 4700 126 4748 281
rect 3748 102 4748 126
rect 3748 99 4747 102
rect 3748 97 3783 99
rect 912 74 1214 76
rect 718 45 797 49
rect 718 36 4829 45
rect 718 32 4792 36
rect 718 11 757 32
rect 786 15 4792 32
rect 4821 15 4829 36
rect 786 11 4829 15
rect 718 3 4829 11
rect 718 -8 797 3
rect 2384 -47 2443 -31
rect 1669 -90 1779 -76
rect 1669 -93 1747 -90
rect 1669 -120 1673 -93
rect 1702 -117 1747 -93
rect 1776 -117 1779 -90
rect 1702 -120 1779 -117
rect 1669 -135 1779 -120
rect 2384 -89 2403 -47
rect 2435 -89 2443 -47
rect 2384 -105 2443 -89
rect 2384 -125 2405 -105
rect 2425 -125 2443 -105
rect 2384 -130 2443 -125
rect 2472 -50 2532 -30
rect 2472 -113 2484 -50
rect 2515 -113 2532 -50
rect 2472 -128 2532 -113
rect 2398 -133 2433 -130
rect 1954 -198 1986 -191
rect 1954 -218 1961 -198
rect 1982 -218 1986 -198
rect 1954 -283 1986 -218
rect 2324 -283 2364 -282
rect 1954 -285 2366 -283
rect 1954 -311 2334 -285
rect 2360 -311 2366 -285
rect 1954 -319 2366 -311
rect 1954 -347 1986 -319
rect 2399 -339 2433 -133
rect 1954 -367 1959 -347
rect 1980 -367 1986 -347
rect 1954 -374 1986 -367
rect 2154 -348 2212 -341
rect 2154 -368 2165 -348
rect 2199 -368 2212 -348
rect 1668 -445 1779 -423
rect 1668 -465 1676 -445
rect 1695 -465 1753 -445
rect 1772 -465 1779 -445
rect 1668 -482 1779 -465
rect 2154 -518 2212 -368
rect 2377 -344 2433 -339
rect 2377 -364 2384 -344
rect 2404 -364 2433 -344
rect 2377 -371 2433 -364
rect 2377 -372 2412 -371
rect 2472 -405 2527 -128
rect 2472 -426 2486 -405
rect 2513 -426 2527 -405
rect 2472 -436 2527 -426
<< via1 >>
rect 2485 4620 2516 4673
rect 2405 4232 2436 4285
rect 2403 -89 2435 -47
rect 2484 -113 2515 -50
<< metal2 >>
rect 2473 4673 2521 4692
rect 2473 4620 2485 4673
rect 2516 4620 2521 4673
rect 2394 4285 2442 4300
rect 2394 4232 2405 4285
rect 2436 4232 2442 4285
rect 2394 -31 2442 4232
rect 2473 -30 2521 4620
rect 2384 -47 2443 -31
rect 2384 -89 2403 -47
rect 2435 -89 2443 -47
rect 2384 -130 2443 -89
rect 2472 -50 2532 -30
rect 2472 -113 2484 -50
rect 2515 -113 2532 -50
rect 2472 -128 2532 -113
<< labels >>
rlabel locali 290 8525 312 8540 1 d0
rlabel metal1 459 8748 487 8753 1 vdd
rlabel metal1 456 8355 490 8361 1 gnd
rlabel locali 1227 8277 1255 8298 1 d1
rlabel metal1 1394 8111 1428 8117 1 gnd
rlabel metal1 1397 8504 1425 8509 1 vdd
rlabel locali 289 7971 311 7986 1 d0
rlabel metal1 458 8194 486 8199 1 vdd
rlabel metal1 455 7801 489 7807 1 gnd
rlabel locali 110 8810 138 8818 1 vref
rlabel locali 291 7422 313 7437 1 d0
rlabel metal1 460 7645 488 7650 1 vdd
rlabel metal1 457 7252 491 7258 1 gnd
rlabel locali 1228 7174 1256 7195 1 d1
rlabel metal1 1395 7008 1429 7014 1 gnd
rlabel metal1 1398 7401 1426 7406 1 vdd
rlabel locali 290 6868 312 6883 1 d0
rlabel metal1 459 7091 487 7096 1 vdd
rlabel metal1 456 6698 490 6704 1 gnd
rlabel metal1 1538 7912 1566 7917 1 vdd
rlabel metal1 1535 7519 1569 7525 1 gnd
rlabel locali 1366 7684 1387 7703 1 d2
rlabel locali 291 6319 313 6334 1 d0
rlabel metal1 460 6542 488 6547 1 vdd
rlabel metal1 457 6149 491 6155 1 gnd
rlabel locali 1228 6071 1256 6092 1 d1
rlabel metal1 1395 5905 1429 5911 1 gnd
rlabel metal1 1398 6298 1426 6303 1 vdd
rlabel locali 290 5765 312 5780 1 d0
rlabel metal1 459 5988 487 5993 1 vdd
rlabel metal1 456 5595 490 5601 1 gnd
rlabel locali 292 5216 314 5231 1 d0
rlabel metal1 461 5439 489 5444 1 vdd
rlabel metal1 458 5046 492 5052 1 gnd
rlabel locali 1229 4968 1257 4989 1 d1
rlabel metal1 1396 4802 1430 4808 1 gnd
rlabel metal1 1399 5195 1427 5200 1 vdd
rlabel locali 291 4662 313 4677 1 d0
rlabel metal1 460 4885 488 4890 1 vdd
rlabel metal1 457 4492 491 4498 1 gnd
rlabel metal1 1539 5706 1567 5711 1 vdd
rlabel metal1 1536 5313 1570 5319 1 gnd
rlabel locali 1367 5478 1388 5497 1 d2
rlabel metal1 1508 6822 1536 6827 1 vdd
rlabel metal1 1505 6429 1539 6435 1 gnd
rlabel locali 1338 6598 1364 6615 1 d3
rlabel locali 1340 2186 1366 2203 1 d3
rlabel metal1 1507 2017 1541 2023 1 gnd
rlabel metal1 1510 2410 1538 2415 1 vdd
rlabel locali 1369 1066 1390 1085 1 d2
rlabel metal1 1538 901 1572 907 1 gnd
rlabel metal1 1541 1294 1569 1299 1 vdd
rlabel metal1 459 80 493 86 1 gnd
rlabel metal1 462 473 490 478 1 vdd
rlabel locali 293 250 315 265 1 d0
rlabel metal1 1401 783 1429 788 1 vdd
rlabel metal1 1398 390 1432 396 1 gnd
rlabel locali 1231 556 1259 577 1 d1
rlabel metal1 460 634 494 640 1 gnd
rlabel metal1 463 1027 491 1032 1 vdd
rlabel locali 294 804 316 819 1 d0
rlabel metal1 458 1183 492 1189 1 gnd
rlabel metal1 461 1576 489 1581 1 vdd
rlabel locali 292 1353 314 1368 1 d0
rlabel metal1 1400 1886 1428 1891 1 vdd
rlabel metal1 1397 1493 1431 1499 1 gnd
rlabel locali 1230 1659 1258 1680 1 d1
rlabel metal1 459 1737 493 1743 1 gnd
rlabel metal1 462 2130 490 2135 1 vdd
rlabel locali 293 1907 315 1922 1 d0
rlabel locali 1368 3272 1389 3291 1 d2
rlabel metal1 1537 3107 1571 3113 1 gnd
rlabel metal1 1540 3500 1568 3505 1 vdd
rlabel metal1 458 2286 492 2292 1 gnd
rlabel metal1 461 2679 489 2684 1 vdd
rlabel locali 292 2456 314 2471 1 d0
rlabel metal1 1400 2989 1428 2994 1 vdd
rlabel metal1 1397 2596 1431 2602 1 gnd
rlabel locali 1230 2762 1258 2783 1 d1
rlabel metal1 459 2840 493 2846 1 gnd
rlabel metal1 462 3233 490 3238 1 vdd
rlabel locali 293 3010 315 3025 1 d0
rlabel metal1 457 3389 491 3395 1 gnd
rlabel metal1 460 3782 488 3787 1 vdd
rlabel locali 291 3559 313 3574 1 d0
rlabel metal1 1399 4092 1427 4097 1 vdd
rlabel metal1 1396 3699 1430 3705 1 gnd
rlabel locali 1229 3865 1257 3886 1 d1
rlabel metal1 458 3943 492 3949 1 gnd
rlabel metal1 461 4336 489 4341 1 vdd
rlabel locali 292 4113 314 4128 1 d0
rlabel metal1 1508 4622 1536 4627 1 vdd
rlabel metal1 1505 4229 1539 4235 1 gnd
rlabel locali 1332 4391 1367 4417 1 d4
rlabel locali 4621 371 4643 386 5 d0
rlabel metal1 4446 158 4474 163 5 vdd
rlabel metal1 4443 550 4477 556 5 gnd
rlabel locali 3678 613 3706 634 5 d1
rlabel metal1 3505 794 3539 800 5 gnd
rlabel metal1 3508 402 3536 407 5 vdd
rlabel locali 4622 925 4644 940 5 d0
rlabel metal1 4447 712 4475 717 5 vdd
rlabel metal1 4444 1104 4478 1110 5 gnd
rlabel locali 4620 1474 4642 1489 5 d0
rlabel metal1 4445 1261 4473 1266 5 vdd
rlabel metal1 4442 1653 4476 1659 5 gnd
rlabel locali 3677 1716 3705 1737 5 d1
rlabel metal1 3504 1897 3538 1903 5 gnd
rlabel metal1 3507 1505 3535 1510 5 vdd
rlabel locali 4621 2028 4643 2043 5 d0
rlabel metal1 4446 1815 4474 1820 5 vdd
rlabel metal1 4443 2207 4477 2213 5 gnd
rlabel metal1 3367 994 3395 999 5 vdd
rlabel metal1 3364 1386 3398 1392 5 gnd
rlabel locali 3546 1208 3567 1227 5 d2
rlabel locali 4620 2577 4642 2592 5 d0
rlabel metal1 4445 2364 4473 2369 5 vdd
rlabel metal1 4442 2756 4476 2762 5 gnd
rlabel locali 3677 2819 3705 2840 5 d1
rlabel metal1 3504 3000 3538 3006 5 gnd
rlabel metal1 3507 2608 3535 2613 5 vdd
rlabel locali 4621 3131 4643 3146 5 d0
rlabel metal1 4446 2918 4474 2923 5 vdd
rlabel metal1 4443 3310 4477 3316 5 gnd
rlabel locali 4619 3680 4641 3695 5 d0
rlabel metal1 4444 3467 4472 3472 5 vdd
rlabel metal1 4441 3859 4475 3865 5 gnd
rlabel locali 3676 3922 3704 3943 5 d1
rlabel metal1 3503 4103 3537 4109 5 gnd
rlabel metal1 3506 3711 3534 3716 5 vdd
rlabel locali 4620 4234 4642 4249 5 d0
rlabel metal1 4445 4021 4473 4026 5 vdd
rlabel metal1 4442 4413 4476 4419 5 gnd
rlabel metal1 3366 3200 3394 3205 5 vdd
rlabel metal1 3363 3592 3397 3598 5 gnd
rlabel locali 3545 3414 3566 3433 5 d2
rlabel metal1 3397 2084 3425 2089 5 vdd
rlabel metal1 3394 2476 3428 2482 5 gnd
rlabel locali 3569 2296 3595 2313 5 d3
rlabel locali 3567 6708 3593 6725 5 d3
rlabel metal1 3392 6888 3426 6894 5 gnd
rlabel metal1 3395 6496 3423 6501 5 vdd
rlabel locali 3543 7826 3564 7845 5 d2
rlabel metal1 3361 8004 3395 8010 5 gnd
rlabel metal1 3364 7612 3392 7617 5 vdd
rlabel metal1 4440 8825 4474 8831 5 gnd
rlabel metal1 4443 8433 4471 8438 5 vdd
rlabel locali 4618 8646 4640 8661 5 d0
rlabel metal1 3504 8123 3532 8128 5 vdd
rlabel metal1 3501 8515 3535 8521 5 gnd
rlabel locali 3674 8334 3702 8355 5 d1
rlabel metal1 4439 8271 4473 8277 5 gnd
rlabel metal1 4442 7879 4470 7884 5 vdd
rlabel locali 4617 8092 4639 8107 5 d0
rlabel metal1 4441 7722 4475 7728 5 gnd
rlabel metal1 4444 7330 4472 7335 5 vdd
rlabel locali 4619 7543 4641 7558 5 d0
rlabel metal1 3505 7020 3533 7025 5 vdd
rlabel metal1 3502 7412 3536 7418 5 gnd
rlabel locali 3675 7231 3703 7252 5 d1
rlabel metal1 4440 7168 4474 7174 5 gnd
rlabel metal1 4443 6776 4471 6781 5 vdd
rlabel locali 4618 6989 4640 7004 5 d0
rlabel locali 3544 5620 3565 5639 5 d2
rlabel metal1 3362 5798 3396 5804 5 gnd
rlabel metal1 3365 5406 3393 5411 5 vdd
rlabel metal1 4441 6619 4475 6625 5 gnd
rlabel metal1 4444 6227 4472 6232 5 vdd
rlabel locali 4619 6440 4641 6455 5 d0
rlabel metal1 3505 5917 3533 5922 5 vdd
rlabel metal1 3502 6309 3536 6315 5 gnd
rlabel locali 3675 6128 3703 6149 5 d1
rlabel metal1 4440 6065 4474 6071 5 gnd
rlabel metal1 4443 5673 4471 5678 5 vdd
rlabel locali 4618 5886 4640 5901 5 d0
rlabel metal1 4442 5516 4476 5522 5 gnd
rlabel metal1 4445 5124 4473 5129 5 vdd
rlabel locali 4620 5337 4642 5352 5 d0
rlabel metal1 3506 4814 3534 4819 5 vdd
rlabel metal1 3503 5206 3537 5212 5 gnd
rlabel locali 3676 5025 3704 5046 5 d1
rlabel metal1 4441 4962 4475 4968 5 gnd
rlabel metal1 4444 4570 4472 4575 5 vdd
rlabel locali 4619 4783 4641 4798 5 d0
rlabel metal1 3397 4284 3425 4289 5 vdd
rlabel metal1 3394 4676 3428 4682 5 gnd
rlabel locali 3566 4494 3601 4520 5 d4
rlabel locali 2170 -274 2192 -259 1 vout
rlabel metal1 1709 -86 1737 -81 1 vdd
rlabel metal1 1706 -479 1740 -473 1 gnd
rlabel locali 1535 -315 1563 -293 1 d5
<< end >>
