magic
tech sky130A
timestamp 1620561391
<< nwell >>
rect 318 2085 645 2159
rect 318 1935 1129 2085
rect 1256 1841 1583 1915
rect 1256 1691 2067 1841
rect 317 1531 644 1605
rect 317 1381 1128 1531
rect 1397 1249 1724 1323
rect 1397 1099 2208 1249
rect 319 982 646 1056
rect 319 832 1130 982
rect 1257 738 1584 812
rect 1257 588 2068 738
rect 318 428 645 502
rect 318 278 1129 428
rect 1367 159 1694 233
rect 1367 9 2178 159
rect 319 -121 646 -47
rect 319 -271 1130 -121
rect 1257 -365 1584 -291
rect 1257 -515 2068 -365
rect 318 -675 645 -601
rect 318 -825 1129 -675
rect 1398 -957 1725 -883
rect 1398 -1107 2209 -957
rect 320 -1224 647 -1150
rect 320 -1374 1131 -1224
rect 1258 -1468 1585 -1394
rect 1258 -1618 2069 -1468
rect 319 -1778 646 -1704
rect 319 -1928 1130 -1778
<< nmos >>
rect 382 1834 432 1876
rect 595 1834 645 1876
rect 803 1834 853 1876
rect 1011 1834 1061 1876
rect 1320 1590 1370 1632
rect 1533 1590 1583 1632
rect 1741 1590 1791 1632
rect 1949 1590 1999 1632
rect 381 1280 431 1322
rect 594 1280 644 1322
rect 802 1280 852 1322
rect 1010 1280 1060 1322
rect 1461 998 1511 1040
rect 1674 998 1724 1040
rect 1882 998 1932 1040
rect 2090 998 2140 1040
rect 383 731 433 773
rect 596 731 646 773
rect 804 731 854 773
rect 1012 731 1062 773
rect 1321 487 1371 529
rect 1534 487 1584 529
rect 1742 487 1792 529
rect 1950 487 2000 529
rect 382 177 432 219
rect 595 177 645 219
rect 803 177 853 219
rect 1011 177 1061 219
rect 1431 -92 1481 -50
rect 1644 -92 1694 -50
rect 1852 -92 1902 -50
rect 2060 -92 2110 -50
rect 383 -372 433 -330
rect 596 -372 646 -330
rect 804 -372 854 -330
rect 1012 -372 1062 -330
rect 1321 -616 1371 -574
rect 1534 -616 1584 -574
rect 1742 -616 1792 -574
rect 1950 -616 2000 -574
rect 382 -926 432 -884
rect 595 -926 645 -884
rect 803 -926 853 -884
rect 1011 -926 1061 -884
rect 1462 -1208 1512 -1166
rect 1675 -1208 1725 -1166
rect 1883 -1208 1933 -1166
rect 2091 -1208 2141 -1166
rect 384 -1475 434 -1433
rect 597 -1475 647 -1433
rect 805 -1475 855 -1433
rect 1013 -1475 1063 -1433
rect 1322 -1719 1372 -1677
rect 1535 -1719 1585 -1677
rect 1743 -1719 1793 -1677
rect 1951 -1719 2001 -1677
rect 383 -2029 433 -1987
rect 596 -2029 646 -1987
rect 804 -2029 854 -1987
rect 1012 -2029 1062 -1987
<< pmos >>
rect 382 1953 432 2053
rect 595 1953 645 2053
rect 803 1953 853 2053
rect 1011 1953 1061 2053
rect 1320 1709 1370 1809
rect 1533 1709 1583 1809
rect 1741 1709 1791 1809
rect 1949 1709 1999 1809
rect 381 1399 431 1499
rect 594 1399 644 1499
rect 802 1399 852 1499
rect 1010 1399 1060 1499
rect 1461 1117 1511 1217
rect 1674 1117 1724 1217
rect 1882 1117 1932 1217
rect 2090 1117 2140 1217
rect 383 850 433 950
rect 596 850 646 950
rect 804 850 854 950
rect 1012 850 1062 950
rect 1321 606 1371 706
rect 1534 606 1584 706
rect 1742 606 1792 706
rect 1950 606 2000 706
rect 382 296 432 396
rect 595 296 645 396
rect 803 296 853 396
rect 1011 296 1061 396
rect 1431 27 1481 127
rect 1644 27 1694 127
rect 1852 27 1902 127
rect 2060 27 2110 127
rect 383 -253 433 -153
rect 596 -253 646 -153
rect 804 -253 854 -153
rect 1012 -253 1062 -153
rect 1321 -497 1371 -397
rect 1534 -497 1584 -397
rect 1742 -497 1792 -397
rect 1950 -497 2000 -397
rect 382 -807 432 -707
rect 595 -807 645 -707
rect 803 -807 853 -707
rect 1011 -807 1061 -707
rect 1462 -1089 1512 -989
rect 1675 -1089 1725 -989
rect 1883 -1089 1933 -989
rect 2091 -1089 2141 -989
rect 384 -1356 434 -1256
rect 597 -1356 647 -1256
rect 805 -1356 855 -1256
rect 1013 -1356 1063 -1256
rect 1322 -1600 1372 -1500
rect 1535 -1600 1585 -1500
rect 1743 -1600 1793 -1500
rect 1951 -1600 2001 -1500
rect 383 -1910 433 -1810
rect 596 -1910 646 -1810
rect 804 -1910 854 -1810
rect 1012 -1910 1062 -1810
<< ndiff >>
rect 333 1866 382 1876
rect 333 1846 344 1866
rect 364 1846 382 1866
rect 333 1834 382 1846
rect 432 1870 476 1876
rect 432 1850 447 1870
rect 467 1850 476 1870
rect 432 1834 476 1850
rect 546 1866 595 1876
rect 546 1846 557 1866
rect 577 1846 595 1866
rect 546 1834 595 1846
rect 645 1870 689 1876
rect 645 1850 660 1870
rect 680 1850 689 1870
rect 645 1834 689 1850
rect 754 1866 803 1876
rect 754 1846 765 1866
rect 785 1846 803 1866
rect 754 1834 803 1846
rect 853 1870 897 1876
rect 853 1850 868 1870
rect 888 1850 897 1870
rect 853 1834 897 1850
rect 967 1870 1011 1876
rect 967 1850 976 1870
rect 996 1850 1011 1870
rect 967 1834 1011 1850
rect 1061 1866 1110 1876
rect 1061 1846 1079 1866
rect 1099 1846 1110 1866
rect 1061 1834 1110 1846
rect 1271 1622 1320 1632
rect 1271 1602 1282 1622
rect 1302 1602 1320 1622
rect 1271 1590 1320 1602
rect 1370 1626 1414 1632
rect 1370 1606 1385 1626
rect 1405 1606 1414 1626
rect 1370 1590 1414 1606
rect 1484 1622 1533 1632
rect 1484 1602 1495 1622
rect 1515 1602 1533 1622
rect 1484 1590 1533 1602
rect 1583 1626 1627 1632
rect 1583 1606 1598 1626
rect 1618 1606 1627 1626
rect 1583 1590 1627 1606
rect 1692 1622 1741 1632
rect 1692 1602 1703 1622
rect 1723 1602 1741 1622
rect 1692 1590 1741 1602
rect 1791 1626 1835 1632
rect 1791 1606 1806 1626
rect 1826 1606 1835 1626
rect 1791 1590 1835 1606
rect 1905 1626 1949 1632
rect 1905 1606 1914 1626
rect 1934 1606 1949 1626
rect 1905 1590 1949 1606
rect 1999 1622 2048 1632
rect 1999 1602 2017 1622
rect 2037 1602 2048 1622
rect 1999 1590 2048 1602
rect 332 1312 381 1322
rect 332 1292 343 1312
rect 363 1292 381 1312
rect 332 1280 381 1292
rect 431 1316 475 1322
rect 431 1296 446 1316
rect 466 1296 475 1316
rect 431 1280 475 1296
rect 545 1312 594 1322
rect 545 1292 556 1312
rect 576 1292 594 1312
rect 545 1280 594 1292
rect 644 1316 688 1322
rect 644 1296 659 1316
rect 679 1296 688 1316
rect 644 1280 688 1296
rect 753 1312 802 1322
rect 753 1292 764 1312
rect 784 1292 802 1312
rect 753 1280 802 1292
rect 852 1316 896 1322
rect 852 1296 867 1316
rect 887 1296 896 1316
rect 852 1280 896 1296
rect 966 1316 1010 1322
rect 966 1296 975 1316
rect 995 1296 1010 1316
rect 966 1280 1010 1296
rect 1060 1312 1109 1322
rect 1060 1292 1078 1312
rect 1098 1292 1109 1312
rect 1060 1280 1109 1292
rect 1412 1030 1461 1040
rect 1412 1010 1423 1030
rect 1443 1010 1461 1030
rect 1412 998 1461 1010
rect 1511 1034 1555 1040
rect 1511 1014 1526 1034
rect 1546 1014 1555 1034
rect 1511 998 1555 1014
rect 1625 1030 1674 1040
rect 1625 1010 1636 1030
rect 1656 1010 1674 1030
rect 1625 998 1674 1010
rect 1724 1034 1768 1040
rect 1724 1014 1739 1034
rect 1759 1014 1768 1034
rect 1724 998 1768 1014
rect 1833 1030 1882 1040
rect 1833 1010 1844 1030
rect 1864 1010 1882 1030
rect 1833 998 1882 1010
rect 1932 1034 1976 1040
rect 1932 1014 1947 1034
rect 1967 1014 1976 1034
rect 1932 998 1976 1014
rect 2046 1034 2090 1040
rect 2046 1014 2055 1034
rect 2075 1014 2090 1034
rect 2046 998 2090 1014
rect 2140 1030 2189 1040
rect 2140 1010 2158 1030
rect 2178 1010 2189 1030
rect 2140 998 2189 1010
rect 334 763 383 773
rect 334 743 345 763
rect 365 743 383 763
rect 334 731 383 743
rect 433 767 477 773
rect 433 747 448 767
rect 468 747 477 767
rect 433 731 477 747
rect 547 763 596 773
rect 547 743 558 763
rect 578 743 596 763
rect 547 731 596 743
rect 646 767 690 773
rect 646 747 661 767
rect 681 747 690 767
rect 646 731 690 747
rect 755 763 804 773
rect 755 743 766 763
rect 786 743 804 763
rect 755 731 804 743
rect 854 767 898 773
rect 854 747 869 767
rect 889 747 898 767
rect 854 731 898 747
rect 968 767 1012 773
rect 968 747 977 767
rect 997 747 1012 767
rect 968 731 1012 747
rect 1062 763 1111 773
rect 1062 743 1080 763
rect 1100 743 1111 763
rect 1062 731 1111 743
rect 1272 519 1321 529
rect 1272 499 1283 519
rect 1303 499 1321 519
rect 1272 487 1321 499
rect 1371 523 1415 529
rect 1371 503 1386 523
rect 1406 503 1415 523
rect 1371 487 1415 503
rect 1485 519 1534 529
rect 1485 499 1496 519
rect 1516 499 1534 519
rect 1485 487 1534 499
rect 1584 523 1628 529
rect 1584 503 1599 523
rect 1619 503 1628 523
rect 1584 487 1628 503
rect 1693 519 1742 529
rect 1693 499 1704 519
rect 1724 499 1742 519
rect 1693 487 1742 499
rect 1792 523 1836 529
rect 1792 503 1807 523
rect 1827 503 1836 523
rect 1792 487 1836 503
rect 1906 523 1950 529
rect 1906 503 1915 523
rect 1935 503 1950 523
rect 1906 487 1950 503
rect 2000 519 2049 529
rect 2000 499 2018 519
rect 2038 499 2049 519
rect 2000 487 2049 499
rect 333 209 382 219
rect 333 189 344 209
rect 364 189 382 209
rect 333 177 382 189
rect 432 213 476 219
rect 432 193 447 213
rect 467 193 476 213
rect 432 177 476 193
rect 546 209 595 219
rect 546 189 557 209
rect 577 189 595 209
rect 546 177 595 189
rect 645 213 689 219
rect 645 193 660 213
rect 680 193 689 213
rect 645 177 689 193
rect 754 209 803 219
rect 754 189 765 209
rect 785 189 803 209
rect 754 177 803 189
rect 853 213 897 219
rect 853 193 868 213
rect 888 193 897 213
rect 853 177 897 193
rect 967 213 1011 219
rect 967 193 976 213
rect 996 193 1011 213
rect 967 177 1011 193
rect 1061 209 1110 219
rect 1061 189 1079 209
rect 1099 189 1110 209
rect 1061 177 1110 189
rect 1382 -60 1431 -50
rect 1382 -80 1393 -60
rect 1413 -80 1431 -60
rect 1382 -92 1431 -80
rect 1481 -56 1525 -50
rect 1481 -76 1496 -56
rect 1516 -76 1525 -56
rect 1481 -92 1525 -76
rect 1595 -60 1644 -50
rect 1595 -80 1606 -60
rect 1626 -80 1644 -60
rect 1595 -92 1644 -80
rect 1694 -56 1738 -50
rect 1694 -76 1709 -56
rect 1729 -76 1738 -56
rect 1694 -92 1738 -76
rect 1803 -60 1852 -50
rect 1803 -80 1814 -60
rect 1834 -80 1852 -60
rect 1803 -92 1852 -80
rect 1902 -56 1946 -50
rect 1902 -76 1917 -56
rect 1937 -76 1946 -56
rect 1902 -92 1946 -76
rect 2016 -56 2060 -50
rect 2016 -76 2025 -56
rect 2045 -76 2060 -56
rect 2016 -92 2060 -76
rect 2110 -60 2159 -50
rect 2110 -80 2128 -60
rect 2148 -80 2159 -60
rect 2110 -92 2159 -80
rect 334 -340 383 -330
rect 334 -360 345 -340
rect 365 -360 383 -340
rect 334 -372 383 -360
rect 433 -336 477 -330
rect 433 -356 448 -336
rect 468 -356 477 -336
rect 433 -372 477 -356
rect 547 -340 596 -330
rect 547 -360 558 -340
rect 578 -360 596 -340
rect 547 -372 596 -360
rect 646 -336 690 -330
rect 646 -356 661 -336
rect 681 -356 690 -336
rect 646 -372 690 -356
rect 755 -340 804 -330
rect 755 -360 766 -340
rect 786 -360 804 -340
rect 755 -372 804 -360
rect 854 -336 898 -330
rect 854 -356 869 -336
rect 889 -356 898 -336
rect 854 -372 898 -356
rect 968 -336 1012 -330
rect 968 -356 977 -336
rect 997 -356 1012 -336
rect 968 -372 1012 -356
rect 1062 -340 1111 -330
rect 1062 -360 1080 -340
rect 1100 -360 1111 -340
rect 1062 -372 1111 -360
rect 1272 -584 1321 -574
rect 1272 -604 1283 -584
rect 1303 -604 1321 -584
rect 1272 -616 1321 -604
rect 1371 -580 1415 -574
rect 1371 -600 1386 -580
rect 1406 -600 1415 -580
rect 1371 -616 1415 -600
rect 1485 -584 1534 -574
rect 1485 -604 1496 -584
rect 1516 -604 1534 -584
rect 1485 -616 1534 -604
rect 1584 -580 1628 -574
rect 1584 -600 1599 -580
rect 1619 -600 1628 -580
rect 1584 -616 1628 -600
rect 1693 -584 1742 -574
rect 1693 -604 1704 -584
rect 1724 -604 1742 -584
rect 1693 -616 1742 -604
rect 1792 -580 1836 -574
rect 1792 -600 1807 -580
rect 1827 -600 1836 -580
rect 1792 -616 1836 -600
rect 1906 -580 1950 -574
rect 1906 -600 1915 -580
rect 1935 -600 1950 -580
rect 1906 -616 1950 -600
rect 2000 -584 2049 -574
rect 2000 -604 2018 -584
rect 2038 -604 2049 -584
rect 2000 -616 2049 -604
rect 333 -894 382 -884
rect 333 -914 344 -894
rect 364 -914 382 -894
rect 333 -926 382 -914
rect 432 -890 476 -884
rect 432 -910 447 -890
rect 467 -910 476 -890
rect 432 -926 476 -910
rect 546 -894 595 -884
rect 546 -914 557 -894
rect 577 -914 595 -894
rect 546 -926 595 -914
rect 645 -890 689 -884
rect 645 -910 660 -890
rect 680 -910 689 -890
rect 645 -926 689 -910
rect 754 -894 803 -884
rect 754 -914 765 -894
rect 785 -914 803 -894
rect 754 -926 803 -914
rect 853 -890 897 -884
rect 853 -910 868 -890
rect 888 -910 897 -890
rect 853 -926 897 -910
rect 967 -890 1011 -884
rect 967 -910 976 -890
rect 996 -910 1011 -890
rect 967 -926 1011 -910
rect 1061 -894 1110 -884
rect 1061 -914 1079 -894
rect 1099 -914 1110 -894
rect 1061 -926 1110 -914
rect 1413 -1176 1462 -1166
rect 1413 -1196 1424 -1176
rect 1444 -1196 1462 -1176
rect 1413 -1208 1462 -1196
rect 1512 -1172 1556 -1166
rect 1512 -1192 1527 -1172
rect 1547 -1192 1556 -1172
rect 1512 -1208 1556 -1192
rect 1626 -1176 1675 -1166
rect 1626 -1196 1637 -1176
rect 1657 -1196 1675 -1176
rect 1626 -1208 1675 -1196
rect 1725 -1172 1769 -1166
rect 1725 -1192 1740 -1172
rect 1760 -1192 1769 -1172
rect 1725 -1208 1769 -1192
rect 1834 -1176 1883 -1166
rect 1834 -1196 1845 -1176
rect 1865 -1196 1883 -1176
rect 1834 -1208 1883 -1196
rect 1933 -1172 1977 -1166
rect 1933 -1192 1948 -1172
rect 1968 -1192 1977 -1172
rect 1933 -1208 1977 -1192
rect 2047 -1172 2091 -1166
rect 2047 -1192 2056 -1172
rect 2076 -1192 2091 -1172
rect 2047 -1208 2091 -1192
rect 2141 -1176 2190 -1166
rect 2141 -1196 2159 -1176
rect 2179 -1196 2190 -1176
rect 2141 -1208 2190 -1196
rect 335 -1443 384 -1433
rect 335 -1463 346 -1443
rect 366 -1463 384 -1443
rect 335 -1475 384 -1463
rect 434 -1439 478 -1433
rect 434 -1459 449 -1439
rect 469 -1459 478 -1439
rect 434 -1475 478 -1459
rect 548 -1443 597 -1433
rect 548 -1463 559 -1443
rect 579 -1463 597 -1443
rect 548 -1475 597 -1463
rect 647 -1439 691 -1433
rect 647 -1459 662 -1439
rect 682 -1459 691 -1439
rect 647 -1475 691 -1459
rect 756 -1443 805 -1433
rect 756 -1463 767 -1443
rect 787 -1463 805 -1443
rect 756 -1475 805 -1463
rect 855 -1439 899 -1433
rect 855 -1459 870 -1439
rect 890 -1459 899 -1439
rect 855 -1475 899 -1459
rect 969 -1439 1013 -1433
rect 969 -1459 978 -1439
rect 998 -1459 1013 -1439
rect 969 -1475 1013 -1459
rect 1063 -1443 1112 -1433
rect 1063 -1463 1081 -1443
rect 1101 -1463 1112 -1443
rect 1063 -1475 1112 -1463
rect 1273 -1687 1322 -1677
rect 1273 -1707 1284 -1687
rect 1304 -1707 1322 -1687
rect 1273 -1719 1322 -1707
rect 1372 -1683 1416 -1677
rect 1372 -1703 1387 -1683
rect 1407 -1703 1416 -1683
rect 1372 -1719 1416 -1703
rect 1486 -1687 1535 -1677
rect 1486 -1707 1497 -1687
rect 1517 -1707 1535 -1687
rect 1486 -1719 1535 -1707
rect 1585 -1683 1629 -1677
rect 1585 -1703 1600 -1683
rect 1620 -1703 1629 -1683
rect 1585 -1719 1629 -1703
rect 1694 -1687 1743 -1677
rect 1694 -1707 1705 -1687
rect 1725 -1707 1743 -1687
rect 1694 -1719 1743 -1707
rect 1793 -1683 1837 -1677
rect 1793 -1703 1808 -1683
rect 1828 -1703 1837 -1683
rect 1793 -1719 1837 -1703
rect 1907 -1683 1951 -1677
rect 1907 -1703 1916 -1683
rect 1936 -1703 1951 -1683
rect 1907 -1719 1951 -1703
rect 2001 -1687 2050 -1677
rect 2001 -1707 2019 -1687
rect 2039 -1707 2050 -1687
rect 2001 -1719 2050 -1707
rect 334 -1997 383 -1987
rect 334 -2017 345 -1997
rect 365 -2017 383 -1997
rect 334 -2029 383 -2017
rect 433 -1993 477 -1987
rect 433 -2013 448 -1993
rect 468 -2013 477 -1993
rect 433 -2029 477 -2013
rect 547 -1997 596 -1987
rect 547 -2017 558 -1997
rect 578 -2017 596 -1997
rect 547 -2029 596 -2017
rect 646 -1993 690 -1987
rect 646 -2013 661 -1993
rect 681 -2013 690 -1993
rect 646 -2029 690 -2013
rect 755 -1997 804 -1987
rect 755 -2017 766 -1997
rect 786 -2017 804 -1997
rect 755 -2029 804 -2017
rect 854 -1993 898 -1987
rect 854 -2013 869 -1993
rect 889 -2013 898 -1993
rect 854 -2029 898 -2013
rect 968 -1993 1012 -1987
rect 968 -2013 977 -1993
rect 997 -2013 1012 -1993
rect 968 -2029 1012 -2013
rect 1062 -1997 1111 -1987
rect 1062 -2017 1080 -1997
rect 1100 -2017 1111 -1997
rect 1062 -2029 1111 -2017
<< pdiff >>
rect 338 2015 382 2053
rect 338 1995 350 2015
rect 370 1995 382 2015
rect 338 1953 382 1995
rect 432 2015 474 2053
rect 432 1995 446 2015
rect 466 1995 474 2015
rect 432 1953 474 1995
rect 551 2015 595 2053
rect 551 1995 563 2015
rect 583 1995 595 2015
rect 551 1953 595 1995
rect 645 2015 687 2053
rect 645 1995 659 2015
rect 679 1995 687 2015
rect 645 1953 687 1995
rect 759 2015 803 2053
rect 759 1995 771 2015
rect 791 1995 803 2015
rect 759 1953 803 1995
rect 853 2015 895 2053
rect 853 1995 867 2015
rect 887 1995 895 2015
rect 853 1953 895 1995
rect 969 2015 1011 2053
rect 969 1995 977 2015
rect 997 1995 1011 2015
rect 969 1953 1011 1995
rect 1061 2022 1106 2053
rect 1061 2015 1105 2022
rect 1061 1995 1073 2015
rect 1093 1995 1105 2015
rect 1061 1953 1105 1995
rect 1276 1771 1320 1809
rect 1276 1751 1288 1771
rect 1308 1751 1320 1771
rect 1276 1709 1320 1751
rect 1370 1771 1412 1809
rect 1370 1751 1384 1771
rect 1404 1751 1412 1771
rect 1370 1709 1412 1751
rect 1489 1771 1533 1809
rect 1489 1751 1501 1771
rect 1521 1751 1533 1771
rect 1489 1709 1533 1751
rect 1583 1771 1625 1809
rect 1583 1751 1597 1771
rect 1617 1751 1625 1771
rect 1583 1709 1625 1751
rect 1697 1771 1741 1809
rect 1697 1751 1709 1771
rect 1729 1751 1741 1771
rect 1697 1709 1741 1751
rect 1791 1771 1833 1809
rect 1791 1751 1805 1771
rect 1825 1751 1833 1771
rect 1791 1709 1833 1751
rect 1907 1771 1949 1809
rect 1907 1751 1915 1771
rect 1935 1751 1949 1771
rect 1907 1709 1949 1751
rect 1999 1778 2044 1809
rect 1999 1771 2043 1778
rect 1999 1751 2011 1771
rect 2031 1751 2043 1771
rect 1999 1709 2043 1751
rect 337 1461 381 1499
rect 337 1441 349 1461
rect 369 1441 381 1461
rect 337 1399 381 1441
rect 431 1461 473 1499
rect 431 1441 445 1461
rect 465 1441 473 1461
rect 431 1399 473 1441
rect 550 1461 594 1499
rect 550 1441 562 1461
rect 582 1441 594 1461
rect 550 1399 594 1441
rect 644 1461 686 1499
rect 644 1441 658 1461
rect 678 1441 686 1461
rect 644 1399 686 1441
rect 758 1461 802 1499
rect 758 1441 770 1461
rect 790 1441 802 1461
rect 758 1399 802 1441
rect 852 1461 894 1499
rect 852 1441 866 1461
rect 886 1441 894 1461
rect 852 1399 894 1441
rect 968 1461 1010 1499
rect 968 1441 976 1461
rect 996 1441 1010 1461
rect 968 1399 1010 1441
rect 1060 1468 1105 1499
rect 1060 1461 1104 1468
rect 1060 1441 1072 1461
rect 1092 1441 1104 1461
rect 1060 1399 1104 1441
rect 1417 1179 1461 1217
rect 1417 1159 1429 1179
rect 1449 1159 1461 1179
rect 1417 1117 1461 1159
rect 1511 1179 1553 1217
rect 1511 1159 1525 1179
rect 1545 1159 1553 1179
rect 1511 1117 1553 1159
rect 1630 1179 1674 1217
rect 1630 1159 1642 1179
rect 1662 1159 1674 1179
rect 1630 1117 1674 1159
rect 1724 1179 1766 1217
rect 1724 1159 1738 1179
rect 1758 1159 1766 1179
rect 1724 1117 1766 1159
rect 1838 1179 1882 1217
rect 1838 1159 1850 1179
rect 1870 1159 1882 1179
rect 1838 1117 1882 1159
rect 1932 1179 1974 1217
rect 1932 1159 1946 1179
rect 1966 1159 1974 1179
rect 1932 1117 1974 1159
rect 2048 1179 2090 1217
rect 2048 1159 2056 1179
rect 2076 1159 2090 1179
rect 2048 1117 2090 1159
rect 2140 1186 2185 1217
rect 2140 1179 2184 1186
rect 2140 1159 2152 1179
rect 2172 1159 2184 1179
rect 2140 1117 2184 1159
rect 339 912 383 950
rect 339 892 351 912
rect 371 892 383 912
rect 339 850 383 892
rect 433 912 475 950
rect 433 892 447 912
rect 467 892 475 912
rect 433 850 475 892
rect 552 912 596 950
rect 552 892 564 912
rect 584 892 596 912
rect 552 850 596 892
rect 646 912 688 950
rect 646 892 660 912
rect 680 892 688 912
rect 646 850 688 892
rect 760 912 804 950
rect 760 892 772 912
rect 792 892 804 912
rect 760 850 804 892
rect 854 912 896 950
rect 854 892 868 912
rect 888 892 896 912
rect 854 850 896 892
rect 970 912 1012 950
rect 970 892 978 912
rect 998 892 1012 912
rect 970 850 1012 892
rect 1062 919 1107 950
rect 1062 912 1106 919
rect 1062 892 1074 912
rect 1094 892 1106 912
rect 1062 850 1106 892
rect 1277 668 1321 706
rect 1277 648 1289 668
rect 1309 648 1321 668
rect 1277 606 1321 648
rect 1371 668 1413 706
rect 1371 648 1385 668
rect 1405 648 1413 668
rect 1371 606 1413 648
rect 1490 668 1534 706
rect 1490 648 1502 668
rect 1522 648 1534 668
rect 1490 606 1534 648
rect 1584 668 1626 706
rect 1584 648 1598 668
rect 1618 648 1626 668
rect 1584 606 1626 648
rect 1698 668 1742 706
rect 1698 648 1710 668
rect 1730 648 1742 668
rect 1698 606 1742 648
rect 1792 668 1834 706
rect 1792 648 1806 668
rect 1826 648 1834 668
rect 1792 606 1834 648
rect 1908 668 1950 706
rect 1908 648 1916 668
rect 1936 648 1950 668
rect 1908 606 1950 648
rect 2000 675 2045 706
rect 2000 668 2044 675
rect 2000 648 2012 668
rect 2032 648 2044 668
rect 2000 606 2044 648
rect 338 358 382 396
rect 338 338 350 358
rect 370 338 382 358
rect 338 296 382 338
rect 432 358 474 396
rect 432 338 446 358
rect 466 338 474 358
rect 432 296 474 338
rect 551 358 595 396
rect 551 338 563 358
rect 583 338 595 358
rect 551 296 595 338
rect 645 358 687 396
rect 645 338 659 358
rect 679 338 687 358
rect 645 296 687 338
rect 759 358 803 396
rect 759 338 771 358
rect 791 338 803 358
rect 759 296 803 338
rect 853 358 895 396
rect 853 338 867 358
rect 887 338 895 358
rect 853 296 895 338
rect 969 358 1011 396
rect 969 338 977 358
rect 997 338 1011 358
rect 969 296 1011 338
rect 1061 365 1106 396
rect 1061 358 1105 365
rect 1061 338 1073 358
rect 1093 338 1105 358
rect 1061 296 1105 338
rect 1387 89 1431 127
rect 1387 69 1399 89
rect 1419 69 1431 89
rect 1387 27 1431 69
rect 1481 89 1523 127
rect 1481 69 1495 89
rect 1515 69 1523 89
rect 1481 27 1523 69
rect 1600 89 1644 127
rect 1600 69 1612 89
rect 1632 69 1644 89
rect 1600 27 1644 69
rect 1694 89 1736 127
rect 1694 69 1708 89
rect 1728 69 1736 89
rect 1694 27 1736 69
rect 1808 89 1852 127
rect 1808 69 1820 89
rect 1840 69 1852 89
rect 1808 27 1852 69
rect 1902 89 1944 127
rect 1902 69 1916 89
rect 1936 69 1944 89
rect 1902 27 1944 69
rect 2018 89 2060 127
rect 2018 69 2026 89
rect 2046 69 2060 89
rect 2018 27 2060 69
rect 2110 96 2155 127
rect 2110 89 2154 96
rect 2110 69 2122 89
rect 2142 69 2154 89
rect 2110 27 2154 69
rect 339 -191 383 -153
rect 339 -211 351 -191
rect 371 -211 383 -191
rect 339 -253 383 -211
rect 433 -191 475 -153
rect 433 -211 447 -191
rect 467 -211 475 -191
rect 433 -253 475 -211
rect 552 -191 596 -153
rect 552 -211 564 -191
rect 584 -211 596 -191
rect 552 -253 596 -211
rect 646 -191 688 -153
rect 646 -211 660 -191
rect 680 -211 688 -191
rect 646 -253 688 -211
rect 760 -191 804 -153
rect 760 -211 772 -191
rect 792 -211 804 -191
rect 760 -253 804 -211
rect 854 -191 896 -153
rect 854 -211 868 -191
rect 888 -211 896 -191
rect 854 -253 896 -211
rect 970 -191 1012 -153
rect 970 -211 978 -191
rect 998 -211 1012 -191
rect 970 -253 1012 -211
rect 1062 -184 1107 -153
rect 1062 -191 1106 -184
rect 1062 -211 1074 -191
rect 1094 -211 1106 -191
rect 1062 -253 1106 -211
rect 1277 -435 1321 -397
rect 1277 -455 1289 -435
rect 1309 -455 1321 -435
rect 1277 -497 1321 -455
rect 1371 -435 1413 -397
rect 1371 -455 1385 -435
rect 1405 -455 1413 -435
rect 1371 -497 1413 -455
rect 1490 -435 1534 -397
rect 1490 -455 1502 -435
rect 1522 -455 1534 -435
rect 1490 -497 1534 -455
rect 1584 -435 1626 -397
rect 1584 -455 1598 -435
rect 1618 -455 1626 -435
rect 1584 -497 1626 -455
rect 1698 -435 1742 -397
rect 1698 -455 1710 -435
rect 1730 -455 1742 -435
rect 1698 -497 1742 -455
rect 1792 -435 1834 -397
rect 1792 -455 1806 -435
rect 1826 -455 1834 -435
rect 1792 -497 1834 -455
rect 1908 -435 1950 -397
rect 1908 -455 1916 -435
rect 1936 -455 1950 -435
rect 1908 -497 1950 -455
rect 2000 -428 2045 -397
rect 2000 -435 2044 -428
rect 2000 -455 2012 -435
rect 2032 -455 2044 -435
rect 2000 -497 2044 -455
rect 338 -745 382 -707
rect 338 -765 350 -745
rect 370 -765 382 -745
rect 338 -807 382 -765
rect 432 -745 474 -707
rect 432 -765 446 -745
rect 466 -765 474 -745
rect 432 -807 474 -765
rect 551 -745 595 -707
rect 551 -765 563 -745
rect 583 -765 595 -745
rect 551 -807 595 -765
rect 645 -745 687 -707
rect 645 -765 659 -745
rect 679 -765 687 -745
rect 645 -807 687 -765
rect 759 -745 803 -707
rect 759 -765 771 -745
rect 791 -765 803 -745
rect 759 -807 803 -765
rect 853 -745 895 -707
rect 853 -765 867 -745
rect 887 -765 895 -745
rect 853 -807 895 -765
rect 969 -745 1011 -707
rect 969 -765 977 -745
rect 997 -765 1011 -745
rect 969 -807 1011 -765
rect 1061 -738 1106 -707
rect 1061 -745 1105 -738
rect 1061 -765 1073 -745
rect 1093 -765 1105 -745
rect 1061 -807 1105 -765
rect 1418 -1027 1462 -989
rect 1418 -1047 1430 -1027
rect 1450 -1047 1462 -1027
rect 1418 -1089 1462 -1047
rect 1512 -1027 1554 -989
rect 1512 -1047 1526 -1027
rect 1546 -1047 1554 -1027
rect 1512 -1089 1554 -1047
rect 1631 -1027 1675 -989
rect 1631 -1047 1643 -1027
rect 1663 -1047 1675 -1027
rect 1631 -1089 1675 -1047
rect 1725 -1027 1767 -989
rect 1725 -1047 1739 -1027
rect 1759 -1047 1767 -1027
rect 1725 -1089 1767 -1047
rect 1839 -1027 1883 -989
rect 1839 -1047 1851 -1027
rect 1871 -1047 1883 -1027
rect 1839 -1089 1883 -1047
rect 1933 -1027 1975 -989
rect 1933 -1047 1947 -1027
rect 1967 -1047 1975 -1027
rect 1933 -1089 1975 -1047
rect 2049 -1027 2091 -989
rect 2049 -1047 2057 -1027
rect 2077 -1047 2091 -1027
rect 2049 -1089 2091 -1047
rect 2141 -1020 2186 -989
rect 2141 -1027 2185 -1020
rect 2141 -1047 2153 -1027
rect 2173 -1047 2185 -1027
rect 2141 -1089 2185 -1047
rect 340 -1294 384 -1256
rect 340 -1314 352 -1294
rect 372 -1314 384 -1294
rect 340 -1356 384 -1314
rect 434 -1294 476 -1256
rect 434 -1314 448 -1294
rect 468 -1314 476 -1294
rect 434 -1356 476 -1314
rect 553 -1294 597 -1256
rect 553 -1314 565 -1294
rect 585 -1314 597 -1294
rect 553 -1356 597 -1314
rect 647 -1294 689 -1256
rect 647 -1314 661 -1294
rect 681 -1314 689 -1294
rect 647 -1356 689 -1314
rect 761 -1294 805 -1256
rect 761 -1314 773 -1294
rect 793 -1314 805 -1294
rect 761 -1356 805 -1314
rect 855 -1294 897 -1256
rect 855 -1314 869 -1294
rect 889 -1314 897 -1294
rect 855 -1356 897 -1314
rect 971 -1294 1013 -1256
rect 971 -1314 979 -1294
rect 999 -1314 1013 -1294
rect 971 -1356 1013 -1314
rect 1063 -1287 1108 -1256
rect 1063 -1294 1107 -1287
rect 1063 -1314 1075 -1294
rect 1095 -1314 1107 -1294
rect 1063 -1356 1107 -1314
rect 1278 -1538 1322 -1500
rect 1278 -1558 1290 -1538
rect 1310 -1558 1322 -1538
rect 1278 -1600 1322 -1558
rect 1372 -1538 1414 -1500
rect 1372 -1558 1386 -1538
rect 1406 -1558 1414 -1538
rect 1372 -1600 1414 -1558
rect 1491 -1538 1535 -1500
rect 1491 -1558 1503 -1538
rect 1523 -1558 1535 -1538
rect 1491 -1600 1535 -1558
rect 1585 -1538 1627 -1500
rect 1585 -1558 1599 -1538
rect 1619 -1558 1627 -1538
rect 1585 -1600 1627 -1558
rect 1699 -1538 1743 -1500
rect 1699 -1558 1711 -1538
rect 1731 -1558 1743 -1538
rect 1699 -1600 1743 -1558
rect 1793 -1538 1835 -1500
rect 1793 -1558 1807 -1538
rect 1827 -1558 1835 -1538
rect 1793 -1600 1835 -1558
rect 1909 -1538 1951 -1500
rect 1909 -1558 1917 -1538
rect 1937 -1558 1951 -1538
rect 1909 -1600 1951 -1558
rect 2001 -1531 2046 -1500
rect 2001 -1538 2045 -1531
rect 2001 -1558 2013 -1538
rect 2033 -1558 2045 -1538
rect 2001 -1600 2045 -1558
rect 339 -1848 383 -1810
rect 339 -1868 351 -1848
rect 371 -1868 383 -1848
rect 339 -1910 383 -1868
rect 433 -1848 475 -1810
rect 433 -1868 447 -1848
rect 467 -1868 475 -1848
rect 433 -1910 475 -1868
rect 552 -1848 596 -1810
rect 552 -1868 564 -1848
rect 584 -1868 596 -1848
rect 552 -1910 596 -1868
rect 646 -1848 688 -1810
rect 646 -1868 660 -1848
rect 680 -1868 688 -1848
rect 646 -1910 688 -1868
rect 760 -1848 804 -1810
rect 760 -1868 772 -1848
rect 792 -1868 804 -1848
rect 760 -1910 804 -1868
rect 854 -1848 896 -1810
rect 854 -1868 868 -1848
rect 888 -1868 896 -1848
rect 854 -1910 896 -1868
rect 970 -1848 1012 -1810
rect 970 -1868 978 -1848
rect 998 -1868 1012 -1848
rect 970 -1910 1012 -1868
rect 1062 -1841 1107 -1810
rect 1062 -1848 1106 -1841
rect 1062 -1868 1074 -1848
rect 1094 -1868 1106 -1848
rect 1062 -1910 1106 -1868
<< ndiffc >>
rect 116 2131 134 2149
rect 118 2032 136 2050
rect 116 1944 134 1962
rect 118 1845 136 1863
rect 344 1846 364 1866
rect 447 1850 467 1870
rect 557 1846 577 1866
rect 660 1850 680 1870
rect 765 1846 785 1866
rect 868 1850 888 1870
rect 976 1850 996 1870
rect 1079 1846 1099 1866
rect 116 1715 134 1733
rect 118 1616 136 1634
rect 1282 1602 1302 1622
rect 1385 1606 1405 1626
rect 1495 1602 1515 1622
rect 1598 1606 1618 1626
rect 1703 1602 1723 1622
rect 1806 1606 1826 1626
rect 1914 1606 1934 1626
rect 2017 1602 2037 1622
rect 116 1485 134 1503
rect 118 1386 136 1404
rect 343 1292 363 1312
rect 446 1296 466 1316
rect 556 1292 576 1312
rect 659 1296 679 1316
rect 764 1292 784 1312
rect 867 1296 887 1316
rect 975 1296 995 1316
rect 1078 1292 1098 1312
rect 117 1028 135 1046
rect 1423 1010 1443 1030
rect 1526 1014 1546 1034
rect 1636 1010 1656 1030
rect 1739 1014 1759 1034
rect 1844 1010 1864 1030
rect 1947 1014 1967 1034
rect 2055 1014 2075 1034
rect 2158 1010 2178 1030
rect 119 929 137 947
rect 117 841 135 859
rect 119 742 137 760
rect 345 743 365 763
rect 448 747 468 767
rect 558 743 578 763
rect 661 747 681 767
rect 766 743 786 763
rect 869 747 889 767
rect 977 747 997 767
rect 1080 743 1100 763
rect 117 612 135 630
rect 119 513 137 531
rect 1283 499 1303 519
rect 1386 503 1406 523
rect 1496 499 1516 519
rect 1599 503 1619 523
rect 1704 499 1724 519
rect 1807 503 1827 523
rect 1915 503 1935 523
rect 2018 499 2038 519
rect 117 382 135 400
rect 119 283 137 301
rect 344 189 364 209
rect 447 193 467 213
rect 557 189 577 209
rect 660 193 680 213
rect 765 189 785 209
rect 868 193 888 213
rect 976 193 996 213
rect 1079 189 1099 209
rect 117 -75 135 -57
rect 1393 -80 1413 -60
rect 1496 -76 1516 -56
rect 1606 -80 1626 -60
rect 1709 -76 1729 -56
rect 1814 -80 1834 -60
rect 1917 -76 1937 -56
rect 2025 -76 2045 -56
rect 2128 -80 2148 -60
rect 119 -174 137 -156
rect 117 -262 135 -244
rect 119 -361 137 -343
rect 345 -360 365 -340
rect 448 -356 468 -336
rect 558 -360 578 -340
rect 661 -356 681 -336
rect 766 -360 786 -340
rect 869 -356 889 -336
rect 977 -356 997 -336
rect 1080 -360 1100 -340
rect 117 -491 135 -473
rect 119 -590 137 -572
rect 1283 -604 1303 -584
rect 1386 -600 1406 -580
rect 1496 -604 1516 -584
rect 1599 -600 1619 -580
rect 1704 -604 1724 -584
rect 1807 -600 1827 -580
rect 1915 -600 1935 -580
rect 2018 -604 2038 -584
rect 117 -721 135 -703
rect 119 -820 137 -802
rect 344 -914 364 -894
rect 447 -910 467 -890
rect 557 -914 577 -894
rect 660 -910 680 -890
rect 765 -914 785 -894
rect 868 -910 888 -890
rect 976 -910 996 -890
rect 1079 -914 1099 -894
rect 118 -1178 136 -1160
rect 1424 -1196 1444 -1176
rect 1527 -1192 1547 -1172
rect 1637 -1196 1657 -1176
rect 1740 -1192 1760 -1172
rect 1845 -1196 1865 -1176
rect 1948 -1192 1968 -1172
rect 2056 -1192 2076 -1172
rect 2159 -1196 2179 -1176
rect 120 -1277 138 -1259
rect 118 -1365 136 -1347
rect 120 -1464 138 -1446
rect 346 -1463 366 -1443
rect 449 -1459 469 -1439
rect 559 -1463 579 -1443
rect 662 -1459 682 -1439
rect 767 -1463 787 -1443
rect 870 -1459 890 -1439
rect 978 -1459 998 -1439
rect 1081 -1463 1101 -1443
rect 118 -1594 136 -1576
rect 120 -1693 138 -1675
rect 1284 -1707 1304 -1687
rect 1387 -1703 1407 -1683
rect 1497 -1707 1517 -1687
rect 1600 -1703 1620 -1683
rect 1705 -1707 1725 -1687
rect 1808 -1703 1828 -1683
rect 1916 -1703 1936 -1683
rect 2019 -1707 2039 -1687
rect 118 -1824 136 -1806
rect 120 -1923 138 -1905
rect 345 -2017 365 -1997
rect 448 -2013 468 -1993
rect 558 -2017 578 -1997
rect 661 -2013 681 -1993
rect 766 -2017 786 -1997
rect 869 -2013 889 -1993
rect 977 -2013 997 -1993
rect 1080 -2017 1100 -1997
<< pdiffc >>
rect 350 1995 370 2015
rect 446 1995 466 2015
rect 563 1995 583 2015
rect 659 1995 679 2015
rect 771 1995 791 2015
rect 867 1995 887 2015
rect 977 1995 997 2015
rect 1073 1995 1093 2015
rect 1288 1751 1308 1771
rect 1384 1751 1404 1771
rect 1501 1751 1521 1771
rect 1597 1751 1617 1771
rect 1709 1751 1729 1771
rect 1805 1751 1825 1771
rect 1915 1751 1935 1771
rect 2011 1751 2031 1771
rect 349 1441 369 1461
rect 445 1441 465 1461
rect 562 1441 582 1461
rect 658 1441 678 1461
rect 770 1441 790 1461
rect 866 1441 886 1461
rect 976 1441 996 1461
rect 1072 1441 1092 1461
rect 1429 1159 1449 1179
rect 1525 1159 1545 1179
rect 1642 1159 1662 1179
rect 1738 1159 1758 1179
rect 1850 1159 1870 1179
rect 1946 1159 1966 1179
rect 2056 1159 2076 1179
rect 2152 1159 2172 1179
rect 351 892 371 912
rect 447 892 467 912
rect 564 892 584 912
rect 660 892 680 912
rect 772 892 792 912
rect 868 892 888 912
rect 978 892 998 912
rect 1074 892 1094 912
rect 1289 648 1309 668
rect 1385 648 1405 668
rect 1502 648 1522 668
rect 1598 648 1618 668
rect 1710 648 1730 668
rect 1806 648 1826 668
rect 1916 648 1936 668
rect 2012 648 2032 668
rect 350 338 370 358
rect 446 338 466 358
rect 563 338 583 358
rect 659 338 679 358
rect 771 338 791 358
rect 867 338 887 358
rect 977 338 997 358
rect 1073 338 1093 358
rect 1399 69 1419 89
rect 1495 69 1515 89
rect 1612 69 1632 89
rect 1708 69 1728 89
rect 1820 69 1840 89
rect 1916 69 1936 89
rect 2026 69 2046 89
rect 2122 69 2142 89
rect 351 -211 371 -191
rect 447 -211 467 -191
rect 564 -211 584 -191
rect 660 -211 680 -191
rect 772 -211 792 -191
rect 868 -211 888 -191
rect 978 -211 998 -191
rect 1074 -211 1094 -191
rect 1289 -455 1309 -435
rect 1385 -455 1405 -435
rect 1502 -455 1522 -435
rect 1598 -455 1618 -435
rect 1710 -455 1730 -435
rect 1806 -455 1826 -435
rect 1916 -455 1936 -435
rect 2012 -455 2032 -435
rect 350 -765 370 -745
rect 446 -765 466 -745
rect 563 -765 583 -745
rect 659 -765 679 -745
rect 771 -765 791 -745
rect 867 -765 887 -745
rect 977 -765 997 -745
rect 1073 -765 1093 -745
rect 1430 -1047 1450 -1027
rect 1526 -1047 1546 -1027
rect 1643 -1047 1663 -1027
rect 1739 -1047 1759 -1027
rect 1851 -1047 1871 -1027
rect 1947 -1047 1967 -1027
rect 2057 -1047 2077 -1027
rect 2153 -1047 2173 -1027
rect 352 -1314 372 -1294
rect 448 -1314 468 -1294
rect 565 -1314 585 -1294
rect 661 -1314 681 -1294
rect 773 -1314 793 -1294
rect 869 -1314 889 -1294
rect 979 -1314 999 -1294
rect 1075 -1314 1095 -1294
rect 1290 -1558 1310 -1538
rect 1386 -1558 1406 -1538
rect 1503 -1558 1523 -1538
rect 1599 -1558 1619 -1538
rect 1711 -1558 1731 -1538
rect 1807 -1558 1827 -1538
rect 1917 -1558 1937 -1538
rect 2013 -1558 2033 -1538
rect 351 -1868 371 -1848
rect 447 -1868 467 -1848
rect 564 -1868 584 -1848
rect 660 -1868 680 -1848
rect 772 -1868 792 -1848
rect 868 -1868 888 -1848
rect 978 -1868 998 -1848
rect 1074 -1868 1094 -1848
<< psubdiff >>
rect 418 1779 529 1793
rect 418 1749 459 1779
rect 487 1749 529 1779
rect 418 1734 529 1749
rect 1356 1535 1467 1549
rect 1356 1505 1397 1535
rect 1425 1505 1467 1535
rect 1356 1490 1467 1505
rect 417 1225 528 1239
rect 417 1195 458 1225
rect 486 1195 528 1225
rect 417 1180 528 1195
rect 1497 943 1608 957
rect 1497 913 1538 943
rect 1566 913 1608 943
rect 1497 898 1608 913
rect 419 676 530 690
rect 419 646 460 676
rect 488 646 530 676
rect 419 631 530 646
rect 1357 432 1468 446
rect 1357 402 1398 432
rect 1426 402 1468 432
rect 1357 387 1468 402
rect 418 122 529 136
rect 418 92 459 122
rect 487 92 529 122
rect 418 78 529 92
rect 1467 -147 1578 -133
rect 1467 -177 1508 -147
rect 1536 -177 1578 -147
rect 1467 -192 1578 -177
rect 419 -427 530 -413
rect 419 -457 460 -427
rect 488 -457 530 -427
rect 419 -472 530 -457
rect 1357 -671 1468 -657
rect 1357 -701 1398 -671
rect 1426 -701 1468 -671
rect 1357 -716 1468 -701
rect 418 -981 529 -967
rect 418 -1011 459 -981
rect 487 -1011 529 -981
rect 418 -1026 529 -1011
rect 1498 -1263 1609 -1249
rect 1498 -1293 1539 -1263
rect 1567 -1293 1609 -1263
rect 1498 -1308 1609 -1293
rect 420 -1530 531 -1516
rect 420 -1560 461 -1530
rect 489 -1560 531 -1530
rect 420 -1575 531 -1560
rect 1358 -1774 1469 -1760
rect 1358 -1804 1399 -1774
rect 1427 -1804 1469 -1774
rect 1358 -1819 1469 -1804
rect 419 -2084 530 -2070
rect 419 -2114 460 -2084
rect 488 -2114 530 -2084
rect 419 -2129 530 -2114
<< nsubdiff >>
rect 419 2126 529 2140
rect 419 2096 462 2126
rect 490 2096 529 2126
rect 419 2081 529 2096
rect 1357 1882 1467 1896
rect 1357 1852 1400 1882
rect 1428 1852 1467 1882
rect 1357 1837 1467 1852
rect 418 1572 528 1586
rect 418 1542 461 1572
rect 489 1542 528 1572
rect 418 1527 528 1542
rect 1498 1290 1608 1304
rect 1498 1260 1541 1290
rect 1569 1260 1608 1290
rect 1498 1245 1608 1260
rect 420 1023 530 1037
rect 420 993 463 1023
rect 491 993 530 1023
rect 420 978 530 993
rect 1358 779 1468 793
rect 1358 749 1401 779
rect 1429 749 1468 779
rect 1358 734 1468 749
rect 419 469 529 483
rect 419 439 462 469
rect 490 439 529 469
rect 419 424 529 439
rect 1468 200 1578 214
rect 1468 170 1511 200
rect 1539 170 1578 200
rect 1468 155 1578 170
rect 420 -80 530 -66
rect 420 -110 463 -80
rect 491 -110 530 -80
rect 420 -125 530 -110
rect 1358 -324 1468 -310
rect 1358 -354 1401 -324
rect 1429 -354 1468 -324
rect 1358 -369 1468 -354
rect 419 -634 529 -620
rect 419 -664 462 -634
rect 490 -664 529 -634
rect 419 -679 529 -664
rect 1499 -916 1609 -902
rect 1499 -946 1542 -916
rect 1570 -946 1609 -916
rect 1499 -961 1609 -946
rect 421 -1183 531 -1169
rect 421 -1213 464 -1183
rect 492 -1213 531 -1183
rect 421 -1228 531 -1213
rect 1359 -1427 1469 -1413
rect 1359 -1457 1402 -1427
rect 1430 -1457 1469 -1427
rect 1359 -1472 1469 -1457
rect 420 -1737 530 -1723
rect 420 -1767 463 -1737
rect 491 -1767 530 -1737
rect 420 -1782 530 -1767
<< psubdiffcont >>
rect 459 1749 487 1779
rect 1397 1505 1425 1535
rect 458 1195 486 1225
rect 1538 913 1566 943
rect 460 646 488 676
rect 1398 402 1426 432
rect 459 92 487 122
rect 1508 -177 1536 -147
rect 460 -457 488 -427
rect 1398 -701 1426 -671
rect 459 -1011 487 -981
rect 1539 -1293 1567 -1263
rect 461 -1560 489 -1530
rect 1399 -1804 1427 -1774
rect 460 -2114 488 -2084
<< nsubdiffcont >>
rect 462 2096 490 2126
rect 1400 1852 1428 1882
rect 461 1542 489 1572
rect 1541 1260 1569 1290
rect 463 993 491 1023
rect 1401 749 1429 779
rect 462 439 490 469
rect 1511 170 1539 200
rect 463 -110 491 -80
rect 1401 -354 1429 -324
rect 462 -664 490 -634
rect 1542 -946 1570 -916
rect 464 -1213 492 -1183
rect 1402 -1457 1430 -1427
rect 463 -1767 491 -1737
<< poly >>
rect 382 2053 432 2066
rect 595 2053 645 2066
rect 803 2053 853 2066
rect 1011 2053 1061 2066
rect 382 1925 432 1953
rect 382 1905 395 1925
rect 415 1905 432 1925
rect 382 1876 432 1905
rect 595 1924 645 1953
rect 595 1900 606 1924
rect 630 1900 645 1924
rect 595 1876 645 1900
rect 803 1929 853 1953
rect 803 1905 815 1929
rect 839 1905 853 1929
rect 803 1876 853 1905
rect 1011 1927 1061 1953
rect 1011 1901 1029 1927
rect 1055 1901 1061 1927
rect 1011 1876 1061 1901
rect 382 1818 432 1834
rect 595 1818 645 1834
rect 803 1818 853 1834
rect 1011 1818 1061 1834
rect 1320 1809 1370 1822
rect 1533 1809 1583 1822
rect 1741 1809 1791 1822
rect 1949 1809 1999 1822
rect 1320 1681 1370 1709
rect 1320 1661 1333 1681
rect 1353 1661 1370 1681
rect 1320 1632 1370 1661
rect 1533 1680 1583 1709
rect 1533 1656 1544 1680
rect 1568 1656 1583 1680
rect 1533 1632 1583 1656
rect 1741 1685 1791 1709
rect 1741 1661 1753 1685
rect 1777 1661 1791 1685
rect 1741 1632 1791 1661
rect 1949 1683 1999 1709
rect 1949 1657 1967 1683
rect 1993 1657 1999 1683
rect 1949 1632 1999 1657
rect 1320 1574 1370 1590
rect 1533 1574 1583 1590
rect 1741 1574 1791 1590
rect 1949 1574 1999 1590
rect 381 1499 431 1512
rect 594 1499 644 1512
rect 802 1499 852 1512
rect 1010 1499 1060 1512
rect 381 1371 431 1399
rect 381 1351 394 1371
rect 414 1351 431 1371
rect 381 1322 431 1351
rect 594 1370 644 1399
rect 594 1346 605 1370
rect 629 1346 644 1370
rect 594 1322 644 1346
rect 802 1375 852 1399
rect 802 1351 814 1375
rect 838 1351 852 1375
rect 802 1322 852 1351
rect 1010 1373 1060 1399
rect 1010 1347 1028 1373
rect 1054 1347 1060 1373
rect 1010 1322 1060 1347
rect 381 1264 431 1280
rect 594 1264 644 1280
rect 802 1264 852 1280
rect 1010 1264 1060 1280
rect 1461 1217 1511 1230
rect 1674 1217 1724 1230
rect 1882 1217 1932 1230
rect 2090 1217 2140 1230
rect 1461 1089 1511 1117
rect 1461 1069 1474 1089
rect 1494 1069 1511 1089
rect 1461 1040 1511 1069
rect 1674 1088 1724 1117
rect 1674 1064 1685 1088
rect 1709 1064 1724 1088
rect 1674 1040 1724 1064
rect 1882 1093 1932 1117
rect 1882 1069 1894 1093
rect 1918 1069 1932 1093
rect 1882 1040 1932 1069
rect 2090 1091 2140 1117
rect 2090 1065 2108 1091
rect 2134 1065 2140 1091
rect 2090 1040 2140 1065
rect 1461 982 1511 998
rect 1674 982 1724 998
rect 1882 982 1932 998
rect 2090 982 2140 998
rect 383 950 433 963
rect 596 950 646 963
rect 804 950 854 963
rect 1012 950 1062 963
rect 383 822 433 850
rect 383 802 396 822
rect 416 802 433 822
rect 383 773 433 802
rect 596 821 646 850
rect 596 797 607 821
rect 631 797 646 821
rect 596 773 646 797
rect 804 826 854 850
rect 804 802 816 826
rect 840 802 854 826
rect 804 773 854 802
rect 1012 824 1062 850
rect 1012 798 1030 824
rect 1056 798 1062 824
rect 1012 773 1062 798
rect 383 715 433 731
rect 596 715 646 731
rect 804 715 854 731
rect 1012 715 1062 731
rect 1321 706 1371 719
rect 1534 706 1584 719
rect 1742 706 1792 719
rect 1950 706 2000 719
rect 1321 578 1371 606
rect 1321 558 1334 578
rect 1354 558 1371 578
rect 1321 529 1371 558
rect 1534 577 1584 606
rect 1534 553 1545 577
rect 1569 553 1584 577
rect 1534 529 1584 553
rect 1742 582 1792 606
rect 1742 558 1754 582
rect 1778 558 1792 582
rect 1742 529 1792 558
rect 1950 580 2000 606
rect 1950 554 1968 580
rect 1994 554 2000 580
rect 1950 529 2000 554
rect 1321 471 1371 487
rect 1534 471 1584 487
rect 1742 471 1792 487
rect 1950 471 2000 487
rect 382 396 432 409
rect 595 396 645 409
rect 803 396 853 409
rect 1011 396 1061 409
rect 382 268 432 296
rect 382 248 395 268
rect 415 248 432 268
rect 382 219 432 248
rect 595 267 645 296
rect 595 243 606 267
rect 630 243 645 267
rect 595 219 645 243
rect 803 272 853 296
rect 803 248 815 272
rect 839 248 853 272
rect 803 219 853 248
rect 1011 270 1061 296
rect 1011 244 1029 270
rect 1055 244 1061 270
rect 1011 219 1061 244
rect 382 161 432 177
rect 595 161 645 177
rect 803 161 853 177
rect 1011 161 1061 177
rect 1431 127 1481 140
rect 1644 127 1694 140
rect 1852 127 1902 140
rect 2060 127 2110 140
rect 1431 -1 1481 27
rect 1431 -21 1444 -1
rect 1464 -21 1481 -1
rect 1431 -50 1481 -21
rect 1644 -2 1694 27
rect 1644 -26 1655 -2
rect 1679 -26 1694 -2
rect 1644 -50 1694 -26
rect 1852 3 1902 27
rect 1852 -21 1864 3
rect 1888 -21 1902 3
rect 1852 -50 1902 -21
rect 2060 1 2110 27
rect 2060 -25 2078 1
rect 2104 -25 2110 1
rect 2060 -50 2110 -25
rect 1431 -108 1481 -92
rect 1644 -108 1694 -92
rect 1852 -108 1902 -92
rect 2060 -108 2110 -92
rect 383 -153 433 -140
rect 596 -153 646 -140
rect 804 -153 854 -140
rect 1012 -153 1062 -140
rect 383 -281 433 -253
rect 383 -301 396 -281
rect 416 -301 433 -281
rect 383 -330 433 -301
rect 596 -282 646 -253
rect 596 -306 607 -282
rect 631 -306 646 -282
rect 596 -330 646 -306
rect 804 -277 854 -253
rect 804 -301 816 -277
rect 840 -301 854 -277
rect 804 -330 854 -301
rect 1012 -279 1062 -253
rect 1012 -305 1030 -279
rect 1056 -305 1062 -279
rect 1012 -330 1062 -305
rect 383 -388 433 -372
rect 596 -388 646 -372
rect 804 -388 854 -372
rect 1012 -388 1062 -372
rect 1321 -397 1371 -384
rect 1534 -397 1584 -384
rect 1742 -397 1792 -384
rect 1950 -397 2000 -384
rect 1321 -525 1371 -497
rect 1321 -545 1334 -525
rect 1354 -545 1371 -525
rect 1321 -574 1371 -545
rect 1534 -526 1584 -497
rect 1534 -550 1545 -526
rect 1569 -550 1584 -526
rect 1534 -574 1584 -550
rect 1742 -521 1792 -497
rect 1742 -545 1754 -521
rect 1778 -545 1792 -521
rect 1742 -574 1792 -545
rect 1950 -523 2000 -497
rect 1950 -549 1968 -523
rect 1994 -549 2000 -523
rect 1950 -574 2000 -549
rect 1321 -632 1371 -616
rect 1534 -632 1584 -616
rect 1742 -632 1792 -616
rect 1950 -632 2000 -616
rect 382 -707 432 -694
rect 595 -707 645 -694
rect 803 -707 853 -694
rect 1011 -707 1061 -694
rect 382 -835 432 -807
rect 382 -855 395 -835
rect 415 -855 432 -835
rect 382 -884 432 -855
rect 595 -836 645 -807
rect 595 -860 606 -836
rect 630 -860 645 -836
rect 595 -884 645 -860
rect 803 -831 853 -807
rect 803 -855 815 -831
rect 839 -855 853 -831
rect 803 -884 853 -855
rect 1011 -833 1061 -807
rect 1011 -859 1029 -833
rect 1055 -859 1061 -833
rect 1011 -884 1061 -859
rect 382 -942 432 -926
rect 595 -942 645 -926
rect 803 -942 853 -926
rect 1011 -942 1061 -926
rect 1462 -989 1512 -976
rect 1675 -989 1725 -976
rect 1883 -989 1933 -976
rect 2091 -989 2141 -976
rect 1462 -1117 1512 -1089
rect 1462 -1137 1475 -1117
rect 1495 -1137 1512 -1117
rect 1462 -1166 1512 -1137
rect 1675 -1118 1725 -1089
rect 1675 -1142 1686 -1118
rect 1710 -1142 1725 -1118
rect 1675 -1166 1725 -1142
rect 1883 -1113 1933 -1089
rect 1883 -1137 1895 -1113
rect 1919 -1137 1933 -1113
rect 1883 -1166 1933 -1137
rect 2091 -1115 2141 -1089
rect 2091 -1141 2109 -1115
rect 2135 -1141 2141 -1115
rect 2091 -1166 2141 -1141
rect 1462 -1224 1512 -1208
rect 1675 -1224 1725 -1208
rect 1883 -1224 1933 -1208
rect 2091 -1224 2141 -1208
rect 384 -1256 434 -1243
rect 597 -1256 647 -1243
rect 805 -1256 855 -1243
rect 1013 -1256 1063 -1243
rect 384 -1384 434 -1356
rect 384 -1404 397 -1384
rect 417 -1404 434 -1384
rect 384 -1433 434 -1404
rect 597 -1385 647 -1356
rect 597 -1409 608 -1385
rect 632 -1409 647 -1385
rect 597 -1433 647 -1409
rect 805 -1380 855 -1356
rect 805 -1404 817 -1380
rect 841 -1404 855 -1380
rect 805 -1433 855 -1404
rect 1013 -1382 1063 -1356
rect 1013 -1408 1031 -1382
rect 1057 -1408 1063 -1382
rect 1013 -1433 1063 -1408
rect 384 -1491 434 -1475
rect 597 -1491 647 -1475
rect 805 -1491 855 -1475
rect 1013 -1491 1063 -1475
rect 1322 -1500 1372 -1487
rect 1535 -1500 1585 -1487
rect 1743 -1500 1793 -1487
rect 1951 -1500 2001 -1487
rect 1322 -1628 1372 -1600
rect 1322 -1648 1335 -1628
rect 1355 -1648 1372 -1628
rect 1322 -1677 1372 -1648
rect 1535 -1629 1585 -1600
rect 1535 -1653 1546 -1629
rect 1570 -1653 1585 -1629
rect 1535 -1677 1585 -1653
rect 1743 -1624 1793 -1600
rect 1743 -1648 1755 -1624
rect 1779 -1648 1793 -1624
rect 1743 -1677 1793 -1648
rect 1951 -1626 2001 -1600
rect 1951 -1652 1969 -1626
rect 1995 -1652 2001 -1626
rect 1951 -1677 2001 -1652
rect 1322 -1735 1372 -1719
rect 1535 -1735 1585 -1719
rect 1743 -1735 1793 -1719
rect 1951 -1735 2001 -1719
rect 383 -1810 433 -1797
rect 596 -1810 646 -1797
rect 804 -1810 854 -1797
rect 1012 -1810 1062 -1797
rect 383 -1938 433 -1910
rect 383 -1958 396 -1938
rect 416 -1958 433 -1938
rect 383 -1987 433 -1958
rect 596 -1939 646 -1910
rect 596 -1963 607 -1939
rect 631 -1963 646 -1939
rect 596 -1987 646 -1963
rect 804 -1934 854 -1910
rect 804 -1958 816 -1934
rect 840 -1958 854 -1934
rect 804 -1987 854 -1958
rect 1012 -1936 1062 -1910
rect 1012 -1962 1030 -1936
rect 1056 -1962 1062 -1936
rect 1012 -1987 1062 -1962
rect 383 -2045 433 -2029
rect 596 -2045 646 -2029
rect 804 -2045 854 -2029
rect 1012 -2045 1062 -2029
<< polycont >>
rect 395 1905 415 1925
rect 606 1900 630 1924
rect 815 1905 839 1929
rect 1029 1901 1055 1927
rect 1333 1661 1353 1681
rect 1544 1656 1568 1680
rect 1753 1661 1777 1685
rect 1967 1657 1993 1683
rect 394 1351 414 1371
rect 605 1346 629 1370
rect 814 1351 838 1375
rect 1028 1347 1054 1373
rect 1474 1069 1494 1089
rect 1685 1064 1709 1088
rect 1894 1069 1918 1093
rect 2108 1065 2134 1091
rect 396 802 416 822
rect 607 797 631 821
rect 816 802 840 826
rect 1030 798 1056 824
rect 1334 558 1354 578
rect 1545 553 1569 577
rect 1754 558 1778 582
rect 1968 554 1994 580
rect 395 248 415 268
rect 606 243 630 267
rect 815 248 839 272
rect 1029 244 1055 270
rect 1444 -21 1464 -1
rect 1655 -26 1679 -2
rect 1864 -21 1888 3
rect 2078 -25 2104 1
rect 396 -301 416 -281
rect 607 -306 631 -282
rect 816 -301 840 -277
rect 1030 -305 1056 -279
rect 1334 -545 1354 -525
rect 1545 -550 1569 -526
rect 1754 -545 1778 -521
rect 1968 -549 1994 -523
rect 395 -855 415 -835
rect 606 -860 630 -836
rect 815 -855 839 -831
rect 1029 -859 1055 -833
rect 1475 -1137 1495 -1117
rect 1686 -1142 1710 -1118
rect 1895 -1137 1919 -1113
rect 2109 -1141 2135 -1115
rect 397 -1404 417 -1384
rect 608 -1409 632 -1385
rect 817 -1404 841 -1380
rect 1031 -1408 1057 -1382
rect 1335 -1648 1355 -1628
rect 1546 -1653 1570 -1629
rect 1755 -1648 1779 -1624
rect 1969 -1652 1995 -1626
rect 396 -1958 416 -1938
rect 607 -1963 631 -1939
rect 816 -1958 840 -1934
rect 1030 -1962 1056 -1936
<< ndiffres >>
rect 95 2149 152 2168
rect 95 2146 116 2149
rect 1 2131 116 2146
rect 134 2131 152 2149
rect 1 2108 152 2131
rect 1 2072 43 2108
rect 0 2071 100 2072
rect 0 2050 156 2071
rect 0 2032 118 2050
rect 136 2032 156 2050
rect 0 2028 156 2032
rect 95 2012 156 2028
rect 95 1962 152 1981
rect 95 1959 116 1962
rect 1 1944 116 1959
rect 134 1944 152 1962
rect 1 1921 152 1944
rect 1 1885 43 1921
rect 0 1884 100 1885
rect 0 1863 156 1884
rect 0 1845 118 1863
rect 136 1845 156 1863
rect 0 1841 156 1845
rect 95 1825 156 1841
rect 95 1733 152 1752
rect 95 1730 116 1733
rect 1 1715 116 1730
rect 134 1715 152 1733
rect 1 1692 152 1715
rect 1 1656 43 1692
rect 0 1655 100 1656
rect 0 1634 156 1655
rect 0 1616 118 1634
rect 136 1616 156 1634
rect 0 1612 156 1616
rect 95 1596 156 1612
rect 95 1503 152 1522
rect 95 1500 116 1503
rect 1 1485 116 1500
rect 134 1485 152 1503
rect 1 1462 152 1485
rect 1 1426 43 1462
rect 0 1425 100 1426
rect 0 1404 156 1425
rect 0 1386 118 1404
rect 136 1386 156 1404
rect 0 1382 156 1386
rect 95 1366 156 1382
rect 96 1046 153 1065
rect 96 1043 117 1046
rect 2 1028 117 1043
rect 135 1028 153 1046
rect 2 1005 153 1028
rect 2 969 44 1005
rect 1 968 101 969
rect 1 947 157 968
rect 1 929 119 947
rect 137 929 157 947
rect 1 925 157 929
rect 96 909 157 925
rect 96 859 153 878
rect 96 856 117 859
rect 2 841 117 856
rect 135 841 153 859
rect 2 818 153 841
rect 2 782 44 818
rect 1 781 101 782
rect 1 760 157 781
rect 1 742 119 760
rect 137 742 157 760
rect 1 738 157 742
rect 96 722 157 738
rect 96 630 153 649
rect 96 627 117 630
rect 2 612 117 627
rect 135 612 153 630
rect 2 589 153 612
rect 2 553 44 589
rect 1 552 101 553
rect 1 531 157 552
rect 1 513 119 531
rect 137 513 157 531
rect 1 509 157 513
rect 96 493 157 509
rect 96 400 153 419
rect 96 397 117 400
rect 2 382 117 397
rect 135 382 153 400
rect 2 359 153 382
rect 2 323 44 359
rect 1 322 101 323
rect 1 301 157 322
rect 1 283 119 301
rect 137 283 157 301
rect 1 279 157 283
rect 96 263 157 279
rect 96 -57 153 -38
rect 96 -60 117 -57
rect 2 -75 117 -60
rect 135 -75 153 -57
rect 2 -98 153 -75
rect 2 -134 44 -98
rect 1 -135 101 -134
rect 1 -156 157 -135
rect 1 -174 119 -156
rect 137 -174 157 -156
rect 1 -178 157 -174
rect 96 -194 157 -178
rect 96 -244 153 -225
rect 96 -247 117 -244
rect 2 -262 117 -247
rect 135 -262 153 -244
rect 2 -285 153 -262
rect 2 -321 44 -285
rect 1 -322 101 -321
rect 1 -343 157 -322
rect 1 -361 119 -343
rect 137 -361 157 -343
rect 1 -365 157 -361
rect 96 -381 157 -365
rect 96 -473 153 -454
rect 96 -476 117 -473
rect 2 -491 117 -476
rect 135 -491 153 -473
rect 2 -514 153 -491
rect 2 -550 44 -514
rect 1 -551 101 -550
rect 1 -572 157 -551
rect 1 -590 119 -572
rect 137 -590 157 -572
rect 1 -594 157 -590
rect 96 -610 157 -594
rect 96 -703 153 -684
rect 96 -706 117 -703
rect 2 -721 117 -706
rect 135 -721 153 -703
rect 2 -744 153 -721
rect 2 -780 44 -744
rect 1 -781 101 -780
rect 1 -802 157 -781
rect 1 -820 119 -802
rect 137 -820 157 -802
rect 1 -824 157 -820
rect 96 -840 157 -824
rect 97 -1160 154 -1141
rect 97 -1163 118 -1160
rect 3 -1178 118 -1163
rect 136 -1178 154 -1160
rect 3 -1201 154 -1178
rect 3 -1237 45 -1201
rect 2 -1238 102 -1237
rect 2 -1259 158 -1238
rect 2 -1277 120 -1259
rect 138 -1277 158 -1259
rect 2 -1281 158 -1277
rect 97 -1297 158 -1281
rect 97 -1347 154 -1328
rect 97 -1350 118 -1347
rect 3 -1365 118 -1350
rect 136 -1365 154 -1347
rect 3 -1388 154 -1365
rect 3 -1424 45 -1388
rect 2 -1425 102 -1424
rect 2 -1446 158 -1425
rect 2 -1464 120 -1446
rect 138 -1464 158 -1446
rect 2 -1468 158 -1464
rect 97 -1484 158 -1468
rect 97 -1576 154 -1557
rect 97 -1579 118 -1576
rect 3 -1594 118 -1579
rect 136 -1594 154 -1576
rect 3 -1617 154 -1594
rect 3 -1653 45 -1617
rect 2 -1654 102 -1653
rect 2 -1675 158 -1654
rect 2 -1693 120 -1675
rect 138 -1693 158 -1675
rect 2 -1697 158 -1693
rect 97 -1713 158 -1697
rect 97 -1806 154 -1787
rect 97 -1809 118 -1806
rect 3 -1824 118 -1809
rect 136 -1824 154 -1806
rect 3 -1847 154 -1824
rect 3 -1883 45 -1847
rect 2 -1884 102 -1883
rect 2 -1905 158 -1884
rect 2 -1923 120 -1905
rect 138 -1923 158 -1905
rect 2 -1927 158 -1923
rect 97 -1943 158 -1927
<< locali >>
rect 105 2151 144 2208
rect 105 2149 153 2151
rect 105 2131 116 2149
rect 134 2131 153 2149
rect 105 2122 153 2131
rect 106 2121 153 2122
rect 419 2126 529 2140
rect 419 2123 462 2126
rect 419 2118 423 2123
rect 341 2096 423 2118
rect 452 2096 462 2123
rect 490 2099 497 2126
rect 526 2118 529 2126
rect 526 2099 591 2118
rect 490 2096 591 2099
rect 341 2094 591 2096
rect 109 2058 146 2059
rect 105 2055 146 2058
rect 105 2050 147 2055
rect 105 2032 118 2050
rect 136 2032 147 2050
rect 105 2018 147 2032
rect 185 2018 232 2022
rect 105 2012 232 2018
rect 105 1983 193 2012
rect 222 1983 232 2012
rect 341 2015 378 2094
rect 419 2081 529 2094
rect 493 2025 524 2026
rect 341 1995 350 2015
rect 370 1995 378 2015
rect 341 1985 378 1995
rect 437 2015 524 2025
rect 437 1995 446 2015
rect 466 1995 524 2015
rect 437 1986 524 1995
rect 437 1985 474 1986
rect 105 1979 232 1983
rect 105 1962 144 1979
rect 185 1978 232 1979
rect 105 1944 116 1962
rect 134 1944 144 1962
rect 105 1935 144 1944
rect 106 1934 143 1935
rect 493 1933 524 1986
rect 554 2015 591 2094
rect 762 2091 1155 2111
rect 1175 2091 1178 2111
rect 762 2086 1178 2091
rect 762 2085 1103 2086
rect 706 2025 737 2026
rect 554 1995 563 2015
rect 583 1995 591 2015
rect 554 1985 591 1995
rect 650 2018 737 2025
rect 650 2015 711 2018
rect 650 1995 659 2015
rect 679 1998 711 2015
rect 732 1998 737 2018
rect 679 1995 737 1998
rect 650 1988 737 1995
rect 762 2015 799 2085
rect 1065 2084 1102 2085
rect 914 2025 950 2026
rect 762 1995 771 2015
rect 791 1995 799 2015
rect 650 1986 706 1988
rect 650 1985 687 1986
rect 762 1985 799 1995
rect 858 2015 1006 2025
rect 1106 2022 1202 2024
rect 858 1995 867 2015
rect 887 1995 977 2015
rect 997 1995 1006 2015
rect 858 1986 1006 1995
rect 1064 2015 1202 2022
rect 1064 1995 1073 2015
rect 1093 1995 1202 2015
rect 1064 1986 1202 1995
rect 858 1985 895 1986
rect 914 1934 950 1986
rect 969 1985 1006 1986
rect 1065 1985 1102 1986
rect 385 1932 426 1933
rect 277 1925 426 1932
rect 277 1905 395 1925
rect 415 1905 426 1925
rect 277 1897 426 1905
rect 493 1929 852 1933
rect 493 1924 815 1929
rect 493 1900 606 1924
rect 630 1905 815 1924
rect 839 1905 852 1929
rect 630 1900 852 1905
rect 493 1897 852 1900
rect 914 1897 949 1934
rect 1017 1931 1117 1934
rect 1017 1927 1084 1931
rect 1017 1901 1029 1927
rect 1055 1905 1084 1927
rect 1110 1905 1117 1931
rect 1055 1901 1117 1905
rect 1017 1897 1117 1901
rect 493 1876 524 1897
rect 914 1876 950 1897
rect 336 1875 373 1876
rect 110 1872 144 1873
rect 109 1863 146 1872
rect 109 1845 118 1863
rect 136 1845 146 1863
rect 109 1835 146 1845
rect 335 1866 373 1875
rect 335 1846 344 1866
rect 364 1846 373 1866
rect 335 1838 373 1846
rect 439 1870 524 1876
rect 549 1875 586 1876
rect 439 1850 447 1870
rect 467 1850 524 1870
rect 439 1842 524 1850
rect 548 1866 586 1875
rect 548 1846 557 1866
rect 577 1846 586 1866
rect 439 1841 475 1842
rect 548 1838 586 1846
rect 652 1870 737 1876
rect 757 1875 794 1876
rect 652 1850 660 1870
rect 680 1869 737 1870
rect 680 1850 709 1869
rect 652 1849 709 1850
rect 730 1849 737 1869
rect 652 1842 737 1849
rect 756 1866 794 1875
rect 756 1846 765 1866
rect 785 1846 794 1866
rect 652 1841 688 1842
rect 756 1838 794 1846
rect 860 1870 1004 1876
rect 860 1850 868 1870
rect 888 1869 976 1870
rect 888 1850 919 1869
rect 860 1849 919 1850
rect 944 1850 976 1869
rect 996 1850 1004 1870
rect 944 1849 1004 1850
rect 860 1842 1004 1849
rect 860 1841 896 1842
rect 968 1841 1004 1842
rect 1070 1875 1107 1876
rect 1070 1874 1108 1875
rect 1070 1866 1134 1874
rect 1070 1846 1079 1866
rect 1099 1852 1134 1866
rect 1154 1852 1157 1872
rect 1099 1847 1157 1852
rect 1099 1846 1134 1847
rect 110 1807 144 1835
rect 336 1809 373 1838
rect 337 1807 373 1809
rect 549 1807 586 1838
rect 110 1806 282 1807
rect 110 1774 296 1806
rect 337 1785 586 1807
rect 757 1806 794 1838
rect 1070 1834 1134 1846
rect 1174 1808 1201 1986
rect 1357 1882 1467 1896
rect 1357 1879 1400 1882
rect 1357 1874 1361 1879
rect 1033 1806 1201 1808
rect 757 1800 1201 1806
rect 110 1742 144 1774
rect 106 1733 144 1742
rect 106 1715 116 1733
rect 134 1715 144 1733
rect 106 1709 144 1715
rect 262 1711 296 1774
rect 418 1779 529 1785
rect 418 1771 459 1779
rect 418 1751 426 1771
rect 445 1751 459 1771
rect 418 1749 459 1751
rect 487 1771 529 1779
rect 487 1751 503 1771
rect 522 1751 529 1771
rect 487 1749 529 1751
rect 418 1734 529 1749
rect 756 1780 1201 1800
rect 756 1711 794 1780
rect 1033 1779 1201 1780
rect 1279 1852 1361 1874
rect 1390 1852 1400 1879
rect 1428 1855 1435 1882
rect 1464 1874 1467 1882
rect 1464 1855 1529 1874
rect 1428 1852 1529 1855
rect 1279 1850 1529 1852
rect 1279 1771 1316 1850
rect 1357 1837 1467 1850
rect 1431 1781 1462 1782
rect 1279 1751 1288 1771
rect 1308 1751 1316 1771
rect 1279 1741 1316 1751
rect 1375 1771 1462 1781
rect 1375 1751 1384 1771
rect 1404 1751 1462 1771
rect 1375 1742 1462 1751
rect 1375 1741 1412 1742
rect 106 1705 143 1709
rect 262 1700 794 1711
rect 261 1684 794 1700
rect 1431 1689 1462 1742
rect 1492 1771 1529 1850
rect 1700 1847 2093 1867
rect 2113 1847 2116 1867
rect 1700 1842 2116 1847
rect 1700 1841 2041 1842
rect 1644 1781 1675 1782
rect 1492 1751 1501 1771
rect 1521 1751 1529 1771
rect 1492 1741 1529 1751
rect 1588 1774 1675 1781
rect 1588 1771 1649 1774
rect 1588 1751 1597 1771
rect 1617 1754 1649 1771
rect 1670 1754 1675 1774
rect 1617 1751 1675 1754
rect 1588 1744 1675 1751
rect 1700 1771 1737 1841
rect 2003 1840 2040 1841
rect 1852 1781 1888 1782
rect 1700 1751 1709 1771
rect 1729 1751 1737 1771
rect 1588 1742 1644 1744
rect 1588 1741 1625 1742
rect 1700 1741 1737 1751
rect 1796 1771 1944 1781
rect 2044 1778 2140 1780
rect 1796 1751 1805 1771
rect 1825 1751 1915 1771
rect 1935 1751 1944 1771
rect 1796 1742 1944 1751
rect 2002 1771 2140 1778
rect 2002 1751 2011 1771
rect 2031 1751 2140 1771
rect 2002 1742 2140 1751
rect 1796 1741 1833 1742
rect 1852 1690 1888 1742
rect 1907 1741 1944 1742
rect 2003 1741 2040 1742
rect 1323 1688 1364 1689
rect 261 1683 775 1684
rect 1215 1681 1364 1688
rect 1215 1661 1333 1681
rect 1353 1661 1364 1681
rect 1215 1653 1364 1661
rect 1431 1685 1790 1689
rect 1431 1680 1753 1685
rect 1431 1656 1544 1680
rect 1568 1661 1753 1680
rect 1777 1661 1790 1685
rect 1568 1656 1790 1661
rect 1431 1653 1790 1656
rect 1852 1653 1887 1690
rect 1955 1687 2055 1690
rect 1955 1683 2022 1687
rect 1955 1657 1967 1683
rect 1993 1661 2022 1683
rect 2048 1661 2055 1687
rect 1993 1657 2055 1661
rect 1955 1653 2055 1657
rect 109 1642 146 1643
rect 107 1634 147 1642
rect 107 1616 118 1634
rect 136 1616 147 1634
rect 1431 1632 1462 1653
rect 1852 1632 1888 1653
rect 1274 1631 1311 1632
rect 107 1568 147 1616
rect 1273 1622 1311 1631
rect 1273 1602 1282 1622
rect 1302 1602 1311 1622
rect 1273 1594 1311 1602
rect 1377 1626 1462 1632
rect 1487 1631 1524 1632
rect 1377 1606 1385 1626
rect 1405 1606 1462 1626
rect 1377 1598 1462 1606
rect 1486 1622 1524 1631
rect 1486 1602 1495 1622
rect 1515 1602 1524 1622
rect 1377 1597 1413 1598
rect 1486 1594 1524 1602
rect 1590 1626 1675 1632
rect 1695 1631 1732 1632
rect 1590 1606 1598 1626
rect 1618 1625 1675 1626
rect 1618 1606 1647 1625
rect 1590 1605 1647 1606
rect 1668 1605 1675 1625
rect 1590 1598 1675 1605
rect 1694 1622 1732 1631
rect 1694 1602 1703 1622
rect 1723 1602 1732 1622
rect 1590 1597 1626 1598
rect 1694 1594 1732 1602
rect 1798 1626 1942 1632
rect 1798 1606 1806 1626
rect 1826 1609 1862 1626
rect 1882 1609 1914 1626
rect 1826 1606 1914 1609
rect 1934 1606 1942 1626
rect 1798 1598 1942 1606
rect 1798 1597 1834 1598
rect 1906 1597 1942 1598
rect 2008 1631 2045 1632
rect 2008 1630 2046 1631
rect 2008 1622 2072 1630
rect 2008 1602 2017 1622
rect 2037 1608 2072 1622
rect 2092 1608 2095 1628
rect 2037 1603 2095 1608
rect 2037 1602 2072 1603
rect 418 1572 528 1586
rect 418 1569 461 1572
rect 107 1561 232 1568
rect 418 1564 422 1569
rect 107 1542 199 1561
rect 224 1542 232 1561
rect 107 1532 232 1542
rect 340 1542 422 1564
rect 451 1542 461 1569
rect 489 1545 496 1572
rect 525 1564 528 1572
rect 1274 1565 1311 1594
rect 525 1545 590 1564
rect 1275 1563 1311 1565
rect 1487 1563 1524 1594
rect 1695 1567 1732 1594
rect 2008 1590 2072 1602
rect 489 1542 590 1545
rect 340 1540 590 1542
rect 107 1512 147 1532
rect 106 1503 147 1512
rect 106 1485 116 1503
rect 134 1485 147 1503
rect 106 1476 147 1485
rect 106 1475 143 1476
rect 340 1461 377 1540
rect 418 1527 528 1540
rect 492 1471 523 1472
rect 340 1441 349 1461
rect 369 1441 377 1461
rect 340 1431 377 1441
rect 436 1461 523 1471
rect 436 1441 445 1461
rect 465 1441 523 1461
rect 436 1432 523 1441
rect 436 1431 473 1432
rect 109 1409 146 1413
rect 106 1404 146 1409
rect 106 1386 118 1404
rect 136 1386 146 1404
rect 106 1206 146 1386
rect 492 1379 523 1432
rect 553 1461 590 1540
rect 761 1537 1154 1557
rect 1174 1537 1177 1557
rect 1275 1541 1524 1563
rect 1693 1562 1734 1567
rect 2112 1564 2139 1742
rect 1971 1562 2139 1564
rect 1693 1556 2139 1562
rect 761 1532 1177 1537
rect 1356 1535 1467 1541
rect 761 1531 1102 1532
rect 705 1471 736 1472
rect 553 1441 562 1461
rect 582 1441 590 1461
rect 553 1431 590 1441
rect 649 1464 736 1471
rect 649 1461 710 1464
rect 649 1441 658 1461
rect 678 1444 710 1461
rect 731 1444 736 1464
rect 678 1441 736 1444
rect 649 1434 736 1441
rect 761 1461 798 1531
rect 1064 1530 1101 1531
rect 1356 1527 1397 1535
rect 1356 1507 1364 1527
rect 1383 1507 1397 1527
rect 1356 1505 1397 1507
rect 1425 1527 1467 1535
rect 1425 1507 1441 1527
rect 1460 1507 1467 1527
rect 1693 1534 1699 1556
rect 1725 1536 2139 1556
rect 1725 1534 1734 1536
rect 1971 1535 2139 1536
rect 1693 1525 1734 1534
rect 1425 1505 1467 1507
rect 1356 1490 1467 1505
rect 913 1471 949 1472
rect 761 1441 770 1461
rect 790 1441 798 1461
rect 649 1432 705 1434
rect 649 1431 686 1432
rect 761 1431 798 1441
rect 857 1461 1005 1471
rect 1105 1468 1201 1470
rect 857 1441 866 1461
rect 886 1441 976 1461
rect 996 1441 1005 1461
rect 857 1432 1005 1441
rect 1063 1461 1201 1468
rect 1063 1441 1072 1461
rect 1092 1441 1201 1461
rect 1063 1432 1201 1441
rect 857 1431 894 1432
rect 913 1380 949 1432
rect 968 1431 1005 1432
rect 1064 1431 1101 1432
rect 384 1378 425 1379
rect 276 1371 425 1378
rect 276 1351 394 1371
rect 414 1351 425 1371
rect 276 1343 425 1351
rect 492 1375 851 1379
rect 492 1370 814 1375
rect 492 1346 605 1370
rect 629 1351 814 1370
rect 838 1351 851 1375
rect 629 1346 851 1351
rect 492 1343 851 1346
rect 913 1343 948 1380
rect 1016 1377 1116 1380
rect 1016 1373 1083 1377
rect 1016 1347 1028 1373
rect 1054 1351 1083 1373
rect 1109 1351 1116 1377
rect 1054 1347 1116 1351
rect 1016 1343 1116 1347
rect 492 1322 523 1343
rect 913 1322 949 1343
rect 335 1321 372 1322
rect 334 1312 372 1321
rect 334 1292 343 1312
rect 363 1292 372 1312
rect 334 1284 372 1292
rect 438 1316 523 1322
rect 548 1321 585 1322
rect 438 1296 446 1316
rect 466 1296 523 1316
rect 438 1288 523 1296
rect 547 1312 585 1321
rect 547 1292 556 1312
rect 576 1292 585 1312
rect 438 1287 474 1288
rect 547 1284 585 1292
rect 651 1316 736 1322
rect 756 1321 793 1322
rect 651 1296 659 1316
rect 679 1315 736 1316
rect 679 1296 708 1315
rect 651 1295 708 1296
rect 729 1295 736 1315
rect 651 1288 736 1295
rect 755 1312 793 1321
rect 755 1292 764 1312
rect 784 1292 793 1312
rect 651 1287 687 1288
rect 755 1284 793 1292
rect 859 1316 1003 1322
rect 859 1296 867 1316
rect 887 1313 975 1316
rect 887 1296 918 1313
rect 859 1293 918 1296
rect 941 1296 975 1313
rect 995 1296 1003 1316
rect 941 1293 1003 1296
rect 859 1288 1003 1293
rect 859 1287 895 1288
rect 967 1287 1003 1288
rect 1069 1321 1106 1322
rect 1069 1320 1107 1321
rect 1069 1312 1133 1320
rect 1069 1292 1078 1312
rect 1098 1298 1133 1312
rect 1153 1298 1156 1318
rect 1098 1293 1156 1298
rect 1098 1292 1133 1293
rect 335 1255 372 1284
rect 336 1253 372 1255
rect 548 1253 585 1284
rect 336 1231 585 1253
rect 756 1252 793 1284
rect 1069 1280 1133 1292
rect 1173 1254 1200 1432
rect 1498 1290 1608 1304
rect 1498 1287 1541 1290
rect 1498 1282 1502 1287
rect 1032 1252 1200 1254
rect 756 1249 1200 1252
rect 417 1225 528 1231
rect 417 1217 458 1225
rect 106 1162 145 1206
rect 417 1197 425 1217
rect 444 1197 458 1217
rect 417 1195 458 1197
rect 486 1217 528 1225
rect 486 1197 502 1217
rect 521 1197 528 1217
rect 486 1195 528 1197
rect 417 1180 528 1195
rect 754 1226 1200 1249
rect 106 1138 146 1162
rect 446 1138 493 1140
rect 754 1138 792 1226
rect 1032 1225 1200 1226
rect 1420 1260 1502 1282
rect 1531 1260 1541 1287
rect 1569 1263 1576 1290
rect 1605 1282 1608 1290
rect 1605 1263 1670 1282
rect 1569 1260 1670 1263
rect 1420 1258 1670 1260
rect 1420 1179 1457 1258
rect 1498 1245 1608 1258
rect 1572 1189 1603 1190
rect 1420 1159 1429 1179
rect 1449 1159 1457 1179
rect 1420 1149 1457 1159
rect 1516 1179 1603 1189
rect 1516 1159 1525 1179
rect 1545 1159 1603 1179
rect 1516 1150 1603 1159
rect 1516 1149 1553 1150
rect 106 1105 792 1138
rect 106 1048 145 1105
rect 754 1103 792 1105
rect 1572 1097 1603 1150
rect 1633 1179 1670 1258
rect 1841 1271 2234 1275
rect 1841 1254 1860 1271
rect 1880 1255 2234 1271
rect 2254 1255 2257 1275
rect 1880 1254 2257 1255
rect 1841 1250 2257 1254
rect 1841 1249 2182 1250
rect 1785 1189 1816 1190
rect 1633 1159 1642 1179
rect 1662 1159 1670 1179
rect 1633 1149 1670 1159
rect 1729 1182 1816 1189
rect 1729 1179 1790 1182
rect 1729 1159 1738 1179
rect 1758 1162 1790 1179
rect 1811 1162 1816 1182
rect 1758 1159 1816 1162
rect 1729 1152 1816 1159
rect 1841 1179 1878 1249
rect 2144 1248 2181 1249
rect 1993 1189 2029 1190
rect 1841 1159 1850 1179
rect 1870 1159 1878 1179
rect 1729 1150 1785 1152
rect 1729 1149 1766 1150
rect 1841 1149 1878 1159
rect 1937 1179 2085 1189
rect 2185 1186 2281 1188
rect 1937 1159 1946 1179
rect 1966 1159 2056 1179
rect 2076 1159 2085 1179
rect 1937 1150 2085 1159
rect 2143 1179 2281 1186
rect 2143 1159 2152 1179
rect 2172 1159 2281 1179
rect 2143 1150 2281 1159
rect 1937 1149 1974 1150
rect 1993 1098 2029 1150
rect 2048 1149 2085 1150
rect 2144 1149 2181 1150
rect 1464 1096 1505 1097
rect 1356 1089 1505 1096
rect 1356 1069 1474 1089
rect 1494 1069 1505 1089
rect 1356 1061 1505 1069
rect 1572 1093 1931 1097
rect 1572 1088 1894 1093
rect 1572 1064 1685 1088
rect 1709 1069 1894 1088
rect 1918 1069 1931 1093
rect 1709 1064 1931 1069
rect 1572 1061 1931 1064
rect 1993 1061 2028 1098
rect 2096 1095 2196 1098
rect 2096 1091 2163 1095
rect 2096 1065 2108 1091
rect 2134 1069 2163 1091
rect 2189 1069 2196 1095
rect 2134 1065 2196 1069
rect 2096 1061 2196 1065
rect 106 1046 154 1048
rect 106 1028 117 1046
rect 135 1028 154 1046
rect 1572 1040 1603 1061
rect 1993 1040 2029 1061
rect 1415 1039 1452 1040
rect 106 1019 154 1028
rect 107 1018 154 1019
rect 420 1023 530 1037
rect 420 1020 463 1023
rect 420 1015 424 1020
rect 342 993 424 1015
rect 453 993 463 1020
rect 491 996 498 1023
rect 527 1015 530 1023
rect 1414 1030 1452 1039
rect 527 996 592 1015
rect 1414 1010 1423 1030
rect 1443 1010 1452 1030
rect 491 993 592 996
rect 342 991 592 993
rect 110 955 147 956
rect 106 952 147 955
rect 106 947 148 952
rect 106 929 119 947
rect 137 929 148 947
rect 106 915 148 929
rect 186 915 233 919
rect 106 909 233 915
rect 106 880 194 909
rect 223 880 233 909
rect 342 912 379 991
rect 420 978 530 991
rect 494 922 525 923
rect 342 892 351 912
rect 371 892 379 912
rect 342 882 379 892
rect 438 912 525 922
rect 438 892 447 912
rect 467 892 525 912
rect 438 883 525 892
rect 438 882 475 883
rect 106 876 233 880
rect 106 859 145 876
rect 186 875 233 876
rect 106 841 117 859
rect 135 841 145 859
rect 106 832 145 841
rect 107 831 144 832
rect 494 830 525 883
rect 555 912 592 991
rect 763 988 1156 1008
rect 1176 988 1179 1008
rect 1414 1002 1452 1010
rect 1518 1034 1603 1040
rect 1628 1039 1665 1040
rect 1518 1014 1526 1034
rect 1546 1014 1603 1034
rect 1518 1006 1603 1014
rect 1627 1030 1665 1039
rect 1627 1010 1636 1030
rect 1656 1010 1665 1030
rect 1518 1005 1554 1006
rect 1627 1002 1665 1010
rect 1731 1034 1816 1040
rect 1836 1039 1873 1040
rect 1731 1014 1739 1034
rect 1759 1033 1816 1034
rect 1759 1014 1788 1033
rect 1731 1013 1788 1014
rect 1809 1013 1816 1033
rect 1731 1006 1816 1013
rect 1835 1030 1873 1039
rect 1835 1010 1844 1030
rect 1864 1010 1873 1030
rect 1731 1005 1767 1006
rect 1835 1002 1873 1010
rect 1939 1034 2083 1040
rect 1939 1014 1947 1034
rect 1967 1032 2055 1034
rect 1967 1014 1996 1032
rect 1939 1011 1996 1014
rect 2023 1014 2055 1032
rect 2075 1014 2083 1034
rect 2023 1011 2083 1014
rect 1939 1006 2083 1011
rect 1939 1005 1975 1006
rect 2047 1005 2083 1006
rect 2149 1039 2186 1040
rect 2149 1038 2187 1039
rect 2149 1030 2213 1038
rect 2149 1010 2158 1030
rect 2178 1016 2213 1030
rect 2233 1016 2236 1036
rect 2178 1011 2236 1016
rect 2178 1010 2213 1011
rect 763 983 1179 988
rect 763 982 1104 983
rect 707 922 738 923
rect 555 892 564 912
rect 584 892 592 912
rect 555 882 592 892
rect 651 915 738 922
rect 651 912 712 915
rect 651 892 660 912
rect 680 895 712 912
rect 733 895 738 915
rect 680 892 738 895
rect 651 885 738 892
rect 763 912 800 982
rect 1066 981 1103 982
rect 1415 973 1452 1002
rect 1416 971 1452 973
rect 1628 971 1665 1002
rect 1416 949 1665 971
rect 1836 970 1873 1002
rect 2149 998 2213 1010
rect 2253 972 2280 1150
rect 2112 970 2280 972
rect 1833 963 2280 970
rect 1497 943 1608 949
rect 1497 935 1538 943
rect 915 922 951 923
rect 763 892 772 912
rect 792 892 800 912
rect 651 883 707 885
rect 651 882 688 883
rect 763 882 800 892
rect 859 912 1007 922
rect 1107 919 1203 921
rect 859 892 868 912
rect 888 892 978 912
rect 998 892 1007 912
rect 859 883 1007 892
rect 1065 912 1203 919
rect 1065 892 1074 912
rect 1094 892 1203 912
rect 1497 915 1505 935
rect 1524 915 1538 935
rect 1497 913 1538 915
rect 1566 935 1608 943
rect 1566 915 1582 935
rect 1601 915 1608 935
rect 1833 936 1858 963
rect 1889 944 2280 963
rect 1889 936 1938 944
rect 2112 943 2280 944
rect 1833 934 1938 936
rect 1566 913 1608 915
rect 1497 898 1608 913
rect 1065 883 1203 892
rect 859 882 896 883
rect 915 831 951 883
rect 970 882 1007 883
rect 1066 882 1103 883
rect 386 829 427 830
rect 278 822 427 829
rect 278 802 396 822
rect 416 802 427 822
rect 278 794 427 802
rect 494 826 853 830
rect 494 821 816 826
rect 494 797 607 821
rect 631 802 816 821
rect 840 802 853 826
rect 631 797 853 802
rect 494 794 853 797
rect 915 794 950 831
rect 1018 828 1118 831
rect 1018 824 1085 828
rect 1018 798 1030 824
rect 1056 802 1085 824
rect 1111 802 1118 828
rect 1056 798 1118 802
rect 1018 794 1118 798
rect 494 773 525 794
rect 915 773 951 794
rect 337 772 374 773
rect 111 769 145 770
rect 110 760 147 769
rect 110 742 119 760
rect 137 742 147 760
rect 110 732 147 742
rect 336 763 374 772
rect 336 743 345 763
rect 365 743 374 763
rect 336 735 374 743
rect 440 767 525 773
rect 550 772 587 773
rect 440 747 448 767
rect 468 747 525 767
rect 440 739 525 747
rect 549 763 587 772
rect 549 743 558 763
rect 578 743 587 763
rect 440 738 476 739
rect 549 735 587 743
rect 653 767 738 773
rect 758 772 795 773
rect 653 747 661 767
rect 681 766 738 767
rect 681 747 710 766
rect 653 746 710 747
rect 731 746 738 766
rect 653 739 738 746
rect 757 763 795 772
rect 757 743 766 763
rect 786 743 795 763
rect 653 738 689 739
rect 757 735 795 743
rect 861 767 1005 773
rect 861 747 869 767
rect 889 766 977 767
rect 889 747 920 766
rect 861 746 920 747
rect 945 747 977 766
rect 997 747 1005 767
rect 945 746 1005 747
rect 861 739 1005 746
rect 861 738 897 739
rect 969 738 1005 739
rect 1071 772 1108 773
rect 1071 771 1109 772
rect 1071 763 1135 771
rect 1071 743 1080 763
rect 1100 749 1135 763
rect 1155 749 1158 769
rect 1100 744 1158 749
rect 1100 743 1135 744
rect 111 704 145 732
rect 337 706 374 735
rect 338 704 374 706
rect 550 704 587 735
rect 111 703 283 704
rect 111 671 297 703
rect 338 682 587 704
rect 758 703 795 735
rect 1071 731 1135 743
rect 1175 705 1202 883
rect 1358 779 1468 793
rect 1358 776 1401 779
rect 1358 771 1362 776
rect 1034 703 1202 705
rect 758 697 1202 703
rect 111 639 145 671
rect 107 630 145 639
rect 107 612 117 630
rect 135 612 145 630
rect 107 606 145 612
rect 263 608 297 671
rect 419 676 530 682
rect 419 668 460 676
rect 419 648 427 668
rect 446 648 460 668
rect 419 646 460 648
rect 488 668 530 676
rect 488 648 504 668
rect 523 648 530 668
rect 488 646 530 648
rect 419 631 530 646
rect 757 677 1202 697
rect 757 608 795 677
rect 1034 676 1202 677
rect 1280 749 1362 771
rect 1391 749 1401 776
rect 1429 752 1436 779
rect 1465 771 1468 779
rect 1465 752 1530 771
rect 1429 749 1530 752
rect 1280 747 1530 749
rect 1280 668 1317 747
rect 1358 734 1468 747
rect 1432 678 1463 679
rect 1280 648 1289 668
rect 1309 648 1317 668
rect 1280 638 1317 648
rect 1376 668 1463 678
rect 1376 648 1385 668
rect 1405 648 1463 668
rect 1376 639 1463 648
rect 1376 638 1413 639
rect 107 602 144 606
rect 263 597 795 608
rect 262 581 795 597
rect 1432 586 1463 639
rect 1493 668 1530 747
rect 1701 757 2094 764
rect 1701 740 1709 757
rect 1741 744 2094 757
rect 2114 744 2117 764
rect 1741 740 2117 744
rect 1701 739 2117 740
rect 1701 738 2042 739
rect 1645 678 1676 679
rect 1493 648 1502 668
rect 1522 648 1530 668
rect 1493 638 1530 648
rect 1589 671 1676 678
rect 1589 668 1650 671
rect 1589 648 1598 668
rect 1618 651 1650 668
rect 1671 651 1676 671
rect 1618 648 1676 651
rect 1589 641 1676 648
rect 1701 668 1738 738
rect 2004 737 2041 738
rect 1853 678 1889 679
rect 1701 648 1710 668
rect 1730 648 1738 668
rect 1589 639 1645 641
rect 1589 638 1626 639
rect 1701 638 1738 648
rect 1797 668 1945 678
rect 2045 675 2141 677
rect 1797 648 1806 668
rect 1826 663 1916 668
rect 1826 648 1861 663
rect 1797 639 1861 648
rect 1797 638 1834 639
rect 1853 622 1861 639
rect 1882 648 1916 663
rect 1936 648 1945 668
rect 1882 639 1945 648
rect 2003 668 2141 675
rect 2003 648 2012 668
rect 2032 648 2141 668
rect 2003 639 2141 648
rect 1882 622 1889 639
rect 1908 638 1945 639
rect 2004 638 2041 639
rect 1853 587 1889 622
rect 1324 585 1365 586
rect 262 580 776 581
rect 1216 578 1365 585
rect 1216 558 1334 578
rect 1354 558 1365 578
rect 1216 550 1365 558
rect 1432 582 1791 586
rect 1432 577 1754 582
rect 1432 553 1545 577
rect 1569 558 1754 577
rect 1778 558 1791 582
rect 1569 553 1791 558
rect 1432 550 1791 553
rect 1853 550 1888 587
rect 1956 584 2056 587
rect 1956 580 2023 584
rect 1956 554 1968 580
rect 1994 558 2023 580
rect 2049 558 2056 584
rect 1994 554 2056 558
rect 1956 550 2056 554
rect 110 539 147 540
rect 108 531 148 539
rect 108 513 119 531
rect 137 513 148 531
rect 1432 529 1463 550
rect 1853 529 1889 550
rect 1275 528 1312 529
rect 108 465 148 513
rect 1274 519 1312 528
rect 1274 499 1283 519
rect 1303 499 1312 519
rect 1274 491 1312 499
rect 1378 523 1463 529
rect 1488 528 1525 529
rect 1378 503 1386 523
rect 1406 503 1463 523
rect 1378 495 1463 503
rect 1487 519 1525 528
rect 1487 499 1496 519
rect 1516 499 1525 519
rect 1378 494 1414 495
rect 1487 491 1525 499
rect 1591 523 1676 529
rect 1696 528 1733 529
rect 1591 503 1599 523
rect 1619 522 1676 523
rect 1619 503 1648 522
rect 1591 502 1648 503
rect 1669 502 1676 522
rect 1591 495 1676 502
rect 1695 519 1733 528
rect 1695 499 1704 519
rect 1724 499 1733 519
rect 1591 494 1627 495
rect 1695 491 1733 499
rect 1799 523 1943 529
rect 1799 503 1807 523
rect 1827 503 1915 523
rect 1935 503 1943 523
rect 1799 495 1943 503
rect 1799 494 1835 495
rect 1907 494 1943 495
rect 2009 528 2046 529
rect 2009 527 2047 528
rect 2009 519 2073 527
rect 2009 499 2018 519
rect 2038 505 2073 519
rect 2093 505 2096 525
rect 2038 500 2096 505
rect 2038 499 2073 500
rect 419 469 529 483
rect 419 466 462 469
rect 108 458 233 465
rect 419 461 423 466
rect 108 439 200 458
rect 225 439 233 458
rect 108 429 233 439
rect 341 439 423 461
rect 452 439 462 466
rect 490 442 497 469
rect 526 461 529 469
rect 1275 462 1312 491
rect 526 442 591 461
rect 1276 460 1312 462
rect 1488 460 1525 491
rect 1696 464 1733 491
rect 2009 487 2073 499
rect 490 439 591 442
rect 341 437 591 439
rect 108 409 148 429
rect 107 400 148 409
rect 107 382 117 400
rect 135 382 148 400
rect 107 373 148 382
rect 107 372 144 373
rect 341 358 378 437
rect 419 424 529 437
rect 493 368 524 369
rect 341 338 350 358
rect 370 338 378 358
rect 341 328 378 338
rect 437 358 524 368
rect 437 338 446 358
rect 466 338 524 358
rect 437 329 524 338
rect 437 328 474 329
rect 110 306 147 310
rect 107 301 147 306
rect 107 283 119 301
rect 137 283 147 301
rect 107 103 147 283
rect 493 276 524 329
rect 554 358 591 437
rect 762 434 1155 454
rect 1175 434 1178 454
rect 1276 438 1525 460
rect 1694 459 1735 464
rect 2113 461 2140 639
rect 1972 459 2140 461
rect 1694 453 2140 459
rect 762 429 1178 434
rect 1357 432 1468 438
rect 762 428 1103 429
rect 706 368 737 369
rect 554 338 563 358
rect 583 338 591 358
rect 554 328 591 338
rect 650 361 737 368
rect 650 358 711 361
rect 650 338 659 358
rect 679 341 711 358
rect 732 341 737 361
rect 679 338 737 341
rect 650 331 737 338
rect 762 358 799 428
rect 1065 427 1102 428
rect 1357 424 1398 432
rect 1357 404 1365 424
rect 1384 404 1398 424
rect 1357 402 1398 404
rect 1426 424 1468 432
rect 1426 404 1442 424
rect 1461 404 1468 424
rect 1694 431 1700 453
rect 1726 433 2140 453
rect 1726 431 1735 433
rect 1972 432 2140 433
rect 1694 422 1735 431
rect 1426 402 1468 404
rect 1357 387 1468 402
rect 914 368 950 369
rect 762 338 771 358
rect 791 338 799 358
rect 650 329 706 331
rect 650 328 687 329
rect 762 328 799 338
rect 858 358 1006 368
rect 1106 365 1202 367
rect 858 338 867 358
rect 887 338 977 358
rect 997 338 1006 358
rect 858 329 1006 338
rect 1064 358 1202 365
rect 1064 338 1073 358
rect 1093 338 1202 358
rect 1064 329 1202 338
rect 858 328 895 329
rect 914 277 950 329
rect 969 328 1006 329
rect 1065 328 1102 329
rect 385 275 426 276
rect 277 268 426 275
rect 277 248 395 268
rect 415 248 426 268
rect 277 240 426 248
rect 493 272 852 276
rect 493 267 815 272
rect 493 243 606 267
rect 630 248 815 267
rect 839 248 852 272
rect 630 243 852 248
rect 493 240 852 243
rect 914 240 949 277
rect 1017 274 1117 277
rect 1017 270 1084 274
rect 1017 244 1029 270
rect 1055 248 1084 270
rect 1110 248 1117 274
rect 1055 244 1117 248
rect 1017 240 1117 244
rect 493 219 524 240
rect 914 219 950 240
rect 336 218 373 219
rect 335 209 373 218
rect 335 189 344 209
rect 364 189 373 209
rect 335 181 373 189
rect 439 213 524 219
rect 549 218 586 219
rect 439 193 447 213
rect 467 193 524 213
rect 439 185 524 193
rect 548 209 586 218
rect 548 189 557 209
rect 577 189 586 209
rect 439 184 475 185
rect 548 181 586 189
rect 652 213 737 219
rect 757 218 794 219
rect 652 193 660 213
rect 680 212 737 213
rect 680 193 709 212
rect 652 192 709 193
rect 730 192 737 212
rect 652 185 737 192
rect 756 209 794 218
rect 756 189 765 209
rect 785 189 794 209
rect 652 184 688 185
rect 756 181 794 189
rect 860 213 1004 219
rect 860 193 868 213
rect 888 210 976 213
rect 888 193 919 210
rect 860 190 919 193
rect 942 193 976 210
rect 996 193 1004 213
rect 942 190 1004 193
rect 860 185 1004 190
rect 860 184 896 185
rect 968 184 1004 185
rect 1070 218 1107 219
rect 1070 217 1108 218
rect 1070 209 1134 217
rect 1070 189 1079 209
rect 1099 195 1134 209
rect 1154 195 1157 215
rect 1099 190 1157 195
rect 1099 189 1134 190
rect 336 152 373 181
rect 337 150 373 152
rect 549 150 586 181
rect 337 128 586 150
rect 757 149 794 181
rect 1070 177 1134 189
rect 1174 151 1201 329
rect 1468 200 1578 214
rect 1468 197 1511 200
rect 1468 192 1472 197
rect 1033 149 1201 151
rect 757 146 1201 149
rect 418 122 529 128
rect 418 114 459 122
rect 107 59 146 103
rect 418 94 426 114
rect 445 94 459 114
rect 418 92 459 94
rect 487 114 529 122
rect 487 94 503 114
rect 522 94 529 114
rect 487 92 529 94
rect 418 78 529 92
rect 755 123 1201 146
rect 107 35 147 59
rect 447 35 494 37
rect 755 35 793 123
rect 1033 122 1201 123
rect 1390 170 1472 192
rect 1501 170 1511 197
rect 1539 173 1546 200
rect 1575 192 1578 200
rect 1575 173 1640 192
rect 1539 170 1640 173
rect 1390 168 1640 170
rect 1390 89 1427 168
rect 1468 155 1578 168
rect 1542 99 1573 100
rect 1390 69 1399 89
rect 1419 69 1427 89
rect 1390 59 1427 69
rect 1486 89 1573 99
rect 1486 69 1495 89
rect 1515 69 1573 89
rect 1486 60 1573 69
rect 1486 59 1523 60
rect 107 2 793 35
rect 1542 7 1573 60
rect 1603 89 1640 168
rect 1811 165 2204 185
rect 2224 165 2227 185
rect 1811 160 2227 165
rect 1811 159 2152 160
rect 1755 99 1786 100
rect 1603 69 1612 89
rect 1632 69 1640 89
rect 1603 59 1640 69
rect 1699 92 1786 99
rect 1699 89 1760 92
rect 1699 69 1708 89
rect 1728 72 1760 89
rect 1781 72 1786 92
rect 1728 69 1786 72
rect 1699 62 1786 69
rect 1811 89 1848 159
rect 2114 158 2151 159
rect 1963 99 1999 100
rect 1811 69 1820 89
rect 1840 69 1848 89
rect 1699 60 1755 62
rect 1699 59 1736 60
rect 1811 59 1848 69
rect 1907 89 2055 99
rect 2155 96 2251 98
rect 1907 69 1916 89
rect 1936 69 2026 89
rect 2046 69 2055 89
rect 1907 60 2055 69
rect 2113 89 2251 96
rect 2113 69 2122 89
rect 2142 69 2251 89
rect 2113 60 2251 69
rect 1907 59 1944 60
rect 1963 8 1999 60
rect 2018 59 2055 60
rect 2114 59 2151 60
rect 1434 6 1475 7
rect 106 -55 145 2
rect 755 0 793 2
rect 1326 -1 1475 6
rect 1326 -21 1444 -1
rect 1464 -21 1475 -1
rect 1326 -29 1475 -21
rect 1542 3 1901 7
rect 1542 -2 1864 3
rect 1542 -26 1655 -2
rect 1679 -21 1864 -2
rect 1888 -21 1901 3
rect 1679 -26 1901 -21
rect 1542 -29 1901 -26
rect 1963 -29 1998 8
rect 2066 5 2166 8
rect 2066 1 2133 5
rect 2066 -25 2078 1
rect 2104 -21 2133 1
rect 2159 -21 2166 5
rect 2104 -25 2166 -21
rect 2066 -29 2166 -25
rect 1542 -50 1573 -29
rect 1963 -50 1999 -29
rect 1385 -51 1422 -50
rect 106 -57 154 -55
rect 106 -75 117 -57
rect 135 -75 154 -57
rect 1384 -60 1422 -51
rect 106 -84 154 -75
rect 107 -85 154 -84
rect 420 -80 530 -66
rect 420 -83 463 -80
rect 420 -88 424 -83
rect 342 -110 424 -88
rect 453 -110 463 -83
rect 491 -107 498 -80
rect 527 -88 530 -80
rect 1384 -80 1393 -60
rect 1413 -80 1422 -60
rect 1384 -88 1422 -80
rect 1488 -56 1573 -50
rect 1598 -51 1635 -50
rect 1488 -76 1496 -56
rect 1516 -76 1573 -56
rect 1488 -84 1573 -76
rect 1597 -60 1635 -51
rect 1597 -80 1606 -60
rect 1626 -80 1635 -60
rect 1488 -85 1524 -84
rect 1597 -88 1635 -80
rect 1701 -56 1786 -50
rect 1806 -51 1843 -50
rect 1701 -76 1709 -56
rect 1729 -57 1786 -56
rect 1729 -76 1758 -57
rect 1701 -77 1758 -76
rect 1779 -77 1786 -57
rect 1701 -84 1786 -77
rect 1805 -60 1843 -51
rect 1805 -80 1814 -60
rect 1834 -80 1843 -60
rect 1701 -85 1737 -84
rect 1805 -88 1843 -80
rect 1909 -56 2053 -50
rect 1909 -76 1917 -56
rect 1937 -76 2025 -56
rect 2045 -76 2053 -56
rect 1909 -84 2053 -76
rect 1909 -85 1945 -84
rect 2017 -85 2053 -84
rect 2119 -51 2156 -50
rect 2119 -52 2157 -51
rect 2119 -60 2183 -52
rect 2119 -80 2128 -60
rect 2148 -74 2183 -60
rect 2203 -74 2206 -54
rect 2148 -79 2206 -74
rect 2148 -80 2183 -79
rect 527 -107 592 -88
rect 491 -110 592 -107
rect 342 -112 592 -110
rect 110 -148 147 -147
rect 106 -151 147 -148
rect 106 -156 148 -151
rect 106 -174 119 -156
rect 137 -174 148 -156
rect 106 -188 148 -174
rect 186 -188 233 -184
rect 106 -194 233 -188
rect 106 -223 194 -194
rect 223 -223 233 -194
rect 342 -191 379 -112
rect 420 -125 530 -112
rect 494 -181 525 -180
rect 342 -211 351 -191
rect 371 -211 379 -191
rect 342 -221 379 -211
rect 438 -191 525 -181
rect 438 -211 447 -191
rect 467 -211 525 -191
rect 438 -220 525 -211
rect 438 -221 475 -220
rect 106 -227 233 -223
rect 106 -244 145 -227
rect 186 -228 233 -227
rect 106 -262 117 -244
rect 135 -262 145 -244
rect 106 -271 145 -262
rect 107 -272 144 -271
rect 494 -273 525 -220
rect 555 -191 592 -112
rect 763 -115 1156 -95
rect 1176 -115 1179 -95
rect 763 -120 1179 -115
rect 1385 -117 1422 -88
rect 1386 -119 1422 -117
rect 1598 -119 1635 -88
rect 763 -121 1104 -120
rect 707 -181 738 -180
rect 555 -211 564 -191
rect 584 -211 592 -191
rect 555 -221 592 -211
rect 651 -188 738 -181
rect 651 -191 712 -188
rect 651 -211 660 -191
rect 680 -208 712 -191
rect 733 -208 738 -188
rect 680 -211 738 -208
rect 651 -218 738 -211
rect 763 -191 800 -121
rect 1066 -122 1103 -121
rect 1386 -141 1635 -119
rect 1806 -120 1843 -88
rect 2119 -92 2183 -80
rect 2223 -110 2250 60
rect 2171 -118 2250 -110
rect 2082 -120 2250 -118
rect 1806 -127 2250 -120
rect 1467 -147 1578 -141
rect 1806 -146 2176 -127
rect 2082 -147 2176 -146
rect 1467 -155 1508 -147
rect 1467 -175 1475 -155
rect 1494 -175 1508 -155
rect 1467 -177 1508 -175
rect 1536 -155 1578 -147
rect 1536 -175 1552 -155
rect 1571 -175 1578 -155
rect 2171 -156 2176 -147
rect 2224 -147 2250 -127
rect 2224 -156 2241 -147
rect 2171 -165 2241 -156
rect 1536 -177 1578 -175
rect 915 -181 951 -180
rect 763 -211 772 -191
rect 792 -211 800 -191
rect 651 -220 707 -218
rect 651 -221 688 -220
rect 763 -221 800 -211
rect 859 -191 1007 -181
rect 1107 -184 1203 -182
rect 859 -211 868 -191
rect 888 -211 978 -191
rect 998 -211 1007 -191
rect 859 -220 1007 -211
rect 1065 -191 1203 -184
rect 1065 -211 1074 -191
rect 1094 -211 1203 -191
rect 1467 -192 1578 -177
rect 1065 -220 1203 -211
rect 859 -221 896 -220
rect 915 -272 951 -220
rect 970 -221 1007 -220
rect 1066 -221 1103 -220
rect 386 -274 427 -273
rect 278 -281 427 -274
rect 278 -301 396 -281
rect 416 -301 427 -281
rect 278 -309 427 -301
rect 494 -277 853 -273
rect 494 -282 816 -277
rect 494 -306 607 -282
rect 631 -301 816 -282
rect 840 -301 853 -277
rect 631 -306 853 -301
rect 494 -309 853 -306
rect 915 -309 950 -272
rect 1018 -275 1118 -272
rect 1018 -279 1085 -275
rect 1018 -305 1030 -279
rect 1056 -301 1085 -279
rect 1111 -301 1118 -275
rect 1056 -305 1118 -301
rect 1018 -309 1118 -305
rect 494 -330 525 -309
rect 915 -330 951 -309
rect 337 -331 374 -330
rect 111 -334 145 -333
rect 110 -343 147 -334
rect 110 -361 119 -343
rect 137 -361 147 -343
rect 110 -371 147 -361
rect 336 -340 374 -331
rect 336 -360 345 -340
rect 365 -360 374 -340
rect 336 -368 374 -360
rect 440 -336 525 -330
rect 550 -331 587 -330
rect 440 -356 448 -336
rect 468 -356 525 -336
rect 440 -364 525 -356
rect 549 -340 587 -331
rect 549 -360 558 -340
rect 578 -360 587 -340
rect 440 -365 476 -364
rect 549 -368 587 -360
rect 653 -336 738 -330
rect 758 -331 795 -330
rect 653 -356 661 -336
rect 681 -337 738 -336
rect 681 -356 710 -337
rect 653 -357 710 -356
rect 731 -357 738 -337
rect 653 -364 738 -357
rect 757 -340 795 -331
rect 757 -360 766 -340
rect 786 -360 795 -340
rect 653 -365 689 -364
rect 757 -368 795 -360
rect 861 -336 1005 -330
rect 861 -356 869 -336
rect 889 -337 977 -336
rect 889 -356 920 -337
rect 861 -357 920 -356
rect 945 -356 977 -337
rect 997 -356 1005 -336
rect 945 -357 1005 -356
rect 861 -364 1005 -357
rect 861 -365 897 -364
rect 969 -365 1005 -364
rect 1071 -331 1108 -330
rect 1071 -332 1109 -331
rect 1071 -340 1135 -332
rect 1071 -360 1080 -340
rect 1100 -354 1135 -340
rect 1155 -354 1158 -334
rect 1100 -359 1158 -354
rect 1100 -360 1135 -359
rect 111 -399 145 -371
rect 337 -397 374 -368
rect 338 -399 374 -397
rect 550 -399 587 -368
rect 111 -400 283 -399
rect 111 -432 297 -400
rect 338 -421 587 -399
rect 758 -400 795 -368
rect 1071 -372 1135 -360
rect 1175 -398 1202 -220
rect 1358 -324 1468 -310
rect 1358 -327 1401 -324
rect 1358 -332 1362 -327
rect 1034 -400 1202 -398
rect 758 -406 1202 -400
rect 111 -464 145 -432
rect 107 -473 145 -464
rect 107 -491 117 -473
rect 135 -491 145 -473
rect 107 -497 145 -491
rect 263 -495 297 -432
rect 419 -427 530 -421
rect 419 -435 460 -427
rect 419 -455 427 -435
rect 446 -455 460 -435
rect 419 -457 460 -455
rect 488 -435 530 -427
rect 488 -455 504 -435
rect 523 -455 530 -435
rect 488 -457 530 -455
rect 419 -472 530 -457
rect 757 -426 1202 -406
rect 757 -495 795 -426
rect 1034 -427 1202 -426
rect 1280 -354 1362 -332
rect 1391 -354 1401 -327
rect 1429 -351 1436 -324
rect 1465 -332 1468 -324
rect 1465 -351 1530 -332
rect 1429 -354 1530 -351
rect 1280 -356 1530 -354
rect 1280 -435 1317 -356
rect 1358 -369 1468 -356
rect 1432 -425 1463 -424
rect 1280 -455 1289 -435
rect 1309 -455 1317 -435
rect 1280 -465 1317 -455
rect 1376 -435 1463 -425
rect 1376 -455 1385 -435
rect 1405 -455 1463 -435
rect 1376 -464 1463 -455
rect 1376 -465 1413 -464
rect 107 -501 144 -497
rect 263 -506 795 -495
rect 262 -522 795 -506
rect 1432 -517 1463 -464
rect 1493 -435 1530 -356
rect 1701 -359 2094 -339
rect 2114 -359 2117 -339
rect 1701 -364 2117 -359
rect 1701 -365 2042 -364
rect 1645 -425 1676 -424
rect 1493 -455 1502 -435
rect 1522 -455 1530 -435
rect 1493 -465 1530 -455
rect 1589 -432 1676 -425
rect 1589 -435 1650 -432
rect 1589 -455 1598 -435
rect 1618 -452 1650 -435
rect 1671 -452 1676 -432
rect 1618 -455 1676 -452
rect 1589 -462 1676 -455
rect 1701 -435 1738 -365
rect 2004 -366 2041 -365
rect 1853 -425 1889 -424
rect 1701 -455 1710 -435
rect 1730 -455 1738 -435
rect 1589 -464 1645 -462
rect 1589 -465 1626 -464
rect 1701 -465 1738 -455
rect 1797 -435 1945 -425
rect 2045 -428 2141 -426
rect 1797 -455 1806 -435
rect 1826 -455 1916 -435
rect 1936 -455 1945 -435
rect 1797 -464 1945 -455
rect 2003 -435 2141 -428
rect 2003 -455 2012 -435
rect 2032 -455 2141 -435
rect 2003 -464 2141 -455
rect 1797 -465 1834 -464
rect 1853 -516 1889 -464
rect 1908 -465 1945 -464
rect 2004 -465 2041 -464
rect 1324 -518 1365 -517
rect 262 -523 776 -522
rect 1216 -525 1365 -518
rect 1216 -545 1334 -525
rect 1354 -545 1365 -525
rect 1216 -553 1365 -545
rect 1432 -521 1791 -517
rect 1432 -526 1754 -521
rect 1432 -550 1545 -526
rect 1569 -545 1754 -526
rect 1778 -545 1791 -521
rect 1569 -550 1791 -545
rect 1432 -553 1791 -550
rect 1853 -553 1888 -516
rect 1956 -519 2056 -516
rect 1956 -523 2023 -519
rect 1956 -549 1968 -523
rect 1994 -545 2023 -523
rect 2049 -545 2056 -519
rect 1994 -549 2056 -545
rect 1956 -553 2056 -549
rect 110 -564 147 -563
rect 108 -572 148 -564
rect 108 -590 119 -572
rect 137 -590 148 -572
rect 1432 -574 1463 -553
rect 1853 -574 1889 -553
rect 1275 -575 1312 -574
rect 108 -638 148 -590
rect 1274 -584 1312 -575
rect 1274 -604 1283 -584
rect 1303 -604 1312 -584
rect 1274 -612 1312 -604
rect 1378 -580 1463 -574
rect 1488 -575 1525 -574
rect 1378 -600 1386 -580
rect 1406 -600 1463 -580
rect 1378 -608 1463 -600
rect 1487 -584 1525 -575
rect 1487 -604 1496 -584
rect 1516 -604 1525 -584
rect 1378 -609 1414 -608
rect 1487 -612 1525 -604
rect 1591 -580 1676 -574
rect 1696 -575 1733 -574
rect 1591 -600 1599 -580
rect 1619 -581 1676 -580
rect 1619 -600 1648 -581
rect 1591 -601 1648 -600
rect 1669 -601 1676 -581
rect 1591 -608 1676 -601
rect 1695 -584 1733 -575
rect 1695 -604 1704 -584
rect 1724 -604 1733 -584
rect 1591 -609 1627 -608
rect 1695 -612 1733 -604
rect 1799 -580 1943 -574
rect 1799 -600 1807 -580
rect 1827 -597 1863 -580
rect 1883 -597 1915 -580
rect 1827 -600 1915 -597
rect 1935 -600 1943 -580
rect 1799 -608 1943 -600
rect 1799 -609 1835 -608
rect 1907 -609 1943 -608
rect 2009 -575 2046 -574
rect 2009 -576 2047 -575
rect 2009 -584 2073 -576
rect 2009 -604 2018 -584
rect 2038 -598 2073 -584
rect 2093 -598 2096 -578
rect 2038 -603 2096 -598
rect 2038 -604 2073 -603
rect 419 -634 529 -620
rect 419 -637 462 -634
rect 108 -645 233 -638
rect 419 -642 423 -637
rect 108 -664 200 -645
rect 225 -664 233 -645
rect 108 -674 233 -664
rect 341 -664 423 -642
rect 452 -664 462 -637
rect 490 -661 497 -634
rect 526 -642 529 -634
rect 1275 -641 1312 -612
rect 526 -661 591 -642
rect 1276 -643 1312 -641
rect 1488 -643 1525 -612
rect 1696 -639 1733 -612
rect 2009 -616 2073 -604
rect 490 -664 591 -661
rect 341 -666 591 -664
rect 108 -694 148 -674
rect 107 -703 148 -694
rect 107 -721 117 -703
rect 135 -721 148 -703
rect 107 -730 148 -721
rect 107 -731 144 -730
rect 341 -745 378 -666
rect 419 -679 529 -666
rect 493 -735 524 -734
rect 341 -765 350 -745
rect 370 -765 378 -745
rect 341 -775 378 -765
rect 437 -745 524 -735
rect 437 -765 446 -745
rect 466 -765 524 -745
rect 437 -774 524 -765
rect 437 -775 474 -774
rect 110 -797 147 -793
rect 107 -802 147 -797
rect 107 -820 119 -802
rect 137 -820 147 -802
rect 107 -1000 147 -820
rect 493 -827 524 -774
rect 554 -745 591 -666
rect 762 -669 1155 -649
rect 1175 -669 1178 -649
rect 1276 -665 1525 -643
rect 1694 -644 1735 -639
rect 2113 -642 2140 -464
rect 1972 -644 2140 -642
rect 1694 -650 2140 -644
rect 762 -674 1178 -669
rect 1357 -671 1468 -665
rect 762 -675 1103 -674
rect 706 -735 737 -734
rect 554 -765 563 -745
rect 583 -765 591 -745
rect 554 -775 591 -765
rect 650 -742 737 -735
rect 650 -745 711 -742
rect 650 -765 659 -745
rect 679 -762 711 -745
rect 732 -762 737 -742
rect 679 -765 737 -762
rect 650 -772 737 -765
rect 762 -745 799 -675
rect 1065 -676 1102 -675
rect 1357 -679 1398 -671
rect 1357 -699 1365 -679
rect 1384 -699 1398 -679
rect 1357 -701 1398 -699
rect 1426 -679 1468 -671
rect 1426 -699 1442 -679
rect 1461 -699 1468 -679
rect 1694 -672 1700 -650
rect 1726 -670 2140 -650
rect 1726 -672 1735 -670
rect 1972 -671 2140 -670
rect 1694 -681 1735 -672
rect 1426 -701 1468 -699
rect 1357 -716 1468 -701
rect 914 -735 950 -734
rect 762 -765 771 -745
rect 791 -765 799 -745
rect 650 -774 706 -772
rect 650 -775 687 -774
rect 762 -775 799 -765
rect 858 -745 1006 -735
rect 1106 -738 1202 -736
rect 858 -765 867 -745
rect 887 -765 977 -745
rect 997 -765 1006 -745
rect 858 -774 1006 -765
rect 1064 -745 1202 -738
rect 1064 -765 1073 -745
rect 1093 -765 1202 -745
rect 1064 -774 1202 -765
rect 858 -775 895 -774
rect 914 -826 950 -774
rect 969 -775 1006 -774
rect 1065 -775 1102 -774
rect 385 -828 426 -827
rect 277 -835 426 -828
rect 277 -855 395 -835
rect 415 -855 426 -835
rect 277 -863 426 -855
rect 493 -831 852 -827
rect 493 -836 815 -831
rect 493 -860 606 -836
rect 630 -855 815 -836
rect 839 -855 852 -831
rect 630 -860 852 -855
rect 493 -863 852 -860
rect 914 -863 949 -826
rect 1017 -829 1117 -826
rect 1017 -833 1084 -829
rect 1017 -859 1029 -833
rect 1055 -855 1084 -833
rect 1110 -855 1117 -829
rect 1055 -859 1117 -855
rect 1017 -863 1117 -859
rect 493 -884 524 -863
rect 914 -884 950 -863
rect 336 -885 373 -884
rect 335 -894 373 -885
rect 335 -914 344 -894
rect 364 -914 373 -894
rect 335 -922 373 -914
rect 439 -890 524 -884
rect 549 -885 586 -884
rect 439 -910 447 -890
rect 467 -910 524 -890
rect 439 -918 524 -910
rect 548 -894 586 -885
rect 548 -914 557 -894
rect 577 -914 586 -894
rect 439 -919 475 -918
rect 548 -922 586 -914
rect 652 -890 737 -884
rect 757 -885 794 -884
rect 652 -910 660 -890
rect 680 -891 737 -890
rect 680 -910 709 -891
rect 652 -911 709 -910
rect 730 -911 737 -891
rect 652 -918 737 -911
rect 756 -894 794 -885
rect 756 -914 765 -894
rect 785 -914 794 -894
rect 652 -919 688 -918
rect 756 -922 794 -914
rect 860 -890 1004 -884
rect 860 -910 868 -890
rect 888 -893 976 -890
rect 888 -910 919 -893
rect 860 -913 919 -910
rect 942 -910 976 -893
rect 996 -910 1004 -890
rect 942 -913 1004 -910
rect 860 -918 1004 -913
rect 860 -919 896 -918
rect 968 -919 1004 -918
rect 1070 -885 1107 -884
rect 1070 -886 1108 -885
rect 1070 -894 1134 -886
rect 1070 -914 1079 -894
rect 1099 -908 1134 -894
rect 1154 -908 1157 -888
rect 1099 -913 1157 -908
rect 1099 -914 1134 -913
rect 336 -951 373 -922
rect 337 -953 373 -951
rect 549 -953 586 -922
rect 337 -975 586 -953
rect 757 -954 794 -922
rect 1070 -926 1134 -914
rect 1174 -952 1201 -774
rect 1499 -916 1609 -902
rect 1499 -919 1542 -916
rect 1499 -924 1503 -919
rect 1033 -954 1201 -952
rect 757 -957 1201 -954
rect 418 -981 529 -975
rect 418 -989 459 -981
rect 107 -1044 146 -1000
rect 418 -1009 426 -989
rect 445 -1009 459 -989
rect 418 -1011 459 -1009
rect 487 -989 529 -981
rect 487 -1009 503 -989
rect 522 -1009 529 -989
rect 487 -1011 529 -1009
rect 418 -1026 529 -1011
rect 755 -980 1201 -957
rect 107 -1068 147 -1044
rect 447 -1068 494 -1066
rect 755 -1068 793 -980
rect 1033 -981 1201 -980
rect 1421 -946 1503 -924
rect 1532 -946 1542 -919
rect 1570 -943 1577 -916
rect 1606 -924 1609 -916
rect 1606 -943 1671 -924
rect 1570 -946 1671 -943
rect 1421 -948 1671 -946
rect 1421 -1027 1458 -948
rect 1499 -961 1609 -948
rect 1573 -1017 1604 -1016
rect 1421 -1047 1430 -1027
rect 1450 -1047 1458 -1027
rect 1421 -1057 1458 -1047
rect 1517 -1027 1604 -1017
rect 1517 -1047 1526 -1027
rect 1546 -1047 1604 -1027
rect 1517 -1056 1604 -1047
rect 1517 -1057 1554 -1056
rect 107 -1101 793 -1068
rect 107 -1158 146 -1101
rect 755 -1103 793 -1101
rect 1573 -1109 1604 -1056
rect 1634 -1027 1671 -948
rect 1842 -935 2235 -931
rect 1842 -952 1861 -935
rect 1881 -951 2235 -935
rect 2255 -951 2258 -931
rect 1881 -952 2258 -951
rect 1842 -956 2258 -952
rect 1842 -957 2183 -956
rect 1786 -1017 1817 -1016
rect 1634 -1047 1643 -1027
rect 1663 -1047 1671 -1027
rect 1634 -1057 1671 -1047
rect 1730 -1024 1817 -1017
rect 1730 -1027 1791 -1024
rect 1730 -1047 1739 -1027
rect 1759 -1044 1791 -1027
rect 1812 -1044 1817 -1024
rect 1759 -1047 1817 -1044
rect 1730 -1054 1817 -1047
rect 1842 -1027 1879 -957
rect 2145 -958 2182 -957
rect 1994 -1017 2030 -1016
rect 1842 -1047 1851 -1027
rect 1871 -1047 1879 -1027
rect 1730 -1056 1786 -1054
rect 1730 -1057 1767 -1056
rect 1842 -1057 1879 -1047
rect 1938 -1027 2086 -1017
rect 2254 -1018 2283 -1017
rect 2186 -1020 2283 -1018
rect 1938 -1047 1947 -1027
rect 1967 -1031 2057 -1027
rect 1967 -1047 2000 -1031
rect 1938 -1056 2000 -1047
rect 1938 -1057 1975 -1056
rect 1994 -1069 2000 -1056
rect 2023 -1047 2057 -1031
rect 2077 -1047 2086 -1027
rect 2023 -1056 2086 -1047
rect 2144 -1027 2283 -1020
rect 2144 -1047 2153 -1027
rect 2173 -1047 2283 -1027
rect 2144 -1056 2283 -1047
rect 2023 -1069 2030 -1056
rect 2049 -1057 2086 -1056
rect 2145 -1057 2182 -1056
rect 1994 -1108 2030 -1069
rect 1465 -1110 1506 -1109
rect 1357 -1117 1506 -1110
rect 1357 -1137 1475 -1117
rect 1495 -1137 1506 -1117
rect 1357 -1145 1506 -1137
rect 1573 -1113 1932 -1109
rect 1573 -1118 1895 -1113
rect 1573 -1142 1686 -1118
rect 1710 -1137 1895 -1118
rect 1919 -1137 1932 -1113
rect 1710 -1142 1932 -1137
rect 1573 -1145 1932 -1142
rect 1994 -1145 2029 -1108
rect 2097 -1111 2197 -1108
rect 2097 -1115 2164 -1111
rect 2097 -1141 2109 -1115
rect 2135 -1137 2164 -1115
rect 2190 -1137 2197 -1111
rect 2135 -1141 2197 -1137
rect 2097 -1145 2197 -1141
rect 107 -1160 155 -1158
rect 107 -1178 118 -1160
rect 136 -1178 155 -1160
rect 1573 -1166 1604 -1145
rect 1994 -1166 2030 -1145
rect 1416 -1167 1453 -1166
rect 107 -1187 155 -1178
rect 108 -1188 155 -1187
rect 421 -1183 531 -1169
rect 421 -1186 464 -1183
rect 421 -1191 425 -1186
rect 343 -1213 425 -1191
rect 454 -1213 464 -1186
rect 492 -1210 499 -1183
rect 528 -1191 531 -1183
rect 1415 -1176 1453 -1167
rect 528 -1210 593 -1191
rect 1415 -1196 1424 -1176
rect 1444 -1196 1453 -1176
rect 492 -1213 593 -1210
rect 343 -1215 593 -1213
rect 111 -1251 148 -1250
rect 107 -1254 148 -1251
rect 107 -1259 149 -1254
rect 107 -1277 120 -1259
rect 138 -1277 149 -1259
rect 107 -1291 149 -1277
rect 187 -1291 234 -1287
rect 107 -1297 234 -1291
rect 107 -1326 195 -1297
rect 224 -1326 234 -1297
rect 343 -1294 380 -1215
rect 421 -1228 531 -1215
rect 495 -1284 526 -1283
rect 343 -1314 352 -1294
rect 372 -1314 380 -1294
rect 343 -1324 380 -1314
rect 439 -1294 526 -1284
rect 439 -1314 448 -1294
rect 468 -1314 526 -1294
rect 439 -1323 526 -1314
rect 439 -1324 476 -1323
rect 107 -1330 234 -1326
rect 107 -1347 146 -1330
rect 187 -1331 234 -1330
rect 107 -1365 118 -1347
rect 136 -1365 146 -1347
rect 107 -1374 146 -1365
rect 108 -1375 145 -1374
rect 495 -1376 526 -1323
rect 556 -1294 593 -1215
rect 764 -1218 1157 -1198
rect 1177 -1218 1180 -1198
rect 1415 -1204 1453 -1196
rect 1519 -1172 1604 -1166
rect 1629 -1167 1666 -1166
rect 1519 -1192 1527 -1172
rect 1547 -1192 1604 -1172
rect 1519 -1200 1604 -1192
rect 1628 -1176 1666 -1167
rect 1628 -1196 1637 -1176
rect 1657 -1196 1666 -1176
rect 1519 -1201 1555 -1200
rect 1628 -1204 1666 -1196
rect 1732 -1172 1817 -1166
rect 1837 -1167 1874 -1166
rect 1732 -1192 1740 -1172
rect 1760 -1173 1817 -1172
rect 1760 -1192 1789 -1173
rect 1732 -1193 1789 -1192
rect 1810 -1193 1817 -1173
rect 1732 -1200 1817 -1193
rect 1836 -1176 1874 -1167
rect 1836 -1196 1845 -1176
rect 1865 -1196 1874 -1176
rect 1732 -1201 1768 -1200
rect 1836 -1204 1874 -1196
rect 1940 -1172 2084 -1166
rect 1940 -1192 1948 -1172
rect 1968 -1192 2056 -1172
rect 2076 -1192 2084 -1172
rect 1940 -1200 2084 -1192
rect 1940 -1201 1976 -1200
rect 2048 -1201 2084 -1200
rect 2150 -1167 2187 -1166
rect 2150 -1168 2188 -1167
rect 2150 -1176 2214 -1168
rect 2150 -1196 2159 -1176
rect 2179 -1190 2214 -1176
rect 2234 -1190 2237 -1170
rect 2179 -1195 2237 -1190
rect 2179 -1196 2214 -1195
rect 764 -1223 1180 -1218
rect 764 -1224 1105 -1223
rect 708 -1284 739 -1283
rect 556 -1314 565 -1294
rect 585 -1314 593 -1294
rect 556 -1324 593 -1314
rect 652 -1291 739 -1284
rect 652 -1294 713 -1291
rect 652 -1314 661 -1294
rect 681 -1311 713 -1294
rect 734 -1311 739 -1291
rect 681 -1314 739 -1311
rect 652 -1321 739 -1314
rect 764 -1294 801 -1224
rect 1067 -1225 1104 -1224
rect 1416 -1233 1453 -1204
rect 1417 -1235 1453 -1233
rect 1629 -1235 1666 -1204
rect 1417 -1257 1666 -1235
rect 1837 -1236 1874 -1204
rect 2150 -1208 2214 -1196
rect 2254 -1234 2283 -1056
rect 2113 -1236 2283 -1234
rect 1834 -1243 2283 -1236
rect 1498 -1263 1609 -1257
rect 1498 -1271 1539 -1263
rect 916 -1284 952 -1283
rect 764 -1314 773 -1294
rect 793 -1314 801 -1294
rect 652 -1323 708 -1321
rect 652 -1324 689 -1323
rect 764 -1324 801 -1314
rect 860 -1294 1008 -1284
rect 1108 -1287 1204 -1285
rect 860 -1314 869 -1294
rect 889 -1314 979 -1294
rect 999 -1314 1008 -1294
rect 860 -1323 1008 -1314
rect 1066 -1294 1204 -1287
rect 1066 -1314 1075 -1294
rect 1095 -1314 1204 -1294
rect 1498 -1291 1506 -1271
rect 1525 -1291 1539 -1271
rect 1498 -1293 1539 -1291
rect 1567 -1271 1609 -1263
rect 1567 -1291 1583 -1271
rect 1602 -1291 1609 -1271
rect 1834 -1270 1859 -1243
rect 1890 -1262 2283 -1243
rect 1890 -1270 1939 -1262
rect 2113 -1263 2283 -1262
rect 1834 -1272 1939 -1270
rect 1567 -1293 1609 -1291
rect 1498 -1308 1609 -1293
rect 1066 -1323 1204 -1314
rect 860 -1324 897 -1323
rect 916 -1375 952 -1323
rect 971 -1324 1008 -1323
rect 1067 -1324 1104 -1323
rect 387 -1377 428 -1376
rect 279 -1384 428 -1377
rect 279 -1404 397 -1384
rect 417 -1404 428 -1384
rect 279 -1412 428 -1404
rect 495 -1380 854 -1376
rect 495 -1385 817 -1380
rect 495 -1409 608 -1385
rect 632 -1404 817 -1385
rect 841 -1404 854 -1380
rect 632 -1409 854 -1404
rect 495 -1412 854 -1409
rect 916 -1412 951 -1375
rect 1019 -1378 1119 -1375
rect 1019 -1382 1086 -1378
rect 1019 -1408 1031 -1382
rect 1057 -1404 1086 -1382
rect 1112 -1404 1119 -1378
rect 1057 -1408 1119 -1404
rect 1019 -1412 1119 -1408
rect 495 -1433 526 -1412
rect 916 -1433 952 -1412
rect 338 -1434 375 -1433
rect 112 -1437 146 -1436
rect 111 -1446 148 -1437
rect 111 -1464 120 -1446
rect 138 -1464 148 -1446
rect 111 -1474 148 -1464
rect 337 -1443 375 -1434
rect 337 -1463 346 -1443
rect 366 -1463 375 -1443
rect 337 -1471 375 -1463
rect 441 -1439 526 -1433
rect 551 -1434 588 -1433
rect 441 -1459 449 -1439
rect 469 -1459 526 -1439
rect 441 -1467 526 -1459
rect 550 -1443 588 -1434
rect 550 -1463 559 -1443
rect 579 -1463 588 -1443
rect 441 -1468 477 -1467
rect 550 -1471 588 -1463
rect 654 -1439 739 -1433
rect 759 -1434 796 -1433
rect 654 -1459 662 -1439
rect 682 -1440 739 -1439
rect 682 -1459 711 -1440
rect 654 -1460 711 -1459
rect 732 -1460 739 -1440
rect 654 -1467 739 -1460
rect 758 -1443 796 -1434
rect 758 -1463 767 -1443
rect 787 -1463 796 -1443
rect 654 -1468 690 -1467
rect 758 -1471 796 -1463
rect 862 -1439 1006 -1433
rect 862 -1459 870 -1439
rect 890 -1440 978 -1439
rect 890 -1459 921 -1440
rect 862 -1460 921 -1459
rect 946 -1459 978 -1440
rect 998 -1459 1006 -1439
rect 946 -1460 1006 -1459
rect 862 -1467 1006 -1460
rect 862 -1468 898 -1467
rect 970 -1468 1006 -1467
rect 1072 -1434 1109 -1433
rect 1072 -1435 1110 -1434
rect 1072 -1443 1136 -1435
rect 1072 -1463 1081 -1443
rect 1101 -1457 1136 -1443
rect 1156 -1457 1159 -1437
rect 1101 -1462 1159 -1457
rect 1101 -1463 1136 -1462
rect 112 -1502 146 -1474
rect 338 -1500 375 -1471
rect 339 -1502 375 -1500
rect 551 -1502 588 -1471
rect 112 -1503 284 -1502
rect 112 -1535 298 -1503
rect 339 -1524 588 -1502
rect 759 -1503 796 -1471
rect 1072 -1475 1136 -1463
rect 1176 -1501 1203 -1323
rect 1359 -1427 1469 -1413
rect 1359 -1430 1402 -1427
rect 1359 -1435 1363 -1430
rect 1035 -1503 1203 -1501
rect 759 -1509 1203 -1503
rect 112 -1567 146 -1535
rect 108 -1576 146 -1567
rect 108 -1594 118 -1576
rect 136 -1594 146 -1576
rect 108 -1600 146 -1594
rect 264 -1598 298 -1535
rect 420 -1530 531 -1524
rect 420 -1538 461 -1530
rect 420 -1558 428 -1538
rect 447 -1558 461 -1538
rect 420 -1560 461 -1558
rect 489 -1538 531 -1530
rect 489 -1558 505 -1538
rect 524 -1558 531 -1538
rect 489 -1560 531 -1558
rect 420 -1575 531 -1560
rect 758 -1529 1203 -1509
rect 758 -1598 796 -1529
rect 1035 -1530 1203 -1529
rect 1281 -1457 1363 -1435
rect 1392 -1457 1402 -1430
rect 1430 -1454 1437 -1427
rect 1466 -1435 1469 -1427
rect 1466 -1454 1531 -1435
rect 1430 -1457 1531 -1454
rect 1281 -1459 1531 -1457
rect 1281 -1538 1318 -1459
rect 1359 -1472 1469 -1459
rect 1433 -1528 1464 -1527
rect 1281 -1558 1290 -1538
rect 1310 -1558 1318 -1538
rect 1281 -1568 1318 -1558
rect 1377 -1538 1464 -1528
rect 1377 -1558 1386 -1538
rect 1406 -1558 1464 -1538
rect 1377 -1567 1464 -1558
rect 1377 -1568 1414 -1567
rect 108 -1604 145 -1600
rect 264 -1609 796 -1598
rect 263 -1625 796 -1609
rect 1433 -1620 1464 -1567
rect 1494 -1538 1531 -1459
rect 1702 -1449 2095 -1442
rect 1702 -1466 1710 -1449
rect 1742 -1462 2095 -1449
rect 2115 -1462 2118 -1442
rect 1742 -1466 2118 -1462
rect 1702 -1467 2118 -1466
rect 1702 -1468 2043 -1467
rect 1646 -1528 1677 -1527
rect 1494 -1558 1503 -1538
rect 1523 -1558 1531 -1538
rect 1494 -1568 1531 -1558
rect 1590 -1535 1677 -1528
rect 1590 -1538 1651 -1535
rect 1590 -1558 1599 -1538
rect 1619 -1555 1651 -1538
rect 1672 -1555 1677 -1535
rect 1619 -1558 1677 -1555
rect 1590 -1565 1677 -1558
rect 1702 -1538 1739 -1468
rect 2005 -1469 2042 -1468
rect 1854 -1528 1890 -1527
rect 1702 -1558 1711 -1538
rect 1731 -1558 1739 -1538
rect 1590 -1567 1646 -1565
rect 1590 -1568 1627 -1567
rect 1702 -1568 1739 -1558
rect 1798 -1538 1946 -1528
rect 2046 -1531 2142 -1529
rect 1798 -1558 1807 -1538
rect 1827 -1543 1917 -1538
rect 1827 -1558 1862 -1543
rect 1798 -1567 1862 -1558
rect 1798 -1568 1835 -1567
rect 1854 -1584 1862 -1567
rect 1883 -1558 1917 -1543
rect 1937 -1558 1946 -1538
rect 1883 -1567 1946 -1558
rect 2004 -1538 2142 -1531
rect 2004 -1558 2013 -1538
rect 2033 -1558 2142 -1538
rect 2004 -1567 2142 -1558
rect 1883 -1584 1890 -1567
rect 1909 -1568 1946 -1567
rect 2005 -1568 2042 -1567
rect 1854 -1619 1890 -1584
rect 1325 -1621 1366 -1620
rect 263 -1626 777 -1625
rect 1217 -1628 1366 -1621
rect 1217 -1648 1335 -1628
rect 1355 -1648 1366 -1628
rect 1217 -1656 1366 -1648
rect 1433 -1624 1792 -1620
rect 1433 -1629 1755 -1624
rect 1433 -1653 1546 -1629
rect 1570 -1648 1755 -1629
rect 1779 -1648 1792 -1624
rect 1570 -1653 1792 -1648
rect 1433 -1656 1792 -1653
rect 1854 -1656 1889 -1619
rect 1957 -1622 2057 -1619
rect 1957 -1626 2024 -1622
rect 1957 -1652 1969 -1626
rect 1995 -1648 2024 -1626
rect 2050 -1648 2057 -1622
rect 1995 -1652 2057 -1648
rect 1957 -1656 2057 -1652
rect 111 -1667 148 -1666
rect 109 -1675 149 -1667
rect 109 -1693 120 -1675
rect 138 -1693 149 -1675
rect 1433 -1677 1464 -1656
rect 1854 -1677 1890 -1656
rect 1276 -1678 1313 -1677
rect 109 -1741 149 -1693
rect 1275 -1687 1313 -1678
rect 1275 -1707 1284 -1687
rect 1304 -1707 1313 -1687
rect 1275 -1715 1313 -1707
rect 1379 -1683 1464 -1677
rect 1489 -1678 1526 -1677
rect 1379 -1703 1387 -1683
rect 1407 -1703 1464 -1683
rect 1379 -1711 1464 -1703
rect 1488 -1687 1526 -1678
rect 1488 -1707 1497 -1687
rect 1517 -1707 1526 -1687
rect 1379 -1712 1415 -1711
rect 1488 -1715 1526 -1707
rect 1592 -1683 1677 -1677
rect 1697 -1678 1734 -1677
rect 1592 -1703 1600 -1683
rect 1620 -1684 1677 -1683
rect 1620 -1703 1649 -1684
rect 1592 -1704 1649 -1703
rect 1670 -1704 1677 -1684
rect 1592 -1711 1677 -1704
rect 1696 -1687 1734 -1678
rect 1696 -1707 1705 -1687
rect 1725 -1707 1734 -1687
rect 1592 -1712 1628 -1711
rect 1696 -1715 1734 -1707
rect 1800 -1683 1944 -1677
rect 1800 -1703 1808 -1683
rect 1828 -1703 1916 -1683
rect 1936 -1703 1944 -1683
rect 1800 -1711 1944 -1703
rect 1800 -1712 1836 -1711
rect 1908 -1712 1944 -1711
rect 2010 -1678 2047 -1677
rect 2010 -1679 2048 -1678
rect 2010 -1687 2074 -1679
rect 2010 -1707 2019 -1687
rect 2039 -1701 2074 -1687
rect 2094 -1701 2097 -1681
rect 2039 -1706 2097 -1701
rect 2039 -1707 2074 -1706
rect 420 -1737 530 -1723
rect 420 -1740 463 -1737
rect 109 -1748 234 -1741
rect 420 -1745 424 -1740
rect 109 -1767 201 -1748
rect 226 -1767 234 -1748
rect 109 -1777 234 -1767
rect 342 -1767 424 -1745
rect 453 -1767 463 -1740
rect 491 -1764 498 -1737
rect 527 -1745 530 -1737
rect 1276 -1744 1313 -1715
rect 527 -1764 592 -1745
rect 1277 -1746 1313 -1744
rect 1489 -1746 1526 -1715
rect 1697 -1742 1734 -1715
rect 2010 -1719 2074 -1707
rect 491 -1767 592 -1764
rect 342 -1769 592 -1767
rect 109 -1797 149 -1777
rect 108 -1806 149 -1797
rect 108 -1824 118 -1806
rect 136 -1824 149 -1806
rect 108 -1833 149 -1824
rect 108 -1834 145 -1833
rect 342 -1848 379 -1769
rect 420 -1782 530 -1769
rect 494 -1838 525 -1837
rect 342 -1868 351 -1848
rect 371 -1868 379 -1848
rect 342 -1878 379 -1868
rect 438 -1848 525 -1838
rect 438 -1868 447 -1848
rect 467 -1868 525 -1848
rect 438 -1877 525 -1868
rect 438 -1878 475 -1877
rect 111 -1900 148 -1896
rect 108 -1905 148 -1900
rect 108 -1923 120 -1905
rect 138 -1923 148 -1905
rect 108 -2103 148 -1923
rect 494 -1930 525 -1877
rect 555 -1848 592 -1769
rect 763 -1772 1156 -1752
rect 1176 -1772 1179 -1752
rect 1277 -1768 1526 -1746
rect 1695 -1747 1736 -1742
rect 2114 -1745 2141 -1567
rect 1973 -1747 2141 -1745
rect 1695 -1753 2141 -1747
rect 763 -1777 1179 -1772
rect 1358 -1774 1469 -1768
rect 763 -1778 1104 -1777
rect 707 -1838 738 -1837
rect 555 -1868 564 -1848
rect 584 -1868 592 -1848
rect 555 -1878 592 -1868
rect 651 -1845 738 -1838
rect 651 -1848 712 -1845
rect 651 -1868 660 -1848
rect 680 -1865 712 -1848
rect 733 -1865 738 -1845
rect 680 -1868 738 -1865
rect 651 -1875 738 -1868
rect 763 -1848 800 -1778
rect 1066 -1779 1103 -1778
rect 1358 -1782 1399 -1774
rect 1358 -1802 1366 -1782
rect 1385 -1802 1399 -1782
rect 1358 -1804 1399 -1802
rect 1427 -1782 1469 -1774
rect 1427 -1802 1443 -1782
rect 1462 -1802 1469 -1782
rect 1695 -1775 1701 -1753
rect 1727 -1773 2141 -1753
rect 1727 -1775 1736 -1773
rect 1973 -1774 2141 -1773
rect 1695 -1784 1736 -1775
rect 1427 -1804 1469 -1802
rect 1358 -1819 1469 -1804
rect 915 -1838 951 -1837
rect 763 -1868 772 -1848
rect 792 -1868 800 -1848
rect 651 -1877 707 -1875
rect 651 -1878 688 -1877
rect 763 -1878 800 -1868
rect 859 -1848 1007 -1838
rect 1107 -1841 1203 -1839
rect 859 -1868 868 -1848
rect 888 -1868 978 -1848
rect 998 -1868 1007 -1848
rect 859 -1877 1007 -1868
rect 1065 -1848 1203 -1841
rect 1065 -1868 1074 -1848
rect 1094 -1868 1203 -1848
rect 1065 -1877 1203 -1868
rect 859 -1878 896 -1877
rect 915 -1929 951 -1877
rect 970 -1878 1007 -1877
rect 1066 -1878 1103 -1877
rect 386 -1931 427 -1930
rect 278 -1938 427 -1931
rect 278 -1958 396 -1938
rect 416 -1958 427 -1938
rect 278 -1966 427 -1958
rect 494 -1934 853 -1930
rect 494 -1939 816 -1934
rect 494 -1963 607 -1939
rect 631 -1958 816 -1939
rect 840 -1958 853 -1934
rect 631 -1963 853 -1958
rect 494 -1966 853 -1963
rect 915 -1966 950 -1929
rect 1018 -1932 1118 -1929
rect 1018 -1936 1085 -1932
rect 1018 -1962 1030 -1936
rect 1056 -1958 1085 -1936
rect 1111 -1958 1118 -1932
rect 1056 -1962 1118 -1958
rect 1018 -1966 1118 -1962
rect 494 -1987 525 -1966
rect 915 -1987 951 -1966
rect 337 -1988 374 -1987
rect 336 -1997 374 -1988
rect 336 -2017 345 -1997
rect 365 -2017 374 -1997
rect 336 -2025 374 -2017
rect 440 -1993 525 -1987
rect 550 -1988 587 -1987
rect 440 -2013 448 -1993
rect 468 -2013 525 -1993
rect 440 -2021 525 -2013
rect 549 -1997 587 -1988
rect 549 -2017 558 -1997
rect 578 -2017 587 -1997
rect 440 -2022 476 -2021
rect 549 -2025 587 -2017
rect 653 -1993 738 -1987
rect 758 -1988 795 -1987
rect 653 -2013 661 -1993
rect 681 -1994 738 -1993
rect 681 -2013 710 -1994
rect 653 -2014 710 -2013
rect 731 -2014 738 -1994
rect 653 -2021 738 -2014
rect 757 -1997 795 -1988
rect 757 -2017 766 -1997
rect 786 -2017 795 -1997
rect 653 -2022 689 -2021
rect 757 -2025 795 -2017
rect 861 -1993 1005 -1987
rect 861 -2013 869 -1993
rect 889 -1996 977 -1993
rect 889 -2013 920 -1996
rect 861 -2016 920 -2013
rect 943 -2013 977 -1996
rect 997 -2013 1005 -1993
rect 943 -2016 1005 -2013
rect 861 -2021 1005 -2016
rect 861 -2022 897 -2021
rect 969 -2022 1005 -2021
rect 1071 -1988 1108 -1987
rect 1071 -1989 1109 -1988
rect 1071 -1997 1135 -1989
rect 1071 -2017 1080 -1997
rect 1100 -2011 1135 -1997
rect 1155 -2011 1158 -1991
rect 1100 -2016 1158 -2011
rect 1100 -2017 1135 -2016
rect 337 -2054 374 -2025
rect 338 -2056 374 -2054
rect 550 -2056 587 -2025
rect 338 -2078 587 -2056
rect 758 -2057 795 -2025
rect 1071 -2029 1135 -2017
rect 1175 -2055 1202 -1877
rect 1034 -2057 1202 -2055
rect 758 -2060 1202 -2057
rect 419 -2084 530 -2078
rect 419 -2092 460 -2084
rect 108 -2147 147 -2103
rect 419 -2112 427 -2092
rect 446 -2112 460 -2092
rect 419 -2114 460 -2112
rect 488 -2092 530 -2084
rect 488 -2112 504 -2092
rect 523 -2112 530 -2092
rect 488 -2113 530 -2112
rect 756 -2083 1202 -2060
rect 488 -2114 531 -2113
rect 108 -2171 148 -2147
rect 419 -2153 531 -2114
rect 448 -2171 495 -2153
rect 756 -2171 794 -2083
rect 1034 -2084 1202 -2083
rect 108 -2204 794 -2171
rect 756 -2206 794 -2204
<< viali >>
rect 423 2096 452 2123
rect 497 2099 526 2126
rect 193 1983 222 2012
rect 1155 2091 1175 2111
rect 711 1998 732 2018
rect 1084 1905 1110 1931
rect 709 1849 730 1869
rect 919 1849 944 1869
rect 1134 1852 1154 1872
rect 426 1751 445 1771
rect 503 1751 522 1771
rect 1361 1852 1390 1879
rect 1435 1855 1464 1882
rect 2093 1847 2113 1867
rect 1649 1754 1670 1774
rect 2022 1661 2048 1687
rect 1647 1605 1668 1625
rect 1862 1609 1882 1626
rect 2072 1608 2092 1628
rect 199 1542 224 1561
rect 422 1542 451 1569
rect 496 1545 525 1572
rect 1154 1537 1174 1557
rect 710 1444 731 1464
rect 1364 1507 1383 1527
rect 1441 1507 1460 1527
rect 1699 1534 1725 1556
rect 1083 1351 1109 1377
rect 708 1295 729 1315
rect 918 1293 941 1313
rect 1133 1298 1153 1318
rect 425 1197 444 1217
rect 502 1197 521 1217
rect 1502 1260 1531 1287
rect 1576 1263 1605 1290
rect 1860 1254 1880 1271
rect 2234 1255 2254 1275
rect 1790 1162 1811 1182
rect 2163 1069 2189 1095
rect 424 993 453 1020
rect 498 996 527 1023
rect 194 880 223 909
rect 1156 988 1176 1008
rect 1788 1013 1809 1033
rect 1996 1011 2023 1032
rect 2213 1016 2233 1036
rect 712 895 733 915
rect 1505 915 1524 935
rect 1582 915 1601 935
rect 1858 936 1889 963
rect 1085 802 1111 828
rect 710 746 731 766
rect 920 746 945 766
rect 1135 749 1155 769
rect 427 648 446 668
rect 504 648 523 668
rect 1362 749 1391 776
rect 1436 752 1465 779
rect 1709 740 1741 757
rect 2094 744 2114 764
rect 1650 651 1671 671
rect 1861 622 1882 663
rect 2023 558 2049 584
rect 1648 502 1669 522
rect 2073 505 2093 525
rect 200 439 225 458
rect 423 439 452 466
rect 497 442 526 469
rect 1155 434 1175 454
rect 711 341 732 361
rect 1365 404 1384 424
rect 1442 404 1461 424
rect 1700 431 1726 453
rect 1084 248 1110 274
rect 709 192 730 212
rect 919 190 942 210
rect 1134 195 1154 215
rect 426 94 445 114
rect 503 94 522 114
rect 1472 170 1501 197
rect 1546 173 1575 200
rect 2204 165 2224 185
rect 1760 72 1781 92
rect 2133 -21 2159 5
rect 424 -110 453 -83
rect 498 -107 527 -80
rect 1758 -77 1779 -57
rect 2183 -74 2203 -54
rect 194 -223 223 -194
rect 1156 -115 1176 -95
rect 712 -208 733 -188
rect 1475 -175 1494 -155
rect 1552 -175 1571 -155
rect 2176 -156 2224 -127
rect 1085 -301 1111 -275
rect 710 -357 731 -337
rect 920 -357 945 -337
rect 1135 -354 1155 -334
rect 427 -455 446 -435
rect 504 -455 523 -435
rect 1362 -354 1391 -327
rect 1436 -351 1465 -324
rect 2094 -359 2114 -339
rect 1650 -452 1671 -432
rect 2023 -545 2049 -519
rect 1648 -601 1669 -581
rect 1863 -597 1883 -580
rect 2073 -598 2093 -578
rect 200 -664 225 -645
rect 423 -664 452 -637
rect 497 -661 526 -634
rect 1155 -669 1175 -649
rect 711 -762 732 -742
rect 1365 -699 1384 -679
rect 1442 -699 1461 -679
rect 1700 -672 1726 -650
rect 1084 -855 1110 -829
rect 709 -911 730 -891
rect 919 -913 942 -893
rect 1134 -908 1154 -888
rect 426 -1009 445 -989
rect 503 -1009 522 -989
rect 1503 -946 1532 -919
rect 1577 -943 1606 -916
rect 1861 -952 1881 -935
rect 2235 -951 2255 -931
rect 1791 -1044 1812 -1024
rect 2000 -1069 2023 -1031
rect 2164 -1137 2190 -1111
rect 425 -1213 454 -1186
rect 499 -1210 528 -1183
rect 195 -1326 224 -1297
rect 1157 -1218 1177 -1198
rect 1789 -1193 1810 -1173
rect 2214 -1190 2234 -1170
rect 713 -1311 734 -1291
rect 1506 -1291 1525 -1271
rect 1583 -1291 1602 -1271
rect 1859 -1270 1890 -1243
rect 1086 -1404 1112 -1378
rect 711 -1460 732 -1440
rect 921 -1460 946 -1440
rect 1136 -1457 1156 -1437
rect 428 -1558 447 -1538
rect 505 -1558 524 -1538
rect 1363 -1457 1392 -1430
rect 1437 -1454 1466 -1427
rect 1710 -1466 1742 -1449
rect 2095 -1462 2115 -1442
rect 1651 -1555 1672 -1535
rect 1862 -1584 1883 -1543
rect 2024 -1648 2050 -1622
rect 1649 -1704 1670 -1684
rect 2074 -1701 2094 -1681
rect 201 -1767 226 -1748
rect 424 -1767 453 -1740
rect 498 -1764 527 -1737
rect 1156 -1772 1176 -1752
rect 712 -1865 733 -1845
rect 1366 -1802 1385 -1782
rect 1443 -1802 1462 -1782
rect 1701 -1775 1727 -1753
rect 1085 -1958 1111 -1932
rect 710 -2014 731 -1994
rect 920 -2016 943 -1996
rect 1135 -2011 1155 -1991
rect 427 -2112 446 -2092
rect 504 -2112 523 -2092
<< metal1 >>
rect 1150 2194 1185 2196
rect 186 2191 1185 2194
rect 185 2167 1185 2191
rect 185 2012 233 2167
rect 419 2126 529 2140
rect 419 2123 497 2126
rect 419 2096 423 2123
rect 452 2099 497 2123
rect 526 2099 529 2126
rect 1150 2116 1185 2167
rect 452 2096 529 2099
rect 419 2081 529 2096
rect 1148 2111 1185 2116
rect 1148 2091 1155 2111
rect 1175 2091 1185 2111
rect 1148 2084 1185 2091
rect 1148 2083 1183 2084
rect 185 1983 193 2012
rect 222 1983 233 2012
rect 185 1978 233 1983
rect 704 2018 736 2025
rect 704 1998 711 2018
rect 732 1998 736 2018
rect 704 1933 736 1998
rect 1074 1933 1114 1934
rect 704 1931 1116 1933
rect 704 1905 1084 1931
rect 1110 1905 1116 1931
rect 704 1897 1116 1905
rect 704 1869 736 1897
rect 1149 1877 1183 2083
rect 2087 1950 2121 1951
rect 1218 1915 2122 1950
rect 704 1849 709 1869
rect 730 1849 736 1869
rect 704 1842 736 1849
rect 911 1869 950 1875
rect 911 1849 919 1869
rect 944 1849 950 1869
rect 911 1842 950 1849
rect 1127 1872 1183 1877
rect 1127 1852 1134 1872
rect 1154 1852 1183 1872
rect 1127 1845 1183 1852
rect 1127 1844 1162 1845
rect 919 1796 950 1842
rect 418 1771 529 1793
rect 418 1751 426 1771
rect 445 1751 503 1771
rect 522 1751 529 1771
rect 918 1779 950 1796
rect 1219 1779 1256 1915
rect 1357 1882 1467 1896
rect 1357 1879 1435 1882
rect 1357 1852 1361 1879
rect 1390 1855 1435 1879
rect 1464 1855 1467 1882
rect 2087 1872 2121 1915
rect 1390 1852 1467 1855
rect 1357 1837 1467 1852
rect 2086 1867 2121 1872
rect 2086 1847 2093 1867
rect 2113 1847 2121 1867
rect 2086 1839 2121 1847
rect 918 1766 1256 1779
rect 418 1734 529 1751
rect 919 1747 1256 1766
rect 1198 1746 1256 1747
rect 1642 1774 1674 1781
rect 1642 1754 1649 1774
rect 1670 1754 1674 1774
rect 1642 1689 1674 1754
rect 2012 1689 2052 1690
rect 1642 1687 2054 1689
rect 1642 1661 2022 1687
rect 2048 1661 2054 1687
rect 1642 1653 2054 1661
rect 188 1614 1184 1640
rect 1642 1625 1674 1653
rect 190 1561 232 1614
rect 190 1542 199 1561
rect 224 1542 232 1561
rect 190 1532 232 1542
rect 418 1572 528 1586
rect 418 1569 496 1572
rect 418 1542 422 1569
rect 451 1545 496 1569
rect 525 1545 528 1572
rect 1148 1562 1182 1614
rect 1642 1605 1647 1625
rect 1668 1605 1674 1625
rect 1642 1598 1674 1605
rect 1852 1626 1890 1636
rect 2087 1633 2121 1839
rect 1852 1609 1862 1626
rect 1882 1609 1890 1626
rect 1693 1566 1734 1567
rect 451 1542 528 1545
rect 418 1527 528 1542
rect 1147 1557 1182 1562
rect 1147 1537 1154 1557
rect 1174 1537 1182 1557
rect 1692 1556 1734 1566
rect 1147 1529 1182 1537
rect 703 1464 735 1471
rect 703 1444 710 1464
rect 731 1444 735 1464
rect 703 1379 735 1444
rect 1073 1379 1113 1380
rect 703 1377 1115 1379
rect 703 1351 1083 1377
rect 1109 1351 1115 1377
rect 703 1343 1115 1351
rect 703 1315 735 1343
rect 1148 1323 1182 1529
rect 1356 1527 1467 1549
rect 1356 1507 1364 1527
rect 1383 1507 1441 1527
rect 1460 1507 1467 1527
rect 1356 1490 1467 1507
rect 1692 1534 1699 1556
rect 1725 1534 1734 1556
rect 1692 1525 1734 1534
rect 909 1320 952 1322
rect 703 1295 708 1315
rect 729 1295 735 1315
rect 703 1288 735 1295
rect 908 1313 952 1320
rect 908 1293 918 1313
rect 941 1293 952 1313
rect 908 1289 952 1293
rect 1126 1318 1182 1323
rect 1126 1298 1133 1318
rect 1153 1298 1182 1318
rect 1126 1291 1182 1298
rect 1238 1459 1271 1460
rect 1692 1459 1729 1525
rect 1238 1430 1729 1459
rect 1126 1290 1161 1291
rect 417 1217 528 1239
rect 417 1197 425 1217
rect 444 1197 502 1217
rect 521 1197 528 1217
rect 417 1180 528 1197
rect 908 1208 950 1289
rect 1238 1210 1271 1430
rect 1692 1428 1729 1430
rect 1498 1290 1608 1304
rect 1498 1287 1576 1290
rect 1498 1260 1502 1287
rect 1531 1263 1576 1287
rect 1605 1263 1608 1290
rect 1531 1260 1608 1263
rect 1498 1245 1608 1260
rect 1852 1271 1890 1609
rect 2065 1628 2121 1633
rect 2065 1608 2072 1628
rect 2092 1608 2121 1628
rect 2065 1601 2121 1608
rect 2065 1600 2100 1601
rect 2230 1280 2262 1281
rect 1852 1254 1860 1271
rect 1880 1254 1890 1271
rect 1852 1248 1890 1254
rect 2227 1275 2262 1280
rect 2227 1255 2234 1275
rect 2254 1255 2262 1275
rect 2227 1247 2262 1255
rect 1210 1208 1271 1210
rect 908 1179 1271 1208
rect 1783 1182 1815 1189
rect 908 1177 1210 1179
rect 1783 1162 1790 1182
rect 1811 1162 1815 1182
rect 1783 1097 1815 1162
rect 2153 1097 2193 1098
rect 1783 1095 2195 1097
rect 1151 1091 1186 1093
rect 187 1088 1186 1091
rect 186 1064 1186 1088
rect 186 909 234 1064
rect 420 1023 530 1037
rect 420 1020 498 1023
rect 420 993 424 1020
rect 453 996 498 1020
rect 527 996 530 1023
rect 1151 1013 1186 1064
rect 453 993 530 996
rect 420 978 530 993
rect 1149 1008 1186 1013
rect 1149 988 1156 1008
rect 1176 988 1186 1008
rect 1783 1069 2163 1095
rect 2189 1069 2195 1095
rect 1783 1061 2195 1069
rect 1783 1033 1815 1061
rect 1783 1013 1788 1033
rect 1809 1013 1815 1033
rect 1783 1006 1815 1013
rect 1989 1032 2031 1043
rect 2228 1041 2262 1247
rect 1989 1011 1996 1032
rect 2023 1011 2031 1032
rect 1149 981 1186 988
rect 1149 980 1184 981
rect 186 880 194 909
rect 223 880 234 909
rect 186 875 234 880
rect 705 915 737 922
rect 705 895 712 915
rect 733 895 737 915
rect 705 830 737 895
rect 1075 830 1115 831
rect 705 828 1117 830
rect 705 802 1085 828
rect 1111 802 1117 828
rect 705 794 1117 802
rect 705 766 737 794
rect 1150 774 1184 980
rect 1854 963 1893 970
rect 1497 935 1608 957
rect 1497 915 1505 935
rect 1524 915 1582 935
rect 1601 915 1608 935
rect 1497 898 1608 915
rect 1854 936 1858 963
rect 1889 936 1893 963
rect 1701 847 1754 851
rect 1219 812 1754 847
rect 705 746 710 766
rect 731 746 737 766
rect 705 739 737 746
rect 912 766 951 772
rect 912 746 920 766
rect 945 746 951 766
rect 912 739 951 746
rect 1128 769 1184 774
rect 1128 749 1135 769
rect 1155 749 1184 769
rect 1128 742 1184 749
rect 1128 741 1163 742
rect 920 693 951 739
rect 419 668 530 690
rect 419 648 427 668
rect 446 648 504 668
rect 523 648 530 668
rect 919 676 951 693
rect 1220 676 1257 812
rect 1358 779 1468 793
rect 1358 776 1436 779
rect 1358 749 1362 776
rect 1391 752 1436 776
rect 1465 752 1468 779
rect 1391 749 1468 752
rect 1358 734 1468 749
rect 1700 765 1754 812
rect 1700 757 1753 765
rect 1700 740 1709 757
rect 1741 740 1753 757
rect 1700 737 1753 740
rect 919 663 1257 676
rect 419 631 530 648
rect 920 644 1257 663
rect 1199 643 1257 644
rect 1643 671 1675 678
rect 1643 651 1650 671
rect 1671 651 1675 671
rect 1643 586 1675 651
rect 1854 663 1893 936
rect 1989 840 2031 1011
rect 2206 1036 2262 1041
rect 2206 1016 2213 1036
rect 2233 1016 2262 1036
rect 2206 1009 2262 1016
rect 2206 1008 2241 1009
rect 1989 806 2233 840
rect 2196 798 2233 806
rect 2089 765 2123 776
rect 2087 764 2123 765
rect 2087 744 2094 764
rect 2114 744 2123 764
rect 2087 736 2123 744
rect 1854 622 1861 663
rect 1882 622 1893 663
rect 1854 607 1893 622
rect 2013 586 2053 587
rect 1643 584 2055 586
rect 1643 558 2023 584
rect 2049 558 2055 584
rect 1643 550 2055 558
rect 189 511 1185 537
rect 1643 522 1675 550
rect 2088 530 2122 736
rect 191 458 233 511
rect 191 439 200 458
rect 225 439 233 458
rect 191 429 233 439
rect 419 469 529 483
rect 419 466 497 469
rect 419 439 423 466
rect 452 442 497 466
rect 526 442 529 469
rect 1149 459 1183 511
rect 1643 502 1648 522
rect 1669 502 1675 522
rect 1643 495 1675 502
rect 2066 525 2122 530
rect 2066 505 2073 525
rect 2093 505 2122 525
rect 2066 498 2122 505
rect 2066 497 2101 498
rect 1694 463 1735 464
rect 452 439 529 442
rect 419 424 529 439
rect 1148 454 1183 459
rect 1148 434 1155 454
rect 1175 434 1183 454
rect 1693 453 1735 463
rect 1148 426 1183 434
rect 704 361 736 368
rect 704 341 711 361
rect 732 341 736 361
rect 704 276 736 341
rect 1074 276 1114 277
rect 704 274 1116 276
rect 704 248 1084 274
rect 1110 248 1116 274
rect 704 240 1116 248
rect 704 212 736 240
rect 1149 220 1183 426
rect 1357 424 1468 446
rect 1357 404 1365 424
rect 1384 404 1442 424
rect 1461 404 1468 424
rect 1357 387 1468 404
rect 1693 431 1700 453
rect 1726 431 1735 453
rect 1693 422 1735 431
rect 910 217 953 219
rect 704 192 709 212
rect 730 192 736 212
rect 704 185 736 192
rect 909 210 953 217
rect 909 190 919 210
rect 942 190 953 210
rect 909 186 953 190
rect 1127 215 1183 220
rect 1127 195 1134 215
rect 1154 195 1183 215
rect 1127 188 1183 195
rect 1239 356 1272 357
rect 1693 356 1730 422
rect 1239 327 1730 356
rect 1127 187 1162 188
rect 418 114 529 136
rect 418 94 426 114
rect 445 94 503 114
rect 522 94 529 114
rect 418 78 529 94
rect 909 105 951 186
rect 1239 107 1272 327
rect 1693 325 1730 327
rect 1468 200 1578 214
rect 1468 197 1546 200
rect 1468 170 1472 197
rect 1501 173 1546 197
rect 1575 173 1578 200
rect 1501 170 1578 173
rect 1468 155 1578 170
rect 2196 185 2234 798
rect 2196 165 2204 185
rect 2224 165 2234 185
rect 2196 158 2234 165
rect 2197 157 2232 158
rect 1211 105 1272 107
rect 909 76 1272 105
rect 1753 92 1785 99
rect 909 74 1211 76
rect 1753 72 1760 92
rect 1781 72 1785 92
rect 1753 7 1785 72
rect 2123 7 2163 8
rect 1753 5 2165 7
rect 1151 -12 1186 -10
rect 187 -15 1186 -12
rect 186 -39 1186 -15
rect 186 -194 234 -39
rect 420 -80 530 -66
rect 420 -83 498 -80
rect 420 -110 424 -83
rect 453 -107 498 -83
rect 527 -107 530 -80
rect 1151 -90 1186 -39
rect 1753 -21 2133 5
rect 2159 -21 2165 5
rect 1753 -29 2165 -21
rect 1753 -57 1785 -29
rect 2198 -49 2232 157
rect 1753 -77 1758 -57
rect 1779 -77 1785 -57
rect 1753 -84 1785 -77
rect 2176 -54 2232 -49
rect 2176 -74 2183 -54
rect 2203 -74 2232 -54
rect 2176 -81 2232 -74
rect 2176 -82 2211 -81
rect 453 -110 530 -107
rect 420 -125 530 -110
rect 1149 -95 1186 -90
rect 1149 -115 1156 -95
rect 1176 -115 1186 -95
rect 1149 -122 1186 -115
rect 2171 -120 2241 -110
rect 1149 -123 1184 -122
rect 186 -223 194 -194
rect 223 -223 234 -194
rect 186 -228 234 -223
rect 705 -188 737 -181
rect 705 -208 712 -188
rect 733 -208 737 -188
rect 705 -273 737 -208
rect 1075 -273 1115 -272
rect 705 -275 1117 -273
rect 705 -301 1085 -275
rect 1111 -301 1117 -275
rect 705 -309 1117 -301
rect 705 -337 737 -309
rect 1150 -329 1184 -123
rect 2169 -127 2241 -120
rect 1467 -155 1578 -133
rect 1467 -175 1475 -155
rect 1494 -175 1552 -155
rect 1571 -175 1578 -155
rect 1467 -192 1578 -175
rect 2169 -156 2176 -127
rect 2224 -156 2241 -127
rect 2169 -165 2241 -156
rect 2088 -256 2122 -255
rect 1219 -291 2123 -256
rect 705 -357 710 -337
rect 731 -357 737 -337
rect 705 -364 737 -357
rect 912 -337 951 -331
rect 912 -357 920 -337
rect 945 -357 951 -337
rect 912 -364 951 -357
rect 1128 -334 1184 -329
rect 1128 -354 1135 -334
rect 1155 -354 1184 -334
rect 1128 -361 1184 -354
rect 1128 -362 1163 -361
rect 920 -410 951 -364
rect 419 -435 530 -413
rect 419 -455 427 -435
rect 446 -455 504 -435
rect 523 -455 530 -435
rect 919 -427 951 -410
rect 1220 -427 1257 -291
rect 1358 -324 1468 -310
rect 1358 -327 1436 -324
rect 1358 -354 1362 -327
rect 1391 -351 1436 -327
rect 1465 -351 1468 -324
rect 2088 -334 2122 -291
rect 1391 -354 1468 -351
rect 1358 -369 1468 -354
rect 2087 -339 2122 -334
rect 2087 -359 2094 -339
rect 2114 -359 2122 -339
rect 2087 -367 2122 -359
rect 919 -440 1257 -427
rect 419 -472 530 -455
rect 920 -459 1257 -440
rect 1199 -460 1257 -459
rect 1643 -432 1675 -425
rect 1643 -452 1650 -432
rect 1671 -452 1675 -432
rect 1643 -517 1675 -452
rect 2013 -517 2053 -516
rect 1643 -519 2055 -517
rect 1643 -545 2023 -519
rect 2049 -545 2055 -519
rect 1643 -553 2055 -545
rect 189 -592 1185 -566
rect 1643 -581 1675 -553
rect 191 -645 233 -592
rect 191 -664 200 -645
rect 225 -664 233 -645
rect 191 -674 233 -664
rect 419 -634 529 -620
rect 419 -637 497 -634
rect 419 -664 423 -637
rect 452 -661 497 -637
rect 526 -661 529 -634
rect 1149 -644 1183 -592
rect 1643 -601 1648 -581
rect 1669 -601 1675 -581
rect 1643 -608 1675 -601
rect 1853 -580 1891 -570
rect 2088 -573 2122 -367
rect 1853 -597 1863 -580
rect 1883 -597 1891 -580
rect 1694 -640 1735 -639
rect 452 -664 529 -661
rect 419 -679 529 -664
rect 1148 -649 1183 -644
rect 1148 -669 1155 -649
rect 1175 -669 1183 -649
rect 1693 -650 1735 -640
rect 1148 -677 1183 -669
rect 704 -742 736 -735
rect 704 -762 711 -742
rect 732 -762 736 -742
rect 704 -827 736 -762
rect 1074 -827 1114 -826
rect 704 -829 1116 -827
rect 704 -855 1084 -829
rect 1110 -855 1116 -829
rect 704 -863 1116 -855
rect 704 -891 736 -863
rect 1149 -883 1183 -677
rect 1357 -679 1468 -657
rect 1357 -699 1365 -679
rect 1384 -699 1442 -679
rect 1461 -699 1468 -679
rect 1357 -716 1468 -699
rect 1693 -672 1700 -650
rect 1726 -672 1735 -650
rect 1693 -681 1735 -672
rect 910 -886 953 -884
rect 704 -911 709 -891
rect 730 -911 736 -891
rect 704 -918 736 -911
rect 909 -893 953 -886
rect 909 -913 919 -893
rect 942 -913 953 -893
rect 909 -917 953 -913
rect 1127 -888 1183 -883
rect 1127 -908 1134 -888
rect 1154 -908 1183 -888
rect 1127 -915 1183 -908
rect 1239 -747 1272 -746
rect 1693 -747 1730 -681
rect 1239 -776 1730 -747
rect 1127 -916 1162 -915
rect 418 -989 529 -967
rect 418 -1009 426 -989
rect 445 -1009 503 -989
rect 522 -1009 529 -989
rect 418 -1026 529 -1009
rect 909 -998 951 -917
rect 1239 -996 1272 -776
rect 1693 -778 1730 -776
rect 1499 -916 1609 -902
rect 1499 -919 1577 -916
rect 1499 -946 1503 -919
rect 1532 -943 1577 -919
rect 1606 -943 1609 -916
rect 1532 -946 1609 -943
rect 1499 -961 1609 -946
rect 1853 -935 1891 -597
rect 2066 -578 2122 -573
rect 2066 -598 2073 -578
rect 2093 -598 2122 -578
rect 2066 -605 2122 -598
rect 2066 -606 2101 -605
rect 1988 -706 2032 -702
rect 2169 -706 2219 -165
rect 1988 -739 2219 -706
rect 1988 -741 2195 -739
rect 1988 -895 2032 -741
rect 1853 -952 1861 -935
rect 1881 -952 1891 -935
rect 1853 -958 1891 -952
rect 1211 -998 1272 -996
rect 909 -1027 1272 -998
rect 1784 -1024 1816 -1017
rect 909 -1029 1211 -1027
rect 1784 -1044 1791 -1024
rect 1812 -1044 1816 -1024
rect 1784 -1109 1816 -1044
rect 1994 -1031 2032 -895
rect 2231 -926 2262 -925
rect 2228 -931 2262 -926
rect 2228 -951 2235 -931
rect 2255 -951 2262 -931
rect 2228 -959 2262 -951
rect 1994 -1069 2000 -1031
rect 2023 -1069 2032 -1031
rect 1994 -1079 2032 -1069
rect 2229 -1017 2262 -959
rect 2154 -1109 2194 -1108
rect 1784 -1111 2196 -1109
rect 1152 -1115 1187 -1113
rect 188 -1118 1187 -1115
rect 187 -1142 1187 -1118
rect 187 -1297 235 -1142
rect 421 -1183 531 -1169
rect 421 -1186 499 -1183
rect 421 -1213 425 -1186
rect 454 -1210 499 -1186
rect 528 -1210 531 -1183
rect 1152 -1193 1187 -1142
rect 454 -1213 531 -1210
rect 421 -1228 531 -1213
rect 1150 -1198 1187 -1193
rect 1150 -1218 1157 -1198
rect 1177 -1218 1187 -1198
rect 1784 -1137 2164 -1111
rect 2190 -1137 2196 -1111
rect 1784 -1145 2196 -1137
rect 1784 -1173 1816 -1145
rect 2229 -1165 2265 -1017
rect 1784 -1193 1789 -1173
rect 1810 -1193 1816 -1173
rect 1784 -1200 1816 -1193
rect 2207 -1170 2265 -1165
rect 2207 -1190 2214 -1170
rect 2234 -1190 2265 -1170
rect 2207 -1197 2265 -1190
rect 2207 -1198 2242 -1197
rect 1150 -1225 1187 -1218
rect 1150 -1226 1185 -1225
rect 187 -1326 195 -1297
rect 224 -1326 235 -1297
rect 187 -1331 235 -1326
rect 706 -1291 738 -1284
rect 706 -1311 713 -1291
rect 734 -1311 738 -1291
rect 706 -1376 738 -1311
rect 1076 -1376 1116 -1375
rect 706 -1378 1118 -1376
rect 706 -1404 1086 -1378
rect 1112 -1404 1118 -1378
rect 706 -1412 1118 -1404
rect 706 -1440 738 -1412
rect 1151 -1432 1185 -1226
rect 1855 -1243 1894 -1236
rect 1498 -1271 1609 -1249
rect 1498 -1291 1506 -1271
rect 1525 -1291 1583 -1271
rect 1602 -1291 1609 -1271
rect 1498 -1308 1609 -1291
rect 1855 -1270 1859 -1243
rect 1890 -1270 1894 -1243
rect 1702 -1359 1755 -1355
rect 1220 -1394 1755 -1359
rect 706 -1460 711 -1440
rect 732 -1460 738 -1440
rect 706 -1467 738 -1460
rect 913 -1440 952 -1434
rect 913 -1460 921 -1440
rect 946 -1460 952 -1440
rect 913 -1467 952 -1460
rect 1129 -1437 1185 -1432
rect 1129 -1457 1136 -1437
rect 1156 -1457 1185 -1437
rect 1129 -1464 1185 -1457
rect 1129 -1465 1164 -1464
rect 921 -1513 952 -1467
rect 420 -1538 531 -1516
rect 420 -1558 428 -1538
rect 447 -1558 505 -1538
rect 524 -1558 531 -1538
rect 920 -1530 952 -1513
rect 1221 -1530 1258 -1394
rect 1359 -1427 1469 -1413
rect 1359 -1430 1437 -1427
rect 1359 -1457 1363 -1430
rect 1392 -1454 1437 -1430
rect 1466 -1454 1469 -1427
rect 1392 -1457 1469 -1454
rect 1359 -1472 1469 -1457
rect 1701 -1441 1755 -1394
rect 1701 -1449 1754 -1441
rect 1701 -1466 1710 -1449
rect 1742 -1466 1754 -1449
rect 1701 -1469 1754 -1466
rect 920 -1543 1258 -1530
rect 420 -1575 531 -1558
rect 921 -1562 1258 -1543
rect 1200 -1563 1258 -1562
rect 1644 -1535 1676 -1528
rect 1644 -1555 1651 -1535
rect 1672 -1555 1676 -1535
rect 1644 -1620 1676 -1555
rect 1855 -1543 1894 -1270
rect 2090 -1441 2124 -1430
rect 2088 -1442 2124 -1441
rect 2088 -1462 2095 -1442
rect 2115 -1462 2124 -1442
rect 2088 -1470 2124 -1462
rect 1855 -1584 1862 -1543
rect 1883 -1584 1894 -1543
rect 1855 -1599 1894 -1584
rect 2014 -1620 2054 -1619
rect 1644 -1622 2056 -1620
rect 1644 -1648 2024 -1622
rect 2050 -1648 2056 -1622
rect 1644 -1656 2056 -1648
rect 190 -1695 1186 -1669
rect 1644 -1684 1676 -1656
rect 2089 -1676 2123 -1470
rect 192 -1748 234 -1695
rect 192 -1767 201 -1748
rect 226 -1767 234 -1748
rect 192 -1777 234 -1767
rect 420 -1737 530 -1723
rect 420 -1740 498 -1737
rect 420 -1767 424 -1740
rect 453 -1764 498 -1740
rect 527 -1764 530 -1737
rect 1150 -1747 1184 -1695
rect 1644 -1704 1649 -1684
rect 1670 -1704 1676 -1684
rect 1644 -1711 1676 -1704
rect 2067 -1681 2123 -1676
rect 2067 -1701 2074 -1681
rect 2094 -1701 2123 -1681
rect 2067 -1708 2123 -1701
rect 2067 -1709 2102 -1708
rect 1695 -1743 1736 -1742
rect 453 -1767 530 -1764
rect 420 -1782 530 -1767
rect 1149 -1752 1184 -1747
rect 1149 -1772 1156 -1752
rect 1176 -1772 1184 -1752
rect 1694 -1753 1736 -1743
rect 1149 -1780 1184 -1772
rect 705 -1845 737 -1838
rect 705 -1865 712 -1845
rect 733 -1865 737 -1845
rect 705 -1930 737 -1865
rect 1075 -1930 1115 -1929
rect 705 -1932 1117 -1930
rect 705 -1958 1085 -1932
rect 1111 -1958 1117 -1932
rect 705 -1966 1117 -1958
rect 705 -1994 737 -1966
rect 1150 -1986 1184 -1780
rect 1358 -1782 1469 -1760
rect 1358 -1802 1366 -1782
rect 1385 -1802 1443 -1782
rect 1462 -1802 1469 -1782
rect 1358 -1819 1469 -1802
rect 1694 -1775 1701 -1753
rect 1727 -1775 1736 -1753
rect 1694 -1784 1736 -1775
rect 911 -1989 954 -1987
rect 705 -2014 710 -1994
rect 731 -2014 737 -1994
rect 705 -2021 737 -2014
rect 910 -1996 954 -1989
rect 910 -2016 920 -1996
rect 943 -2016 954 -1996
rect 910 -2020 954 -2016
rect 1128 -1991 1184 -1986
rect 1128 -2011 1135 -1991
rect 1155 -2011 1184 -1991
rect 1128 -2018 1184 -2011
rect 1240 -1850 1273 -1849
rect 1694 -1850 1731 -1784
rect 1240 -1879 1731 -1850
rect 1128 -2019 1163 -2018
rect 419 -2092 530 -2070
rect 419 -2112 427 -2092
rect 446 -2112 504 -2092
rect 523 -2112 530 -2092
rect 419 -2129 530 -2112
rect 910 -2101 952 -2020
rect 1240 -2099 1273 -1879
rect 1694 -1881 1731 -1879
rect 1212 -2101 1273 -2099
rect 910 -2130 1273 -2101
rect 910 -2132 1212 -2130
<< labels >>
rlabel locali 290 1907 312 1922 1 d0
rlabel metal1 459 2130 487 2135 1 vdd
rlabel metal1 456 1737 490 1743 1 gnd
rlabel locali 1227 1659 1255 1680 1 d1
rlabel metal1 1394 1493 1428 1499 1 gnd
rlabel metal1 1397 1886 1425 1891 1 vdd
rlabel locali 289 1353 311 1368 1 d0
rlabel metal1 458 1576 486 1581 1 vdd
rlabel metal1 455 1183 489 1189 1 gnd
rlabel locali 110 2192 138 2200 1 vref
rlabel locali 291 804 313 819 1 d0
rlabel metal1 460 1027 488 1032 1 vdd
rlabel metal1 457 634 491 640 1 gnd
rlabel locali 1228 556 1256 577 1 d1
rlabel metal1 1395 390 1429 396 1 gnd
rlabel metal1 1398 783 1426 788 1 vdd
rlabel locali 290 250 312 265 1 d0
rlabel metal1 459 473 487 478 1 vdd
rlabel metal1 456 80 490 86 1 gnd
rlabel metal1 1538 1294 1566 1299 1 vdd
rlabel metal1 1535 901 1569 907 1 gnd
rlabel locali 1366 1066 1387 1085 1 d2
rlabel locali 291 -299 313 -284 1 d0
rlabel metal1 460 -76 488 -71 1 vdd
rlabel metal1 457 -469 491 -463 1 gnd
rlabel locali 1228 -547 1256 -526 1 d1
rlabel metal1 1395 -713 1429 -707 1 gnd
rlabel metal1 1398 -320 1426 -315 1 vdd
rlabel locali 290 -853 312 -838 1 d0
rlabel metal1 459 -630 487 -625 1 vdd
rlabel metal1 456 -1023 490 -1017 1 gnd
rlabel locali 292 -1402 314 -1387 1 d0
rlabel metal1 461 -1179 489 -1174 1 vdd
rlabel metal1 458 -1572 492 -1566 1 gnd
rlabel locali 1229 -1650 1257 -1629 1 d1
rlabel metal1 1396 -1816 1430 -1810 1 gnd
rlabel metal1 1399 -1423 1427 -1418 1 vdd
rlabel locali 291 -1956 313 -1941 1 d0
rlabel metal1 460 -1733 488 -1728 1 vdd
rlabel metal1 457 -2126 491 -2120 1 gnd
rlabel metal1 1539 -912 1567 -907 1 vdd
rlabel metal1 1536 -1305 1570 -1299 1 gnd
rlabel locali 1367 -1140 1388 -1121 1 d2
rlabel locali 1969 16 1991 31 1 vout
rlabel metal1 1508 204 1536 209 1 vdd
rlabel metal1 1505 -189 1539 -183 1 gnd
rlabel locali 1338 -20 1364 -3 1 d3
<< end >>
