* SPICE3 file created from 9bit_DAC.ext - technology: sky130A

.option scale=10000u

X0 a_31071_8063# a_30650_8063# a_30334_8173# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1 a_39098_4304# a_39094_4481# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2 a_15943_951# a_16674_1261# a_16882_1261# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3 a_12776_8427# a_13029_8414# a_12807_7311# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4 a_853_7523# a_432_7523# a_117_7728# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5 vdd d0 a_4080_2612# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6 a_34038_5543# a_34043_4817# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7 a_10150_3967# a_10677_4219# a_10885_4219# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8 a_854_4214# a_433_4214# a_119_3962# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9 a_11825_2323# a_11758_1731# a_11836_2847# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X10 a_26098_3687# a_25677_3687# a_25361_3797# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X11 a_6864_7414# a_6567_8385# a_6848_7874# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X12 a_7938_8048# a_8195_7858# a_7797_8640# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X13 vdd d0 a_24267_1490# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X14 a_35392_2240# a_35393_1783# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X15 vdd a_14111_2617# a_13903_2617# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X16 vdd a_33215_8395# a_33007_8395# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X17 gnd d1 a_28383_2324# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X18 a_12919_2320# a_13903_2617# a_13854_2807# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X19 a_8878_3392# a_8883_2666# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X20 gnd a_9132_8717# a_8924_8717# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X21 a_19317_134# a_19208_134# vout vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X22 a_6738_387# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X23 a_35708_3692# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X24 a_5173_6666# a_5701_6461# a_5909_6461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X25 a_21041_4749# a_20620_4749# a_20304_4859# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X26 a_23074_2296# a_24058_2593# a_24013_2606# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X27 a_2778_2894# a_3031_2881# a_2774_5271# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X28 a_12778_4015# a_12963_4513# a_12918_4526# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X29 vdd a_33218_1777# a_33010_1777# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X30 a_10149_4654# a_10149_4424# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X31 a_30074_191# a_29965_191# a_19317_134# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X32 a_20620_5852# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X33 a_27989_4032# a_28174_4530# a_28125_4720# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X34 a_117_7958# a_117_7728# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X35 a_10884_6425# a_10463_6425# a_10148_6630# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X36 a_25675_5339# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X37 a_21981_1196# a_21560_1196# a_21043_1440# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X38 gnd d0 a_19167_1001# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X39 a_15942_5917# a_15521_5917# a_15205_5798# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X40 a_13859_1527# a_13855_1704# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X41 a_5909_9221# a_6639_8977# a_6847_8977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X42 vdd d1 a_28381_6736# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X43 a_8884_1563# a_9137_1550# a_7945_1253# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X44 a_5176_1151# a_5178_1052# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X45 a_15940_9226# a_15519_9226# a_15203_9336# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X46 a_855_3111# a_434_3111# a_119_3316# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X47 a_35392_3573# a_35921_3692# a_36129_3692# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X48 gnd d0 a_34295_7010# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X49 a_13856_4282# a_13852_4459# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X50 a_24007_8298# a_24010_7567# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X51 a_39095_2275# a_39352_2085# a_38157_2519# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X52 vdd a_29322_3737# a_29114_3737# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X53 gnd d0 a_14110_5926# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X54 a_11823_6735# a_11402_6735# a_10884_6425# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X55 vdd a_23325_6695# a_23117_6695# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X56 a_25891_1481# a_25678_1481# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X57 a_27987_8444# a_28172_8942# a_28127_8955# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X58 a_38045_7510# a_38064_6230# a_38019_6243# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X59 a_26614_5649# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X60 a_16769_392# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X61 a_35392_3802# a_35392_3573# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X62 a_34040_2788# a_34297_2598# a_33105_2301# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X63 a_11713_351# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X64 a_26612_8958# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X65 vdd d0 a_24262_8657# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X66 a_31069_8612# a_30648_8612# a_30334_8360# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X67 a_3820_7763# a_3825_7037# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X68 a_8878_6152# a_9135_5962# a_7943_5665# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X69 gnd a_33357_5597# a_33149_5597# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X70 a_1895_346# a_1682_346# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X71 a_12134_351# a_14876_331# a_9888_210# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X72 a_28125_5823# a_29112_5389# a_29067_5402# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X73 a_5174_4460# a_5175_4003# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X74 a_2888_3418# a_3141_3405# a_2743_4187# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X75 a_20622_1440# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X76 a_10886_2013# a_10465_2013# a_10150_2218# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X77 a_38047_3098# a_38304_2908# a_38047_5298# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X78 gnd d3 a_33246_7279# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X79 gnd d1 a_18226_6760# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X80 a_5490_3152# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X81 a_25677_927# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X82 a_12772_8604# a_13029_8414# a_12807_7311# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X83 a_5909_7564# a_6640_7874# a_6848_7874# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X84 a_27045_7276# a_26754_6160# a_27034_6752# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X85 a_5053_326# a_4632_326# a_4954_326# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X86 gnd d0 a_29323_1531# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X87 a_15944_1505# a_15523_1505# a_15207_1386# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X88 a_5911_4809# a_6641_4565# a_6849_4565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X89 vdd d2 a_33217_3983# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X90 gnd d1 a_3139_6714# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X91 gnd a_29322_977# a_29114_977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X92 a_31590_2304# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X93 vdd d1 a_28383_2324# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X94 a_15204_7130# a_15204_6901# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X95 a_28130_2337# a_29114_2634# a_29065_2824# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X96 a_11824_5632# a_11403_5632# a_10886_5876# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X97 a_855_4768# a_434_4768# a_118_4878# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X98 vdd a_8087_2922# a_7879_2922# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X99 a_30649_9166# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X100 a_26966_8366# a_26753_8366# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X101 a_15519_6466# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X102 a_29066_6505# a_29319_6492# a_28124_6926# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X103 a_11834_5059# a_11725_5059# a_11933_5059# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X104 a_32959_6379# a_33149_5597# a_33104_5610# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X105 a_27989_4032# a_28174_4530# a_28129_4543# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X106 a_15207_1615# a_15207_1386# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X107 a_11825_2323# a_11404_2323# a_10886_2013# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X108 a_26616_1237# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X109 a_29068_2093# a_29064_2270# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X110 a_119_2859# a_119_2672# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X111 a_26095_6442# a_25674_6442# a_25359_6647# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X112 vdd d0 a_29321_5943# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X113 a_24008_3332# a_24013_2606# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X114 gnd a_33359_1185# a_33151_1185# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X115 a_21697_8325# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X116 a_8880_1740# a_9137_1550# a_7945_1253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X117 a_37066_5654# a_36998_6165# a_37076_7281# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X118 a_20304_5503# a_20832_5298# a_21040_5298# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X119 a_16895_7419# a_16598_8390# a_16878_8982# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X120 a_5911_3152# a_6642_3462# a_6850_3462# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X121 gnd d3 a_33248_2867# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X122 a_2776_7306# a_2790_8409# a_2741_8599# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X123 vdd d0 a_34295_7010# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X124 vdd a_24265_5902# a_24057_5902# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X125 a_7939_5842# a_8926_5408# a_8877_5598# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X126 a_18911_1745# a_18914_1014# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X127 a_20303_8355# a_20303_8168# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X128 a_2741_8599# a_2931_7817# a_2882_8007# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X129 a_36127_7001# a_35706_7001# a_35390_6882# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X130 a_15205_4924# a_15205_4695# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X131 a_10465_4773# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X132 vdd a_9134_4305# a_8926_4305# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X133 a_10150_3967# a_10150_3780# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X134 a_20834_3646# a_20621_3646# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X135 a_5702_5358# a_5489_5358# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X136 a_20832_6955# a_20619_6955# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X137 a_1805_2842# a_1514_1726# a_1794_2318# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X138 a_5703_2049# a_5490_2049# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X139 a_31700_2828# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X140 a_10677_5322# a_10464_5322# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X141 a_6537_5095# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X142 a_31802_4510# a_31589_4510# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X143 a_26968_3954# a_26755_3954# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X144 a_3823_2802# a_3826_2071# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X145 vdd d1 a_18226_6760# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X146 vdd d0 a_29323_1531# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X147 a_11834_5059# a_11514_2847# a_11836_2847# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X148 a_15733_8123# a_15520_8123# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X149 vdd d1 a_3139_6714# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X150 a_21699_3913# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X151 a_16458_7879# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X152 vdd d2 a_13030_6208# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X153 a_6641_5668# a_6428_5668# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X154 a_28020_5116# a_28273_5103# a_27246_368# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X155 a_25362_1591# a_25362_1362# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X156 a_12777_6221# a_12962_6719# a_12913_6909# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X157 vdd a_13170_6719# a_12962_6719# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X158 a_2778_2894# a_2792_3997# a_2743_4187# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X159 a_2748_1804# a_3001_1791# a_2774_3071# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X160 a_28130_2337# a_29114_2634# a_29069_2647# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X161 vdd a_24267_1490# a_24059_1490# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X162 a_7941_1430# a_8928_996# a_8879_1186# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X163 a_30336_2845# a_30336_2658# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X164 a_10148_8192# a_10677_8082# a_10885_8082# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X165 a_5704_946# a_5491_946# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X166 a_645_9180# a_432_9180# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X167 a_15941_4260# a_15520_4260# a_15206_4008# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X168 a_21040_5298# a_20619_5298# a_20304_5503# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X169 vdd a_33359_1185# a_33151_1185# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X170 a_10677_6979# a_10464_6979# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X171 gnd a_19167_1001# a_18959_1001# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X172 vdd d1 a_18228_2348# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X173 a_7943_5665# a_8196_5652# a_7798_6434# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X174 vdd d1 a_3141_2302# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X175 a_38049_7333# a_38063_8436# a_38014_8626# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X176 a_6643_1256# a_6430_1256# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X177 a_39096_2829# a_39353_2639# a_38161_2342# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X178 gnd a_34295_7010# a_34087_7010# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X179 a_21557_6711# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X180 a_32119_5040# a_31698_5040# a_32020_5040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X181 a_36127_4241# a_36858_4551# a_37066_4551# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X182 a_1724_8344# a_1511_8344# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X183 a_3824_6483# a_4077_6470# a_2882_6904# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X184 a_21868_327# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X185 vdd d0 a_19166_5967# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X186 a_20304_5962# a_20304_5733# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X187 a_11824_4529# a_11757_3937# a_11841_2966# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X188 vdd a_24262_8657# a_24054_8657# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X189 vdd a_14110_4823# a_13902_4823# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X190 vdd d0 a_24266_3696# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X191 a_10678_5876# a_10465_5876# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X192 a_21042_886# a_20621_886# a_20306_1091# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X193 a_25678_1481# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X194 a_8879_2843# a_8882_2112# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X195 a_27045_5076# a_26725_2864# a_27047_2864# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X196 gnd a_33246_7279# a_33038_7279# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X197 gnd a_18226_6760# a_18018_6760# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X198 a_35707_5898# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X199 a_10679_2567# a_10466_2567# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X200 a_5172_8872# a_5700_8667# a_5908_8667# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X201 gnd a_29323_1531# a_29115_1531# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X202 a_7945_1253# a_8198_1240# a_7800_2022# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X203 vdd a_33217_3983# a_33009_3983# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X204 a_16880_5673# a_16459_5673# a_15942_5917# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X205 a_30862_9166# a_30649_9166# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X206 a_24007_8298# a_24264_8108# a_23072_7811# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X207 a_27988_6238# a_28173_6736# a_28124_6926# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X208 a_38051_2921# a_38065_4024# a_38016_4214# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X209 a_18914_3774# a_18910_3951# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X210 a_16881_2364# a_16460_2364# a_15942_2054# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X211 a_38015_6420# a_38205_5638# a_38160_5651# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X212 vdd a_28383_3427# a_28175_3427# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X213 gnd d0 a_19166_3207# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X214 a_117_8187# a_117_7958# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X215 a_18911_6529# a_18907_6706# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X216 gnd d0 a_24263_6451# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X217 a_26753_8366# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X218 a_2778_5094# a_2821_7293# a_2772_7483# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X219 a_1726_3932# a_1513_3932# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X220 a_8883_3769# a_9136_3756# a_7944_3459# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X221 a_25359_8209# a_25359_7980# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X222 a_854_5317# a_433_5317# a_118_5522# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X223 gnd d3 a_38304_2908# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X224 gnd d0 a_34294_9216# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X225 a_117_7084# a_646_6974# a_854_6974# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X226 gnd d2 a_33218_1777# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X227 a_6859_7295# a_6568_6179# a_6849_5668# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X228 a_7939_5842# a_8196_5652# a_7798_6434# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X229 a_35920_2035# a_35707_2035# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X230 a_855_2008# a_434_2008# a_120_1756# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X231 a_20304_5962# a_20833_5852# a_21041_5852# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X232 a_38049_7333# a_38063_8436# a_38018_8449# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X233 a_25890_3687# a_25677_3687# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X234 a_5173_7312# a_5701_7564# a_5909_7564# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X235 a_35709_1486# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X236 gnd a_33248_2867# a_33040_2867# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X237 vdd d2 a_2998_8409# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X238 a_5174_4460# a_5702_4255# a_5910_4255# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X239 a_34039_4994# a_34296_4804# a_33104_4507# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X240 a_20302_9042# a_20831_9161# a_21039_9161# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X241 a_37065_7860# a_36644_7860# a_36126_7550# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X242 vdd a_34295_7010# a_34087_7010# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X243 a_6861_2883# a_6570_1767# a_6850_2359# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X244 a_38158_8960# a_39142_9257# gnd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X245 a_30863_8063# a_30650_8063# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X246 a_31070_6406# a_31801_6716# a_32009_6716# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X247 a_30335_5738# a_30335_5508# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X248 a_16882_1261# a_16461_1261# a_15944_1505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X249 a_28124_8029# a_29111_7595# a_29066_7608# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X250 a_3820_6660# a_4077_6470# a_2882_6904# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X251 a_10885_4219# a_10464_4219# a_10149_4424# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X252 a_20621_3646# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X253 a_19317_134# a_29752_191# a_30074_191# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X254 a_11836_2847# a_11545_1731# a_11826_1220# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X255 a_27990_1826# a_28175_2324# a_28126_2514# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X256 a_7797_8640# a_7987_7858# a_7942_7871# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X257 a_5704_2603# a_5491_2603# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X258 a_16568_5100# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X259 gnd d0 a_29322_3737# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X260 a_5490_2049# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X261 a_16890_5100# a_16570_2888# a_16892_2888# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X262 a_10464_5322# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X263 a_26755_3954# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X264 a_31899_332# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X265 gnd d2 a_13029_8414# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X266 a_5909_6461# a_5488_6461# a_5174_6209# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X267 a_25360_6003# a_25360_5774# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X268 a_32320_332# a_35062_312# a_30074_191# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X269 a_21669_2823# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X270 a_2774_5271# a_2823_2881# a_2774_3071# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X271 a_15941_7020# a_15520_7020# a_15204_7130# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X272 a_21994_7354# a_21880_7235# a_21994_5154# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X273 a_118_5752# a_647_5871# a_855_5871# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X274 a_15205_4695# a_15734_4814# a_15942_4814# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X275 vdd a_18226_6760# a_18018_6760# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X276 a_35393_1367# a_35922_1486# a_36130_1486# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X277 a_856_905# a_435_905# a_120_1110# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X278 vdd a_29323_1531# a_29115_1531# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X279 a_7941_1430# a_8198_1240# a_7800_2022# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X280 a_119_2672# a_648_2562# a_856_2562# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X281 a_25358_8853# a_25359_8396# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X282 a_11823_7838# a_11402_7838# a_10885_8082# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X283 a_15520_8123# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X284 a_29065_8711# a_29318_8698# a_28123_9132# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X285 a_32958_8585# a_33148_7803# a_33103_7816# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X286 a_27988_6238# a_28173_6736# a_28128_6749# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X287 a_11824_4529# a_11403_4529# a_10885_4219# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X288 a_38051_2921# a_38065_4024# a_38020_4037# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X289 a_5175_2900# a_5703_3152# a_5911_3152# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X290 a_6750_7295# a_6537_7295# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X291 a_7945_1253# a_8929_1550# a_8880_1740# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X292 a_26094_8648# a_25673_8648# a_25358_8853# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X293 a_33103_6713# a_34087_7010# a_34038_7200# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X294 vdd d0 a_24263_6451# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X295 a_31072_1994# a_31803_2304# a_32011_2304# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X296 a_39093_7790# a_39350_7600# a_38155_8034# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X297 a_32221_332# a_33040_5067# a_32995_5080# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X298 a_8879_3946# a_9136_3756# a_7944_3459# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X299 a_2889_1212# a_3142_1199# a_2744_1981# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X300 a_3822_2248# a_4079_2058# a_2884_2492# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X301 a_5491_946# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X302 a_5910_5358# a_6641_5668# a_6849_5668# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X303 gnd d1 a_18227_4554# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X304 a_432_9180# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X305 vdd d0 a_34294_9216# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X306 a_34038_4440# a_34044_3714# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X307 a_5912_2603# a_6642_2359# a_6850_2359# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X308 a_31944_1712# a_31731_1712# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X309 a_19208_134# a_18995_134# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X310 a_36126_9207# a_35705_9207# a_35389_9088# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X311 a_10464_6979# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X312 a_13852_7219# a_14109_7029# a_12917_6732# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X313 a_8882_4872# a_8878_5049# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X314 a_8878_2289# a_8884_1563# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X315 gnd a_13171_4513# a_12963_4513# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X316 a_37175_5081# a_36754_5081# a_37076_5081# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X317 vdd a_18228_2348# a_18020_2348# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X318 a_7943_5665# a_8927_5962# a_8882_5975# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X319 a_2743_4187# a_2933_3405# a_2884_3595# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X320 gnd a_39349_8703# a_39141_8703# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X321 a_7832_7347# a_8085_7334# a_7834_5135# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X322 a_15519_7569# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X323 a_10676_7528# a_10463_7528# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X324 a_26967_6160# a_26754_6160# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X325 a_11825_3426# a_11404_3426# a_10887_3670# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X326 a_27990_1826# a_28175_2324# a_28130_2337# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X327 a_117_6855# a_117_6625# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X328 a_6430_1256# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X329 vdd d1 a_18225_8966# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X330 a_35390_8401# a_35917_8653# a_36125_8653# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X331 a_39097_7613# a_39093_7790# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X332 a_6752_2883# a_6539_2883# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X333 a_26096_4236# a_25675_4236# a_25360_4441# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X334 vdd d0 a_24265_2039# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X335 a_1511_8344# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X336 a_21698_6119# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X337 a_35391_5549# a_35391_5092# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X338 a_21041_1989# a_20620_1989# a_20306_1737# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X339 a_39095_3378# a_39352_3188# a_38157_3622# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X340 vdd d2 a_13029_8414# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X341 vdd a_19166_5967# a_18958_5967# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X342 a_37067_3448# a_36999_3959# a_37083_2988# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X343 vdd a_13169_8925# a_12961_8925# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X344 a_5912_946# a_6643_1256# a_6851_1256# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X345 vdd a_24266_3696# a_24058_3696# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X346 a_32022_2828# a_31913_2828# a_32020_5040# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X347 a_36127_8104# a_35706_8104# a_35390_8214# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X348 a_11933_5059# a_11512_5059# a_11839_5178# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X349 a_29063_8339# a_29320_8149# a_28128_7852# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X350 a_24007_7195# a_24010_6464# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X351 a_10465_5876# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X352 a_10148_7963# a_10148_7733# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X353 a_25887_6442# a_25674_6442# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X354 gnd a_28382_5633# a_28174_5633# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X355 a_35392_2699# a_35392_2470# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X356 a_10466_2567# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X357 a_25890_927# a_25677_927# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X358 gnd d3 a_28271_7315# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X359 a_15940_6466# a_15519_6466# a_15205_6214# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X360 gnd d0 a_29319_6492# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X361 a_7945_1253# a_8929_1550# a_8884_1563# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X362 a_33103_6713# a_34087_7010# a_34042_7023# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X363 a_10678_3116# a_10465_3116# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X364 a_6782_3973# a_6569_3973# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X365 gnd a_39351_4291# a_39143_4291# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X366 gnd d0 a_19167_3761# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X367 a_7834_2935# a_8087_2922# a_7830_5312# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X368 a_3820_6660# a_3826_5934# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X369 a_20618_6401# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X370 a_1696_2842# a_1483_2842# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X371 vdd d1 a_18227_4554# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X372 gnd a_19166_3207# a_18958_3207# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X373 a_35919_7001# a_35706_7001# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X374 a_35392_3989# a_35919_4241# a_36127_4241# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X375 gnd a_14111_2617# a_13903_2617# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X376 a_13855_7591# a_13851_7768# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X377 gnd a_24263_6451# a_24055_6451# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X378 a_854_6974# a_1584_6730# a_1792_6730# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X379 a_25360_6003# a_25889_5893# a_26097_5893# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X380 a_1513_3932# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X381 a_26826_6752# a_26613_6752# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X382 vdd d2 a_13031_4002# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X383 vdd d0 a_29322_977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X384 a_39095_5035# a_39352_4845# a_38160_4548# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X385 a_29065_1167# a_29322_977# a_28127_1411# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X386 a_17976_1258# a_18960_1555# a_18911_1745# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X387 gnd a_38304_2908# a_38096_2908# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X388 gnd a_34294_9216# a_34086_9216# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X389 vdd a_13171_4513# a_12963_4513# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X390 gnd a_33218_1777# a_33010_1777# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X391 gnd d1 a_33356_6700# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X392 a_36126_6447# a_36857_6757# a_37065_6757# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X393 a_10467_1464# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X394 a_3823_8689# a_4076_8676# a_2881_9110# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X395 a_7828_7524# a_8085_7334# a_7834_5135# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X396 a_38016_4214# a_38206_3432# a_38157_3622# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X397 a_117_7728# a_645_7523# a_853_7523# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X398 gnd a_28384_1221# a_28176_1221# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X399 vdd a_2998_8409# a_2790_8409# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X400 a_5173_7769# a_5173_7312# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X401 a_15941_5363# a_15520_5363# a_15205_5568# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X402 vdd d4 a_38304_5108# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X403 a_30650_8063# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X404 a_24008_2229# a_24014_1503# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X405 gnd d0 a_29321_2080# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X406 a_15942_2054# a_15521_2054# a_15207_1802# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X407 a_25677_3687# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X408 a_34040_3891# a_34043_3160# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X409 a_27050_7395# a_26936_7276# a_27050_5195# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X410 a_5491_2603# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X411 a_7944_3459# a_8197_3446# a_7799_4228# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X412 gnd a_29322_3737# a_29114_3737# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X413 a_6951_387# a_6738_387# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X414 a_35171_312# a_36955_373# a_37175_5081# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X415 a_10885_8082# a_10464_8082# a_10148_7963# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X416 a_25362_1591# a_25891_1481# a_26099_1481# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X417 a_26828_2340# a_26615_2340# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X418 a_38014_8626# a_38204_7844# a_38159_7857# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X419 vdd a_28382_5633# a_28174_5633# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X420 a_27144_5076# a_26723_5076# a_27050_5195# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X421 a_10150_2864# a_10150_2677# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X422 a_22088_5035# a_22081_327# a_22289_327# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X423 a_38159_6754# a_39143_7051# a_39094_7241# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X424 a_29067_5402# a_29063_5579# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X425 a_21558_4505# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X426 gnd d0 a_24262_8657# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X427 vdd d0 a_34294_7559# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X428 vdd d3 a_28271_7315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X429 a_36128_2035# a_36859_2345# a_37067_2345# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X430 a_1725_6138# a_1512_6138# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X431 a_7798_6434# a_7988_5652# a_7939_5842# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X432 a_3825_4277# a_4078_4264# a_2883_4698# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X433 vdd d0 a_19167_3761# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X434 gnd d1 a_13173_1204# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X435 a_25361_3338# a_25361_2881# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X436 a_119_3316# a_647_3111# a_855_3111# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X437 a_36126_7550# a_35705_7550# a_35390_7298# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X438 vdd a_3000_3997# a_2792_3997# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X439 a_15943_951# a_15522_951# a_15207_1156# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X440 a_37000_1753# a_36787_1753# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X441 vdd a_24263_6451# a_24055_6451# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X442 a_13855_9248# a_14108_9235# a_12916_8938# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X443 a_11725_7259# a_11512_7259# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X444 gnd d0 a_34296_4804# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X445 a_10679_3670# a_10466_3670# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X446 a_10679_910# a_10466_910# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X447 a_16457_8982# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X448 a_35389_9317# a_35389_9088# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X449 gnd a_18227_4554# a_18019_4554# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X450 a_20832_4195# a_20619_4195# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X451 a_17976_1258# a_18960_1555# a_18915_1568# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X452 a_25239_307# a_24818_307# a_22289_327# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X453 vdd a_34294_9216# a_34086_9216# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X454 a_2882_6904# a_3869_6470# a_3820_6660# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X455 a_32962_8408# a_33215_8395# a_32993_7292# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X456 a_16881_3467# a_16460_3467# a_15943_3711# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X457 a_31731_1712# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X458 a_38047_3098# a_38066_1818# a_38017_2008# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X459 a_3819_8866# a_4076_8676# a_2881_9110# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X460 a_11841_2966# a_11544_3937# a_11825_3426# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X461 a_38016_4214# a_38206_3432# a_38161_3445# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X462 a_5703_4809# a_5490_4809# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X463 vdd a_28384_1221# a_28176_1221# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X464 a_16982_392# a_16769_392# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X465 a_3822_6111# a_3825_5380# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X466 vdd d0 a_24266_936# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X467 gnd d1 a_8195_7858# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X468 gnd d0 a_24264_4245# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X469 a_24009_1126# a_24266_936# a_23071_1370# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X470 vdd d0 a_29321_2080# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X471 a_26938_2864# a_26725_2864# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X472 a_5908_8667# a_5487_8667# a_5173_8415# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X473 a_10463_7528# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X474 a_26754_6160# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X475 vdd d0 a_34296_3147# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X476 vdd a_18225_8966# a_18017_8966# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X477 a_118_4878# a_647_4768# a_855_4768# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X478 a_32112_332# a_31899_332# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X479 a_20306_1550# a_20306_1321# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X480 a_37078_2869# a_36969_2869# a_37076_5081# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X481 a_7940_3636# a_8197_3446# a_7799_4228# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X482 a_120_1340# a_120_1110# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X483 a_17861_3117# a_17880_1837# a_17835_1850# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X484 gnd a_3139_7817# a_2931_7817# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X485 vdd a_24265_2039# a_24057_2039# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X486 a_20303_7709# a_20303_7252# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X487 a_5174_5106# a_5702_5358# a_5910_5358# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X488 a_5175_2254# a_5703_2049# a_5911_2049# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X489 a_20303_6836# a_20832_6955# a_21040_6955# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X490 a_37066_5654# a_36645_5654# a_36127_5344# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X491 a_7944_3459# a_8928_3756# a_8879_3946# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X492 a_38047_5298# a_38096_2908# a_38047_3098# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X493 a_33102_8919# a_34086_9216# a_34037_9406# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X494 a_38159_6754# a_39143_7051# a_39098_7064# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X495 a_32964_3996# a_33217_3983# a_32995_2880# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X496 a_23072_6708# a_23325_6695# a_22932_6197# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X497 a_31071_4200# a_31802_4510# a_32010_4510# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X498 a_25674_6442# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X499 a_3821_4454# a_4078_4264# a_2883_4698# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X500 a_5704_3706# a_5491_3706# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X501 a_24010_1680# a_24013_949# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X502 a_37064_8963# a_36643_8963# a_36126_9207# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X503 a_7798_6434# a_7988_5652# a_7943_5665# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X504 a_8877_8358# a_8880_7627# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X505 a_20304_4859# a_20304_4630# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X506 a_15204_8233# a_15733_8123# a_15941_8123# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X507 a_5909_7564# a_5488_7564# a_5173_7769# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X508 a_21772_2299# a_21559_2299# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X509 a_10465_3116# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X510 a_31943_3918# a_31730_3918# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X511 a_21039_9161# a_20618_9161# a_20302_9271# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X512 gnd a_19167_3761# a_18959_3761# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X513 a_13851_9425# a_14108_9235# a_12916_8938# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X514 a_36857_7860# a_36644_7860# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X515 a_119_3546# a_648_3665# a_856_3665# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X516 a_30337_1096# a_30865_891# a_31073_891# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X517 a_15206_2489# a_15735_2608# a_15943_2608# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X518 a_1483_2842# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X519 a_1808_7373# a_1694_7254# a_1808_5173# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X520 gnd a_13170_6719# a_12962_6719# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X521 a_32009_6716# a_31588_6716# a_31071_6960# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X522 vdd a_18227_4554# a_18019_4554# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X523 a_35706_7001# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X524 a_1585_4524# a_1372_4524# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X525 a_36128_4795# a_35707_4795# a_35391_4676# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X526 a_2882_6904# a_3869_6470# a_3824_6483# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X527 a_29068_5956# a_29321_5943# a_28129_5646# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X528 a_26613_6752# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X529 a_18914_2671# a_18910_2848# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X530 a_37068_1242# a_36647_1242# a_36129_932# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X531 a_6848_7874# a_6427_7874# a_5909_7564# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X532 a_27052_2983# a_26755_3954# a_27036_3443# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X533 a_2746_6216# a_2999_6203# a_2772_7483# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X534 gnd a_33356_6700# a_33148_6700# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X535 vdd d0 a_24264_4245# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X536 a_23074_2296# a_23327_2283# a_22934_1785# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X537 a_39094_5584# a_39351_5394# a_38156_5828# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X538 a_30337_1326# a_30337_1096# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X539 a_25359_7106# a_25359_6877# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X540 vdd a_38304_5108# a_38096_5108# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X541 gnd d1 a_18228_2348# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X542 gnd d3 a_13060_7298# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X543 gnd d1 a_38411_8947# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X544 a_25886_8648# a_25673_8648# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X545 a_39100_2652# a_39353_2639# a_38161_2342# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X546 a_7944_3459# a_8928_3756# a_8883_3769# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X547 a_33102_8919# a_34086_9216# a_34041_9229# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X548 a_2744_1981# a_2934_1199# a_2885_1389# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X549 a_31072_3097# a_30651_3097# a_30336_2845# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X550 gnd a_39350_6497# a_39142_6497# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X551 a_11826_1220# a_11405_1220# a_10888_1464# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X552 a_6781_6179# a_6568_6179# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X553 a_8881_4318# a_9134_4305# a_7939_4739# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X554 a_30335_4635# a_30335_4405# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X555 a_26615_2340# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X556 a_20617_8607# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X557 a_7800_2022# a_8057_1832# a_7830_3112# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X558 a_11756_6143# a_11543_6143# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X559 a_35918_9207# a_35705_9207# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X560 a_35391_6195# a_35918_6447# a_36126_6447# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X561 a_26097_2030# a_25676_2030# a_25361_2235# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X562 gnd a_24262_8657# a_24054_8657# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X563 vdd a_34294_7559# a_34086_7559# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X564 a_1512_6138# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X565 a_39094_7241# a_39097_6510# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X566 a_36967_5081# a_36754_5081# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X567 a_26825_8958# a_26612_8958# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X568 vdd a_19167_3761# a_18959_3761# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X569 gnd a_13173_1204# a_12965_1204# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X570 a_7834_5135# a_7877_7334# a_7828_7524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X571 a_35920_4795# a_35707_4795# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X572 gnd d3 a_13062_2886# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X573 a_30333_9276# a_30862_9166# a_31070_9166# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X574 vdd d0 a_14109_7029# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X575 a_36128_5898# a_35707_5898# a_35391_6008# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X576 a_2745_8422# a_2930_8920# a_2881_9110# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X577 a_10466_3670# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X578 a_11512_7259# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X579 a_39099_5961# a_39095_6138# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X580 a_38015_6420# a_38205_5638# a_38156_5828# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X581 a_31698_5040# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X582 gnd a_34296_4804# a_34088_4804# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X583 a_5701_6461# a_5488_6461# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X584 a_25888_4236# a_25675_4236# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X585 gnd a_28383_3427# a_28175_3427# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X586 a_15940_7569# a_15519_7569# a_15204_7774# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X587 a_30335_4635# a_30864_4754# a_31072_4754# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X588 a_24014_1503# a_24267_1490# a_23075_1193# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X589 gnd a_3029_7293# a_2821_7293# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X590 gnd d0 a_34295_5353# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X591 gnd d0 a_29320_4286# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X592 vdd d2 a_28243_1813# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X593 a_17861_5317# a_18118_5127# a_17091_392# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X594 gnd d0 a_19168_1555# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X595 a_23070_2473# a_23327_2283# a_22934_1785# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X596 a_22931_8403# a_23116_8901# a_23067_9091# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X597 a_20619_4195# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X598 a_35919_8104# a_35706_8104# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X599 a_5490_4809# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X600 a_15205_5568# a_15205_5111# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X601 a_9779_210# a_9566_210# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X602 a_35393_1783# a_35920_2035# a_36128_2035# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X603 a_853_7523# a_1584_7833# a_1792_7833# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X604 gnd a_8195_7858# a_7987_7858# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X605 gnd a_24264_4245# a_24056_4245# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X606 a_26725_2864# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X607 vdd a_34296_3147# a_34088_3147# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X608 gnd d0 a_39351_8154# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X609 a_26826_7855# a_26613_7855# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X610 a_855_4768# a_1585_4524# a_1793_4524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X611 a_25361_3797# a_25890_3687# a_26098_3687# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X612 a_6640_6771# a_6427_6771# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X613 a_26827_4546# a_26614_4546# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X614 a_30334_7944# a_30863_8063# a_31071_8063# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X615 a_36955_373# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X616 a_7830_5312# a_7879_2922# a_7830_3112# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X617 a_12916_8938# a_13169_8925# a_12776_8427# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X618 a_38158_8960# a_39142_9257# a_39093_9447# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X619 gnd d1 a_33357_4494# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X620 a_38017_2008# a_38207_1226# a_38158_1416# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X621 a_5489_8118# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X622 a_118_5522# a_646_5317# a_854_5317# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X623 a_13851_7768# a_14108_7578# a_12913_8012# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X624 vdd a_2999_6203# a_2791_6203# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X625 a_13857_5939# a_13853_6116# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X626 a_646_8077# a_433_8077# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X627 a_15942_3157# a_15521_3157# a_15206_3362# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X628 gnd d0 a_34297_941# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X629 gnd a_3031_2881# a_2823_2881# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X630 a_34037_7749# a_34042_7023# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X631 a_3822_5008# a_4079_4818# a_2887_4521# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X632 a_35391_4446# a_35392_3989# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X633 a_5491_3706# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X634 a_37277_373# a_38096_5108# a_38051_5121# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X635 a_2881_9110# a_3868_8676# a_3819_8866# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X636 a_7834_5135# a_7877_7334# a_7832_7347# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X637 a_855_3111# a_1586_3421# a_1794_3421# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X638 a_31730_3918# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X639 a_32025_5159# a_31698_7240# a_32025_7359# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X640 a_26828_3443# a_26615_3443# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X641 a_6859_7295# a_6750_7295# a_6864_5214# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X642 a_24818_307# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X643 a_1372_4524# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X644 a_38160_4548# a_39144_4845# a_39095_5035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X645 a_21559_2299# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X646 vdd d0 a_29320_4286# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X647 vdd d0 a_34295_5353# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X648 a_32221_332# a_33040_5067# a_32991_5257# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X649 a_7799_4228# a_7989_3446# a_7940_3636# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X650 vdd d0 a_19168_1555# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X651 a_3826_2071# a_4079_2058# a_2884_2492# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X652 a_36127_5344# a_35706_5344# a_35391_5092# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X653 vdd d0 a_24265_4799# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X654 a_26936_5076# a_26723_5076# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X655 vdd d0 a_39351_8154# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X656 vdd a_24264_4245# a_24056_4245# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X657 a_33099_7993# a_34086_7559# a_34041_7572# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X658 a_13856_7042# a_14109_7029# a_12917_6732# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X659 a_22927_8580# a_23184_8390# a_22962_7287# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X660 gnd d0 a_34297_2598# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X661 gnd a_3141_3405# a_2933_3405# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X662 gnd a_18228_2348# a_18020_2348# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X663 a_30074_191# a_34849_312# a_35171_312# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X664 a_35918_7550# a_35705_7550# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X665 a_32963_6202# a_33216_6189# a_32989_7469# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X666 a_5175_3816# a_5175_3587# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X667 a_25673_8648# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X668 a_117_7271# a_117_7084# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X669 a_38017_2008# a_38207_1226# a_38162_1239# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X670 a_33104_4507# a_34088_4804# a_34039_4994# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X671 a_6861_2883# a_6752_2883# a_6859_5095# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X672 a_31073_3651# a_30652_3651# a_30336_3532# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X673 a_5173_6666# a_5174_6209# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X674 gnd d0 a_24265_2039# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X675 a_10676_9185# a_10463_9185# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X676 a_34040_2788# a_34043_2057# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X677 a_26098_2584# a_25677_2584# a_25361_2694# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X678 a_35705_9207# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X679 a_2886_7830# a_3870_8127# a_3825_8140# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X680 a_1584_6730# a_1371_6730# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X681 a_15203_9336# a_15203_9107# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X682 a_2881_9110# a_3868_8676# a_3823_8689# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X683 a_10148_8379# a_10148_8192# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X684 gnd d2 a_13032_1796# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X685 a_29067_8162# a_29320_8149# a_28128_7852# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X686 a_36754_5081# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X687 a_33101_3581# a_34088_3147# a_34043_3160# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X688 a_26612_8958# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X689 a_37067_3448# a_36646_3448# a_36128_3138# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X690 gnd a_13062_2886# a_12854_2886# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X691 a_6850_3462# a_6782_3973# a_6866_3002# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X692 a_2745_8422# a_2998_8409# a_2776_7306# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X693 a_16568_7300# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X694 a_118_5065# a_118_4878# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X695 a_23073_4502# a_23326_4489# a_22933_3991# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X696 a_28123_9132# a_29110_8698# a_29065_8711# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X697 a_24007_5538# a_24012_4812# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X698 a_5705_1500# a_5492_1500# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X699 a_25675_4236# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X700 a_7799_4228# a_7989_3446# a_7944_3459# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X701 a_25361_2235# a_25362_1778# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X702 a_15942_4814# a_15521_4814# a_15205_4695# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X703 gnd a_34295_5353# a_34087_5353# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X704 vdd a_28243_1813# a_28035_1813# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X705 a_32025_7359# a_31728_8330# a_32009_7819# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X706 a_38155_8034# a_39142_7600# a_39093_7790# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X707 a_37076_5081# a_36967_5081# a_37175_5081# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X708 gnd a_19168_1555# a_18960_1555# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X709 a_27987_8444# a_28240_8431# a_28018_7328# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X710 a_36858_5654# a_36645_5654# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X711 a_15943_951# a_15522_951# a_15209_1057# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X712 a_35706_8104# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X713 a_35390_6882# a_35390_6652# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X714 a_120_1340# a_649_1459# a_857_1459# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X715 a_15522_951# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X716 a_36129_2589# a_35708_2589# a_35392_2470# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X717 a_1586_2318# a_1373_2318# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X718 a_17972_8979# a_18225_8966# a_17832_8468# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X719 a_36856_8963# a_36643_8963# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X720 gnd d0 a_14110_4823# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X721 a_5704_946# a_5491_946# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X722 a_21770_7814# a_21557_7814# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X723 a_26613_7855# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X724 a_24005_8847# a_24011_8121# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X725 a_31589_5613# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X726 a_26614_4546# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X727 a_11755_8349# a_11542_8349# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X728 a_6849_5668# a_6428_5668# a_5910_5358# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X729 a_3822_5008# a_3825_4277# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X730 a_27047_2864# a_26756_1748# a_27037_1237# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X731 a_31587_8922# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X732 a_8878_5049# a_9135_4859# a_7943_4562# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X733 gnd a_33357_4494# a_33149_4494# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X734 a_27144_5076# a_27137_368# a_25140_307# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X735 a_2888_2315# a_3141_2302# a_2748_1804# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X736 a_1808_5173# a_1481_7254# a_1803_7254# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X737 gnd a_3001_1791# a_2793_1791# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X738 a_15943_3711# a_15522_3711# a_15206_3821# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X739 a_6847_8977# a_6426_8977# a_5909_9221# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X740 a_433_8077# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X741 a_5909_6461# a_6640_6771# a_6848_6771# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X742 a_25361_3797# a_25361_3568# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X743 gnd a_34297_941# a_34089_941# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X744 a_20832_6955# a_20619_6955# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X745 a_5700_8667# a_5487_8667# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X746 a_20303_6606# a_20304_6149# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X747 a_26968_3954# a_26755_3954# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X748 a_30339_997# a_30865_891# a_31073_891# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X749 a_15518_8672# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X750 a_24013_3709# a_24266_3696# a_23074_3399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X751 a_10675_8631# a_10462_8631# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X752 gnd d0 a_34294_7559# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X753 a_26615_3443# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X754 a_21772_3402# a_21559_3402# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X755 a_8882_2112# a_9135_2099# a_7940_2533# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X756 a_17861_5317# a_17910_2927# a_17865_2940# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X757 a_21699_3913# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X758 a_13856_5385# a_14109_5372# a_12914_5806# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X759 gnd d1 a_3138_8920# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X760 vdd d0 a_34296_5907# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X761 vdd d0 a_29321_4840# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X762 a_37067_2345# a_37000_1753# a_37078_2869# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X763 a_10151_1345# a_10151_1115# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X764 vdd a_34295_5353# a_34087_5353# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X765 a_5172_9102# a_5172_8872# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X766 a_20304_4400# a_20832_4195# a_21040_4195# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X767 a_31074_1445# a_31804_1201# a_32012_1201# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X768 vdd a_19168_1555# a_18960_1555# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X769 a_18912_8186# a_19165_8173# a_17973_7876# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X770 a_27983_8621# a_28240_8431# a_28018_7328# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X771 a_22190_327# a_23009_5062# a_22960_5252# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X772 a_30864_3097# a_30651_3097# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X773 vdd a_24265_4799# a_24057_4799# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X774 a_35921_2589# a_35708_2589# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X775 a_20833_5852# a_20620_5852# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X776 a_26723_5076# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X777 a_7939_4739# a_8926_4305# a_8877_4495# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X778 a_11836_2847# a_11727_2847# a_11834_5059# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X779 a_21880_5035# a_21667_5035# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X780 a_7830_3112# a_7849_1832# a_7804_1845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X781 a_5174_4919# a_5703_4809# a_5911_4809# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X782 gnd a_34297_2598# a_34089_2598# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X783 a_20834_2543# a_20621_2543# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X784 a_5702_4255# a_5489_4255# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X785 a_13858_973# a_13854_1150# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X786 a_25889_2030# a_25676_2030# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X787 a_8879_8730# a_8875_8907# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X788 a_30336_2429# a_30865_2548# a_31073_2548# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X789 a_35705_7550# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X790 gnd d0 a_34296_3147# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X791 vdd a_18088_1837# a_17880_1837# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X792 a_25360_4671# a_25360_4441# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X793 a_15733_7020# a_15520_7020# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X794 a_854_5317# a_1585_5627# a_1793_5627# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X795 gnd a_24265_2039# a_24057_2039# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X796 a_6640_7874# a_6427_7874# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X797 gnd d0 a_39352_5948# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X798 a_26827_5649# a_26614_5649# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X799 a_856_2562# a_1586_2318# a_1794_2318# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X800 a_16458_6776# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X801 a_33100_5787# a_34087_5353# a_34038_5543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X802 a_10463_9185# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X803 a_23068_7988# a_23325_7798# a_22927_8580# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X804 a_21880_7235# a_21667_7235# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X805 a_6641_4565# a_6428_4565# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X806 a_27985_4209# a_28242_4019# a_28020_2916# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X807 a_1371_6730# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X808 gnd a_13032_1796# a_12824_1796# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X809 gnd d1 a_33358_2288# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X810 a_13852_5562# a_14109_5372# a_12914_5806# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X811 a_17830_4233# a_18020_3451# a_17971_3641# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X812 a_21042_2543# a_21772_2299# a_21980_2299# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X813 a_37081_7400# a_36784_8371# a_37065_7860# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X814 a_21040_4195# a_20619_4195# a_20304_4400# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X815 a_25358_9312# a_25887_9202# a_26095_9202# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X816 gnd d2 a_23184_8390# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X817 gnd d2 a_38272_6230# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X818 a_5492_1500# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X819 a_18908_8363# a_19165_8173# a_17973_7876# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X820 a_29062_7785# a_29319_7595# a_28124_8029# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X821 a_2887_5624# a_3871_5921# a_3822_6111# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X822 a_22190_327# a_23009_5062# a_22964_5075# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X823 a_15206_4008# a_15206_3821# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X824 a_15207_1156# a_15209_1057# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X825 a_856_905# a_1587_1215# a_1795_1215# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X826 a_26829_1237# a_26616_1237# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X827 a_38018_8449# a_38203_8947# a_38158_8960# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X828 a_6642_3462# a_6429_3462# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X829 a_22929_4168# a_23186_3978# a_22964_2875# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X830 a_33102_1375# a_34089_941# a_34040_1131# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X831 a_1726_3932# a_1513_3932# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X832 a_21042_886# a_20621_886# a_20308_992# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X833 gnd d1 a_13169_8925# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X834 a_30334_7944# a_30334_7714# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X835 a_31072_5857# a_30651_5857# a_30335_5738# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X836 a_20621_886# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X837 a_20302_9042# a_20302_8812# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X838 a_28128_7852# a_28381_7839# a_27983_8621# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X839 a_1373_2318# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X840 a_5910_8118# a_5489_8118# a_5173_7999# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X841 a_23073_5605# a_24057_5902# a_24008_6092# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X842 a_31070_9166# a_30649_9166# a_30333_9276# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X843 a_852_8626# a_431_8626# a_116_8831# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X844 a_26097_4790# a_25676_4790# a_25360_4900# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X845 a_36128_3138# a_35707_3138# a_35392_2886# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X846 vdd d0 a_24266_2593# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X847 a_7937_9151# a_8194_8961# a_7801_8463# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X848 a_15205_4465# a_15206_4008# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X849 a_6864_5214# a_6537_7295# a_6864_7414# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X850 a_10678_4773# a_10465_4773# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X851 a_33100_5787# a_34087_5353# a_34042_5366# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X852 a_26096_8099# a_25675_8099# a_25359_7980# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X853 a_35707_4795# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X854 a_30336_2199# a_30864_1994# a_31072_1994# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X855 a_24009_8670# a_24005_8847# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X856 vdd a_39350_7600# a_39142_7600# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X857 a_32991_5257# a_33248_5067# a_32221_332# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X858 a_8877_5598# a_9134_5408# a_7939_5842# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X859 a_6849_5668# a_6781_6179# a_6859_7295# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X860 a_35919_5344# a_35706_5344# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X861 a_26755_3954# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X862 a_21980_2299# a_21559_2299# a_21042_2543# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X863 gnd d0 a_19166_2104# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X864 a_33105_2301# a_34089_2598# a_34040_2788# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X865 vdd d0 a_4078_8127# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X866 a_31074_1445# a_30653_1445# a_30337_1326# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X867 a_17830_4233# a_18020_3451# a_17975_3464# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X868 gnd d1 a_8194_8961# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X869 a_10462_8631# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X870 a_20831_7504# a_20618_7504# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X871 a_22962_7287# a_22976_8390# a_22931_8403# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X872 gnd a_34294_7559# a_34086_7559# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X873 a_8883_2666# a_9136_2653# a_7944_2356# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X874 a_34037_6646# a_34043_5920# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X875 vdd d2 a_38272_6230# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X876 a_854_4214# a_433_4214# a_118_4419# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X877 a_35391_4676# a_35920_4795# a_36128_4795# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X878 a_11826_1220# a_11758_1731# a_11836_2847# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X879 gnd a_3138_8920# a_2930_8920# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X880 vdd a_34296_5907# a_34088_5907# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X881 a_7939_4739# a_8196_4549# a_7803_4051# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X882 a_29065_1167# a_25364_1033# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X883 gnd d0 a_14109_7029# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X884 a_5174_6209# a_5701_6461# a_5909_6461# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X885 a_25890_2584# a_25677_2584# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X886 a_30865_3651# a_30652_3651# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X887 a_31588_7819# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X888 vdd d0 a_29320_5389# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X889 a_30651_3097# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X890 a_20620_5852# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X891 a_35708_932# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X892 a_17865_5140# a_18118_5127# a_17091_392# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X893 a_2887_4521# a_3140_4508# a_2747_4010# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X894 a_20621_2543# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X895 a_28124_6926# a_29111_6492# a_29066_6505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X896 a_12778_4015# a_13031_4002# a_12809_2899# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X897 a_25676_2030# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X898 vdd a_29320_8149# a_29112_8149# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X899 a_35390_7755# a_35390_7298# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X900 gnd d0 a_29322_2634# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X901 a_15943_2608# a_15522_2608# a_15206_2489# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X902 gnd a_34296_3147# a_34088_3147# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X903 a_38156_5828# a_39143_5394# a_39094_5584# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X904 a_27988_6238# a_28241_6225# a_28014_7505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X905 a_36859_3448# a_36646_3448# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X906 a_35707_5898# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X907 vdd d1 a_33357_5597# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X908 a_30336_2845# a_30864_3097# a_31072_3097# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X909 a_15520_7020# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X910 a_11823_6735# a_11402_6735# a_10885_6979# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X911 gnd a_39352_5948# a_39144_5948# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X912 a_21771_5608# a_21558_5608# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X913 a_26614_5649# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X914 a_15206_3592# a_15206_3362# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X915 a_5175_2713# a_5175_2484# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X916 a_32963_6202# a_33148_6700# a_33103_6713# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X917 a_11713_351# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X918 a_13855_7591# a_14108_7578# a_12913_8012# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X919 a_14985_331# a_14876_331# a_9888_210# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X920 a_3819_8866# a_3825_8140# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X921 a_31069_8612# a_30648_8612# a_30333_8817# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X922 a_1895_346# a_1682_346# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X923 a_37066_4551# a_36999_3959# a_37083_2988# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X924 a_39093_6687# a_39350_6497# a_38155_6931# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X925 gnd a_33358_2288# a_33150_2288# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X926 a_8879_2843# a_9136_2653# a_7944_2356# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X927 a_5053_326# a_4632_326# a_2103_346# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X928 a_15944_1505# a_15523_1505# a_15207_1615# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X929 a_5910_4255# a_6641_4565# a_6849_4565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X930 a_18913_3220# a_18909_3397# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X931 a_15204_6901# a_15204_6671# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X932 a_38158_1416# a_39145_982# a_39096_1172# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X933 vdd d3 a_18118_2927# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X934 a_10148_7276# a_10148_7089# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X935 gnd a_38272_6230# a_38064_6230# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X936 a_20833_4749# a_20620_4749# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X937 a_25140_307# a_26924_368# a_27246_368# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X938 vdd d0 a_4080_955# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X939 a_27990_1826# a_28243_1813# a_28016_3093# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X940 a_6782_3973# a_6569_3973# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X941 a_26969_1748# a_26756_1748# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X942 a_7943_4562# a_8927_4859# a_8882_4872# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X943 a_2748_1804# a_2933_2302# a_2884_2492# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X944 a_15519_6466# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X945 a_11825_2323# a_11404_2323# a_10887_2567# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X946 a_10676_6425# a_10463_6425# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X947 a_32010_5613# a_31589_5613# a_31071_5303# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X948 a_26616_1237# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X949 a_1513_3932# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X950 a_24007_4435# a_24013_3709# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X951 a_34039_6097# a_34042_5366# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X952 vdd d0 a_29322_2634# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X953 a_16890_5100# a_16570_2888# a_16897_3007# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X954 vdd d0 a_34297_3701# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X955 a_15732_9226# a_15519_9226# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X956 a_33099_7993# a_34086_7559# a_34037_7749# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X957 a_27984_6415# a_28241_6225# a_28014_7505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X958 a_8880_7627# a_9133_7614# a_7938_8048# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X959 a_31698_7240# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X960 a_18913_5980# a_19166_5967# a_17974_5670# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X961 vdd a_24266_2593# a_24058_2593# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X962 a_36127_7001# a_35706_7001# a_35390_7111# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X963 a_7940_2533# a_8927_2099# a_8878_2289# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X964 a_28020_2916# a_28273_2903# a_28016_5293# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X965 a_24010_9224# a_24263_9211# a_23071_8914# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X966 a_33104_5610# a_34088_5907# a_34043_5920# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X967 a_10465_4773# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X968 a_20834_3646# a_20621_3646# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X969 a_22934_1785# a_23187_1772# a_22960_3052# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X970 a_10147_9295# a_10676_9185# a_10884_9185# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X971 a_38019_6243# a_38204_6741# a_38155_6931# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X972 gnd a_28382_4530# a_28174_4530# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X973 a_5703_2049# a_5490_2049# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X974 vdd d0 a_9134_8168# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X975 a_10677_5322# a_10464_5322# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X976 a_25360_5544# a_25360_5087# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X977 a_25031_307# a_24818_307# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X978 a_5053_326# a_9779_210# a_9987_210# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X979 a_35706_5344# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X980 a_32012_1201# a_31591_1201# a_31073_891# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X981 a_10678_2013# a_10465_2013# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X982 a_17973_7876# a_18957_8173# a_18908_8363# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X983 gnd d0 a_14109_5372# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X984 a_33102_8919# a_33355_8906# a_32962_8408# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X985 gnd d2 a_38271_8436# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X986 a_16897_3007# a_16600_3978# a_16880_4570# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X987 gnd a_19166_2104# a_18958_2104# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X988 vdd a_4078_8127# a_3870_8127# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X989 a_11834_5059# a_11514_2847# a_11841_2966# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X990 a_2886_7830# a_3870_8127# a_3821_8317# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X991 a_15733_8123# a_15520_8123# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X992 a_7942_6768# a_8195_6755# a_7802_6257# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X993 gnd a_8194_8961# a_7986_8961# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X994 a_25360_4900# a_25889_4790# a_26097_4790# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X995 a_6641_5668# a_6428_5668# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X996 a_25361_2694# a_25361_2465# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X997 vdd a_38272_6230# a_38064_6230# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X998 a_16459_4570# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X999 a_33101_3581# a_34088_3147# a_34039_3337# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1000 a_6642_2359# a_6429_2359# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1001 a_11616_5632# a_11403_5632# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1002 a_23069_5782# a_23326_5592# a_22928_6374# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1003 a_647_5871# a_434_5871# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1004 a_5488_9221# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1005 a_3821_8317# a_3824_7586# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1006 a_23072_7811# a_24056_8108# a_24007_8298# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1007 a_30334_8173# a_30334_7944# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1008 a_117_6625# a_645_6420# a_853_6420# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1009 a_8884_1563# a_8880_1740# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1010 a_30652_3651# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1011 a_20302_9271# a_20302_9042# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1012 a_11614_8941# a_11401_8941# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1013 a_34041_6469# a_34037_6646# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1014 a_17831_2027# a_18021_1245# a_17972_1435# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1015 a_8881_4318# a_8877_4495# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1016 a_37076_7281# a_36785_6165# a_37066_5654# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1017 a_21041_1989# a_20620_1989# a_20305_2194# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1018 a_25677_2584# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1019 gnd d2 a_23185_6184# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1020 a_119_3546# a_119_3316# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1021 gnd d2 a_38273_4024# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1022 gnd d0 a_14111_960# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1023 vdd d1 a_38413_5638# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1024 a_25362_1132# a_25890_927# a_26098_927# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1025 gnd a_29322_2634# a_29114_2634# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1026 a_7944_2356# a_8197_2343# a_7804_1845# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1027 a_8876_7804# a_9133_7614# a_7938_8048# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1028 a_21040_8058# a_21770_7814# a_21978_7814# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1029 a_24006_9401# a_24263_9211# a_23071_8914# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1030 a_24006_9401# a_24009_8670# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1031 a_18912_7083# a_18908_7260# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1032 a_22930_1962# a_23187_1772# a_22960_3052# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1033 a_6643_1256# a_6430_1256# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1034 a_38019_6243# a_38204_6741# a_38159_6754# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1035 vdd a_33357_5597# a_33149_5597# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1036 vdd a_28382_4530# a_28174_4530# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1037 a_11618_1220# a_11405_1220# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1038 a_1727_1726# a_1514_1726# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1039 a_36997_8371# a_36784_8371# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1040 a_24009_3886# a_24012_3155# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1041 a_30649_7509# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1042 a_17973_7876# a_18957_8173# a_18912_8186# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1043 a_20303_7065# a_20303_6836# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1044 a_31071_6960# a_30650_6960# a_30334_7070# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1045 vdd d0 a_14109_5372# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1046 vdd d0 a_19167_2658# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1047 vdd d2 a_38271_8436# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1048 a_18911_7632# a_18907_7809# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1049 a_853_6420# a_432_6420# a_117_6625# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1050 gnd a_29321_5943# a_29113_5943# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1051 a_31728_8330# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1052 a_22964_2875# a_22978_3978# a_22933_3991# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1053 a_7938_6945# a_8195_6755# a_7802_6257# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1054 vdd d0 a_39350_9257# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1055 a_20303_7065# a_20832_6955# a_21040_6955# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1056 a_17829_6439# a_18086_6249# a_17859_7529# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1057 a_25360_5774# a_25889_5893# a_26097_5893# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1058 gnd d4 a_8087_5122# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1059 a_10679_2567# a_10466_2567# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1060 a_27045_5076# a_26725_2864# a_27052_2983# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1061 a_5173_8415# a_5700_8667# a_5908_8667# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1062 a_30864_5857# a_30651_5857# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1063 a_35391_5092# a_35391_4905# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1064 a_3822_3351# a_3827_2625# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1065 vdd d0 a_29319_7595# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1066 a_35708_2589# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1067 vdd a_39351_5394# a_39143_5394# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1068 a_37064_8963# a_36643_8963# a_36125_8653# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1069 a_8878_3392# a_9135_3202# a_7940_3636# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1070 a_30862_9166# a_30649_9166# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1071 a_18913_4877# a_18909_5054# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1072 a_16881_2364# a_16460_2364# a_15943_2608# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1073 vdd a_18118_2927# a_17910_2927# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1074 a_21042_3646# a_21772_3402# a_21980_3402# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1075 a_3823_8689# a_3819_8866# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1076 a_20620_4749# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1077 a_25889_4790# a_25676_4790# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1078 a_7801_8463# a_7986_8961# a_7941_8974# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1079 a_12777_6221# a_13030_6208# a_12803_7488# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1080 a_38021_1831# a_38206_2329# a_38161_2342# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1081 a_6958_5095# a_6951_387# a_4954_326# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1082 a_26756_1748# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1083 a_17831_2027# a_18021_1245# a_17976_1258# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1084 a_10463_6425# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1085 a_28016_5293# a_28065_2903# a_28020_2916# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1086 a_2776_7306# a_2790_8409# a_2745_8422# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1087 a_25888_8099# a_25675_8099# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1088 a_25359_7980# a_25359_7750# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1089 vdd d2 a_23185_6184# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1090 a_7939_5842# a_8926_5408# a_8881_5421# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1091 vdd d2 a_38273_4024# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1092 a_35392_2470# a_35921_2589# a_36129_2589# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1093 a_855_2008# a_434_2008# a_119_2213# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1094 vdd d1 a_33356_7803# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1095 a_6859_7295# a_6568_6179# a_6848_6771# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1096 a_20304_5733# a_20833_5852# a_21041_5852# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1097 a_21994_5154# a_21880_5035# a_22088_5035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1098 vdd a_29322_2634# a_29114_2634# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1099 a_7940_2533# a_8197_2343# a_7804_1845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1100 vdd a_34297_3701# a_34089_3701# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1101 a_38160_5651# a_39144_5948# a_39099_5961# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1102 a_32960_4173# a_33150_3391# a_33101_3581# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1103 a_20619_8058# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1104 a_5175_4003# a_5702_4255# a_5910_4255# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1105 a_15206_2905# a_15206_2718# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1106 a_32962_8408# a_33147_8906# a_33102_8919# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1107 a_30866_1445# a_30653_1445# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1108 a_7944_2356# a_8928_2653# a_8879_2843# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1109 gnd d3 a_38302_7320# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1110 a_24011_4258# a_24007_4435# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1111 a_37066_4551# a_36645_4551# a_36127_4241# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1112 a_20621_3646# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1113 a_6750_5095# a_6537_5095# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1114 a_856_905# a_435_905# a_122_1011# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1115 a_11836_2847# a_11545_1731# a_11825_2323# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1116 a_5704_2603# a_5491_2603# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1117 a_7803_4051# a_7988_4549# a_7943_4562# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1118 a_5490_2049# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1119 vdd a_9134_8168# a_8926_8168# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1120 a_10464_5322# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1121 a_15204_7130# a_15733_7020# a_15941_7020# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1122 a_5909_6461# a_5488_6461# a_5173_6666# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1123 a_31899_332# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1124 a_2778_2894# a_2792_3997# a_2747_4010# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1125 a_35171_312# a_35062_312# a_30074_191# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1126 a_10465_2013# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1127 a_21989_7235# a_21880_7235# a_21994_5154# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1128 vdd d4 a_8087_5122# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1129 a_38157_3622# a_39144_3188# a_39095_3378# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1130 a_27989_4032# a_28242_4019# a_28020_2916# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1131 a_17091_392# a_16982_392# a_14985_331# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1132 a_119_2443# a_648_2562# a_856_2562# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1133 vdd d1 a_33358_3391# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1134 a_15520_8123# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1135 a_16672_5673# a_16459_5673# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1136 a_2747_4010# a_2932_4508# a_2883_4698# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1137 a_39098_8167# a_39094_8344# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1138 a_29068_4853# a_29321_4840# a_28129_4543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1139 a_11824_4529# a_11403_4529# a_10886_4773# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1140 a_12809_2899# a_12823_4002# a_12774_4192# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1141 a_4954_326# a_6738_387# a_6958_5095# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1142 a_11933_5059# a_11926_351# a_12134_351# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1143 a_32964_3996# a_33149_4494# a_33104_4507# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1144 vdd a_34297_941# a_34089_941# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1145 gnd d0 a_9135_5962# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1146 a_2103_346# a_1682_346# a_2004_346# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1147 a_11403_5632# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1148 a_6848_6771# a_6427_6771# a_5909_6461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1149 a_434_5871# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1150 a_11401_8941# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1151 a_15204_7774# a_15204_7317# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1152 a_24012_5915# a_24008_6092# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1153 a_39094_4481# a_39351_4291# a_38156_4725# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1154 a_25361_2881# a_25361_2694# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1155 gnd a_4079_5921# a_3871_5921# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1156 a_31944_1712# a_31731_1712# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1157 a_5911_2049# a_6642_2359# a_6850_2359# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1158 a_36126_9207# a_35705_9207# a_35389_9317# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1159 vdd d0 a_19164_7619# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1160 a_30334_8360# a_30334_8173# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1161 gnd a_38273_4024# a_38065_4024# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1162 a_2887_5624# a_3140_5611# a_2742_6393# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1163 vdd a_38413_5638# a_38205_5638# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1164 a_6783_1767# a_6570_1767# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1165 a_16674_1261# a_16461_1261# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1166 a_7944_2356# a_8928_2653# a_8883_2666# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1167 gnd d0 a_34293_8662# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1168 a_10676_7528# a_10463_7528# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1169 vdd d3 a_38302_7320# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1170 a_3828_1522# a_4081_1509# a_2889_1212# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1171 a_10677_4219# a_10464_4219# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1172 a_32011_3407# a_31590_3407# a_31072_3097# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1173 a_29062_9442# a_29065_8711# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1174 a_6430_1256# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1175 a_1514_1726# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1176 a_11405_1220# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1177 a_36784_8371# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1178 vdd d0 a_34298_1495# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1179 a_17832_8468# a_18085_8455# a_17863_7352# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1180 a_25359_7106# a_25888_6996# a_26096_6996# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1181 a_16881_2364# a_16814_1772# a_16892_2888# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1182 vdd a_19167_2658# a_18959_2658# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1183 gnd d1 a_38414_3432# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1184 a_32995_5080# a_33248_5067# a_32221_332# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1185 a_11615_7838# a_11402_7838# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1186 a_5173_8228# a_5173_7999# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1187 vdd d0 a_19166_3207# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1188 a_20835_1440# a_20622_1440# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1189 a_21989_5035# a_21669_2823# a_21991_2823# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1190 a_10466_2567# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1191 a_33105_3404# a_34089_3701# a_34044_3714# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1192 a_116_8831# a_644_8626# a_852_8626# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1193 a_30651_5857# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1194 a_38020_4037# a_38205_4535# a_38156_4725# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1195 gnd a_28383_2324# a_28175_2324# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1196 a_20304_4400# a_20305_3943# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1197 a_15206_2489# a_15206_2259# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1198 gnd d0 a_4078_8127# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1199 a_20303_7709# a_20831_7504# a_21039_7504# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1200 a_15940_6466# a_15519_6466# a_15204_6671# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1201 a_10678_3116# a_10465_3116# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1202 a_29063_7236# a_29066_6505# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1203 gnd d0 a_34295_4250# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1204 a_17974_5670# a_18958_5967# a_18909_6157# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1205 a_25676_4790# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1206 a_35707_3138# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1207 a_7938_8048# a_8925_7614# a_8876_7804# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1208 gnd d0 a_14110_3166# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1209 vdd d1 a_38412_7844# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1210 a_35919_7001# a_35706_7001# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1211 a_7943_4562# a_8196_4549# a_7803_4051# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1212 a_22960_3052# a_22979_1772# a_22930_1962# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1213 a_10884_9185# a_10463_9185# a_10147_9066# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1214 a_39092_8893# a_39098_8167# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1215 gnd d0 a_39351_7051# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1216 a_15734_5917# a_15521_5917# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1217 a_27050_5195# a_26936_5076# a_27144_5076# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1218 a_17834_4056# a_18087_4043# a_17865_2940# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1219 a_25675_8099# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1220 a_26826_6752# a_26613_6752# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1221 a_29068_5956# a_29064_6133# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1222 a_17970_5847# a_18227_5657# a_17829_6439# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1223 a_18913_2117# a_18909_2294# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1224 a_25361_2694# a_25890_2584# a_26098_2584# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1225 vdd a_33356_7803# a_33148_7803# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1226 vdd a_38273_4024# a_38065_4024# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1227 a_120_1110# a_648_905# a_856_905# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1228 a_2883_5801# a_3140_5611# a_2742_6393# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1229 a_11617_3426# a_11404_3426# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1230 vref a_116_9290# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1231 vdd d0 a_34293_8662# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1232 a_117_7271# a_645_7523# a_853_7523# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1233 a_648_3665# a_435_3665# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1234 a_5489_7015# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1235 a_30653_1445# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1236 a_36125_8653# a_35704_8653# a_35390_8401# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1237 a_7802_6257# a_7987_6755# a_7938_6945# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1238 vdd d0 a_19166_4864# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1239 a_118_4419# a_646_4214# a_854_4214# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1240 gnd d1 a_13172_2307# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1241 gnd a_29320_8149# a_29112_8149# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1242 a_646_6974# a_433_6974# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1243 a_15942_2054# a_15521_2054# a_15206_2259# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1244 vdd d3 a_33248_2867# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1245 gnd a_38302_7320# a_38094_7320# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1246 a_32991_3057# a_33010_1777# a_32965_1790# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1247 a_17828_8645# a_18085_8455# a_17863_7352# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1248 a_34039_4994# a_34042_4263# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1249 a_18908_8363# a_18911_7632# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1250 a_25359_7980# a_25888_8099# a_26096_8099# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1251 a_5491_2603# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1252 a_2741_8599# a_2931_7817# a_2886_7830# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1253 a_27045_7276# a_26936_7276# a_27050_5195# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1254 gnd d2 a_2999_6203# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1255 gnd d2 a_23186_3978# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1256 gnd d2 a_38274_1818# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1257 vdd d1 a_38414_3432# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1258 a_29061_8888# a_29318_8698# a_28123_9132# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1259 a_11725_5059# a_11512_5059# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1260 a_38161_3445# a_39145_3742# a_39096_3932# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1261 a_21041_5852# a_21771_5608# a_21979_5608# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1262 a_16880_4570# a_16459_4570# a_15942_4814# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1263 a_13850_8871# a_13856_8145# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1264 a_24007_7195# a_24264_7005# a_23072_6708# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1265 a_22190_327# a_22081_327# a_22289_327# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1266 a_38020_4037# a_38205_4535# a_38160_4548# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1267 vdd a_28383_2324# a_28175_2324# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1268 a_21038_8607# a_21769_8917# a_21977_8917# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1269 a_31071_6960# a_30650_6960# a_30334_6841# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1270 a_2885_1389# a_3142_1199# a_2744_1981# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1271 vdd a_33358_3391# a_33150_3391# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1272 a_3820_9420# a_3823_8689# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1273 a_28127_8955# a_28380_8942# a_27987_8444# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1274 gnd a_28240_8431# a_28032_8431# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1275 a_36998_6165# a_36785_6165# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1276 vdd d0 a_34295_4250# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1277 a_34043_5920# a_34296_5907# a_33104_5610# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1278 a_119_2859# a_647_3111# a_855_3111# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1279 a_7938_8048# a_8925_7614# a_8880_7627# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1280 a_36127_4241# a_35706_4241# a_35392_3989# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1281 a_35921_932# a_35708_932# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1282 a_7804_1845# a_7989_2343# a_7940_2533# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1283 vdd d0 a_14110_3166# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1284 a_21910_8325# a_21697_8325# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1285 gnd a_9135_5962# a_8927_5962# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1286 a_21978_7814# a_21557_7814# a_21039_7504# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1287 a_31729_6124# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1288 a_37000_1753# a_36787_1753# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1289 a_22960_3052# a_22979_1772# a_22934_1785# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1290 a_11725_7259# a_11512_7259# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1291 vdd d0 a_39351_7051# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1292 a_20304_4859# a_20833_4749# a_21041_4749# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1293 a_17830_4233# a_18087_4043# a_17865_2940# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1294 a_35389_9088# a_35389_8858# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1295 a_6849_4565# a_6782_3973# a_6866_3002# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1296 a_18910_1191# a_15209_1057# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1297 a_10148_6630# a_10149_6173# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1298 a_31731_1712# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1299 gnd a_3141_2302# a_2933_2302# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1300 a_37065_6757# a_36644_6757# a_36126_6447# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1301 a_8879_1186# a_9136_996# a_7941_1430# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1302 a_15207_1802# a_15207_1615# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1303 vdd a_19164_7619# a_18956_7619# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1304 a_30863_6960# a_30650_6960# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1305 a_5703_4809# a_5490_4809# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1306 a_15733_5363# a_15520_5363# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1307 a_3821_7214# a_3824_6483# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1308 a_7802_6257# a_7987_6755# a_7942_6768# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1309 a_17859_7529# a_17878_6249# a_17833_6262# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1310 a_6570_1767# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1311 a_10463_7528# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1312 a_16461_1261# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1313 a_26938_2864# a_26725_2864# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1314 a_15203_9336# a_15732_9226# a_15940_9226# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1315 a_5908_8667# a_5487_8667# a_5172_8872# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1316 gnd a_34293_8662# a_34085_8662# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1317 vdd a_38302_7320# a_38094_7320# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1318 a_2772_7483# a_2791_6203# a_2746_6216# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1319 a_29062_6682# a_29068_5956# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1320 a_10464_4219# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1321 a_36856_8963# a_36643_8963# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1322 a_118_4649# a_647_4768# a_855_4768# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1323 a_7940_3636# a_8927_3202# a_8882_3215# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1324 a_38051_5121# a_38304_5108# a_37277_373# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1325 a_119_2443# a_119_2213# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1326 a_16671_7879# a_16458_7879# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1327 gnd d0 a_19165_5413# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1328 a_1808_5173# a_1694_5054# a_1902_5054# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1329 vdd a_34298_1495# a_34090_1495# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1330 a_39099_3201# a_39095_3378# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1331 a_29067_7059# a_29320_7046# a_28128_6749# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1332 a_12803_7488# a_12822_6208# a_12773_6398# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1333 a_32961_1967# a_33151_1185# a_33102_1375# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1334 a_38161_3445# a_39145_3742# a_39100_3755# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1335 a_35393_1137# a_35395_1038# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1336 a_31587_8922# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1337 a_5176_1797# a_5703_2049# a_5911_2049# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1338 gnd a_38414_3432# a_38206_3432# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1339 gnd d0 a_9134_8168# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1340 a_37066_5654# a_36645_5654# a_36128_5898# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1341 a_11402_7838# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1342 a_25359_7750# a_25887_7545# a_26095_7545# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1343 a_37067_2345# a_36646_2345# a_36128_2035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1344 a_6847_8977# a_6426_8977# a_5908_8667# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1345 vdd a_28240_8431# a_28032_8431# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1346 vdd a_19166_3207# a_18958_3207# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1347 a_32119_5040# a_32112_332# a_32320_332# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1348 a_20622_1440# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1349 a_24009_2783# a_24012_2052# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1350 a_8880_7627# a_8876_7804# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1351 a_7804_1845# a_7989_2343# a_7944_2356# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1352 gnd a_4078_8127# a_3870_8127# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1353 a_15204_8004# a_15733_8123# a_15941_8123# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1354 a_22960_3052# a_23217_2862# a_22960_5252# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1355 gnd a_34295_4250# a_34087_4250# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1356 a_10465_3116# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1357 a_38051_5121# a_38094_7320# a_38045_7510# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1358 gnd d0 a_14111_3720# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1359 a_1803_7254# a_1694_7254# a_1808_5173# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1360 a_648_905# a_435_905# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1361 a_35706_7001# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1362 a_3826_4831# a_3822_5008# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1363 a_36858_4551# a_36645_4551# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1364 a_3822_2248# a_3828_1522# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1365 a_13852_8322# a_13855_7591# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1366 vdd a_38412_7844# a_38204_7844# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1367 a_21040_8058# a_20619_8058# a_20303_7939# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1368 a_15521_5917# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1369 a_16673_3467# a_16460_3467# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1370 gnd d2 a_8054_8450# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1371 a_21770_6711# a_21557_6711# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1372 a_26613_6752# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1373 a_4845_326# a_4632_326# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1374 a_31589_4510# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1375 a_13854_8694# a_14107_8681# a_12912_9115# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1376 a_17859_7529# a_18116_7339# a_17865_5140# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1377 a_37068_1242# a_36647_1242# a_36130_1486# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1378 a_6848_7874# a_6427_7874# a_5910_8118# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1379 a_11404_3426# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1380 a_25361_3338# a_25889_3133# a_26097_3133# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1381 a_6849_4565# a_6428_4565# a_5910_4255# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1382 vdd a_34293_8662# a_34085_8662# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1383 a_435_3665# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1384 vdd a_19166_4864# a_18958_4864# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1385 a_25359_6877# a_25359_6647# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1386 a_24007_5538# a_24264_5348# a_23069_5782# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1387 gnd d1 a_38413_5638# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1388 a_37076_5081# a_36756_2869# a_37078_2869# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1389 gnd a_13172_2307# a_12964_2307# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1390 a_433_6974# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1391 a_34040_1131# a_34297_941# a_33102_1375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1392 vdd a_33248_2867# a_33040_2867# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1393 a_5175_3357# a_5175_2900# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1394 vdd d0 a_19165_5413# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1395 a_17975_3464# a_18228_3451# a_17830_4233# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1396 a_29063_7236# a_29320_7046# a_28128_6749# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1397 a_32961_1967# a_33151_1185# a_33106_1198# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1398 gnd a_38274_1818# a_38066_1818# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1399 a_11512_5059# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1400 vdd a_38414_3432# a_38206_3432# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1401 gnd d1 a_23324_8901# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1402 a_24013_2606# a_24266_2593# a_23074_2296# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1403 a_20306_1550# a_20835_1440# a_21043_1440# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1404 gnd d0 a_34294_6456# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1405 a_14876_331# a_14663_331# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1406 gnd d0 a_19167_2658# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1407 a_35918_9207# a_35705_9207# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1408 a_11756_6143# a_11543_6143# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1409 a_36785_6165# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1410 gnd d0 a_39350_9257# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1411 a_17833_6262# a_18086_6249# a_17859_7529# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1412 vdd a_34295_4250# a_34087_4250# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1413 a_120_1756# a_120_1569# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1414 a_33098_9096# a_34085_8662# a_34036_8852# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1415 a_17969_8053# a_18226_7863# a_17828_8645# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1416 a_38051_5121# a_38094_7320# a_38049_7333# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1417 a_2742_6393# a_2932_5611# a_2883_5801# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1418 vdd d0 a_14111_3720# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1419 gnd a_28381_7839# a_28173_7839# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1420 a_18912_7083# a_19165_7070# a_17973_6773# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1421 gnd d1 a_38415_1226# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1422 a_2889_1212# a_3873_1509# a_3824_1699# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1423 a_30333_9047# a_30862_9166# a_31070_9166# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1424 vdd d2 a_8054_8450# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1425 a_11512_7259# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1426 vdd d0 a_19167_1001# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1427 a_24010_7567# a_24006_7744# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1428 a_854_8077# a_433_8077# a_117_7958# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1429 a_38021_1831# a_38206_2329# a_38157_2519# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1430 a_645_9180# a_432_9180# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1431 a_13850_8871# a_14107_8681# a_12912_9115# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1432 a_17863_7352# a_17877_8455# a_17828_8645# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1433 a_22928_6374# a_23118_5592# a_23069_5782# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1434 a_15941_4260# a_15520_4260# a_15205_4465# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1435 a_16892_2888# a_16601_1772# a_16882_1261# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1436 a_10679_910# a_10466_910# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1437 a_30650_6960# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1438 gnd d0 a_34296_2044# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1439 a_5490_4809# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1440 a_15520_5363# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1441 a_24012_4812# a_24008_4989# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1442 a_9987_210# a_9566_210# a_9888_210# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1443 a_9566_210# d7 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1444 a_3824_1699# a_3827_968# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1445 a_2774_3071# a_2793_1791# a_2744_1981# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1446 a_21882_2823# a_21669_2823# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1447 a_26725_2864# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1448 a_854_4214# a_1585_4524# a_1793_4524# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1449 gnd d0 a_39352_4845# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1450 a_17835_1850# a_18088_1837# a_17861_3117# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1451 a_6640_6771# a_6427_6771# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1452 a_26827_4546# a_26614_4546# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1453 a_33100_4684# a_34087_4250# a_34038_4440# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1454 a_17971_3641# a_18228_3451# a_17830_4233# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1455 a_21039_7504# a_20618_7504# a_20303_7252# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1456 a_32119_5040# a_31698_5040# a_32025_5159# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1457 a_36955_373# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1458 a_30334_7257# a_30334_7070# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1459 a_2884_3595# a_3141_3405# a_2743_4187# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1460 a_6859_5095# a_6750_5095# a_6958_5095# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1461 gnd a_19165_5413# a_18957_5413# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1462 a_5489_8118# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1463 vdd d0 a_34294_6456# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1464 vdd d2 a_8056_4038# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1465 a_649_1459# a_436_1459# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1466 a_118_5065# a_646_5317# a_854_5317# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1467 a_36126_6447# a_35705_6447# a_35391_6195# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1468 a_7803_4051# a_7988_4549# a_7939_4739# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1469 a_119_2213# a_647_2008# a_855_2008# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1470 gnd a_9134_8168# a_8926_8168# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1471 a_16781_7300# a_16568_7300# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1472 a_13852_4459# a_14109_4269# a_12914_4703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1473 a_17865_2940# a_17879_4043# a_17830_4233# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1474 a_32991_5257# a_33040_2867# a_32991_3057# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1475 a_33098_9096# a_34085_8662# a_34040_8675# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1476 a_2742_6393# a_2932_5611# a_2887_5624# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1477 gnd d2 a_3000_3997# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1478 a_15942_5917# a_16672_5673# a_16880_5673# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1479 vdd d1 a_38415_1226# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1480 a_8875_8907# a_9132_8717# a_7937_9151# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1481 a_18908_7260# a_19165_7070# a_17973_6773# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1482 a_29062_6682# a_29319_6492# a_28124_6926# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1483 gnd a_3140_4508# a_2932_4508# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1484 gnd a_13031_4002# a_12823_4002# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1485 a_35917_8653# a_35704_8653# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1486 a_5173_7125# a_5173_6896# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1487 a_38162_1239# a_39146_1536# a_39097_1726# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1488 a_24818_307# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1489 a_15732_7569# a_15519_7569# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1490 a_17863_7352# a_17877_8455# a_17832_8468# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1491 a_31072_4754# a_30651_4754# a_30335_4635# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1492 gnd a_8054_8450# a_7846_8450# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1493 gnd a_28241_6225# a_28033_6225# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1494 a_16460_3467# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1495 a_30648_8612# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1496 a_5910_7015# a_5489_7015# a_5173_6896# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1497 a_16811_8390# a_16598_8390# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1498 vdd d3 a_13060_7298# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1499 a_36127_5344# a_35706_5344# a_35391_5549# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1500 a_122_1011# a_648_905# a_856_905# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1501 vdd d0 a_34296_2044# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1502 a_24010_7567# a_24263_7554# a_23068_7988# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1503 a_21911_6119# a_21698_6119# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1504 a_36128_2035# a_35707_2035# a_35393_1783# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1505 a_1792_7833# a_1371_7833# a_853_7523# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1506 a_21979_5608# a_21558_5608# a_21040_5298# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1507 gnd d0 a_19164_7619# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1508 a_21977_8917# a_21556_8917# a_21039_9161# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1509 a_30863_6960# a_30650_6960# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1510 a_33100_4684# a_34087_4250# a_34042_4263# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1511 a_2744_1981# a_2934_1199# a_2889_1212# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1512 gnd a_38413_5638# a_38205_5638# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1513 a_6850_2359# a_6783_1767# a_6861_2883# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1514 a_37065_7860# a_36644_7860# a_36127_8104# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1515 vdd a_39350_6497# a_39142_6497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1516 a_25362_1362# a_25362_1132# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1517 a_30074_191# a_34849_312# a_32320_332# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1518 gnd d1 a_13172_3410# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1519 a_14985_331# a_16769_392# a_16989_5100# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1520 vdd a_19165_5413# a_18957_5413# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1521 a_35919_4241# a_35706_4241# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1522 gnd d0 a_39350_7600# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1523 a_15734_3157# a_15521_3157# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1524 a_31073_3651# a_30652_3651# a_30336_3761# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1525 gnd a_23324_8901# a_23116_8901# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1526 a_16568_5100# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1527 a_17835_1850# a_18020_2348# a_17975_2361# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1528 a_5911_5912# a_5490_5912# a_5174_6022# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1529 a_17865_2940# a_17879_4043# a_17834_4056# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1530 gnd a_34294_6456# a_34086_6456# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1531 a_20831_6401# a_20618_6401# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1532 a_38154_9137# a_39141_8703# a_39092_8893# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1533 a_28016_5293# a_28273_5103# a_27246_368# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1534 a_36129_932# a_35708_932# a_35393_1137# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1535 a_2744_1981# a_3001_1791# a_2774_3071# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1536 gnd a_19167_2658# a_18959_2658# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1537 a_35705_9207# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1538 a_36857_6757# a_36644_6757# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1539 a_18912_5426# a_18908_5603# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1540 a_7941_1430# a_8928_996# a_8883_1009# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1541 a_24012_3155# a_24265_3142# a_23070_3576# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1542 a_5488_7564# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1543 a_1794_3421# a_1373_3421# a_855_3111# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1544 vdd d1 a_13170_7822# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1545 a_20618_9161# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1546 a_38162_1239# a_39146_1536# a_39101_1549# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1547 a_31588_6716# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1548 gnd a_38415_1226# a_38207_1226# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1549 a_10680_1464# a_10467_1464# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1550 a_37067_3448# a_36646_3448# a_36129_3692# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1551 a_25360_5544# a_25888_5339# a_26096_5339# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1552 vdd a_8054_8450# a_7846_8450# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1553 vdd a_28241_6225# a_28033_6225# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1554 vdd a_19167_1001# a_18959_1001# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1555 a_34849_312# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1556 a_34038_8303# a_34041_7572# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1557 a_27034_6752# a_26967_6160# a_27045_7276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1558 a_24006_7744# a_24263_7554# a_23068_7988# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1559 a_1902_5054# a_1481_5054# a_1803_5054# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1560 a_15942_4814# a_15521_4814# a_15205_4924# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1561 a_432_9180# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1562 a_2774_3071# a_3031_2881# a_2774_5271# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1563 a_10466_910# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1564 vout a_18995_134# a_19317_134# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1565 a_22964_5075# a_23007_7274# a_22958_7464# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1566 a_17974_5670# a_18227_5657# a_17829_6439# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1567 gnd d0 a_14112_1514# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1568 gnd a_34296_2044# a_34088_2044# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1569 a_36858_5654# a_36645_5654# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1570 a_38156_4725# a_39143_4291# a_39094_4481# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1571 a_38047_3098# a_38066_1818# a_38021_1831# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1572 a_36859_2345# a_36646_2345# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1573 a_30337_1742# a_30864_1994# a_31072_1994# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1574 a_24012_4812# a_24265_4799# a_23073_4502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1575 vdd d1 a_13172_3410# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1576 a_21770_7814# a_21557_7814# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1577 gnd d2 a_8055_6244# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1578 a_8882_5975# a_8878_6152# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1579 gnd a_39352_4845# a_39144_4845# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1580 a_20305_3756# a_20834_3646# a_21042_3646# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1581 a_116_8831# a_117_8374# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1582 vdd d1 a_8195_7858# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1583 a_31589_5613# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1584 a_21771_4505# a_21558_4505# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1585 a_26614_4546# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1586 a_11755_8349# a_11542_8349# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1587 a_13855_6488# a_14108_6475# a_12913_6909# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1588 a_6849_5668# a_6428_5668# a_5911_5912# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1589 a_32991_3057# a_33010_1777# a_32961_1967# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1590 a_27047_2864# a_26756_1748# a_27036_2340# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1591 a_1808_5173# a_1481_7254# a_1808_7373# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1592 gnd d4 a_23217_5062# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1593 vdd a_8056_4038# a_7848_4038# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1594 a_27246_368# a_27137_368# a_25140_307# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1595 vdd a_3139_7817# a_2931_7817# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1596 vdd a_34294_6456# a_34086_6456# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1597 a_436_1459# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1598 vdd d0 a_14110_5926# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1599 a_18911_9289# a_19164_9276# a_17972_8979# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1600 a_24008_3332# a_24265_3142# a_23070_3576# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1601 a_8880_9284# a_8876_9461# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1602 a_17976_1258# a_18229_1245# a_17831_2027# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1603 a_22960_5252# a_23009_2862# a_22960_3052# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1604 a_17865_5140# a_17908_7339# a_17863_7352# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1605 a_34039_3337# a_34044_2611# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1606 vdd a_38415_1226# a_38207_1226# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1607 a_10675_8631# a_10462_8631# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1608 a_22927_8580# a_23117_7798# a_23068_7988# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1609 a_2778_5094# a_2821_7293# a_2776_7306# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1610 a_16897_3007# a_16600_3978# a_16881_3467# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1611 a_8883_3769# a_8879_3946# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1612 a_38159_7857# a_38412_7844# a_38014_8626# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1613 gnd d2 a_8057_1832# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1614 a_21772_3402# a_21559_3402# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1615 a_34040_8675# a_34036_8852# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1616 a_35704_8653# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1617 a_10148_7089# a_10148_6860# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1618 a_32010_4510# a_31589_4510# a_31071_4200# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1619 a_39096_1172# a_35395_1038# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1620 a_36969_2869# a_36756_2869# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1621 a_21977_8917# a_21910_8325# a_21994_7354# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1622 a_11757_3937# a_11544_3937# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1623 a_37068_1242# a_37000_1753# a_37078_2869# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1624 a_8880_6524# a_8876_6701# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1625 vdd d0 a_34297_2598# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1626 a_853_6420# a_1584_6730# a_1792_6730# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1627 vdd a_34296_2044# a_34088_2044# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1628 a_5173_7312# a_5173_7125# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1629 a_22964_5075# a_23007_7274# a_22962_7287# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1630 a_33099_6890# a_34086_6456# a_34037_6646# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1631 a_31073_891# a_31804_1201# a_32012_1201# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1632 vdd d0 a_14112_1514# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1633 a_31071_5303# a_30650_5303# a_30335_5051# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1634 a_23067_9091# a_23324_8901# a_22931_8403# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1635 a_6780_8385# a_6567_8385# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1636 a_8880_6524# a_9133_6511# a_7938_6945# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1637 a_32959_6379# a_33216_6189# a_32989_7469# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1638 a_18913_4877# a_19166_4864# a_17974_4567# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1639 a_18911_9289# a_18907_9466# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1640 a_11614_8941# a_11401_8941# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1641 a_30334_6841# a_30863_6960# a_31071_6960# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1642 a_21880_5035# a_21667_5035# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1643 gnd a_19164_7619# a_18956_7619# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1644 a_13852_7219# a_13855_6488# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1645 a_12809_5099# a_13062_5086# a_12035_351# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1646 a_20834_2543# a_20621_2543# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1647 vdd d2 a_8055_6244# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1648 a_5174_4690# a_5703_4809# a_5911_4809# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1649 a_30650_6960# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1650 a_15205_5568# a_15733_5363# a_15941_5363# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1651 a_33103_7816# a_33356_7803# a_32958_8585# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1652 gnd d0 a_4077_9230# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1653 a_13851_6665# a_14108_6475# a_12913_6909# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1654 a_17859_7529# a_17878_6249# a_17829_6439# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1655 gnd a_13172_3410# a_12964_3410# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1656 a_22929_4168# a_23119_3386# a_23070_3576# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1657 a_6537_7295# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1658 vdd d4 a_23217_5062# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1659 a_35393_1596# a_35393_1367# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1660 a_35706_4241# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1661 a_17973_6773# a_18957_7070# a_18908_7260# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1662 a_15735_3711# a_15522_3711# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1663 a_37081_5200# a_36754_7281# a_37081_7400# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1664 a_29068_3196# a_29321_3183# a_28126_3617# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1665 a_15521_3157# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1666 vdd d1 a_38411_8947# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1667 a_15941_8123# a_16671_7879# a_16879_7879# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1668 a_18907_9466# a_19164_9276# a_17972_8979# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1669 a_2886_6727# a_3870_7024# a_3821_7214# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1670 gnd a_13030_6208# a_12822_6208# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1671 a_3821_5557# a_3826_4831# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1672 a_6850_3462# a_6429_3462# a_5911_3152# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1673 a_37175_5081# a_37168_373# a_35171_312# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1674 a_32989_7469# a_33246_7279# a_32995_5080# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1675 a_5175_2254# a_5176_1797# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1676 a_855_2008# a_1586_2318# a_1794_2318# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1677 a_6641_4565# a_6428_4565# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1678 a_17972_1435# a_18229_1245# a_17831_2027# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1679 a_33101_2478# a_34088_2044# a_34039_2234# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1680 a_26828_2340# a_26615_2340# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1681 gnd d0 a_24265_5902# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1682 a_10150_3780# a_10679_3670# a_10887_3670# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1683 a_17828_8645# a_18018_7863# a_17969_8053# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1684 a_23069_4679# a_23326_4489# a_22933_3991# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1685 a_2741_8599# a_2998_8409# a_2776_7306# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1686 a_36644_7860# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1687 a_36126_7550# a_35705_7550# a_35390_7755# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1688 a_23072_6708# a_24056_7005# a_24007_7195# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1689 gnd a_29319_9252# a_29111_9252# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1690 a_33105_3404# a_33358_3391# a_32960_4173# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1691 a_29064_5030# a_29067_4299# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1692 a_13853_2253# a_13859_1527# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1693 a_37081_7400# a_36784_8371# a_37064_8963# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1694 a_25358_9083# a_25887_9202# a_26095_9202# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1695 a_33099_6890# a_34086_6456# a_34041_6469# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1696 a_2743_4187# a_2933_3405# a_2888_3418# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1697 a_6958_5095# a_6537_5095# a_6864_5214# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1698 a_15943_3711# a_16673_3467# a_16881_3467# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1699 vdd a_39349_8703# a_39141_8703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1700 a_8876_6701# a_9133_6511# a_7938_6945# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1701 a_22289_327# a_25031_307# a_25239_307# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1702 a_21040_6955# a_21770_6711# a_21978_6711# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1703 gnd d1 a_13171_5616# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1704 vdd d0 a_39353_982# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1705 a_35918_6447# a_35705_6447# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1706 a_12805_5276# a_13062_5086# a_12035_351# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1707 gnd a_14112_1514# a_13904_1514# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1708 a_24010_6464# a_24006_6641# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1709 a_39096_1172# a_39353_982# a_38158_1416# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1710 a_17863_7352# a_18116_7339# a_17865_5140# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1711 a_31072_5857# a_30651_5857# a_30335_5967# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1712 vdd d0 a_4077_9230# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1713 a_31073_2548# a_30652_2548# a_30336_2429# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1714 a_5910_8118# a_5489_8118# a_5173_8228# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1715 gnd a_8055_6244# a_7847_6244# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1716 vdd a_13172_3410# a_12964_3410# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1717 a_35392_2470# a_35392_2240# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1718 a_22929_4168# a_23119_3386# a_23074_3399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1719 a_20830_8607# a_20617_8607# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1720 vdd a_8195_7858# a_7987_7858# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1721 a_16812_6184# a_16599_6184# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1722 a_30649_6406# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1723 a_7937_9151# a_8924_8717# a_8879_8730# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1724 a_17973_6773# a_18957_7070# a_18912_7083# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1725 vdd d0 a_14109_4269# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1726 a_36128_3138# a_35707_3138# a_35392_3343# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1727 a_24011_5361# a_24264_5348# a_23069_5782# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1728 gnd a_29321_4840# a_29113_4840# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1729 a_29064_3373# a_29321_3183# a_28126_3617# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1730 a_1793_5627# a_1372_5627# a_854_5317# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1731 gnd a_23217_5062# a_23009_5062# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1732 a_32320_332# a_31899_332# a_32221_332# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1733 a_2886_6727# a_3870_7024# a_3825_7037# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1734 a_11543_6143# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1735 a_1791_8936# a_1370_8936# a_853_9180# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1736 a_30864_4754# a_30651_4754# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1737 a_33101_2478# a_34088_2044# a_34043_2057# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1738 vdd d0 a_29319_6492# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1739 vdd a_39351_4291# a_39143_4291# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1740 a_35390_8214# a_35390_7985# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1741 a_35919_5344# a_35706_5344# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1742 a_8878_2289# a_9135_2099# a_7940_2533# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1743 gnd d1 a_8196_5652# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1744 a_5176_1381# a_5176_1151# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1745 a_27033_8958# a_26966_8366# a_27050_7395# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1746 gnd d0 a_39351_5394# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1747 a_31074_1445# a_30653_1445# a_30337_1555# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1748 a_17865_2940# a_18118_2927# a_17861_5317# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1749 vdd a_29319_9252# a_29111_9252# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1750 a_10462_8631# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1751 a_20831_7504# a_20618_7504# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1752 gnd a_3140_5611# a_2932_5611# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1753 a_25360_5087# a_25360_4900# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1754 gnd a_8057_1832# a_7849_1832# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1755 a_36756_2869# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1756 a_36857_7860# a_36644_7860# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1757 a_38155_6931# a_39142_6497# a_39093_6687# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1758 gnd a_4081_1509# a_3873_1509# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1759 vdd d1 a_33356_6700# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1760 a_24013_949# a_24266_936# a_23071_1370# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1761 a_34043_3160# a_34039_3337# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1762 a_16670_8982# a_16457_8982# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1763 a_5489_5358# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1764 a_32011_2304# a_31944_1712# a_32022_2828# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1765 a_1795_1215# a_1374_1215# a_856_905# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1766 vdd d1 a_13171_5616# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1767 a_8883_1009# a_8879_1186# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1768 vdd a_34297_2598# a_34089_2598# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1769 a_31911_7240# a_31698_7240# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1770 a_30865_3651# a_30652_3651# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1771 a_31588_7819# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1772 a_5174_4690# a_5174_4460# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1773 vdd a_14112_1514# a_13904_1514# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1774 gnd d0 a_9133_9271# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1775 a_11401_8941# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1776 vdd a_8055_6244# a_7847_6244# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1777 gnd d1 a_8198_1240# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1778 a_20621_2543# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1779 gnd d0 a_39353_982# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1780 gnd a_4077_9230# a_3869_9230# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1781 a_15943_2608# a_15522_2608# a_15206_2718# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1782 a_21996_2942# a_21882_2823# a_21989_5035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1783 a_20833_3092# a_20620_3092# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1784 vdd a_23217_5062# a_23009_5062# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1785 a_15522_3711# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1786 a_20305_3756# a_20305_3527# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1787 a_38157_2519# a_39144_2085# a_39095_2275# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1788 a_36859_3448# a_36646_3448# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1789 a_16672_4570# a_16459_4570# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1790 vdd d1 a_33358_2288# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1791 a_15204_8004# a_15204_7774# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1792 a_30334_6611# a_30335_6154# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1793 a_21771_5608# a_21558_5608# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1794 gnd d2 a_8056_4038# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1795 vdd d1 a_13173_1204# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1796 vdd d1 a_8196_5652# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1797 a_26615_2340# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1798 a_16895_7419# a_16781_7300# a_16895_5219# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1799 gnd a_24265_5902# a_24057_5902# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1800 a_2774_5271# a_2823_2881# a_2778_2894# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1801 a_34037_9406# a_34040_8675# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1802 a_13856_4282# a_14109_4269# a_12914_4703# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1803 gnd d4 a_3031_5081# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1804 vdd d0 a_34296_4804# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1805 a_18915_1568# a_18911_1745# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1806 vdd a_3140_5611# a_2932_5611# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1807 a_3825_5380# a_3821_5557# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1808 a_31070_7509# a_30649_7509# a_30334_7257# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1809 gnd d1 a_38412_6741# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1810 a_30865_891# a_30652_891# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1811 a_8879_8730# a_9132_8717# a_7937_9151# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1812 a_32958_8585# a_33215_8395# a_32993_7292# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1813 a_18912_4323# a_18908_4500# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1814 a_31698_5040# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1815 a_20833_4749# a_20620_4749# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1816 a_20306_1321# a_20306_1091# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1817 a_25140_307# a_26924_368# a_27144_5076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1818 a_32961_1967# a_33218_1777# a_32991_3057# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1819 a_15204_7774# a_15732_7569# a_15940_7569# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1820 a_15205_5111# a_15205_4924# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1821 a_26969_1748# a_26756_1748# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1822 a_3827_2625# a_3823_2802# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1823 a_5911_3152# a_5490_3152# a_5175_2900# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1824 vdd d0 a_9133_9271# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1825 a_10676_6425# a_10463_6425# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1826 a_16878_8982# a_16811_8390# a_16895_7419# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1827 a_32010_5613# a_31589_5613# a_31072_5857# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1828 a_21773_1196# a_21560_1196# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1829 a_35705_6447# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1830 vdd d1 a_8198_1240# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1831 a_32011_2304# a_31590_2304# a_31072_1994# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1832 a_17972_8979# a_18956_9276# a_18907_9466# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1833 a_15734_5917# a_15521_5917# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1834 a_2883_5801# a_3870_5367# a_3825_5380# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1835 a_1791_8936# a_1724_8344# a_1808_7373# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1836 a_21978_6711# a_21911_6119# a_21989_7235# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1837 a_29067_5402# a_29320_5389# a_28125_5823# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1838 vdd a_4077_9230# a_3869_9230# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1839 a_24013_949# a_24009_1126# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1840 a_15732_9226# a_15519_9226# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1841 a_30334_7070# a_30863_6960# a_31071_6960# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1842 a_20304_4630# a_20304_4400# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1843 a_36129_3692# a_35708_3692# a_35392_3802# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1844 gnd a_28380_8942# a_28172_8942# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1845 a_29065_3927# a_29322_3737# a_28130_3440# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1846 gnd d0 a_24264_8108# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1847 a_10149_5986# a_10678_5876# a_10886_5876# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1848 a_38157_2519# a_39144_2085# a_39099_2098# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1849 a_23068_6885# a_23325_6695# a_22932_6197# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1850 a_11615_6735# a_11402_6735# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1851 a_39095_6138# a_39098_5407# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1852 gnd d1 a_18229_1245# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1853 a_646_6974# a_433_6974# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1854 a_853_9180# a_432_9180# a_116_9061# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1855 a_16599_6184# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1856 a_33105_2301# a_34089_2598# a_34044_2611# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1857 a_30651_4754# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1858 gnd d0 a_4078_7024# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1859 a_20303_6606# a_20831_6401# a_21039_6401# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1860 a_33104_5610# a_33357_5597# a_32959_6379# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1861 a_25031_307# a_24818_307# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1862 a_17835_1850# a_18020_2348# a_17971_2538# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1863 a_35706_5344# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1864 a_30863_5303# a_30650_5303# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1865 a_32012_1201# a_31591_1201# a_31074_1445# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1866 a_10678_2013# a_10465_2013# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1867 gnd a_8196_5652# a_7988_5652# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1868 vdd d4 a_3031_5081# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1869 a_35707_2035# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1870 a_7938_6945# a_8925_6511# a_8876_6701# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1871 a_17974_4567# a_18958_4864# a_18909_5054# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1872 a_15736_1505# a_15523_1505# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1873 gnd d0 a_14110_2063# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1874 gnd d3 a_8085_7334# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1875 a_29069_990# a_29322_977# a_28127_1411# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1876 vdd d1 a_38412_6741# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1877 a_12035_351# a_12854_5086# a_12805_5276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1878 a_2887_4521# a_3871_4818# a_3822_5008# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1879 a_6851_1256# a_6430_1256# a_5912_946# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1880 a_21039_9161# a_21769_8917# a_21977_8917# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1881 a_10147_8836# a_10148_8379# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1882 a_6642_2359# a_6429_2359# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1883 a_7830_3112# a_8087_2922# a_7830_5312# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1884 vdd a_33356_6700# a_33148_6700# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1885 a_11616_5632# a_11403_5632# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1886 a_10151_1574# a_10680_1464# a_10888_1464# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1887 a_2742_6393# a_2999_6203# a_2772_7483# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1888 a_647_5871# a_434_5871# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1889 a_2883_4698# a_3140_4508# a_2747_4010# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1890 a_11617_2323# a_11404_2323# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1891 a_36645_5654# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1892 a_5488_9221# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1893 a_36967_7281# a_36754_7281# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1894 a_8883_2666# a_8879_2843# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1895 a_648_2562# a_435_2562# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1896 a_30652_3651# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1897 a_16879_7879# a_16458_7879# a_15940_7569# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1898 a_17972_8979# a_18956_9276# a_18911_9289# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1899 a_36643_8963# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1900 gnd a_9133_9271# a_8925_9271# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1901 gnd a_29320_7046# a_29112_7046# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1902 a_33106_1198# a_33359_1185# a_32961_1967# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1903 a_27052_2983# a_26938_2864# a_27045_5076# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1904 a_29061_8888# a_29067_8162# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1905 a_35708_932# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1906 a_37076_7281# a_36785_6165# a_37065_6757# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1907 a_10887_3670# a_10466_3670# a_10150_3551# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1908 gnd a_8198_1240# a_7990_1240# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1909 a_11542_8349# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1910 a_25359_6877# a_25888_6996# a_26096_6996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1911 a_3824_9243# a_3820_9420# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1912 a_24008_6092# a_24265_5902# a_23073_5605# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1913 gnd a_39353_982# a_39145_982# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1914 gnd d3 a_8087_2922# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1915 vdd d1 a_38414_2329# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1916 a_21039_7504# a_21770_7814# a_21978_7814# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1917 a_8877_4495# a_9134_4305# a_7939_4739# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1918 a_35392_3343# a_35392_2886# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1919 a_20620_3092# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1920 a_35918_7550# a_35705_7550# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1921 vdd d1 a_18229_1245# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1922 a_21041_4749# a_21771_4505# a_21979_4505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1923 vdd d3 a_28273_2903# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1924 a_1727_1726# a_1514_1726# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1925 a_15731_8672# a_15518_8672# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1926 vdd a_33358_2288# a_33150_2288# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1927 a_36997_8371# a_36784_8371# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1928 vdd d0 a_4078_7024# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1929 a_36647_1242# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1930 vdd a_13173_1204# a_12965_1204# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1931 a_30649_7509# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1932 gnd a_8056_4038# a_7848_4038# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1933 a_12917_7835# a_13170_7822# a_12772_8604# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1934 vdd a_8196_5652# a_7988_5652# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1935 vdd d0 a_39352_5948# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1936 a_7938_6945# a_8925_6511# a_8880_6524# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1937 vdd d0 a_14110_2063# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1938 a_11727_2847# a_11514_2847# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1939 vdd d1 a_33355_8906# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1940 vdd d3 a_8085_7334# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1941 a_21978_6711# a_21557_6711# a_21039_6401# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1942 a_37168_373# a_36955_373# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1943 a_5176_1610# a_5705_1500# a_5913_1500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1944 a_12035_351# a_12854_5086# a_12809_5099# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1945 gnd d0 a_19163_8722# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1946 vdd a_34296_4804# a_34088_4804# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1947 a_17865_5140# a_17908_7339# a_17859_7529# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1948 a_30864_5857# a_30651_5857# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1949 a_27246_368# a_28065_5103# a_28016_5293# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1950 a_29752_191# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1951 a_24010_1680# a_24267_1490# a_23075_1193# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1952 a_30865_2548# a_30652_2548# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1953 a_6567_8385# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1954 vdd a_3029_7293# a_2821_7293# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1955 gnd a_38412_6741# a_38204_6741# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1956 a_21996_2942# a_21699_3913# a_21979_4505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1957 a_39094_5584# a_39099_4858# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1958 a_21041_3092# a_21772_3402# a_21980_3402# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1959 a_20620_4749# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1960 gnd d1 a_8197_3446# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1961 a_26756_1748# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1962 a_15733_4260# a_15520_4260# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1963 gnd d0 a_39352_3188# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1964 vdd a_29320_7046# a_29112_7046# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1965 vdd a_9133_9271# a_8925_9271# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1966 a_10463_6425# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1967 a_118_6168# a_118_5981# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1968 a_20832_5298# a_20619_5298# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1969 a_33102_1375# a_33359_1185# a_32961_1967# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1970 a_25358_9083# a_25358_8853# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1971 a_32025_7359# a_31728_8330# a_32008_8922# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1972 a_21560_1196# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1973 a_18914_1014# a_19167_1001# a_17972_1435# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1974 a_15521_5917# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1975 vdd a_8198_1240# a_7990_1240# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1976 a_5174_5563# a_5174_5106# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1977 a_7940_2533# a_8927_2099# a_8882_2112# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1978 a_6848_7874# a_6780_8385# a_6864_7414# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1979 vdd d1 a_33357_4494# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1980 a_3827_968# a_4080_955# a_2885_1389# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1981 a_16671_6776# a_16458_6776# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1982 a_21989_5035# a_21880_5035# a_22088_5035# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1983 a_20619_8058# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1984 a_10886_5876# a_11616_5632# a_11824_5632# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1985 gnd d0 a_19165_4310# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1986 a_34041_1685# a_34044_954# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1987 a_18906_8912# a_18912_8186# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1988 a_28124_8029# a_28381_7839# a_27983_8621# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1989 a_30866_1445# a_30653_1445# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1990 a_35393_1137# a_35921_932# a_36129_932# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1991 a_38161_2342# a_39145_2639# a_39100_2652# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1992 a_15204_8233# a_15204_8004# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1993 gnd a_24264_8108# a_24056_8108# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1994 a_13857_5939# a_14110_5926# a_12918_5629# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1995 a_10883_8631# a_11614_8941# a_11822_8941# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1996 gnd d0 a_9134_7065# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1997 a_37066_4551# a_36645_4551# a_36128_4795# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1998 a_11402_6735# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1999 a_25359_6647# a_25887_6442# a_26095_6442# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2000 a_433_6974# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2001 a_13852_5562# a_13857_4836# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2002 a_2884_3595# a_3871_3161# a_3822_3351# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2003 a_24005_8847# a_24262_8657# a_23067_9091# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2004 gnd a_4078_7024# a_3870_7024# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2005 a_645_7523# a_432_7523# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2006 a_20834_886# a_20621_886# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2007 a_10465_2013# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2008 a_1810_2961# a_1696_2842# a_1803_5054# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2009 a_30650_5303# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2010 vdd d0 a_19163_8722# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2011 a_12917_7835# a_13901_8132# a_13852_8322# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2012 a_32993_7292# a_33246_7279# a_32995_5080# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2013 a_17973_6773# a_18226_6760# a_17833_6262# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2014 a_32960_4173# a_33217_3983# a_32995_2880# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2015 a_29070_1544# a_29323_1531# a_28131_1234# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2016 a_15523_1505# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2017 vdd a_38412_6741# a_38204_6741# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2018 a_16672_5673# a_16459_5673# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2019 a_5910_5358# a_5489_5358# a_5174_5106# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2020 gnd a_23184_8390# a_22976_8390# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2021 a_23072_7811# a_24056_8108# a_24011_8121# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2022 a_12035_351# a_11926_351# a_12134_351# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2023 a_10888_1464# a_11618_1220# a_11826_1220# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2024 a_16673_2364# a_16460_2364# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2025 a_26924_368# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2026 a_28126_3617# a_28383_3427# a_27985_4209# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2027 a_35391_5779# a_35391_5549# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2028 vdd d1 a_8197_3446# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2029 a_2103_346# a_1682_346# a_1902_5054# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2030 a_10150_3321# a_10150_2864# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2031 a_6848_6771# a_6427_6771# a_5910_7015# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2032 a_11403_5632# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2033 a_434_5871# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2034 a_25361_2235# a_25889_2030# a_26097_2030# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2035 a_11404_2323# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2036 a_435_2562# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2037 a_36754_7281# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2038 vdd a_3141_3405# a_2933_3405# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2039 a_29064_6133# a_29321_5943# a_28129_5646# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2040 gnd d1 a_38413_4535# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2041 a_3823_3905# a_3826_3174# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2042 a_34043_2057# a_34039_2234# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2043 a_647_3111# a_434_3111# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2044 a_16895_5219# a_16568_7300# a_16890_7300# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2045 vdd d0 a_4078_5367# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2046 a_32020_7240# a_31729_6124# a_32010_5613# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2047 a_33104_4507# a_34088_4804# a_34043_4817# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2048 vdd d0 a_19165_4310# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2049 a_32995_2880# a_33248_2867# a_32991_5257# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2050 a_29064_3373# a_29069_2647# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2051 a_29066_9265# a_30333_9276# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2052 a_16598_8390# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2053 a_15203_9107# a_15203_8877# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2054 a_6783_1767# a_6570_1767# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2055 a_16674_1261# a_16461_1261# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2056 vdd a_38414_2329# a_38206_2329# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2057 a_20302_8812# a_20830_8607# a_21038_8607# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2058 vdd d0 a_9134_7065# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2059 a_11758_1731# a_11545_1731# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2060 a_35705_7550# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2061 a_30862_7509# a_30649_7509# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2062 a_16879_6776# a_16812_6184# a_16890_7300# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2063 a_10677_4219# a_10464_4219# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2064 vdd a_28273_2903# a_28065_2903# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2065 a_32011_3407# a_31590_3407# a_31073_3651# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2066 a_20304_5503# a_20304_5046# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2067 a_36130_1486# a_35709_1486# a_35393_1367# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2068 a_7937_9151# a_8924_8717# a_8875_8907# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2069 gnd d0 a_14109_4269# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2070 a_2884_3595# a_3871_3161# a_3826_3174# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2071 a_1514_1726# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2072 a_16783_2888# a_16570_2888# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2073 a_36784_8371# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2074 a_1792_6730# a_1725_6138# a_1803_7254# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2075 vdd d2 a_13032_1796# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2076 vdd a_4078_7024# a_3870_7024# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2077 a_15733_7020# a_15520_7020# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2078 a_16882_1261# a_16814_1772# a_16892_2888# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2079 a_21994_5154# a_21667_7235# a_21989_7235# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2080 a_12917_7835# a_13901_8132# a_13856_8145# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2081 a_17969_6950# a_18226_6760# a_17833_6262# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2082 vdd a_39352_5948# a_39144_5948# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2083 vdd d0 a_14111_2617# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2084 a_29066_1721# a_29323_1531# a_28131_1234# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2085 a_20305_2653# a_20305_2424# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2086 a_11514_2847# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2087 vdd a_33355_8906# a_33147_8906# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2088 a_16895_7419# a_16598_8390# a_16879_7879# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2089 a_5173_7999# a_5173_7769# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2090 a_11615_7838# a_11402_7838# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2091 a_12773_6398# a_13030_6208# a_12803_7488# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2092 a_11616_4529# a_11403_4529# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2093 a_35921_3692# a_35708_3692# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2094 gnd a_19163_8722# a_18955_8722# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2095 a_21989_5035# a_21669_2823# a_21996_2942# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2096 a_117_8374# a_644_8626# a_852_8626# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2097 a_1808_7373# a_1511_8344# a_1792_7833# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2098 a_10148_6860# a_10677_6979# a_10885_6979# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2099 a_30651_5857# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2100 a_647_4768# a_434_4768# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2101 a_34044_3714# a_34040_3891# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2102 a_30652_2548# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2103 a_20303_7252# a_20831_7504# a_21039_7504# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2104 a_38155_8034# a_39142_7600# a_39097_7613# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2105 a_35707_3138# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2106 a_10886_5876# a_10465_5876# a_10149_5757# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2107 gnd a_8197_3446# a_7989_3446# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2108 vdd d3 a_13062_2886# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2109 a_2745_8422# a_2930_8920# a_2885_8933# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2110 a_3825_4277# a_3821_4454# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2111 gnd d0 a_39353_3742# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2112 a_15520_4260# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2113 gnd a_39352_3188# a_39144_3188# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2114 a_30336_3761# a_30336_3532# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2115 a_15940_9226# a_16670_8982# a_16878_8982# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2116 a_27045_5076# a_26936_5076# a_27144_5076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2117 vdd d1 a_38413_4535# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2118 a_32025_7359# a_31911_7240# a_32025_5159# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2119 a_17971_2538# a_18228_2348# a_17835_1850# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2120 a_21039_6401# a_20618_6401# a_20304_6149# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2121 a_25361_3568# a_25361_3338# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2122 vdd a_33357_4494# a_33149_4494# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2123 a_11617_3426# a_11404_3426# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2124 a_39096_8716# a_39349_8703# a_38154_9137# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2125 a_16890_7300# a_16599_6184# a_16879_6776# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2126 vdd a_3001_1791# a_2793_1791# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2127 a_2884_2492# a_3141_2302# a_2748_1804# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2128 gnd a_19165_4310# a_18957_4310# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2129 a_648_3665# a_435_3665# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2130 a_36646_3448# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2131 a_5489_7015# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2132 a_119_3962# a_646_4214# a_854_4214# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2133 a_30653_1445# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2134 a_36125_8653# a_35704_8653# a_35389_8858# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2135 a_30334_7070# a_30334_6841# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2136 a_20305_2840# a_20833_3092# a_21041_3092# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2137 a_21977_8917# a_21556_8917# a_21038_8607# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2138 gnd a_9134_7065# a_8926_7065# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2139 a_5175_3816# a_5704_3706# a_5912_3706# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2140 a_25890_927# a_25677_927# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2141 a_20833_1989# a_20620_1989# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2142 a_38157_3622# a_39144_3188# a_39099_3201# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2143 a_18909_6157# a_19166_5967# a_17974_5670# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2144 a_37083_2988# a_36786_3959# a_37066_4551# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2145 a_10888_1464# a_10467_1464# a_10151_1345# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2146 a_7830_5312# a_7879_2922# a_7834_2935# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2147 a_12912_9115# a_13169_8925# a_12776_8427# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2148 a_11725_5059# a_11512_5059# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2149 a_2747_4010# a_2932_4508# a_2887_4521# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2150 a_24009_3886# a_24266_3696# a_23074_3399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2151 a_15942_4814# a_16672_4570# a_16880_4570# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2152 a_15204_8420# a_15204_8233# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2153 a_28128_7852# a_29112_8149# a_29067_8162# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2154 a_432_7523# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2155 a_20621_886# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2156 vdd a_19163_8722# a_18955_8722# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2157 a_21040_5298# a_21771_5608# a_21979_5608# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2158 a_28129_5646# a_28382_5633# a_27984_6415# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2159 a_39095_5035# a_39098_4304# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2160 a_5175_2900# a_5175_2713# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2161 a_5911_5912# a_5490_5912# a_5174_5793# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2162 vdd a_3031_2881# a_2823_2881# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2163 a_15732_6466# a_15519_6466# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2164 a_36998_6165# a_36785_6165# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2165 a_16460_2364# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2166 a_18913_3220# a_19166_3207# a_17971_3641# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2167 a_36127_4241# a_35706_4241# a_35391_4446# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2168 vdd a_8197_3446# a_7989_3446# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2169 vdd d0 a_39353_3742# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2170 a_21910_8325# a_21697_8325# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2171 a_20303_7939# a_20303_7709# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2172 a_21978_7814# a_21557_7814# a_21040_8058# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2173 a_24010_6464# a_24263_6451# a_23068_6885# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2174 gnd d0 a_4079_5921# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2175 a_7939_4739# a_8926_4305# a_8881_4318# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2176 gnd d1 a_33359_1185# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2177 a_31729_6124# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2178 a_26097_5893# a_25676_5893# a_25360_5774# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2179 a_1792_6730# a_1371_6730# a_853_6420# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2180 a_21979_4505# a_21558_4505# a_21040_4195# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2181 gnd d0 a_4077_7573# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2182 a_10885_8082# a_11615_7838# a_11823_7838# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2183 gnd d0 a_19164_6516# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2184 a_20304_4630# a_20833_4749# a_21041_4749# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2185 a_38051_2921# a_38304_2908# a_38047_5298# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2186 a_38160_4548# a_39144_4845# a_39099_4858# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2187 a_32965_1790# a_33218_1777# a_32991_3057# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2188 a_32965_1790# a_33150_2288# a_33101_2478# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2189 a_29965_191# a_29752_191# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2190 a_24014_1503# a_24010_1680# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2191 a_3824_1699# a_4081_1509# a_2889_1212# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2192 a_6568_6179# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2193 a_37065_6757# a_36644_6757# a_36127_7001# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2194 gnd a_38413_4535# a_38205_4535# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2195 a_25358_8853# a_25886_8648# a_26094_8648# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2196 a_8881_8181# a_8877_8358# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2197 a_434_3111# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2198 a_12772_8604# a_12962_7822# a_12913_8012# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2199 a_21042_886# a_21773_1196# a_21981_1196# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2200 a_28131_1234# a_28384_1221# a_27986_2003# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2201 vdd a_4078_5367# a_3870_5367# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2202 vdd a_19165_4310# a_18957_4310# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2203 a_2883_5801# a_3870_5367# a_3821_5557# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2204 a_15733_5363# a_15520_5363# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2205 a_5913_1500# a_5492_1500# a_5176_1381# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2206 a_16461_1261# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2207 a_15734_2054# a_15521_2054# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2208 a_6570_1767# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2209 a_15203_9107# a_15732_9226# a_15940_9226# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2210 vdd a_9134_7065# a_8926_7065# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2211 a_10464_4219# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2212 a_21912_3913# a_21699_3913# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2213 a_29069_3750# a_29322_3737# a_28130_3440# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2214 a_16570_2888# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2215 a_10677_8082# a_10464_8082# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2216 a_16671_7879# a_16458_7879# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2217 a_26099_1481# a_25678_1481# a_25362_1362# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2218 vdd a_13032_1796# a_12824_1796# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2219 a_5488_6461# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2220 a_1803_5054# a_1694_5054# a_1902_5054# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2221 gnd a_29319_7595# a_29111_7595# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2222 a_15520_7020# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2223 vdd d1 a_13170_6719# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2224 a_10887_3670# a_11617_3426# a_11825_3426# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2225 a_28125_5823# a_28382_5633# a_27984_6415# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2226 a_25359_7293# a_25887_7545# a_26095_7545# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2227 a_11402_7838# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2228 gnd d0 a_9135_4859# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2229 a_17972_1435# a_18959_1001# a_18910_1191# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2230 a_37067_2345# a_36646_2345# a_36129_2589# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2231 vdd d2 a_23184_8390# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2232 a_30335_5508# a_30863_5303# a_31071_5303# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2233 a_11403_4529# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2234 a_25360_4441# a_25888_4236# a_26096_4236# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2235 a_434_4768# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2236 a_32221_332# a_32112_332# a_32320_332# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2237 a_6864_7414# a_6567_8385# a_6847_8977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2238 a_15735_951# a_15522_951# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2239 a_1682_346# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2240 a_2885_1389# a_3872_955# a_3823_1145# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2241 vdd d1 a_33359_1185# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2242 a_2103_346# a_4845_326# a_5053_326# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2243 a_24006_6641# a_24263_6451# a_23068_6885# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2244 a_20305_2840# a_20305_2653# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2245 a_646_5317# a_433_5317# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2246 gnd a_4079_4818# a_3871_4818# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2247 a_35708_3692# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2248 a_3824_9243# a_5172_9331# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2249 a_35390_8214# a_35919_8104# a_36127_8104# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2250 a_37081_7400# a_36967_7281# a_37081_5200# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2251 a_33106_1198# a_34090_1495# a_34041_1685# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2252 vdd d0 a_4077_7573# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2253 vdd d0 a_19164_6516# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2254 a_12918_5629# a_13902_5926# a_13853_6116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2255 a_17974_4567# a_18227_4554# a_17834_4056# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2256 a_36858_4551# a_36645_4551# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2257 vdd a_13062_2886# a_12854_2886# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2258 gnd a_39353_3742# a_39145_3742# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2259 a_26096_8099# a_26826_7855# a_27034_7855# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2260 a_32993_7292# a_33007_8395# a_32958_8585# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2261 a_21040_8058# a_20619_8058# a_20303_8168# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2262 gnd a_23185_6184# a_22977_6184# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2263 vdd a_38413_4535# a_38205_4535# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2264 a_16673_3467# a_16460_3467# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2265 a_11757_3937# a_11544_3937# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2266 a_20305_2653# a_20834_2543# a_21042_2543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2267 vdd d1 a_13172_2307# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2268 a_21770_6711# a_21557_6711# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2269 a_28127_1411# a_28384_1221# a_27986_2003# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2270 a_4845_326# a_4632_326# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2271 gnd a_29321_3183# a_29113_3183# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2272 a_39094_4481# a_39100_3755# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2273 a_1803_5054# a_1483_2842# a_1805_2842# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2274 a_11404_3426# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2275 a_25361_2881# a_25889_3133# a_26097_3133# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2276 a_6849_4565# a_6428_4565# a_5911_4809# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2277 a_435_3665# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2278 a_17968_9156# a_18225_8966# a_17832_8468# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2279 vdd d0 a_14110_4823# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2280 a_2746_6216# a_2931_6714# a_2882_6904# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2281 a_2885_1389# a_3872_955# a_3827_968# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2282 a_37076_5081# a_36756_2869# a_37083_2988# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2283 a_2886_7830# a_3139_7817# a_2741_8599# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2284 a_25891_1481# a_25678_1481# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2285 gnd d1 a_38414_2329# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2286 a_24008_2229# a_24265_2039# a_23070_2473# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2287 a_20620_1989# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2288 gnd d1 a_23326_5592# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2289 a_35920_5898# a_35707_5898# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2290 a_34040_1131# a_30339_997# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2291 vdd d0 a_19166_2104# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2292 a_15203_8877# a_15731_8672# a_15939_8672# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2293 gnd a_8087_5122# a_7879_5122# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2294 a_11512_5059# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2295 a_26098_3687# a_26828_3443# a_27036_3443# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2296 a_22932_6197# a_23117_6695# a_23068_6885# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2297 a_32995_2880# a_33009_3983# a_32960_4173# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2298 a_10149_6173# a_10149_5986# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2299 a_15205_5798# a_15205_5568# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2300 a_9888_210# a_9779_210# a_9987_210# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2301 a_14876_331# a_14663_331# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2302 a_28018_7328# a_28271_7315# a_28020_5116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2303 a_13852_4459# a_13858_3733# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2304 a_20619_5298# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2305 a_36785_6165# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2306 a_18914_3774# a_19167_3761# a_17975_3464# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2307 a_17970_4744# a_18227_4554# a_17834_4056# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2308 a_3827_3728# a_4080_3715# a_2888_3418# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2309 a_31071_4200# a_30650_4200# a_30336_3948# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2310 a_12916_1394# a_13903_960# a_13858_973# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2311 vdd a_39353_3742# a_39145_3742# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2312 a_21038_8607# a_20617_8607# a_20303_8355# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2313 a_28129_5646# a_29113_5943# a_29064_6133# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2314 vdd a_23185_6184# a_22977_6184# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2315 gnd d1 a_23328_1180# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2316 a_35922_1486# a_35709_1486# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2317 a_854_8077# a_433_8077# a_117_8187# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2318 gnd a_4077_7573# a_3869_7573# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2319 gnd a_19164_6516# a_18956_6516# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2320 a_12774_4192# a_13031_4002# a_12809_2899# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2321 vdd a_29321_3183# a_29113_3183# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2322 vdd d1 a_3138_8920# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2323 a_118_6168# a_645_6420# a_853_6420# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2324 a_1803_7254# a_1512_6138# a_1793_5627# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2325 a_15205_4465# a_15733_4260# a_15941_4260# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2326 a_35391_4676# a_35391_4446# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2327 a_33103_6713# a_33356_6700# a_32963_6202# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2328 a_20304_5046# a_20832_5298# a_21040_5298# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2329 a_16892_2888# a_16601_1772# a_16881_2364# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2330 a_10150_2218# a_10151_1761# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2331 a_38156_5828# a_39143_5394# a_39098_5407# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2332 a_22934_1785# a_23119_2283# a_23070_2473# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2333 a_24010_9224# a_25358_9312# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2334 a_852_8626# a_1583_8936# a_1791_8936# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2335 a_118_5522# a_118_5065# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2336 a_16781_5100# a_16568_5100# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2337 a_38047_5298# a_38304_5108# a_37277_373# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2338 a_2746_6216# a_2931_6714# a_2886_6727# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2339 a_15520_5363# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2340 gnd d0 a_39354_1536# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2341 a_12803_7488# a_12822_6208# a_12777_6221# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2342 a_29068_2093# a_29321_2080# a_28126_2514# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2343 a_15521_2054# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2344 a_15941_7020# a_16671_6776# a_16879_6776# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2345 a_21882_2823# a_21669_2823# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2346 a_10885_6979# a_10464_6979# a_10148_7089# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2347 gnd d0 a_9135_3202# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2348 a_38161_2342# a_39145_2639# a_39096_2829# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2349 a_21039_7504# a_20618_7504# a_20303_7709# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2350 a_29068_4853# a_29064_5030# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2351 a_29064_2270# a_29070_1544# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2352 a_119_2672# a_119_2443# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2353 a_10464_8082# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2354 vdd a_8087_5122# a_7879_5122# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2355 a_11618_1220# a_11405_1220# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2356 a_39096_3932# a_39099_3201# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2357 gnd a_4079_3161# a_3871_3161# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2358 a_649_1459# a_436_1459# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2359 a_16878_8982# a_16457_8982# a_15939_8672# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2360 a_36126_6447# a_35705_6447# a_35390_6652# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2361 a_120_1756# a_647_2008# a_855_2008# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2362 a_24009_8670# a_24262_8657# a_23067_9091# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2363 a_28014_7505# a_28271_7315# a_28020_5116# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2364 a_31728_8330# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2365 gnd a_9135_4859# a_8927_4859# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2366 a_1791_8936# a_1370_8936# a_852_8626# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2367 a_18910_3951# a_19167_3761# a_17975_3464# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2368 a_12920_1217# a_13173_1204# a_12775_1986# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2369 gnd a_14109_8132# a_13901_8132# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2370 a_20303_8168# a_20303_7939# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2371 a_34042_5366# a_34038_5543# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2372 a_10150_3780# a_10150_3551# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2373 a_15522_951# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2374 a_21041_3092# a_20620_3092# a_20305_2840# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2375 a_15941_5363# a_16672_5673# a_16880_5673# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2376 a_3823_3905# a_4080_3715# a_2888_3418# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2377 a_2748_1804# a_2933_2302# a_2888_2315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2378 a_10148_7963# a_10677_8082# a_10885_8082# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2379 a_18908_7260# a_18911_6529# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2380 a_8882_3215# a_8878_3392# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2381 a_15943_2608# a_16673_2364# a_16881_2364# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2382 a_433_5317# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2383 gnd d1 a_13171_4513# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2384 a_35917_8653# a_35704_8653# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2385 a_5173_6896# a_5173_6666# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2386 vdd d1 a_23328_1180# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2387 a_28130_3440# a_28383_3427# a_27985_4209# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2388 vdd a_4077_7573# a_3869_7573# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2389 vdd a_19164_6516# a_18956_6516# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2390 a_15732_7569# a_15519_7569# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2391 a_5912_3706# a_5491_3706# a_5175_3587# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2392 a_23075_1193# a_24059_1490# a_24010_1680# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2393 a_34044_2611# a_34040_2788# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2394 a_6859_5095# a_6539_2883# a_6861_2883# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2395 gnd d0 a_39349_8703# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2396 a_2776_7306# a_3029_7293# a_2778_5094# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2397 a_17974_5670# a_18958_5967# a_18913_5980# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2398 a_31072_4754# a_30651_4754# a_30335_4864# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2399 a_16460_3467# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2400 a_18913_5980# a_18909_6157# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2401 a_36999_3959# a_36786_3959# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2402 a_22934_1785# a_23119_2283# a_23074_2296# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2403 a_30648_8612# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2404 a_5910_7015# a_5489_7015# a_5173_7125# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2405 a_13854_3910# a_13857_3179# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2406 vdd a_13172_2307# a_12964_2307# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2407 a_2887_5624# a_3871_5921# a_3826_5934# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2408 a_36128_2035# a_35707_2035# a_35392_2240# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2409 a_21911_6119# a_21698_6119# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2410 a_21979_5608# a_21558_5608# a_21041_5852# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2411 a_24011_4258# a_24264_4245# a_23069_4679# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2412 vdd d0 a_39354_1536# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2413 a_13854_1150# a_10153_1016# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2414 a_1792_7833# a_1371_7833# a_854_8077# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2415 a_29064_2270# a_29321_2080# a_28126_2514# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2416 a_26098_3687# a_25677_3687# a_25361_3568# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2417 a_5487_8667# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2418 a_1793_4524# a_1372_4524# a_854_4214# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2419 a_30336_2658# a_30336_2429# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2420 vdd d1 a_13169_8925# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2421 gnd d0 a_4078_5367# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2422 a_6851_1256# a_6783_1767# a_6861_2883# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2423 a_30333_8817# a_30334_8360# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2424 a_34042_8126# a_34295_8113# a_33103_7816# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2425 a_6738_387# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2426 gnd a_38414_2329# a_38206_2329# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2427 a_25361_2465# a_25361_2235# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2428 a_35392_3989# a_35392_3802# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2429 a_17971_3641# a_18958_3207# a_18909_3397# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2430 a_30334_7714# a_30862_7509# a_31070_7509# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2431 gnd a_23326_5592# a_23118_5592# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2432 a_35919_4241# a_35706_4241# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2433 vdd a_4079_3161# a_3871_3161# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2434 a_25239_307# a_29965_191# a_19317_134# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2435 vdd a_19166_2104# a_18958_2104# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2436 gnd d3 a_23215_7274# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2437 a_25889_5893# a_25676_5893# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2438 a_16897_3007# a_16783_2888# a_16890_5100# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2439 a_15734_3157# a_15521_3157# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2440 a_32008_8922# a_31941_8330# a_32025_7359# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2441 gnd d0 a_39351_4291# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2442 vdd d2 a_23186_3978# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2443 a_21981_1196# a_21560_1196# a_21042_886# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2444 a_3824_7586# a_3820_7763# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2445 a_20831_6401# a_20618_6401# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2446 vdd d2 a_38274_1818# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2447 a_15204_6901# a_15733_7020# a_15941_7020# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2448 vdd a_14109_8132# a_13901_8132# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2449 a_2889_1212# a_3873_1509# a_3828_1522# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2450 gnd d1 a_28381_7839# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2451 a_36857_6757# a_36644_6757# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2452 gnd d0 a_14111_2617# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2453 a_5488_7564# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2454 a_1794_3421# a_1373_3421# a_856_3665# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2455 a_35392_3802# a_35921_3692# a_36129_3692# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2456 a_5489_4255# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2457 a_29066_1721# a_29069_990# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2458 a_20618_9161# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2459 a_15204_7317# a_15204_7130# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2460 gnd a_29320_5389# a_29112_5389# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2461 vdd d1 a_13171_4513# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2462 vdd d1 a_8194_8961# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2463 a_31588_6716# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2464 a_16769_392# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2465 a_10680_1464# a_10467_1464# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2466 a_25360_5087# a_25888_5339# a_26096_5339# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2467 gnd a_23328_1180# a_23120_1180# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2468 a_34849_312# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2469 vdd a_3138_8920# a_2930_8920# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2470 gnd d3 a_23217_2862# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2471 a_24012_3155# a_24008_3332# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2472 a_12807_7311# a_12821_8414# a_12772_8604# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2473 a_6427_7874# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2474 a_1902_5054# a_1481_5054# a_1808_5173# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2475 a_20303_6836# a_20303_6606# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2476 a_24007_4435# a_24264_4245# a_23069_4679# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2477 a_25890_3687# a_25677_3687# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2478 a_21667_7235# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2479 a_35709_1486# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2480 vout a_18995_134# a_9987_210# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2481 gnd d1 a_23325_7798# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2482 a_17975_2361# a_18228_2348# a_17835_1850# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2483 a_34041_9229# a_34037_9406# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2484 a_12807_7311# a_13060_7298# a_12809_5099# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2485 gnd a_39354_1536# a_39146_1536# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2486 a_36859_2345# a_36646_2345# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2487 a_26097_5893# a_26827_5649# a_27035_5649# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2488 a_19317_134# a_29752_191# a_25239_307# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2489 a_34038_8303# a_34295_8113# a_33103_7816# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2490 a_32989_7469# a_33008_6189# a_32959_6379# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2491 gnd a_23186_3978# a_22978_3978# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2492 a_20305_3527# a_20834_3646# a_21042_3646# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2493 a_38158_8960# a_38411_8947# a_38018_8449# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2494 a_8881_7078# a_8877_7255# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2495 a_21771_4505# a_21558_4505# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2496 gnd a_9135_3202# a_8927_3202# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2497 a_26094_8648# a_26825_8958# a_27033_8958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2498 vdd d1 a_8196_4549# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2499 vdd d3 a_23215_7274# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2500 a_25364_1033# a_25890_927# a_26098_927# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2501 a_11405_1220# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2502 a_20305_2194# a_20833_1989# a_21041_1989# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2503 vdd d2 a_3000_3997# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2504 a_436_1459# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2505 a_27034_7855# a_26613_7855# a_26095_7545# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2506 vdd a_3140_4508# a_2932_4508# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2507 a_31070_6406# a_30649_6406# a_30335_6154# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2508 a_6429_3462# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2509 a_28128_7852# a_29112_8149# a_29063_8339# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2510 a_16670_8982# a_16457_8982# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2511 a_25362_1778# a_25362_1591# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2512 gnd d1 a_23327_3386# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2513 a_30337_1096# a_30339_997# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2514 a_11926_351# a_11713_351# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2515 a_15204_6671# a_15732_6466# a_15940_6466# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2516 a_26099_1481# a_26829_1237# a_27037_1237# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2517 a_9888_210# a_14663_331# a_14985_331# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2518 a_12809_2899# a_13062_2886# a_12805_5276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2519 a_22933_3991# a_23118_4489# a_23069_4679# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2520 a_36969_2869# a_36756_2869# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2521 a_35704_8653# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2522 a_30861_8612# a_30648_8612# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2523 vdd a_23328_1180# a_23120_1180# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2524 a_21978_7814# a_21910_8325# a_21994_7354# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2525 a_15734_4814# a_15521_4814# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2526 a_6537_5095# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2527 a_12807_7311# a_12821_8414# a_12776_8427# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2528 a_29067_4299# a_29320_4286# a_28125_4720# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2529 gnd d1 a_18226_7863# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2530 a_29063_8339# a_29066_7608# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2531 a_36786_3959# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2532 a_27986_2003# a_28243_1813# a_28016_3093# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2533 a_32960_4173# a_33150_3391# a_33105_3404# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2534 a_15939_8672# a_15518_8672# a_15204_8420# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2535 a_28018_7328# a_28032_8431# a_27983_8621# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2536 a_37175_5081# a_36754_5081# a_37081_5200# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2537 a_18915_1568# a_19168_1555# a_17976_1258# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2538 gnd d0 a_9134_5408# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2539 a_31071_5303# a_30650_5303# a_30335_5508# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2540 a_27036_3443# a_26615_3443# a_26097_3133# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2541 gnd d1 a_3139_7817# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2542 vdd a_39354_1536# a_39146_1536# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2543 vdd a_29322_977# a_29114_977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2544 a_17832_8468# a_18017_8966# a_17968_9156# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2545 gnd d0 a_24264_7005# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2546 a_10149_4883# a_10678_4773# a_10886_4773# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2547 gnd a_13170_7822# a_12962_7822# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2548 a_39098_8167# a_39351_8154# a_38159_7857# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2549 a_36643_8963# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2550 a_8876_7804# a_8881_7078# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2551 gnd a_4078_5367# a_3870_5367# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2552 a_15205_5111# a_15733_5363# a_15941_5363# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2553 a_17975_3464# a_18959_3761# a_18910_3951# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2554 a_33104_4507# a_33357_4494# a_32964_3996# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2555 a_1694_7254# a_1481_7254# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2556 a_2888_3418# a_3872_3715# a_3823_3905# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2557 a_35706_4241# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2558 a_15735_3711# a_15522_3711# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2559 a_30863_4200# a_30650_4200# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2560 a_15207_1386# a_15207_1156# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2561 a_20305_3297# a_20305_2840# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2562 a_6639_8977# a_6426_8977# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2563 gnd a_23215_7274# a_23007_7274# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2564 a_25676_5893# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2565 a_21040_5298# a_20619_5298# a_20304_5046# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2566 a_21980_3402# a_21912_3913# a_21996_2942# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2567 a_15521_3157# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2568 a_15940_7569# a_16671_7879# a_16879_7879# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2569 a_29064_6133# a_29067_5402# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2570 a_12809_2899# a_12823_4002# a_12778_4015# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2571 a_6850_3462# a_6429_3462# a_5912_3706# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2572 vdd a_38274_1818# a_38066_1818# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2573 a_37277_373# a_37168_373# a_35171_312# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2574 gnd d1 a_13170_6719# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2575 gnd d0 a_9136_996# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2576 vdd d1 a_23327_3386# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2577 a_31073_891# a_30652_891# a_30337_1096# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2578 a_23074_3399# a_24058_3696# a_24009_3886# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2579 a_39093_7790# a_39098_7064# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2580 a_18914_1014# a_18910_1191# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2581 a_36645_4551# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2582 a_15205_4695# a_15205_4465# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2583 vdd a_8194_8961# a_7986_8961# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2584 gnd a_4080_955# a_3872_955# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2585 a_16879_6776# a_16458_6776# a_15940_6466# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2586 a_37078_2869# a_36787_1753# a_37068_1242# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2587 a_117_8374# a_117_8187# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2588 vdd a_28381_7839# a_28173_7839# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2589 gnd d2 a_23187_1772# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2590 a_29063_4476# a_29320_4286# a_28125_4720# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2591 a_18911_1745# a_19168_1555# a_17976_1258# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2592 a_28018_7328# a_28032_8431# a_27987_8444# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2593 gnd a_14110_5926# a_13902_5926# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2594 a_21996_2942# a_21699_3913# a_21980_3402# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2595 a_25678_1481# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2596 a_10887_910# a_10466_910# a_10153_1016# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2597 gnd a_23217_2862# a_23009_2862# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2598 a_24008_4989# a_24265_4799# a_23073_4502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2599 a_15942_3157# a_16673_3467# a_16881_3467# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2600 a_10466_910# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2601 a_25140_307# a_25031_307# a_25239_307# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2602 a_39094_8344# a_39351_8154# a_38159_7857# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2603 a_21039_6401# a_21770_6711# a_21978_6711# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2604 gnd a_23325_7798# a_23117_7798# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2605 a_35918_6447# a_35705_6447# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2606 gnd d1 a_8195_6755# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2607 a_34044_3714# a_34297_3701# a_33105_3404# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2608 gnd d0 a_39350_6497# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2609 a_17975_3464# a_18959_3761# a_18914_3774# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2610 a_12775_1986# a_12965_1204# a_12916_1394# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2611 a_31073_2548# a_30652_2548# a_30336_2658# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2612 a_20830_8607# a_20617_8607# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2613 a_13851_7768# a_13856_7042# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2614 a_30649_6406# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2615 vdd a_24266_936# a_24058_936# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2616 a_6951_387# a_6738_387# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2617 gnd a_3139_6714# a_2931_6714# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2618 vdd a_8196_4549# a_7988_4549# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2619 a_2888_3418# a_3872_3715# a_3827_3728# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2620 a_10885_8082# a_10464_8082# a_10148_8192# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2621 a_118_4419# a_119_3962# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2622 a_25362_1362# a_25891_1481# a_26099_1481# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2623 a_17831_2027# a_18088_1837# a_17861_3117# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2624 vdd a_23215_7274# a_23007_7274# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2625 a_1793_5627# a_1372_5627# a_855_5871# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2626 a_35391_6008# a_35920_5898# a_36128_5898# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2627 a_32320_332# a_31899_332# a_32119_5040# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2628 a_24012_2052# a_24265_2039# a_23070_2473# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2629 a_1794_2318# a_1373_2318# a_855_2008# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2630 a_10884_9185# a_11614_8941# a_11822_8941# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2631 a_11543_6143# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2632 a_28020_2916# a_28034_4019# a_27989_4032# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2633 a_22927_8580# a_23117_7798# a_23072_7811# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2634 a_30864_4754# a_30651_4754# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2635 a_31911_5040# a_31698_5040# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2636 a_12779_1809# a_13032_1796# a_12805_3076# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2637 a_35390_7985# a_35390_7755# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2638 a_39096_2829# a_39099_2098# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2639 a_32991_5257# a_33040_2867# a_32995_2880# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2640 vdd a_29321_5943# a_29113_5943# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2641 gnd a_23327_3386# a_23119_3386# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2642 a_10149_5527# a_10149_5070# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2643 gnd d1 a_8197_2343# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2644 a_27034_7855# a_26966_8366# a_27050_7395# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2645 gnd d3 a_3029_7293# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2646 a_32009_6716# a_31942_6124# a_32020_7240# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2647 gnd d0 a_39352_2085# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2648 a_20832_4195# a_20619_4195# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2649 vdd d2 a_23187_1772# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2650 a_36756_2869# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2651 a_26095_9202# a_25674_9202# a_25358_9083# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2652 a_15521_4814# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2653 a_34042_4263# a_34038_4440# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2654 a_32012_1201# a_31944_1712# a_32022_2828# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2655 a_10150_2677# a_10150_2448# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2656 a_5489_5358# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2657 a_35393_1596# a_35922_1486# a_36130_1486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2658 a_7800_2022# a_7990_1240# a_7941_1430# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2659 a_1795_1215# a_1374_1215# a_857_1459# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2660 gnd a_18226_7863# a_18018_7863# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2661 a_118_5981# a_118_5752# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2662 a_29063_5579# a_29068_4853# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2663 a_18995_134# d8 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2664 a_8882_2112# a_8878_2289# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2665 a_20619_6955# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2666 a_20306_1091# a_20308_992# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2667 gnd a_9134_5408# a_8926_5408# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2668 vdd d1 a_8195_6755# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2669 vdd d2 a_18086_6249# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2670 a_3826_5934# a_3822_6111# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2671 a_31589_4510# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2672 a_27983_8621# a_28173_7839# a_28124_8029# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2673 gnd a_24264_7005# a_24056_7005# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2674 a_13857_4836# a_14110_4823# a_12918_4526# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2675 a_5702_8118# a_5489_8118# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2676 a_6750_7295# a_6537_7295# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2677 vdd d2 a_2999_6203# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2678 a_16895_5219# a_16781_5100# a_16989_5100# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2679 a_13854_2807# a_13857_2076# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2680 vdd a_3139_6714# a_2931_6714# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2681 a_10149_5527# a_10677_5322# a_10885_5322# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2682 a_27036_3443# a_26968_3954# a_27052_2983# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2683 gnd d3 a_3031_2881# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2684 vdd a_13030_6208# a_12822_6208# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2685 a_6428_5668# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2686 a_21991_2823# a_21882_2823# a_21989_5035# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2687 a_1481_7254# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2688 a_645_6420# a_432_6420# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2689 a_117_8187# a_646_8077# a_854_8077# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2690 a_21041_5852# a_20620_5852# a_20304_5733# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2691 a_15522_3711# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2692 a_30650_4200# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2693 a_6426_8977# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2694 a_31072_1994# a_30651_1994# a_30337_1742# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2695 a_5910_4255# a_5489_4255# a_5175_4003# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2696 a_12912_9115# a_13899_8681# a_13850_8871# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2697 a_20306_1321# a_20835_1440# a_21043_1440# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2698 a_34043_5920# a_34039_6097# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2699 gnd d0 a_9137_1550# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2700 a_35392_2886# a_35392_2699# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2701 a_3827_3728# a_3823_3905# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2702 gnd a_9136_996# a_8928_996# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2703 a_21772_2299# a_21559_2299# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2704 vdd a_23327_3386# a_23119_3386# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2705 vdd d1 a_8197_2343# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2706 a_5178_1052# a_5704_946# a_5912_946# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2707 vdd d0 a_39352_2085# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2708 a_3824_6483# a_3820_6660# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2709 a_12809_5099# a_12852_7298# a_12803_7488# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2710 a_8879_1186# a_5178_1052# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2711 a_31070_7509# a_30649_7509# a_30334_7714# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2712 a_27035_5649# a_26614_5649# a_26096_5339# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2713 a_36128_4795# a_35707_4795# a_35391_4905# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2714 vdd a_3141_2302# a_2933_2302# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2715 a_29064_5030# a_29321_4840# a_28129_4543# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2716 a_2885_8933# a_3138_8920# a_2745_8422# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2717 a_10148_7089# a_10677_6979# a_10885_6979# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2718 a_15205_5798# a_15734_5917# a_15942_5917# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2719 a_27033_8958# a_26612_8958# a_26095_9202# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2720 a_39093_9447# a_39096_8716# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2721 a_7800_2022# a_7990_1240# a_7945_1253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2722 vdd d0 a_9135_5962# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2723 a_25360_5774# a_25360_5544# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2724 gnd d1 a_3141_3405# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2725 a_21043_1440# a_20622_1440# a_20306_1321# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2726 a_15204_7317# a_15732_7569# a_15940_7569# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2727 vdd d3 a_38304_2908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2728 a_5911_3152# a_5490_3152# a_5175_3357# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2729 a_5176_1797# a_5176_1610# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2730 vdd a_4079_5921# a_3871_5921# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2731 a_35705_6447# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2732 a_30862_6406# a_30649_6406# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2733 a_18908_5603# a_18913_4877# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2734 a_32011_2304# a_31590_2304# a_31073_2548# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2735 gnd a_8195_6755# a_7987_6755# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2736 a_2884_2492# a_3871_2058# a_3826_2071# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2737 a_1792_7833# a_1724_8344# a_1808_7373# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2738 a_21979_5608# a_21911_6119# a_21989_7235# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2739 a_15735_2608# a_15522_2608# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2740 a_9987_210# a_9566_210# a_5053_326# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2741 a_24012_2052# a_24008_2229# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2742 a_9566_210# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2743 a_6850_2359# a_6429_2359# a_5911_2049# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2744 a_28014_7505# a_28033_6225# a_27984_6415# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2745 a_12805_5276# a_12854_2886# a_12805_3076# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2746 a_27037_1237# a_26616_1237# a_26098_927# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2747 a_31072_3097# a_30651_3097# a_30336_3302# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2748 a_12917_6732# a_13901_7029# a_13856_7042# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2749 a_855_5871# a_434_5871# a_118_5752# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2750 a_10149_5757# a_10678_5876# a_10886_5876# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2751 a_10150_2677# a_10679_2567# a_10887_2567# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2752 a_11615_6735# a_11402_6735# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2753 a_39099_5961# a_39352_5948# a_38160_5651# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2754 a_12912_9115# a_13899_8681# a_13854_8694# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2755 a_36644_6757# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2756 vdd d0 a_9137_1550# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2757 a_30651_4754# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2758 a_37083_2988# a_36786_3959# a_37067_3448# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2759 a_16781_7300# a_16568_7300# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2760 a_20304_6149# a_20831_6401# a_21039_6401# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2761 a_36967_5081# a_36754_5081# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2762 a_33105_2301# a_33358_2288# a_32965_1790# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2763 a_38155_6931# a_39142_6497# a_39097_6510# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2764 a_30863_5303# a_30650_5303# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2765 vdd a_4081_1509# a_3873_1509# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2766 a_35707_2035# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2767 a_10886_4773# a_10465_4773# a_10149_4654# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2768 a_15736_1505# a_15523_1505# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2769 gnd a_8197_2343# a_7989_2343# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2770 a_24010_9224# a_24006_9401# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2771 a_1794_3421# a_1726_3932# a_1810_2961# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2772 gnd d0 a_4081_1509# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2773 a_25677_3687# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2774 a_6851_1256# a_6430_1256# a_5913_1500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2775 gnd a_39352_2085# a_39144_2085# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2776 a_34041_9229# a_35389_9317# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2777 a_38019_6243# a_38272_6230# a_38045_7510# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2778 a_24013_3709# a_24009_3886# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2779 a_28016_3093# a_28035_1813# a_27986_2003# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2780 a_10151_1345# a_10680_1464# a_10888_1464# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2781 gnd d2 a_18085_8455# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2782 a_36645_5654# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2783 a_11617_2323# a_11404_2323# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2784 a_31802_5613# a_31589_5613# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2785 a_648_2562# a_435_2562# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2786 a_36646_2345# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2787 a_16879_7879# a_16458_7879# a_15941_8123# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2788 vdd a_8195_6755# a_7987_6755# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2789 a_30335_6154# a_30335_5967# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2790 a_31800_8922# a_31587_8922# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2791 gnd a_13029_8414# a_12821_8414# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2792 gnd d4 a_28273_5103# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2793 a_25361_3568# a_25890_3687# a_26098_3687# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2794 a_20303_7252# a_20303_7065# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2795 gnd d2 a_3001_1791# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2796 a_5175_2713# a_5704_2603# a_5912_2603# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2797 a_27047_2864# a_26938_2864# a_27045_5076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2798 a_16783_2888# a_16570_2888# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2799 a_30865_891# a_30652_891# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2800 a_11542_8349# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2801 a_28014_7505# a_28033_6225# a_27988_6238# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2802 a_28127_1411# a_29114_977# a_29069_990# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2803 a_21991_2823# a_21700_1707# a_21981_1196# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2804 a_20306_1737# a_20306_1550# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2805 a_24009_2783# a_24266_2593# a_23074_2296# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2806 a_28016_5293# a_28065_2903# a_28016_3093# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2807 a_23071_8914# a_24055_9211# a_24006_9401# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2808 a_432_6420# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2809 a_21040_4195# a_21771_4505# a_21979_4505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2810 a_28129_4543# a_28382_4530# a_27989_4032# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2811 a_15731_8672# a_15518_8672# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2812 a_8876_6701# a_8882_5975# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2813 gnd d1 a_8196_4549# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2814 gnd d2 a_18087_4043# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2815 a_34045_1508# a_34298_1495# a_33106_1198# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2816 a_21912_3913# a_21699_3913# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2817 a_31804_1201# a_31591_1201# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2818 a_36647_1242# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2819 a_16982_392# a_16769_392# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2820 gnd a_9137_1550# a_8929_1550# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2821 a_32962_8408# a_33147_8906# a_33098_9096# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2822 a_16813_3978# a_16600_3978# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2823 a_20305_2194# a_20306_1737# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2824 a_18913_2117# a_19166_2104# a_17971_2538# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2825 a_3821_8317# a_4078_8127# a_2886_7830# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2826 a_20304_5046# a_20304_4859# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2827 a_37168_373# a_36955_373# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2828 vdd d0 a_39353_2639# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2829 vdd a_8197_2343# a_7989_2343# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2830 a_11727_2847# a_11514_2847# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2831 a_21978_6711# a_21557_6711# a_21040_6955# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2832 a_15939_8672# a_16670_8982# a_16878_8982# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2833 a_26097_4790# a_25676_4790# a_25360_4671# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2834 vdd a_39352_2085# a_39144_2085# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2835 a_28123_9132# a_28380_8942# a_27987_8444# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2836 gnd d0 a_4077_6470# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2837 a_10885_6979# a_11615_6735# a_11823_6735# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2838 a_38015_6420# a_38272_6230# a_38045_7510# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2839 a_11544_3937# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2840 a_22289_327# a_21868_327# a_22190_327# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2841 a_22928_6374# a_23118_5592# a_23073_5605# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2842 a_3827_968# a_3823_1145# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2843 a_30865_2548# a_30652_2548# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2844 vdd d2 a_18085_8455# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2845 a_30333_8817# a_30861_8612# a_31069_8612# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2846 a_39093_6687# a_39099_5961# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2847 vdd a_9135_5962# a_8927_5962# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2848 a_29063_5579# a_29320_5389# a_28125_5823# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2849 a_10148_7733# a_10676_7528# a_10884_7528# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2850 vdd a_38304_2908# a_38096_2908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2851 a_27035_5649# a_26967_6160# a_27045_7276# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2852 a_2883_4698# a_3870_4264# a_3821_4454# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2853 a_2774_3071# a_2793_1791# a_2748_1804# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2854 a_30336_3302# a_30336_2845# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2855 vdd a_13029_8414# a_12821_8414# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2856 a_644_8626# a_431_8626# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2857 a_20833_1989# a_20620_1989# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2858 vdd d0 a_24264_8108# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2859 a_12916_8938# a_13900_9235# a_13851_9425# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2860 gnd d1 a_28380_8942# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2861 a_12805_3076# a_12824_1796# a_12775_1986# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2862 a_29069_2647# a_29322_2634# a_28130_2337# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2863 a_15522_2608# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2864 a_16671_6776# a_16458_6776# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2865 gnd d0 a_34296_5907# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2866 a_23071_8914# a_24055_9211# a_24010_9224# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2867 gnd a_28271_7315# a_28063_7315# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2868 a_10885_5322# a_11616_5632# a_11824_5632# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2869 gnd d0 a_9136_3756# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2870 gnd a_29319_6492# a_29111_6492# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2871 a_5912_946# a_5491_946# a_5178_1052# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2872 a_10887_2567# a_11617_2323# a_11825_2323# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2873 a_33100_5787# a_33357_5597# a_32959_6379# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2874 a_28125_4720# a_28382_4530# a_27989_4032# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2875 a_6569_3973# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2876 a_5491_946# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2877 a_25887_9202# a_25674_9202# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2878 a_11402_6735# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2879 a_25360_6190# a_25887_6442# a_26095_6442# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2880 vdd d2 a_18087_4043# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2881 a_23071_1370# a_24058_936# a_24013_949# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2882 gnd a_4080_3715# a_3872_3715# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2883 a_30335_4405# a_30863_4200# a_31071_4200# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2884 vdd a_9137_1550# a_8929_1550# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2885 a_13851_6665# a_13857_5939# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2886 a_10150_3321# a_10678_3116# a_10886_3116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2887 a_36754_5081# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2888 vdd a_13031_4002# a_12823_4002# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2889 a_1805_2842# a_1696_2842# a_1803_5054# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2890 a_645_7523# a_432_7523# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2891 a_35390_7111# a_35919_7001# a_36127_7001# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2892 a_26097_5893# a_25676_5893# a_25360_6003# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2893 a_30650_5303# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2894 a_646_4214# a_433_4214# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2895 a_21042_3646# a_20621_3646# a_20305_3527# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2896 a_15523_1505# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2897 a_29066_9265# a_29062_9442# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2898 vdd d0 a_4077_6470# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2899 a_12918_4526# a_13902_4823# a_13853_5013# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2900 a_5910_5358# a_5489_5358# a_5174_5563# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2901 a_26096_6996# a_26826_6752# a_27034_6752# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2902 a_8878_6152# a_8881_5421# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2903 a_16989_5100# a_16568_5100# a_16890_5100# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2904 a_5911_2049# a_5490_2049# a_5176_1797# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2905 a_16673_2364# a_16460_2364# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2906 a_21040_6955# a_20619_6955# a_20303_7065# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2907 a_10885_5322# a_10464_5322# a_10149_5070# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2908 a_17861_3117# a_18118_2927# a_17861_5317# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2909 a_26924_368# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2910 gnd a_29321_2080# a_29113_2080# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2911 a_32010_4510# a_31589_4510# a_31072_4754# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2912 a_2883_4698# a_3870_4264# a_3825_4277# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2913 a_10149_4424# a_10150_3967# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2914 a_117_7728# a_117_7271# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2915 a_11404_2323# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2916 a_15941_8123# a_15520_8123# a_15204_8004# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2917 a_30864_1994# a_30651_1994# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2918 a_435_2562# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2919 gnd d0 a_29318_8698# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2920 a_10148_8192# a_10148_7963# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2921 a_31073_891# a_30652_891# a_30339_997# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2922 a_36129_2589# a_35708_2589# a_35392_2699# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2923 a_12916_8938# a_13900_9235# a_13855_9248# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2924 gnd a_28273_5103# a_28065_5103# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2925 a_29065_2824# a_29322_2634# a_28130_2337# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2926 a_22088_5035# a_21667_5035# a_21989_5035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2927 a_647_3111# a_434_3111# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2928 a_16570_2888# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2929 a_28127_8955# a_29111_9252# a_29062_9442# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2930 a_35920_4795# a_35707_4795# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2931 a_30652_891# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2932 vdd d0 a_39350_7600# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2933 vdd a_28271_7315# a_28063_7315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2934 a_32020_7240# a_31729_6124# a_32009_6716# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2935 a_118_4878# a_118_4649# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2936 a_29063_4476# a_29069_3750# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2937 vdd d0 a_9136_3756# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2938 gnd d1 a_3142_1199# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2939 a_853_9180# a_1583_8936# a_1791_8936# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2940 a_34042_7023# a_34038_7200# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2941 a_5912_946# a_5491_946# a_5176_1151# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2942 a_26098_2584# a_26828_2340# a_27036_2340# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2943 a_20303_8355# a_20830_8607# a_21038_8607# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2944 a_36860_1242# a_36647_1242# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2945 a_11758_1731# a_11545_1731# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2946 a_38154_9137# a_39141_8703# a_39096_8716# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2947 a_30862_7509# a_30649_7509# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2948 vdd a_4080_3715# a_3872_3715# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2949 a_36787_1753# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2950 a_8877_8358# a_9134_8168# a_7942_7871# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2951 a_10885_6979# a_10464_6979# a_10148_6860# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2952 gnd a_8196_4549# a_7988_4549# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2953 a_1793_5627# a_1725_6138# a_1803_7254# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2954 a_38047_5298# a_38096_2908# a_38051_2921# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2955 a_20619_4195# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2956 a_34041_7572# a_34037_7749# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2957 a_10149_5986# a_10149_5757# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2958 a_31591_1201# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2959 a_38018_8449# a_38271_8436# a_38049_7333# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2960 a_21994_5154# a_21667_7235# a_21994_7354# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2961 a_16600_3978# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2962 a_8881_5421# a_8877_5598# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2963 a_28020_2916# a_28034_4019# a_27985_4209# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2964 a_11514_2847# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2965 a_32025_5159# a_31911_5040# a_32119_5040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2966 a_10150_3551# a_10679_3670# a_10887_3670# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2967 vdd a_39353_2639# a_39145_2639# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2968 a_3827_2625# a_4080_2612# a_2888_2315# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2969 a_11839_7378# a_11725_7259# a_11839_5178# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2970 a_856_3665# a_435_3665# a_119_3546# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2971 a_35390_8401# a_35390_8214# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2972 a_36644_7860# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2973 a_28129_4543# a_29113_4840# a_29064_5030# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2974 a_11616_4529# a_11403_4529# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2975 a_31801_7819# a_31588_7819# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2976 a_5174_6209# a_5174_6022# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2977 a_647_4768# a_434_4768# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2978 a_1808_7373# a_1511_8344# a_1791_8936# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2979 a_854_6974# a_433_6974# a_117_7084# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2980 gnd a_4077_6470# a_3869_6470# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2981 a_34043_4817# a_34039_4994# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2982 vdd a_29321_2080# a_29113_2080# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2983 vdd d0 a_39352_3188# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2984 a_18912_8186# a_18908_8363# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2985 vdd a_4080_955# a_3872_955# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2986 a_30652_2548# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2987 a_13853_6116# a_13856_5385# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2988 a_20305_3943# a_20832_4195# a_21040_4195# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2989 a_38156_4725# a_39143_4291# a_39098_4304# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2990 a_30864_3097# a_30651_3097# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2991 vdd d0 a_29320_8149# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2992 a_10886_5876# a_10465_5876# a_10149_5986# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2993 a_3826_5934# a_4079_5921# a_2887_5624# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2994 a_10887_2567# a_10466_2567# a_10150_2448# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2995 a_39100_3755# a_39096_3932# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2996 a_431_8626# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2997 a_20620_1989# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2998 a_28127_8955# a_29111_9252# a_29066_9265# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2999 vdd a_24264_8108# a_24056_8108# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3000 a_35920_5898# a_35707_5898# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3001 a_38020_4037# a_38273_4024# a_38051_2921# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3002 a_13858_973# a_14111_960# a_12916_1394# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3003 a_28128_6749# a_28381_6736# a_27988_6238# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3004 a_39097_6510# a_39093_6687# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3005 a_38156_5828# a_38413_5638# a_38015_6420# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3006 a_36999_3959# a_36786_3959# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3007 a_21039_6401# a_20618_6401# a_20303_6606# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3008 a_5173_8228# a_5702_8118# a_5910_8118# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3009 gnd d2 a_18086_6249# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3010 a_6864_7414# a_6750_7295# a_6864_5214# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3011 gnd a_34296_5907# a_34088_5907# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3012 a_5175_4003# a_5175_3816# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3013 a_36646_3448# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3014 gnd a_9136_3756# a_8928_3756# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3015 a_21559_2299# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3016 a_31803_3407# a_31590_3407# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3017 a_1810_2961# a_1513_3932# a_1793_4524# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3018 a_17091_392# a_17910_5127# a_17865_5140# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3019 a_18908_4500# a_18914_3774# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3020 vdd a_14111_960# a_13903_960# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3021 a_15206_3362# a_15734_3157# a_15942_3157# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3022 vdd d0 a_39352_4845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3023 a_5175_3587# a_5704_3706# a_5912_3706# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3024 a_25674_9202# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3025 a_10148_6860# a_10148_6630# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3026 a_26096_6996# a_25675_6996# a_25359_6877# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3027 a_10888_1464# a_10467_1464# a_10151_1574# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3028 a_18910_2848# a_19167_2658# a_17975_2361# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3029 gnd d0 a_4076_8676# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3030 a_38014_8626# a_38271_8436# a_38049_7333# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3031 a_29065_3927# a_29068_3196# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3032 a_13855_9248# a_15203_9336# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3033 a_432_7523# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3034 a_36127_8104# a_36857_7860# a_37065_7860# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3035 a_13858_3733# a_13854_3910# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3036 a_3823_2802# a_4080_2612# a_2888_2315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3037 a_39093_9447# a_39350_9257# a_38158_8960# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3038 a_12776_8427# a_12961_8925# a_12912_9115# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3039 a_433_4214# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3040 a_21041_1989# a_21772_2299# a_21980_2299# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3041 a_28130_2337# a_28383_2324# a_27990_1826# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3042 vdd a_4077_6470# a_3869_6470# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3043 a_13855_6488# a_13851_6665# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3044 a_5912_2603# a_5491_2603# a_5175_2484# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3045 a_15732_6466# a_15519_6466# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3046 gnd d2 a_18088_1837# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3047 a_12913_8012# a_13900_7578# a_13855_7591# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3048 a_16460_2364# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3049 gnd a_13060_7298# a_12852_7298# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3050 a_24011_5361# a_24007_5538# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3051 a_21913_1707# a_21700_1707# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3052 a_2887_4521# a_3871_4818# a_3826_4831# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3053 a_35393_1367# a_35393_1137# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3054 gnd a_38411_8947# a_38203_8947# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3055 a_21979_4505# a_21558_4505# a_21041_4749# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3056 a_10676_9185# a_10463_9185# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3057 a_17829_6439# a_18019_5657# a_17974_5670# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3058 a_30651_1994# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3059 a_26098_2584# a_25677_2584# a_25361_2465# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3060 a_10884_7528# a_11615_7838# a_11823_7838# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3061 a_25360_6190# a_25360_6003# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3062 gnd a_29318_8698# a_29110_8698# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3063 a_31911_7240# a_31698_7240# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3064 gnd d0 a_4078_4264# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3065 a_10886_4773# a_11616_4529# a_11824_4529# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3066 a_38016_4214# a_38273_4024# a_38051_2921# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3067 a_33099_7993# a_33356_7803# a_32958_8585# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3068 a_28124_6926# a_28381_6736# a_27988_6238# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3069 a_6568_6179# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3070 a_24013_2606# a_24009_2783# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3071 a_25359_8396# a_25886_8648# a_26094_8648# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3072 a_34042_7023# a_34295_7010# a_33103_6713# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3073 a_434_3111# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3074 a_17971_2538# a_18958_2104# a_18909_2294# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3075 gnd d0 a_14108_9235# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3076 a_30334_6611# a_30862_6406# a_31070_6406# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3077 vdd a_9136_3756# a_8928_3756# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3078 gnd a_3142_1199# a_2934_1199# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3079 vdd a_4079_2058# a_3871_2058# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3080 a_16878_8982# a_16457_8982# a_15940_9226# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3081 a_25889_4790# a_25676_4790# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3082 a_29070_1544# a_29066_1721# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3083 a_15734_2054# a_15521_2054# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3084 a_2884_2492# a_3871_2058# a_3822_2248# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3085 a_38049_7333# a_38302_7320# a_38051_5121# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3086 a_35707_4795# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3087 a_35389_9317# a_35918_9207# a_36126_9207# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3088 gnd d2 a_33215_8395# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3089 a_26096_8099# a_25675_8099# a_25359_8209# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3090 a_11823_6735# a_11756_6143# a_11834_7259# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3091 a_15206_3821# a_15206_3592# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3092 vdd a_14109_7029# a_13901_7029# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3093 vdd d0 a_4076_8676# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3094 a_12917_6732# a_13901_7029# a_13852_7219# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3095 a_29067_4299# a_29063_4476# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3096 a_37081_5200# a_36967_5081# a_37175_5081# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3097 a_35062_312# a_34849_312# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3098 a_26095_9202# a_26825_8958# a_27033_8958# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3099 a_5488_6461# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3100 a_16672_4570# a_16459_4570# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3101 a_25361_3984# a_25361_3797# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3102 a_10884_7528# a_10463_7528# a_10148_7276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3103 a_23072_6708# a_24056_7005# a_24011_7018# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3104 a_10886_3116# a_11617_3426# a_11825_3426# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3105 gnd a_8085_7334# a_7877_7334# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3106 gnd a_29320_4286# a_29112_4286# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3107 a_28126_2514# a_28383_2324# a_27990_1826# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3108 a_33101_3581# a_33358_3391# a_32960_4173# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3109 a_27987_8444# a_28172_8942# a_28123_9132# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3110 a_16890_7300# a_16781_7300# a_16895_5219# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3111 a_25361_3984# a_25888_4236# a_26096_4236# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3112 a_18910_3951# a_18913_3220# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3113 a_6859_5095# a_6539_2883# a_6866_3002# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3114 a_5701_9221# a_5488_9221# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3115 a_33104_5610# a_34088_5907# a_34039_6097# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3116 a_30335_5051# a_30863_5303# a_31071_5303# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3117 a_11403_4529# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3118 a_434_4768# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3119 a_5175_3587# a_5175_3357# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3120 vdd a_39352_3188# a_39144_3188# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3121 gnd a_39351_8154# a_39143_8154# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3122 a_1682_346# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3123 a_8882_5975# a_9135_5962# a_7943_5665# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3124 a_4954_326# a_4845_326# a_5053_326# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3125 a_6427_6771# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3126 a_25890_2584# a_25677_2584# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3127 a_35390_7985# a_35919_8104# a_36127_8104# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3128 a_646_5317# a_433_5317# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3129 a_116_9290# a_645_9180# a_853_9180# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3130 gnd d2 a_33217_3983# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3131 a_647_2008# a_434_2008# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3132 a_30651_3097# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3133 gnd d1 a_23325_6695# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3134 vdd d0 a_4078_4264# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3135 a_26095_7545# a_26826_7855# a_27034_7855# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3136 a_18907_7809# a_19164_7619# a_17969_8053# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3137 a_31072_5857# a_31802_5613# a_32010_5613# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3138 a_26097_4790# a_26827_4546# a_27035_4546# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3139 a_34038_7200# a_34295_7010# a_33103_6713# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3140 a_20305_2424# a_20834_2543# a_21042_2543# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3141 a_6866_3002# a_6569_3973# a_6849_4565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3142 a_10886_3116# a_10465_3116# a_10150_2864# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3143 gnd a_8087_2922# a_7879_2922# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3144 vdd d0 a_14108_9235# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3145 a_1803_5054# a_1483_2842# a_1810_2961# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3146 a_36786_3959# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3147 a_31069_8612# a_31800_8922# a_32008_8922# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3148 a_16892_2888# a_16783_2888# a_16890_5100# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3149 a_38045_7510# a_38302_7320# a_38051_5121# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3150 a_25889_5893# a_25676_5893# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3151 a_30335_5508# a_30335_5051# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3152 a_30336_2199# a_30337_1742# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3153 gnd d0 a_29321_5943# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3154 a_31590_3407# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3155 a_15206_3821# a_15735_3711# a_15943_3711# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3156 a_15735_951# a_15522_951# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3157 a_31941_8330# a_31728_8330# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3158 a_27034_6752# a_26613_6752# a_26095_6442# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3159 vdd a_39352_4845# a_39144_4845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3160 a_648_905# a_435_905# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3161 a_28128_6749# a_29112_7046# a_29063_7236# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3162 a_35921_2589# a_35708_2589# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3163 a_32027_2947# a_31730_3918# a_32010_4510# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3164 gnd d1 a_23327_2283# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3165 a_853_9180# a_432_9180# a_116_9290# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3166 gnd a_4076_8676# a_3868_8676# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3167 a_15204_8420# a_15731_8672# a_15939_8672# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3168 vdd a_8085_7334# a_7877_7334# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3169 vdd d0 a_39351_5394# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3170 vdd a_29320_4286# a_29112_4286# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3171 a_38161_3445# a_38414_3432# a_38016_4214# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3172 a_26095_7545# a_25674_7545# a_25359_7293# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3173 a_26097_3133# a_26828_3443# a_27036_3443# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3174 a_6639_8977# a_6426_8977# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3175 a_18909_3397# a_19166_3207# a_17971_3641# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3176 a_21979_4505# a_21912_3913# a_21996_2942# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3177 a_16881_3467# a_16813_3978# a_16897_3007# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3178 a_3828_1522# a_3824_1699# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3179 a_3825_8140# a_4078_8127# a_2886_7830# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3180 vdd a_39351_8154# a_39143_8154# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3181 gnd d0 a_39353_2639# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3182 a_22960_5252# a_23009_2862# a_22964_2875# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3183 a_32965_1790# a_33150_2288# a_33105_2301# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3184 a_21700_1707# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3185 a_13857_3179# a_14110_3166# a_12915_3600# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3186 a_38155_8034# a_38412_7844# a_38014_8626# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3187 gnd d0 a_9134_4305# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3188 a_27036_2340# a_26615_2340# a_26097_2030# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3189 a_21038_8607# a_20617_8607# a_20302_8812# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3190 vdd d2 a_8057_1832# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3191 a_10463_9185# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3192 a_20832_8058# a_20619_8058# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3193 a_857_1459# a_436_1459# a_120_1340# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3194 a_20305_3527# a_20305_3297# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3195 a_39098_7064# a_39351_7051# a_38159_6754# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3196 a_8878_5049# a_8881_4318# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3197 a_7942_7871# a_8926_8168# a_8881_8181# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3198 a_1803_7254# a_1512_6138# a_1792_6730# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3199 gnd a_4078_4264# a_3870_4264# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3200 a_6539_2883# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3201 a_35390_7755# a_35918_7550# a_36126_7550# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3202 a_39097_1726# a_39100_995# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3203 a_26097_3133# a_25676_3133# a_25361_2881# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3204 a_12914_5806# a_13901_5372# a_13852_5562# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3205 a_20306_1737# a_20833_1989# a_21041_1989# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3206 gnd a_14108_9235# a_13900_9235# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3207 a_11839_5178# a_11512_7259# a_11834_7259# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3208 a_117_6625# a_118_6168# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3209 a_18909_5054# a_19166_4864# a_17974_4567# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3210 a_10887_3670# a_10466_3670# a_10150_3780# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3211 a_12919_2320# a_13172_2307# a_12779_1809# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3212 a_2888_2315# a_3872_2612# a_3823_2802# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3213 a_23069_5782# a_24056_5348# a_24011_5361# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3214 a_32991_3057# a_33248_2867# a_32991_5257# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3215 a_15940_6466# a_16671_6776# a_16879_6776# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3216 a_25676_4790# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3217 a_21040_4195# a_20619_4195# a_20305_3943# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3218 a_15521_2054# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3219 a_10147_9066# a_10676_9185# a_10884_9185# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3220 gnd d0 a_24267_1490# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3221 gnd a_33215_8395# a_33007_8395# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3222 a_28128_6749# a_29112_7046# a_29067_7059# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3223 vdd d4 a_18118_5127# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3224 a_38021_1831# a_38274_1818# a_38047_3098# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3225 vdd d1 a_23327_2283# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3226 vdd a_4076_8676# a_3868_8676# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3227 a_5911_4809# a_5490_4809# a_5174_4690# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3228 a_38157_3622# a_38414_3432# a_38016_4214# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3229 a_23074_2296# a_24058_2593# a_24009_2783# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3230 a_10148_7733# a_10148_7276# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3231 a_22081_327# a_21868_327# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3232 gnd d0 a_4079_4818# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3233 a_12916_1394# a_13903_960# a_13854_1150# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3234 a_5176_1381# a_5705_1500# a_5913_1500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3235 a_17828_8645# a_18018_7863# a_17973_7876# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3236 a_10149_4883# a_10149_4654# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3237 gnd a_14110_4823# a_13902_4823# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3238 a_13853_3356# a_14110_3166# a_12915_3600# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3239 a_21557_7814# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3240 a_29062_7785# a_29067_7059# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3241 a_6864_5214# a_6537_7295# a_6859_7295# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3242 vdd d0 a_14108_7578# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3243 a_15942_2054# a_16673_2364# a_16881_2364# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3244 a_34041_9229# a_34294_9216# a_33102_8919# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3245 a_39094_7241# a_39351_7051# a_38159_6754# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3246 a_433_5317# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3247 a_36128_5898# a_36858_5654# a_37066_5654# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3248 a_3825_8140# a_3821_8317# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3249 a_35390_7298# a_35390_7111# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3250 gnd a_23325_6695# a_23117_6695# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3251 gnd a_33217_3983# a_33009_3983# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3252 a_434_2008# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3253 a_5174_5106# a_5174_4919# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3254 a_5912_3706# a_5491_3706# a_5175_3816# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3255 a_36125_8653# a_36856_8963# a_37064_8963# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3256 vdd a_4078_4264# a_3870_4264# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3257 a_25888_6996# a_25675_6996# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3258 a_15733_4260# a_15520_4260# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3259 a_16814_1772# a_16601_1772# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3260 a_13853_5013# a_13856_4282# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3261 a_21980_2299# a_21559_2299# a_21041_1989# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3262 a_17975_2361# a_18959_2658# a_18914_2671# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3263 a_12914_5806# a_13901_5372# a_13856_5385# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3264 a_11822_8941# a_11755_8349# a_11839_7378# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3265 vdd a_14108_9235# a_13900_9235# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3266 a_2888_2315# a_3872_2612# a_3827_2625# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3267 a_20619_6955# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3268 a_25676_5893# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3269 a_11545_1731# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3270 a_39100_2652# a_39096_2829# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3271 a_5487_8667# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3272 a_27050_5195# a_26723_7276# a_27045_7276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3273 a_1793_4524# a_1372_4524# a_855_4768# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3274 a_35391_4905# a_35920_4795# a_36128_4795# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3275 a_20834_886# a_20621_886# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3276 a_21559_3402# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3277 a_18912_5426# a_19165_5413# a_17970_5847# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3278 a_27035_4546# a_26968_3954# a_27052_2983# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3279 a_36130_1486# a_36860_1242# a_37068_1242# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3280 a_435_905# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3281 a_30334_7257# a_30862_7509# a_31070_7509# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3282 vdd a_29321_4840# a_29113_4840# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3283 gnd a_23327_2283# a_23119_2283# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3284 a_10147_8836# a_10675_8631# a_10883_8631# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3285 a_8881_8181# a_9134_8168# a_7942_7871# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3286 a_6426_8977# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3287 a_35920_3138# a_35707_3138# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3288 a_35708_2589# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3289 gnd d2 a_33216_6189# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3290 a_21667_5035# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3291 a_116_9061# a_116_8831# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3292 gnd a_39353_2639# a_39145_2639# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3293 a_31071_8063# a_31801_7819# a_32009_7819# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3294 a_5489_4255# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3295 a_13858_3733# a_14111_3720# a_12919_3423# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3296 a_29065_2824# a_29068_2093# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3297 a_13858_2630# a_13854_2807# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3298 a_34037_9406# a_34294_9216# a_33102_8919# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3299 a_7060_387# a_6951_387# a_4954_326# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3300 a_10887_910# a_11618_1220# a_11826_1220# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3301 a_30336_3302# a_30864_3097# a_31072_3097# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3302 gnd a_9134_4305# a_8926_4305# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3303 vdd a_8057_1832# a_7849_1832# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3304 a_1902_5054# a_1895_346# a_2103_346# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3305 a_7801_8463# a_8054_8450# a_7832_7347# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3306 a_25888_8099# a_25675_8099# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3307 a_18907_7809# a_18912_7083# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3308 a_11834_7259# a_11543_6143# a_11824_5632# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3309 a_5702_7015# a_5489_7015# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3310 a_25362_1778# a_25889_2030# a_26097_2030# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3311 gnd d0 a_29320_8149# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3312 a_15205_6027# a_15734_5917# a_15942_5917# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3313 a_23068_7988# a_24055_7554# a_24006_7744# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3314 a_27033_8958# a_26612_8958# a_26094_8648# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3315 a_1584_7833# a_1371_7833# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3316 a_6427_7874# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3317 a_21667_7235# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3318 a_6428_4565# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3319 a_35391_5779# a_35920_5898# a_36128_5898# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3320 a_24011_8121# a_24007_8298# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3321 a_21769_8917# a_21556_8917# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3322 a_16895_5219# a_16568_7300# a_16895_7419# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3323 gnd d1 a_23326_4489# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3324 a_38160_5651# a_38413_5638# a_38015_6420# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3325 a_120_1110# a_122_1011# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3326 a_26096_5339# a_26827_5649# a_27035_5649# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3327 a_18908_5603# a_19165_5413# a_17970_5847# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3328 gnd a_24267_1490# a_24059_1490# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3329 a_31073_3651# a_31803_3407# a_32011_3407# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3330 a_7943_5665# a_8927_5962# a_8878_6152# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3331 vdd a_18118_5127# a_17910_5127# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3332 gnd d0 a_4079_3161# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3333 vdd a_23327_2283# a_23119_2283# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3334 gnd d2 a_28240_8431# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3335 a_17091_392# a_17910_5127# a_17861_5317# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3336 a_23071_8914# a_23324_8901# a_22931_8403# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3337 a_5703_5912# a_5490_5912# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3338 a_27246_368# a_28065_5103# a_28020_5116# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3339 gnd d1 a_18225_8966# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3340 a_3823_1145# a_4080_955# a_2885_1389# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3341 a_18914_2671# a_19167_2658# a_17975_2361# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3342 a_27034_7855# a_26613_7855# a_26096_8099# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3343 a_15207_1615# a_15736_1505# a_15944_1505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3344 a_15206_2718# a_15206_2489# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3345 a_23070_3576# a_24057_3142# a_24008_3332# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3346 a_17969_8053# a_18956_7619# a_18911_7632# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3347 a_31070_6406# a_30649_6406# a_30334_6611# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3348 a_31942_6124# a_31729_6124# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3349 a_27035_4546# a_26614_4546# a_26096_4236# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3350 a_6429_3462# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3351 a_1586_3421# a_1373_3421# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3352 gnd a_13169_8925# a_12961_8925# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3353 gnd a_39350_9257# a_38158_8960# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3354 a_32008_8922# a_31587_8922# a_31070_9166# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3355 a_13854_3910# a_14111_3720# a_12919_3423# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3356 vdd d0 a_9135_4859# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3357 a_11926_351# a_11713_351# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3358 gnd d1 a_3141_2302# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3359 a_15205_6214# a_15732_6466# a_15940_6466# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3360 a_38162_1239# a_38415_1226# a_38017_2008# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3361 a_26096_5339# a_25675_5339# a_25360_5087# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3362 a_26098_927# a_26829_1237# a_27037_1237# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3363 a_34044_954# a_34040_1131# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3364 a_9888_210# a_14663_331# a_12134_351# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3365 vdd a_14108_7578# a_13900_7578# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3366 a_7797_8640# a_8054_8450# a_7832_7347# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3367 a_12913_8012# a_13900_7578# a_13851_7768# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3368 a_1793_4524# a_1726_3932# a_1810_2961# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3369 a_18910_1191# a_19167_1001# a_17972_1435# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3370 a_21980_2299# a_21913_1707# a_21991_2823# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3371 a_18910_2848# a_18913_2117# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3372 a_30861_8612# a_30648_8612# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3373 vdd a_4079_4818# a_3871_4818# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3374 a_18911_9289# a_20302_9271# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3375 a_27045_7276# a_26754_6160# a_27035_5649# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3376 a_15734_4814# a_15521_4814# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3377 a_5175_2484# a_5175_2254# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3378 a_23068_7988# a_24055_7554# a_24010_7567# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3379 a_1694_5054# a_1481_5054# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3380 a_10149_5070# a_10149_4883# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3381 a_25675_6996# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3382 a_15520_4260# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3383 vdd d0 a_14111_960# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3384 a_16601_1772# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3385 a_29066_7608# a_29062_7785# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3386 gnd d0 a_24266_3696# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3387 a_13854_1150# a_14111_960# a_12916_1394# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3388 a_15939_8672# a_15518_8672# a_15203_8877# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3389 a_17829_6439# a_18019_5657# a_17970_5847# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3390 a_25887_7545# a_25674_7545# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3391 a_32020_7240# a_31911_7240# a_32025_5159# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3392 a_27137_368# a_26924_368# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3393 a_27036_3443# a_26615_3443# a_26098_3687# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3394 a_31072_1994# a_30651_1994# a_30336_2199# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3395 gnd d0 a_9135_2099# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3396 a_17971_3641# a_18958_3207# a_18913_3220# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3397 a_10149_4654# a_10678_4773# a_10886_4773# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3398 a_23073_4502# a_24057_4799# a_24008_4989# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3399 a_31800_8922# a_31587_8922# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3400 a_39099_4858# a_39352_4845# a_38160_4548# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3401 a_20618_7504# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3402 vdd d0 a_4079_3161# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3403 gnd a_4079_2058# a_3871_2058# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3404 vdd d2 a_28240_8431# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3405 a_35391_5549# a_35919_5344# a_36127_5344# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3406 gnd d0 a_19165_8173# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3407 vdd a_28380_8942# a_28172_8942# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3408 a_1694_7254# a_1481_7254# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3409 a_7799_4228# a_8056_4038# a_7834_2935# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3410 a_30335_4405# a_30336_3948# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3411 a_12915_3600# a_13902_3166# a_13853_3356# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3412 a_2882_8007# a_3139_7817# a_2741_8599# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3413 gnd a_14109_7029# a_13901_7029# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3414 a_34037_7749# a_34294_7559# a_33099_7993# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3415 a_23070_3576# a_24057_3142# a_24012_3155# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3416 vdd a_23184_8390# a_22976_8390# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3417 a_25677_2584# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3418 vdd a_29320_5389# a_29112_5389# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3419 a_15941_4260# a_16672_4570# a_16880_4570# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3420 a_3826_3174# a_3822_3351# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3421 gnd a_33216_6189# a_33008_6189# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3422 a_2747_4010# a_3000_3997# a_2778_2894# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3423 a_25889_3133# a_25676_3133# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3424 a_38158_1416# a_38415_1226# a_38017_2008# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3425 a_5172_9331# a_5701_9221# a_5909_9221# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3426 a_38014_8626# a_38204_7844# a_38155_8034# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3427 a_34043_4817# a_34296_4804# a_33104_4507# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3428 a_16813_3978# a_16600_3978# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3429 a_30336_3761# a_30865_3651# a_31073_3651# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3430 a_17974_4567# a_18958_4864# a_18913_4877# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3431 a_31802_4510# a_31589_4510# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3432 a_36645_4551# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3433 a_12779_1809# a_12964_2307# a_12915_2497# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3434 a_21994_7354# a_21697_8325# a_21978_7814# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3435 a_16879_6776# a_16458_6776# a_15941_7020# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3436 a_10884_9185# a_10463_9185# a_10147_9295# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3437 a_28124_8029# a_29111_7595# a_29062_7785# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3438 vdd d2 a_28242_4019# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3439 a_37078_2869# a_36787_1753# a_37067_2345# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3440 a_25675_8099# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3441 vdd d1 a_23325_7798# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3442 a_11544_3937# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3443 a_25361_2465# a_25890_2584# a_26098_2584# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3444 a_1792_6730# a_1371_6730# a_854_6974# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3445 a_7942_7871# a_8195_7858# a_7797_8640# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3446 a_12803_7488# a_13060_7298# a_12809_5099# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3447 a_32989_7469# a_33008_6189# a_32963_6202# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3448 a_30335_5967# a_30335_5738# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3449 a_34039_3337# a_34296_3147# a_33101_3581# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3450 a_22931_8403# a_23116_8901# a_23071_8914# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3451 a_1371_7833# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3452 a_21558_5608# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3453 a_18911_7632# a_19164_7619# a_17969_8053# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3454 a_20305_2424# a_20305_2194# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3455 a_36129_3692# a_36859_3448# a_37067_3448# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3456 a_21556_8917# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3457 gnd a_23326_4489# a_23118_4489# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3458 a_32020_5040# a_31700_2828# a_32022_2828# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3459 a_5913_1500# a_5492_1500# a_5176_1610# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3460 a_32958_8585# a_33148_7803# a_33099_7993# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3461 a_12919_3423# a_13172_3410# a_12774_4192# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3462 vdd d0 a_19165_8173# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3463 vdd d3 a_8087_2922# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3464 a_12915_3600# a_13902_3166# a_13857_3179# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3465 a_39097_7613# a_39350_7600# a_38155_8034# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3466 a_26098_927# a_25677_927# a_25364_1033# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3467 a_18909_2294# a_18915_1568# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3468 a_28126_3617# a_29113_3183# a_29064_3373# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3469 a_5490_5912# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3470 a_20308_992# a_20834_886# a_21042_886# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3471 gnd a_18225_8966# a_18017_8966# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3472 a_32995_5080# a_33038_7279# a_32993_7292# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3473 a_6569_3973# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3474 a_35392_2699# a_35921_2589# a_36129_2589# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3475 a_1794_2318# a_1373_2318# a_856_2562# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3476 a_116_9290# a_116_9061# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3477 a_30336_3532# a_30336_3302# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3478 a_25358_9312# a_25358_9083# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3479 a_22933_3991# a_23118_4489# a_23073_4502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3480 a_1373_3421# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3481 a_12913_8012# a_13170_7822# a_12772_8604# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3482 a_11839_7378# a_11542_8349# a_11823_7838# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3483 a_27036_2340# a_26969_1748# a_27047_2864# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3484 vdd a_9135_4859# a_8927_4859# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3485 a_15519_9226# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3486 a_29066_9265# a_29319_9252# a_28127_8955# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3487 a_26936_7276# a_26723_7276# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3488 a_10148_6630# a_10676_6425# a_10884_6425# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3489 a_6750_5095# a_6537_5095# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3490 a_32010_5613# a_31942_6124# a_32020_7240# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3491 vdd d0 a_9134_5408# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3492 vdd d4 a_33248_5067# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3493 a_26095_9202# a_25674_9202# a_25358_9312# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3494 a_30334_6841# a_30334_6611# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3495 a_21040_6955# a_20619_6955# a_20303_6836# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3496 a_17970_5847# a_18957_5413# a_18908_5603# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3497 a_15521_4814# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3498 a_39092_8893# a_39349_8703# a_38154_9137# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3499 a_20303_8168# a_20832_8058# a_21040_8058# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3500 a_1481_5054# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3501 a_435_905# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3502 a_18995_134# d8 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3503 a_16989_5100# a_16982_392# a_14985_331# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3504 a_117_7084# a_117_6855# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3505 gnd a_24266_3696# a_24058_3696# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3506 a_13859_1527# a_14112_1514# a_12920_1217# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3507 a_10883_8631# a_10462_8631# a_10148_8379# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3508 gnd d0 a_9136_2653# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3509 a_7942_7871# a_8926_8168# a_8877_8358# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3510 a_25674_7545# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3511 a_3825_7037# a_3821_7214# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3512 a_21980_3402# a_21559_3402# a_21041_3092# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3513 a_4954_326# a_6738_387# a_7060_387# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3514 gnd a_9135_2099# a_8927_2099# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3515 gnd a_38271_8436# a_38063_8436# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3516 gnd a_14109_5372# a_13901_5372# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3517 a_4632_326# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3518 a_5702_8118# a_5489_8118# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3519 a_7802_6257# a_8055_6244# a_7828_7524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3520 a_12915_3600# a_13172_3410# a_12774_4192# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3521 a_10149_5070# a_10677_5322# a_10885_5322# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3522 gnd a_4080_2612# a_3872_2612# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3523 a_23069_5782# a_24056_5348# a_24007_5538# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3524 a_10150_2218# a_10678_2013# a_10886_2013# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3525 a_32009_7819# a_31588_7819# a_31070_7509# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3526 a_6428_5668# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3527 a_12919_3423# a_13903_3720# a_13854_3910# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3528 a_28126_3617# a_29113_3183# a_29068_3196# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3529 gnd a_19165_8173# a_18957_8173# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3530 a_1585_5627# a_1372_5627# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3531 a_22964_5075# a_23217_5062# a_22190_327# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3532 a_6429_2359# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3533 a_117_7958# a_646_8077# a_854_8077# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3534 a_1481_7254# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3535 a_13853_6116# a_14110_5926# a_12918_5629# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3536 a_21041_5852# a_20620_5852# a_20304_5962# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3537 a_1583_8936# a_1370_8936# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3538 gnd d4 a_18118_5127# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3539 gnd d1 a_3140_4508# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3540 a_21042_2543# a_20621_2543# a_20305_2424# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3541 a_7832_7347# a_7846_8450# a_7797_8640# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3542 gnd d2 a_13031_4002# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3543 a_5173_8415# a_5173_8228# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3544 a_5910_4255# a_5489_4255# a_5174_4460# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3545 gnd d0 a_4080_955# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3546 a_25676_3133# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3547 a_27050_7395# a_26753_8366# a_27034_7855# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3548 a_29062_9442# a_29319_9252# a_28127_8955# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3549 gnd d2 a_28241_6225# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3550 a_16600_3978# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3551 gnd a_14111_960# a_13903_960# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3552 a_14663_331# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3553 vdd d1 a_28381_7839# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3554 gnd a_28381_6736# a_28173_6736# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3555 a_7804_1845# a_8057_1832# a_7830_3112# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3556 a_39095_3378# a_39100_2652# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3557 a_15941_7020# a_15520_7020# a_15204_6901# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3558 a_27035_5649# a_26614_5649# a_26097_5893# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3559 a_34042_5366# a_34295_5353# a_33100_5787# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3560 a_23071_1370# a_24058_936# a_24009_1126# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3561 a_13856_8145# a_13852_8322# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3562 a_17970_5847# a_18957_5413# a_18912_5426# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3563 a_31071_4200# a_30650_4200# a_30335_4405# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3564 vdd a_28242_4019# a_28034_4019# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3565 a_32022_2828# a_31731_1712# a_32012_1201# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3566 gnd d0 a_14108_7578# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3567 vdd a_23325_7798# a_23117_7798# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3568 a_854_6974# a_433_6974# a_117_6855# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3569 a_12134_351# a_11713_351# a_12035_351# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3570 a_1587_1215# a_1374_1215# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3571 a_39096_8716# a_39092_8893# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3572 vdd d0 a_34297_941# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3573 a_13855_1704# a_14112_1514# a_12920_1217# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3574 a_35390_6652# a_35391_6195# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3575 vdd d0 a_39350_6497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3576 vdd d0 a_9136_2653# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3577 a_15206_4008# a_15733_4260# a_15941_4260# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3578 vdd a_38271_8436# a_38063_8436# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3579 vdd a_14109_5372# a_13901_5372# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3580 a_17975_2361# a_18959_2658# a_18910_2848# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3581 a_18907_6706# a_18913_5980# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3582 a_7798_6434# a_8055_6244# a_7828_7524# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3583 a_1794_2318# a_1727_1726# a_1805_2842# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3584 a_37064_8963# a_36997_8371# a_37081_7400# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3585 a_30862_6406# a_30649_6406# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3586 a_16781_5100# a_16568_5100# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3587 vdd a_4080_2612# a_3872_2612# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3588 a_10147_9066# a_10147_8836# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3589 a_15735_2608# a_15522_2608# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3590 a_3824_9243# a_4077_9230# a_2885_8933# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3591 vdd a_39350_9257# a_39142_9257# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3592 gnd d2 a_28243_1813# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3593 a_12919_3423# a_13903_3720# a_13858_3733# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3594 vdd d1 a_28383_3427# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3595 vdd a_19165_8173# a_18957_8173# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3596 vdd a_29319_7595# a_29111_7595# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3597 a_22960_5252# a_23217_5062# a_22190_327# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3598 a_6850_2359# a_6429_2359# a_5912_2603# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3599 a_5701_7564# a_5488_7564# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3600 a_24011_7018# a_24007_7195# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3601 a_25888_5339# a_25675_5339# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3602 vdd a_23186_3978# a_22978_3978# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3603 a_27037_1237# a_26616_1237# a_26099_1481# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3604 a_34044_954# a_34297_941# a_33102_1375# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3605 a_13853_3356# a_13858_2630# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3606 a_38154_9137# a_38411_8947# a_38018_8449# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3607 a_855_5871# a_434_5871# a_118_5981# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3608 a_20831_9161# a_20618_9161# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3609 a_7832_7347# a_7846_8450# a_7801_8463# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3610 a_1810_2961# a_1513_3932# a_1794_3421# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3611 a_17972_1435# a_18959_1001# a_18914_1014# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3612 a_10150_2448# a_10679_2567# a_10887_2567# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3613 a_856_2562# a_435_2562# a_119_2443# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3614 a_30335_5967# a_30864_5857# a_31072_5857# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3615 a_31801_6716# a_31588_6716# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3616 a_36644_6757# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3617 a_26967_6160# a_26754_6160# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3618 a_13854_8694# a_13850_8871# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3619 a_24012_5915# a_24265_5902# a_23073_5605# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3620 vdd d2 a_28241_6225# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3621 a_35392_3343# a_35920_3138# a_36128_3138# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3622 gnd d0 a_9133_7614# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3623 gnd d0 a_19166_5967# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3624 a_25360_4671# a_25889_4790# a_26097_4790# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3625 a_33106_1198# a_34090_1495# a_34045_1508# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3626 vdd a_28381_6736# a_28173_6736# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3627 a_5174_6022# a_5174_5793# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3628 gnd d3 a_28273_2903# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3629 gnd d0 a_24263_9211# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3630 a_30864_1994# a_30651_1994# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3631 a_35392_3573# a_35392_3343# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3632 a_10886_4773# a_10465_4773# a_10149_4883# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3633 a_32993_7292# a_33007_8395# a_32962_8408# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3634 a_26723_7276# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3635 a_34038_5543# a_34295_5353# a_33100_5787# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3636 a_10151_1115# a_10153_1016# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3637 a_25359_8396# a_25359_8209# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3638 a_25359_8209# a_25888_8099# a_26096_8099# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3639 vdd a_33248_5067# a_33040_5067# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3640 a_5172_8872# a_5173_8415# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3641 vdd a_9134_5408# a_8926_5408# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3642 a_5703_3152# a_5490_3152# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3643 gnd d1 a_33355_8906# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3644 a_7834_2935# a_7848_4038# a_7803_4051# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3645 a_5173_7125# a_5702_7015# a_5910_7015# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3646 a_12918_5629# a_13171_5616# a_12773_6398# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3647 a_31802_5613# a_31589_5613# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3648 a_30337_1555# a_30866_1445# a_31074_1445# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3649 a_34044_2611# a_34297_2598# a_33105_2301# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3650 a_36646_2345# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3651 a_120_1569# a_120_1340# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3652 a_31803_2304# a_31590_2304# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3653 gnd a_9136_2653# a_8928_2653# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3654 a_29069_3750# a_29065_3927# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3655 a_21989_7235# a_21698_6119# a_21979_5608# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3656 a_28125_5823# a_29112_5389# a_29063_5579# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3657 a_15206_2259# a_15734_2054# a_15942_2054# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3658 a_3820_9420# a_4077_9230# a_2885_8933# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3659 vdd d1 a_3139_7817# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3660 vdd d1 a_23326_5592# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3661 a_5175_2484# a_5704_2603# a_5912_2603# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3662 a_10151_1115# a_10679_910# a_10887_910# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3663 a_29066_6505# a_29062_6682# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3664 a_16459_5673# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3665 a_22930_1962# a_23120_1180# a_23071_1370# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3666 a_21991_2823# a_21700_1707# a_21980_2299# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3667 a_28130_3440# a_29114_3737# a_29069_3750# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3668 a_5909_9221# a_5488_9221# a_5172_9102# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3669 a_24006_7744# a_24011_7018# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3670 a_25360_4441# a_25361_3984# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3671 a_22932_6197# a_23117_6695# a_23072_6708# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3672 a_1372_5627# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3673 gnd a_18118_5127# a_17910_5127# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3674 a_1370_8936# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3675 a_18909_6157# a_18912_5426# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3676 a_5174_5793# a_5703_5912# a_5911_5912# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3677 a_32959_6379# a_33149_5597# a_33100_5787# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3678 a_32009_7819# a_31941_8330# a_32025_7359# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3679 a_5174_5793# a_5174_5563# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3680 a_7797_8640# a_7987_7858# a_7938_8048# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3681 vdd d0 a_9133_7614# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3682 a_12809_5099# a_12852_7298# a_12807_7311# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3683 a_31804_1201# a_31591_1201# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3684 vdd d0 a_24263_9211# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3685 a_39098_5407# a_39351_5394# a_38156_5828# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3686 a_34045_1508# a_34041_1685# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3687 a_15209_1057# a_15735_951# a_15943_951# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3688 a_17969_8053# a_18956_7619# a_18907_7809# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3689 a_28127_1411# a_29114_977# a_29065_1167# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3690 a_31913_2828# a_31700_2828# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3691 a_10884_6425# a_11615_6735# a_11823_6735# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3692 a_22289_327# a_21868_327# a_22088_5035# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3693 a_12774_4192# a_12964_3410# a_12915_3600# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3694 a_3826_2071# a_3822_2248# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3695 a_33099_6890# a_33356_6700# a_32963_6202# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3696 a_30337_1555# a_30337_1326# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3697 gnd a_14108_7578# a_13900_7578# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3698 a_1374_1215# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3699 a_30334_8360# a_30861_8612# a_31069_8612# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3700 a_12914_5806# a_13171_5616# a_12773_6398# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3701 a_31071_8063# a_30650_8063# a_30334_7944# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3702 vdd d0 a_4079_5921# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3703 a_15944_1505# a_16674_1261# a_16882_1261# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3704 a_10148_7276# a_10676_7528# a_10884_7528# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3705 a_30334_7714# a_30334_7257# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3706 vdd a_9136_2653# a_8928_2653# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3707 a_8880_9284# a_9133_9271# a_7941_8974# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3708 a_853_7523# a_432_7523# a_117_7271# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3709 a_10149_4424# a_10677_4219# a_10885_4219# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3710 a_20302_8812# a_20303_8355# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3711 gnd d1 a_28382_5633# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3712 a_32011_3407# a_31943_3918# a_32027_2947# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3713 a_644_8626# a_431_8626# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3714 vdd d0 a_9135_3202# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3715 a_26096_6996# a_25675_6996# a_25359_7106# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3716 a_10679_3670# a_10466_3670# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3717 a_23073_5605# a_24057_5902# a_24012_5915# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3718 a_9987_210# a_19208_134# vout gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3719 a_12772_8604# a_12962_7822# a_12917_7835# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3720 a_21041_4749# a_20620_4749# a_20304_4630# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3721 a_22930_1962# a_23120_1180# a_23075_1193# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3722 a_39100_995# a_39353_982# a_38158_1416# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3723 a_15522_2608# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3724 gnd d2 a_13030_6208# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3725 a_30335_4864# a_30335_4635# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3726 a_6866_3002# a_6569_3973# a_6850_3462# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3727 gnd a_28243_1813# a_28035_1813# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3728 a_10150_3551# a_10150_3321# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3729 a_31070_9166# a_31800_8922# a_32008_8922# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3730 a_10884_6425# a_10463_6425# a_10149_6173# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3731 a_10886_2013# a_11617_2323# a_11825_2323# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3732 a_25675_5339# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3733 a_33101_2478# a_33358_2288# a_32965_1790# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3734 a_25887_9202# a_25674_9202# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3735 a_15205_6214# a_15205_6027# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3736 gnd a_14110_3166# a_13902_3166# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3737 a_26754_6160# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3738 a_7803_4051# a_8056_4038# a_7834_2935# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3739 a_12916_1394# a_13173_1204# a_12775_1986# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3740 vdd d0 a_4081_1509# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3741 a_15940_9226# a_15519_9226# a_15203_9107# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3742 gnd d0 a_29319_9252# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3743 a_10150_2864# a_10678_3116# a_10886_3116# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3744 a_34041_7572# a_34294_7559# a_33099_7993# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3745 gnd a_39351_7051# a_39143_7051# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3746 a_855_3111# a_434_3111# a_119_2859# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3747 a_13857_3179# a_13853_3356# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3748 gnd d1 a_28384_1221# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3749 a_12920_1217# a_13904_1514# a_13855_1704# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3750 a_32027_2947# a_31730_3918# a_32011_3407# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3751 gnd a_9133_7614# a_8925_7614# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3752 gnd a_19166_5967# a_18958_5967# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3753 a_2778_5094# a_3031_5081# a_2004_346# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3754 a_35390_6882# a_35919_7001# a_36127_7001# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3755 a_646_4214# a_433_4214# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3756 gnd a_28273_2903# a_28065_2903# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3757 gnd a_24263_9211# a_24055_9211# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3758 a_34039_6097# a_34296_5907# a_33104_5610# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3759 a_21042_3646# a_20621_3646# a_20305_3756# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3760 gnd a_23187_1772# a_22979_1772# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3761 a_30651_1994# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3762 vdd d0 a_39349_8703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3763 a_38159_6754# a_38412_6741# a_38019_6243# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3764 a_23075_1193# a_24059_1490# a_24014_1503# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3765 a_30336_2429# a_30336_2199# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3766 a_2772_7483# a_3029_7293# a_2778_5094# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3767 a_8877_7255# a_8880_6524# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3768 a_7828_7524# a_7847_6244# a_7798_6434# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3769 a_26095_6442# a_26826_6752# a_27034_6752# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3770 a_20304_5733# a_20304_5503# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3771 a_16880_4570# a_16813_3978# a_16897_3007# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3772 a_12774_4192# a_12964_3410# a_12919_3423# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3773 a_5911_2049# a_5490_2049# a_5175_2254# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3774 a_10885_5322# a_10464_5322# a_10149_5527# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3775 a_31072_4754# a_31802_4510# a_32010_4510# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3776 a_10886_2013# a_10465_2013# a_10151_1761# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3777 a_34042_8126# a_34038_8303# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3778 a_5490_3152# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3779 a_5910_8118# a_6640_7874# a_6848_7874# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3780 a_8876_9461# a_9133_9271# a_7941_8974# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3781 gnd a_33355_8906# a_33147_8906# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3782 gnd d2 a_28242_4019# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3783 gnd a_2999_6203# a_2791_6203# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3784 a_12918_5629# a_13902_5926# a_13857_5939# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3785 vdd d1 a_28382_5633# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3786 a_10147_9295# a_10147_9066# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3787 a_15941_8123# a_15520_8123# a_15204_8233# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3788 a_31590_2304# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3789 gnd d0 a_29321_4840# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3790 a_34043_3160# a_34296_3147# a_33101_3581# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3791 a_22088_5035# a_21667_5035# a_21994_5154# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3792 vdd a_23326_5592# a_23118_5592# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3793 a_855_4768# a_434_4768# a_118_4649# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3794 a_30649_9166# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3795 a_27983_8621# a_28173_7839# a_28128_7852# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3796 a_11824_5632# a_11403_5632# a_10885_5322# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3797 a_26966_8366# a_26753_8366# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3798 a_11839_5178# a_11725_5059# a_11933_5059# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3799 vdd d0 a_39351_4291# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3800 a_11822_8941# a_11401_8941# a_10884_9185# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3801 a_24011_8121# a_24264_8108# a_23072_7811# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3802 a_29069_990# a_29065_1167# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3803 a_7830_3112# a_7849_1832# a_7800_2022# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3804 a_26095_6442# a_25674_6442# a_25360_6190# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3805 a_13851_9425# a_13854_8694# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3806 a_36860_1242# a_36647_1242# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3807 vdd a_14110_3166# a_13902_3166# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3808 a_15206_3362# a_15206_2905# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3809 a_21697_8325# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3810 a_30863_4200# a_30650_4200# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3811 a_36787_1753# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3812 vdd d0 a_29319_9252# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3813 a_23067_9091# a_24054_8657# a_24009_8670# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3814 a_37065_6757# a_36998_6165# a_37076_7281# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3815 a_3825_7037# a_4078_7024# a_2886_6727# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3816 a_39098_7064# a_39094_7241# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3817 vdd a_39351_7051# a_39143_7051# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3818 a_5912_3706# a_6642_3462# a_6850_3462# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3819 a_33102_1375# a_34089_941# a_34044_954# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3820 gnd d1 a_3140_5611# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3821 vdd d1 a_28384_1221# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3822 a_31591_1201# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3823 a_12920_1217# a_13904_1514# a_13859_1527# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3824 vdd a_9133_7614# a_8925_7614# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3825 a_32995_5080# a_33038_7279# a_32989_7469# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3826 a_17833_6262# a_18018_6760# a_17969_6950# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3827 a_2774_5271# a_3031_5081# a_2004_346# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3828 a_28131_1234# a_29115_1531# a_29066_1721# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3829 vdd a_24263_9211# a_24055_9211# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3830 a_32995_2880# a_33009_3983# a_32964_3996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3831 a_39101_1549# a_39097_1726# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3832 vdd a_23187_1772# a_22979_1772# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3833 a_13857_2076# a_14110_2063# a_12915_2497# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3834 a_11834_7259# a_11725_7259# a_11839_5178# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3835 a_38155_6931# a_38412_6741# a_38019_6243# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3836 a_5702_5358# a_5489_5358# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3837 a_856_3665# a_435_3665# a_119_3775# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3838 a_22931_8403# a_23184_8390# a_22962_7287# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3839 a_7828_7524# a_7847_6244# a_7802_6257# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3840 a_1805_2842# a_1514_1726# a_1795_1215# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3841 a_31700_2828# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3842 gnd d2 a_2998_8409# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3843 a_31801_7819# a_31588_7819# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3844 a_15204_6671# a_15205_6214# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3845 a_11826_1220# a_11405_1220# a_10887_910# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3846 a_27985_4209# a_28175_3427# a_28130_3440# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3847 a_2885_8933# a_3869_9230# a_3820_9420# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3848 a_6864_5214# a_6750_5095# a_6958_5095# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3849 a_26097_2030# a_25676_2030# a_25362_1778# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3850 gnd d4 a_33248_5067# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3851 a_16458_7879# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3852 vdd a_18086_6249# a_17878_6249# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3853 a_39095_2275# a_39101_1549# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3854 a_28129_5646# a_29113_5943# a_29068_5956# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3855 a_39099_4858# a_39095_5035# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3856 a_10887_2567# a_10466_2567# a_10150_2677# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3857 a_13856_7042# a_13852_7219# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3858 a_431_8626# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3859 a_36126_9207# a_36856_8963# a_37064_8963# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3860 a_30337_1742# a_30337_1555# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3861 vdd a_9135_3202# a_8927_3202# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3862 a_10466_3670# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3863 a_34036_8852# a_34042_8126# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3864 a_6537_7295# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3865 a_24009_1126# a_20308_992# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3866 vdd a_39353_982# a_39145_982# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3867 a_38157_2519# a_38414_2329# a_38021_1831# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3868 a_5173_7999# a_5702_8118# a_5910_8118# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3869 gnd d0 a_4080_3715# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3870 a_28016_3093# a_28273_2903# a_28016_5293# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3871 a_31803_3407# a_31590_3407# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3872 vdd d1 a_18227_5657# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3873 a_15206_2905# a_15734_3157# a_15942_3157# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3874 gnd a_14111_3720# a_13903_3720# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3875 a_9779_210# a_9566_210# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3876 a_25674_9202# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3877 a_3821_7214# a_4078_7024# a_2886_6727# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3878 vdd d1 a_3140_5611# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3879 a_30335_5051# a_30335_4864# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3880 a_17833_6262# a_18018_6760# a_17973_6773# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3881 a_7941_8974# a_8194_8961# a_7801_8463# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3882 a_39095_6138# a_39352_5948# a_38160_5651# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3883 a_28131_1234# a_29115_1531# a_29070_1544# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3884 a_5176_1610# a_5176_1381# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3885 a_17861_3117# a_17880_1837# a_17831_2027# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3886 a_12773_6398# a_12963_5616# a_12914_5806# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3887 a_13857_4836# a_13853_5013# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3888 a_13853_2253# a_14110_2063# a_12915_2497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3889 a_33098_9096# a_33355_8906# a_32962_8408# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3890 a_21557_6711# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3891 a_18910_8735# a_19163_8722# a_17968_9156# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3892 a_31911_5040# a_31698_5040# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3893 a_433_4214# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3894 a_36128_4795# a_36858_4551# a_37066_4551# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3895 a_1724_8344# a_1511_8344# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3896 a_21868_327# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3897 a_2885_8933# a_3869_9230# a_3824_9243# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3898 a_14985_331# a_16769_392# a_17091_392# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3899 a_5912_2603# a_5491_2603# a_5175_2713# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3900 a_6539_2883# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3901 vdd d0 a_29318_8698# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3902 a_12914_4703# a_13901_4269# a_13856_4282# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3903 a_8880_1740# a_8883_1009# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3904 a_21913_1707# a_21700_1707# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3905 a_10678_5876# a_10465_5876# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3906 vdd d0 a_24264_7005# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3907 a_5174_4919# a_5174_4690# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3908 a_39099_3201# a_39352_3188# a_38157_3622# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3909 gnd a_28242_4019# a_28034_4019# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3910 a_25359_7293# a_25359_7106# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3911 a_32025_5159# a_31698_7240# a_32020_7240# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3912 a_16880_5673# a_16459_5673# a_15941_5363# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3913 vdd d1 a_3142_1199# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3914 a_10885_4219# a_11616_4529# a_11824_4529# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3915 a_119_3316# a_119_2859# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3916 a_33100_4684# a_33357_4494# a_32964_3996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3917 a_16812_6184# a_16599_6184# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3918 a_18912_4323# a_19165_4310# a_17970_4744# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3919 a_26753_8366# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3920 a_30335_6154# a_30862_6406# a_31070_6406# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3921 a_16890_5100# a_16781_5100# a_16989_5100# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3922 vdd d0 a_4080_3715# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3923 a_8880_9284# a_10147_9295# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3924 gnd a_39350_9257# a_39142_9257# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3925 a_8881_7078# a_9134_7065# a_7942_6768# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3926 a_854_5317# a_433_5317# a_118_5065# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3927 vdd a_14111_3720# a_13903_3720# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3928 a_29069_2647# a_29065_2824# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3929 a_21769_8917# a_21556_8917# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3930 gnd d1 a_28383_3427# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3931 a_645_6420# a_432_6420# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3932 a_35920_2035# a_35707_2035# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3933 a_35389_9088# a_35918_9207# a_36126_9207# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3934 a_11824_5632# a_11756_6143# a_11834_7259# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3935 vdd d0 a_9136_996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3936 a_5173_7769# a_5701_7564# a_5909_7564# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3937 a_30650_4200# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3938 a_23074_3399# a_24058_3696# a_24013_3709# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3939 a_20302_9271# a_20831_9161# a_21039_9161# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3940 a_24006_6641# a_24012_5915# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3941 a_12773_6398# a_12963_5616# a_12918_5629# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3942 a_5176_1151# a_5704_946# a_5912_946# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3943 a_35062_312# a_34849_312# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3944 a_30863_8063# a_30650_8063# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3945 a_16882_1261# a_16461_1261# a_15943_951# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3946 a_6861_2883# a_6570_1767# a_6851_1256# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3947 a_18906_8912# a_19163_8722# a_17968_9156# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3948 a_10884_7528# a_10463_7528# a_10148_7733# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3949 a_31071_6960# a_31801_6716# a_32009_6716# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3950 a_27984_6415# a_28174_5633# a_28125_5823# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3951 a_7941_8974# a_8925_9271# a_8876_9461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3952 a_5703_5912# a_5490_5912# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3953 a_10885_4219# a_10464_4219# a_10150_3967# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3954 a_10151_1574# a_10151_1345# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3955 a_5701_9221# a_5488_9221# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3956 a_25888_6996# a_25675_6996# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3957 gnd d4 a_38304_5108# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3958 a_18909_5054# a_18912_4323# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3959 gnd a_2998_8409# a_2790_8409# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3960 gnd a_18085_8455# a_17877_8455# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3961 gnd d0 a_34295_8113# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3962 gnd d0 a_29320_7046# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3963 a_15205_4924# a_15734_4814# a_15942_4814# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3964 a_21669_2823# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3965 a_23068_6885# a_24055_6451# a_24006_6641# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3966 a_118_5981# a_647_5871# a_855_5871# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3967 a_10153_1016# a_10679_910# a_10887_910# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3968 a_32008_8922# a_31587_8922# a_31069_8612# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3969 a_1584_6730# a_1371_6730# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3970 a_6427_6771# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3971 a_35921_932# a_35708_932# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3972 gnd a_33248_5067# a_33040_5067# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3973 a_13855_1704# a_13858_973# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3974 a_11823_7838# a_11402_7838# a_10884_7528# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3975 a_25359_7750# a_25359_7293# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3976 a_30652_891# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3977 a_647_2008# a_434_2008# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3978 a_21043_1440# a_20622_1440# a_20306_1550# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3979 a_34040_3891# a_34297_3701# a_33105_3404# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3980 a_5175_3357# a_5703_3152# a_5911_3152# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3981 a_38160_4548# a_38413_4535# a_38020_4037# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3982 a_7834_2935# a_7848_4038# a_7799_4228# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3983 a_15207_1156# a_15735_951# a_15943_951# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3984 a_12775_1986# a_12965_1204# a_12920_1217# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3985 a_26094_8648# a_25673_8648# a_25359_8396# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3986 a_31071_5303# a_31802_5613# a_32010_5613# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3987 a_26096_4236# a_26827_4546# a_27035_4546# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3988 a_18908_4500# a_19165_4310# a_17970_4744# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3989 a_27986_2003# a_28176_1221# a_28127_1411# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3990 a_31073_2548# a_31803_2304# a_32011_2304# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3991 vdd d3 a_23217_2862# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3992 a_10886_3116# a_10465_3116# a_10150_3321# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3993 a_16568_7300# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3994 a_3821_5557# a_4078_5367# a_2883_5801# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3995 a_5705_1500# a_5492_1500# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3996 a_25360_4900# a_25360_4671# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3997 a_5911_5912# a_6641_5668# a_6849_5668# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3998 a_2004_346# a_2823_5081# a_2774_5271# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3999 a_39099_2098# a_39095_2275# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4000 a_8877_7255# a_9134_7065# a_7942_6768# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4001 gnd a_3000_3997# a_2792_3997# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4002 a_19208_134# a_18995_134# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4003 a_35393_1783# a_35393_1596# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4004 a_31590_3407# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4005 a_15942_5917# a_15521_5917# a_15205_6027# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4006 gnd a_18087_4043# a_17879_4043# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4007 a_15206_3592# a_15735_3711# a_15943_3711# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4008 a_5908_8667# a_6639_8977# a_6847_8977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4009 a_27034_6752# a_26613_6752# a_26096_6996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4010 vdd a_18227_5657# a_18019_5657# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4011 a_28130_3440# a_29114_3737# a_29065_3927# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4012 a_12775_1986# a_13032_1796# a_12805_3076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4013 gnd d0 a_14107_8681# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4014 vdd d3 a_18116_7339# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4015 a_15519_7569# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4016 a_29066_7608# a_29319_7595# a_28124_8029# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4017 a_27984_6415# a_28174_5633# a_28129_5646# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4018 a_11825_3426# a_11404_3426# a_10886_3116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4019 a_10150_2448# a_10150_2218# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4020 a_6780_8385# a_6567_8385# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4021 a_13854_2807# a_14111_2617# a_12919_2320# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4022 a_7941_8974# a_8925_9271# a_8880_9284# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4023 vdd d3 a_3029_7293# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4024 a_16598_8390# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4025 a_26095_7545# a_25674_7545# a_25359_7750# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4026 a_118_5752# a_118_5522# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4027 a_35389_8858# a_35917_8653# a_36125_8653# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4028 a_39094_8344# a_39097_7613# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4029 vdd a_13060_7298# a_12852_7298# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4030 vdd d0 a_24264_5348# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4031 a_26096_4236# a_25675_4236# a_25361_3984# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4032 a_12913_6909# a_13900_6475# a_13851_6665# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4033 a_1511_8344# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4034 a_21698_6119# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4035 vdd a_18085_8455# a_17877_8455# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4036 gnd d1 a_18228_3451# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4037 vdd d0 a_34295_8113# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4038 vdd d0 a_29320_7046# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4039 a_23068_6885# a_24055_6451# a_24010_6464# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4040 a_3826_4831# a_4079_4818# a_2887_4521# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4041 a_5913_1500# a_6643_1256# a_6851_1256# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4042 a_13857_2076# a_13853_2253# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4043 a_32027_2947# a_31913_2828# a_32020_5040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4044 vdd a_29318_8698# a_29110_8698# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4045 a_36127_8104# a_35706_8104# a_35390_7985# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4046 a_11933_5059# a_11512_5059# a_11834_5059# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4047 a_37081_5200# a_36754_7281# a_37076_7281# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4048 a_24008_6092# a_24011_5361# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4049 a_17834_4056# a_18019_4554# a_17970_4744# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4050 a_21700_1707# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4051 gnd d0 a_24266_2593# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4052 a_12805_3076# a_13062_2886# a_12805_5276# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4053 a_10465_5876# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4054 a_39100_3755# a_39353_3742# a_38161_3445# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4055 vdd a_24264_7005# a_24056_7005# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4056 a_25887_6442# a_25674_6442# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4057 a_38156_4725# a_38413_4535# a_38020_4037# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4058 a_857_1459# a_436_1459# a_120_1569# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4059 a_20832_8058# a_20619_8058# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4060 a_22932_6197# a_23185_6184# a_22958_7464# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4061 gnd a_39350_7600# a_39142_7600# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4062 vdd a_3142_1199# a_2934_1199# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4063 a_27986_2003# a_28176_1221# a_28131_1234# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4064 vdd d1 a_18226_7863# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4065 a_20618_6401# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4066 vdd d0 a_4079_2058# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4067 a_1696_2842# a_1483_2842# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4068 a_26097_3133# a_25676_3133# a_25361_3338# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4069 a_2004_346# a_2823_5081# a_2778_5094# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4070 a_35391_4446# a_35919_4241# a_36127_4241# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4071 gnd d0 a_19165_7070# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4072 a_12915_2497# a_13902_2063# a_13853_2253# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4073 a_17832_8468# a_18017_8966# a_17972_8979# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4074 a_11839_5178# a_11512_7259# a_11839_7378# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4075 vdd a_18087_4043# a_17879_4043# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4076 a_22962_7287# a_22976_8390# a_22927_8580# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4077 vdd a_13170_7822# a_12962_7822# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4078 a_23070_2473# a_24057_2039# a_24012_2052# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4079 a_21556_8917# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4080 vdd d0 a_14107_8681# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4081 a_432_6420# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4082 a_36127_7001# a_36857_6757# a_37065_6757# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4083 vdd a_9136_996# a_8928_996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4084 a_6958_5095# a_6537_5095# a_6859_5095# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4085 a_10467_1464# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4086 a_25889_2030# a_25676_2030# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4087 a_7834_5135# a_8087_5122# a_7060_387# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4088 a_5911_4809# a_5490_4809# a_5174_4919# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4089 a_15941_5363# a_15520_5363# a_15205_5111# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4090 a_30650_8063# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4091 a_22081_327# a_21868_327# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4092 a_12913_6909# a_13900_6475# a_13855_6488# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4093 a_5490_5912# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4094 a_15206_2259# a_15207_1802# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4095 a_28020_5116# a_28063_7315# a_28014_7505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4096 a_28124_6926# a_29111_6492# a_29062_6682# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4097 vdd d1 a_18228_3451# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4098 a_30333_9047# a_30333_8817# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4099 a_25675_6996# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4100 gnd a_38304_5108# a_38096_5108# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4101 a_35171_312# a_36955_373# a_37277_373# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4102 vdd d1 a_3141_3405# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4103 a_17834_4056# a_18019_4554# a_17974_4567# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4104 gnd a_34295_8113# a_34087_8113# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4105 a_20304_6149# a_20304_5962# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4106 a_27144_5076# a_26723_5076# a_27045_5076# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4107 a_39096_3932# a_39353_3742# a_38161_3445# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4108 a_21557_7814# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4109 a_10151_1761# a_10151_1574# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4110 a_1371_6730# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4111 a_36127_5344# a_36858_5654# a_37066_5654# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4112 a_21558_4505# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4113 a_16811_8390# a_16598_8390# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4114 a_18911_6529# a_19164_6516# a_17969_6950# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4115 a_22928_6374# a_23185_6184# a_22958_7464# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4116 a_434_2008# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4117 a_3824_7586# a_4077_7573# a_2882_8007# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4118 a_36129_2589# a_36859_2345# a_37067_2345# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4119 a_1725_6138# a_1512_6138# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4120 a_20306_1091# a_20834_886# a_21042_886# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4121 a_16814_1772# a_16601_1772# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4122 a_32963_6202# a_33148_6700# a_33099_6890# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4123 vdd a_14110_5926# a_13902_5926# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4124 a_7801_8463# a_7986_8961# a_7937_9151# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4125 vdd d0 a_9132_8717# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4126 vdd d0 a_19165_7070# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4127 a_8877_5598# a_8882_4872# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4128 a_12915_2497# a_13902_2063# a_13857_2076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4129 vdd a_23217_2862# a_23009_2862# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4130 a_11823_7838# a_11755_8349# a_11839_7378# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4131 a_5492_1500# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4132 a_17968_9156# a_18955_8722# a_18906_8912# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4133 a_25239_307# a_24818_307# a_25140_307# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4134 a_28126_2514# a_29113_2080# a_29064_2270# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4135 a_11545_1731# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4136 a_27050_5195# a_26723_7276# a_27050_7395# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4137 a_10677_6979# a_10464_6979# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4138 a_16881_3467# a_16460_3467# a_15942_3157# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4139 a_20305_3943# a_20305_3756# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4140 a_38158_1416# a_39145_982# a_39100_995# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4141 a_21559_3402# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4142 gnd d0 a_24263_7554# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4143 vdd a_18116_7339# a_17908_7339# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4144 a_7830_5312# a_8087_5122# a_7060_387# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4145 gnd a_14107_8681# a_13899_8681# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4146 a_12913_6909# a_13170_6719# a_12777_6221# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4147 a_36129_932# a_36860_1242# a_37068_1242# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4148 a_8875_8907# a_8881_8181# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4149 a_30336_3948# a_30863_4200# a_31071_4200# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4150 a_3826_3174# a_4079_3161# a_2884_3595# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4151 a_10148_8379# a_10675_8631# a_10883_8631# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4152 a_23067_9091# a_24054_8657# a_24005_8847# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4153 a_28020_5116# a_28063_7315# a_28018_7328# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4154 a_37083_2988# a_36969_2869# a_37076_5081# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4155 a_1583_8936# a_1370_8936# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4156 vdd a_24264_5348# a_24056_5348# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4157 a_8882_4872# a_9135_4859# a_7943_4562# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4158 a_32112_332# a_31899_332# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4159 a_35920_3138# a_35707_3138# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4160 a_13856_8145# a_14109_8132# a_12917_7835# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4161 a_6567_8385# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4162 a_35391_6008# a_35391_5779# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4163 a_11825_3426# a_11757_3937# a_11841_2966# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4164 a_20833_3092# a_20620_3092# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4165 gnd d0 a_34297_3701# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4166 a_5174_5563# a_5702_5358# a_5910_5358# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4167 a_21667_5035# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4168 gnd a_18228_3451# a_18020_3451# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4169 vdd a_34295_8113# a_34087_8113# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4170 a_17970_4744# a_18957_4310# a_18908_4500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4171 a_31070_7509# a_31801_7819# a_32009_7819# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4172 a_16989_5100# a_16568_5100# a_16895_5219# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4173 vdd d2 a_18088_1837# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4174 a_35389_8858# a_35390_8401# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4175 a_3820_7763# a_4077_7573# a_2882_8007# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4176 a_18907_6706# a_19164_6516# a_17969_6950# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4177 gnd a_24266_2593# a_24058_2593# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4178 a_27985_4209# a_28175_3427# a_28126_3617# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4179 a_7942_6768# a_8926_7065# a_8877_7255# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4180 vdd d4 a_28273_5103# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4181 a_5704_3706# a_5491_3706# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4182 a_25674_6442# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4183 vdd d2 a_3001_1791# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4184 a_6752_2883# a_6539_2883# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4185 a_2004_346# a_1895_346# a_2103_346# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4186 gnd d0 a_24265_3142# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4187 a_5702_7015# a_5489_7015# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4188 a_11834_7259# a_11543_6143# a_11823_6735# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4189 a_12915_2497# a_13172_2307# a_12779_1809# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4190 vdd a_38411_8947# a_38203_8947# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4191 a_5909_7564# a_5488_7564# a_5173_7312# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4192 a_17861_5317# a_17910_2927# a_17861_3117# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4193 gnd a_18086_6249# a_17878_6249# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4194 a_21039_9161# a_20618_9161# a_20302_9042# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4195 a_34040_8675# a_34293_8662# a_33098_9096# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4196 vdd a_18226_7863# a_18018_7863# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4197 a_15206_2718# a_15735_2608# a_15943_2608# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4198 a_1483_2842# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4199 a_1584_7833# a_1371_7833# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4200 a_23069_4679# a_24056_4245# a_24007_4435# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4201 a_119_3775# a_648_3665# a_856_3665# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4202 a_28126_2514# a_29113_2080# a_29068_2093# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4203 a_17968_9156# a_18955_8722# a_18910_8735# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4204 a_32009_6716# a_31588_6716# a_31070_6406# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4205 a_1585_4524# a_1372_4524# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4206 a_6428_4565# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4207 gnd a_19165_7070# a_18957_7070# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4208 a_117_6855# a_646_6974# a_854_6974# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4209 a_37277_373# a_38096_5108# a_38047_5298# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4210 a_13853_5013# a_14110_4823# a_12918_4526# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4211 a_34041_1685# a_34298_1495# a_33106_1198# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4212 a_119_2213# a_120_1756# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4213 a_33103_7816# a_34087_8113# a_34038_8303# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4214 a_38161_2342# a_38414_2329# a_38021_1831# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4215 vdd a_14107_8681# a_13899_8681# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4216 vdd d0 a_24263_7554# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4217 a_23073_5605# a_23326_5592# a_22928_6374# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4218 a_26097_2030# a_26828_2340# a_27036_2340# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4219 a_31072_3097# a_31803_3407# a_32011_3407# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4220 a_10887_910# a_10466_910# a_10151_1115# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4221 a_18909_2294# a_19166_2104# a_17971_2538# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4222 vdd d3 a_3031_2881# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4223 a_29067_8162# a_29063_8339# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4224 a_3822_3351# a_4079_3161# a_2884_3595# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4225 gnd d1 a_18227_5657# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4226 a_25676_2030# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4227 a_21773_1196# a_21560_1196# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4228 a_13852_8322# a_14109_8132# a_12917_7835# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4229 gnd d0 a_24265_4799# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4230 a_15207_1386# a_15736_1505# a_15944_1505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4231 a_31942_6124# a_31729_6124# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4232 gnd a_13171_5616# a_12963_5616# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4233 a_27035_4546# a_26614_4546# a_26097_4790# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4234 gnd a_18088_1837# a_17880_1837# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4235 vdd a_18228_3451# a_18020_3451# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4236 a_25886_8648# a_25673_8648# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4237 a_34042_4263# a_34295_4250# a_33100_4684# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4238 a_1586_3421# a_1373_3421# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4239 a_32020_5040# a_31911_5040# a_32119_5040# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4240 a_17970_4744# a_18957_4310# a_18912_4323# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4241 a_36129_3692# a_35708_3692# a_35392_3573# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4242 gnd d0 a_14108_6475# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4243 a_34038_7200# a_34041_6469# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4244 a_6781_6179# a_6568_6179# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4245 a_20617_8607# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4246 a_7942_6768# a_8926_7065# a_8881_7078# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4247 a_16599_6184# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4248 a_26096_5339# a_25675_5339# a_25360_5544# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4249 a_35390_6652# a_35918_6447# a_36126_6447# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4250 a_23075_1193# a_23328_1180# a_22930_1962# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4251 vdd d0 a_24265_3142# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4252 gnd d0 a_19164_9276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4253 vdd a_14109_4269# a_13901_4269# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4254 a_119_3775# a_119_3546# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4255 a_21981_1196# a_21913_1707# a_21991_2823# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4256 a_2881_9110# a_3138_8920# a_2745_8422# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4257 a_1512_6138# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4258 a_12914_4703# a_13901_4269# a_13852_4459# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4259 a_12805_3076# a_12824_1796# a_12779_1809# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4260 a_1694_5054# a_1481_5054# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4261 a_34036_8852# a_34293_8662# a_33098_9096# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4262 a_16601_1772# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4263 a_29065_8711# a_29061_8888# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4264 a_23069_4679# a_24056_4245# a_24011_4258# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4265 vdd a_19165_7070# a_18957_7070# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4266 a_12919_2320# a_13903_2617# a_13858_2630# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4267 vdd a_9132_8717# a_8924_8717# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4268 gnd d1 a_38412_7844# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4269 vdd a_29319_6492# a_29111_6492# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4270 a_25887_7545# a_25674_7545# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4271 a_25359_6647# a_25360_6190# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4272 a_39101_1549# a_39354_1536# a_38162_1239# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4273 a_27137_368# a_26924_368# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4274 a_5701_6461# a_5488_6461# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4275 a_25888_4236# a_25675_4236# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4276 a_16880_5673# a_16812_6184# a_16890_7300# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4277 a_33103_7816# a_34087_8113# a_34042_8126# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4278 a_15940_7569# a_15519_7569# a_15204_7317# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4279 gnd d0 a_29319_7595# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4280 a_10464_6979# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4281 a_22933_3991# a_23186_3978# a_22964_2875# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4282 a_36130_1486# a_35709_1486# a_35393_1596# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4283 a_38018_8449# a_38203_8947# a_38154_9137# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4284 gnd a_39351_5394# a_39143_5394# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4285 a_30335_4864# a_30864_4754# a_31072_4754# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4286 a_8882_3215# a_9135_3202# a_7940_3636# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4287 a_20618_7504# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4288 a_28123_9132# a_29110_8698# a_29061_8888# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4289 a_35919_8104# a_35706_8104# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4290 a_35391_5092# a_35919_5344# a_36127_5344# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4291 a_26098_927# a_25677_927# a_25362_1132# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4292 gnd a_24263_7554# a_24055_7554# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4293 a_36967_7281# a_36754_7281# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4294 vdd d2 a_33216_6189# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4295 a_35392_2240# a_35920_2035# a_36128_2035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4296 a_12805_5276# a_12854_2886# a_12809_2899# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4297 vdd d1 a_23324_8901# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4298 a_854_8077# a_1584_7833# a_1792_7833# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4299 gnd d0 a_9133_6511# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4300 gnd d0 a_19166_4864# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4301 a_26826_7855# a_26613_7855# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4302 a_34039_2234# a_34045_1508# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4303 a_16457_8982# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4304 gnd d4 a_13062_5086# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4305 a_30333_9276# a_30333_9047# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4306 a_22958_7464# a_22977_6184# a_22928_6374# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4307 vdd a_13171_5616# a_12963_5616# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4308 a_35921_3692# a_35708_3692# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4309 a_31698_7240# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4310 a_34038_4440# a_34295_4250# a_33100_4684# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4311 a_1370_8936# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4312 a_30334_8173# a_30863_8063# a_31071_8063# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4313 gnd d1 a_33356_7803# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4314 a_36126_7550# a_36857_7860# a_37065_7860# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4315 vdd d0 a_14108_6475# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4316 a_5174_6022# a_5703_5912# a_5911_5912# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4317 gnd a_34297_3701# a_34089_3701# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4318 a_20620_3092# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4319 a_25889_3133# a_25676_3133# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4320 a_5172_9102# a_5701_9221# a_5909_9221# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4321 a_646_8077# a_433_8077# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4322 a_118_4649# a_118_4419# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4323 gnd d0 a_29321_3183# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4324 a_15942_3157# a_15521_3157# a_15206_2905# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4325 a_30336_3532# a_30865_3651# a_31073_3651# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4326 a_39098_5407# a_39094_5584# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4327 a_12918_4526# a_13171_4513# a_12778_4015# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4328 a_23071_1370# a_23328_1180# a_22930_1962# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4329 vdd d0 a_19164_9276# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4330 a_21994_7354# a_21697_8325# a_21977_8917# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4331 vdd d3 a_33246_7279# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4332 vdd a_28273_5103# a_28065_5103# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4333 a_5491_3706# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4334 a_28125_4720# a_29112_4286# a_29063_4476# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4335 a_35395_1038# a_35921_932# a_36129_932# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4336 a_28016_3093# a_28035_1813# a_27990_1826# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4337 gnd a_24265_3142# a_24057_3142# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4338 vdd d1 a_23326_4489# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4339 a_856_3665# a_1586_3421# a_1794_3421# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4340 a_18909_3397# a_18914_2671# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4341 a_7060_387# a_7879_5122# a_7830_5312# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4342 a_16459_4570# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4343 a_24008_4989# a_24011_4258# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4344 a_26828_3443# a_26615_3443# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4345 a_10149_5757# a_10149_5527# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4346 a_39097_1726# a_39354_1536# a_38162_1239# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4347 a_1371_7833# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4348 a_38159_7857# a_39143_8154# a_39094_8344# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4349 a_21558_5608# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4350 a_1372_4524# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4351 a_29752_191# d7 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4352 a_36128_3138# a_36859_3448# a_37067_3448# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4353 gnd d1 a_33358_3391# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4354 a_18910_8735# a_18906_8912# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4355 a_32020_5040# a_31700_2828# a_32027_2947# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4356 a_3825_5380# a_4078_5367# a_2883_5801# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4357 a_32010_4510# a_31943_3918# a_32027_2947# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4358 gnd a_3031_5081# a_2823_5081# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4359 a_3821_4454# a_3827_3728# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4360 a_32964_3996# a_33149_4494# a_33100_4684# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4361 vdd a_24263_7554# a_24055_7554# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4362 vdd d0 a_9133_6511# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4363 a_26936_5076# a_26723_5076# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4364 a_22962_7287# a_23215_7274# a_22964_5075# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4365 a_13856_5385# a_13852_5562# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4366 a_20832_5298# a_20619_5298# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4367 vdd d4 a_13062_5086# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4368 gnd a_18227_5657# a_18019_5657# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4369 a_39098_4304# a_39351_4291# a_38156_4725# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4370 a_17969_6950# a_18956_6516# a_18907_6706# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4371 a_22958_7464# a_22977_6184# a_22932_6197# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4372 a_21560_1196# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4373 a_38017_2008# a_38274_1818# a_38047_3098# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4374 a_2882_8007# a_3869_7573# a_3820_7763# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4375 gnd d3 a_18116_7339# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4376 a_6847_8977# a_6780_8385# a_6864_7414# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4377 gnd a_24265_4799# a_24057_4799# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4378 a_13858_2630# a_14111_2617# a_12919_2320# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4379 a_25673_8648# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4380 a_1373_3421# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4381 gnd d0 a_24264_5348# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4382 a_11839_7378# a_11542_8349# a_11822_8941# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4383 gnd a_14108_6475# a_13900_6475# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4384 a_12914_4703# a_13171_4513# a_12778_4015# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4385 a_27037_1237# a_26969_1748# a_27047_2864# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4386 vdd d0 a_29321_3183# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4387 vdd d0 a_4079_4818# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4388 a_15519_9226# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4389 a_26936_7276# a_26723_7276# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4390 a_10149_6173# a_10676_6425# a_10884_6425# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4391 a_853_6420# a_432_6420# a_118_6168# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4392 a_28125_4720# a_29112_4286# a_29067_4299# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4393 gnd d1 a_28382_4530# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4394 vdd a_24265_3142# a_24057_3142# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4395 gnd a_19164_9276# a_18956_9276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4396 a_29965_191# a_29752_191# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4397 vdd d0 a_9135_2099# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4398 a_116_9061# a_645_9180# a_853_9180# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4399 gnd d0 a_34298_1495# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4400 a_22964_2875# a_23217_2862# a_22960_5252# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4401 a_1481_5054# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4402 a_7060_387# a_7879_5122# a_7834_5135# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4403 a_23073_4502# a_24057_4799# a_24012_4812# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4404 gnd a_18229_1245# a_18021_1245# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4405 a_20303_7939# a_20832_8058# a_21040_8058# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4406 a_12777_6221# a_12962_6719# a_12917_6732# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4407 a_38159_7857# a_39143_8154# a_39098_8167# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4408 gnd d3 a_18118_2927# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4409 a_23072_7811# a_23325_7798# a_22927_8580# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4410 a_10883_8631# a_10462_8631# a_10147_8836# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4411 gnd a_38412_7844# a_38204_7844# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4412 a_119_3962# a_119_3775# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4413 a_29068_3196# a_29064_3373# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4414 a_25674_7545# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4415 a_21980_3402# a_21559_3402# a_21042_3646# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4416 a_33105_3404# a_34089_3701# a_34040_3891# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4417 vdd a_3031_5081# a_2823_5081# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4418 a_7943_4562# a_8927_4859# a_8878_5049# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4419 a_25675_4236# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4420 a_25362_1132# a_25364_1033# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4421 gnd d0 a_4079_2058# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4422 a_4632_326# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4423 vdd d1 a_28380_8942# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4424 a_11841_2966# a_11544_3937# a_11824_4529# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4425 gnd d0 a_24266_936# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4426 gnd a_14110_2063# a_13902_2063# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4427 gnd a_39093_9447# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4428 a_10677_8082# a_10464_8082# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4429 a_2886_6727# a_3139_6714# a_2746_6216# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4430 a_8877_4495# a_8883_3769# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4431 a_31941_8330# a_31728_8330# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4432 a_22958_7464# a_23215_7274# a_22964_5075# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4433 a_26099_1481# a_25678_1481# a_25362_1591# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4434 a_10151_1761# a_10678_2013# a_10886_2013# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4435 a_35706_8104# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4436 a_32009_7819# a_31588_7819# a_31071_8063# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4437 a_36754_7281# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4438 a_35390_7111# a_35390_6882# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4439 a_34041_6469# a_34294_6456# a_33099_6890# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4440 a_1585_5627# a_1372_5627# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4441 a_120_1569# a_649_1459# a_857_1459# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4442 a_23070_2473# a_24057_2039# a_24008_2229# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4443 gnd d0 a_14109_8132# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4444 a_2882_8007# a_3869_7573# a_3824_7586# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4445 a_17969_6950# a_18956_6516# a_18911_6529# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4446 a_15205_6027# a_15205_5798# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4447 vdd a_33216_6189# a_33008_6189# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4448 a_36128_5898# a_35707_5898# a_35391_5779# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4449 a_6429_2359# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4450 a_1586_2318# a_1373_2318# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4451 a_11822_8941# a_11401_8941# a_10883_8631# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4452 vdd a_23324_8901# a_23116_8901# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4453 gnd a_9133_6511# a_8925_6511# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4454 gnd a_19166_4864# a_18958_4864# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4455 a_2743_4187# a_3000_3997# a_2778_2894# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4456 a_26613_7855# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4457 gnd a_13062_5086# a_12854_5086# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4458 a_36129_932# a_35708_932# a_35395_1038# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4459 a_21042_2543# a_20621_2543# a_20305_2653# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4460 a_12779_1809# a_12964_2307# a_12919_2320# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4461 a_15203_8877# a_15204_8420# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4462 gnd a_33356_7803# a_33148_7803# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4463 a_23074_3399# a_23327_3386# a_22929_4168# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4464 vdd a_14108_6475# a_13900_6475# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4465 a_27050_7395# a_26753_8366# a_27033_8958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4466 a_25676_3133# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4467 a_15943_3711# a_15522_3711# a_15206_3592# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4468 a_14663_331# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4469 a_5910_7015# a_6640_6771# a_6848_6771# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4470 a_433_8077# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4471 a_37076_7281# a_36967_7281# a_37081_5200# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4472 vdd a_19164_9276# a_18956_9276# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4473 a_12918_4526# a_13902_4823# a_13857_4836# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4474 vdd d1 a_28382_4530# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4475 vdd a_33246_7279# a_33038_7279# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4476 a_13855_9248# a_13851_9425# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4477 a_5700_8667# a_5487_8667# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4478 a_35391_4905# a_35391_4676# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4479 a_31943_3918# a_31730_3918# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4480 a_30336_3948# a_30336_3761# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4481 vdd a_18229_1245# a_18021_1245# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4482 a_32022_2828# a_31731_1712# a_32011_2304# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4483 a_1587_1215# a_1374_1215# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4484 a_34043_2057# a_34296_2044# a_33101_2478# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4485 a_27036_2340# a_26615_2340# a_26098_2584# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4486 a_16879_7879# a_16811_8390# a_16895_7419# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4487 a_17973_7876# a_18226_7863# a_17828_8645# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4488 a_12134_351# a_11713_351# a_11933_5059# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4489 a_17971_2538# a_18958_2104# a_18913_2117# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4490 a_15518_8672# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4491 vdd a_23326_4489# a_23118_4489# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4492 a_8881_5421# a_9134_5408# a_7939_5842# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4493 a_26615_3443# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4494 a_24011_7018# a_24264_7005# a_23072_6708# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4495 a_35390_7298# a_35918_7550# a_36126_7550# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4496 vdd d2 a_33215_8395# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4497 gnd a_33358_3391# a_33150_3391# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4498 gnd d0 a_9132_8717# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4499 a_1795_1215# a_1727_1726# a_1805_2842# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4500 vdd a_14110_2063# a_13902_2063# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4501 a_5172_9331# a_5172_9102# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4502 a_37065_7860# a_36997_8371# a_37081_7400# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4503 a_2882_6904# a_3139_6714# a_2746_6216# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4504 a_27052_2983# a_26755_3954# a_27035_4546# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4505 a_34037_6646# a_34294_6456# a_33099_6890# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4506 vdd d2 a_33218_1777# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4507 vdd d0 a_14109_8132# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4508 vdd a_9133_6511# a_8925_6511# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4509 a_20833_5852# a_20620_5852# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4510 a_26723_5076# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4511 a_11841_2966# a_11727_2847# a_11834_5059# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4512 a_5701_7564# a_5488_7564# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4513 a_25888_5339# a_25675_5339# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4514 vdd a_13062_5086# a_12854_5086# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4515 a_5702_4255# a_5489_4255# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4516 a_20831_9161# a_20618_9161# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4517 a_856_2562# a_435_2562# a_119_2672# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4518 a_8876_9461# a_8879_8730# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4519 gnd a_18116_7339# a_17908_7339# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4520 a_30335_5738# a_30864_5857# a_31072_5857# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4521 gnd d0 a_29320_5389# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4522 a_12917_6732# a_13170_6719# a_12777_6221# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4523 a_31801_6716# a_31588_6716# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4524 a_30336_2658# a_30865_2548# a_31073_2548# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4525 a_23070_3576# a_23327_3386# a_22929_4168# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4526 a_20619_5298# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4527 a_8883_1009# a_9136_996# a_7941_1430# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4528 a_29067_7059# a_29063_7236# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4529 a_16890_7300# a_16599_6184# a_16880_5673# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4530 a_8879_3946# a_8882_3215# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4531 a_35392_2886# a_35920_3138# a_36128_3138# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4532 vdd d0 a_29322_3737# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4533 gnd a_24264_5348# a_24056_5348# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4534 vdd d1 a_23325_6695# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4535 a_855_5871# a_1585_5627# a_1793_5627# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4536 a_20305_3297# a_20833_3092# a_21041_3092# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4537 a_6640_7874# a_6427_7874# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4538 a_16458_6776# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4539 a_26827_5649# a_26614_5649# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4540 a_26723_7276# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4541 a_21880_7235# a_21667_7235# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4542 a_2772_7483# a_2791_6203# a_2742_6393# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4543 a_28129_4543# a_29113_4840# a_29068_4853# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4544 a_22964_2875# a_22978_3978# a_22929_4168# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4545 a_35922_1486# a_35709_1486# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4546 a_7940_3636# a_8927_3202# a_8878_3392# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4547 a_34039_2234# a_34296_2044# a_33101_2478# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4548 a_26825_8958# a_26612_8958# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4549 gnd d1 a_33357_5597# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4550 a_20835_1440# a_20622_1440# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4551 vdd a_9135_2099# a_8927_2099# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4552 a_5703_3152# a_5490_3152# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4553 gnd a_34298_1495# a_34090_1495# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4554 a_6866_3002# a_6752_2883# a_6859_5095# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4555 a_18907_9466# a_18910_8735# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4556 a_5173_6896# a_5702_7015# a_5910_7015# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4557 a_30337_1326# a_30866_1445# a_31074_1445# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4558 gnd d0 a_29322_977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4559 gnd a_18118_2927# a_17910_2927# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4560 a_3822_6111# a_4079_5921# a_2887_5624# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4561 a_31803_2304# a_31590_2304# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4562 gnd d0 a_4080_2612# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4563 a_21989_7235# a_21698_6119# a_21978_6711# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4564 a_39097_6510# a_39350_6497# a_38155_6931# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4565 a_3823_1145# a_122_1011# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4566 a_15207_1802# a_15734_2054# a_15942_2054# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4567 gnd a_24266_936# a_24058_936# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4568 vdd d1 a_3140_4508# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4569 a_16459_5673# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4570 a_857_1459# a_1587_1215# a_1795_1215# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4571 a_10464_8082# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4572 a_6642_3462# a_6429_3462# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4573 a_26829_1237# a_26616_1237# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4574 a_25677_927# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4575 a_5909_9221# a_5488_9221# a_5172_9331# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4576 a_12778_4015# a_12963_4513# a_12914_4703# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4577 a_1372_5627# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4578 a_38160_5651# a_39144_5948# a_39095_6138# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4579 a_1373_2318# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4580 a_31070_9166# a_30649_9166# a_30333_9047# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4581 a_21043_1440# a_21773_1196# a_21981_1196# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4582 a_852_8626# a_431_8626# a_117_8374# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4583 a_35391_6195# a_35391_6008# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4584 vdd d0 a_24265_5902# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4585 gnd d1 a_28381_6736# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4586 a_21041_3092# a_20620_3092# a_20305_3297# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4587 vdd d0 a_9134_4305# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4588 a_39100_995# a_39096_1172# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4589 a_10678_4773# a_10465_4773# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4590 a_39099_2098# a_39352_2085# a_38157_2519# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4591 a_12776_8427# a_12961_8925# a_12916_8938# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4592 a_31913_2828# a_31700_2828# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4593 a_6848_6771# a_6781_6179# a_6859_7295# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4594 a_38045_7510# a_38064_6230# a_38015_6420# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4595 a_16880_4570# a_16459_4570# a_15941_4260# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4596 a_31730_3918# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4597 gnd d1 a_13170_7822# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4598 a_1374_1215# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4599 gnd a_14109_4269# a_13901_4269# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
C0 a_37175_5081# a_37277_373# 8.08fF
C1 a_16989_5100# a_17091_392# 8.08fF
C2 a_1902_5054# a_2004_346# 8.08fF
C3 a_22088_5035# a_22190_327# 8.08fF
C4 a_32119_5040# a_32221_332# 8.08fF
C5 a_11933_5059# a_12035_351# 8.08fF
C6 vdd d2 2.11fF
C7 a_25239_307# a_25140_307# 3.47fF
C8 vdd d0 8.45fF
C9 a_6958_5095# a_7060_387# 8.08fF
C10 a_5053_326# a_4954_326# 3.47fF
C11 a_27144_5076# a_27246_368# 8.08fF
C12 vdd d1 4.22fF
C13 a_35171_312# gnd 3.40fF
C14 a_30074_191# gnd 6.50fF
C15 a_32320_332# gnd 4.59fF
C16 d5 gnd 2.50fF
C17 a_25140_307# gnd 3.40fF
C18 a_25239_307# gnd 7.14fF
C19 a_22289_327# gnd 4.59fF
C20 a_14985_331# gnd 3.40fF
C21 a_9888_210# gnd 6.50fF
C22 a_9987_210# gnd 11.31fF
C23 a_12134_351# gnd 4.59fF
C24 a_4954_326# gnd 3.40fF
C25 a_5053_326# gnd 7.14fF
C26 a_2103_346# gnd 4.59fF
C27 a_39096_1172# gnd 2.22fF
C28 a_35395_1038# gnd 6.43fF
C29 d0 gnd 95.26fF
C30 a_34040_1131# gnd 2.22fF
C31 a_30339_997# gnd 6.43fF
C32 a_39100_995# gnd 2.38fF
C33 a_35393_1137# gnd 2.23fF
C34 a_34044_954# gnd 2.38fF
C35 a_38158_1416# gnd 2.38fF
C36 d1 gnd 49.89fF
C37 a_36129_932# gnd 2.52fF
C38 a_29065_1167# gnd 2.22fF
C39 a_25364_1033# gnd 6.43fF
C40 a_24009_1126# gnd 2.22fF
C41 a_20308_992# gnd 6.43fF
C42 a_30337_1096# gnd 2.23fF
C43 a_33102_1375# gnd 2.38fF
C44 a_31073_891# gnd 2.52fF
C45 a_29069_990# gnd 2.38fF
C46 a_25362_1132# gnd 2.23fF
C47 a_24013_949# gnd 2.38fF
C48 a_35393_1367# gnd 2.38fF
C49 a_36130_1486# gnd 2.18fF
C50 a_28127_1411# gnd 2.38fF
C51 a_26098_927# gnd 2.52fF
C52 a_20306_1091# gnd 2.23fF
C53 a_18910_1191# gnd 2.22fF
C54 a_15209_1057# gnd 6.43fF
C55 a_13854_1150# gnd 2.22fF
C56 a_10153_1016# gnd 6.43fF
C57 a_23071_1370# gnd 2.38fF
C58 a_21042_886# gnd 2.52fF
C59 a_18914_1014# gnd 2.38fF
C60 a_35393_1596# gnd 2.28fF
C61 a_30337_1326# gnd 2.38fF
C62 a_31074_1445# gnd 2.18fF
C63 a_30337_1555# gnd 2.28fF
C64 a_38162_1239# gnd 2.52fF
C65 a_39097_1726# gnd 2.23fF
C66 a_33106_1198# gnd 2.52fF
C67 a_34041_1685# gnd 2.23fF
C68 a_25362_1362# gnd 2.38fF
C69 a_26099_1481# gnd 2.18fF
C70 a_15207_1156# gnd 2.23fF
C71 a_13858_973# gnd 2.38fF
C72 a_17972_1435# gnd 2.38fF
C73 a_15943_951# gnd 2.52fF
C74 a_8879_1186# gnd 2.22fF
C75 a_5178_1052# gnd 6.43fF
C76 a_3823_1145# gnd 2.22fF
C77 a_122_1011# gnd 6.43fF
C78 a_10151_1115# gnd 2.23fF
C79 a_12916_1394# gnd 2.38fF
C80 a_10887_910# gnd 2.52fF
C81 a_8883_1009# gnd 2.38fF
C82 a_5176_1151# gnd 2.23fF
C83 a_3827_968# gnd 2.38fF
C84 a_25362_1591# gnd 2.28fF
C85 a_20306_1321# gnd 2.38fF
C86 a_21043_1440# gnd 2.18fF
C87 a_20306_1550# gnd 2.28fF
C88 a_39101_1549# gnd 2.49fF
C89 a_28131_1234# gnd 2.52fF
C90 a_29066_1721# gnd 2.23fF
C91 a_23075_1193# gnd 2.52fF
C92 a_24010_1680# gnd 2.23fF
C93 d2 gnd 25.13fF
C94 a_34045_1508# gnd 2.49fF
C95 a_29070_1544# gnd 2.49fF
C96 a_15207_1386# gnd 2.38fF
C97 a_15944_1505# gnd 2.18fF
C98 a_7941_1430# gnd 2.38fF
C99 a_5912_946# gnd 2.52fF
C100 a_120_1110# gnd 2.23fF
C101 a_2885_1389# gnd 2.38fF
C102 a_856_905# gnd 2.52fF
C103 a_15207_1615# gnd 2.28fF
C104 a_10151_1345# gnd 2.38fF
C105 a_10888_1464# gnd 2.18fF
C106 a_10151_1574# gnd 2.28fF
C107 a_17976_1258# gnd 2.52fF
C108 a_18911_1745# gnd 2.23fF
C109 a_12920_1217# gnd 2.52fF
C110 a_13855_1704# gnd 2.23fF
C111 a_5176_1381# gnd 2.38fF
C112 a_5913_1500# gnd 2.18fF
C113 a_5176_1610# gnd 2.28fF
C114 a_120_1340# gnd 2.38fF
C115 a_857_1459# gnd 2.18fF
C116 a_120_1569# gnd 2.28fF
C117 a_24014_1503# gnd 2.49fF
C118 a_39095_2275# gnd 2.28fF
C119 a_35393_1783# gnd 2.49fF
C120 a_34039_2234# gnd 2.28fF
C121 a_30337_1742# gnd 2.49fF
C122 a_39099_2098# gnd 2.38fF
C123 a_35392_2240# gnd 2.23fF
C124 a_34043_2057# gnd 2.38fF
C125 a_38157_2519# gnd 2.18fF
C126 a_36128_2035# gnd 2.52fF
C127 a_29064_2270# gnd 2.28fF
C128 a_25362_1778# gnd 2.49fF
C129 a_18915_1568# gnd 2.49fF
C130 a_7945_1253# gnd 2.52fF
C131 a_8880_1740# gnd 2.23fF
C132 a_2889_1212# gnd 2.52fF
C133 a_3824_1699# gnd 2.23fF
C134 a_13859_1527# gnd 2.49fF
C135 a_24008_2229# gnd 2.28fF
C136 a_20306_1737# gnd 2.49fF
C137 a_8884_1563# gnd 2.49fF
C138 a_3828_1522# gnd 2.49fF
C139 a_30336_2199# gnd 2.23fF
C140 a_33101_2478# gnd 2.18fF
C141 a_31072_1994# gnd 2.52fF
C142 a_29068_2093# gnd 2.38fF
C143 a_25361_2235# gnd 2.23fF
C144 a_24012_2052# gnd 2.38fF
C145 a_35392_2470# gnd 2.38fF
C146 a_36129_2589# gnd 2.45fF
C147 a_28126_2514# gnd 2.18fF
C148 a_26097_2030# gnd 2.52fF
C149 a_20305_2194# gnd 2.23fF
C150 a_18909_2294# gnd 2.28fF
C151 a_15207_1802# gnd 2.49fF
C152 a_13853_2253# gnd 2.28fF
C153 a_10151_1761# gnd 2.49fF
C154 a_23070_2473# gnd 2.18fF
C155 a_21041_1989# gnd 2.52fF
C156 a_18913_2117# gnd 2.38fF
C157 a_35392_2699# gnd 2.28fF
C158 a_30336_2429# gnd 2.38fF
C159 a_31073_2548# gnd 2.45fF
C160 a_30336_2658# gnd 2.28fF
C161 a_38161_2342# gnd 2.52fF
C162 a_39096_2829# gnd 2.23fF
C163 a_33105_2301# gnd 2.52fF
C164 a_34040_2788# gnd 2.23fF
C165 a_25361_2465# gnd 2.38fF
C166 a_26098_2584# gnd 2.45fF
C167 a_15206_2259# gnd 2.23fF
C168 a_13857_2076# gnd 2.38fF
C169 a_17971_2538# gnd 2.18fF
C170 a_15942_2054# gnd 2.52fF
C171 a_8878_2289# gnd 2.28fF
C172 a_5176_1797# gnd 2.49fF
C173 a_3822_2248# gnd 2.28fF
C174 a_120_1756# gnd 2.49fF
C175 a_10150_2218# gnd 2.23fF
C176 a_12915_2497# gnd 2.18fF
C177 a_10886_2013# gnd 2.52fF
C178 a_8882_2112# gnd 2.38fF
C179 a_5175_2254# gnd 2.23fF
C180 a_3826_2071# gnd 2.38fF
C181 a_25361_2694# gnd 2.28fF
C182 a_20305_2424# gnd 2.38fF
C183 a_21042_2543# gnd 2.45fF
C184 a_20305_2653# gnd 2.28fF
C185 a_28130_2337# gnd 2.52fF
C186 a_29065_2824# gnd 2.23fF
C187 a_23074_2296# gnd 2.52fF
C188 a_24009_2783# gnd 2.23fF
C189 a_15206_2489# gnd 2.38fF
C190 a_15943_2608# gnd 2.45fF
C191 a_7940_2533# gnd 2.18fF
C192 a_5911_2049# gnd 2.52fF
C193 a_119_2213# gnd 2.23fF
C194 a_2884_2492# gnd 2.18fF
C195 a_855_2008# gnd 2.52fF
C196 a_15206_2718# gnd 2.28fF
C197 a_10150_2448# gnd 2.38fF
C198 a_10887_2567# gnd 2.45fF
C199 a_10150_2677# gnd 2.28fF
C200 a_37078_2869# gnd 2.28fF
C201 a_32022_2828# gnd 2.28fF
C202 a_17975_2361# gnd 2.52fF
C203 a_18910_2848# gnd 2.23fF
C204 a_39100_2652# gnd 2.49fF
C205 d3 gnd 11.35fF
C206 a_34044_2611# gnd 2.49fF
C207 a_38047_3098# gnd 2.04fF
C208 a_32991_3057# gnd 2.04fF
C209 a_27047_2864# gnd 2.28fF
C210 a_21991_2823# gnd 2.28fF
C211 a_12919_2320# gnd 2.52fF
C212 a_13854_2807# gnd 2.23fF
C213 a_5175_2484# gnd 2.38fF
C214 a_5912_2603# gnd 2.45fF
C215 a_5175_2713# gnd 2.28fF
C216 a_119_2443# gnd 2.38fF
C217 a_856_2562# gnd 2.45fF
C218 a_119_2672# gnd 2.28fF
C219 a_29069_2647# gnd 2.49fF
C220 a_39095_3378# gnd 2.28fF
C221 a_35392_2886# gnd 2.49fF
C222 a_24013_2606# gnd 2.49fF
C223 a_28016_3093# gnd 2.04fF
C224 a_7944_2356# gnd 2.52fF
C225 a_8879_2843# gnd 2.23fF
C226 a_2888_2315# gnd 2.52fF
C227 a_3823_2802# gnd 2.23fF
C228 a_22960_3052# gnd 2.04fF
C229 a_16892_2888# gnd 2.28fF
C230 a_11836_2847# gnd 2.28fF
C231 a_34039_3337# gnd 2.28fF
C232 a_30336_2845# gnd 2.49fF
C233 a_39099_3201# gnd 2.38fF
C234 a_35392_3343# gnd 2.23fF
C235 a_34043_3160# gnd 2.38fF
C236 a_38157_3622# gnd 2.45fF
C237 a_36128_3138# gnd 2.52fF
C238 a_29064_3373# gnd 2.28fF
C239 a_25361_2881# gnd 2.49fF
C240 a_18914_2671# gnd 2.49fF
C241 a_24008_3332# gnd 2.28fF
C242 a_20305_2840# gnd 2.49fF
C243 a_13858_2630# gnd 2.49fF
C244 a_17861_3117# gnd 2.04fF
C245 a_12805_3076# gnd 2.04fF
C246 a_6861_2883# gnd 2.28fF
C247 a_1805_2842# gnd 2.28fF
C248 a_8883_2666# gnd 2.49fF
C249 a_30336_3302# gnd 2.23fF
C250 a_33101_3581# gnd 2.45fF
C251 a_31072_3097# gnd 2.52fF
C252 a_29068_3196# gnd 2.38fF
C253 a_25361_3338# gnd 2.23fF
C254 a_24012_3155# gnd 2.38fF
C255 a_35392_3573# gnd 2.38fF
C256 a_36129_3692# gnd 2.18fF
C257 a_28126_3617# gnd 2.45fF
C258 a_26097_3133# gnd 2.52fF
C259 a_20305_3297# gnd 2.23fF
C260 a_18909_3397# gnd 2.28fF
C261 a_15206_2905# gnd 2.49fF
C262 a_3827_2625# gnd 2.49fF
C263 a_7830_3112# gnd 2.04fF
C264 a_2774_3071# gnd 2.04fF
C265 a_13853_3356# gnd 2.28fF
C266 a_10150_2864# gnd 2.49fF
C267 a_23070_3576# gnd 2.45fF
C268 a_21041_3092# gnd 2.52fF
C269 a_18913_3220# gnd 2.38fF
C270 a_35392_3802# gnd 2.28fF
C271 a_30336_3532# gnd 2.38fF
C272 a_31073_3651# gnd 2.18fF
C273 a_30336_3761# gnd 2.28fF
C274 a_38161_3445# gnd 2.52fF
C275 a_39096_3932# gnd 2.23fF
C276 a_33105_3404# gnd 2.52fF
C277 a_34040_3891# gnd 2.23fF
C278 a_25361_3568# gnd 2.38fF
C279 a_26098_3687# gnd 2.18fF
C280 a_15206_3362# gnd 2.23fF
C281 a_13857_3179# gnd 2.38fF
C282 a_17971_3641# gnd 2.45fF
C283 a_15942_3157# gnd 2.52fF
C284 a_8878_3392# gnd 2.28fF
C285 a_5175_2900# gnd 2.49fF
C286 a_3822_3351# gnd 2.28fF
C287 a_119_2859# gnd 2.49fF
C288 a_10150_3321# gnd 2.23fF
C289 a_12915_3600# gnd 2.45fF
C290 a_10886_3116# gnd 2.52fF
C291 a_8882_3215# gnd 2.38fF
C292 a_5175_3357# gnd 2.23fF
C293 a_3826_3174# gnd 2.38fF
C294 a_25361_3797# gnd 2.28fF
C295 a_20305_3527# gnd 2.38fF
C296 a_21042_3646# gnd 2.18fF
C297 a_20305_3756# gnd 2.28fF
C298 a_39100_3755# gnd 2.49fF
C299 a_37083_2988# gnd 2.45fF
C300 a_28130_3440# gnd 2.52fF
C301 a_29065_3927# gnd 2.23fF
C302 a_23074_3399# gnd 2.52fF
C303 a_24009_3886# gnd 2.23fF
C304 a_34044_3714# gnd 2.49fF
C305 a_32027_2947# gnd 2.45fF
C306 a_38051_2921# gnd 2.34fF
C307 a_32995_2880# gnd 2.34fF
C308 a_29069_3750# gnd 2.49fF
C309 a_27052_2983# gnd 2.45fF
C310 a_15206_3592# gnd 2.38fF
C311 a_15943_3711# gnd 2.18fF
C312 a_7940_3636# gnd 2.45fF
C313 a_5911_3152# gnd 2.52fF
C314 a_119_3316# gnd 2.23fF
C315 a_2884_3595# gnd 2.45fF
C316 a_855_3111# gnd 2.52fF
C317 a_15206_3821# gnd 2.28fF
C318 a_10150_3551# gnd 2.38fF
C319 a_10887_3670# gnd 2.18fF
C320 a_10150_3780# gnd 2.28fF
C321 a_17975_3464# gnd 2.52fF
C322 a_18910_3951# gnd 2.23fF
C323 a_12919_3423# gnd 2.52fF
C324 a_13854_3910# gnd 2.23fF
C325 a_5175_3587# gnd 2.38fF
C326 a_5912_3706# gnd 2.18fF
C327 a_5175_3816# gnd 2.28fF
C328 a_119_3546# gnd 2.38fF
C329 a_856_3665# gnd 2.18fF
C330 a_119_3775# gnd 2.28fF
C331 a_24013_3709# gnd 2.49fF
C332 a_21996_2942# gnd 2.45fF
C333 a_39094_4481# gnd 2.28fF
C334 a_35392_3989# gnd 2.49fF
C335 a_28020_2916# gnd 2.34fF
C336 a_22964_2875# gnd 2.34fF
C337 a_34038_4440# gnd 2.28fF
C338 a_30336_3948# gnd 2.49fF
C339 a_39098_4304# gnd 2.38fF
C340 a_35391_4446# gnd 2.23fF
C341 a_34042_4263# gnd 2.38fF
C342 a_38156_4725# gnd 2.18fF
C343 a_36127_4241# gnd 2.52fF
C344 a_29063_4476# gnd 2.28fF
C345 a_25361_3984# gnd 2.49fF
C346 a_18914_3774# gnd 2.49fF
C347 a_16897_3007# gnd 2.45fF
C348 a_7944_3459# gnd 2.52fF
C349 a_8879_3946# gnd 2.23fF
C350 a_2888_3418# gnd 2.52fF
C351 a_3823_3905# gnd 2.23fF
C352 a_13858_3733# gnd 2.49fF
C353 a_11841_2966# gnd 2.45fF
C354 a_24007_4435# gnd 2.28fF
C355 a_20305_3943# gnd 2.49fF
C356 a_17865_2940# gnd 2.34fF
C357 a_12809_2899# gnd 2.34fF
C358 a_8883_3769# gnd 2.49fF
C359 a_6866_3002# gnd 2.45fF
C360 a_3827_3728# gnd 2.49fF
C361 a_1810_2961# gnd 2.45fF
C362 a_30335_4405# gnd 2.23fF
C363 a_33100_4684# gnd 2.18fF
C364 a_31071_4200# gnd 2.52fF
C365 a_29067_4299# gnd 2.38fF
C366 a_25360_4441# gnd 2.23fF
C367 a_24011_4258# gnd 2.38fF
C368 a_35391_4676# gnd 2.38fF
C369 a_36128_4795# gnd 2.45fF
C370 a_28125_4720# gnd 2.18fF
C371 a_26096_4236# gnd 2.52fF
C372 a_20304_4400# gnd 2.23fF
C373 a_18908_4500# gnd 2.28fF
C374 a_15206_4008# gnd 2.49fF
C375 a_7834_2935# gnd 2.34fF
C376 a_2778_2894# gnd 2.34fF
C377 a_13852_4459# gnd 2.28fF
C378 a_10150_3967# gnd 2.49fF
C379 a_23069_4679# gnd 2.18fF
C380 a_21040_4195# gnd 2.52fF
C381 a_18912_4323# gnd 2.38fF
C382 a_35391_4905# gnd 2.28fF
C383 a_30335_4635# gnd 2.38fF
C384 a_31072_4754# gnd 2.45fF
C385 a_30335_4864# gnd 2.28fF
C386 a_38160_4548# gnd 2.52fF
C387 a_39095_5035# gnd 2.23fF
C388 a_33104_4507# gnd 2.52fF
C389 a_34039_4994# gnd 2.23fF
C390 a_25360_4671# gnd 2.38fF
C391 a_26097_4790# gnd 2.45fF
C392 a_15205_4465# gnd 2.23fF
C393 a_13856_4282# gnd 2.38fF
C394 a_17970_4744# gnd 2.18fF
C395 a_15941_4260# gnd 2.52fF
C396 a_8877_4495# gnd 2.28fF
C397 a_5175_4003# gnd 2.49fF
C398 a_3821_4454# gnd 2.28fF
C399 a_119_3962# gnd 2.49fF
C400 a_10149_4424# gnd 2.23fF
C401 a_12914_4703# gnd 2.18fF
C402 a_10885_4219# gnd 2.52fF
C403 a_8881_4318# gnd 2.38fF
C404 a_5174_4460# gnd 2.23fF
C405 a_3825_4277# gnd 2.38fF
C406 a_25360_4900# gnd 2.28fF
C407 a_20304_4630# gnd 2.38fF
C408 a_21041_4749# gnd 2.45fF
C409 a_20304_4859# gnd 2.28fF
C410 a_28129_4543# gnd 2.52fF
C411 a_29064_5030# gnd 2.23fF
C412 a_39099_4858# gnd 2.50fF
C413 a_37277_373# gnd 6.48fF
C414 a_37076_5081# gnd 3.68fF
C415 a_37175_5081# gnd 5.48fF
C416 d4 gnd 5.88fF
C417 a_34043_4817# gnd 2.50fF
C418 a_38047_5298# gnd 3.32fF
C419 a_32221_332# gnd 6.48fF
C420 a_32020_5040# gnd 3.68fF
C421 a_32119_5040# gnd 5.48fF
C422 a_23073_4502# gnd 2.52fF
C423 a_24008_4989# gnd 2.23fF
C424 a_15205_4695# gnd 2.38fF
C425 a_15942_4814# gnd 2.45fF
C426 a_7939_4739# gnd 2.18fF
C427 a_5910_4255# gnd 2.52fF
C428 a_118_4419# gnd 2.23fF
C429 a_2883_4698# gnd 2.18fF
C430 a_854_4214# gnd 2.52fF
C431 a_15205_4924# gnd 2.28fF
C432 a_10149_4654# gnd 2.38fF
C433 a_10886_4773# gnd 2.45fF
C434 a_10149_4883# gnd 2.28fF
C435 a_17974_4567# gnd 2.52fF
C436 a_18909_5054# gnd 2.23fF
C437 a_32991_5257# gnd 3.32fF
C438 a_29068_4853# gnd 2.50fF
C439 a_39094_5584# gnd 2.28fF
C440 a_35391_5092# gnd 2.50fF
C441 a_27246_368# gnd 6.48fF
C442 a_27045_5076# gnd 3.68fF
C443 a_27144_5076# gnd 5.48fF
C444 a_24012_4812# gnd 2.50fF
C445 a_28016_5293# gnd 3.32fF
C446 a_22190_327# gnd 6.48fF
C447 a_21989_5035# gnd 3.68fF
C448 a_22088_5035# gnd 5.48fF
C449 a_12918_4526# gnd 2.52fF
C450 a_13853_5013# gnd 2.23fF
C451 a_5174_4690# gnd 2.38fF
C452 a_5911_4809# gnd 2.45fF
C453 a_5174_4919# gnd 2.28fF
C454 a_118_4649# gnd 2.38fF
C455 a_855_4768# gnd 2.45fF
C456 a_118_4878# gnd 2.28fF
C457 a_7943_4562# gnd 2.52fF
C458 a_8878_5049# gnd 2.23fF
C459 a_22960_5252# gnd 3.32fF
C460 a_34038_5543# gnd 2.28fF
C461 a_30335_5051# gnd 2.50fF
C462 a_39098_5407# gnd 2.38fF
C463 a_35391_5549# gnd 2.23fF
C464 a_34042_5366# gnd 2.38fF
C465 a_38156_5828# gnd 2.45fF
C466 a_36127_5344# gnd 2.52fF
C467 a_29063_5579# gnd 2.28fF
C468 a_25360_5087# gnd 2.50fF
C469 a_18913_4877# gnd 2.50fF
C470 a_24007_5538# gnd 2.28fF
C471 a_20304_5046# gnd 2.50fF
C472 a_17091_392# gnd 6.48fF
C473 a_16890_5100# gnd 3.68fF
C474 a_16989_5100# gnd 5.48fF
C475 a_13857_4836# gnd 2.50fF
C476 a_17861_5317# gnd 3.32fF
C477 a_12035_351# gnd 6.48fF
C478 a_11834_5059# gnd 3.68fF
C479 a_11933_5059# gnd 5.48fF
C480 a_2887_4521# gnd 2.52fF
C481 a_3822_5008# gnd 2.23fF
C482 a_12805_5276# gnd 3.32fF
C483 a_8882_4872# gnd 2.50fF
C484 a_30335_5508# gnd 2.23fF
C485 a_33100_5787# gnd 2.45fF
C486 a_31071_5303# gnd 2.52fF
C487 a_29067_5402# gnd 2.38fF
C488 a_25360_5544# gnd 2.23fF
C489 a_24011_5361# gnd 2.38fF
C490 a_35391_5779# gnd 2.38fF
C491 a_36128_5898# gnd 2.18fF
C492 a_28125_5823# gnd 2.45fF
C493 a_26096_5339# gnd 2.52fF
C494 a_20304_5503# gnd 2.23fF
C495 a_18908_5603# gnd 2.28fF
C496 a_15205_5111# gnd 2.50fF
C497 a_7060_387# gnd 6.48fF
C498 a_6859_5095# gnd 3.68fF
C499 a_6958_5095# gnd 5.48fF
C500 a_3826_4831# gnd 2.50fF
C501 a_7830_5312# gnd 3.32fF
C502 a_2004_346# gnd 6.48fF
C503 a_1803_5054# gnd 3.68fF
C504 a_1902_5054# gnd 5.48fF
C505 a_2774_5271# gnd 3.32fF
C506 a_13852_5562# gnd 2.28fF
C507 a_10149_5070# gnd 2.50fF
C508 a_23069_5782# gnd 2.45fF
C509 a_21040_5298# gnd 2.52fF
C510 a_18912_5426# gnd 2.38fF
C511 a_35391_6008# gnd 2.28fF
C512 a_30335_5738# gnd 2.38fF
C513 a_31072_5857# gnd 2.18fF
C514 a_30335_5967# gnd 2.28fF
C515 a_38160_5651# gnd 2.52fF
C516 a_39095_6138# gnd 2.23fF
C517 a_33104_5610# gnd 2.52fF
C518 a_34039_6097# gnd 2.23fF
C519 a_25360_5774# gnd 2.38fF
C520 a_26097_5893# gnd 2.18fF
C521 a_15205_5568# gnd 2.23fF
C522 a_13856_5385# gnd 2.38fF
C523 a_17970_5847# gnd 2.45fF
C524 a_15941_5363# gnd 2.52fF
C525 a_8877_5598# gnd 2.28fF
C526 a_5174_5106# gnd 2.50fF
C527 a_3821_5557# gnd 2.28fF
C528 a_118_5065# gnd 2.50fF
C529 a_10149_5527# gnd 2.23fF
C530 a_12914_5806# gnd 2.45fF
C531 a_10885_5322# gnd 2.52fF
C532 a_8881_5421# gnd 2.38fF
C533 a_5174_5563# gnd 2.23fF
C534 a_3825_5380# gnd 2.38fF
C535 a_25360_6003# gnd 2.28fF
C536 a_20304_5733# gnd 2.38fF
C537 a_21041_5852# gnd 2.18fF
C538 a_20304_5962# gnd 2.28fF
C539 a_39099_5961# gnd 2.49fF
C540 a_28129_5646# gnd 2.52fF
C541 a_29064_6133# gnd 2.23fF
C542 a_23073_5605# gnd 2.52fF
C543 a_24008_6092# gnd 2.23fF
C544 a_34043_5920# gnd 2.49fF
C545 a_29068_5956# gnd 2.49fF
C546 a_15205_5798# gnd 2.38fF
C547 a_15942_5917# gnd 2.18fF
C548 a_7939_5842# gnd 2.45fF
C549 a_5910_5358# gnd 2.52fF
C550 a_118_5522# gnd 2.23fF
C551 a_2883_5801# gnd 2.45fF
C552 a_854_5317# gnd 2.52fF
C553 a_15205_6027# gnd 2.28fF
C554 a_10149_5757# gnd 2.38fF
C555 a_10886_5876# gnd 2.18fF
C556 a_10149_5986# gnd 2.28fF
C557 a_17974_5670# gnd 2.52fF
C558 a_18909_6157# gnd 2.23fF
C559 a_12918_5629# gnd 2.52fF
C560 a_13853_6116# gnd 2.23fF
C561 a_5174_5793# gnd 2.38fF
C562 a_5911_5912# gnd 2.18fF
C563 a_5174_6022# gnd 2.28fF
C564 a_118_5752# gnd 2.38fF
C565 a_855_5871# gnd 2.18fF
C566 a_118_5981# gnd 2.28fF
C567 a_24012_5915# gnd 2.49fF
C568 a_39093_6687# gnd 2.28fF
C569 a_35391_6195# gnd 2.49fF
C570 a_34037_6646# gnd 2.28fF
C571 a_30335_6154# gnd 2.49fF
C572 a_39097_6510# gnd 2.38fF
C573 a_35390_6652# gnd 2.23fF
C574 a_34041_6469# gnd 2.38fF
C575 a_38155_6931# gnd 2.18fF
C576 a_36126_6447# gnd 2.52fF
C577 a_29062_6682# gnd 2.28fF
C578 a_25360_6190# gnd 2.49fF
C579 a_18913_5980# gnd 2.49fF
C580 a_7943_5665# gnd 2.52fF
C581 a_8878_6152# gnd 2.23fF
C582 a_2887_5624# gnd 2.52fF
C583 a_3822_6111# gnd 2.23fF
C584 a_13857_5939# gnd 2.49fF
C585 a_24006_6641# gnd 2.28fF
C586 a_20304_6149# gnd 2.49fF
C587 a_8882_5975# gnd 2.49fF
C588 a_3826_5934# gnd 2.49fF
C589 a_30334_6611# gnd 2.23fF
C590 a_33099_6890# gnd 2.18fF
C591 a_31070_6406# gnd 2.52fF
C592 a_29066_6505# gnd 2.38fF
C593 a_25359_6647# gnd 2.23fF
C594 a_24010_6464# gnd 2.38fF
C595 a_35390_6882# gnd 2.38fF
C596 a_36127_7001# gnd 2.45fF
C597 a_28124_6926# gnd 2.18fF
C598 a_26095_6442# gnd 2.52fF
C599 a_20303_6606# gnd 2.23fF
C600 a_18907_6706# gnd 2.28fF
C601 a_15205_6214# gnd 2.49fF
C602 a_13851_6665# gnd 2.28fF
C603 a_10149_6173# gnd 2.49fF
C604 a_23068_6885# gnd 2.18fF
C605 a_21039_6401# gnd 2.52fF
C606 a_18911_6529# gnd 2.38fF
C607 a_35390_7111# gnd 2.28fF
C608 a_30334_6841# gnd 2.38fF
C609 a_31071_6960# gnd 2.45fF
C610 a_30334_7070# gnd 2.28fF
C611 a_38159_6754# gnd 2.52fF
C612 a_39094_7241# gnd 2.23fF
C613 a_33103_6713# gnd 2.52fF
C614 a_34038_7200# gnd 2.23fF
C615 a_25359_6877# gnd 2.38fF
C616 a_26096_6996# gnd 2.45fF
C617 a_15204_6671# gnd 2.23fF
C618 a_13855_6488# gnd 2.38fF
C619 a_17969_6950# gnd 2.18fF
C620 a_15940_6466# gnd 2.52fF
C621 a_8876_6701# gnd 2.28fF
C622 a_5174_6209# gnd 2.49fF
C623 a_3820_6660# gnd 2.28fF
C624 a_118_6168# gnd 2.49fF
C625 a_10148_6630# gnd 2.23fF
C626 a_12913_6909# gnd 2.18fF
C627 a_10884_6425# gnd 2.52fF
C628 a_8880_6524# gnd 2.38fF
C629 a_5173_6666# gnd 2.23fF
C630 a_3824_6483# gnd 2.38fF
C631 a_25359_7106# gnd 2.28fF
C632 a_20303_6836# gnd 2.38fF
C633 a_21040_6955# gnd 2.45fF
C634 a_20303_7065# gnd 2.28fF
C635 a_28128_6749# gnd 2.52fF
C636 a_29063_7236# gnd 2.23fF
C637 a_23072_6708# gnd 2.52fF
C638 a_24007_7195# gnd 2.23fF
C639 a_15204_6901# gnd 2.38fF
C640 a_15941_7020# gnd 2.45fF
C641 a_7938_6945# gnd 2.18fF
C642 a_5909_6461# gnd 2.52fF
C643 a_117_6625# gnd 2.23fF
C644 a_2882_6904# gnd 2.18fF
C645 a_853_6420# gnd 2.52fF
C646 a_15204_7130# gnd 2.28fF
C647 a_10148_6860# gnd 2.38fF
C648 a_10885_6979# gnd 2.45fF
C649 a_10148_7089# gnd 2.28fF
C650 a_37076_7281# gnd 2.34fF
C651 a_37081_5200# gnd 3.32fF
C652 a_32020_7240# gnd 2.34fF
C653 a_32025_5159# gnd 3.32fF
C654 a_17973_6773# gnd 2.52fF
C655 a_18908_7260# gnd 2.23fF
C656 a_39098_7064# gnd 2.49fF
C657 a_38051_5121# gnd 3.68fF
C658 a_34042_7023# gnd 2.49fF
C659 a_38045_7510# gnd 2.45fF
C660 a_32995_5080# gnd 3.68fF
C661 a_32989_7469# gnd 2.45fF
C662 a_27045_7276# gnd 2.34fF
C663 a_27050_5195# gnd 3.32fF
C664 a_21989_7235# gnd 2.34fF
C665 a_21994_5154# gnd 3.32fF
C666 a_12917_6732# gnd 2.52fF
C667 a_13852_7219# gnd 2.23fF
C668 a_5173_6896# gnd 2.38fF
C669 a_5910_7015# gnd 2.45fF
C670 a_5173_7125# gnd 2.28fF
C671 a_117_6855# gnd 2.38fF
C672 a_854_6974# gnd 2.45fF
C673 a_117_7084# gnd 2.28fF
C674 a_29067_7059# gnd 2.49fF
C675 a_39093_7790# gnd 2.28fF
C676 a_35390_7298# gnd 2.49fF
C677 a_28020_5116# gnd 3.68fF
C678 a_24011_7018# gnd 2.49fF
C679 a_28014_7505# gnd 2.45fF
C680 a_22964_5075# gnd 3.68fF
C681 a_7942_6768# gnd 2.52fF
C682 a_8877_7255# gnd 2.23fF
C683 a_2886_6727# gnd 2.52fF
C684 a_3821_7214# gnd 2.23fF
C685 a_22958_7464# gnd 2.45fF
C686 a_16890_7300# gnd 2.34fF
C687 a_16895_5219# gnd 3.32fF
C688 a_11834_7259# gnd 2.34fF
C689 a_11839_5178# gnd 3.32fF
C690 a_34037_7749# gnd 2.28fF
C691 a_30334_7257# gnd 2.49fF
C692 a_39097_7613# gnd 2.38fF
C693 a_35390_7755# gnd 2.23fF
C694 a_34041_7572# gnd 2.38fF
C695 a_38155_8034# gnd 2.45fF
C696 a_36126_7550# gnd 2.52fF
C697 a_29062_7785# gnd 2.28fF
C698 a_25359_7293# gnd 2.49fF
C699 a_18912_7083# gnd 2.49fF
C700 a_24006_7744# gnd 2.28fF
C701 a_20303_7252# gnd 2.49fF
C702 a_17865_5140# gnd 3.68fF
C703 a_13856_7042# gnd 2.49fF
C704 a_17859_7529# gnd 2.45fF
C705 a_12809_5099# gnd 3.68fF
C706 a_12803_7488# gnd 2.45fF
C707 a_6859_7295# gnd 2.34fF
C708 a_6864_5214# gnd 3.32fF
C709 a_1803_7254# gnd 2.34fF
C710 a_1808_5173# gnd 3.32fF
C711 a_8881_7078# gnd 2.49fF
C712 a_30334_7714# gnd 2.23fF
C713 a_33099_7993# gnd 2.45fF
C714 a_31070_7509# gnd 2.52fF
C715 a_29066_7608# gnd 2.38fF
C716 a_25359_7750# gnd 2.23fF
C717 a_24010_7567# gnd 2.38fF
C718 a_35390_7985# gnd 2.38fF
C719 a_36127_8104# gnd 2.18fF
C720 a_28124_8029# gnd 2.45fF
C721 a_26095_7545# gnd 2.52fF
C722 a_20303_7709# gnd 2.23fF
C723 a_18907_7809# gnd 2.28fF
C724 a_15204_7317# gnd 2.49fF
C725 a_7834_5135# gnd 3.68fF
C726 a_3825_7037# gnd 2.49fF
C727 a_7828_7524# gnd 2.45fF
C728 a_2778_5094# gnd 3.68fF
C729 a_2772_7483# gnd 2.45fF
C730 a_13851_7768# gnd 2.28fF
C731 a_10148_7276# gnd 2.49fF
C732 a_23068_7988# gnd 2.45fF
C733 a_21039_7504# gnd 2.52fF
C734 a_18911_7632# gnd 2.38fF
C735 a_35390_8214# gnd 2.28fF
C736 a_30334_7944# gnd 2.38fF
C737 a_31071_8063# gnd 2.18fF
C738 a_30334_8173# gnd 2.28fF
C739 a_38159_7857# gnd 2.52fF
C740 a_39094_8344# gnd 2.23fF
C741 a_33103_7816# gnd 2.52fF
C742 a_34038_8303# gnd 2.23fF
C743 a_25359_7980# gnd 2.38fF
C744 a_26096_8099# gnd 2.18fF
C745 a_15204_7774# gnd 2.23fF
C746 a_13855_7591# gnd 2.38fF
C747 a_17969_8053# gnd 2.45fF
C748 a_15940_7569# gnd 2.52fF
C749 a_8876_7804# gnd 2.28fF
C750 a_5173_7312# gnd 2.49fF
C751 a_3820_7763# gnd 2.28fF
C752 a_117_7271# gnd 2.49fF
C753 a_10148_7733# gnd 2.23fF
C754 a_12913_8012# gnd 2.45fF
C755 a_10884_7528# gnd 2.52fF
C756 a_8880_7627# gnd 2.38fF
C757 a_5173_7769# gnd 2.23fF
C758 a_3824_7586# gnd 2.38fF
C759 a_25359_8209# gnd 2.28fF
C760 a_20303_7939# gnd 2.38fF
C761 a_21040_8058# gnd 2.18fF
C762 a_20303_8168# gnd 2.28fF
C763 a_39098_8167# gnd 2.49fF
C764 a_37081_7400# gnd 2.04fF
C765 a_28128_7852# gnd 2.52fF
C766 a_29063_8339# gnd 2.23fF
C767 a_23072_7811# gnd 2.52fF
C768 a_24007_8298# gnd 2.23fF
C769 a_34042_8126# gnd 2.49fF
C770 a_32025_7359# gnd 2.04fF
C771 a_38049_7333# gnd 2.28fF
C772 a_32993_7292# gnd 2.28fF
C773 a_29067_8162# gnd 2.49fF
C774 a_27050_7395# gnd 2.04fF
C775 a_15204_8004# gnd 2.38fF
C776 a_15941_8123# gnd 2.18fF
C777 a_7938_8048# gnd 2.45fF
C778 a_5909_7564# gnd 2.52fF
C779 a_117_7728# gnd 2.23fF
C780 a_2882_8007# gnd 2.45fF
C781 a_853_7523# gnd 2.52fF
C782 a_15204_8233# gnd 2.28fF
C783 a_10148_7963# gnd 2.38fF
C784 a_10885_8082# gnd 2.18fF
C785 a_10148_8192# gnd 2.28fF
C786 a_17973_7876# gnd 2.52fF
C787 a_18908_8363# gnd 2.23fF
C788 a_12917_7835# gnd 2.52fF
C789 a_13852_8322# gnd 2.23fF
C790 a_5173_7999# gnd 2.38fF
C791 a_5910_8118# gnd 2.18fF
C792 a_5173_8228# gnd 2.28fF
C793 a_117_7958# gnd 2.38fF
C794 a_854_8077# gnd 2.18fF
C795 a_117_8187# gnd 2.28fF
C796 a_24011_8121# gnd 2.49fF
C797 a_21994_7354# gnd 2.04fF
C798 a_39092_8893# gnd 2.28fF
C799 a_35390_8401# gnd 2.49fF
C800 a_28018_7328# gnd 2.28fF
C801 a_22962_7287# gnd 2.28fF
C802 a_34036_8852# gnd 2.28fF
C803 a_30334_8360# gnd 2.49fF
C804 a_39096_8716# gnd 2.38fF
C805 a_35389_8858# gnd 2.23fF
C806 a_34040_8675# gnd 2.38fF
C807 a_38154_9137# gnd 2.18fF
C808 a_36125_8653# gnd 2.52fF
C809 a_29061_8888# gnd 2.28fF
C810 a_25359_8396# gnd 2.49fF
C811 a_18912_8186# gnd 2.49fF
C812 a_16895_7419# gnd 2.04fF
C813 a_7942_7871# gnd 2.52fF
C814 a_8877_8358# gnd 2.23fF
C815 a_2886_7830# gnd 2.52fF
C816 a_3821_8317# gnd 2.23fF
C817 a_13856_8145# gnd 2.49fF
C818 a_11839_7378# gnd 2.04fF
C819 a_24005_8847# gnd 2.28fF
C820 a_20303_8355# gnd 2.49fF
C821 a_17863_7352# gnd 2.28fF
C822 a_12807_7311# gnd 2.28fF
C823 a_8881_8181# gnd 2.49fF
C824 a_6864_7414# gnd 2.04fF
C825 a_3825_8140# gnd 2.49fF
C826 a_1808_7373# gnd 2.04fF
C827 a_30333_8817# gnd 2.23fF
C828 a_33098_9096# gnd 2.18fF
C829 a_31069_8612# gnd 2.52fF
C830 a_29065_8711# gnd 2.38fF
C831 a_25358_8853# gnd 2.23fF
C832 a_24009_8670# gnd 2.38fF
C833 a_35389_9088# gnd 2.38fF
C834 a_36126_9207# gnd 2.38fF
C835 a_28123_9132# gnd 2.18fF
C836 a_26094_8648# gnd 2.52fF
C837 a_20302_8812# gnd 2.23fF
C838 a_18906_8912# gnd 2.28fF
C839 a_15204_8420# gnd 2.49fF
C840 a_7832_7347# gnd 2.28fF
C841 a_2776_7306# gnd 2.28fF
C842 a_13850_8871# gnd 2.28fF
C843 a_10148_8379# gnd 2.49fF
C844 a_23067_9091# gnd 2.18fF
C845 a_21038_8607# gnd 2.52fF
C846 a_18910_8735# gnd 2.38fF
C847 a_35389_9317# gnd 2.22fF
C848 a_30333_9047# gnd 2.38fF
C849 a_31070_9166# gnd 2.38fF
C850 a_30333_9276# gnd 2.22fF
C851 a_38158_8960# gnd 2.79fF
C852 a_39093_9447# gnd 2.75fF
C853 a_33102_8919# gnd 2.52fF
C854 a_34037_9406# gnd 2.23fF
C855 a_25358_9083# gnd 2.38fF
C856 a_26095_9202# gnd 2.38fF
C857 a_15203_8877# gnd 2.23fF
C858 a_13854_8694# gnd 2.38fF
C859 a_17968_9156# gnd 2.18fF
C860 a_15939_8672# gnd 2.52fF
C861 a_8875_8907# gnd 2.28fF
C862 a_5173_8415# gnd 2.49fF
C863 a_3819_8866# gnd 2.28fF
C864 a_117_8374# gnd 2.49fF
C865 a_10147_8836# gnd 2.23fF
C866 a_12912_9115# gnd 2.18fF
C867 a_10883_8631# gnd 2.52fF
C868 a_8879_8730# gnd 2.38fF
C869 a_5172_8872# gnd 2.23fF
C870 a_3823_8689# gnd 2.38fF
C871 a_25358_9312# gnd 2.22fF
C872 a_20302_9042# gnd 2.38fF
C873 a_21039_9161# gnd 2.38fF
C874 a_20302_9271# gnd 2.22fF
C875 a_34041_9229# gnd 2.98fF
C876 a_29066_9265# gnd 2.82fF
C877 a_28127_8955# gnd 2.52fF
C878 a_29062_9442# gnd 2.23fF
C879 a_23071_8914# gnd 2.52fF
C880 a_24006_9401# gnd 2.23fF
C881 a_15203_9107# gnd 2.38fF
C882 a_15940_9226# gnd 2.38fF
C883 a_7937_9151# gnd 2.18fF
C884 a_5908_8667# gnd 2.52fF
C885 a_116_8831# gnd 2.23fF
C886 a_2881_9110# gnd 2.18fF
C887 a_852_8626# gnd 2.52fF
C888 a_15203_9336# gnd 2.22fF
C889 a_10147_9066# gnd 2.38fF
C890 a_10884_9185# gnd 2.38fF
C891 a_10147_9295# gnd 2.22fF
C892 a_24010_9224# gnd 2.98fF
C893 a_18911_9289# gnd 2.97fF
C894 a_17972_8979# gnd 2.52fF
C895 a_18907_9466# gnd 2.23fF
C896 a_12916_8938# gnd 2.52fF
C897 a_13851_9425# gnd 2.23fF
C898 a_5172_9102# gnd 2.38fF
C899 a_5909_9221# gnd 2.38fF
C900 a_5172_9331# gnd 2.22fF
C901 a_116_9061# gnd 2.38fF
C902 a_853_9180# gnd 2.38fF
C903 a_13855_9248# gnd 2.98fF
C904 a_8880_9284# gnd 2.82fF
C905 a_7941_8974# gnd 2.52fF
C906 a_8876_9461# gnd 2.23fF
C907 a_2885_8933# gnd 2.52fF
C908 a_3820_9420# gnd 2.23fF
C909 a_3824_9243# gnd 2.98fF
C910 vdd gnd 950.06fF
