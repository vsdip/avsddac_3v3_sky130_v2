magic
tech sky130A
timestamp 1616169439
<< nwell >>
rect 278 8004 1089 8154
rect 4103 8028 4914 8178
rect 5559 7983 6370 8133
rect 9384 8007 10195 8157
rect 10939 8012 11750 8162
rect 14764 8036 15575 8186
rect 16220 7991 17031 8141
rect 20045 8015 20856 8165
rect 1290 7823 2101 7973
rect 3090 7794 3901 7944
rect 6571 7802 7382 7952
rect 8371 7773 9182 7923
rect 11951 7831 12762 7981
rect 13751 7802 14562 7952
rect 17232 7810 18043 7960
rect 19032 7781 19843 7931
rect 277 7589 1088 7739
rect 4102 7613 4913 7763
rect 5558 7568 6369 7718
rect 9383 7592 10194 7742
rect 10938 7597 11749 7747
rect 14763 7621 15574 7771
rect 16219 7576 17030 7726
rect 20044 7600 20855 7750
rect 1345 7262 2156 7412
rect 3040 7374 3851 7524
rect 6626 7241 7437 7391
rect 8321 7353 9132 7503
rect 12006 7270 12817 7420
rect 13701 7382 14512 7532
rect 17287 7249 18098 7399
rect 18982 7361 19793 7511
rect 283 7023 1094 7173
rect 4108 7047 4919 7197
rect 5564 7002 6375 7152
rect 9389 7026 10200 7176
rect 10944 7031 11755 7181
rect 14769 7055 15580 7205
rect 16225 7010 17036 7160
rect 20050 7034 20861 7184
rect 1295 6842 2106 6992
rect 3095 6813 3906 6963
rect 6576 6821 7387 6971
rect 8376 6792 9187 6942
rect 11956 6850 12767 7000
rect 13756 6821 14567 6971
rect 17237 6829 18048 6979
rect 19037 6800 19848 6950
rect 282 6608 1093 6758
rect 4107 6632 4918 6782
rect 5563 6587 6374 6737
rect 9388 6611 10199 6761
rect 10943 6616 11754 6766
rect 14768 6640 15579 6790
rect 16224 6595 17035 6745
rect 20049 6619 20860 6769
rect 1510 6330 2321 6480
rect 2887 6346 3698 6496
rect 6791 6309 7602 6459
rect 8168 6325 8979 6475
rect 12171 6338 12982 6488
rect 13548 6354 14359 6504
rect 17452 6317 18263 6467
rect 18829 6333 19640 6483
rect 290 6044 1101 6194
rect 4115 6068 4926 6218
rect 5571 6023 6382 6173
rect 9396 6047 10207 6197
rect 10951 6052 11762 6202
rect 14776 6076 15587 6226
rect 16232 6031 17043 6181
rect 20057 6055 20868 6205
rect 1302 5863 2113 6013
rect 3102 5834 3913 5984
rect 6583 5842 7394 5992
rect 8383 5813 9194 5963
rect 11963 5871 12774 6021
rect 13763 5842 14574 5992
rect 17244 5850 18055 6000
rect 19044 5821 19855 5971
rect 289 5629 1100 5779
rect 4114 5653 4925 5803
rect 5570 5608 6381 5758
rect 9395 5632 10206 5782
rect 10950 5637 11761 5787
rect 14775 5661 15586 5811
rect 16231 5616 17042 5766
rect 20056 5640 20867 5790
rect 1357 5302 2168 5452
rect 3052 5414 3863 5564
rect 6638 5281 7449 5431
rect 8333 5393 9144 5543
rect 12018 5310 12829 5460
rect 13713 5422 14524 5572
rect 17299 5289 18110 5439
rect 18994 5401 19805 5551
rect 295 5063 1106 5213
rect 4120 5087 4931 5237
rect 5576 5042 6387 5192
rect 9401 5066 10212 5216
rect 10956 5071 11767 5221
rect 14781 5095 15592 5245
rect 16237 5050 17048 5200
rect 20062 5074 20873 5224
rect 1307 4882 2118 5032
rect 3107 4853 3918 5003
rect 6588 4861 7399 5011
rect 8388 4832 9199 4982
rect 11968 4890 12779 5040
rect 13768 4861 14579 5011
rect 17249 4869 18060 5019
rect 19049 4840 19860 4990
rect 294 4648 1105 4798
rect 4119 4672 4930 4822
rect 5575 4627 6386 4777
rect 9400 4651 10211 4801
rect 10955 4656 11766 4806
rect 14780 4680 15591 4830
rect 16236 4635 17047 4785
rect 20061 4659 20872 4809
rect 1605 4338 2416 4488
rect 2812 4421 3623 4571
rect 6886 4317 7697 4467
rect 8093 4400 8904 4550
rect 12266 4346 13077 4496
rect 13473 4429 14284 4579
rect 17547 4325 18358 4475
rect 18754 4408 19565 4558
rect 298 4087 1109 4237
rect 4123 4111 4934 4261
rect 5579 4066 6390 4216
rect 9404 4090 10215 4240
rect 10959 4095 11770 4245
rect 14784 4119 15595 4269
rect 16240 4074 17051 4224
rect 20065 4098 20876 4248
rect 1310 3906 2121 4056
rect 3110 3877 3921 4027
rect 6591 3885 7402 4035
rect 8391 3856 9202 4006
rect 11971 3914 12782 4064
rect 13771 3885 14582 4035
rect 17252 3893 18063 4043
rect 19052 3864 19863 4014
rect 297 3672 1108 3822
rect 4122 3696 4933 3846
rect 5578 3651 6389 3801
rect 9403 3675 10214 3825
rect 10958 3680 11769 3830
rect 14783 3704 15594 3854
rect 16239 3659 17050 3809
rect 20064 3683 20875 3833
rect 1365 3345 2176 3495
rect 3060 3457 3871 3607
rect 6646 3324 7457 3474
rect 8341 3436 9152 3586
rect 12026 3353 12837 3503
rect 13721 3465 14532 3615
rect 17307 3332 18118 3482
rect 19002 3444 19813 3594
rect 303 3106 1114 3256
rect 4128 3130 4939 3280
rect 5584 3085 6395 3235
rect 9409 3109 10220 3259
rect 10964 3114 11775 3264
rect 14789 3138 15600 3288
rect 16245 3093 17056 3243
rect 20070 3117 20881 3267
rect 1315 2925 2126 3075
rect 3115 2896 3926 3046
rect 6596 2904 7407 3054
rect 8396 2875 9207 3025
rect 11976 2933 12787 3083
rect 13776 2904 14587 3054
rect 17257 2912 18068 3062
rect 19057 2883 19868 3033
rect 302 2691 1113 2841
rect 4127 2715 4938 2865
rect 5583 2670 6394 2820
rect 9408 2694 10219 2844
rect 10963 2699 11774 2849
rect 14788 2723 15599 2873
rect 16244 2678 17055 2828
rect 20069 2702 20880 2852
rect 1530 2413 2341 2563
rect 2907 2429 3718 2579
rect 6811 2392 7622 2542
rect 8188 2408 8999 2558
rect 12191 2421 13002 2571
rect 13568 2437 14379 2587
rect 17472 2400 18283 2550
rect 18849 2416 19660 2566
rect 310 2127 1121 2277
rect 4135 2151 4946 2301
rect 5591 2106 6402 2256
rect 9416 2130 10227 2280
rect 10971 2135 11782 2285
rect 14796 2159 15607 2309
rect 16252 2114 17063 2264
rect 20077 2138 20888 2288
rect 1322 1946 2133 2096
rect 3122 1917 3933 2067
rect 6603 1925 7414 2075
rect 8403 1896 9214 2046
rect 11983 1954 12794 2104
rect 13783 1925 14594 2075
rect 17264 1933 18075 2083
rect 19064 1904 19875 2054
rect 309 1712 1120 1862
rect 4134 1736 4945 1886
rect 5590 1691 6401 1841
rect 9415 1715 10226 1865
rect 10970 1720 11781 1870
rect 14795 1744 15606 1894
rect 16251 1699 17062 1849
rect 20076 1723 20887 1873
rect 1377 1385 2188 1535
rect 3072 1497 3883 1647
rect 6658 1364 7469 1514
rect 8353 1476 9164 1626
rect 12038 1393 12849 1543
rect 13733 1505 14544 1655
rect 17319 1372 18130 1522
rect 19014 1484 19825 1634
rect 315 1146 1126 1296
rect 4140 1170 4951 1320
rect 5596 1125 6407 1275
rect 9421 1149 10232 1299
rect 10976 1154 11787 1304
rect 14801 1178 15612 1328
rect 16257 1133 17068 1283
rect 20082 1157 20893 1307
rect 1327 965 2138 1115
rect 3127 936 3938 1086
rect 6608 944 7419 1094
rect 8408 915 9219 1065
rect 11988 973 12799 1123
rect 13788 944 14599 1094
rect 17269 952 18080 1102
rect 19069 923 19880 1073
rect 314 731 1125 881
rect 4139 755 4950 905
rect 5595 710 6406 860
rect 9420 734 10231 884
rect 10975 739 11786 889
rect 14800 763 15611 913
rect 16256 718 17067 868
rect 20081 742 20892 892
rect 1717 250 2528 400
rect 4807 162 5618 312
rect 6998 229 7809 379
rect 10068 155 10879 305
rect 12378 258 13189 408
rect 15468 170 16279 320
rect 17659 237 18470 387
<< nmos >>
rect 4171 8237 4221 8279
rect 4379 8237 4429 8279
rect 4587 8237 4637 8279
rect 4800 8237 4850 8279
rect 9452 8216 9502 8258
rect 9660 8216 9710 8258
rect 9868 8216 9918 8258
rect 10081 8216 10131 8258
rect 14832 8245 14882 8287
rect 15040 8245 15090 8287
rect 15248 8245 15298 8287
rect 15461 8245 15511 8287
rect 20113 8224 20163 8266
rect 20321 8224 20371 8266
rect 20529 8224 20579 8266
rect 20742 8224 20792 8266
rect 3158 8003 3208 8045
rect 3366 8003 3416 8045
rect 3574 8003 3624 8045
rect 3787 8003 3837 8045
rect 342 7903 392 7945
rect 555 7903 605 7945
rect 763 7903 813 7945
rect 971 7903 1021 7945
rect 8439 7982 8489 8024
rect 8647 7982 8697 8024
rect 8855 7982 8905 8024
rect 9068 7982 9118 8024
rect 5623 7882 5673 7924
rect 5836 7882 5886 7924
rect 6044 7882 6094 7924
rect 6252 7882 6302 7924
rect 4170 7822 4220 7864
rect 4378 7822 4428 7864
rect 4586 7822 4636 7864
rect 4799 7822 4849 7864
rect 1354 7722 1404 7764
rect 1567 7722 1617 7764
rect 1775 7722 1825 7764
rect 1983 7722 2033 7764
rect 13819 8011 13869 8053
rect 14027 8011 14077 8053
rect 14235 8011 14285 8053
rect 14448 8011 14498 8053
rect 11003 7911 11053 7953
rect 11216 7911 11266 7953
rect 11424 7911 11474 7953
rect 11632 7911 11682 7953
rect 9451 7801 9501 7843
rect 9659 7801 9709 7843
rect 9867 7801 9917 7843
rect 10080 7801 10130 7843
rect 6635 7701 6685 7743
rect 6848 7701 6898 7743
rect 7056 7701 7106 7743
rect 7264 7701 7314 7743
rect 19100 7990 19150 8032
rect 19308 7990 19358 8032
rect 19516 7990 19566 8032
rect 19729 7990 19779 8032
rect 16284 7890 16334 7932
rect 16497 7890 16547 7932
rect 16705 7890 16755 7932
rect 16913 7890 16963 7932
rect 14831 7830 14881 7872
rect 15039 7830 15089 7872
rect 15247 7830 15297 7872
rect 15460 7830 15510 7872
rect 3108 7583 3158 7625
rect 3316 7583 3366 7625
rect 3524 7583 3574 7625
rect 3737 7583 3787 7625
rect 341 7488 391 7530
rect 554 7488 604 7530
rect 762 7488 812 7530
rect 970 7488 1020 7530
rect 12015 7730 12065 7772
rect 12228 7730 12278 7772
rect 12436 7730 12486 7772
rect 12644 7730 12694 7772
rect 20112 7809 20162 7851
rect 20320 7809 20370 7851
rect 20528 7809 20578 7851
rect 20741 7809 20791 7851
rect 17296 7709 17346 7751
rect 17509 7709 17559 7751
rect 17717 7709 17767 7751
rect 17925 7709 17975 7751
rect 8389 7562 8439 7604
rect 8597 7562 8647 7604
rect 8805 7562 8855 7604
rect 9018 7562 9068 7604
rect 5622 7467 5672 7509
rect 5835 7467 5885 7509
rect 6043 7467 6093 7509
rect 6251 7467 6301 7509
rect 13769 7591 13819 7633
rect 13977 7591 14027 7633
rect 14185 7591 14235 7633
rect 14398 7591 14448 7633
rect 11002 7496 11052 7538
rect 11215 7496 11265 7538
rect 11423 7496 11473 7538
rect 11631 7496 11681 7538
rect 19050 7570 19100 7612
rect 19258 7570 19308 7612
rect 19466 7570 19516 7612
rect 19679 7570 19729 7612
rect 16283 7475 16333 7517
rect 16496 7475 16546 7517
rect 16704 7475 16754 7517
rect 16912 7475 16962 7517
rect 4176 7256 4226 7298
rect 4384 7256 4434 7298
rect 4592 7256 4642 7298
rect 4805 7256 4855 7298
rect 1409 7161 1459 7203
rect 1622 7161 1672 7203
rect 1830 7161 1880 7203
rect 2038 7161 2088 7203
rect 9457 7235 9507 7277
rect 9665 7235 9715 7277
rect 9873 7235 9923 7277
rect 10086 7235 10136 7277
rect 6690 7140 6740 7182
rect 6903 7140 6953 7182
rect 7111 7140 7161 7182
rect 7319 7140 7369 7182
rect 14837 7264 14887 7306
rect 15045 7264 15095 7306
rect 15253 7264 15303 7306
rect 15466 7264 15516 7306
rect 12070 7169 12120 7211
rect 12283 7169 12333 7211
rect 12491 7169 12541 7211
rect 12699 7169 12749 7211
rect 3163 7022 3213 7064
rect 3371 7022 3421 7064
rect 3579 7022 3629 7064
rect 3792 7022 3842 7064
rect 347 6922 397 6964
rect 560 6922 610 6964
rect 768 6922 818 6964
rect 976 6922 1026 6964
rect 8444 7001 8494 7043
rect 8652 7001 8702 7043
rect 8860 7001 8910 7043
rect 9073 7001 9123 7043
rect 20118 7243 20168 7285
rect 20326 7243 20376 7285
rect 20534 7243 20584 7285
rect 20747 7243 20797 7285
rect 17351 7148 17401 7190
rect 17564 7148 17614 7190
rect 17772 7148 17822 7190
rect 17980 7148 18030 7190
rect 5628 6901 5678 6943
rect 5841 6901 5891 6943
rect 6049 6901 6099 6943
rect 6257 6901 6307 6943
rect 4175 6841 4225 6883
rect 4383 6841 4433 6883
rect 4591 6841 4641 6883
rect 4804 6841 4854 6883
rect 1359 6741 1409 6783
rect 1572 6741 1622 6783
rect 1780 6741 1830 6783
rect 1988 6741 2038 6783
rect 13824 7030 13874 7072
rect 14032 7030 14082 7072
rect 14240 7030 14290 7072
rect 14453 7030 14503 7072
rect 11008 6930 11058 6972
rect 11221 6930 11271 6972
rect 11429 6930 11479 6972
rect 11637 6930 11687 6972
rect 9456 6820 9506 6862
rect 9664 6820 9714 6862
rect 9872 6820 9922 6862
rect 10085 6820 10135 6862
rect 6640 6720 6690 6762
rect 6853 6720 6903 6762
rect 7061 6720 7111 6762
rect 7269 6720 7319 6762
rect 19105 7009 19155 7051
rect 19313 7009 19363 7051
rect 19521 7009 19571 7051
rect 19734 7009 19784 7051
rect 16289 6909 16339 6951
rect 16502 6909 16552 6951
rect 16710 6909 16760 6951
rect 16918 6909 16968 6951
rect 14836 6849 14886 6891
rect 15044 6849 15094 6891
rect 15252 6849 15302 6891
rect 15465 6849 15515 6891
rect 2955 6555 3005 6597
rect 3163 6555 3213 6597
rect 3371 6555 3421 6597
rect 3584 6555 3634 6597
rect 12020 6749 12070 6791
rect 12233 6749 12283 6791
rect 12441 6749 12491 6791
rect 12649 6749 12699 6791
rect 20117 6828 20167 6870
rect 20325 6828 20375 6870
rect 20533 6828 20583 6870
rect 20746 6828 20796 6870
rect 17301 6728 17351 6770
rect 17514 6728 17564 6770
rect 17722 6728 17772 6770
rect 17930 6728 17980 6770
rect 346 6507 396 6549
rect 559 6507 609 6549
rect 767 6507 817 6549
rect 975 6507 1025 6549
rect 8236 6534 8286 6576
rect 8444 6534 8494 6576
rect 8652 6534 8702 6576
rect 8865 6534 8915 6576
rect 5627 6486 5677 6528
rect 5840 6486 5890 6528
rect 6048 6486 6098 6528
rect 6256 6486 6306 6528
rect 13616 6563 13666 6605
rect 13824 6563 13874 6605
rect 14032 6563 14082 6605
rect 14245 6563 14295 6605
rect 11007 6515 11057 6557
rect 11220 6515 11270 6557
rect 11428 6515 11478 6557
rect 11636 6515 11686 6557
rect 18897 6542 18947 6584
rect 19105 6542 19155 6584
rect 19313 6542 19363 6584
rect 19526 6542 19576 6584
rect 4183 6277 4233 6319
rect 4391 6277 4441 6319
rect 4599 6277 4649 6319
rect 4812 6277 4862 6319
rect 16288 6494 16338 6536
rect 16501 6494 16551 6536
rect 16709 6494 16759 6536
rect 16917 6494 16967 6536
rect 1574 6229 1624 6271
rect 1787 6229 1837 6271
rect 1995 6229 2045 6271
rect 2203 6229 2253 6271
rect 9464 6256 9514 6298
rect 9672 6256 9722 6298
rect 9880 6256 9930 6298
rect 10093 6256 10143 6298
rect 6855 6208 6905 6250
rect 7068 6208 7118 6250
rect 7276 6208 7326 6250
rect 7484 6208 7534 6250
rect 14844 6285 14894 6327
rect 15052 6285 15102 6327
rect 15260 6285 15310 6327
rect 15473 6285 15523 6327
rect 12235 6237 12285 6279
rect 12448 6237 12498 6279
rect 12656 6237 12706 6279
rect 12864 6237 12914 6279
rect 20125 6264 20175 6306
rect 20333 6264 20383 6306
rect 20541 6264 20591 6306
rect 20754 6264 20804 6306
rect 3170 6043 3220 6085
rect 3378 6043 3428 6085
rect 3586 6043 3636 6085
rect 3799 6043 3849 6085
rect 354 5943 404 5985
rect 567 5943 617 5985
rect 775 5943 825 5985
rect 983 5943 1033 5985
rect 8451 6022 8501 6064
rect 8659 6022 8709 6064
rect 8867 6022 8917 6064
rect 9080 6022 9130 6064
rect 17516 6216 17566 6258
rect 17729 6216 17779 6258
rect 17937 6216 17987 6258
rect 18145 6216 18195 6258
rect 5635 5922 5685 5964
rect 5848 5922 5898 5964
rect 6056 5922 6106 5964
rect 6264 5922 6314 5964
rect 4182 5862 4232 5904
rect 4390 5862 4440 5904
rect 4598 5862 4648 5904
rect 4811 5862 4861 5904
rect 1366 5762 1416 5804
rect 1579 5762 1629 5804
rect 1787 5762 1837 5804
rect 1995 5762 2045 5804
rect 13831 6051 13881 6093
rect 14039 6051 14089 6093
rect 14247 6051 14297 6093
rect 14460 6051 14510 6093
rect 11015 5951 11065 5993
rect 11228 5951 11278 5993
rect 11436 5951 11486 5993
rect 11644 5951 11694 5993
rect 9463 5841 9513 5883
rect 9671 5841 9721 5883
rect 9879 5841 9929 5883
rect 10092 5841 10142 5883
rect 6647 5741 6697 5783
rect 6860 5741 6910 5783
rect 7068 5741 7118 5783
rect 7276 5741 7326 5783
rect 19112 6030 19162 6072
rect 19320 6030 19370 6072
rect 19528 6030 19578 6072
rect 19741 6030 19791 6072
rect 16296 5930 16346 5972
rect 16509 5930 16559 5972
rect 16717 5930 16767 5972
rect 16925 5930 16975 5972
rect 14843 5870 14893 5912
rect 15051 5870 15101 5912
rect 15259 5870 15309 5912
rect 15472 5870 15522 5912
rect 3120 5623 3170 5665
rect 3328 5623 3378 5665
rect 3536 5623 3586 5665
rect 3749 5623 3799 5665
rect 353 5528 403 5570
rect 566 5528 616 5570
rect 774 5528 824 5570
rect 982 5528 1032 5570
rect 12027 5770 12077 5812
rect 12240 5770 12290 5812
rect 12448 5770 12498 5812
rect 12656 5770 12706 5812
rect 20124 5849 20174 5891
rect 20332 5849 20382 5891
rect 20540 5849 20590 5891
rect 20753 5849 20803 5891
rect 17308 5749 17358 5791
rect 17521 5749 17571 5791
rect 17729 5749 17779 5791
rect 17937 5749 17987 5791
rect 8401 5602 8451 5644
rect 8609 5602 8659 5644
rect 8817 5602 8867 5644
rect 9030 5602 9080 5644
rect 5634 5507 5684 5549
rect 5847 5507 5897 5549
rect 6055 5507 6105 5549
rect 6263 5507 6313 5549
rect 13781 5631 13831 5673
rect 13989 5631 14039 5673
rect 14197 5631 14247 5673
rect 14410 5631 14460 5673
rect 11014 5536 11064 5578
rect 11227 5536 11277 5578
rect 11435 5536 11485 5578
rect 11643 5536 11693 5578
rect 19062 5610 19112 5652
rect 19270 5610 19320 5652
rect 19478 5610 19528 5652
rect 19691 5610 19741 5652
rect 16295 5515 16345 5557
rect 16508 5515 16558 5557
rect 16716 5515 16766 5557
rect 16924 5515 16974 5557
rect 4188 5296 4238 5338
rect 4396 5296 4446 5338
rect 4604 5296 4654 5338
rect 4817 5296 4867 5338
rect 1421 5201 1471 5243
rect 1634 5201 1684 5243
rect 1842 5201 1892 5243
rect 2050 5201 2100 5243
rect 9469 5275 9519 5317
rect 9677 5275 9727 5317
rect 9885 5275 9935 5317
rect 10098 5275 10148 5317
rect 6702 5180 6752 5222
rect 6915 5180 6965 5222
rect 7123 5180 7173 5222
rect 7331 5180 7381 5222
rect 14849 5304 14899 5346
rect 15057 5304 15107 5346
rect 15265 5304 15315 5346
rect 15478 5304 15528 5346
rect 12082 5209 12132 5251
rect 12295 5209 12345 5251
rect 12503 5209 12553 5251
rect 12711 5209 12761 5251
rect 3175 5062 3225 5104
rect 3383 5062 3433 5104
rect 3591 5062 3641 5104
rect 3804 5062 3854 5104
rect 359 4962 409 5004
rect 572 4962 622 5004
rect 780 4962 830 5004
rect 988 4962 1038 5004
rect 8456 5041 8506 5083
rect 8664 5041 8714 5083
rect 8872 5041 8922 5083
rect 9085 5041 9135 5083
rect 20130 5283 20180 5325
rect 20338 5283 20388 5325
rect 20546 5283 20596 5325
rect 20759 5283 20809 5325
rect 17363 5188 17413 5230
rect 17576 5188 17626 5230
rect 17784 5188 17834 5230
rect 17992 5188 18042 5230
rect 5640 4941 5690 4983
rect 5853 4941 5903 4983
rect 6061 4941 6111 4983
rect 6269 4941 6319 4983
rect 4187 4881 4237 4923
rect 4395 4881 4445 4923
rect 4603 4881 4653 4923
rect 4816 4881 4866 4923
rect 1371 4781 1421 4823
rect 1584 4781 1634 4823
rect 1792 4781 1842 4823
rect 2000 4781 2050 4823
rect 13836 5070 13886 5112
rect 14044 5070 14094 5112
rect 14252 5070 14302 5112
rect 14465 5070 14515 5112
rect 11020 4970 11070 5012
rect 11233 4970 11283 5012
rect 11441 4970 11491 5012
rect 11649 4970 11699 5012
rect 9468 4860 9518 4902
rect 9676 4860 9726 4902
rect 9884 4860 9934 4902
rect 10097 4860 10147 4902
rect 6652 4760 6702 4802
rect 6865 4760 6915 4802
rect 7073 4760 7123 4802
rect 7281 4760 7331 4802
rect 19117 5049 19167 5091
rect 19325 5049 19375 5091
rect 19533 5049 19583 5091
rect 19746 5049 19796 5091
rect 16301 4949 16351 4991
rect 16514 4949 16564 4991
rect 16722 4949 16772 4991
rect 16930 4949 16980 4991
rect 14848 4889 14898 4931
rect 15056 4889 15106 4931
rect 15264 4889 15314 4931
rect 15477 4889 15527 4931
rect 2880 4630 2930 4672
rect 3088 4630 3138 4672
rect 3296 4630 3346 4672
rect 3509 4630 3559 4672
rect 12032 4789 12082 4831
rect 12245 4789 12295 4831
rect 12453 4789 12503 4831
rect 12661 4789 12711 4831
rect 20129 4868 20179 4910
rect 20337 4868 20387 4910
rect 20545 4868 20595 4910
rect 20758 4868 20808 4910
rect 17313 4768 17363 4810
rect 17526 4768 17576 4810
rect 17734 4768 17784 4810
rect 17942 4768 17992 4810
rect 358 4547 408 4589
rect 571 4547 621 4589
rect 779 4547 829 4589
rect 987 4547 1037 4589
rect 8161 4609 8211 4651
rect 8369 4609 8419 4651
rect 8577 4609 8627 4651
rect 8790 4609 8840 4651
rect 5639 4526 5689 4568
rect 5852 4526 5902 4568
rect 6060 4526 6110 4568
rect 6268 4526 6318 4568
rect 13541 4638 13591 4680
rect 13749 4638 13799 4680
rect 13957 4638 14007 4680
rect 14170 4638 14220 4680
rect 4191 4320 4241 4362
rect 4399 4320 4449 4362
rect 4607 4320 4657 4362
rect 4820 4320 4870 4362
rect 1669 4237 1719 4279
rect 1882 4237 1932 4279
rect 2090 4237 2140 4279
rect 2298 4237 2348 4279
rect 11019 4555 11069 4597
rect 11232 4555 11282 4597
rect 11440 4555 11490 4597
rect 11648 4555 11698 4597
rect 9472 4299 9522 4341
rect 9680 4299 9730 4341
rect 9888 4299 9938 4341
rect 10101 4299 10151 4341
rect 18822 4617 18872 4659
rect 19030 4617 19080 4659
rect 19238 4617 19288 4659
rect 19451 4617 19501 4659
rect 16300 4534 16350 4576
rect 16513 4534 16563 4576
rect 16721 4534 16771 4576
rect 16929 4534 16979 4576
rect 6950 4216 7000 4258
rect 7163 4216 7213 4258
rect 7371 4216 7421 4258
rect 7579 4216 7629 4258
rect 14852 4328 14902 4370
rect 15060 4328 15110 4370
rect 15268 4328 15318 4370
rect 15481 4328 15531 4370
rect 12330 4245 12380 4287
rect 12543 4245 12593 4287
rect 12751 4245 12801 4287
rect 12959 4245 13009 4287
rect 20133 4307 20183 4349
rect 20341 4307 20391 4349
rect 20549 4307 20599 4349
rect 20762 4307 20812 4349
rect 3178 4086 3228 4128
rect 3386 4086 3436 4128
rect 3594 4086 3644 4128
rect 3807 4086 3857 4128
rect 362 3986 412 4028
rect 575 3986 625 4028
rect 783 3986 833 4028
rect 991 3986 1041 4028
rect 8459 4065 8509 4107
rect 8667 4065 8717 4107
rect 8875 4065 8925 4107
rect 9088 4065 9138 4107
rect 17611 4224 17661 4266
rect 17824 4224 17874 4266
rect 18032 4224 18082 4266
rect 18240 4224 18290 4266
rect 5643 3965 5693 4007
rect 5856 3965 5906 4007
rect 6064 3965 6114 4007
rect 6272 3965 6322 4007
rect 4190 3905 4240 3947
rect 4398 3905 4448 3947
rect 4606 3905 4656 3947
rect 4819 3905 4869 3947
rect 1374 3805 1424 3847
rect 1587 3805 1637 3847
rect 1795 3805 1845 3847
rect 2003 3805 2053 3847
rect 13839 4094 13889 4136
rect 14047 4094 14097 4136
rect 14255 4094 14305 4136
rect 14468 4094 14518 4136
rect 11023 3994 11073 4036
rect 11236 3994 11286 4036
rect 11444 3994 11494 4036
rect 11652 3994 11702 4036
rect 9471 3884 9521 3926
rect 9679 3884 9729 3926
rect 9887 3884 9937 3926
rect 10100 3884 10150 3926
rect 6655 3784 6705 3826
rect 6868 3784 6918 3826
rect 7076 3784 7126 3826
rect 7284 3784 7334 3826
rect 19120 4073 19170 4115
rect 19328 4073 19378 4115
rect 19536 4073 19586 4115
rect 19749 4073 19799 4115
rect 16304 3973 16354 4015
rect 16517 3973 16567 4015
rect 16725 3973 16775 4015
rect 16933 3973 16983 4015
rect 14851 3913 14901 3955
rect 15059 3913 15109 3955
rect 15267 3913 15317 3955
rect 15480 3913 15530 3955
rect 3128 3666 3178 3708
rect 3336 3666 3386 3708
rect 3544 3666 3594 3708
rect 3757 3666 3807 3708
rect 361 3571 411 3613
rect 574 3571 624 3613
rect 782 3571 832 3613
rect 990 3571 1040 3613
rect 12035 3813 12085 3855
rect 12248 3813 12298 3855
rect 12456 3813 12506 3855
rect 12664 3813 12714 3855
rect 20132 3892 20182 3934
rect 20340 3892 20390 3934
rect 20548 3892 20598 3934
rect 20761 3892 20811 3934
rect 17316 3792 17366 3834
rect 17529 3792 17579 3834
rect 17737 3792 17787 3834
rect 17945 3792 17995 3834
rect 8409 3645 8459 3687
rect 8617 3645 8667 3687
rect 8825 3645 8875 3687
rect 9038 3645 9088 3687
rect 5642 3550 5692 3592
rect 5855 3550 5905 3592
rect 6063 3550 6113 3592
rect 6271 3550 6321 3592
rect 13789 3674 13839 3716
rect 13997 3674 14047 3716
rect 14205 3674 14255 3716
rect 14418 3674 14468 3716
rect 11022 3579 11072 3621
rect 11235 3579 11285 3621
rect 11443 3579 11493 3621
rect 11651 3579 11701 3621
rect 19070 3653 19120 3695
rect 19278 3653 19328 3695
rect 19486 3653 19536 3695
rect 19699 3653 19749 3695
rect 16303 3558 16353 3600
rect 16516 3558 16566 3600
rect 16724 3558 16774 3600
rect 16932 3558 16982 3600
rect 4196 3339 4246 3381
rect 4404 3339 4454 3381
rect 4612 3339 4662 3381
rect 4825 3339 4875 3381
rect 1429 3244 1479 3286
rect 1642 3244 1692 3286
rect 1850 3244 1900 3286
rect 2058 3244 2108 3286
rect 9477 3318 9527 3360
rect 9685 3318 9735 3360
rect 9893 3318 9943 3360
rect 10106 3318 10156 3360
rect 6710 3223 6760 3265
rect 6923 3223 6973 3265
rect 7131 3223 7181 3265
rect 7339 3223 7389 3265
rect 14857 3347 14907 3389
rect 15065 3347 15115 3389
rect 15273 3347 15323 3389
rect 15486 3347 15536 3389
rect 12090 3252 12140 3294
rect 12303 3252 12353 3294
rect 12511 3252 12561 3294
rect 12719 3252 12769 3294
rect 3183 3105 3233 3147
rect 3391 3105 3441 3147
rect 3599 3105 3649 3147
rect 3812 3105 3862 3147
rect 367 3005 417 3047
rect 580 3005 630 3047
rect 788 3005 838 3047
rect 996 3005 1046 3047
rect 8464 3084 8514 3126
rect 8672 3084 8722 3126
rect 8880 3084 8930 3126
rect 9093 3084 9143 3126
rect 20138 3326 20188 3368
rect 20346 3326 20396 3368
rect 20554 3326 20604 3368
rect 20767 3326 20817 3368
rect 17371 3231 17421 3273
rect 17584 3231 17634 3273
rect 17792 3231 17842 3273
rect 18000 3231 18050 3273
rect 5648 2984 5698 3026
rect 5861 2984 5911 3026
rect 6069 2984 6119 3026
rect 6277 2984 6327 3026
rect 4195 2924 4245 2966
rect 4403 2924 4453 2966
rect 4611 2924 4661 2966
rect 4824 2924 4874 2966
rect 1379 2824 1429 2866
rect 1592 2824 1642 2866
rect 1800 2824 1850 2866
rect 2008 2824 2058 2866
rect 13844 3113 13894 3155
rect 14052 3113 14102 3155
rect 14260 3113 14310 3155
rect 14473 3113 14523 3155
rect 11028 3013 11078 3055
rect 11241 3013 11291 3055
rect 11449 3013 11499 3055
rect 11657 3013 11707 3055
rect 9476 2903 9526 2945
rect 9684 2903 9734 2945
rect 9892 2903 9942 2945
rect 10105 2903 10155 2945
rect 6660 2803 6710 2845
rect 6873 2803 6923 2845
rect 7081 2803 7131 2845
rect 7289 2803 7339 2845
rect 19125 3092 19175 3134
rect 19333 3092 19383 3134
rect 19541 3092 19591 3134
rect 19754 3092 19804 3134
rect 16309 2992 16359 3034
rect 16522 2992 16572 3034
rect 16730 2992 16780 3034
rect 16938 2992 16988 3034
rect 14856 2932 14906 2974
rect 15064 2932 15114 2974
rect 15272 2932 15322 2974
rect 15485 2932 15535 2974
rect 2975 2638 3025 2680
rect 3183 2638 3233 2680
rect 3391 2638 3441 2680
rect 3604 2638 3654 2680
rect 12040 2832 12090 2874
rect 12253 2832 12303 2874
rect 12461 2832 12511 2874
rect 12669 2832 12719 2874
rect 20137 2911 20187 2953
rect 20345 2911 20395 2953
rect 20553 2911 20603 2953
rect 20766 2911 20816 2953
rect 17321 2811 17371 2853
rect 17534 2811 17584 2853
rect 17742 2811 17792 2853
rect 17950 2811 18000 2853
rect 366 2590 416 2632
rect 579 2590 629 2632
rect 787 2590 837 2632
rect 995 2590 1045 2632
rect 8256 2617 8306 2659
rect 8464 2617 8514 2659
rect 8672 2617 8722 2659
rect 8885 2617 8935 2659
rect 5647 2569 5697 2611
rect 5860 2569 5910 2611
rect 6068 2569 6118 2611
rect 6276 2569 6326 2611
rect 13636 2646 13686 2688
rect 13844 2646 13894 2688
rect 14052 2646 14102 2688
rect 14265 2646 14315 2688
rect 11027 2598 11077 2640
rect 11240 2598 11290 2640
rect 11448 2598 11498 2640
rect 11656 2598 11706 2640
rect 18917 2625 18967 2667
rect 19125 2625 19175 2667
rect 19333 2625 19383 2667
rect 19546 2625 19596 2667
rect 4203 2360 4253 2402
rect 4411 2360 4461 2402
rect 4619 2360 4669 2402
rect 4832 2360 4882 2402
rect 16308 2577 16358 2619
rect 16521 2577 16571 2619
rect 16729 2577 16779 2619
rect 16937 2577 16987 2619
rect 1594 2312 1644 2354
rect 1807 2312 1857 2354
rect 2015 2312 2065 2354
rect 2223 2312 2273 2354
rect 9484 2339 9534 2381
rect 9692 2339 9742 2381
rect 9900 2339 9950 2381
rect 10113 2339 10163 2381
rect 6875 2291 6925 2333
rect 7088 2291 7138 2333
rect 7296 2291 7346 2333
rect 7504 2291 7554 2333
rect 14864 2368 14914 2410
rect 15072 2368 15122 2410
rect 15280 2368 15330 2410
rect 15493 2368 15543 2410
rect 12255 2320 12305 2362
rect 12468 2320 12518 2362
rect 12676 2320 12726 2362
rect 12884 2320 12934 2362
rect 20145 2347 20195 2389
rect 20353 2347 20403 2389
rect 20561 2347 20611 2389
rect 20774 2347 20824 2389
rect 3190 2126 3240 2168
rect 3398 2126 3448 2168
rect 3606 2126 3656 2168
rect 3819 2126 3869 2168
rect 374 2026 424 2068
rect 587 2026 637 2068
rect 795 2026 845 2068
rect 1003 2026 1053 2068
rect 8471 2105 8521 2147
rect 8679 2105 8729 2147
rect 8887 2105 8937 2147
rect 9100 2105 9150 2147
rect 17536 2299 17586 2341
rect 17749 2299 17799 2341
rect 17957 2299 18007 2341
rect 18165 2299 18215 2341
rect 5655 2005 5705 2047
rect 5868 2005 5918 2047
rect 6076 2005 6126 2047
rect 6284 2005 6334 2047
rect 4202 1945 4252 1987
rect 4410 1945 4460 1987
rect 4618 1945 4668 1987
rect 4831 1945 4881 1987
rect 1386 1845 1436 1887
rect 1599 1845 1649 1887
rect 1807 1845 1857 1887
rect 2015 1845 2065 1887
rect 13851 2134 13901 2176
rect 14059 2134 14109 2176
rect 14267 2134 14317 2176
rect 14480 2134 14530 2176
rect 11035 2034 11085 2076
rect 11248 2034 11298 2076
rect 11456 2034 11506 2076
rect 11664 2034 11714 2076
rect 9483 1924 9533 1966
rect 9691 1924 9741 1966
rect 9899 1924 9949 1966
rect 10112 1924 10162 1966
rect 6667 1824 6717 1866
rect 6880 1824 6930 1866
rect 7088 1824 7138 1866
rect 7296 1824 7346 1866
rect 19132 2113 19182 2155
rect 19340 2113 19390 2155
rect 19548 2113 19598 2155
rect 19761 2113 19811 2155
rect 16316 2013 16366 2055
rect 16529 2013 16579 2055
rect 16737 2013 16787 2055
rect 16945 2013 16995 2055
rect 14863 1953 14913 1995
rect 15071 1953 15121 1995
rect 15279 1953 15329 1995
rect 15492 1953 15542 1995
rect 3140 1706 3190 1748
rect 3348 1706 3398 1748
rect 3556 1706 3606 1748
rect 3769 1706 3819 1748
rect 373 1611 423 1653
rect 586 1611 636 1653
rect 794 1611 844 1653
rect 1002 1611 1052 1653
rect 12047 1853 12097 1895
rect 12260 1853 12310 1895
rect 12468 1853 12518 1895
rect 12676 1853 12726 1895
rect 20144 1932 20194 1974
rect 20352 1932 20402 1974
rect 20560 1932 20610 1974
rect 20773 1932 20823 1974
rect 17328 1832 17378 1874
rect 17541 1832 17591 1874
rect 17749 1832 17799 1874
rect 17957 1832 18007 1874
rect 8421 1685 8471 1727
rect 8629 1685 8679 1727
rect 8837 1685 8887 1727
rect 9050 1685 9100 1727
rect 5654 1590 5704 1632
rect 5867 1590 5917 1632
rect 6075 1590 6125 1632
rect 6283 1590 6333 1632
rect 13801 1714 13851 1756
rect 14009 1714 14059 1756
rect 14217 1714 14267 1756
rect 14430 1714 14480 1756
rect 11034 1619 11084 1661
rect 11247 1619 11297 1661
rect 11455 1619 11505 1661
rect 11663 1619 11713 1661
rect 19082 1693 19132 1735
rect 19290 1693 19340 1735
rect 19498 1693 19548 1735
rect 19711 1693 19761 1735
rect 16315 1598 16365 1640
rect 16528 1598 16578 1640
rect 16736 1598 16786 1640
rect 16944 1598 16994 1640
rect 4208 1379 4258 1421
rect 4416 1379 4466 1421
rect 4624 1379 4674 1421
rect 4837 1379 4887 1421
rect 1441 1284 1491 1326
rect 1654 1284 1704 1326
rect 1862 1284 1912 1326
rect 2070 1284 2120 1326
rect 9489 1358 9539 1400
rect 9697 1358 9747 1400
rect 9905 1358 9955 1400
rect 10118 1358 10168 1400
rect 6722 1263 6772 1305
rect 6935 1263 6985 1305
rect 7143 1263 7193 1305
rect 7351 1263 7401 1305
rect 14869 1387 14919 1429
rect 15077 1387 15127 1429
rect 15285 1387 15335 1429
rect 15498 1387 15548 1429
rect 12102 1292 12152 1334
rect 12315 1292 12365 1334
rect 12523 1292 12573 1334
rect 12731 1292 12781 1334
rect 3195 1145 3245 1187
rect 3403 1145 3453 1187
rect 3611 1145 3661 1187
rect 3824 1145 3874 1187
rect 379 1045 429 1087
rect 592 1045 642 1087
rect 800 1045 850 1087
rect 1008 1045 1058 1087
rect 8476 1124 8526 1166
rect 8684 1124 8734 1166
rect 8892 1124 8942 1166
rect 9105 1124 9155 1166
rect 20150 1366 20200 1408
rect 20358 1366 20408 1408
rect 20566 1366 20616 1408
rect 20779 1366 20829 1408
rect 17383 1271 17433 1313
rect 17596 1271 17646 1313
rect 17804 1271 17854 1313
rect 18012 1271 18062 1313
rect 5660 1024 5710 1066
rect 5873 1024 5923 1066
rect 6081 1024 6131 1066
rect 6289 1024 6339 1066
rect 4207 964 4257 1006
rect 4415 964 4465 1006
rect 4623 964 4673 1006
rect 4836 964 4886 1006
rect 1391 864 1441 906
rect 1604 864 1654 906
rect 1812 864 1862 906
rect 2020 864 2070 906
rect 13856 1153 13906 1195
rect 14064 1153 14114 1195
rect 14272 1153 14322 1195
rect 14485 1153 14535 1195
rect 11040 1053 11090 1095
rect 11253 1053 11303 1095
rect 11461 1053 11511 1095
rect 11669 1053 11719 1095
rect 9488 943 9538 985
rect 9696 943 9746 985
rect 9904 943 9954 985
rect 10117 943 10167 985
rect 6672 843 6722 885
rect 6885 843 6935 885
rect 7093 843 7143 885
rect 7301 843 7351 885
rect 19137 1132 19187 1174
rect 19345 1132 19395 1174
rect 19553 1132 19603 1174
rect 19766 1132 19816 1174
rect 16321 1032 16371 1074
rect 16534 1032 16584 1074
rect 16742 1032 16792 1074
rect 16950 1032 17000 1074
rect 14868 972 14918 1014
rect 15076 972 15126 1014
rect 15284 972 15334 1014
rect 15497 972 15547 1014
rect 12052 872 12102 914
rect 12265 872 12315 914
rect 12473 872 12523 914
rect 12681 872 12731 914
rect 20149 951 20199 993
rect 20357 951 20407 993
rect 20565 951 20615 993
rect 20778 951 20828 993
rect 17333 851 17383 893
rect 17546 851 17596 893
rect 17754 851 17804 893
rect 17962 851 18012 893
rect 378 630 428 672
rect 591 630 641 672
rect 799 630 849 672
rect 1007 630 1057 672
rect 5659 609 5709 651
rect 5872 609 5922 651
rect 6080 609 6130 651
rect 6288 609 6338 651
rect 11039 638 11089 680
rect 11252 638 11302 680
rect 11460 638 11510 680
rect 11668 638 11718 680
rect 16320 617 16370 659
rect 16533 617 16583 659
rect 16741 617 16791 659
rect 16949 617 16999 659
rect 1781 149 1831 191
rect 1994 149 2044 191
rect 2202 149 2252 191
rect 2410 149 2460 191
rect 7062 128 7112 170
rect 7275 128 7325 170
rect 7483 128 7533 170
rect 7691 128 7741 170
rect 4871 61 4921 103
rect 5084 61 5134 103
rect 5292 61 5342 103
rect 5500 61 5550 103
rect 12442 157 12492 199
rect 12655 157 12705 199
rect 12863 157 12913 199
rect 13071 157 13121 199
rect 17723 136 17773 178
rect 17936 136 17986 178
rect 18144 136 18194 178
rect 18352 136 18402 178
rect 10132 54 10182 96
rect 10345 54 10395 96
rect 10553 54 10603 96
rect 10761 54 10811 96
rect 15532 69 15582 111
rect 15745 69 15795 111
rect 15953 69 16003 111
rect 16161 69 16211 111
<< pmos >>
rect 342 8022 392 8122
rect 555 8022 605 8122
rect 763 8022 813 8122
rect 971 8022 1021 8122
rect 4171 8060 4221 8160
rect 4379 8060 4429 8160
rect 4587 8060 4637 8160
rect 4800 8060 4850 8160
rect 1354 7841 1404 7941
rect 1567 7841 1617 7941
rect 1775 7841 1825 7941
rect 1983 7841 2033 7941
rect 5623 8001 5673 8101
rect 5836 8001 5886 8101
rect 6044 8001 6094 8101
rect 6252 8001 6302 8101
rect 9452 8039 9502 8139
rect 9660 8039 9710 8139
rect 9868 8039 9918 8139
rect 10081 8039 10131 8139
rect 3158 7826 3208 7926
rect 3366 7826 3416 7926
rect 3574 7826 3624 7926
rect 3787 7826 3837 7926
rect 11003 8030 11053 8130
rect 11216 8030 11266 8130
rect 11424 8030 11474 8130
rect 11632 8030 11682 8130
rect 14832 8068 14882 8168
rect 15040 8068 15090 8168
rect 15248 8068 15298 8168
rect 15461 8068 15511 8168
rect 6635 7820 6685 7920
rect 6848 7820 6898 7920
rect 7056 7820 7106 7920
rect 7264 7820 7314 7920
rect 341 7607 391 7707
rect 554 7607 604 7707
rect 762 7607 812 7707
rect 970 7607 1020 7707
rect 4170 7645 4220 7745
rect 4378 7645 4428 7745
rect 4586 7645 4636 7745
rect 4799 7645 4849 7745
rect 8439 7805 8489 7905
rect 8647 7805 8697 7905
rect 8855 7805 8905 7905
rect 9068 7805 9118 7905
rect 12015 7849 12065 7949
rect 12228 7849 12278 7949
rect 12436 7849 12486 7949
rect 12644 7849 12694 7949
rect 16284 8009 16334 8109
rect 16497 8009 16547 8109
rect 16705 8009 16755 8109
rect 16913 8009 16963 8109
rect 20113 8047 20163 8147
rect 20321 8047 20371 8147
rect 20529 8047 20579 8147
rect 20742 8047 20792 8147
rect 13819 7834 13869 7934
rect 14027 7834 14077 7934
rect 14235 7834 14285 7934
rect 14448 7834 14498 7934
rect 5622 7586 5672 7686
rect 5835 7586 5885 7686
rect 6043 7586 6093 7686
rect 6251 7586 6301 7686
rect 9451 7624 9501 7724
rect 9659 7624 9709 7724
rect 9867 7624 9917 7724
rect 10080 7624 10130 7724
rect 17296 7828 17346 7928
rect 17509 7828 17559 7928
rect 17717 7828 17767 7928
rect 17925 7828 17975 7928
rect 11002 7615 11052 7715
rect 11215 7615 11265 7715
rect 11423 7615 11473 7715
rect 11631 7615 11681 7715
rect 14831 7653 14881 7753
rect 15039 7653 15089 7753
rect 15247 7653 15297 7753
rect 15460 7653 15510 7753
rect 19100 7813 19150 7913
rect 19308 7813 19358 7913
rect 19516 7813 19566 7913
rect 19729 7813 19779 7913
rect 3108 7406 3158 7506
rect 3316 7406 3366 7506
rect 3524 7406 3574 7506
rect 3737 7406 3787 7506
rect 8389 7385 8439 7485
rect 8597 7385 8647 7485
rect 8805 7385 8855 7485
rect 9018 7385 9068 7485
rect 16283 7594 16333 7694
rect 16496 7594 16546 7694
rect 16704 7594 16754 7694
rect 16912 7594 16962 7694
rect 20112 7632 20162 7732
rect 20320 7632 20370 7732
rect 20528 7632 20578 7732
rect 20741 7632 20791 7732
rect 13769 7414 13819 7514
rect 13977 7414 14027 7514
rect 14185 7414 14235 7514
rect 14398 7414 14448 7514
rect 19050 7393 19100 7493
rect 19258 7393 19308 7493
rect 19466 7393 19516 7493
rect 19679 7393 19729 7493
rect 1409 7280 1459 7380
rect 1622 7280 1672 7380
rect 1830 7280 1880 7380
rect 2038 7280 2088 7380
rect 6690 7259 6740 7359
rect 6903 7259 6953 7359
rect 7111 7259 7161 7359
rect 7319 7259 7369 7359
rect 347 7041 397 7141
rect 560 7041 610 7141
rect 768 7041 818 7141
rect 976 7041 1026 7141
rect 4176 7079 4226 7179
rect 4384 7079 4434 7179
rect 4592 7079 4642 7179
rect 4805 7079 4855 7179
rect 12070 7288 12120 7388
rect 12283 7288 12333 7388
rect 12491 7288 12541 7388
rect 12699 7288 12749 7388
rect 17351 7267 17401 7367
rect 17564 7267 17614 7367
rect 17772 7267 17822 7367
rect 17980 7267 18030 7367
rect 1359 6860 1409 6960
rect 1572 6860 1622 6960
rect 1780 6860 1830 6960
rect 1988 6860 2038 6960
rect 5628 7020 5678 7120
rect 5841 7020 5891 7120
rect 6049 7020 6099 7120
rect 6257 7020 6307 7120
rect 9457 7058 9507 7158
rect 9665 7058 9715 7158
rect 9873 7058 9923 7158
rect 10086 7058 10136 7158
rect 3163 6845 3213 6945
rect 3371 6845 3421 6945
rect 3579 6845 3629 6945
rect 3792 6845 3842 6945
rect 11008 7049 11058 7149
rect 11221 7049 11271 7149
rect 11429 7049 11479 7149
rect 11637 7049 11687 7149
rect 14837 7087 14887 7187
rect 15045 7087 15095 7187
rect 15253 7087 15303 7187
rect 15466 7087 15516 7187
rect 6640 6839 6690 6939
rect 6853 6839 6903 6939
rect 7061 6839 7111 6939
rect 7269 6839 7319 6939
rect 346 6626 396 6726
rect 559 6626 609 6726
rect 767 6626 817 6726
rect 975 6626 1025 6726
rect 4175 6664 4225 6764
rect 4383 6664 4433 6764
rect 4591 6664 4641 6764
rect 4804 6664 4854 6764
rect 8444 6824 8494 6924
rect 8652 6824 8702 6924
rect 8860 6824 8910 6924
rect 9073 6824 9123 6924
rect 12020 6868 12070 6968
rect 12233 6868 12283 6968
rect 12441 6868 12491 6968
rect 12649 6868 12699 6968
rect 16289 7028 16339 7128
rect 16502 7028 16552 7128
rect 16710 7028 16760 7128
rect 16918 7028 16968 7128
rect 20118 7066 20168 7166
rect 20326 7066 20376 7166
rect 20534 7066 20584 7166
rect 20747 7066 20797 7166
rect 13824 6853 13874 6953
rect 14032 6853 14082 6953
rect 14240 6853 14290 6953
rect 14453 6853 14503 6953
rect 5627 6605 5677 6705
rect 5840 6605 5890 6705
rect 6048 6605 6098 6705
rect 6256 6605 6306 6705
rect 9456 6643 9506 6743
rect 9664 6643 9714 6743
rect 9872 6643 9922 6743
rect 10085 6643 10135 6743
rect 17301 6847 17351 6947
rect 17514 6847 17564 6947
rect 17722 6847 17772 6947
rect 17930 6847 17980 6947
rect 11007 6634 11057 6734
rect 11220 6634 11270 6734
rect 11428 6634 11478 6734
rect 11636 6634 11686 6734
rect 14836 6672 14886 6772
rect 15044 6672 15094 6772
rect 15252 6672 15302 6772
rect 15465 6672 15515 6772
rect 19105 6832 19155 6932
rect 19313 6832 19363 6932
rect 19521 6832 19571 6932
rect 19734 6832 19784 6932
rect 1574 6348 1624 6448
rect 1787 6348 1837 6448
rect 1995 6348 2045 6448
rect 2203 6348 2253 6448
rect 2955 6378 3005 6478
rect 3163 6378 3213 6478
rect 3371 6378 3421 6478
rect 3584 6378 3634 6478
rect 16288 6613 16338 6713
rect 16501 6613 16551 6713
rect 16709 6613 16759 6713
rect 16917 6613 16967 6713
rect 20117 6651 20167 6751
rect 20325 6651 20375 6751
rect 20533 6651 20583 6751
rect 20746 6651 20796 6751
rect 6855 6327 6905 6427
rect 7068 6327 7118 6427
rect 7276 6327 7326 6427
rect 7484 6327 7534 6427
rect 8236 6357 8286 6457
rect 8444 6357 8494 6457
rect 8652 6357 8702 6457
rect 8865 6357 8915 6457
rect 12235 6356 12285 6456
rect 12448 6356 12498 6456
rect 12656 6356 12706 6456
rect 12864 6356 12914 6456
rect 13616 6386 13666 6486
rect 13824 6386 13874 6486
rect 14032 6386 14082 6486
rect 14245 6386 14295 6486
rect 354 6062 404 6162
rect 567 6062 617 6162
rect 775 6062 825 6162
rect 983 6062 1033 6162
rect 4183 6100 4233 6200
rect 4391 6100 4441 6200
rect 4599 6100 4649 6200
rect 4812 6100 4862 6200
rect 17516 6335 17566 6435
rect 17729 6335 17779 6435
rect 17937 6335 17987 6435
rect 18145 6335 18195 6435
rect 18897 6365 18947 6465
rect 19105 6365 19155 6465
rect 19313 6365 19363 6465
rect 19526 6365 19576 6465
rect 1366 5881 1416 5981
rect 1579 5881 1629 5981
rect 1787 5881 1837 5981
rect 1995 5881 2045 5981
rect 5635 6041 5685 6141
rect 5848 6041 5898 6141
rect 6056 6041 6106 6141
rect 6264 6041 6314 6141
rect 9464 6079 9514 6179
rect 9672 6079 9722 6179
rect 9880 6079 9930 6179
rect 10093 6079 10143 6179
rect 3170 5866 3220 5966
rect 3378 5866 3428 5966
rect 3586 5866 3636 5966
rect 3799 5866 3849 5966
rect 11015 6070 11065 6170
rect 11228 6070 11278 6170
rect 11436 6070 11486 6170
rect 11644 6070 11694 6170
rect 14844 6108 14894 6208
rect 15052 6108 15102 6208
rect 15260 6108 15310 6208
rect 15473 6108 15523 6208
rect 6647 5860 6697 5960
rect 6860 5860 6910 5960
rect 7068 5860 7118 5960
rect 7276 5860 7326 5960
rect 353 5647 403 5747
rect 566 5647 616 5747
rect 774 5647 824 5747
rect 982 5647 1032 5747
rect 4182 5685 4232 5785
rect 4390 5685 4440 5785
rect 4598 5685 4648 5785
rect 4811 5685 4861 5785
rect 8451 5845 8501 5945
rect 8659 5845 8709 5945
rect 8867 5845 8917 5945
rect 9080 5845 9130 5945
rect 12027 5889 12077 5989
rect 12240 5889 12290 5989
rect 12448 5889 12498 5989
rect 12656 5889 12706 5989
rect 16296 6049 16346 6149
rect 16509 6049 16559 6149
rect 16717 6049 16767 6149
rect 16925 6049 16975 6149
rect 20125 6087 20175 6187
rect 20333 6087 20383 6187
rect 20541 6087 20591 6187
rect 20754 6087 20804 6187
rect 13831 5874 13881 5974
rect 14039 5874 14089 5974
rect 14247 5874 14297 5974
rect 14460 5874 14510 5974
rect 5634 5626 5684 5726
rect 5847 5626 5897 5726
rect 6055 5626 6105 5726
rect 6263 5626 6313 5726
rect 9463 5664 9513 5764
rect 9671 5664 9721 5764
rect 9879 5664 9929 5764
rect 10092 5664 10142 5764
rect 17308 5868 17358 5968
rect 17521 5868 17571 5968
rect 17729 5868 17779 5968
rect 17937 5868 17987 5968
rect 11014 5655 11064 5755
rect 11227 5655 11277 5755
rect 11435 5655 11485 5755
rect 11643 5655 11693 5755
rect 14843 5693 14893 5793
rect 15051 5693 15101 5793
rect 15259 5693 15309 5793
rect 15472 5693 15522 5793
rect 19112 5853 19162 5953
rect 19320 5853 19370 5953
rect 19528 5853 19578 5953
rect 19741 5853 19791 5953
rect 3120 5446 3170 5546
rect 3328 5446 3378 5546
rect 3536 5446 3586 5546
rect 3749 5446 3799 5546
rect 8401 5425 8451 5525
rect 8609 5425 8659 5525
rect 8817 5425 8867 5525
rect 9030 5425 9080 5525
rect 16295 5634 16345 5734
rect 16508 5634 16558 5734
rect 16716 5634 16766 5734
rect 16924 5634 16974 5734
rect 20124 5672 20174 5772
rect 20332 5672 20382 5772
rect 20540 5672 20590 5772
rect 20753 5672 20803 5772
rect 13781 5454 13831 5554
rect 13989 5454 14039 5554
rect 14197 5454 14247 5554
rect 14410 5454 14460 5554
rect 19062 5433 19112 5533
rect 19270 5433 19320 5533
rect 19478 5433 19528 5533
rect 19691 5433 19741 5533
rect 1421 5320 1471 5420
rect 1634 5320 1684 5420
rect 1842 5320 1892 5420
rect 2050 5320 2100 5420
rect 6702 5299 6752 5399
rect 6915 5299 6965 5399
rect 7123 5299 7173 5399
rect 7331 5299 7381 5399
rect 359 5081 409 5181
rect 572 5081 622 5181
rect 780 5081 830 5181
rect 988 5081 1038 5181
rect 4188 5119 4238 5219
rect 4396 5119 4446 5219
rect 4604 5119 4654 5219
rect 4817 5119 4867 5219
rect 12082 5328 12132 5428
rect 12295 5328 12345 5428
rect 12503 5328 12553 5428
rect 12711 5328 12761 5428
rect 17363 5307 17413 5407
rect 17576 5307 17626 5407
rect 17784 5307 17834 5407
rect 17992 5307 18042 5407
rect 1371 4900 1421 5000
rect 1584 4900 1634 5000
rect 1792 4900 1842 5000
rect 2000 4900 2050 5000
rect 5640 5060 5690 5160
rect 5853 5060 5903 5160
rect 6061 5060 6111 5160
rect 6269 5060 6319 5160
rect 9469 5098 9519 5198
rect 9677 5098 9727 5198
rect 9885 5098 9935 5198
rect 10098 5098 10148 5198
rect 3175 4885 3225 4985
rect 3383 4885 3433 4985
rect 3591 4885 3641 4985
rect 3804 4885 3854 4985
rect 11020 5089 11070 5189
rect 11233 5089 11283 5189
rect 11441 5089 11491 5189
rect 11649 5089 11699 5189
rect 14849 5127 14899 5227
rect 15057 5127 15107 5227
rect 15265 5127 15315 5227
rect 15478 5127 15528 5227
rect 6652 4879 6702 4979
rect 6865 4879 6915 4979
rect 7073 4879 7123 4979
rect 7281 4879 7331 4979
rect 358 4666 408 4766
rect 571 4666 621 4766
rect 779 4666 829 4766
rect 987 4666 1037 4766
rect 4187 4704 4237 4804
rect 4395 4704 4445 4804
rect 4603 4704 4653 4804
rect 4816 4704 4866 4804
rect 8456 4864 8506 4964
rect 8664 4864 8714 4964
rect 8872 4864 8922 4964
rect 9085 4864 9135 4964
rect 12032 4908 12082 5008
rect 12245 4908 12295 5008
rect 12453 4908 12503 5008
rect 12661 4908 12711 5008
rect 16301 5068 16351 5168
rect 16514 5068 16564 5168
rect 16722 5068 16772 5168
rect 16930 5068 16980 5168
rect 20130 5106 20180 5206
rect 20338 5106 20388 5206
rect 20546 5106 20596 5206
rect 20759 5106 20809 5206
rect 13836 4893 13886 4993
rect 14044 4893 14094 4993
rect 14252 4893 14302 4993
rect 14465 4893 14515 4993
rect 5639 4645 5689 4745
rect 5852 4645 5902 4745
rect 6060 4645 6110 4745
rect 6268 4645 6318 4745
rect 9468 4683 9518 4783
rect 9676 4683 9726 4783
rect 9884 4683 9934 4783
rect 10097 4683 10147 4783
rect 17313 4887 17363 4987
rect 17526 4887 17576 4987
rect 17734 4887 17784 4987
rect 17942 4887 17992 4987
rect 11019 4674 11069 4774
rect 11232 4674 11282 4774
rect 11440 4674 11490 4774
rect 11648 4674 11698 4774
rect 14848 4712 14898 4812
rect 15056 4712 15106 4812
rect 15264 4712 15314 4812
rect 15477 4712 15527 4812
rect 19117 4872 19167 4972
rect 19325 4872 19375 4972
rect 19533 4872 19583 4972
rect 19746 4872 19796 4972
rect 1669 4356 1719 4456
rect 1882 4356 1932 4456
rect 2090 4356 2140 4456
rect 2298 4356 2348 4456
rect 2880 4453 2930 4553
rect 3088 4453 3138 4553
rect 3296 4453 3346 4553
rect 3509 4453 3559 4553
rect 16300 4653 16350 4753
rect 16513 4653 16563 4753
rect 16721 4653 16771 4753
rect 16929 4653 16979 4753
rect 20129 4691 20179 4791
rect 20337 4691 20387 4791
rect 20545 4691 20595 4791
rect 20758 4691 20808 4791
rect 6950 4335 7000 4435
rect 7163 4335 7213 4435
rect 7371 4335 7421 4435
rect 7579 4335 7629 4435
rect 8161 4432 8211 4532
rect 8369 4432 8419 4532
rect 8577 4432 8627 4532
rect 8790 4432 8840 4532
rect 12330 4364 12380 4464
rect 12543 4364 12593 4464
rect 12751 4364 12801 4464
rect 12959 4364 13009 4464
rect 13541 4461 13591 4561
rect 13749 4461 13799 4561
rect 13957 4461 14007 4561
rect 14170 4461 14220 4561
rect 362 4105 412 4205
rect 575 4105 625 4205
rect 783 4105 833 4205
rect 991 4105 1041 4205
rect 4191 4143 4241 4243
rect 4399 4143 4449 4243
rect 4607 4143 4657 4243
rect 4820 4143 4870 4243
rect 17611 4343 17661 4443
rect 17824 4343 17874 4443
rect 18032 4343 18082 4443
rect 18240 4343 18290 4443
rect 18822 4440 18872 4540
rect 19030 4440 19080 4540
rect 19238 4440 19288 4540
rect 19451 4440 19501 4540
rect 1374 3924 1424 4024
rect 1587 3924 1637 4024
rect 1795 3924 1845 4024
rect 2003 3924 2053 4024
rect 5643 4084 5693 4184
rect 5856 4084 5906 4184
rect 6064 4084 6114 4184
rect 6272 4084 6322 4184
rect 9472 4122 9522 4222
rect 9680 4122 9730 4222
rect 9888 4122 9938 4222
rect 10101 4122 10151 4222
rect 3178 3909 3228 4009
rect 3386 3909 3436 4009
rect 3594 3909 3644 4009
rect 3807 3909 3857 4009
rect 11023 4113 11073 4213
rect 11236 4113 11286 4213
rect 11444 4113 11494 4213
rect 11652 4113 11702 4213
rect 14852 4151 14902 4251
rect 15060 4151 15110 4251
rect 15268 4151 15318 4251
rect 15481 4151 15531 4251
rect 6655 3903 6705 4003
rect 6868 3903 6918 4003
rect 7076 3903 7126 4003
rect 7284 3903 7334 4003
rect 361 3690 411 3790
rect 574 3690 624 3790
rect 782 3690 832 3790
rect 990 3690 1040 3790
rect 4190 3728 4240 3828
rect 4398 3728 4448 3828
rect 4606 3728 4656 3828
rect 4819 3728 4869 3828
rect 8459 3888 8509 3988
rect 8667 3888 8717 3988
rect 8875 3888 8925 3988
rect 9088 3888 9138 3988
rect 12035 3932 12085 4032
rect 12248 3932 12298 4032
rect 12456 3932 12506 4032
rect 12664 3932 12714 4032
rect 16304 4092 16354 4192
rect 16517 4092 16567 4192
rect 16725 4092 16775 4192
rect 16933 4092 16983 4192
rect 20133 4130 20183 4230
rect 20341 4130 20391 4230
rect 20549 4130 20599 4230
rect 20762 4130 20812 4230
rect 13839 3917 13889 4017
rect 14047 3917 14097 4017
rect 14255 3917 14305 4017
rect 14468 3917 14518 4017
rect 5642 3669 5692 3769
rect 5855 3669 5905 3769
rect 6063 3669 6113 3769
rect 6271 3669 6321 3769
rect 9471 3707 9521 3807
rect 9679 3707 9729 3807
rect 9887 3707 9937 3807
rect 10100 3707 10150 3807
rect 17316 3911 17366 4011
rect 17529 3911 17579 4011
rect 17737 3911 17787 4011
rect 17945 3911 17995 4011
rect 11022 3698 11072 3798
rect 11235 3698 11285 3798
rect 11443 3698 11493 3798
rect 11651 3698 11701 3798
rect 14851 3736 14901 3836
rect 15059 3736 15109 3836
rect 15267 3736 15317 3836
rect 15480 3736 15530 3836
rect 19120 3896 19170 3996
rect 19328 3896 19378 3996
rect 19536 3896 19586 3996
rect 19749 3896 19799 3996
rect 3128 3489 3178 3589
rect 3336 3489 3386 3589
rect 3544 3489 3594 3589
rect 3757 3489 3807 3589
rect 8409 3468 8459 3568
rect 8617 3468 8667 3568
rect 8825 3468 8875 3568
rect 9038 3468 9088 3568
rect 16303 3677 16353 3777
rect 16516 3677 16566 3777
rect 16724 3677 16774 3777
rect 16932 3677 16982 3777
rect 20132 3715 20182 3815
rect 20340 3715 20390 3815
rect 20548 3715 20598 3815
rect 20761 3715 20811 3815
rect 13789 3497 13839 3597
rect 13997 3497 14047 3597
rect 14205 3497 14255 3597
rect 14418 3497 14468 3597
rect 19070 3476 19120 3576
rect 19278 3476 19328 3576
rect 19486 3476 19536 3576
rect 19699 3476 19749 3576
rect 1429 3363 1479 3463
rect 1642 3363 1692 3463
rect 1850 3363 1900 3463
rect 2058 3363 2108 3463
rect 6710 3342 6760 3442
rect 6923 3342 6973 3442
rect 7131 3342 7181 3442
rect 7339 3342 7389 3442
rect 367 3124 417 3224
rect 580 3124 630 3224
rect 788 3124 838 3224
rect 996 3124 1046 3224
rect 4196 3162 4246 3262
rect 4404 3162 4454 3262
rect 4612 3162 4662 3262
rect 4825 3162 4875 3262
rect 12090 3371 12140 3471
rect 12303 3371 12353 3471
rect 12511 3371 12561 3471
rect 12719 3371 12769 3471
rect 17371 3350 17421 3450
rect 17584 3350 17634 3450
rect 17792 3350 17842 3450
rect 18000 3350 18050 3450
rect 1379 2943 1429 3043
rect 1592 2943 1642 3043
rect 1800 2943 1850 3043
rect 2008 2943 2058 3043
rect 5648 3103 5698 3203
rect 5861 3103 5911 3203
rect 6069 3103 6119 3203
rect 6277 3103 6327 3203
rect 9477 3141 9527 3241
rect 9685 3141 9735 3241
rect 9893 3141 9943 3241
rect 10106 3141 10156 3241
rect 3183 2928 3233 3028
rect 3391 2928 3441 3028
rect 3599 2928 3649 3028
rect 3812 2928 3862 3028
rect 11028 3132 11078 3232
rect 11241 3132 11291 3232
rect 11449 3132 11499 3232
rect 11657 3132 11707 3232
rect 14857 3170 14907 3270
rect 15065 3170 15115 3270
rect 15273 3170 15323 3270
rect 15486 3170 15536 3270
rect 6660 2922 6710 3022
rect 6873 2922 6923 3022
rect 7081 2922 7131 3022
rect 7289 2922 7339 3022
rect 366 2709 416 2809
rect 579 2709 629 2809
rect 787 2709 837 2809
rect 995 2709 1045 2809
rect 4195 2747 4245 2847
rect 4403 2747 4453 2847
rect 4611 2747 4661 2847
rect 4824 2747 4874 2847
rect 8464 2907 8514 3007
rect 8672 2907 8722 3007
rect 8880 2907 8930 3007
rect 9093 2907 9143 3007
rect 12040 2951 12090 3051
rect 12253 2951 12303 3051
rect 12461 2951 12511 3051
rect 12669 2951 12719 3051
rect 16309 3111 16359 3211
rect 16522 3111 16572 3211
rect 16730 3111 16780 3211
rect 16938 3111 16988 3211
rect 20138 3149 20188 3249
rect 20346 3149 20396 3249
rect 20554 3149 20604 3249
rect 20767 3149 20817 3249
rect 13844 2936 13894 3036
rect 14052 2936 14102 3036
rect 14260 2936 14310 3036
rect 14473 2936 14523 3036
rect 5647 2688 5697 2788
rect 5860 2688 5910 2788
rect 6068 2688 6118 2788
rect 6276 2688 6326 2788
rect 9476 2726 9526 2826
rect 9684 2726 9734 2826
rect 9892 2726 9942 2826
rect 10105 2726 10155 2826
rect 17321 2930 17371 3030
rect 17534 2930 17584 3030
rect 17742 2930 17792 3030
rect 17950 2930 18000 3030
rect 11027 2717 11077 2817
rect 11240 2717 11290 2817
rect 11448 2717 11498 2817
rect 11656 2717 11706 2817
rect 14856 2755 14906 2855
rect 15064 2755 15114 2855
rect 15272 2755 15322 2855
rect 15485 2755 15535 2855
rect 19125 2915 19175 3015
rect 19333 2915 19383 3015
rect 19541 2915 19591 3015
rect 19754 2915 19804 3015
rect 1594 2431 1644 2531
rect 1807 2431 1857 2531
rect 2015 2431 2065 2531
rect 2223 2431 2273 2531
rect 2975 2461 3025 2561
rect 3183 2461 3233 2561
rect 3391 2461 3441 2561
rect 3604 2461 3654 2561
rect 16308 2696 16358 2796
rect 16521 2696 16571 2796
rect 16729 2696 16779 2796
rect 16937 2696 16987 2796
rect 20137 2734 20187 2834
rect 20345 2734 20395 2834
rect 20553 2734 20603 2834
rect 20766 2734 20816 2834
rect 6875 2410 6925 2510
rect 7088 2410 7138 2510
rect 7296 2410 7346 2510
rect 7504 2410 7554 2510
rect 8256 2440 8306 2540
rect 8464 2440 8514 2540
rect 8672 2440 8722 2540
rect 8885 2440 8935 2540
rect 12255 2439 12305 2539
rect 12468 2439 12518 2539
rect 12676 2439 12726 2539
rect 12884 2439 12934 2539
rect 13636 2469 13686 2569
rect 13844 2469 13894 2569
rect 14052 2469 14102 2569
rect 14265 2469 14315 2569
rect 374 2145 424 2245
rect 587 2145 637 2245
rect 795 2145 845 2245
rect 1003 2145 1053 2245
rect 4203 2183 4253 2283
rect 4411 2183 4461 2283
rect 4619 2183 4669 2283
rect 4832 2183 4882 2283
rect 17536 2418 17586 2518
rect 17749 2418 17799 2518
rect 17957 2418 18007 2518
rect 18165 2418 18215 2518
rect 18917 2448 18967 2548
rect 19125 2448 19175 2548
rect 19333 2448 19383 2548
rect 19546 2448 19596 2548
rect 1386 1964 1436 2064
rect 1599 1964 1649 2064
rect 1807 1964 1857 2064
rect 2015 1964 2065 2064
rect 5655 2124 5705 2224
rect 5868 2124 5918 2224
rect 6076 2124 6126 2224
rect 6284 2124 6334 2224
rect 9484 2162 9534 2262
rect 9692 2162 9742 2262
rect 9900 2162 9950 2262
rect 10113 2162 10163 2262
rect 3190 1949 3240 2049
rect 3398 1949 3448 2049
rect 3606 1949 3656 2049
rect 3819 1949 3869 2049
rect 11035 2153 11085 2253
rect 11248 2153 11298 2253
rect 11456 2153 11506 2253
rect 11664 2153 11714 2253
rect 14864 2191 14914 2291
rect 15072 2191 15122 2291
rect 15280 2191 15330 2291
rect 15493 2191 15543 2291
rect 6667 1943 6717 2043
rect 6880 1943 6930 2043
rect 7088 1943 7138 2043
rect 7296 1943 7346 2043
rect 373 1730 423 1830
rect 586 1730 636 1830
rect 794 1730 844 1830
rect 1002 1730 1052 1830
rect 4202 1768 4252 1868
rect 4410 1768 4460 1868
rect 4618 1768 4668 1868
rect 4831 1768 4881 1868
rect 8471 1928 8521 2028
rect 8679 1928 8729 2028
rect 8887 1928 8937 2028
rect 9100 1928 9150 2028
rect 12047 1972 12097 2072
rect 12260 1972 12310 2072
rect 12468 1972 12518 2072
rect 12676 1972 12726 2072
rect 16316 2132 16366 2232
rect 16529 2132 16579 2232
rect 16737 2132 16787 2232
rect 16945 2132 16995 2232
rect 20145 2170 20195 2270
rect 20353 2170 20403 2270
rect 20561 2170 20611 2270
rect 20774 2170 20824 2270
rect 13851 1957 13901 2057
rect 14059 1957 14109 2057
rect 14267 1957 14317 2057
rect 14480 1957 14530 2057
rect 5654 1709 5704 1809
rect 5867 1709 5917 1809
rect 6075 1709 6125 1809
rect 6283 1709 6333 1809
rect 9483 1747 9533 1847
rect 9691 1747 9741 1847
rect 9899 1747 9949 1847
rect 10112 1747 10162 1847
rect 17328 1951 17378 2051
rect 17541 1951 17591 2051
rect 17749 1951 17799 2051
rect 17957 1951 18007 2051
rect 11034 1738 11084 1838
rect 11247 1738 11297 1838
rect 11455 1738 11505 1838
rect 11663 1738 11713 1838
rect 14863 1776 14913 1876
rect 15071 1776 15121 1876
rect 15279 1776 15329 1876
rect 15492 1776 15542 1876
rect 19132 1936 19182 2036
rect 19340 1936 19390 2036
rect 19548 1936 19598 2036
rect 19761 1936 19811 2036
rect 3140 1529 3190 1629
rect 3348 1529 3398 1629
rect 3556 1529 3606 1629
rect 3769 1529 3819 1629
rect 8421 1508 8471 1608
rect 8629 1508 8679 1608
rect 8837 1508 8887 1608
rect 9050 1508 9100 1608
rect 16315 1717 16365 1817
rect 16528 1717 16578 1817
rect 16736 1717 16786 1817
rect 16944 1717 16994 1817
rect 20144 1755 20194 1855
rect 20352 1755 20402 1855
rect 20560 1755 20610 1855
rect 20773 1755 20823 1855
rect 13801 1537 13851 1637
rect 14009 1537 14059 1637
rect 14217 1537 14267 1637
rect 14430 1537 14480 1637
rect 19082 1516 19132 1616
rect 19290 1516 19340 1616
rect 19498 1516 19548 1616
rect 19711 1516 19761 1616
rect 1441 1403 1491 1503
rect 1654 1403 1704 1503
rect 1862 1403 1912 1503
rect 2070 1403 2120 1503
rect 6722 1382 6772 1482
rect 6935 1382 6985 1482
rect 7143 1382 7193 1482
rect 7351 1382 7401 1482
rect 379 1164 429 1264
rect 592 1164 642 1264
rect 800 1164 850 1264
rect 1008 1164 1058 1264
rect 4208 1202 4258 1302
rect 4416 1202 4466 1302
rect 4624 1202 4674 1302
rect 4837 1202 4887 1302
rect 12102 1411 12152 1511
rect 12315 1411 12365 1511
rect 12523 1411 12573 1511
rect 12731 1411 12781 1511
rect 17383 1390 17433 1490
rect 17596 1390 17646 1490
rect 17804 1390 17854 1490
rect 18012 1390 18062 1490
rect 1391 983 1441 1083
rect 1604 983 1654 1083
rect 1812 983 1862 1083
rect 2020 983 2070 1083
rect 5660 1143 5710 1243
rect 5873 1143 5923 1243
rect 6081 1143 6131 1243
rect 6289 1143 6339 1243
rect 9489 1181 9539 1281
rect 9697 1181 9747 1281
rect 9905 1181 9955 1281
rect 10118 1181 10168 1281
rect 3195 968 3245 1068
rect 3403 968 3453 1068
rect 3611 968 3661 1068
rect 3824 968 3874 1068
rect 11040 1172 11090 1272
rect 11253 1172 11303 1272
rect 11461 1172 11511 1272
rect 11669 1172 11719 1272
rect 14869 1210 14919 1310
rect 15077 1210 15127 1310
rect 15285 1210 15335 1310
rect 15498 1210 15548 1310
rect 6672 962 6722 1062
rect 6885 962 6935 1062
rect 7093 962 7143 1062
rect 7301 962 7351 1062
rect 378 749 428 849
rect 591 749 641 849
rect 799 749 849 849
rect 1007 749 1057 849
rect 4207 787 4257 887
rect 4415 787 4465 887
rect 4623 787 4673 887
rect 4836 787 4886 887
rect 8476 947 8526 1047
rect 8684 947 8734 1047
rect 8892 947 8942 1047
rect 9105 947 9155 1047
rect 12052 991 12102 1091
rect 12265 991 12315 1091
rect 12473 991 12523 1091
rect 12681 991 12731 1091
rect 16321 1151 16371 1251
rect 16534 1151 16584 1251
rect 16742 1151 16792 1251
rect 16950 1151 17000 1251
rect 20150 1189 20200 1289
rect 20358 1189 20408 1289
rect 20566 1189 20616 1289
rect 20779 1189 20829 1289
rect 13856 976 13906 1076
rect 14064 976 14114 1076
rect 14272 976 14322 1076
rect 14485 976 14535 1076
rect 5659 728 5709 828
rect 5872 728 5922 828
rect 6080 728 6130 828
rect 6288 728 6338 828
rect 9488 766 9538 866
rect 9696 766 9746 866
rect 9904 766 9954 866
rect 10117 766 10167 866
rect 17333 970 17383 1070
rect 17546 970 17596 1070
rect 17754 970 17804 1070
rect 17962 970 18012 1070
rect 11039 757 11089 857
rect 11252 757 11302 857
rect 11460 757 11510 857
rect 11668 757 11718 857
rect 14868 795 14918 895
rect 15076 795 15126 895
rect 15284 795 15334 895
rect 15497 795 15547 895
rect 19137 955 19187 1055
rect 19345 955 19395 1055
rect 19553 955 19603 1055
rect 19766 955 19816 1055
rect 16320 736 16370 836
rect 16533 736 16583 836
rect 16741 736 16791 836
rect 16949 736 16999 836
rect 20149 774 20199 874
rect 20357 774 20407 874
rect 20565 774 20615 874
rect 20778 774 20828 874
rect 1781 268 1831 368
rect 1994 268 2044 368
rect 2202 268 2252 368
rect 2410 268 2460 368
rect 4871 180 4921 280
rect 5084 180 5134 280
rect 5292 180 5342 280
rect 5500 180 5550 280
rect 7062 247 7112 347
rect 7275 247 7325 347
rect 7483 247 7533 347
rect 7691 247 7741 347
rect 12442 276 12492 376
rect 12655 276 12705 376
rect 12863 276 12913 376
rect 13071 276 13121 376
rect 10132 173 10182 273
rect 10345 173 10395 273
rect 10553 173 10603 273
rect 10761 173 10811 273
rect 15532 188 15582 288
rect 15745 188 15795 288
rect 15953 188 16003 288
rect 16161 188 16211 288
rect 17723 255 17773 355
rect 17936 255 17986 355
rect 18144 255 18194 355
rect 18352 255 18402 355
<< ndiff >>
rect 4122 8267 4171 8279
rect 4122 8247 4133 8267
rect 4153 8247 4171 8267
rect 4122 8237 4171 8247
rect 4221 8263 4265 8279
rect 4221 8243 4236 8263
rect 4256 8243 4265 8263
rect 4221 8237 4265 8243
rect 4335 8263 4379 8279
rect 4335 8243 4344 8263
rect 4364 8243 4379 8263
rect 4335 8237 4379 8243
rect 4429 8267 4478 8279
rect 4429 8247 4447 8267
rect 4467 8247 4478 8267
rect 4429 8237 4478 8247
rect 4543 8263 4587 8279
rect 4543 8243 4552 8263
rect 4572 8243 4587 8263
rect 4543 8237 4587 8243
rect 4637 8267 4686 8279
rect 4637 8247 4655 8267
rect 4675 8247 4686 8267
rect 4637 8237 4686 8247
rect 4756 8263 4800 8279
rect 4756 8243 4765 8263
rect 4785 8243 4800 8263
rect 4756 8237 4800 8243
rect 4850 8267 4899 8279
rect 4850 8247 4868 8267
rect 4888 8247 4899 8267
rect 4850 8237 4899 8247
rect 9403 8246 9452 8258
rect 9403 8226 9414 8246
rect 9434 8226 9452 8246
rect 9403 8216 9452 8226
rect 9502 8242 9546 8258
rect 9502 8222 9517 8242
rect 9537 8222 9546 8242
rect 9502 8216 9546 8222
rect 9616 8242 9660 8258
rect 9616 8222 9625 8242
rect 9645 8222 9660 8242
rect 9616 8216 9660 8222
rect 9710 8246 9759 8258
rect 9710 8226 9728 8246
rect 9748 8226 9759 8246
rect 9710 8216 9759 8226
rect 9824 8242 9868 8258
rect 9824 8222 9833 8242
rect 9853 8222 9868 8242
rect 9824 8216 9868 8222
rect 9918 8246 9967 8258
rect 9918 8226 9936 8246
rect 9956 8226 9967 8246
rect 9918 8216 9967 8226
rect 10037 8242 10081 8258
rect 10037 8222 10046 8242
rect 10066 8222 10081 8242
rect 10037 8216 10081 8222
rect 10131 8246 10180 8258
rect 10131 8226 10149 8246
rect 10169 8226 10180 8246
rect 10131 8216 10180 8226
rect 14783 8275 14832 8287
rect 14783 8255 14794 8275
rect 14814 8255 14832 8275
rect 14783 8245 14832 8255
rect 14882 8271 14926 8287
rect 14882 8251 14897 8271
rect 14917 8251 14926 8271
rect 14882 8245 14926 8251
rect 14996 8271 15040 8287
rect 14996 8251 15005 8271
rect 15025 8251 15040 8271
rect 14996 8245 15040 8251
rect 15090 8275 15139 8287
rect 15090 8255 15108 8275
rect 15128 8255 15139 8275
rect 15090 8245 15139 8255
rect 15204 8271 15248 8287
rect 15204 8251 15213 8271
rect 15233 8251 15248 8271
rect 15204 8245 15248 8251
rect 15298 8275 15347 8287
rect 15298 8255 15316 8275
rect 15336 8255 15347 8275
rect 15298 8245 15347 8255
rect 15417 8271 15461 8287
rect 15417 8251 15426 8271
rect 15446 8251 15461 8271
rect 15417 8245 15461 8251
rect 15511 8275 15560 8287
rect 15511 8255 15529 8275
rect 15549 8255 15560 8275
rect 15511 8245 15560 8255
rect 20064 8254 20113 8266
rect 20064 8234 20075 8254
rect 20095 8234 20113 8254
rect 20064 8224 20113 8234
rect 20163 8250 20207 8266
rect 20163 8230 20178 8250
rect 20198 8230 20207 8250
rect 20163 8224 20207 8230
rect 20277 8250 20321 8266
rect 20277 8230 20286 8250
rect 20306 8230 20321 8250
rect 20277 8224 20321 8230
rect 20371 8254 20420 8266
rect 20371 8234 20389 8254
rect 20409 8234 20420 8254
rect 20371 8224 20420 8234
rect 20485 8250 20529 8266
rect 20485 8230 20494 8250
rect 20514 8230 20529 8250
rect 20485 8224 20529 8230
rect 20579 8254 20628 8266
rect 20579 8234 20597 8254
rect 20617 8234 20628 8254
rect 20579 8224 20628 8234
rect 20698 8250 20742 8266
rect 20698 8230 20707 8250
rect 20727 8230 20742 8250
rect 20698 8224 20742 8230
rect 20792 8254 20841 8266
rect 20792 8234 20810 8254
rect 20830 8234 20841 8254
rect 20792 8224 20841 8234
rect 3109 8033 3158 8045
rect 3109 8013 3120 8033
rect 3140 8013 3158 8033
rect 3109 8003 3158 8013
rect 3208 8029 3252 8045
rect 3208 8009 3223 8029
rect 3243 8009 3252 8029
rect 3208 8003 3252 8009
rect 3322 8029 3366 8045
rect 3322 8009 3331 8029
rect 3351 8009 3366 8029
rect 3322 8003 3366 8009
rect 3416 8033 3465 8045
rect 3416 8013 3434 8033
rect 3454 8013 3465 8033
rect 3416 8003 3465 8013
rect 3530 8029 3574 8045
rect 3530 8009 3539 8029
rect 3559 8009 3574 8029
rect 3530 8003 3574 8009
rect 3624 8033 3673 8045
rect 3624 8013 3642 8033
rect 3662 8013 3673 8033
rect 3624 8003 3673 8013
rect 3743 8029 3787 8045
rect 3743 8009 3752 8029
rect 3772 8009 3787 8029
rect 3743 8003 3787 8009
rect 3837 8033 3886 8045
rect 3837 8013 3855 8033
rect 3875 8013 3886 8033
rect 3837 8003 3886 8013
rect 293 7935 342 7945
rect 293 7915 304 7935
rect 324 7915 342 7935
rect 293 7903 342 7915
rect 392 7939 436 7945
rect 392 7919 407 7939
rect 427 7919 436 7939
rect 392 7903 436 7919
rect 506 7935 555 7945
rect 506 7915 517 7935
rect 537 7915 555 7935
rect 506 7903 555 7915
rect 605 7939 649 7945
rect 605 7919 620 7939
rect 640 7919 649 7939
rect 605 7903 649 7919
rect 714 7935 763 7945
rect 714 7915 725 7935
rect 745 7915 763 7935
rect 714 7903 763 7915
rect 813 7939 857 7945
rect 813 7919 828 7939
rect 848 7919 857 7939
rect 813 7903 857 7919
rect 927 7939 971 7945
rect 927 7919 936 7939
rect 956 7919 971 7939
rect 927 7903 971 7919
rect 1021 7935 1070 7945
rect 1021 7915 1039 7935
rect 1059 7915 1070 7935
rect 1021 7903 1070 7915
rect 8390 8012 8439 8024
rect 8390 7992 8401 8012
rect 8421 7992 8439 8012
rect 8390 7982 8439 7992
rect 8489 8008 8533 8024
rect 8489 7988 8504 8008
rect 8524 7988 8533 8008
rect 8489 7982 8533 7988
rect 8603 8008 8647 8024
rect 8603 7988 8612 8008
rect 8632 7988 8647 8008
rect 8603 7982 8647 7988
rect 8697 8012 8746 8024
rect 8697 7992 8715 8012
rect 8735 7992 8746 8012
rect 8697 7982 8746 7992
rect 8811 8008 8855 8024
rect 8811 7988 8820 8008
rect 8840 7988 8855 8008
rect 8811 7982 8855 7988
rect 8905 8012 8954 8024
rect 8905 7992 8923 8012
rect 8943 7992 8954 8012
rect 8905 7982 8954 7992
rect 9024 8008 9068 8024
rect 9024 7988 9033 8008
rect 9053 7988 9068 8008
rect 9024 7982 9068 7988
rect 9118 8012 9167 8024
rect 9118 7992 9136 8012
rect 9156 7992 9167 8012
rect 13770 8041 13819 8053
rect 9118 7982 9167 7992
rect 5574 7914 5623 7924
rect 5574 7894 5585 7914
rect 5605 7894 5623 7914
rect 5574 7882 5623 7894
rect 5673 7918 5717 7924
rect 5673 7898 5688 7918
rect 5708 7898 5717 7918
rect 5673 7882 5717 7898
rect 5787 7914 5836 7924
rect 5787 7894 5798 7914
rect 5818 7894 5836 7914
rect 5787 7882 5836 7894
rect 5886 7918 5930 7924
rect 5886 7898 5901 7918
rect 5921 7898 5930 7918
rect 5886 7882 5930 7898
rect 5995 7914 6044 7924
rect 5995 7894 6006 7914
rect 6026 7894 6044 7914
rect 5995 7882 6044 7894
rect 6094 7918 6138 7924
rect 6094 7898 6109 7918
rect 6129 7898 6138 7918
rect 6094 7882 6138 7898
rect 6208 7918 6252 7924
rect 6208 7898 6217 7918
rect 6237 7898 6252 7918
rect 6208 7882 6252 7898
rect 6302 7914 6351 7924
rect 6302 7894 6320 7914
rect 6340 7894 6351 7914
rect 6302 7882 6351 7894
rect 4121 7852 4170 7864
rect 4121 7832 4132 7852
rect 4152 7832 4170 7852
rect 4121 7822 4170 7832
rect 4220 7848 4264 7864
rect 4220 7828 4235 7848
rect 4255 7828 4264 7848
rect 4220 7822 4264 7828
rect 4334 7848 4378 7864
rect 4334 7828 4343 7848
rect 4363 7828 4378 7848
rect 4334 7822 4378 7828
rect 4428 7852 4477 7864
rect 4428 7832 4446 7852
rect 4466 7832 4477 7852
rect 4428 7822 4477 7832
rect 4542 7848 4586 7864
rect 4542 7828 4551 7848
rect 4571 7828 4586 7848
rect 4542 7822 4586 7828
rect 4636 7852 4685 7864
rect 4636 7832 4654 7852
rect 4674 7832 4685 7852
rect 4636 7822 4685 7832
rect 4755 7848 4799 7864
rect 4755 7828 4764 7848
rect 4784 7828 4799 7848
rect 4755 7822 4799 7828
rect 4849 7852 4898 7864
rect 4849 7832 4867 7852
rect 4887 7832 4898 7852
rect 4849 7822 4898 7832
rect 1305 7754 1354 7764
rect 1305 7734 1316 7754
rect 1336 7734 1354 7754
rect 1305 7722 1354 7734
rect 1404 7758 1448 7764
rect 1404 7738 1419 7758
rect 1439 7738 1448 7758
rect 1404 7722 1448 7738
rect 1518 7754 1567 7764
rect 1518 7734 1529 7754
rect 1549 7734 1567 7754
rect 1518 7722 1567 7734
rect 1617 7758 1661 7764
rect 1617 7738 1632 7758
rect 1652 7738 1661 7758
rect 1617 7722 1661 7738
rect 1726 7754 1775 7764
rect 1726 7734 1737 7754
rect 1757 7734 1775 7754
rect 1726 7722 1775 7734
rect 1825 7758 1869 7764
rect 1825 7738 1840 7758
rect 1860 7738 1869 7758
rect 1825 7722 1869 7738
rect 1939 7758 1983 7764
rect 1939 7738 1948 7758
rect 1968 7738 1983 7758
rect 1939 7722 1983 7738
rect 2033 7754 2082 7764
rect 2033 7734 2051 7754
rect 2071 7734 2082 7754
rect 13770 8021 13781 8041
rect 13801 8021 13819 8041
rect 13770 8011 13819 8021
rect 13869 8037 13913 8053
rect 13869 8017 13884 8037
rect 13904 8017 13913 8037
rect 13869 8011 13913 8017
rect 13983 8037 14027 8053
rect 13983 8017 13992 8037
rect 14012 8017 14027 8037
rect 13983 8011 14027 8017
rect 14077 8041 14126 8053
rect 14077 8021 14095 8041
rect 14115 8021 14126 8041
rect 14077 8011 14126 8021
rect 14191 8037 14235 8053
rect 14191 8017 14200 8037
rect 14220 8017 14235 8037
rect 14191 8011 14235 8017
rect 14285 8041 14334 8053
rect 14285 8021 14303 8041
rect 14323 8021 14334 8041
rect 14285 8011 14334 8021
rect 14404 8037 14448 8053
rect 14404 8017 14413 8037
rect 14433 8017 14448 8037
rect 14404 8011 14448 8017
rect 14498 8041 14547 8053
rect 14498 8021 14516 8041
rect 14536 8021 14547 8041
rect 14498 8011 14547 8021
rect 10954 7943 11003 7953
rect 10954 7923 10965 7943
rect 10985 7923 11003 7943
rect 10954 7911 11003 7923
rect 11053 7947 11097 7953
rect 11053 7927 11068 7947
rect 11088 7927 11097 7947
rect 11053 7911 11097 7927
rect 11167 7943 11216 7953
rect 11167 7923 11178 7943
rect 11198 7923 11216 7943
rect 11167 7911 11216 7923
rect 11266 7947 11310 7953
rect 11266 7927 11281 7947
rect 11301 7927 11310 7947
rect 11266 7911 11310 7927
rect 11375 7943 11424 7953
rect 11375 7923 11386 7943
rect 11406 7923 11424 7943
rect 11375 7911 11424 7923
rect 11474 7947 11518 7953
rect 11474 7927 11489 7947
rect 11509 7927 11518 7947
rect 11474 7911 11518 7927
rect 11588 7947 11632 7953
rect 11588 7927 11597 7947
rect 11617 7927 11632 7947
rect 11588 7911 11632 7927
rect 11682 7943 11731 7953
rect 11682 7923 11700 7943
rect 11720 7923 11731 7943
rect 11682 7911 11731 7923
rect 2033 7722 2082 7734
rect 19051 8020 19100 8032
rect 9402 7831 9451 7843
rect 9402 7811 9413 7831
rect 9433 7811 9451 7831
rect 9402 7801 9451 7811
rect 9501 7827 9545 7843
rect 9501 7807 9516 7827
rect 9536 7807 9545 7827
rect 9501 7801 9545 7807
rect 9615 7827 9659 7843
rect 9615 7807 9624 7827
rect 9644 7807 9659 7827
rect 9615 7801 9659 7807
rect 9709 7831 9758 7843
rect 9709 7811 9727 7831
rect 9747 7811 9758 7831
rect 9709 7801 9758 7811
rect 9823 7827 9867 7843
rect 9823 7807 9832 7827
rect 9852 7807 9867 7827
rect 9823 7801 9867 7807
rect 9917 7831 9966 7843
rect 9917 7811 9935 7831
rect 9955 7811 9966 7831
rect 9917 7801 9966 7811
rect 10036 7827 10080 7843
rect 10036 7807 10045 7827
rect 10065 7807 10080 7827
rect 10036 7801 10080 7807
rect 10130 7831 10179 7843
rect 10130 7811 10148 7831
rect 10168 7811 10179 7831
rect 10130 7801 10179 7811
rect 6586 7733 6635 7743
rect 6586 7713 6597 7733
rect 6617 7713 6635 7733
rect 6586 7701 6635 7713
rect 6685 7737 6729 7743
rect 6685 7717 6700 7737
rect 6720 7717 6729 7737
rect 6685 7701 6729 7717
rect 6799 7733 6848 7743
rect 6799 7713 6810 7733
rect 6830 7713 6848 7733
rect 6799 7701 6848 7713
rect 6898 7737 6942 7743
rect 6898 7717 6913 7737
rect 6933 7717 6942 7737
rect 6898 7701 6942 7717
rect 7007 7733 7056 7743
rect 7007 7713 7018 7733
rect 7038 7713 7056 7733
rect 7007 7701 7056 7713
rect 7106 7737 7150 7743
rect 7106 7717 7121 7737
rect 7141 7717 7150 7737
rect 7106 7701 7150 7717
rect 7220 7737 7264 7743
rect 7220 7717 7229 7737
rect 7249 7717 7264 7737
rect 7220 7701 7264 7717
rect 7314 7733 7363 7743
rect 7314 7713 7332 7733
rect 7352 7713 7363 7733
rect 19051 8000 19062 8020
rect 19082 8000 19100 8020
rect 19051 7990 19100 8000
rect 19150 8016 19194 8032
rect 19150 7996 19165 8016
rect 19185 7996 19194 8016
rect 19150 7990 19194 7996
rect 19264 8016 19308 8032
rect 19264 7996 19273 8016
rect 19293 7996 19308 8016
rect 19264 7990 19308 7996
rect 19358 8020 19407 8032
rect 19358 8000 19376 8020
rect 19396 8000 19407 8020
rect 19358 7990 19407 8000
rect 19472 8016 19516 8032
rect 19472 7996 19481 8016
rect 19501 7996 19516 8016
rect 19472 7990 19516 7996
rect 19566 8020 19615 8032
rect 19566 8000 19584 8020
rect 19604 8000 19615 8020
rect 19566 7990 19615 8000
rect 19685 8016 19729 8032
rect 19685 7996 19694 8016
rect 19714 7996 19729 8016
rect 19685 7990 19729 7996
rect 19779 8020 19828 8032
rect 19779 8000 19797 8020
rect 19817 8000 19828 8020
rect 19779 7990 19828 8000
rect 16235 7922 16284 7932
rect 16235 7902 16246 7922
rect 16266 7902 16284 7922
rect 16235 7890 16284 7902
rect 16334 7926 16378 7932
rect 16334 7906 16349 7926
rect 16369 7906 16378 7926
rect 16334 7890 16378 7906
rect 16448 7922 16497 7932
rect 16448 7902 16459 7922
rect 16479 7902 16497 7922
rect 16448 7890 16497 7902
rect 16547 7926 16591 7932
rect 16547 7906 16562 7926
rect 16582 7906 16591 7926
rect 16547 7890 16591 7906
rect 16656 7922 16705 7932
rect 16656 7902 16667 7922
rect 16687 7902 16705 7922
rect 16656 7890 16705 7902
rect 16755 7926 16799 7932
rect 16755 7906 16770 7926
rect 16790 7906 16799 7926
rect 16755 7890 16799 7906
rect 16869 7926 16913 7932
rect 16869 7906 16878 7926
rect 16898 7906 16913 7926
rect 16869 7890 16913 7906
rect 16963 7922 17012 7932
rect 16963 7902 16981 7922
rect 17001 7902 17012 7922
rect 16963 7890 17012 7902
rect 14782 7860 14831 7872
rect 14782 7840 14793 7860
rect 14813 7840 14831 7860
rect 14782 7830 14831 7840
rect 14881 7856 14925 7872
rect 14881 7836 14896 7856
rect 14916 7836 14925 7856
rect 14881 7830 14925 7836
rect 14995 7856 15039 7872
rect 14995 7836 15004 7856
rect 15024 7836 15039 7856
rect 14995 7830 15039 7836
rect 15089 7860 15138 7872
rect 15089 7840 15107 7860
rect 15127 7840 15138 7860
rect 15089 7830 15138 7840
rect 15203 7856 15247 7872
rect 15203 7836 15212 7856
rect 15232 7836 15247 7856
rect 15203 7830 15247 7836
rect 15297 7860 15346 7872
rect 15297 7840 15315 7860
rect 15335 7840 15346 7860
rect 15297 7830 15346 7840
rect 15416 7856 15460 7872
rect 15416 7836 15425 7856
rect 15445 7836 15460 7856
rect 15416 7830 15460 7836
rect 15510 7860 15559 7872
rect 15510 7840 15528 7860
rect 15548 7840 15559 7860
rect 15510 7830 15559 7840
rect 11966 7762 12015 7772
rect 7314 7701 7363 7713
rect 3059 7613 3108 7625
rect 3059 7593 3070 7613
rect 3090 7593 3108 7613
rect 3059 7583 3108 7593
rect 3158 7609 3202 7625
rect 3158 7589 3173 7609
rect 3193 7589 3202 7609
rect 3158 7583 3202 7589
rect 3272 7609 3316 7625
rect 3272 7589 3281 7609
rect 3301 7589 3316 7609
rect 3272 7583 3316 7589
rect 3366 7613 3415 7625
rect 3366 7593 3384 7613
rect 3404 7593 3415 7613
rect 3366 7583 3415 7593
rect 3480 7609 3524 7625
rect 3480 7589 3489 7609
rect 3509 7589 3524 7609
rect 3480 7583 3524 7589
rect 3574 7613 3623 7625
rect 3574 7593 3592 7613
rect 3612 7593 3623 7613
rect 3574 7583 3623 7593
rect 3693 7609 3737 7625
rect 3693 7589 3702 7609
rect 3722 7589 3737 7609
rect 3693 7583 3737 7589
rect 3787 7613 3836 7625
rect 3787 7593 3805 7613
rect 3825 7593 3836 7613
rect 3787 7583 3836 7593
rect 292 7520 341 7530
rect 292 7500 303 7520
rect 323 7500 341 7520
rect 292 7488 341 7500
rect 391 7524 435 7530
rect 391 7504 406 7524
rect 426 7504 435 7524
rect 391 7488 435 7504
rect 505 7520 554 7530
rect 505 7500 516 7520
rect 536 7500 554 7520
rect 505 7488 554 7500
rect 604 7524 648 7530
rect 604 7504 619 7524
rect 639 7504 648 7524
rect 604 7488 648 7504
rect 713 7520 762 7530
rect 713 7500 724 7520
rect 744 7500 762 7520
rect 713 7488 762 7500
rect 812 7524 856 7530
rect 812 7504 827 7524
rect 847 7504 856 7524
rect 812 7488 856 7504
rect 926 7524 970 7530
rect 926 7504 935 7524
rect 955 7504 970 7524
rect 926 7488 970 7504
rect 1020 7520 1069 7530
rect 1020 7500 1038 7520
rect 1058 7500 1069 7520
rect 11966 7742 11977 7762
rect 11997 7742 12015 7762
rect 11966 7730 12015 7742
rect 12065 7766 12109 7772
rect 12065 7746 12080 7766
rect 12100 7746 12109 7766
rect 12065 7730 12109 7746
rect 12179 7762 12228 7772
rect 12179 7742 12190 7762
rect 12210 7742 12228 7762
rect 12179 7730 12228 7742
rect 12278 7766 12322 7772
rect 12278 7746 12293 7766
rect 12313 7746 12322 7766
rect 12278 7730 12322 7746
rect 12387 7762 12436 7772
rect 12387 7742 12398 7762
rect 12418 7742 12436 7762
rect 12387 7730 12436 7742
rect 12486 7766 12530 7772
rect 12486 7746 12501 7766
rect 12521 7746 12530 7766
rect 12486 7730 12530 7746
rect 12600 7766 12644 7772
rect 12600 7746 12609 7766
rect 12629 7746 12644 7766
rect 12600 7730 12644 7746
rect 12694 7762 12743 7772
rect 12694 7742 12712 7762
rect 12732 7742 12743 7762
rect 12694 7730 12743 7742
rect 20063 7839 20112 7851
rect 20063 7819 20074 7839
rect 20094 7819 20112 7839
rect 20063 7809 20112 7819
rect 20162 7835 20206 7851
rect 20162 7815 20177 7835
rect 20197 7815 20206 7835
rect 20162 7809 20206 7815
rect 20276 7835 20320 7851
rect 20276 7815 20285 7835
rect 20305 7815 20320 7835
rect 20276 7809 20320 7815
rect 20370 7839 20419 7851
rect 20370 7819 20388 7839
rect 20408 7819 20419 7839
rect 20370 7809 20419 7819
rect 20484 7835 20528 7851
rect 20484 7815 20493 7835
rect 20513 7815 20528 7835
rect 20484 7809 20528 7815
rect 20578 7839 20627 7851
rect 20578 7819 20596 7839
rect 20616 7819 20627 7839
rect 20578 7809 20627 7819
rect 20697 7835 20741 7851
rect 20697 7815 20706 7835
rect 20726 7815 20741 7835
rect 20697 7809 20741 7815
rect 20791 7839 20840 7851
rect 20791 7819 20809 7839
rect 20829 7819 20840 7839
rect 20791 7809 20840 7819
rect 17247 7741 17296 7751
rect 17247 7721 17258 7741
rect 17278 7721 17296 7741
rect 17247 7709 17296 7721
rect 17346 7745 17390 7751
rect 17346 7725 17361 7745
rect 17381 7725 17390 7745
rect 17346 7709 17390 7725
rect 17460 7741 17509 7751
rect 17460 7721 17471 7741
rect 17491 7721 17509 7741
rect 17460 7709 17509 7721
rect 17559 7745 17603 7751
rect 17559 7725 17574 7745
rect 17594 7725 17603 7745
rect 17559 7709 17603 7725
rect 17668 7741 17717 7751
rect 17668 7721 17679 7741
rect 17699 7721 17717 7741
rect 17668 7709 17717 7721
rect 17767 7745 17811 7751
rect 17767 7725 17782 7745
rect 17802 7725 17811 7745
rect 17767 7709 17811 7725
rect 17881 7745 17925 7751
rect 17881 7725 17890 7745
rect 17910 7725 17925 7745
rect 17881 7709 17925 7725
rect 17975 7741 18024 7751
rect 17975 7721 17993 7741
rect 18013 7721 18024 7741
rect 17975 7709 18024 7721
rect 13720 7621 13769 7633
rect 8340 7592 8389 7604
rect 1020 7488 1069 7500
rect 8340 7572 8351 7592
rect 8371 7572 8389 7592
rect 8340 7562 8389 7572
rect 8439 7588 8483 7604
rect 8439 7568 8454 7588
rect 8474 7568 8483 7588
rect 8439 7562 8483 7568
rect 8553 7588 8597 7604
rect 8553 7568 8562 7588
rect 8582 7568 8597 7588
rect 8553 7562 8597 7568
rect 8647 7592 8696 7604
rect 8647 7572 8665 7592
rect 8685 7572 8696 7592
rect 8647 7562 8696 7572
rect 8761 7588 8805 7604
rect 8761 7568 8770 7588
rect 8790 7568 8805 7588
rect 8761 7562 8805 7568
rect 8855 7592 8904 7604
rect 8855 7572 8873 7592
rect 8893 7572 8904 7592
rect 8855 7562 8904 7572
rect 8974 7588 9018 7604
rect 8974 7568 8983 7588
rect 9003 7568 9018 7588
rect 8974 7562 9018 7568
rect 9068 7592 9117 7604
rect 9068 7572 9086 7592
rect 9106 7572 9117 7592
rect 9068 7562 9117 7572
rect 5573 7499 5622 7509
rect 5573 7479 5584 7499
rect 5604 7479 5622 7499
rect 5573 7467 5622 7479
rect 5672 7503 5716 7509
rect 5672 7483 5687 7503
rect 5707 7483 5716 7503
rect 5672 7467 5716 7483
rect 5786 7499 5835 7509
rect 5786 7479 5797 7499
rect 5817 7479 5835 7499
rect 5786 7467 5835 7479
rect 5885 7503 5929 7509
rect 5885 7483 5900 7503
rect 5920 7483 5929 7503
rect 5885 7467 5929 7483
rect 5994 7499 6043 7509
rect 5994 7479 6005 7499
rect 6025 7479 6043 7499
rect 5994 7467 6043 7479
rect 6093 7503 6137 7509
rect 6093 7483 6108 7503
rect 6128 7483 6137 7503
rect 6093 7467 6137 7483
rect 6207 7503 6251 7509
rect 6207 7483 6216 7503
rect 6236 7483 6251 7503
rect 6207 7467 6251 7483
rect 6301 7499 6350 7509
rect 6301 7479 6319 7499
rect 6339 7479 6350 7499
rect 13720 7601 13731 7621
rect 13751 7601 13769 7621
rect 13720 7591 13769 7601
rect 13819 7617 13863 7633
rect 13819 7597 13834 7617
rect 13854 7597 13863 7617
rect 13819 7591 13863 7597
rect 13933 7617 13977 7633
rect 13933 7597 13942 7617
rect 13962 7597 13977 7617
rect 13933 7591 13977 7597
rect 14027 7621 14076 7633
rect 14027 7601 14045 7621
rect 14065 7601 14076 7621
rect 14027 7591 14076 7601
rect 14141 7617 14185 7633
rect 14141 7597 14150 7617
rect 14170 7597 14185 7617
rect 14141 7591 14185 7597
rect 14235 7621 14284 7633
rect 14235 7601 14253 7621
rect 14273 7601 14284 7621
rect 14235 7591 14284 7601
rect 14354 7617 14398 7633
rect 14354 7597 14363 7617
rect 14383 7597 14398 7617
rect 14354 7591 14398 7597
rect 14448 7621 14497 7633
rect 14448 7601 14466 7621
rect 14486 7601 14497 7621
rect 14448 7591 14497 7601
rect 6301 7467 6350 7479
rect 10953 7528 11002 7538
rect 10953 7508 10964 7528
rect 10984 7508 11002 7528
rect 10953 7496 11002 7508
rect 11052 7532 11096 7538
rect 11052 7512 11067 7532
rect 11087 7512 11096 7532
rect 11052 7496 11096 7512
rect 11166 7528 11215 7538
rect 11166 7508 11177 7528
rect 11197 7508 11215 7528
rect 11166 7496 11215 7508
rect 11265 7532 11309 7538
rect 11265 7512 11280 7532
rect 11300 7512 11309 7532
rect 11265 7496 11309 7512
rect 11374 7528 11423 7538
rect 11374 7508 11385 7528
rect 11405 7508 11423 7528
rect 11374 7496 11423 7508
rect 11473 7532 11517 7538
rect 11473 7512 11488 7532
rect 11508 7512 11517 7532
rect 11473 7496 11517 7512
rect 11587 7532 11631 7538
rect 11587 7512 11596 7532
rect 11616 7512 11631 7532
rect 11587 7496 11631 7512
rect 11681 7528 11730 7538
rect 11681 7508 11699 7528
rect 11719 7508 11730 7528
rect 19001 7600 19050 7612
rect 11681 7496 11730 7508
rect 19001 7580 19012 7600
rect 19032 7580 19050 7600
rect 19001 7570 19050 7580
rect 19100 7596 19144 7612
rect 19100 7576 19115 7596
rect 19135 7576 19144 7596
rect 19100 7570 19144 7576
rect 19214 7596 19258 7612
rect 19214 7576 19223 7596
rect 19243 7576 19258 7596
rect 19214 7570 19258 7576
rect 19308 7600 19357 7612
rect 19308 7580 19326 7600
rect 19346 7580 19357 7600
rect 19308 7570 19357 7580
rect 19422 7596 19466 7612
rect 19422 7576 19431 7596
rect 19451 7576 19466 7596
rect 19422 7570 19466 7576
rect 19516 7600 19565 7612
rect 19516 7580 19534 7600
rect 19554 7580 19565 7600
rect 19516 7570 19565 7580
rect 19635 7596 19679 7612
rect 19635 7576 19644 7596
rect 19664 7576 19679 7596
rect 19635 7570 19679 7576
rect 19729 7600 19778 7612
rect 19729 7580 19747 7600
rect 19767 7580 19778 7600
rect 19729 7570 19778 7580
rect 16234 7507 16283 7517
rect 16234 7487 16245 7507
rect 16265 7487 16283 7507
rect 16234 7475 16283 7487
rect 16333 7511 16377 7517
rect 16333 7491 16348 7511
rect 16368 7491 16377 7511
rect 16333 7475 16377 7491
rect 16447 7507 16496 7517
rect 16447 7487 16458 7507
rect 16478 7487 16496 7507
rect 16447 7475 16496 7487
rect 16546 7511 16590 7517
rect 16546 7491 16561 7511
rect 16581 7491 16590 7511
rect 16546 7475 16590 7491
rect 16655 7507 16704 7517
rect 16655 7487 16666 7507
rect 16686 7487 16704 7507
rect 16655 7475 16704 7487
rect 16754 7511 16798 7517
rect 16754 7491 16769 7511
rect 16789 7491 16798 7511
rect 16754 7475 16798 7491
rect 16868 7511 16912 7517
rect 16868 7491 16877 7511
rect 16897 7491 16912 7511
rect 16868 7475 16912 7491
rect 16962 7507 17011 7517
rect 16962 7487 16980 7507
rect 17000 7487 17011 7507
rect 16962 7475 17011 7487
rect 4127 7286 4176 7298
rect 4127 7266 4138 7286
rect 4158 7266 4176 7286
rect 4127 7256 4176 7266
rect 4226 7282 4270 7298
rect 4226 7262 4241 7282
rect 4261 7262 4270 7282
rect 4226 7256 4270 7262
rect 4340 7282 4384 7298
rect 4340 7262 4349 7282
rect 4369 7262 4384 7282
rect 4340 7256 4384 7262
rect 4434 7286 4483 7298
rect 4434 7266 4452 7286
rect 4472 7266 4483 7286
rect 4434 7256 4483 7266
rect 4548 7282 4592 7298
rect 4548 7262 4557 7282
rect 4577 7262 4592 7282
rect 4548 7256 4592 7262
rect 4642 7286 4691 7298
rect 4642 7266 4660 7286
rect 4680 7266 4691 7286
rect 4642 7256 4691 7266
rect 4761 7282 4805 7298
rect 4761 7262 4770 7282
rect 4790 7262 4805 7282
rect 4761 7256 4805 7262
rect 4855 7286 4904 7298
rect 4855 7266 4873 7286
rect 4893 7266 4904 7286
rect 4855 7256 4904 7266
rect 1360 7193 1409 7203
rect 1360 7173 1371 7193
rect 1391 7173 1409 7193
rect 1360 7161 1409 7173
rect 1459 7197 1503 7203
rect 1459 7177 1474 7197
rect 1494 7177 1503 7197
rect 1459 7161 1503 7177
rect 1573 7193 1622 7203
rect 1573 7173 1584 7193
rect 1604 7173 1622 7193
rect 1573 7161 1622 7173
rect 1672 7197 1716 7203
rect 1672 7177 1687 7197
rect 1707 7177 1716 7197
rect 1672 7161 1716 7177
rect 1781 7193 1830 7203
rect 1781 7173 1792 7193
rect 1812 7173 1830 7193
rect 1781 7161 1830 7173
rect 1880 7197 1924 7203
rect 1880 7177 1895 7197
rect 1915 7177 1924 7197
rect 1880 7161 1924 7177
rect 1994 7197 2038 7203
rect 1994 7177 2003 7197
rect 2023 7177 2038 7197
rect 1994 7161 2038 7177
rect 2088 7193 2137 7203
rect 2088 7173 2106 7193
rect 2126 7173 2137 7193
rect 9408 7265 9457 7277
rect 2088 7161 2137 7173
rect 9408 7245 9419 7265
rect 9439 7245 9457 7265
rect 9408 7235 9457 7245
rect 9507 7261 9551 7277
rect 9507 7241 9522 7261
rect 9542 7241 9551 7261
rect 9507 7235 9551 7241
rect 9621 7261 9665 7277
rect 9621 7241 9630 7261
rect 9650 7241 9665 7261
rect 9621 7235 9665 7241
rect 9715 7265 9764 7277
rect 9715 7245 9733 7265
rect 9753 7245 9764 7265
rect 9715 7235 9764 7245
rect 9829 7261 9873 7277
rect 9829 7241 9838 7261
rect 9858 7241 9873 7261
rect 9829 7235 9873 7241
rect 9923 7265 9972 7277
rect 9923 7245 9941 7265
rect 9961 7245 9972 7265
rect 9923 7235 9972 7245
rect 10042 7261 10086 7277
rect 10042 7241 10051 7261
rect 10071 7241 10086 7261
rect 10042 7235 10086 7241
rect 10136 7265 10185 7277
rect 10136 7245 10154 7265
rect 10174 7245 10185 7265
rect 10136 7235 10185 7245
rect 14788 7294 14837 7306
rect 6641 7172 6690 7182
rect 6641 7152 6652 7172
rect 6672 7152 6690 7172
rect 6641 7140 6690 7152
rect 6740 7176 6784 7182
rect 6740 7156 6755 7176
rect 6775 7156 6784 7176
rect 6740 7140 6784 7156
rect 6854 7172 6903 7182
rect 6854 7152 6865 7172
rect 6885 7152 6903 7172
rect 6854 7140 6903 7152
rect 6953 7176 6997 7182
rect 6953 7156 6968 7176
rect 6988 7156 6997 7176
rect 6953 7140 6997 7156
rect 7062 7172 7111 7182
rect 7062 7152 7073 7172
rect 7093 7152 7111 7172
rect 7062 7140 7111 7152
rect 7161 7176 7205 7182
rect 7161 7156 7176 7176
rect 7196 7156 7205 7176
rect 7161 7140 7205 7156
rect 7275 7176 7319 7182
rect 7275 7156 7284 7176
rect 7304 7156 7319 7176
rect 7275 7140 7319 7156
rect 7369 7172 7418 7182
rect 7369 7152 7387 7172
rect 7407 7152 7418 7172
rect 14788 7274 14799 7294
rect 14819 7274 14837 7294
rect 14788 7264 14837 7274
rect 14887 7290 14931 7306
rect 14887 7270 14902 7290
rect 14922 7270 14931 7290
rect 14887 7264 14931 7270
rect 15001 7290 15045 7306
rect 15001 7270 15010 7290
rect 15030 7270 15045 7290
rect 15001 7264 15045 7270
rect 15095 7294 15144 7306
rect 15095 7274 15113 7294
rect 15133 7274 15144 7294
rect 15095 7264 15144 7274
rect 15209 7290 15253 7306
rect 15209 7270 15218 7290
rect 15238 7270 15253 7290
rect 15209 7264 15253 7270
rect 15303 7294 15352 7306
rect 15303 7274 15321 7294
rect 15341 7274 15352 7294
rect 15303 7264 15352 7274
rect 15422 7290 15466 7306
rect 15422 7270 15431 7290
rect 15451 7270 15466 7290
rect 15422 7264 15466 7270
rect 15516 7294 15565 7306
rect 15516 7274 15534 7294
rect 15554 7274 15565 7294
rect 15516 7264 15565 7274
rect 12021 7201 12070 7211
rect 12021 7181 12032 7201
rect 12052 7181 12070 7201
rect 12021 7169 12070 7181
rect 12120 7205 12164 7211
rect 12120 7185 12135 7205
rect 12155 7185 12164 7205
rect 12120 7169 12164 7185
rect 12234 7201 12283 7211
rect 12234 7181 12245 7201
rect 12265 7181 12283 7201
rect 12234 7169 12283 7181
rect 12333 7205 12377 7211
rect 12333 7185 12348 7205
rect 12368 7185 12377 7205
rect 12333 7169 12377 7185
rect 12442 7201 12491 7211
rect 12442 7181 12453 7201
rect 12473 7181 12491 7201
rect 12442 7169 12491 7181
rect 12541 7205 12585 7211
rect 12541 7185 12556 7205
rect 12576 7185 12585 7205
rect 12541 7169 12585 7185
rect 12655 7205 12699 7211
rect 12655 7185 12664 7205
rect 12684 7185 12699 7205
rect 12655 7169 12699 7185
rect 12749 7201 12798 7211
rect 12749 7181 12767 7201
rect 12787 7181 12798 7201
rect 20069 7273 20118 7285
rect 12749 7169 12798 7181
rect 7369 7140 7418 7152
rect 3114 7052 3163 7064
rect 3114 7032 3125 7052
rect 3145 7032 3163 7052
rect 3114 7022 3163 7032
rect 3213 7048 3257 7064
rect 3213 7028 3228 7048
rect 3248 7028 3257 7048
rect 3213 7022 3257 7028
rect 3327 7048 3371 7064
rect 3327 7028 3336 7048
rect 3356 7028 3371 7048
rect 3327 7022 3371 7028
rect 3421 7052 3470 7064
rect 3421 7032 3439 7052
rect 3459 7032 3470 7052
rect 3421 7022 3470 7032
rect 3535 7048 3579 7064
rect 3535 7028 3544 7048
rect 3564 7028 3579 7048
rect 3535 7022 3579 7028
rect 3629 7052 3678 7064
rect 3629 7032 3647 7052
rect 3667 7032 3678 7052
rect 3629 7022 3678 7032
rect 3748 7048 3792 7064
rect 3748 7028 3757 7048
rect 3777 7028 3792 7048
rect 3748 7022 3792 7028
rect 3842 7052 3891 7064
rect 3842 7032 3860 7052
rect 3880 7032 3891 7052
rect 3842 7022 3891 7032
rect 298 6954 347 6964
rect 298 6934 309 6954
rect 329 6934 347 6954
rect 298 6922 347 6934
rect 397 6958 441 6964
rect 397 6938 412 6958
rect 432 6938 441 6958
rect 397 6922 441 6938
rect 511 6954 560 6964
rect 511 6934 522 6954
rect 542 6934 560 6954
rect 511 6922 560 6934
rect 610 6958 654 6964
rect 610 6938 625 6958
rect 645 6938 654 6958
rect 610 6922 654 6938
rect 719 6954 768 6964
rect 719 6934 730 6954
rect 750 6934 768 6954
rect 719 6922 768 6934
rect 818 6958 862 6964
rect 818 6938 833 6958
rect 853 6938 862 6958
rect 818 6922 862 6938
rect 932 6958 976 6964
rect 932 6938 941 6958
rect 961 6938 976 6958
rect 932 6922 976 6938
rect 1026 6954 1075 6964
rect 1026 6934 1044 6954
rect 1064 6934 1075 6954
rect 1026 6922 1075 6934
rect 8395 7031 8444 7043
rect 8395 7011 8406 7031
rect 8426 7011 8444 7031
rect 8395 7001 8444 7011
rect 8494 7027 8538 7043
rect 8494 7007 8509 7027
rect 8529 7007 8538 7027
rect 8494 7001 8538 7007
rect 8608 7027 8652 7043
rect 8608 7007 8617 7027
rect 8637 7007 8652 7027
rect 8608 7001 8652 7007
rect 8702 7031 8751 7043
rect 8702 7011 8720 7031
rect 8740 7011 8751 7031
rect 8702 7001 8751 7011
rect 8816 7027 8860 7043
rect 8816 7007 8825 7027
rect 8845 7007 8860 7027
rect 8816 7001 8860 7007
rect 8910 7031 8959 7043
rect 8910 7011 8928 7031
rect 8948 7011 8959 7031
rect 8910 7001 8959 7011
rect 9029 7027 9073 7043
rect 9029 7007 9038 7027
rect 9058 7007 9073 7027
rect 9029 7001 9073 7007
rect 9123 7031 9172 7043
rect 9123 7011 9141 7031
rect 9161 7011 9172 7031
rect 20069 7253 20080 7273
rect 20100 7253 20118 7273
rect 20069 7243 20118 7253
rect 20168 7269 20212 7285
rect 20168 7249 20183 7269
rect 20203 7249 20212 7269
rect 20168 7243 20212 7249
rect 20282 7269 20326 7285
rect 20282 7249 20291 7269
rect 20311 7249 20326 7269
rect 20282 7243 20326 7249
rect 20376 7273 20425 7285
rect 20376 7253 20394 7273
rect 20414 7253 20425 7273
rect 20376 7243 20425 7253
rect 20490 7269 20534 7285
rect 20490 7249 20499 7269
rect 20519 7249 20534 7269
rect 20490 7243 20534 7249
rect 20584 7273 20633 7285
rect 20584 7253 20602 7273
rect 20622 7253 20633 7273
rect 20584 7243 20633 7253
rect 20703 7269 20747 7285
rect 20703 7249 20712 7269
rect 20732 7249 20747 7269
rect 20703 7243 20747 7249
rect 20797 7273 20846 7285
rect 20797 7253 20815 7273
rect 20835 7253 20846 7273
rect 20797 7243 20846 7253
rect 17302 7180 17351 7190
rect 17302 7160 17313 7180
rect 17333 7160 17351 7180
rect 17302 7148 17351 7160
rect 17401 7184 17445 7190
rect 17401 7164 17416 7184
rect 17436 7164 17445 7184
rect 17401 7148 17445 7164
rect 17515 7180 17564 7190
rect 17515 7160 17526 7180
rect 17546 7160 17564 7180
rect 17515 7148 17564 7160
rect 17614 7184 17658 7190
rect 17614 7164 17629 7184
rect 17649 7164 17658 7184
rect 17614 7148 17658 7164
rect 17723 7180 17772 7190
rect 17723 7160 17734 7180
rect 17754 7160 17772 7180
rect 17723 7148 17772 7160
rect 17822 7184 17866 7190
rect 17822 7164 17837 7184
rect 17857 7164 17866 7184
rect 17822 7148 17866 7164
rect 17936 7184 17980 7190
rect 17936 7164 17945 7184
rect 17965 7164 17980 7184
rect 17936 7148 17980 7164
rect 18030 7180 18079 7190
rect 18030 7160 18048 7180
rect 18068 7160 18079 7180
rect 18030 7148 18079 7160
rect 13775 7060 13824 7072
rect 9123 7001 9172 7011
rect 5579 6933 5628 6943
rect 5579 6913 5590 6933
rect 5610 6913 5628 6933
rect 5579 6901 5628 6913
rect 5678 6937 5722 6943
rect 5678 6917 5693 6937
rect 5713 6917 5722 6937
rect 5678 6901 5722 6917
rect 5792 6933 5841 6943
rect 5792 6913 5803 6933
rect 5823 6913 5841 6933
rect 5792 6901 5841 6913
rect 5891 6937 5935 6943
rect 5891 6917 5906 6937
rect 5926 6917 5935 6937
rect 5891 6901 5935 6917
rect 6000 6933 6049 6943
rect 6000 6913 6011 6933
rect 6031 6913 6049 6933
rect 6000 6901 6049 6913
rect 6099 6937 6143 6943
rect 6099 6917 6114 6937
rect 6134 6917 6143 6937
rect 6099 6901 6143 6917
rect 6213 6937 6257 6943
rect 6213 6917 6222 6937
rect 6242 6917 6257 6937
rect 6213 6901 6257 6917
rect 6307 6933 6356 6943
rect 6307 6913 6325 6933
rect 6345 6913 6356 6933
rect 6307 6901 6356 6913
rect 4126 6871 4175 6883
rect 4126 6851 4137 6871
rect 4157 6851 4175 6871
rect 4126 6841 4175 6851
rect 4225 6867 4269 6883
rect 4225 6847 4240 6867
rect 4260 6847 4269 6867
rect 4225 6841 4269 6847
rect 4339 6867 4383 6883
rect 4339 6847 4348 6867
rect 4368 6847 4383 6867
rect 4339 6841 4383 6847
rect 4433 6871 4482 6883
rect 4433 6851 4451 6871
rect 4471 6851 4482 6871
rect 4433 6841 4482 6851
rect 4547 6867 4591 6883
rect 4547 6847 4556 6867
rect 4576 6847 4591 6867
rect 4547 6841 4591 6847
rect 4641 6871 4690 6883
rect 4641 6851 4659 6871
rect 4679 6851 4690 6871
rect 4641 6841 4690 6851
rect 4760 6867 4804 6883
rect 4760 6847 4769 6867
rect 4789 6847 4804 6867
rect 4760 6841 4804 6847
rect 4854 6871 4903 6883
rect 4854 6851 4872 6871
rect 4892 6851 4903 6871
rect 4854 6841 4903 6851
rect 1310 6773 1359 6783
rect 1310 6753 1321 6773
rect 1341 6753 1359 6773
rect 1310 6741 1359 6753
rect 1409 6777 1453 6783
rect 1409 6757 1424 6777
rect 1444 6757 1453 6777
rect 1409 6741 1453 6757
rect 1523 6773 1572 6783
rect 1523 6753 1534 6773
rect 1554 6753 1572 6773
rect 1523 6741 1572 6753
rect 1622 6777 1666 6783
rect 1622 6757 1637 6777
rect 1657 6757 1666 6777
rect 1622 6741 1666 6757
rect 1731 6773 1780 6783
rect 1731 6753 1742 6773
rect 1762 6753 1780 6773
rect 1731 6741 1780 6753
rect 1830 6777 1874 6783
rect 1830 6757 1845 6777
rect 1865 6757 1874 6777
rect 1830 6741 1874 6757
rect 1944 6777 1988 6783
rect 1944 6757 1953 6777
rect 1973 6757 1988 6777
rect 1944 6741 1988 6757
rect 2038 6773 2087 6783
rect 2038 6753 2056 6773
rect 2076 6753 2087 6773
rect 13775 7040 13786 7060
rect 13806 7040 13824 7060
rect 13775 7030 13824 7040
rect 13874 7056 13918 7072
rect 13874 7036 13889 7056
rect 13909 7036 13918 7056
rect 13874 7030 13918 7036
rect 13988 7056 14032 7072
rect 13988 7036 13997 7056
rect 14017 7036 14032 7056
rect 13988 7030 14032 7036
rect 14082 7060 14131 7072
rect 14082 7040 14100 7060
rect 14120 7040 14131 7060
rect 14082 7030 14131 7040
rect 14196 7056 14240 7072
rect 14196 7036 14205 7056
rect 14225 7036 14240 7056
rect 14196 7030 14240 7036
rect 14290 7060 14339 7072
rect 14290 7040 14308 7060
rect 14328 7040 14339 7060
rect 14290 7030 14339 7040
rect 14409 7056 14453 7072
rect 14409 7036 14418 7056
rect 14438 7036 14453 7056
rect 14409 7030 14453 7036
rect 14503 7060 14552 7072
rect 14503 7040 14521 7060
rect 14541 7040 14552 7060
rect 14503 7030 14552 7040
rect 10959 6962 11008 6972
rect 10959 6942 10970 6962
rect 10990 6942 11008 6962
rect 10959 6930 11008 6942
rect 11058 6966 11102 6972
rect 11058 6946 11073 6966
rect 11093 6946 11102 6966
rect 11058 6930 11102 6946
rect 11172 6962 11221 6972
rect 11172 6942 11183 6962
rect 11203 6942 11221 6962
rect 11172 6930 11221 6942
rect 11271 6966 11315 6972
rect 11271 6946 11286 6966
rect 11306 6946 11315 6966
rect 11271 6930 11315 6946
rect 11380 6962 11429 6972
rect 11380 6942 11391 6962
rect 11411 6942 11429 6962
rect 11380 6930 11429 6942
rect 11479 6966 11523 6972
rect 11479 6946 11494 6966
rect 11514 6946 11523 6966
rect 11479 6930 11523 6946
rect 11593 6966 11637 6972
rect 11593 6946 11602 6966
rect 11622 6946 11637 6966
rect 11593 6930 11637 6946
rect 11687 6962 11736 6972
rect 11687 6942 11705 6962
rect 11725 6942 11736 6962
rect 11687 6930 11736 6942
rect 2038 6741 2087 6753
rect 19056 7039 19105 7051
rect 9407 6850 9456 6862
rect 9407 6830 9418 6850
rect 9438 6830 9456 6850
rect 9407 6820 9456 6830
rect 9506 6846 9550 6862
rect 9506 6826 9521 6846
rect 9541 6826 9550 6846
rect 9506 6820 9550 6826
rect 9620 6846 9664 6862
rect 9620 6826 9629 6846
rect 9649 6826 9664 6846
rect 9620 6820 9664 6826
rect 9714 6850 9763 6862
rect 9714 6830 9732 6850
rect 9752 6830 9763 6850
rect 9714 6820 9763 6830
rect 9828 6846 9872 6862
rect 9828 6826 9837 6846
rect 9857 6826 9872 6846
rect 9828 6820 9872 6826
rect 9922 6850 9971 6862
rect 9922 6830 9940 6850
rect 9960 6830 9971 6850
rect 9922 6820 9971 6830
rect 10041 6846 10085 6862
rect 10041 6826 10050 6846
rect 10070 6826 10085 6846
rect 10041 6820 10085 6826
rect 10135 6850 10184 6862
rect 10135 6830 10153 6850
rect 10173 6830 10184 6850
rect 10135 6820 10184 6830
rect 6591 6752 6640 6762
rect 6591 6732 6602 6752
rect 6622 6732 6640 6752
rect 6591 6720 6640 6732
rect 6690 6756 6734 6762
rect 6690 6736 6705 6756
rect 6725 6736 6734 6756
rect 6690 6720 6734 6736
rect 6804 6752 6853 6762
rect 6804 6732 6815 6752
rect 6835 6732 6853 6752
rect 6804 6720 6853 6732
rect 6903 6756 6947 6762
rect 6903 6736 6918 6756
rect 6938 6736 6947 6756
rect 6903 6720 6947 6736
rect 7012 6752 7061 6762
rect 7012 6732 7023 6752
rect 7043 6732 7061 6752
rect 7012 6720 7061 6732
rect 7111 6756 7155 6762
rect 7111 6736 7126 6756
rect 7146 6736 7155 6756
rect 7111 6720 7155 6736
rect 7225 6756 7269 6762
rect 7225 6736 7234 6756
rect 7254 6736 7269 6756
rect 7225 6720 7269 6736
rect 7319 6752 7368 6762
rect 7319 6732 7337 6752
rect 7357 6732 7368 6752
rect 19056 7019 19067 7039
rect 19087 7019 19105 7039
rect 19056 7009 19105 7019
rect 19155 7035 19199 7051
rect 19155 7015 19170 7035
rect 19190 7015 19199 7035
rect 19155 7009 19199 7015
rect 19269 7035 19313 7051
rect 19269 7015 19278 7035
rect 19298 7015 19313 7035
rect 19269 7009 19313 7015
rect 19363 7039 19412 7051
rect 19363 7019 19381 7039
rect 19401 7019 19412 7039
rect 19363 7009 19412 7019
rect 19477 7035 19521 7051
rect 19477 7015 19486 7035
rect 19506 7015 19521 7035
rect 19477 7009 19521 7015
rect 19571 7039 19620 7051
rect 19571 7019 19589 7039
rect 19609 7019 19620 7039
rect 19571 7009 19620 7019
rect 19690 7035 19734 7051
rect 19690 7015 19699 7035
rect 19719 7015 19734 7035
rect 19690 7009 19734 7015
rect 19784 7039 19833 7051
rect 19784 7019 19802 7039
rect 19822 7019 19833 7039
rect 19784 7009 19833 7019
rect 16240 6941 16289 6951
rect 16240 6921 16251 6941
rect 16271 6921 16289 6941
rect 16240 6909 16289 6921
rect 16339 6945 16383 6951
rect 16339 6925 16354 6945
rect 16374 6925 16383 6945
rect 16339 6909 16383 6925
rect 16453 6941 16502 6951
rect 16453 6921 16464 6941
rect 16484 6921 16502 6941
rect 16453 6909 16502 6921
rect 16552 6945 16596 6951
rect 16552 6925 16567 6945
rect 16587 6925 16596 6945
rect 16552 6909 16596 6925
rect 16661 6941 16710 6951
rect 16661 6921 16672 6941
rect 16692 6921 16710 6941
rect 16661 6909 16710 6921
rect 16760 6945 16804 6951
rect 16760 6925 16775 6945
rect 16795 6925 16804 6945
rect 16760 6909 16804 6925
rect 16874 6945 16918 6951
rect 16874 6925 16883 6945
rect 16903 6925 16918 6945
rect 16874 6909 16918 6925
rect 16968 6941 17017 6951
rect 16968 6921 16986 6941
rect 17006 6921 17017 6941
rect 16968 6909 17017 6921
rect 14787 6879 14836 6891
rect 14787 6859 14798 6879
rect 14818 6859 14836 6879
rect 14787 6849 14836 6859
rect 14886 6875 14930 6891
rect 14886 6855 14901 6875
rect 14921 6855 14930 6875
rect 14886 6849 14930 6855
rect 15000 6875 15044 6891
rect 15000 6855 15009 6875
rect 15029 6855 15044 6875
rect 15000 6849 15044 6855
rect 15094 6879 15143 6891
rect 15094 6859 15112 6879
rect 15132 6859 15143 6879
rect 15094 6849 15143 6859
rect 15208 6875 15252 6891
rect 15208 6855 15217 6875
rect 15237 6855 15252 6875
rect 15208 6849 15252 6855
rect 15302 6879 15351 6891
rect 15302 6859 15320 6879
rect 15340 6859 15351 6879
rect 15302 6849 15351 6859
rect 15421 6875 15465 6891
rect 15421 6855 15430 6875
rect 15450 6855 15465 6875
rect 15421 6849 15465 6855
rect 15515 6879 15564 6891
rect 15515 6859 15533 6879
rect 15553 6859 15564 6879
rect 15515 6849 15564 6859
rect 11971 6781 12020 6791
rect 7319 6720 7368 6732
rect 2906 6585 2955 6597
rect 2906 6565 2917 6585
rect 2937 6565 2955 6585
rect 2906 6555 2955 6565
rect 3005 6581 3049 6597
rect 3005 6561 3020 6581
rect 3040 6561 3049 6581
rect 3005 6555 3049 6561
rect 3119 6581 3163 6597
rect 3119 6561 3128 6581
rect 3148 6561 3163 6581
rect 3119 6555 3163 6561
rect 3213 6585 3262 6597
rect 3213 6565 3231 6585
rect 3251 6565 3262 6585
rect 3213 6555 3262 6565
rect 3327 6581 3371 6597
rect 3327 6561 3336 6581
rect 3356 6561 3371 6581
rect 3327 6555 3371 6561
rect 3421 6585 3470 6597
rect 3421 6565 3439 6585
rect 3459 6565 3470 6585
rect 3421 6555 3470 6565
rect 3540 6581 3584 6597
rect 3540 6561 3549 6581
rect 3569 6561 3584 6581
rect 3540 6555 3584 6561
rect 3634 6585 3683 6597
rect 3634 6565 3652 6585
rect 3672 6565 3683 6585
rect 3634 6555 3683 6565
rect 11971 6761 11982 6781
rect 12002 6761 12020 6781
rect 11971 6749 12020 6761
rect 12070 6785 12114 6791
rect 12070 6765 12085 6785
rect 12105 6765 12114 6785
rect 12070 6749 12114 6765
rect 12184 6781 12233 6791
rect 12184 6761 12195 6781
rect 12215 6761 12233 6781
rect 12184 6749 12233 6761
rect 12283 6785 12327 6791
rect 12283 6765 12298 6785
rect 12318 6765 12327 6785
rect 12283 6749 12327 6765
rect 12392 6781 12441 6791
rect 12392 6761 12403 6781
rect 12423 6761 12441 6781
rect 12392 6749 12441 6761
rect 12491 6785 12535 6791
rect 12491 6765 12506 6785
rect 12526 6765 12535 6785
rect 12491 6749 12535 6765
rect 12605 6785 12649 6791
rect 12605 6765 12614 6785
rect 12634 6765 12649 6785
rect 12605 6749 12649 6765
rect 12699 6781 12748 6791
rect 12699 6761 12717 6781
rect 12737 6761 12748 6781
rect 12699 6749 12748 6761
rect 20068 6858 20117 6870
rect 20068 6838 20079 6858
rect 20099 6838 20117 6858
rect 20068 6828 20117 6838
rect 20167 6854 20211 6870
rect 20167 6834 20182 6854
rect 20202 6834 20211 6854
rect 20167 6828 20211 6834
rect 20281 6854 20325 6870
rect 20281 6834 20290 6854
rect 20310 6834 20325 6854
rect 20281 6828 20325 6834
rect 20375 6858 20424 6870
rect 20375 6838 20393 6858
rect 20413 6838 20424 6858
rect 20375 6828 20424 6838
rect 20489 6854 20533 6870
rect 20489 6834 20498 6854
rect 20518 6834 20533 6854
rect 20489 6828 20533 6834
rect 20583 6858 20632 6870
rect 20583 6838 20601 6858
rect 20621 6838 20632 6858
rect 20583 6828 20632 6838
rect 20702 6854 20746 6870
rect 20702 6834 20711 6854
rect 20731 6834 20746 6854
rect 20702 6828 20746 6834
rect 20796 6858 20845 6870
rect 20796 6838 20814 6858
rect 20834 6838 20845 6858
rect 20796 6828 20845 6838
rect 17252 6760 17301 6770
rect 17252 6740 17263 6760
rect 17283 6740 17301 6760
rect 17252 6728 17301 6740
rect 17351 6764 17395 6770
rect 17351 6744 17366 6764
rect 17386 6744 17395 6764
rect 17351 6728 17395 6744
rect 17465 6760 17514 6770
rect 17465 6740 17476 6760
rect 17496 6740 17514 6760
rect 17465 6728 17514 6740
rect 17564 6764 17608 6770
rect 17564 6744 17579 6764
rect 17599 6744 17608 6764
rect 17564 6728 17608 6744
rect 17673 6760 17722 6770
rect 17673 6740 17684 6760
rect 17704 6740 17722 6760
rect 17673 6728 17722 6740
rect 17772 6764 17816 6770
rect 17772 6744 17787 6764
rect 17807 6744 17816 6764
rect 17772 6728 17816 6744
rect 17886 6764 17930 6770
rect 17886 6744 17895 6764
rect 17915 6744 17930 6764
rect 17886 6728 17930 6744
rect 17980 6760 18029 6770
rect 17980 6740 17998 6760
rect 18018 6740 18029 6760
rect 17980 6728 18029 6740
rect 297 6539 346 6549
rect 297 6519 308 6539
rect 328 6519 346 6539
rect 297 6507 346 6519
rect 396 6543 440 6549
rect 396 6523 411 6543
rect 431 6523 440 6543
rect 396 6507 440 6523
rect 510 6539 559 6549
rect 510 6519 521 6539
rect 541 6519 559 6539
rect 510 6507 559 6519
rect 609 6543 653 6549
rect 609 6523 624 6543
rect 644 6523 653 6543
rect 609 6507 653 6523
rect 718 6539 767 6549
rect 718 6519 729 6539
rect 749 6519 767 6539
rect 718 6507 767 6519
rect 817 6543 861 6549
rect 817 6523 832 6543
rect 852 6523 861 6543
rect 817 6507 861 6523
rect 931 6543 975 6549
rect 931 6523 940 6543
rect 960 6523 975 6543
rect 931 6507 975 6523
rect 1025 6539 1074 6549
rect 1025 6519 1043 6539
rect 1063 6519 1074 6539
rect 1025 6507 1074 6519
rect 8187 6564 8236 6576
rect 8187 6544 8198 6564
rect 8218 6544 8236 6564
rect 8187 6534 8236 6544
rect 8286 6560 8330 6576
rect 8286 6540 8301 6560
rect 8321 6540 8330 6560
rect 8286 6534 8330 6540
rect 8400 6560 8444 6576
rect 8400 6540 8409 6560
rect 8429 6540 8444 6560
rect 8400 6534 8444 6540
rect 8494 6564 8543 6576
rect 8494 6544 8512 6564
rect 8532 6544 8543 6564
rect 8494 6534 8543 6544
rect 8608 6560 8652 6576
rect 8608 6540 8617 6560
rect 8637 6540 8652 6560
rect 8608 6534 8652 6540
rect 8702 6564 8751 6576
rect 8702 6544 8720 6564
rect 8740 6544 8751 6564
rect 8702 6534 8751 6544
rect 8821 6560 8865 6576
rect 8821 6540 8830 6560
rect 8850 6540 8865 6560
rect 8821 6534 8865 6540
rect 8915 6564 8964 6576
rect 8915 6544 8933 6564
rect 8953 6544 8964 6564
rect 8915 6534 8964 6544
rect 5578 6518 5627 6528
rect 5578 6498 5589 6518
rect 5609 6498 5627 6518
rect 5578 6486 5627 6498
rect 5677 6522 5721 6528
rect 5677 6502 5692 6522
rect 5712 6502 5721 6522
rect 5677 6486 5721 6502
rect 5791 6518 5840 6528
rect 5791 6498 5802 6518
rect 5822 6498 5840 6518
rect 5791 6486 5840 6498
rect 5890 6522 5934 6528
rect 5890 6502 5905 6522
rect 5925 6502 5934 6522
rect 5890 6486 5934 6502
rect 5999 6518 6048 6528
rect 5999 6498 6010 6518
rect 6030 6498 6048 6518
rect 5999 6486 6048 6498
rect 6098 6522 6142 6528
rect 6098 6502 6113 6522
rect 6133 6502 6142 6522
rect 6098 6486 6142 6502
rect 6212 6522 6256 6528
rect 6212 6502 6221 6522
rect 6241 6502 6256 6522
rect 6212 6486 6256 6502
rect 6306 6518 6355 6528
rect 6306 6498 6324 6518
rect 6344 6498 6355 6518
rect 6306 6486 6355 6498
rect 13567 6593 13616 6605
rect 13567 6573 13578 6593
rect 13598 6573 13616 6593
rect 13567 6563 13616 6573
rect 13666 6589 13710 6605
rect 13666 6569 13681 6589
rect 13701 6569 13710 6589
rect 13666 6563 13710 6569
rect 13780 6589 13824 6605
rect 13780 6569 13789 6589
rect 13809 6569 13824 6589
rect 13780 6563 13824 6569
rect 13874 6593 13923 6605
rect 13874 6573 13892 6593
rect 13912 6573 13923 6593
rect 13874 6563 13923 6573
rect 13988 6589 14032 6605
rect 13988 6569 13997 6589
rect 14017 6569 14032 6589
rect 13988 6563 14032 6569
rect 14082 6593 14131 6605
rect 14082 6573 14100 6593
rect 14120 6573 14131 6593
rect 14082 6563 14131 6573
rect 14201 6589 14245 6605
rect 14201 6569 14210 6589
rect 14230 6569 14245 6589
rect 14201 6563 14245 6569
rect 14295 6593 14344 6605
rect 14295 6573 14313 6593
rect 14333 6573 14344 6593
rect 14295 6563 14344 6573
rect 10958 6547 11007 6557
rect 10958 6527 10969 6547
rect 10989 6527 11007 6547
rect 10958 6515 11007 6527
rect 11057 6551 11101 6557
rect 11057 6531 11072 6551
rect 11092 6531 11101 6551
rect 11057 6515 11101 6531
rect 11171 6547 11220 6557
rect 11171 6527 11182 6547
rect 11202 6527 11220 6547
rect 11171 6515 11220 6527
rect 11270 6551 11314 6557
rect 11270 6531 11285 6551
rect 11305 6531 11314 6551
rect 11270 6515 11314 6531
rect 11379 6547 11428 6557
rect 11379 6527 11390 6547
rect 11410 6527 11428 6547
rect 11379 6515 11428 6527
rect 11478 6551 11522 6557
rect 11478 6531 11493 6551
rect 11513 6531 11522 6551
rect 11478 6515 11522 6531
rect 11592 6551 11636 6557
rect 11592 6531 11601 6551
rect 11621 6531 11636 6551
rect 11592 6515 11636 6531
rect 11686 6547 11735 6557
rect 11686 6527 11704 6547
rect 11724 6527 11735 6547
rect 11686 6515 11735 6527
rect 18848 6572 18897 6584
rect 18848 6552 18859 6572
rect 18879 6552 18897 6572
rect 18848 6542 18897 6552
rect 18947 6568 18991 6584
rect 18947 6548 18962 6568
rect 18982 6548 18991 6568
rect 18947 6542 18991 6548
rect 19061 6568 19105 6584
rect 19061 6548 19070 6568
rect 19090 6548 19105 6568
rect 19061 6542 19105 6548
rect 19155 6572 19204 6584
rect 19155 6552 19173 6572
rect 19193 6552 19204 6572
rect 19155 6542 19204 6552
rect 19269 6568 19313 6584
rect 19269 6548 19278 6568
rect 19298 6548 19313 6568
rect 19269 6542 19313 6548
rect 19363 6572 19412 6584
rect 19363 6552 19381 6572
rect 19401 6552 19412 6572
rect 19363 6542 19412 6552
rect 19482 6568 19526 6584
rect 19482 6548 19491 6568
rect 19511 6548 19526 6568
rect 19482 6542 19526 6548
rect 19576 6572 19625 6584
rect 19576 6552 19594 6572
rect 19614 6552 19625 6572
rect 19576 6542 19625 6552
rect 4134 6307 4183 6319
rect 4134 6287 4145 6307
rect 4165 6287 4183 6307
rect 4134 6277 4183 6287
rect 4233 6303 4277 6319
rect 4233 6283 4248 6303
rect 4268 6283 4277 6303
rect 4233 6277 4277 6283
rect 4347 6303 4391 6319
rect 4347 6283 4356 6303
rect 4376 6283 4391 6303
rect 4347 6277 4391 6283
rect 4441 6307 4490 6319
rect 4441 6287 4459 6307
rect 4479 6287 4490 6307
rect 4441 6277 4490 6287
rect 4555 6303 4599 6319
rect 4555 6283 4564 6303
rect 4584 6283 4599 6303
rect 4555 6277 4599 6283
rect 4649 6307 4698 6319
rect 4649 6287 4667 6307
rect 4687 6287 4698 6307
rect 4649 6277 4698 6287
rect 4768 6303 4812 6319
rect 4768 6283 4777 6303
rect 4797 6283 4812 6303
rect 4768 6277 4812 6283
rect 4862 6307 4911 6319
rect 4862 6287 4880 6307
rect 4900 6287 4911 6307
rect 4862 6277 4911 6287
rect 16239 6526 16288 6536
rect 16239 6506 16250 6526
rect 16270 6506 16288 6526
rect 16239 6494 16288 6506
rect 16338 6530 16382 6536
rect 16338 6510 16353 6530
rect 16373 6510 16382 6530
rect 16338 6494 16382 6510
rect 16452 6526 16501 6536
rect 16452 6506 16463 6526
rect 16483 6506 16501 6526
rect 16452 6494 16501 6506
rect 16551 6530 16595 6536
rect 16551 6510 16566 6530
rect 16586 6510 16595 6530
rect 16551 6494 16595 6510
rect 16660 6526 16709 6536
rect 16660 6506 16671 6526
rect 16691 6506 16709 6526
rect 16660 6494 16709 6506
rect 16759 6530 16803 6536
rect 16759 6510 16774 6530
rect 16794 6510 16803 6530
rect 16759 6494 16803 6510
rect 16873 6530 16917 6536
rect 16873 6510 16882 6530
rect 16902 6510 16917 6530
rect 16873 6494 16917 6510
rect 16967 6526 17016 6536
rect 16967 6506 16985 6526
rect 17005 6506 17016 6526
rect 16967 6494 17016 6506
rect 1525 6261 1574 6271
rect 1525 6241 1536 6261
rect 1556 6241 1574 6261
rect 1525 6229 1574 6241
rect 1624 6265 1668 6271
rect 1624 6245 1639 6265
rect 1659 6245 1668 6265
rect 1624 6229 1668 6245
rect 1738 6261 1787 6271
rect 1738 6241 1749 6261
rect 1769 6241 1787 6261
rect 1738 6229 1787 6241
rect 1837 6265 1881 6271
rect 1837 6245 1852 6265
rect 1872 6245 1881 6265
rect 1837 6229 1881 6245
rect 1946 6261 1995 6271
rect 1946 6241 1957 6261
rect 1977 6241 1995 6261
rect 1946 6229 1995 6241
rect 2045 6265 2089 6271
rect 2045 6245 2060 6265
rect 2080 6245 2089 6265
rect 2045 6229 2089 6245
rect 2159 6265 2203 6271
rect 2159 6245 2168 6265
rect 2188 6245 2203 6265
rect 2159 6229 2203 6245
rect 2253 6261 2302 6271
rect 2253 6241 2271 6261
rect 2291 6241 2302 6261
rect 2253 6229 2302 6241
rect 9415 6286 9464 6298
rect 9415 6266 9426 6286
rect 9446 6266 9464 6286
rect 9415 6256 9464 6266
rect 9514 6282 9558 6298
rect 9514 6262 9529 6282
rect 9549 6262 9558 6282
rect 9514 6256 9558 6262
rect 9628 6282 9672 6298
rect 9628 6262 9637 6282
rect 9657 6262 9672 6282
rect 9628 6256 9672 6262
rect 9722 6286 9771 6298
rect 9722 6266 9740 6286
rect 9760 6266 9771 6286
rect 9722 6256 9771 6266
rect 9836 6282 9880 6298
rect 9836 6262 9845 6282
rect 9865 6262 9880 6282
rect 9836 6256 9880 6262
rect 9930 6286 9979 6298
rect 9930 6266 9948 6286
rect 9968 6266 9979 6286
rect 9930 6256 9979 6266
rect 10049 6282 10093 6298
rect 10049 6262 10058 6282
rect 10078 6262 10093 6282
rect 10049 6256 10093 6262
rect 10143 6286 10192 6298
rect 10143 6266 10161 6286
rect 10181 6266 10192 6286
rect 10143 6256 10192 6266
rect 6806 6240 6855 6250
rect 6806 6220 6817 6240
rect 6837 6220 6855 6240
rect 6806 6208 6855 6220
rect 6905 6244 6949 6250
rect 6905 6224 6920 6244
rect 6940 6224 6949 6244
rect 6905 6208 6949 6224
rect 7019 6240 7068 6250
rect 7019 6220 7030 6240
rect 7050 6220 7068 6240
rect 7019 6208 7068 6220
rect 7118 6244 7162 6250
rect 7118 6224 7133 6244
rect 7153 6224 7162 6244
rect 7118 6208 7162 6224
rect 7227 6240 7276 6250
rect 7227 6220 7238 6240
rect 7258 6220 7276 6240
rect 7227 6208 7276 6220
rect 7326 6244 7370 6250
rect 7326 6224 7341 6244
rect 7361 6224 7370 6244
rect 7326 6208 7370 6224
rect 7440 6244 7484 6250
rect 7440 6224 7449 6244
rect 7469 6224 7484 6244
rect 7440 6208 7484 6224
rect 7534 6240 7583 6250
rect 7534 6220 7552 6240
rect 7572 6220 7583 6240
rect 7534 6208 7583 6220
rect 14795 6315 14844 6327
rect 14795 6295 14806 6315
rect 14826 6295 14844 6315
rect 14795 6285 14844 6295
rect 14894 6311 14938 6327
rect 14894 6291 14909 6311
rect 14929 6291 14938 6311
rect 14894 6285 14938 6291
rect 15008 6311 15052 6327
rect 15008 6291 15017 6311
rect 15037 6291 15052 6311
rect 15008 6285 15052 6291
rect 15102 6315 15151 6327
rect 15102 6295 15120 6315
rect 15140 6295 15151 6315
rect 15102 6285 15151 6295
rect 15216 6311 15260 6327
rect 15216 6291 15225 6311
rect 15245 6291 15260 6311
rect 15216 6285 15260 6291
rect 15310 6315 15359 6327
rect 15310 6295 15328 6315
rect 15348 6295 15359 6315
rect 15310 6285 15359 6295
rect 15429 6311 15473 6327
rect 15429 6291 15438 6311
rect 15458 6291 15473 6311
rect 15429 6285 15473 6291
rect 15523 6315 15572 6327
rect 15523 6295 15541 6315
rect 15561 6295 15572 6315
rect 15523 6285 15572 6295
rect 12186 6269 12235 6279
rect 12186 6249 12197 6269
rect 12217 6249 12235 6269
rect 12186 6237 12235 6249
rect 12285 6273 12329 6279
rect 12285 6253 12300 6273
rect 12320 6253 12329 6273
rect 12285 6237 12329 6253
rect 12399 6269 12448 6279
rect 12399 6249 12410 6269
rect 12430 6249 12448 6269
rect 12399 6237 12448 6249
rect 12498 6273 12542 6279
rect 12498 6253 12513 6273
rect 12533 6253 12542 6273
rect 12498 6237 12542 6253
rect 12607 6269 12656 6279
rect 12607 6249 12618 6269
rect 12638 6249 12656 6269
rect 12607 6237 12656 6249
rect 12706 6273 12750 6279
rect 12706 6253 12721 6273
rect 12741 6253 12750 6273
rect 12706 6237 12750 6253
rect 12820 6273 12864 6279
rect 12820 6253 12829 6273
rect 12849 6253 12864 6273
rect 12820 6237 12864 6253
rect 12914 6269 12963 6279
rect 12914 6249 12932 6269
rect 12952 6249 12963 6269
rect 12914 6237 12963 6249
rect 20076 6294 20125 6306
rect 20076 6274 20087 6294
rect 20107 6274 20125 6294
rect 20076 6264 20125 6274
rect 20175 6290 20219 6306
rect 20175 6270 20190 6290
rect 20210 6270 20219 6290
rect 20175 6264 20219 6270
rect 20289 6290 20333 6306
rect 20289 6270 20298 6290
rect 20318 6270 20333 6290
rect 20289 6264 20333 6270
rect 20383 6294 20432 6306
rect 20383 6274 20401 6294
rect 20421 6274 20432 6294
rect 20383 6264 20432 6274
rect 20497 6290 20541 6306
rect 20497 6270 20506 6290
rect 20526 6270 20541 6290
rect 20497 6264 20541 6270
rect 20591 6294 20640 6306
rect 20591 6274 20609 6294
rect 20629 6274 20640 6294
rect 20591 6264 20640 6274
rect 20710 6290 20754 6306
rect 20710 6270 20719 6290
rect 20739 6270 20754 6290
rect 20710 6264 20754 6270
rect 20804 6294 20853 6306
rect 20804 6274 20822 6294
rect 20842 6274 20853 6294
rect 20804 6264 20853 6274
rect 3121 6073 3170 6085
rect 3121 6053 3132 6073
rect 3152 6053 3170 6073
rect 3121 6043 3170 6053
rect 3220 6069 3264 6085
rect 3220 6049 3235 6069
rect 3255 6049 3264 6069
rect 3220 6043 3264 6049
rect 3334 6069 3378 6085
rect 3334 6049 3343 6069
rect 3363 6049 3378 6069
rect 3334 6043 3378 6049
rect 3428 6073 3477 6085
rect 3428 6053 3446 6073
rect 3466 6053 3477 6073
rect 3428 6043 3477 6053
rect 3542 6069 3586 6085
rect 3542 6049 3551 6069
rect 3571 6049 3586 6069
rect 3542 6043 3586 6049
rect 3636 6073 3685 6085
rect 3636 6053 3654 6073
rect 3674 6053 3685 6073
rect 3636 6043 3685 6053
rect 3755 6069 3799 6085
rect 3755 6049 3764 6069
rect 3784 6049 3799 6069
rect 3755 6043 3799 6049
rect 3849 6073 3898 6085
rect 3849 6053 3867 6073
rect 3887 6053 3898 6073
rect 3849 6043 3898 6053
rect 305 5975 354 5985
rect 305 5955 316 5975
rect 336 5955 354 5975
rect 305 5943 354 5955
rect 404 5979 448 5985
rect 404 5959 419 5979
rect 439 5959 448 5979
rect 404 5943 448 5959
rect 518 5975 567 5985
rect 518 5955 529 5975
rect 549 5955 567 5975
rect 518 5943 567 5955
rect 617 5979 661 5985
rect 617 5959 632 5979
rect 652 5959 661 5979
rect 617 5943 661 5959
rect 726 5975 775 5985
rect 726 5955 737 5975
rect 757 5955 775 5975
rect 726 5943 775 5955
rect 825 5979 869 5985
rect 825 5959 840 5979
rect 860 5959 869 5979
rect 825 5943 869 5959
rect 939 5979 983 5985
rect 939 5959 948 5979
rect 968 5959 983 5979
rect 939 5943 983 5959
rect 1033 5975 1082 5985
rect 1033 5955 1051 5975
rect 1071 5955 1082 5975
rect 1033 5943 1082 5955
rect 8402 6052 8451 6064
rect 8402 6032 8413 6052
rect 8433 6032 8451 6052
rect 8402 6022 8451 6032
rect 8501 6048 8545 6064
rect 8501 6028 8516 6048
rect 8536 6028 8545 6048
rect 8501 6022 8545 6028
rect 8615 6048 8659 6064
rect 8615 6028 8624 6048
rect 8644 6028 8659 6048
rect 8615 6022 8659 6028
rect 8709 6052 8758 6064
rect 8709 6032 8727 6052
rect 8747 6032 8758 6052
rect 8709 6022 8758 6032
rect 8823 6048 8867 6064
rect 8823 6028 8832 6048
rect 8852 6028 8867 6048
rect 8823 6022 8867 6028
rect 8917 6052 8966 6064
rect 8917 6032 8935 6052
rect 8955 6032 8966 6052
rect 8917 6022 8966 6032
rect 9036 6048 9080 6064
rect 9036 6028 9045 6048
rect 9065 6028 9080 6048
rect 9036 6022 9080 6028
rect 9130 6052 9179 6064
rect 9130 6032 9148 6052
rect 9168 6032 9179 6052
rect 17467 6248 17516 6258
rect 17467 6228 17478 6248
rect 17498 6228 17516 6248
rect 17467 6216 17516 6228
rect 17566 6252 17610 6258
rect 17566 6232 17581 6252
rect 17601 6232 17610 6252
rect 17566 6216 17610 6232
rect 17680 6248 17729 6258
rect 17680 6228 17691 6248
rect 17711 6228 17729 6248
rect 17680 6216 17729 6228
rect 17779 6252 17823 6258
rect 17779 6232 17794 6252
rect 17814 6232 17823 6252
rect 17779 6216 17823 6232
rect 17888 6248 17937 6258
rect 17888 6228 17899 6248
rect 17919 6228 17937 6248
rect 17888 6216 17937 6228
rect 17987 6252 18031 6258
rect 17987 6232 18002 6252
rect 18022 6232 18031 6252
rect 17987 6216 18031 6232
rect 18101 6252 18145 6258
rect 18101 6232 18110 6252
rect 18130 6232 18145 6252
rect 18101 6216 18145 6232
rect 18195 6248 18244 6258
rect 18195 6228 18213 6248
rect 18233 6228 18244 6248
rect 18195 6216 18244 6228
rect 13782 6081 13831 6093
rect 9130 6022 9179 6032
rect 5586 5954 5635 5964
rect 5586 5934 5597 5954
rect 5617 5934 5635 5954
rect 5586 5922 5635 5934
rect 5685 5958 5729 5964
rect 5685 5938 5700 5958
rect 5720 5938 5729 5958
rect 5685 5922 5729 5938
rect 5799 5954 5848 5964
rect 5799 5934 5810 5954
rect 5830 5934 5848 5954
rect 5799 5922 5848 5934
rect 5898 5958 5942 5964
rect 5898 5938 5913 5958
rect 5933 5938 5942 5958
rect 5898 5922 5942 5938
rect 6007 5954 6056 5964
rect 6007 5934 6018 5954
rect 6038 5934 6056 5954
rect 6007 5922 6056 5934
rect 6106 5958 6150 5964
rect 6106 5938 6121 5958
rect 6141 5938 6150 5958
rect 6106 5922 6150 5938
rect 6220 5958 6264 5964
rect 6220 5938 6229 5958
rect 6249 5938 6264 5958
rect 6220 5922 6264 5938
rect 6314 5954 6363 5964
rect 6314 5934 6332 5954
rect 6352 5934 6363 5954
rect 6314 5922 6363 5934
rect 4133 5892 4182 5904
rect 4133 5872 4144 5892
rect 4164 5872 4182 5892
rect 4133 5862 4182 5872
rect 4232 5888 4276 5904
rect 4232 5868 4247 5888
rect 4267 5868 4276 5888
rect 4232 5862 4276 5868
rect 4346 5888 4390 5904
rect 4346 5868 4355 5888
rect 4375 5868 4390 5888
rect 4346 5862 4390 5868
rect 4440 5892 4489 5904
rect 4440 5872 4458 5892
rect 4478 5872 4489 5892
rect 4440 5862 4489 5872
rect 4554 5888 4598 5904
rect 4554 5868 4563 5888
rect 4583 5868 4598 5888
rect 4554 5862 4598 5868
rect 4648 5892 4697 5904
rect 4648 5872 4666 5892
rect 4686 5872 4697 5892
rect 4648 5862 4697 5872
rect 4767 5888 4811 5904
rect 4767 5868 4776 5888
rect 4796 5868 4811 5888
rect 4767 5862 4811 5868
rect 4861 5892 4910 5904
rect 4861 5872 4879 5892
rect 4899 5872 4910 5892
rect 4861 5862 4910 5872
rect 1317 5794 1366 5804
rect 1317 5774 1328 5794
rect 1348 5774 1366 5794
rect 1317 5762 1366 5774
rect 1416 5798 1460 5804
rect 1416 5778 1431 5798
rect 1451 5778 1460 5798
rect 1416 5762 1460 5778
rect 1530 5794 1579 5804
rect 1530 5774 1541 5794
rect 1561 5774 1579 5794
rect 1530 5762 1579 5774
rect 1629 5798 1673 5804
rect 1629 5778 1644 5798
rect 1664 5778 1673 5798
rect 1629 5762 1673 5778
rect 1738 5794 1787 5804
rect 1738 5774 1749 5794
rect 1769 5774 1787 5794
rect 1738 5762 1787 5774
rect 1837 5798 1881 5804
rect 1837 5778 1852 5798
rect 1872 5778 1881 5798
rect 1837 5762 1881 5778
rect 1951 5798 1995 5804
rect 1951 5778 1960 5798
rect 1980 5778 1995 5798
rect 1951 5762 1995 5778
rect 2045 5794 2094 5804
rect 2045 5774 2063 5794
rect 2083 5774 2094 5794
rect 13782 6061 13793 6081
rect 13813 6061 13831 6081
rect 13782 6051 13831 6061
rect 13881 6077 13925 6093
rect 13881 6057 13896 6077
rect 13916 6057 13925 6077
rect 13881 6051 13925 6057
rect 13995 6077 14039 6093
rect 13995 6057 14004 6077
rect 14024 6057 14039 6077
rect 13995 6051 14039 6057
rect 14089 6081 14138 6093
rect 14089 6061 14107 6081
rect 14127 6061 14138 6081
rect 14089 6051 14138 6061
rect 14203 6077 14247 6093
rect 14203 6057 14212 6077
rect 14232 6057 14247 6077
rect 14203 6051 14247 6057
rect 14297 6081 14346 6093
rect 14297 6061 14315 6081
rect 14335 6061 14346 6081
rect 14297 6051 14346 6061
rect 14416 6077 14460 6093
rect 14416 6057 14425 6077
rect 14445 6057 14460 6077
rect 14416 6051 14460 6057
rect 14510 6081 14559 6093
rect 14510 6061 14528 6081
rect 14548 6061 14559 6081
rect 14510 6051 14559 6061
rect 10966 5983 11015 5993
rect 10966 5963 10977 5983
rect 10997 5963 11015 5983
rect 10966 5951 11015 5963
rect 11065 5987 11109 5993
rect 11065 5967 11080 5987
rect 11100 5967 11109 5987
rect 11065 5951 11109 5967
rect 11179 5983 11228 5993
rect 11179 5963 11190 5983
rect 11210 5963 11228 5983
rect 11179 5951 11228 5963
rect 11278 5987 11322 5993
rect 11278 5967 11293 5987
rect 11313 5967 11322 5987
rect 11278 5951 11322 5967
rect 11387 5983 11436 5993
rect 11387 5963 11398 5983
rect 11418 5963 11436 5983
rect 11387 5951 11436 5963
rect 11486 5987 11530 5993
rect 11486 5967 11501 5987
rect 11521 5967 11530 5987
rect 11486 5951 11530 5967
rect 11600 5987 11644 5993
rect 11600 5967 11609 5987
rect 11629 5967 11644 5987
rect 11600 5951 11644 5967
rect 11694 5983 11743 5993
rect 11694 5963 11712 5983
rect 11732 5963 11743 5983
rect 11694 5951 11743 5963
rect 2045 5762 2094 5774
rect 19063 6060 19112 6072
rect 9414 5871 9463 5883
rect 9414 5851 9425 5871
rect 9445 5851 9463 5871
rect 9414 5841 9463 5851
rect 9513 5867 9557 5883
rect 9513 5847 9528 5867
rect 9548 5847 9557 5867
rect 9513 5841 9557 5847
rect 9627 5867 9671 5883
rect 9627 5847 9636 5867
rect 9656 5847 9671 5867
rect 9627 5841 9671 5847
rect 9721 5871 9770 5883
rect 9721 5851 9739 5871
rect 9759 5851 9770 5871
rect 9721 5841 9770 5851
rect 9835 5867 9879 5883
rect 9835 5847 9844 5867
rect 9864 5847 9879 5867
rect 9835 5841 9879 5847
rect 9929 5871 9978 5883
rect 9929 5851 9947 5871
rect 9967 5851 9978 5871
rect 9929 5841 9978 5851
rect 10048 5867 10092 5883
rect 10048 5847 10057 5867
rect 10077 5847 10092 5867
rect 10048 5841 10092 5847
rect 10142 5871 10191 5883
rect 10142 5851 10160 5871
rect 10180 5851 10191 5871
rect 10142 5841 10191 5851
rect 6598 5773 6647 5783
rect 6598 5753 6609 5773
rect 6629 5753 6647 5773
rect 6598 5741 6647 5753
rect 6697 5777 6741 5783
rect 6697 5757 6712 5777
rect 6732 5757 6741 5777
rect 6697 5741 6741 5757
rect 6811 5773 6860 5783
rect 6811 5753 6822 5773
rect 6842 5753 6860 5773
rect 6811 5741 6860 5753
rect 6910 5777 6954 5783
rect 6910 5757 6925 5777
rect 6945 5757 6954 5777
rect 6910 5741 6954 5757
rect 7019 5773 7068 5783
rect 7019 5753 7030 5773
rect 7050 5753 7068 5773
rect 7019 5741 7068 5753
rect 7118 5777 7162 5783
rect 7118 5757 7133 5777
rect 7153 5757 7162 5777
rect 7118 5741 7162 5757
rect 7232 5777 7276 5783
rect 7232 5757 7241 5777
rect 7261 5757 7276 5777
rect 7232 5741 7276 5757
rect 7326 5773 7375 5783
rect 7326 5753 7344 5773
rect 7364 5753 7375 5773
rect 19063 6040 19074 6060
rect 19094 6040 19112 6060
rect 19063 6030 19112 6040
rect 19162 6056 19206 6072
rect 19162 6036 19177 6056
rect 19197 6036 19206 6056
rect 19162 6030 19206 6036
rect 19276 6056 19320 6072
rect 19276 6036 19285 6056
rect 19305 6036 19320 6056
rect 19276 6030 19320 6036
rect 19370 6060 19419 6072
rect 19370 6040 19388 6060
rect 19408 6040 19419 6060
rect 19370 6030 19419 6040
rect 19484 6056 19528 6072
rect 19484 6036 19493 6056
rect 19513 6036 19528 6056
rect 19484 6030 19528 6036
rect 19578 6060 19627 6072
rect 19578 6040 19596 6060
rect 19616 6040 19627 6060
rect 19578 6030 19627 6040
rect 19697 6056 19741 6072
rect 19697 6036 19706 6056
rect 19726 6036 19741 6056
rect 19697 6030 19741 6036
rect 19791 6060 19840 6072
rect 19791 6040 19809 6060
rect 19829 6040 19840 6060
rect 19791 6030 19840 6040
rect 16247 5962 16296 5972
rect 16247 5942 16258 5962
rect 16278 5942 16296 5962
rect 16247 5930 16296 5942
rect 16346 5966 16390 5972
rect 16346 5946 16361 5966
rect 16381 5946 16390 5966
rect 16346 5930 16390 5946
rect 16460 5962 16509 5972
rect 16460 5942 16471 5962
rect 16491 5942 16509 5962
rect 16460 5930 16509 5942
rect 16559 5966 16603 5972
rect 16559 5946 16574 5966
rect 16594 5946 16603 5966
rect 16559 5930 16603 5946
rect 16668 5962 16717 5972
rect 16668 5942 16679 5962
rect 16699 5942 16717 5962
rect 16668 5930 16717 5942
rect 16767 5966 16811 5972
rect 16767 5946 16782 5966
rect 16802 5946 16811 5966
rect 16767 5930 16811 5946
rect 16881 5966 16925 5972
rect 16881 5946 16890 5966
rect 16910 5946 16925 5966
rect 16881 5930 16925 5946
rect 16975 5962 17024 5972
rect 16975 5942 16993 5962
rect 17013 5942 17024 5962
rect 16975 5930 17024 5942
rect 14794 5900 14843 5912
rect 14794 5880 14805 5900
rect 14825 5880 14843 5900
rect 14794 5870 14843 5880
rect 14893 5896 14937 5912
rect 14893 5876 14908 5896
rect 14928 5876 14937 5896
rect 14893 5870 14937 5876
rect 15007 5896 15051 5912
rect 15007 5876 15016 5896
rect 15036 5876 15051 5896
rect 15007 5870 15051 5876
rect 15101 5900 15150 5912
rect 15101 5880 15119 5900
rect 15139 5880 15150 5900
rect 15101 5870 15150 5880
rect 15215 5896 15259 5912
rect 15215 5876 15224 5896
rect 15244 5876 15259 5896
rect 15215 5870 15259 5876
rect 15309 5900 15358 5912
rect 15309 5880 15327 5900
rect 15347 5880 15358 5900
rect 15309 5870 15358 5880
rect 15428 5896 15472 5912
rect 15428 5876 15437 5896
rect 15457 5876 15472 5896
rect 15428 5870 15472 5876
rect 15522 5900 15571 5912
rect 15522 5880 15540 5900
rect 15560 5880 15571 5900
rect 15522 5870 15571 5880
rect 11978 5802 12027 5812
rect 7326 5741 7375 5753
rect 3071 5653 3120 5665
rect 3071 5633 3082 5653
rect 3102 5633 3120 5653
rect 3071 5623 3120 5633
rect 3170 5649 3214 5665
rect 3170 5629 3185 5649
rect 3205 5629 3214 5649
rect 3170 5623 3214 5629
rect 3284 5649 3328 5665
rect 3284 5629 3293 5649
rect 3313 5629 3328 5649
rect 3284 5623 3328 5629
rect 3378 5653 3427 5665
rect 3378 5633 3396 5653
rect 3416 5633 3427 5653
rect 3378 5623 3427 5633
rect 3492 5649 3536 5665
rect 3492 5629 3501 5649
rect 3521 5629 3536 5649
rect 3492 5623 3536 5629
rect 3586 5653 3635 5665
rect 3586 5633 3604 5653
rect 3624 5633 3635 5653
rect 3586 5623 3635 5633
rect 3705 5649 3749 5665
rect 3705 5629 3714 5649
rect 3734 5629 3749 5649
rect 3705 5623 3749 5629
rect 3799 5653 3848 5665
rect 3799 5633 3817 5653
rect 3837 5633 3848 5653
rect 3799 5623 3848 5633
rect 304 5560 353 5570
rect 304 5540 315 5560
rect 335 5540 353 5560
rect 304 5528 353 5540
rect 403 5564 447 5570
rect 403 5544 418 5564
rect 438 5544 447 5564
rect 403 5528 447 5544
rect 517 5560 566 5570
rect 517 5540 528 5560
rect 548 5540 566 5560
rect 517 5528 566 5540
rect 616 5564 660 5570
rect 616 5544 631 5564
rect 651 5544 660 5564
rect 616 5528 660 5544
rect 725 5560 774 5570
rect 725 5540 736 5560
rect 756 5540 774 5560
rect 725 5528 774 5540
rect 824 5564 868 5570
rect 824 5544 839 5564
rect 859 5544 868 5564
rect 824 5528 868 5544
rect 938 5564 982 5570
rect 938 5544 947 5564
rect 967 5544 982 5564
rect 938 5528 982 5544
rect 1032 5560 1081 5570
rect 1032 5540 1050 5560
rect 1070 5540 1081 5560
rect 11978 5782 11989 5802
rect 12009 5782 12027 5802
rect 11978 5770 12027 5782
rect 12077 5806 12121 5812
rect 12077 5786 12092 5806
rect 12112 5786 12121 5806
rect 12077 5770 12121 5786
rect 12191 5802 12240 5812
rect 12191 5782 12202 5802
rect 12222 5782 12240 5802
rect 12191 5770 12240 5782
rect 12290 5806 12334 5812
rect 12290 5786 12305 5806
rect 12325 5786 12334 5806
rect 12290 5770 12334 5786
rect 12399 5802 12448 5812
rect 12399 5782 12410 5802
rect 12430 5782 12448 5802
rect 12399 5770 12448 5782
rect 12498 5806 12542 5812
rect 12498 5786 12513 5806
rect 12533 5786 12542 5806
rect 12498 5770 12542 5786
rect 12612 5806 12656 5812
rect 12612 5786 12621 5806
rect 12641 5786 12656 5806
rect 12612 5770 12656 5786
rect 12706 5802 12755 5812
rect 12706 5782 12724 5802
rect 12744 5782 12755 5802
rect 12706 5770 12755 5782
rect 20075 5879 20124 5891
rect 20075 5859 20086 5879
rect 20106 5859 20124 5879
rect 20075 5849 20124 5859
rect 20174 5875 20218 5891
rect 20174 5855 20189 5875
rect 20209 5855 20218 5875
rect 20174 5849 20218 5855
rect 20288 5875 20332 5891
rect 20288 5855 20297 5875
rect 20317 5855 20332 5875
rect 20288 5849 20332 5855
rect 20382 5879 20431 5891
rect 20382 5859 20400 5879
rect 20420 5859 20431 5879
rect 20382 5849 20431 5859
rect 20496 5875 20540 5891
rect 20496 5855 20505 5875
rect 20525 5855 20540 5875
rect 20496 5849 20540 5855
rect 20590 5879 20639 5891
rect 20590 5859 20608 5879
rect 20628 5859 20639 5879
rect 20590 5849 20639 5859
rect 20709 5875 20753 5891
rect 20709 5855 20718 5875
rect 20738 5855 20753 5875
rect 20709 5849 20753 5855
rect 20803 5879 20852 5891
rect 20803 5859 20821 5879
rect 20841 5859 20852 5879
rect 20803 5849 20852 5859
rect 17259 5781 17308 5791
rect 17259 5761 17270 5781
rect 17290 5761 17308 5781
rect 17259 5749 17308 5761
rect 17358 5785 17402 5791
rect 17358 5765 17373 5785
rect 17393 5765 17402 5785
rect 17358 5749 17402 5765
rect 17472 5781 17521 5791
rect 17472 5761 17483 5781
rect 17503 5761 17521 5781
rect 17472 5749 17521 5761
rect 17571 5785 17615 5791
rect 17571 5765 17586 5785
rect 17606 5765 17615 5785
rect 17571 5749 17615 5765
rect 17680 5781 17729 5791
rect 17680 5761 17691 5781
rect 17711 5761 17729 5781
rect 17680 5749 17729 5761
rect 17779 5785 17823 5791
rect 17779 5765 17794 5785
rect 17814 5765 17823 5785
rect 17779 5749 17823 5765
rect 17893 5785 17937 5791
rect 17893 5765 17902 5785
rect 17922 5765 17937 5785
rect 17893 5749 17937 5765
rect 17987 5781 18036 5791
rect 17987 5761 18005 5781
rect 18025 5761 18036 5781
rect 17987 5749 18036 5761
rect 13732 5661 13781 5673
rect 8352 5632 8401 5644
rect 1032 5528 1081 5540
rect 8352 5612 8363 5632
rect 8383 5612 8401 5632
rect 8352 5602 8401 5612
rect 8451 5628 8495 5644
rect 8451 5608 8466 5628
rect 8486 5608 8495 5628
rect 8451 5602 8495 5608
rect 8565 5628 8609 5644
rect 8565 5608 8574 5628
rect 8594 5608 8609 5628
rect 8565 5602 8609 5608
rect 8659 5632 8708 5644
rect 8659 5612 8677 5632
rect 8697 5612 8708 5632
rect 8659 5602 8708 5612
rect 8773 5628 8817 5644
rect 8773 5608 8782 5628
rect 8802 5608 8817 5628
rect 8773 5602 8817 5608
rect 8867 5632 8916 5644
rect 8867 5612 8885 5632
rect 8905 5612 8916 5632
rect 8867 5602 8916 5612
rect 8986 5628 9030 5644
rect 8986 5608 8995 5628
rect 9015 5608 9030 5628
rect 8986 5602 9030 5608
rect 9080 5632 9129 5644
rect 9080 5612 9098 5632
rect 9118 5612 9129 5632
rect 9080 5602 9129 5612
rect 5585 5539 5634 5549
rect 5585 5519 5596 5539
rect 5616 5519 5634 5539
rect 5585 5507 5634 5519
rect 5684 5543 5728 5549
rect 5684 5523 5699 5543
rect 5719 5523 5728 5543
rect 5684 5507 5728 5523
rect 5798 5539 5847 5549
rect 5798 5519 5809 5539
rect 5829 5519 5847 5539
rect 5798 5507 5847 5519
rect 5897 5543 5941 5549
rect 5897 5523 5912 5543
rect 5932 5523 5941 5543
rect 5897 5507 5941 5523
rect 6006 5539 6055 5549
rect 6006 5519 6017 5539
rect 6037 5519 6055 5539
rect 6006 5507 6055 5519
rect 6105 5543 6149 5549
rect 6105 5523 6120 5543
rect 6140 5523 6149 5543
rect 6105 5507 6149 5523
rect 6219 5543 6263 5549
rect 6219 5523 6228 5543
rect 6248 5523 6263 5543
rect 6219 5507 6263 5523
rect 6313 5539 6362 5549
rect 6313 5519 6331 5539
rect 6351 5519 6362 5539
rect 13732 5641 13743 5661
rect 13763 5641 13781 5661
rect 13732 5631 13781 5641
rect 13831 5657 13875 5673
rect 13831 5637 13846 5657
rect 13866 5637 13875 5657
rect 13831 5631 13875 5637
rect 13945 5657 13989 5673
rect 13945 5637 13954 5657
rect 13974 5637 13989 5657
rect 13945 5631 13989 5637
rect 14039 5661 14088 5673
rect 14039 5641 14057 5661
rect 14077 5641 14088 5661
rect 14039 5631 14088 5641
rect 14153 5657 14197 5673
rect 14153 5637 14162 5657
rect 14182 5637 14197 5657
rect 14153 5631 14197 5637
rect 14247 5661 14296 5673
rect 14247 5641 14265 5661
rect 14285 5641 14296 5661
rect 14247 5631 14296 5641
rect 14366 5657 14410 5673
rect 14366 5637 14375 5657
rect 14395 5637 14410 5657
rect 14366 5631 14410 5637
rect 14460 5661 14509 5673
rect 14460 5641 14478 5661
rect 14498 5641 14509 5661
rect 14460 5631 14509 5641
rect 6313 5507 6362 5519
rect 10965 5568 11014 5578
rect 10965 5548 10976 5568
rect 10996 5548 11014 5568
rect 10965 5536 11014 5548
rect 11064 5572 11108 5578
rect 11064 5552 11079 5572
rect 11099 5552 11108 5572
rect 11064 5536 11108 5552
rect 11178 5568 11227 5578
rect 11178 5548 11189 5568
rect 11209 5548 11227 5568
rect 11178 5536 11227 5548
rect 11277 5572 11321 5578
rect 11277 5552 11292 5572
rect 11312 5552 11321 5572
rect 11277 5536 11321 5552
rect 11386 5568 11435 5578
rect 11386 5548 11397 5568
rect 11417 5548 11435 5568
rect 11386 5536 11435 5548
rect 11485 5572 11529 5578
rect 11485 5552 11500 5572
rect 11520 5552 11529 5572
rect 11485 5536 11529 5552
rect 11599 5572 11643 5578
rect 11599 5552 11608 5572
rect 11628 5552 11643 5572
rect 11599 5536 11643 5552
rect 11693 5568 11742 5578
rect 11693 5548 11711 5568
rect 11731 5548 11742 5568
rect 19013 5640 19062 5652
rect 11693 5536 11742 5548
rect 19013 5620 19024 5640
rect 19044 5620 19062 5640
rect 19013 5610 19062 5620
rect 19112 5636 19156 5652
rect 19112 5616 19127 5636
rect 19147 5616 19156 5636
rect 19112 5610 19156 5616
rect 19226 5636 19270 5652
rect 19226 5616 19235 5636
rect 19255 5616 19270 5636
rect 19226 5610 19270 5616
rect 19320 5640 19369 5652
rect 19320 5620 19338 5640
rect 19358 5620 19369 5640
rect 19320 5610 19369 5620
rect 19434 5636 19478 5652
rect 19434 5616 19443 5636
rect 19463 5616 19478 5636
rect 19434 5610 19478 5616
rect 19528 5640 19577 5652
rect 19528 5620 19546 5640
rect 19566 5620 19577 5640
rect 19528 5610 19577 5620
rect 19647 5636 19691 5652
rect 19647 5616 19656 5636
rect 19676 5616 19691 5636
rect 19647 5610 19691 5616
rect 19741 5640 19790 5652
rect 19741 5620 19759 5640
rect 19779 5620 19790 5640
rect 19741 5610 19790 5620
rect 16246 5547 16295 5557
rect 16246 5527 16257 5547
rect 16277 5527 16295 5547
rect 16246 5515 16295 5527
rect 16345 5551 16389 5557
rect 16345 5531 16360 5551
rect 16380 5531 16389 5551
rect 16345 5515 16389 5531
rect 16459 5547 16508 5557
rect 16459 5527 16470 5547
rect 16490 5527 16508 5547
rect 16459 5515 16508 5527
rect 16558 5551 16602 5557
rect 16558 5531 16573 5551
rect 16593 5531 16602 5551
rect 16558 5515 16602 5531
rect 16667 5547 16716 5557
rect 16667 5527 16678 5547
rect 16698 5527 16716 5547
rect 16667 5515 16716 5527
rect 16766 5551 16810 5557
rect 16766 5531 16781 5551
rect 16801 5531 16810 5551
rect 16766 5515 16810 5531
rect 16880 5551 16924 5557
rect 16880 5531 16889 5551
rect 16909 5531 16924 5551
rect 16880 5515 16924 5531
rect 16974 5547 17023 5557
rect 16974 5527 16992 5547
rect 17012 5527 17023 5547
rect 16974 5515 17023 5527
rect 4139 5326 4188 5338
rect 4139 5306 4150 5326
rect 4170 5306 4188 5326
rect 4139 5296 4188 5306
rect 4238 5322 4282 5338
rect 4238 5302 4253 5322
rect 4273 5302 4282 5322
rect 4238 5296 4282 5302
rect 4352 5322 4396 5338
rect 4352 5302 4361 5322
rect 4381 5302 4396 5322
rect 4352 5296 4396 5302
rect 4446 5326 4495 5338
rect 4446 5306 4464 5326
rect 4484 5306 4495 5326
rect 4446 5296 4495 5306
rect 4560 5322 4604 5338
rect 4560 5302 4569 5322
rect 4589 5302 4604 5322
rect 4560 5296 4604 5302
rect 4654 5326 4703 5338
rect 4654 5306 4672 5326
rect 4692 5306 4703 5326
rect 4654 5296 4703 5306
rect 4773 5322 4817 5338
rect 4773 5302 4782 5322
rect 4802 5302 4817 5322
rect 4773 5296 4817 5302
rect 4867 5326 4916 5338
rect 4867 5306 4885 5326
rect 4905 5306 4916 5326
rect 4867 5296 4916 5306
rect 1372 5233 1421 5243
rect 1372 5213 1383 5233
rect 1403 5213 1421 5233
rect 1372 5201 1421 5213
rect 1471 5237 1515 5243
rect 1471 5217 1486 5237
rect 1506 5217 1515 5237
rect 1471 5201 1515 5217
rect 1585 5233 1634 5243
rect 1585 5213 1596 5233
rect 1616 5213 1634 5233
rect 1585 5201 1634 5213
rect 1684 5237 1728 5243
rect 1684 5217 1699 5237
rect 1719 5217 1728 5237
rect 1684 5201 1728 5217
rect 1793 5233 1842 5243
rect 1793 5213 1804 5233
rect 1824 5213 1842 5233
rect 1793 5201 1842 5213
rect 1892 5237 1936 5243
rect 1892 5217 1907 5237
rect 1927 5217 1936 5237
rect 1892 5201 1936 5217
rect 2006 5237 2050 5243
rect 2006 5217 2015 5237
rect 2035 5217 2050 5237
rect 2006 5201 2050 5217
rect 2100 5233 2149 5243
rect 2100 5213 2118 5233
rect 2138 5213 2149 5233
rect 9420 5305 9469 5317
rect 2100 5201 2149 5213
rect 9420 5285 9431 5305
rect 9451 5285 9469 5305
rect 9420 5275 9469 5285
rect 9519 5301 9563 5317
rect 9519 5281 9534 5301
rect 9554 5281 9563 5301
rect 9519 5275 9563 5281
rect 9633 5301 9677 5317
rect 9633 5281 9642 5301
rect 9662 5281 9677 5301
rect 9633 5275 9677 5281
rect 9727 5305 9776 5317
rect 9727 5285 9745 5305
rect 9765 5285 9776 5305
rect 9727 5275 9776 5285
rect 9841 5301 9885 5317
rect 9841 5281 9850 5301
rect 9870 5281 9885 5301
rect 9841 5275 9885 5281
rect 9935 5305 9984 5317
rect 9935 5285 9953 5305
rect 9973 5285 9984 5305
rect 9935 5275 9984 5285
rect 10054 5301 10098 5317
rect 10054 5281 10063 5301
rect 10083 5281 10098 5301
rect 10054 5275 10098 5281
rect 10148 5305 10197 5317
rect 10148 5285 10166 5305
rect 10186 5285 10197 5305
rect 10148 5275 10197 5285
rect 14800 5334 14849 5346
rect 6653 5212 6702 5222
rect 6653 5192 6664 5212
rect 6684 5192 6702 5212
rect 6653 5180 6702 5192
rect 6752 5216 6796 5222
rect 6752 5196 6767 5216
rect 6787 5196 6796 5216
rect 6752 5180 6796 5196
rect 6866 5212 6915 5222
rect 6866 5192 6877 5212
rect 6897 5192 6915 5212
rect 6866 5180 6915 5192
rect 6965 5216 7009 5222
rect 6965 5196 6980 5216
rect 7000 5196 7009 5216
rect 6965 5180 7009 5196
rect 7074 5212 7123 5222
rect 7074 5192 7085 5212
rect 7105 5192 7123 5212
rect 7074 5180 7123 5192
rect 7173 5216 7217 5222
rect 7173 5196 7188 5216
rect 7208 5196 7217 5216
rect 7173 5180 7217 5196
rect 7287 5216 7331 5222
rect 7287 5196 7296 5216
rect 7316 5196 7331 5216
rect 7287 5180 7331 5196
rect 7381 5212 7430 5222
rect 7381 5192 7399 5212
rect 7419 5192 7430 5212
rect 14800 5314 14811 5334
rect 14831 5314 14849 5334
rect 14800 5304 14849 5314
rect 14899 5330 14943 5346
rect 14899 5310 14914 5330
rect 14934 5310 14943 5330
rect 14899 5304 14943 5310
rect 15013 5330 15057 5346
rect 15013 5310 15022 5330
rect 15042 5310 15057 5330
rect 15013 5304 15057 5310
rect 15107 5334 15156 5346
rect 15107 5314 15125 5334
rect 15145 5314 15156 5334
rect 15107 5304 15156 5314
rect 15221 5330 15265 5346
rect 15221 5310 15230 5330
rect 15250 5310 15265 5330
rect 15221 5304 15265 5310
rect 15315 5334 15364 5346
rect 15315 5314 15333 5334
rect 15353 5314 15364 5334
rect 15315 5304 15364 5314
rect 15434 5330 15478 5346
rect 15434 5310 15443 5330
rect 15463 5310 15478 5330
rect 15434 5304 15478 5310
rect 15528 5334 15577 5346
rect 15528 5314 15546 5334
rect 15566 5314 15577 5334
rect 15528 5304 15577 5314
rect 12033 5241 12082 5251
rect 12033 5221 12044 5241
rect 12064 5221 12082 5241
rect 12033 5209 12082 5221
rect 12132 5245 12176 5251
rect 12132 5225 12147 5245
rect 12167 5225 12176 5245
rect 12132 5209 12176 5225
rect 12246 5241 12295 5251
rect 12246 5221 12257 5241
rect 12277 5221 12295 5241
rect 12246 5209 12295 5221
rect 12345 5245 12389 5251
rect 12345 5225 12360 5245
rect 12380 5225 12389 5245
rect 12345 5209 12389 5225
rect 12454 5241 12503 5251
rect 12454 5221 12465 5241
rect 12485 5221 12503 5241
rect 12454 5209 12503 5221
rect 12553 5245 12597 5251
rect 12553 5225 12568 5245
rect 12588 5225 12597 5245
rect 12553 5209 12597 5225
rect 12667 5245 12711 5251
rect 12667 5225 12676 5245
rect 12696 5225 12711 5245
rect 12667 5209 12711 5225
rect 12761 5241 12810 5251
rect 12761 5221 12779 5241
rect 12799 5221 12810 5241
rect 20081 5313 20130 5325
rect 12761 5209 12810 5221
rect 7381 5180 7430 5192
rect 3126 5092 3175 5104
rect 3126 5072 3137 5092
rect 3157 5072 3175 5092
rect 3126 5062 3175 5072
rect 3225 5088 3269 5104
rect 3225 5068 3240 5088
rect 3260 5068 3269 5088
rect 3225 5062 3269 5068
rect 3339 5088 3383 5104
rect 3339 5068 3348 5088
rect 3368 5068 3383 5088
rect 3339 5062 3383 5068
rect 3433 5092 3482 5104
rect 3433 5072 3451 5092
rect 3471 5072 3482 5092
rect 3433 5062 3482 5072
rect 3547 5088 3591 5104
rect 3547 5068 3556 5088
rect 3576 5068 3591 5088
rect 3547 5062 3591 5068
rect 3641 5092 3690 5104
rect 3641 5072 3659 5092
rect 3679 5072 3690 5092
rect 3641 5062 3690 5072
rect 3760 5088 3804 5104
rect 3760 5068 3769 5088
rect 3789 5068 3804 5088
rect 3760 5062 3804 5068
rect 3854 5092 3903 5104
rect 3854 5072 3872 5092
rect 3892 5072 3903 5092
rect 3854 5062 3903 5072
rect 310 4994 359 5004
rect 310 4974 321 4994
rect 341 4974 359 4994
rect 310 4962 359 4974
rect 409 4998 453 5004
rect 409 4978 424 4998
rect 444 4978 453 4998
rect 409 4962 453 4978
rect 523 4994 572 5004
rect 523 4974 534 4994
rect 554 4974 572 4994
rect 523 4962 572 4974
rect 622 4998 666 5004
rect 622 4978 637 4998
rect 657 4978 666 4998
rect 622 4962 666 4978
rect 731 4994 780 5004
rect 731 4974 742 4994
rect 762 4974 780 4994
rect 731 4962 780 4974
rect 830 4998 874 5004
rect 830 4978 845 4998
rect 865 4978 874 4998
rect 830 4962 874 4978
rect 944 4998 988 5004
rect 944 4978 953 4998
rect 973 4978 988 4998
rect 944 4962 988 4978
rect 1038 4994 1087 5004
rect 1038 4974 1056 4994
rect 1076 4974 1087 4994
rect 1038 4962 1087 4974
rect 8407 5071 8456 5083
rect 8407 5051 8418 5071
rect 8438 5051 8456 5071
rect 8407 5041 8456 5051
rect 8506 5067 8550 5083
rect 8506 5047 8521 5067
rect 8541 5047 8550 5067
rect 8506 5041 8550 5047
rect 8620 5067 8664 5083
rect 8620 5047 8629 5067
rect 8649 5047 8664 5067
rect 8620 5041 8664 5047
rect 8714 5071 8763 5083
rect 8714 5051 8732 5071
rect 8752 5051 8763 5071
rect 8714 5041 8763 5051
rect 8828 5067 8872 5083
rect 8828 5047 8837 5067
rect 8857 5047 8872 5067
rect 8828 5041 8872 5047
rect 8922 5071 8971 5083
rect 8922 5051 8940 5071
rect 8960 5051 8971 5071
rect 8922 5041 8971 5051
rect 9041 5067 9085 5083
rect 9041 5047 9050 5067
rect 9070 5047 9085 5067
rect 9041 5041 9085 5047
rect 9135 5071 9184 5083
rect 9135 5051 9153 5071
rect 9173 5051 9184 5071
rect 20081 5293 20092 5313
rect 20112 5293 20130 5313
rect 20081 5283 20130 5293
rect 20180 5309 20224 5325
rect 20180 5289 20195 5309
rect 20215 5289 20224 5309
rect 20180 5283 20224 5289
rect 20294 5309 20338 5325
rect 20294 5289 20303 5309
rect 20323 5289 20338 5309
rect 20294 5283 20338 5289
rect 20388 5313 20437 5325
rect 20388 5293 20406 5313
rect 20426 5293 20437 5313
rect 20388 5283 20437 5293
rect 20502 5309 20546 5325
rect 20502 5289 20511 5309
rect 20531 5289 20546 5309
rect 20502 5283 20546 5289
rect 20596 5313 20645 5325
rect 20596 5293 20614 5313
rect 20634 5293 20645 5313
rect 20596 5283 20645 5293
rect 20715 5309 20759 5325
rect 20715 5289 20724 5309
rect 20744 5289 20759 5309
rect 20715 5283 20759 5289
rect 20809 5313 20858 5325
rect 20809 5293 20827 5313
rect 20847 5293 20858 5313
rect 20809 5283 20858 5293
rect 17314 5220 17363 5230
rect 17314 5200 17325 5220
rect 17345 5200 17363 5220
rect 17314 5188 17363 5200
rect 17413 5224 17457 5230
rect 17413 5204 17428 5224
rect 17448 5204 17457 5224
rect 17413 5188 17457 5204
rect 17527 5220 17576 5230
rect 17527 5200 17538 5220
rect 17558 5200 17576 5220
rect 17527 5188 17576 5200
rect 17626 5224 17670 5230
rect 17626 5204 17641 5224
rect 17661 5204 17670 5224
rect 17626 5188 17670 5204
rect 17735 5220 17784 5230
rect 17735 5200 17746 5220
rect 17766 5200 17784 5220
rect 17735 5188 17784 5200
rect 17834 5224 17878 5230
rect 17834 5204 17849 5224
rect 17869 5204 17878 5224
rect 17834 5188 17878 5204
rect 17948 5224 17992 5230
rect 17948 5204 17957 5224
rect 17977 5204 17992 5224
rect 17948 5188 17992 5204
rect 18042 5220 18091 5230
rect 18042 5200 18060 5220
rect 18080 5200 18091 5220
rect 18042 5188 18091 5200
rect 13787 5100 13836 5112
rect 9135 5041 9184 5051
rect 5591 4973 5640 4983
rect 5591 4953 5602 4973
rect 5622 4953 5640 4973
rect 5591 4941 5640 4953
rect 5690 4977 5734 4983
rect 5690 4957 5705 4977
rect 5725 4957 5734 4977
rect 5690 4941 5734 4957
rect 5804 4973 5853 4983
rect 5804 4953 5815 4973
rect 5835 4953 5853 4973
rect 5804 4941 5853 4953
rect 5903 4977 5947 4983
rect 5903 4957 5918 4977
rect 5938 4957 5947 4977
rect 5903 4941 5947 4957
rect 6012 4973 6061 4983
rect 6012 4953 6023 4973
rect 6043 4953 6061 4973
rect 6012 4941 6061 4953
rect 6111 4977 6155 4983
rect 6111 4957 6126 4977
rect 6146 4957 6155 4977
rect 6111 4941 6155 4957
rect 6225 4977 6269 4983
rect 6225 4957 6234 4977
rect 6254 4957 6269 4977
rect 6225 4941 6269 4957
rect 6319 4973 6368 4983
rect 6319 4953 6337 4973
rect 6357 4953 6368 4973
rect 6319 4941 6368 4953
rect 4138 4911 4187 4923
rect 4138 4891 4149 4911
rect 4169 4891 4187 4911
rect 4138 4881 4187 4891
rect 4237 4907 4281 4923
rect 4237 4887 4252 4907
rect 4272 4887 4281 4907
rect 4237 4881 4281 4887
rect 4351 4907 4395 4923
rect 4351 4887 4360 4907
rect 4380 4887 4395 4907
rect 4351 4881 4395 4887
rect 4445 4911 4494 4923
rect 4445 4891 4463 4911
rect 4483 4891 4494 4911
rect 4445 4881 4494 4891
rect 4559 4907 4603 4923
rect 4559 4887 4568 4907
rect 4588 4887 4603 4907
rect 4559 4881 4603 4887
rect 4653 4911 4702 4923
rect 4653 4891 4671 4911
rect 4691 4891 4702 4911
rect 4653 4881 4702 4891
rect 4772 4907 4816 4923
rect 4772 4887 4781 4907
rect 4801 4887 4816 4907
rect 4772 4881 4816 4887
rect 4866 4911 4915 4923
rect 4866 4891 4884 4911
rect 4904 4891 4915 4911
rect 4866 4881 4915 4891
rect 1322 4813 1371 4823
rect 1322 4793 1333 4813
rect 1353 4793 1371 4813
rect 1322 4781 1371 4793
rect 1421 4817 1465 4823
rect 1421 4797 1436 4817
rect 1456 4797 1465 4817
rect 1421 4781 1465 4797
rect 1535 4813 1584 4823
rect 1535 4793 1546 4813
rect 1566 4793 1584 4813
rect 1535 4781 1584 4793
rect 1634 4817 1678 4823
rect 1634 4797 1649 4817
rect 1669 4797 1678 4817
rect 1634 4781 1678 4797
rect 1743 4813 1792 4823
rect 1743 4793 1754 4813
rect 1774 4793 1792 4813
rect 1743 4781 1792 4793
rect 1842 4817 1886 4823
rect 1842 4797 1857 4817
rect 1877 4797 1886 4817
rect 1842 4781 1886 4797
rect 1956 4817 2000 4823
rect 1956 4797 1965 4817
rect 1985 4797 2000 4817
rect 1956 4781 2000 4797
rect 2050 4813 2099 4823
rect 2050 4793 2068 4813
rect 2088 4793 2099 4813
rect 13787 5080 13798 5100
rect 13818 5080 13836 5100
rect 13787 5070 13836 5080
rect 13886 5096 13930 5112
rect 13886 5076 13901 5096
rect 13921 5076 13930 5096
rect 13886 5070 13930 5076
rect 14000 5096 14044 5112
rect 14000 5076 14009 5096
rect 14029 5076 14044 5096
rect 14000 5070 14044 5076
rect 14094 5100 14143 5112
rect 14094 5080 14112 5100
rect 14132 5080 14143 5100
rect 14094 5070 14143 5080
rect 14208 5096 14252 5112
rect 14208 5076 14217 5096
rect 14237 5076 14252 5096
rect 14208 5070 14252 5076
rect 14302 5100 14351 5112
rect 14302 5080 14320 5100
rect 14340 5080 14351 5100
rect 14302 5070 14351 5080
rect 14421 5096 14465 5112
rect 14421 5076 14430 5096
rect 14450 5076 14465 5096
rect 14421 5070 14465 5076
rect 14515 5100 14564 5112
rect 14515 5080 14533 5100
rect 14553 5080 14564 5100
rect 14515 5070 14564 5080
rect 10971 5002 11020 5012
rect 10971 4982 10982 5002
rect 11002 4982 11020 5002
rect 10971 4970 11020 4982
rect 11070 5006 11114 5012
rect 11070 4986 11085 5006
rect 11105 4986 11114 5006
rect 11070 4970 11114 4986
rect 11184 5002 11233 5012
rect 11184 4982 11195 5002
rect 11215 4982 11233 5002
rect 11184 4970 11233 4982
rect 11283 5006 11327 5012
rect 11283 4986 11298 5006
rect 11318 4986 11327 5006
rect 11283 4970 11327 4986
rect 11392 5002 11441 5012
rect 11392 4982 11403 5002
rect 11423 4982 11441 5002
rect 11392 4970 11441 4982
rect 11491 5006 11535 5012
rect 11491 4986 11506 5006
rect 11526 4986 11535 5006
rect 11491 4970 11535 4986
rect 11605 5006 11649 5012
rect 11605 4986 11614 5006
rect 11634 4986 11649 5006
rect 11605 4970 11649 4986
rect 11699 5002 11748 5012
rect 11699 4982 11717 5002
rect 11737 4982 11748 5002
rect 11699 4970 11748 4982
rect 2050 4781 2099 4793
rect 19068 5079 19117 5091
rect 9419 4890 9468 4902
rect 9419 4870 9430 4890
rect 9450 4870 9468 4890
rect 9419 4860 9468 4870
rect 9518 4886 9562 4902
rect 9518 4866 9533 4886
rect 9553 4866 9562 4886
rect 9518 4860 9562 4866
rect 9632 4886 9676 4902
rect 9632 4866 9641 4886
rect 9661 4866 9676 4886
rect 9632 4860 9676 4866
rect 9726 4890 9775 4902
rect 9726 4870 9744 4890
rect 9764 4870 9775 4890
rect 9726 4860 9775 4870
rect 9840 4886 9884 4902
rect 9840 4866 9849 4886
rect 9869 4866 9884 4886
rect 9840 4860 9884 4866
rect 9934 4890 9983 4902
rect 9934 4870 9952 4890
rect 9972 4870 9983 4890
rect 9934 4860 9983 4870
rect 10053 4886 10097 4902
rect 10053 4866 10062 4886
rect 10082 4866 10097 4886
rect 10053 4860 10097 4866
rect 10147 4890 10196 4902
rect 10147 4870 10165 4890
rect 10185 4870 10196 4890
rect 10147 4860 10196 4870
rect 6603 4792 6652 4802
rect 6603 4772 6614 4792
rect 6634 4772 6652 4792
rect 6603 4760 6652 4772
rect 6702 4796 6746 4802
rect 6702 4776 6717 4796
rect 6737 4776 6746 4796
rect 6702 4760 6746 4776
rect 6816 4792 6865 4802
rect 6816 4772 6827 4792
rect 6847 4772 6865 4792
rect 6816 4760 6865 4772
rect 6915 4796 6959 4802
rect 6915 4776 6930 4796
rect 6950 4776 6959 4796
rect 6915 4760 6959 4776
rect 7024 4792 7073 4802
rect 7024 4772 7035 4792
rect 7055 4772 7073 4792
rect 7024 4760 7073 4772
rect 7123 4796 7167 4802
rect 7123 4776 7138 4796
rect 7158 4776 7167 4796
rect 7123 4760 7167 4776
rect 7237 4796 7281 4802
rect 7237 4776 7246 4796
rect 7266 4776 7281 4796
rect 7237 4760 7281 4776
rect 7331 4792 7380 4802
rect 7331 4772 7349 4792
rect 7369 4772 7380 4792
rect 19068 5059 19079 5079
rect 19099 5059 19117 5079
rect 19068 5049 19117 5059
rect 19167 5075 19211 5091
rect 19167 5055 19182 5075
rect 19202 5055 19211 5075
rect 19167 5049 19211 5055
rect 19281 5075 19325 5091
rect 19281 5055 19290 5075
rect 19310 5055 19325 5075
rect 19281 5049 19325 5055
rect 19375 5079 19424 5091
rect 19375 5059 19393 5079
rect 19413 5059 19424 5079
rect 19375 5049 19424 5059
rect 19489 5075 19533 5091
rect 19489 5055 19498 5075
rect 19518 5055 19533 5075
rect 19489 5049 19533 5055
rect 19583 5079 19632 5091
rect 19583 5059 19601 5079
rect 19621 5059 19632 5079
rect 19583 5049 19632 5059
rect 19702 5075 19746 5091
rect 19702 5055 19711 5075
rect 19731 5055 19746 5075
rect 19702 5049 19746 5055
rect 19796 5079 19845 5091
rect 19796 5059 19814 5079
rect 19834 5059 19845 5079
rect 19796 5049 19845 5059
rect 16252 4981 16301 4991
rect 16252 4961 16263 4981
rect 16283 4961 16301 4981
rect 16252 4949 16301 4961
rect 16351 4985 16395 4991
rect 16351 4965 16366 4985
rect 16386 4965 16395 4985
rect 16351 4949 16395 4965
rect 16465 4981 16514 4991
rect 16465 4961 16476 4981
rect 16496 4961 16514 4981
rect 16465 4949 16514 4961
rect 16564 4985 16608 4991
rect 16564 4965 16579 4985
rect 16599 4965 16608 4985
rect 16564 4949 16608 4965
rect 16673 4981 16722 4991
rect 16673 4961 16684 4981
rect 16704 4961 16722 4981
rect 16673 4949 16722 4961
rect 16772 4985 16816 4991
rect 16772 4965 16787 4985
rect 16807 4965 16816 4985
rect 16772 4949 16816 4965
rect 16886 4985 16930 4991
rect 16886 4965 16895 4985
rect 16915 4965 16930 4985
rect 16886 4949 16930 4965
rect 16980 4981 17029 4991
rect 16980 4961 16998 4981
rect 17018 4961 17029 4981
rect 16980 4949 17029 4961
rect 14799 4919 14848 4931
rect 14799 4899 14810 4919
rect 14830 4899 14848 4919
rect 14799 4889 14848 4899
rect 14898 4915 14942 4931
rect 14898 4895 14913 4915
rect 14933 4895 14942 4915
rect 14898 4889 14942 4895
rect 15012 4915 15056 4931
rect 15012 4895 15021 4915
rect 15041 4895 15056 4915
rect 15012 4889 15056 4895
rect 15106 4919 15155 4931
rect 15106 4899 15124 4919
rect 15144 4899 15155 4919
rect 15106 4889 15155 4899
rect 15220 4915 15264 4931
rect 15220 4895 15229 4915
rect 15249 4895 15264 4915
rect 15220 4889 15264 4895
rect 15314 4919 15363 4931
rect 15314 4899 15332 4919
rect 15352 4899 15363 4919
rect 15314 4889 15363 4899
rect 15433 4915 15477 4931
rect 15433 4895 15442 4915
rect 15462 4895 15477 4915
rect 15433 4889 15477 4895
rect 15527 4919 15576 4931
rect 15527 4899 15545 4919
rect 15565 4899 15576 4919
rect 15527 4889 15576 4899
rect 11983 4821 12032 4831
rect 7331 4760 7380 4772
rect 2831 4660 2880 4672
rect 2831 4640 2842 4660
rect 2862 4640 2880 4660
rect 2831 4630 2880 4640
rect 2930 4656 2974 4672
rect 2930 4636 2945 4656
rect 2965 4636 2974 4656
rect 2930 4630 2974 4636
rect 3044 4656 3088 4672
rect 3044 4636 3053 4656
rect 3073 4636 3088 4656
rect 3044 4630 3088 4636
rect 3138 4660 3187 4672
rect 3138 4640 3156 4660
rect 3176 4640 3187 4660
rect 3138 4630 3187 4640
rect 3252 4656 3296 4672
rect 3252 4636 3261 4656
rect 3281 4636 3296 4656
rect 3252 4630 3296 4636
rect 3346 4660 3395 4672
rect 3346 4640 3364 4660
rect 3384 4640 3395 4660
rect 3346 4630 3395 4640
rect 3465 4656 3509 4672
rect 3465 4636 3474 4656
rect 3494 4636 3509 4656
rect 3465 4630 3509 4636
rect 3559 4660 3608 4672
rect 3559 4640 3577 4660
rect 3597 4640 3608 4660
rect 3559 4630 3608 4640
rect 11983 4801 11994 4821
rect 12014 4801 12032 4821
rect 11983 4789 12032 4801
rect 12082 4825 12126 4831
rect 12082 4805 12097 4825
rect 12117 4805 12126 4825
rect 12082 4789 12126 4805
rect 12196 4821 12245 4831
rect 12196 4801 12207 4821
rect 12227 4801 12245 4821
rect 12196 4789 12245 4801
rect 12295 4825 12339 4831
rect 12295 4805 12310 4825
rect 12330 4805 12339 4825
rect 12295 4789 12339 4805
rect 12404 4821 12453 4831
rect 12404 4801 12415 4821
rect 12435 4801 12453 4821
rect 12404 4789 12453 4801
rect 12503 4825 12547 4831
rect 12503 4805 12518 4825
rect 12538 4805 12547 4825
rect 12503 4789 12547 4805
rect 12617 4825 12661 4831
rect 12617 4805 12626 4825
rect 12646 4805 12661 4825
rect 12617 4789 12661 4805
rect 12711 4821 12760 4831
rect 12711 4801 12729 4821
rect 12749 4801 12760 4821
rect 12711 4789 12760 4801
rect 20080 4898 20129 4910
rect 20080 4878 20091 4898
rect 20111 4878 20129 4898
rect 20080 4868 20129 4878
rect 20179 4894 20223 4910
rect 20179 4874 20194 4894
rect 20214 4874 20223 4894
rect 20179 4868 20223 4874
rect 20293 4894 20337 4910
rect 20293 4874 20302 4894
rect 20322 4874 20337 4894
rect 20293 4868 20337 4874
rect 20387 4898 20436 4910
rect 20387 4878 20405 4898
rect 20425 4878 20436 4898
rect 20387 4868 20436 4878
rect 20501 4894 20545 4910
rect 20501 4874 20510 4894
rect 20530 4874 20545 4894
rect 20501 4868 20545 4874
rect 20595 4898 20644 4910
rect 20595 4878 20613 4898
rect 20633 4878 20644 4898
rect 20595 4868 20644 4878
rect 20714 4894 20758 4910
rect 20714 4874 20723 4894
rect 20743 4874 20758 4894
rect 20714 4868 20758 4874
rect 20808 4898 20857 4910
rect 20808 4878 20826 4898
rect 20846 4878 20857 4898
rect 20808 4868 20857 4878
rect 17264 4800 17313 4810
rect 17264 4780 17275 4800
rect 17295 4780 17313 4800
rect 17264 4768 17313 4780
rect 17363 4804 17407 4810
rect 17363 4784 17378 4804
rect 17398 4784 17407 4804
rect 17363 4768 17407 4784
rect 17477 4800 17526 4810
rect 17477 4780 17488 4800
rect 17508 4780 17526 4800
rect 17477 4768 17526 4780
rect 17576 4804 17620 4810
rect 17576 4784 17591 4804
rect 17611 4784 17620 4804
rect 17576 4768 17620 4784
rect 17685 4800 17734 4810
rect 17685 4780 17696 4800
rect 17716 4780 17734 4800
rect 17685 4768 17734 4780
rect 17784 4804 17828 4810
rect 17784 4784 17799 4804
rect 17819 4784 17828 4804
rect 17784 4768 17828 4784
rect 17898 4804 17942 4810
rect 17898 4784 17907 4804
rect 17927 4784 17942 4804
rect 17898 4768 17942 4784
rect 17992 4800 18041 4810
rect 17992 4780 18010 4800
rect 18030 4780 18041 4800
rect 17992 4768 18041 4780
rect 309 4579 358 4589
rect 309 4559 320 4579
rect 340 4559 358 4579
rect 309 4547 358 4559
rect 408 4583 452 4589
rect 408 4563 423 4583
rect 443 4563 452 4583
rect 408 4547 452 4563
rect 522 4579 571 4589
rect 522 4559 533 4579
rect 553 4559 571 4579
rect 522 4547 571 4559
rect 621 4583 665 4589
rect 621 4563 636 4583
rect 656 4563 665 4583
rect 621 4547 665 4563
rect 730 4579 779 4589
rect 730 4559 741 4579
rect 761 4559 779 4579
rect 730 4547 779 4559
rect 829 4583 873 4589
rect 829 4563 844 4583
rect 864 4563 873 4583
rect 829 4547 873 4563
rect 943 4583 987 4589
rect 943 4563 952 4583
rect 972 4563 987 4583
rect 943 4547 987 4563
rect 1037 4579 1086 4589
rect 1037 4559 1055 4579
rect 1075 4559 1086 4579
rect 1037 4547 1086 4559
rect 8112 4639 8161 4651
rect 8112 4619 8123 4639
rect 8143 4619 8161 4639
rect 8112 4609 8161 4619
rect 8211 4635 8255 4651
rect 8211 4615 8226 4635
rect 8246 4615 8255 4635
rect 8211 4609 8255 4615
rect 8325 4635 8369 4651
rect 8325 4615 8334 4635
rect 8354 4615 8369 4635
rect 8325 4609 8369 4615
rect 8419 4639 8468 4651
rect 8419 4619 8437 4639
rect 8457 4619 8468 4639
rect 8419 4609 8468 4619
rect 8533 4635 8577 4651
rect 8533 4615 8542 4635
rect 8562 4615 8577 4635
rect 8533 4609 8577 4615
rect 8627 4639 8676 4651
rect 8627 4619 8645 4639
rect 8665 4619 8676 4639
rect 8627 4609 8676 4619
rect 8746 4635 8790 4651
rect 8746 4615 8755 4635
rect 8775 4615 8790 4635
rect 8746 4609 8790 4615
rect 8840 4639 8889 4651
rect 8840 4619 8858 4639
rect 8878 4619 8889 4639
rect 8840 4609 8889 4619
rect 5590 4558 5639 4568
rect 5590 4538 5601 4558
rect 5621 4538 5639 4558
rect 5590 4526 5639 4538
rect 5689 4562 5733 4568
rect 5689 4542 5704 4562
rect 5724 4542 5733 4562
rect 5689 4526 5733 4542
rect 5803 4558 5852 4568
rect 5803 4538 5814 4558
rect 5834 4538 5852 4558
rect 5803 4526 5852 4538
rect 5902 4562 5946 4568
rect 5902 4542 5917 4562
rect 5937 4542 5946 4562
rect 5902 4526 5946 4542
rect 6011 4558 6060 4568
rect 6011 4538 6022 4558
rect 6042 4538 6060 4558
rect 6011 4526 6060 4538
rect 6110 4562 6154 4568
rect 6110 4542 6125 4562
rect 6145 4542 6154 4562
rect 6110 4526 6154 4542
rect 6224 4562 6268 4568
rect 6224 4542 6233 4562
rect 6253 4542 6268 4562
rect 6224 4526 6268 4542
rect 6318 4558 6367 4568
rect 6318 4538 6336 4558
rect 6356 4538 6367 4558
rect 6318 4526 6367 4538
rect 13492 4668 13541 4680
rect 13492 4648 13503 4668
rect 13523 4648 13541 4668
rect 13492 4638 13541 4648
rect 13591 4664 13635 4680
rect 13591 4644 13606 4664
rect 13626 4644 13635 4664
rect 13591 4638 13635 4644
rect 13705 4664 13749 4680
rect 13705 4644 13714 4664
rect 13734 4644 13749 4664
rect 13705 4638 13749 4644
rect 13799 4668 13848 4680
rect 13799 4648 13817 4668
rect 13837 4648 13848 4668
rect 13799 4638 13848 4648
rect 13913 4664 13957 4680
rect 13913 4644 13922 4664
rect 13942 4644 13957 4664
rect 13913 4638 13957 4644
rect 14007 4668 14056 4680
rect 14007 4648 14025 4668
rect 14045 4648 14056 4668
rect 14007 4638 14056 4648
rect 14126 4664 14170 4680
rect 14126 4644 14135 4664
rect 14155 4644 14170 4664
rect 14126 4638 14170 4644
rect 14220 4668 14269 4680
rect 14220 4648 14238 4668
rect 14258 4648 14269 4668
rect 14220 4638 14269 4648
rect 4142 4350 4191 4362
rect 4142 4330 4153 4350
rect 4173 4330 4191 4350
rect 4142 4320 4191 4330
rect 4241 4346 4285 4362
rect 4241 4326 4256 4346
rect 4276 4326 4285 4346
rect 4241 4320 4285 4326
rect 4355 4346 4399 4362
rect 4355 4326 4364 4346
rect 4384 4326 4399 4346
rect 4355 4320 4399 4326
rect 4449 4350 4498 4362
rect 4449 4330 4467 4350
rect 4487 4330 4498 4350
rect 4449 4320 4498 4330
rect 4563 4346 4607 4362
rect 4563 4326 4572 4346
rect 4592 4326 4607 4346
rect 4563 4320 4607 4326
rect 4657 4350 4706 4362
rect 4657 4330 4675 4350
rect 4695 4330 4706 4350
rect 4657 4320 4706 4330
rect 4776 4346 4820 4362
rect 4776 4326 4785 4346
rect 4805 4326 4820 4346
rect 4776 4320 4820 4326
rect 4870 4350 4919 4362
rect 4870 4330 4888 4350
rect 4908 4330 4919 4350
rect 4870 4320 4919 4330
rect 1620 4269 1669 4279
rect 1620 4249 1631 4269
rect 1651 4249 1669 4269
rect 1620 4237 1669 4249
rect 1719 4273 1763 4279
rect 1719 4253 1734 4273
rect 1754 4253 1763 4273
rect 1719 4237 1763 4253
rect 1833 4269 1882 4279
rect 1833 4249 1844 4269
rect 1864 4249 1882 4269
rect 1833 4237 1882 4249
rect 1932 4273 1976 4279
rect 1932 4253 1947 4273
rect 1967 4253 1976 4273
rect 1932 4237 1976 4253
rect 2041 4269 2090 4279
rect 2041 4249 2052 4269
rect 2072 4249 2090 4269
rect 2041 4237 2090 4249
rect 2140 4273 2184 4279
rect 2140 4253 2155 4273
rect 2175 4253 2184 4273
rect 2140 4237 2184 4253
rect 2254 4273 2298 4279
rect 2254 4253 2263 4273
rect 2283 4253 2298 4273
rect 2254 4237 2298 4253
rect 2348 4269 2397 4279
rect 2348 4249 2366 4269
rect 2386 4249 2397 4269
rect 2348 4237 2397 4249
rect 10970 4587 11019 4597
rect 10970 4567 10981 4587
rect 11001 4567 11019 4587
rect 10970 4555 11019 4567
rect 11069 4591 11113 4597
rect 11069 4571 11084 4591
rect 11104 4571 11113 4591
rect 11069 4555 11113 4571
rect 11183 4587 11232 4597
rect 11183 4567 11194 4587
rect 11214 4567 11232 4587
rect 11183 4555 11232 4567
rect 11282 4591 11326 4597
rect 11282 4571 11297 4591
rect 11317 4571 11326 4591
rect 11282 4555 11326 4571
rect 11391 4587 11440 4597
rect 11391 4567 11402 4587
rect 11422 4567 11440 4587
rect 11391 4555 11440 4567
rect 11490 4591 11534 4597
rect 11490 4571 11505 4591
rect 11525 4571 11534 4591
rect 11490 4555 11534 4571
rect 11604 4591 11648 4597
rect 11604 4571 11613 4591
rect 11633 4571 11648 4591
rect 11604 4555 11648 4571
rect 11698 4587 11747 4597
rect 11698 4567 11716 4587
rect 11736 4567 11747 4587
rect 11698 4555 11747 4567
rect 9423 4329 9472 4341
rect 9423 4309 9434 4329
rect 9454 4309 9472 4329
rect 9423 4299 9472 4309
rect 9522 4325 9566 4341
rect 9522 4305 9537 4325
rect 9557 4305 9566 4325
rect 9522 4299 9566 4305
rect 9636 4325 9680 4341
rect 9636 4305 9645 4325
rect 9665 4305 9680 4325
rect 9636 4299 9680 4305
rect 9730 4329 9779 4341
rect 9730 4309 9748 4329
rect 9768 4309 9779 4329
rect 9730 4299 9779 4309
rect 9844 4325 9888 4341
rect 9844 4305 9853 4325
rect 9873 4305 9888 4325
rect 9844 4299 9888 4305
rect 9938 4329 9987 4341
rect 9938 4309 9956 4329
rect 9976 4309 9987 4329
rect 9938 4299 9987 4309
rect 10057 4325 10101 4341
rect 10057 4305 10066 4325
rect 10086 4305 10101 4325
rect 10057 4299 10101 4305
rect 10151 4329 10200 4341
rect 10151 4309 10169 4329
rect 10189 4309 10200 4329
rect 10151 4299 10200 4309
rect 18773 4647 18822 4659
rect 18773 4627 18784 4647
rect 18804 4627 18822 4647
rect 18773 4617 18822 4627
rect 18872 4643 18916 4659
rect 18872 4623 18887 4643
rect 18907 4623 18916 4643
rect 18872 4617 18916 4623
rect 18986 4643 19030 4659
rect 18986 4623 18995 4643
rect 19015 4623 19030 4643
rect 18986 4617 19030 4623
rect 19080 4647 19129 4659
rect 19080 4627 19098 4647
rect 19118 4627 19129 4647
rect 19080 4617 19129 4627
rect 19194 4643 19238 4659
rect 19194 4623 19203 4643
rect 19223 4623 19238 4643
rect 19194 4617 19238 4623
rect 19288 4647 19337 4659
rect 19288 4627 19306 4647
rect 19326 4627 19337 4647
rect 19288 4617 19337 4627
rect 19407 4643 19451 4659
rect 19407 4623 19416 4643
rect 19436 4623 19451 4643
rect 19407 4617 19451 4623
rect 19501 4647 19550 4659
rect 19501 4627 19519 4647
rect 19539 4627 19550 4647
rect 19501 4617 19550 4627
rect 16251 4566 16300 4576
rect 16251 4546 16262 4566
rect 16282 4546 16300 4566
rect 16251 4534 16300 4546
rect 16350 4570 16394 4576
rect 16350 4550 16365 4570
rect 16385 4550 16394 4570
rect 16350 4534 16394 4550
rect 16464 4566 16513 4576
rect 16464 4546 16475 4566
rect 16495 4546 16513 4566
rect 16464 4534 16513 4546
rect 16563 4570 16607 4576
rect 16563 4550 16578 4570
rect 16598 4550 16607 4570
rect 16563 4534 16607 4550
rect 16672 4566 16721 4576
rect 16672 4546 16683 4566
rect 16703 4546 16721 4566
rect 16672 4534 16721 4546
rect 16771 4570 16815 4576
rect 16771 4550 16786 4570
rect 16806 4550 16815 4570
rect 16771 4534 16815 4550
rect 16885 4570 16929 4576
rect 16885 4550 16894 4570
rect 16914 4550 16929 4570
rect 16885 4534 16929 4550
rect 16979 4566 17028 4576
rect 16979 4546 16997 4566
rect 17017 4546 17028 4566
rect 16979 4534 17028 4546
rect 6901 4248 6950 4258
rect 6901 4228 6912 4248
rect 6932 4228 6950 4248
rect 6901 4216 6950 4228
rect 7000 4252 7044 4258
rect 7000 4232 7015 4252
rect 7035 4232 7044 4252
rect 7000 4216 7044 4232
rect 7114 4248 7163 4258
rect 7114 4228 7125 4248
rect 7145 4228 7163 4248
rect 7114 4216 7163 4228
rect 7213 4252 7257 4258
rect 7213 4232 7228 4252
rect 7248 4232 7257 4252
rect 7213 4216 7257 4232
rect 7322 4248 7371 4258
rect 7322 4228 7333 4248
rect 7353 4228 7371 4248
rect 7322 4216 7371 4228
rect 7421 4252 7465 4258
rect 7421 4232 7436 4252
rect 7456 4232 7465 4252
rect 7421 4216 7465 4232
rect 7535 4252 7579 4258
rect 7535 4232 7544 4252
rect 7564 4232 7579 4252
rect 7535 4216 7579 4232
rect 7629 4248 7678 4258
rect 7629 4228 7647 4248
rect 7667 4228 7678 4248
rect 7629 4216 7678 4228
rect 14803 4358 14852 4370
rect 14803 4338 14814 4358
rect 14834 4338 14852 4358
rect 14803 4328 14852 4338
rect 14902 4354 14946 4370
rect 14902 4334 14917 4354
rect 14937 4334 14946 4354
rect 14902 4328 14946 4334
rect 15016 4354 15060 4370
rect 15016 4334 15025 4354
rect 15045 4334 15060 4354
rect 15016 4328 15060 4334
rect 15110 4358 15159 4370
rect 15110 4338 15128 4358
rect 15148 4338 15159 4358
rect 15110 4328 15159 4338
rect 15224 4354 15268 4370
rect 15224 4334 15233 4354
rect 15253 4334 15268 4354
rect 15224 4328 15268 4334
rect 15318 4358 15367 4370
rect 15318 4338 15336 4358
rect 15356 4338 15367 4358
rect 15318 4328 15367 4338
rect 15437 4354 15481 4370
rect 15437 4334 15446 4354
rect 15466 4334 15481 4354
rect 15437 4328 15481 4334
rect 15531 4358 15580 4370
rect 15531 4338 15549 4358
rect 15569 4338 15580 4358
rect 15531 4328 15580 4338
rect 12281 4277 12330 4287
rect 12281 4257 12292 4277
rect 12312 4257 12330 4277
rect 12281 4245 12330 4257
rect 12380 4281 12424 4287
rect 12380 4261 12395 4281
rect 12415 4261 12424 4281
rect 12380 4245 12424 4261
rect 12494 4277 12543 4287
rect 12494 4257 12505 4277
rect 12525 4257 12543 4277
rect 12494 4245 12543 4257
rect 12593 4281 12637 4287
rect 12593 4261 12608 4281
rect 12628 4261 12637 4281
rect 12593 4245 12637 4261
rect 12702 4277 12751 4287
rect 12702 4257 12713 4277
rect 12733 4257 12751 4277
rect 12702 4245 12751 4257
rect 12801 4281 12845 4287
rect 12801 4261 12816 4281
rect 12836 4261 12845 4281
rect 12801 4245 12845 4261
rect 12915 4281 12959 4287
rect 12915 4261 12924 4281
rect 12944 4261 12959 4281
rect 12915 4245 12959 4261
rect 13009 4277 13058 4287
rect 13009 4257 13027 4277
rect 13047 4257 13058 4277
rect 13009 4245 13058 4257
rect 20084 4337 20133 4349
rect 20084 4317 20095 4337
rect 20115 4317 20133 4337
rect 20084 4307 20133 4317
rect 20183 4333 20227 4349
rect 20183 4313 20198 4333
rect 20218 4313 20227 4333
rect 20183 4307 20227 4313
rect 20297 4333 20341 4349
rect 20297 4313 20306 4333
rect 20326 4313 20341 4333
rect 20297 4307 20341 4313
rect 20391 4337 20440 4349
rect 20391 4317 20409 4337
rect 20429 4317 20440 4337
rect 20391 4307 20440 4317
rect 20505 4333 20549 4349
rect 20505 4313 20514 4333
rect 20534 4313 20549 4333
rect 20505 4307 20549 4313
rect 20599 4337 20648 4349
rect 20599 4317 20617 4337
rect 20637 4317 20648 4337
rect 20599 4307 20648 4317
rect 20718 4333 20762 4349
rect 20718 4313 20727 4333
rect 20747 4313 20762 4333
rect 20718 4307 20762 4313
rect 20812 4337 20861 4349
rect 20812 4317 20830 4337
rect 20850 4317 20861 4337
rect 20812 4307 20861 4317
rect 3129 4116 3178 4128
rect 3129 4096 3140 4116
rect 3160 4096 3178 4116
rect 3129 4086 3178 4096
rect 3228 4112 3272 4128
rect 3228 4092 3243 4112
rect 3263 4092 3272 4112
rect 3228 4086 3272 4092
rect 3342 4112 3386 4128
rect 3342 4092 3351 4112
rect 3371 4092 3386 4112
rect 3342 4086 3386 4092
rect 3436 4116 3485 4128
rect 3436 4096 3454 4116
rect 3474 4096 3485 4116
rect 3436 4086 3485 4096
rect 3550 4112 3594 4128
rect 3550 4092 3559 4112
rect 3579 4092 3594 4112
rect 3550 4086 3594 4092
rect 3644 4116 3693 4128
rect 3644 4096 3662 4116
rect 3682 4096 3693 4116
rect 3644 4086 3693 4096
rect 3763 4112 3807 4128
rect 3763 4092 3772 4112
rect 3792 4092 3807 4112
rect 3763 4086 3807 4092
rect 3857 4116 3906 4128
rect 3857 4096 3875 4116
rect 3895 4096 3906 4116
rect 3857 4086 3906 4096
rect 313 4018 362 4028
rect 313 3998 324 4018
rect 344 3998 362 4018
rect 313 3986 362 3998
rect 412 4022 456 4028
rect 412 4002 427 4022
rect 447 4002 456 4022
rect 412 3986 456 4002
rect 526 4018 575 4028
rect 526 3998 537 4018
rect 557 3998 575 4018
rect 526 3986 575 3998
rect 625 4022 669 4028
rect 625 4002 640 4022
rect 660 4002 669 4022
rect 625 3986 669 4002
rect 734 4018 783 4028
rect 734 3998 745 4018
rect 765 3998 783 4018
rect 734 3986 783 3998
rect 833 4022 877 4028
rect 833 4002 848 4022
rect 868 4002 877 4022
rect 833 3986 877 4002
rect 947 4022 991 4028
rect 947 4002 956 4022
rect 976 4002 991 4022
rect 947 3986 991 4002
rect 1041 4018 1090 4028
rect 1041 3998 1059 4018
rect 1079 3998 1090 4018
rect 1041 3986 1090 3998
rect 8410 4095 8459 4107
rect 8410 4075 8421 4095
rect 8441 4075 8459 4095
rect 8410 4065 8459 4075
rect 8509 4091 8553 4107
rect 8509 4071 8524 4091
rect 8544 4071 8553 4091
rect 8509 4065 8553 4071
rect 8623 4091 8667 4107
rect 8623 4071 8632 4091
rect 8652 4071 8667 4091
rect 8623 4065 8667 4071
rect 8717 4095 8766 4107
rect 8717 4075 8735 4095
rect 8755 4075 8766 4095
rect 8717 4065 8766 4075
rect 8831 4091 8875 4107
rect 8831 4071 8840 4091
rect 8860 4071 8875 4091
rect 8831 4065 8875 4071
rect 8925 4095 8974 4107
rect 8925 4075 8943 4095
rect 8963 4075 8974 4095
rect 8925 4065 8974 4075
rect 9044 4091 9088 4107
rect 9044 4071 9053 4091
rect 9073 4071 9088 4091
rect 9044 4065 9088 4071
rect 9138 4095 9187 4107
rect 9138 4075 9156 4095
rect 9176 4075 9187 4095
rect 17562 4256 17611 4266
rect 17562 4236 17573 4256
rect 17593 4236 17611 4256
rect 17562 4224 17611 4236
rect 17661 4260 17705 4266
rect 17661 4240 17676 4260
rect 17696 4240 17705 4260
rect 17661 4224 17705 4240
rect 17775 4256 17824 4266
rect 17775 4236 17786 4256
rect 17806 4236 17824 4256
rect 17775 4224 17824 4236
rect 17874 4260 17918 4266
rect 17874 4240 17889 4260
rect 17909 4240 17918 4260
rect 17874 4224 17918 4240
rect 17983 4256 18032 4266
rect 17983 4236 17994 4256
rect 18014 4236 18032 4256
rect 17983 4224 18032 4236
rect 18082 4260 18126 4266
rect 18082 4240 18097 4260
rect 18117 4240 18126 4260
rect 18082 4224 18126 4240
rect 18196 4260 18240 4266
rect 18196 4240 18205 4260
rect 18225 4240 18240 4260
rect 18196 4224 18240 4240
rect 18290 4256 18339 4266
rect 18290 4236 18308 4256
rect 18328 4236 18339 4256
rect 18290 4224 18339 4236
rect 13790 4124 13839 4136
rect 9138 4065 9187 4075
rect 5594 3997 5643 4007
rect 5594 3977 5605 3997
rect 5625 3977 5643 3997
rect 5594 3965 5643 3977
rect 5693 4001 5737 4007
rect 5693 3981 5708 4001
rect 5728 3981 5737 4001
rect 5693 3965 5737 3981
rect 5807 3997 5856 4007
rect 5807 3977 5818 3997
rect 5838 3977 5856 3997
rect 5807 3965 5856 3977
rect 5906 4001 5950 4007
rect 5906 3981 5921 4001
rect 5941 3981 5950 4001
rect 5906 3965 5950 3981
rect 6015 3997 6064 4007
rect 6015 3977 6026 3997
rect 6046 3977 6064 3997
rect 6015 3965 6064 3977
rect 6114 4001 6158 4007
rect 6114 3981 6129 4001
rect 6149 3981 6158 4001
rect 6114 3965 6158 3981
rect 6228 4001 6272 4007
rect 6228 3981 6237 4001
rect 6257 3981 6272 4001
rect 6228 3965 6272 3981
rect 6322 3997 6371 4007
rect 6322 3977 6340 3997
rect 6360 3977 6371 3997
rect 6322 3965 6371 3977
rect 4141 3935 4190 3947
rect 4141 3915 4152 3935
rect 4172 3915 4190 3935
rect 4141 3905 4190 3915
rect 4240 3931 4284 3947
rect 4240 3911 4255 3931
rect 4275 3911 4284 3931
rect 4240 3905 4284 3911
rect 4354 3931 4398 3947
rect 4354 3911 4363 3931
rect 4383 3911 4398 3931
rect 4354 3905 4398 3911
rect 4448 3935 4497 3947
rect 4448 3915 4466 3935
rect 4486 3915 4497 3935
rect 4448 3905 4497 3915
rect 4562 3931 4606 3947
rect 4562 3911 4571 3931
rect 4591 3911 4606 3931
rect 4562 3905 4606 3911
rect 4656 3935 4705 3947
rect 4656 3915 4674 3935
rect 4694 3915 4705 3935
rect 4656 3905 4705 3915
rect 4775 3931 4819 3947
rect 4775 3911 4784 3931
rect 4804 3911 4819 3931
rect 4775 3905 4819 3911
rect 4869 3935 4918 3947
rect 4869 3915 4887 3935
rect 4907 3915 4918 3935
rect 4869 3905 4918 3915
rect 1325 3837 1374 3847
rect 1325 3817 1336 3837
rect 1356 3817 1374 3837
rect 1325 3805 1374 3817
rect 1424 3841 1468 3847
rect 1424 3821 1439 3841
rect 1459 3821 1468 3841
rect 1424 3805 1468 3821
rect 1538 3837 1587 3847
rect 1538 3817 1549 3837
rect 1569 3817 1587 3837
rect 1538 3805 1587 3817
rect 1637 3841 1681 3847
rect 1637 3821 1652 3841
rect 1672 3821 1681 3841
rect 1637 3805 1681 3821
rect 1746 3837 1795 3847
rect 1746 3817 1757 3837
rect 1777 3817 1795 3837
rect 1746 3805 1795 3817
rect 1845 3841 1889 3847
rect 1845 3821 1860 3841
rect 1880 3821 1889 3841
rect 1845 3805 1889 3821
rect 1959 3841 2003 3847
rect 1959 3821 1968 3841
rect 1988 3821 2003 3841
rect 1959 3805 2003 3821
rect 2053 3837 2102 3847
rect 2053 3817 2071 3837
rect 2091 3817 2102 3837
rect 13790 4104 13801 4124
rect 13821 4104 13839 4124
rect 13790 4094 13839 4104
rect 13889 4120 13933 4136
rect 13889 4100 13904 4120
rect 13924 4100 13933 4120
rect 13889 4094 13933 4100
rect 14003 4120 14047 4136
rect 14003 4100 14012 4120
rect 14032 4100 14047 4120
rect 14003 4094 14047 4100
rect 14097 4124 14146 4136
rect 14097 4104 14115 4124
rect 14135 4104 14146 4124
rect 14097 4094 14146 4104
rect 14211 4120 14255 4136
rect 14211 4100 14220 4120
rect 14240 4100 14255 4120
rect 14211 4094 14255 4100
rect 14305 4124 14354 4136
rect 14305 4104 14323 4124
rect 14343 4104 14354 4124
rect 14305 4094 14354 4104
rect 14424 4120 14468 4136
rect 14424 4100 14433 4120
rect 14453 4100 14468 4120
rect 14424 4094 14468 4100
rect 14518 4124 14567 4136
rect 14518 4104 14536 4124
rect 14556 4104 14567 4124
rect 14518 4094 14567 4104
rect 10974 4026 11023 4036
rect 10974 4006 10985 4026
rect 11005 4006 11023 4026
rect 10974 3994 11023 4006
rect 11073 4030 11117 4036
rect 11073 4010 11088 4030
rect 11108 4010 11117 4030
rect 11073 3994 11117 4010
rect 11187 4026 11236 4036
rect 11187 4006 11198 4026
rect 11218 4006 11236 4026
rect 11187 3994 11236 4006
rect 11286 4030 11330 4036
rect 11286 4010 11301 4030
rect 11321 4010 11330 4030
rect 11286 3994 11330 4010
rect 11395 4026 11444 4036
rect 11395 4006 11406 4026
rect 11426 4006 11444 4026
rect 11395 3994 11444 4006
rect 11494 4030 11538 4036
rect 11494 4010 11509 4030
rect 11529 4010 11538 4030
rect 11494 3994 11538 4010
rect 11608 4030 11652 4036
rect 11608 4010 11617 4030
rect 11637 4010 11652 4030
rect 11608 3994 11652 4010
rect 11702 4026 11751 4036
rect 11702 4006 11720 4026
rect 11740 4006 11751 4026
rect 11702 3994 11751 4006
rect 2053 3805 2102 3817
rect 19071 4103 19120 4115
rect 9422 3914 9471 3926
rect 9422 3894 9433 3914
rect 9453 3894 9471 3914
rect 9422 3884 9471 3894
rect 9521 3910 9565 3926
rect 9521 3890 9536 3910
rect 9556 3890 9565 3910
rect 9521 3884 9565 3890
rect 9635 3910 9679 3926
rect 9635 3890 9644 3910
rect 9664 3890 9679 3910
rect 9635 3884 9679 3890
rect 9729 3914 9778 3926
rect 9729 3894 9747 3914
rect 9767 3894 9778 3914
rect 9729 3884 9778 3894
rect 9843 3910 9887 3926
rect 9843 3890 9852 3910
rect 9872 3890 9887 3910
rect 9843 3884 9887 3890
rect 9937 3914 9986 3926
rect 9937 3894 9955 3914
rect 9975 3894 9986 3914
rect 9937 3884 9986 3894
rect 10056 3910 10100 3926
rect 10056 3890 10065 3910
rect 10085 3890 10100 3910
rect 10056 3884 10100 3890
rect 10150 3914 10199 3926
rect 10150 3894 10168 3914
rect 10188 3894 10199 3914
rect 10150 3884 10199 3894
rect 6606 3816 6655 3826
rect 6606 3796 6617 3816
rect 6637 3796 6655 3816
rect 6606 3784 6655 3796
rect 6705 3820 6749 3826
rect 6705 3800 6720 3820
rect 6740 3800 6749 3820
rect 6705 3784 6749 3800
rect 6819 3816 6868 3826
rect 6819 3796 6830 3816
rect 6850 3796 6868 3816
rect 6819 3784 6868 3796
rect 6918 3820 6962 3826
rect 6918 3800 6933 3820
rect 6953 3800 6962 3820
rect 6918 3784 6962 3800
rect 7027 3816 7076 3826
rect 7027 3796 7038 3816
rect 7058 3796 7076 3816
rect 7027 3784 7076 3796
rect 7126 3820 7170 3826
rect 7126 3800 7141 3820
rect 7161 3800 7170 3820
rect 7126 3784 7170 3800
rect 7240 3820 7284 3826
rect 7240 3800 7249 3820
rect 7269 3800 7284 3820
rect 7240 3784 7284 3800
rect 7334 3816 7383 3826
rect 7334 3796 7352 3816
rect 7372 3796 7383 3816
rect 19071 4083 19082 4103
rect 19102 4083 19120 4103
rect 19071 4073 19120 4083
rect 19170 4099 19214 4115
rect 19170 4079 19185 4099
rect 19205 4079 19214 4099
rect 19170 4073 19214 4079
rect 19284 4099 19328 4115
rect 19284 4079 19293 4099
rect 19313 4079 19328 4099
rect 19284 4073 19328 4079
rect 19378 4103 19427 4115
rect 19378 4083 19396 4103
rect 19416 4083 19427 4103
rect 19378 4073 19427 4083
rect 19492 4099 19536 4115
rect 19492 4079 19501 4099
rect 19521 4079 19536 4099
rect 19492 4073 19536 4079
rect 19586 4103 19635 4115
rect 19586 4083 19604 4103
rect 19624 4083 19635 4103
rect 19586 4073 19635 4083
rect 19705 4099 19749 4115
rect 19705 4079 19714 4099
rect 19734 4079 19749 4099
rect 19705 4073 19749 4079
rect 19799 4103 19848 4115
rect 19799 4083 19817 4103
rect 19837 4083 19848 4103
rect 19799 4073 19848 4083
rect 16255 4005 16304 4015
rect 16255 3985 16266 4005
rect 16286 3985 16304 4005
rect 16255 3973 16304 3985
rect 16354 4009 16398 4015
rect 16354 3989 16369 4009
rect 16389 3989 16398 4009
rect 16354 3973 16398 3989
rect 16468 4005 16517 4015
rect 16468 3985 16479 4005
rect 16499 3985 16517 4005
rect 16468 3973 16517 3985
rect 16567 4009 16611 4015
rect 16567 3989 16582 4009
rect 16602 3989 16611 4009
rect 16567 3973 16611 3989
rect 16676 4005 16725 4015
rect 16676 3985 16687 4005
rect 16707 3985 16725 4005
rect 16676 3973 16725 3985
rect 16775 4009 16819 4015
rect 16775 3989 16790 4009
rect 16810 3989 16819 4009
rect 16775 3973 16819 3989
rect 16889 4009 16933 4015
rect 16889 3989 16898 4009
rect 16918 3989 16933 4009
rect 16889 3973 16933 3989
rect 16983 4005 17032 4015
rect 16983 3985 17001 4005
rect 17021 3985 17032 4005
rect 16983 3973 17032 3985
rect 14802 3943 14851 3955
rect 14802 3923 14813 3943
rect 14833 3923 14851 3943
rect 14802 3913 14851 3923
rect 14901 3939 14945 3955
rect 14901 3919 14916 3939
rect 14936 3919 14945 3939
rect 14901 3913 14945 3919
rect 15015 3939 15059 3955
rect 15015 3919 15024 3939
rect 15044 3919 15059 3939
rect 15015 3913 15059 3919
rect 15109 3943 15158 3955
rect 15109 3923 15127 3943
rect 15147 3923 15158 3943
rect 15109 3913 15158 3923
rect 15223 3939 15267 3955
rect 15223 3919 15232 3939
rect 15252 3919 15267 3939
rect 15223 3913 15267 3919
rect 15317 3943 15366 3955
rect 15317 3923 15335 3943
rect 15355 3923 15366 3943
rect 15317 3913 15366 3923
rect 15436 3939 15480 3955
rect 15436 3919 15445 3939
rect 15465 3919 15480 3939
rect 15436 3913 15480 3919
rect 15530 3943 15579 3955
rect 15530 3923 15548 3943
rect 15568 3923 15579 3943
rect 15530 3913 15579 3923
rect 11986 3845 12035 3855
rect 7334 3784 7383 3796
rect 3079 3696 3128 3708
rect 3079 3676 3090 3696
rect 3110 3676 3128 3696
rect 3079 3666 3128 3676
rect 3178 3692 3222 3708
rect 3178 3672 3193 3692
rect 3213 3672 3222 3692
rect 3178 3666 3222 3672
rect 3292 3692 3336 3708
rect 3292 3672 3301 3692
rect 3321 3672 3336 3692
rect 3292 3666 3336 3672
rect 3386 3696 3435 3708
rect 3386 3676 3404 3696
rect 3424 3676 3435 3696
rect 3386 3666 3435 3676
rect 3500 3692 3544 3708
rect 3500 3672 3509 3692
rect 3529 3672 3544 3692
rect 3500 3666 3544 3672
rect 3594 3696 3643 3708
rect 3594 3676 3612 3696
rect 3632 3676 3643 3696
rect 3594 3666 3643 3676
rect 3713 3692 3757 3708
rect 3713 3672 3722 3692
rect 3742 3672 3757 3692
rect 3713 3666 3757 3672
rect 3807 3696 3856 3708
rect 3807 3676 3825 3696
rect 3845 3676 3856 3696
rect 3807 3666 3856 3676
rect 312 3603 361 3613
rect 312 3583 323 3603
rect 343 3583 361 3603
rect 312 3571 361 3583
rect 411 3607 455 3613
rect 411 3587 426 3607
rect 446 3587 455 3607
rect 411 3571 455 3587
rect 525 3603 574 3613
rect 525 3583 536 3603
rect 556 3583 574 3603
rect 525 3571 574 3583
rect 624 3607 668 3613
rect 624 3587 639 3607
rect 659 3587 668 3607
rect 624 3571 668 3587
rect 733 3603 782 3613
rect 733 3583 744 3603
rect 764 3583 782 3603
rect 733 3571 782 3583
rect 832 3607 876 3613
rect 832 3587 847 3607
rect 867 3587 876 3607
rect 832 3571 876 3587
rect 946 3607 990 3613
rect 946 3587 955 3607
rect 975 3587 990 3607
rect 946 3571 990 3587
rect 1040 3603 1089 3613
rect 1040 3583 1058 3603
rect 1078 3583 1089 3603
rect 11986 3825 11997 3845
rect 12017 3825 12035 3845
rect 11986 3813 12035 3825
rect 12085 3849 12129 3855
rect 12085 3829 12100 3849
rect 12120 3829 12129 3849
rect 12085 3813 12129 3829
rect 12199 3845 12248 3855
rect 12199 3825 12210 3845
rect 12230 3825 12248 3845
rect 12199 3813 12248 3825
rect 12298 3849 12342 3855
rect 12298 3829 12313 3849
rect 12333 3829 12342 3849
rect 12298 3813 12342 3829
rect 12407 3845 12456 3855
rect 12407 3825 12418 3845
rect 12438 3825 12456 3845
rect 12407 3813 12456 3825
rect 12506 3849 12550 3855
rect 12506 3829 12521 3849
rect 12541 3829 12550 3849
rect 12506 3813 12550 3829
rect 12620 3849 12664 3855
rect 12620 3829 12629 3849
rect 12649 3829 12664 3849
rect 12620 3813 12664 3829
rect 12714 3845 12763 3855
rect 12714 3825 12732 3845
rect 12752 3825 12763 3845
rect 12714 3813 12763 3825
rect 20083 3922 20132 3934
rect 20083 3902 20094 3922
rect 20114 3902 20132 3922
rect 20083 3892 20132 3902
rect 20182 3918 20226 3934
rect 20182 3898 20197 3918
rect 20217 3898 20226 3918
rect 20182 3892 20226 3898
rect 20296 3918 20340 3934
rect 20296 3898 20305 3918
rect 20325 3898 20340 3918
rect 20296 3892 20340 3898
rect 20390 3922 20439 3934
rect 20390 3902 20408 3922
rect 20428 3902 20439 3922
rect 20390 3892 20439 3902
rect 20504 3918 20548 3934
rect 20504 3898 20513 3918
rect 20533 3898 20548 3918
rect 20504 3892 20548 3898
rect 20598 3922 20647 3934
rect 20598 3902 20616 3922
rect 20636 3902 20647 3922
rect 20598 3892 20647 3902
rect 20717 3918 20761 3934
rect 20717 3898 20726 3918
rect 20746 3898 20761 3918
rect 20717 3892 20761 3898
rect 20811 3922 20860 3934
rect 20811 3902 20829 3922
rect 20849 3902 20860 3922
rect 20811 3892 20860 3902
rect 17267 3824 17316 3834
rect 17267 3804 17278 3824
rect 17298 3804 17316 3824
rect 17267 3792 17316 3804
rect 17366 3828 17410 3834
rect 17366 3808 17381 3828
rect 17401 3808 17410 3828
rect 17366 3792 17410 3808
rect 17480 3824 17529 3834
rect 17480 3804 17491 3824
rect 17511 3804 17529 3824
rect 17480 3792 17529 3804
rect 17579 3828 17623 3834
rect 17579 3808 17594 3828
rect 17614 3808 17623 3828
rect 17579 3792 17623 3808
rect 17688 3824 17737 3834
rect 17688 3804 17699 3824
rect 17719 3804 17737 3824
rect 17688 3792 17737 3804
rect 17787 3828 17831 3834
rect 17787 3808 17802 3828
rect 17822 3808 17831 3828
rect 17787 3792 17831 3808
rect 17901 3828 17945 3834
rect 17901 3808 17910 3828
rect 17930 3808 17945 3828
rect 17901 3792 17945 3808
rect 17995 3824 18044 3834
rect 17995 3804 18013 3824
rect 18033 3804 18044 3824
rect 17995 3792 18044 3804
rect 13740 3704 13789 3716
rect 8360 3675 8409 3687
rect 1040 3571 1089 3583
rect 8360 3655 8371 3675
rect 8391 3655 8409 3675
rect 8360 3645 8409 3655
rect 8459 3671 8503 3687
rect 8459 3651 8474 3671
rect 8494 3651 8503 3671
rect 8459 3645 8503 3651
rect 8573 3671 8617 3687
rect 8573 3651 8582 3671
rect 8602 3651 8617 3671
rect 8573 3645 8617 3651
rect 8667 3675 8716 3687
rect 8667 3655 8685 3675
rect 8705 3655 8716 3675
rect 8667 3645 8716 3655
rect 8781 3671 8825 3687
rect 8781 3651 8790 3671
rect 8810 3651 8825 3671
rect 8781 3645 8825 3651
rect 8875 3675 8924 3687
rect 8875 3655 8893 3675
rect 8913 3655 8924 3675
rect 8875 3645 8924 3655
rect 8994 3671 9038 3687
rect 8994 3651 9003 3671
rect 9023 3651 9038 3671
rect 8994 3645 9038 3651
rect 9088 3675 9137 3687
rect 9088 3655 9106 3675
rect 9126 3655 9137 3675
rect 9088 3645 9137 3655
rect 5593 3582 5642 3592
rect 5593 3562 5604 3582
rect 5624 3562 5642 3582
rect 5593 3550 5642 3562
rect 5692 3586 5736 3592
rect 5692 3566 5707 3586
rect 5727 3566 5736 3586
rect 5692 3550 5736 3566
rect 5806 3582 5855 3592
rect 5806 3562 5817 3582
rect 5837 3562 5855 3582
rect 5806 3550 5855 3562
rect 5905 3586 5949 3592
rect 5905 3566 5920 3586
rect 5940 3566 5949 3586
rect 5905 3550 5949 3566
rect 6014 3582 6063 3592
rect 6014 3562 6025 3582
rect 6045 3562 6063 3582
rect 6014 3550 6063 3562
rect 6113 3586 6157 3592
rect 6113 3566 6128 3586
rect 6148 3566 6157 3586
rect 6113 3550 6157 3566
rect 6227 3586 6271 3592
rect 6227 3566 6236 3586
rect 6256 3566 6271 3586
rect 6227 3550 6271 3566
rect 6321 3582 6370 3592
rect 6321 3562 6339 3582
rect 6359 3562 6370 3582
rect 13740 3684 13751 3704
rect 13771 3684 13789 3704
rect 13740 3674 13789 3684
rect 13839 3700 13883 3716
rect 13839 3680 13854 3700
rect 13874 3680 13883 3700
rect 13839 3674 13883 3680
rect 13953 3700 13997 3716
rect 13953 3680 13962 3700
rect 13982 3680 13997 3700
rect 13953 3674 13997 3680
rect 14047 3704 14096 3716
rect 14047 3684 14065 3704
rect 14085 3684 14096 3704
rect 14047 3674 14096 3684
rect 14161 3700 14205 3716
rect 14161 3680 14170 3700
rect 14190 3680 14205 3700
rect 14161 3674 14205 3680
rect 14255 3704 14304 3716
rect 14255 3684 14273 3704
rect 14293 3684 14304 3704
rect 14255 3674 14304 3684
rect 14374 3700 14418 3716
rect 14374 3680 14383 3700
rect 14403 3680 14418 3700
rect 14374 3674 14418 3680
rect 14468 3704 14517 3716
rect 14468 3684 14486 3704
rect 14506 3684 14517 3704
rect 14468 3674 14517 3684
rect 6321 3550 6370 3562
rect 10973 3611 11022 3621
rect 10973 3591 10984 3611
rect 11004 3591 11022 3611
rect 10973 3579 11022 3591
rect 11072 3615 11116 3621
rect 11072 3595 11087 3615
rect 11107 3595 11116 3615
rect 11072 3579 11116 3595
rect 11186 3611 11235 3621
rect 11186 3591 11197 3611
rect 11217 3591 11235 3611
rect 11186 3579 11235 3591
rect 11285 3615 11329 3621
rect 11285 3595 11300 3615
rect 11320 3595 11329 3615
rect 11285 3579 11329 3595
rect 11394 3611 11443 3621
rect 11394 3591 11405 3611
rect 11425 3591 11443 3611
rect 11394 3579 11443 3591
rect 11493 3615 11537 3621
rect 11493 3595 11508 3615
rect 11528 3595 11537 3615
rect 11493 3579 11537 3595
rect 11607 3615 11651 3621
rect 11607 3595 11616 3615
rect 11636 3595 11651 3615
rect 11607 3579 11651 3595
rect 11701 3611 11750 3621
rect 11701 3591 11719 3611
rect 11739 3591 11750 3611
rect 19021 3683 19070 3695
rect 11701 3579 11750 3591
rect 19021 3663 19032 3683
rect 19052 3663 19070 3683
rect 19021 3653 19070 3663
rect 19120 3679 19164 3695
rect 19120 3659 19135 3679
rect 19155 3659 19164 3679
rect 19120 3653 19164 3659
rect 19234 3679 19278 3695
rect 19234 3659 19243 3679
rect 19263 3659 19278 3679
rect 19234 3653 19278 3659
rect 19328 3683 19377 3695
rect 19328 3663 19346 3683
rect 19366 3663 19377 3683
rect 19328 3653 19377 3663
rect 19442 3679 19486 3695
rect 19442 3659 19451 3679
rect 19471 3659 19486 3679
rect 19442 3653 19486 3659
rect 19536 3683 19585 3695
rect 19536 3663 19554 3683
rect 19574 3663 19585 3683
rect 19536 3653 19585 3663
rect 19655 3679 19699 3695
rect 19655 3659 19664 3679
rect 19684 3659 19699 3679
rect 19655 3653 19699 3659
rect 19749 3683 19798 3695
rect 19749 3663 19767 3683
rect 19787 3663 19798 3683
rect 19749 3653 19798 3663
rect 16254 3590 16303 3600
rect 16254 3570 16265 3590
rect 16285 3570 16303 3590
rect 16254 3558 16303 3570
rect 16353 3594 16397 3600
rect 16353 3574 16368 3594
rect 16388 3574 16397 3594
rect 16353 3558 16397 3574
rect 16467 3590 16516 3600
rect 16467 3570 16478 3590
rect 16498 3570 16516 3590
rect 16467 3558 16516 3570
rect 16566 3594 16610 3600
rect 16566 3574 16581 3594
rect 16601 3574 16610 3594
rect 16566 3558 16610 3574
rect 16675 3590 16724 3600
rect 16675 3570 16686 3590
rect 16706 3570 16724 3590
rect 16675 3558 16724 3570
rect 16774 3594 16818 3600
rect 16774 3574 16789 3594
rect 16809 3574 16818 3594
rect 16774 3558 16818 3574
rect 16888 3594 16932 3600
rect 16888 3574 16897 3594
rect 16917 3574 16932 3594
rect 16888 3558 16932 3574
rect 16982 3590 17031 3600
rect 16982 3570 17000 3590
rect 17020 3570 17031 3590
rect 16982 3558 17031 3570
rect 4147 3369 4196 3381
rect 4147 3349 4158 3369
rect 4178 3349 4196 3369
rect 4147 3339 4196 3349
rect 4246 3365 4290 3381
rect 4246 3345 4261 3365
rect 4281 3345 4290 3365
rect 4246 3339 4290 3345
rect 4360 3365 4404 3381
rect 4360 3345 4369 3365
rect 4389 3345 4404 3365
rect 4360 3339 4404 3345
rect 4454 3369 4503 3381
rect 4454 3349 4472 3369
rect 4492 3349 4503 3369
rect 4454 3339 4503 3349
rect 4568 3365 4612 3381
rect 4568 3345 4577 3365
rect 4597 3345 4612 3365
rect 4568 3339 4612 3345
rect 4662 3369 4711 3381
rect 4662 3349 4680 3369
rect 4700 3349 4711 3369
rect 4662 3339 4711 3349
rect 4781 3365 4825 3381
rect 4781 3345 4790 3365
rect 4810 3345 4825 3365
rect 4781 3339 4825 3345
rect 4875 3369 4924 3381
rect 4875 3349 4893 3369
rect 4913 3349 4924 3369
rect 4875 3339 4924 3349
rect 1380 3276 1429 3286
rect 1380 3256 1391 3276
rect 1411 3256 1429 3276
rect 1380 3244 1429 3256
rect 1479 3280 1523 3286
rect 1479 3260 1494 3280
rect 1514 3260 1523 3280
rect 1479 3244 1523 3260
rect 1593 3276 1642 3286
rect 1593 3256 1604 3276
rect 1624 3256 1642 3276
rect 1593 3244 1642 3256
rect 1692 3280 1736 3286
rect 1692 3260 1707 3280
rect 1727 3260 1736 3280
rect 1692 3244 1736 3260
rect 1801 3276 1850 3286
rect 1801 3256 1812 3276
rect 1832 3256 1850 3276
rect 1801 3244 1850 3256
rect 1900 3280 1944 3286
rect 1900 3260 1915 3280
rect 1935 3260 1944 3280
rect 1900 3244 1944 3260
rect 2014 3280 2058 3286
rect 2014 3260 2023 3280
rect 2043 3260 2058 3280
rect 2014 3244 2058 3260
rect 2108 3276 2157 3286
rect 2108 3256 2126 3276
rect 2146 3256 2157 3276
rect 9428 3348 9477 3360
rect 2108 3244 2157 3256
rect 9428 3328 9439 3348
rect 9459 3328 9477 3348
rect 9428 3318 9477 3328
rect 9527 3344 9571 3360
rect 9527 3324 9542 3344
rect 9562 3324 9571 3344
rect 9527 3318 9571 3324
rect 9641 3344 9685 3360
rect 9641 3324 9650 3344
rect 9670 3324 9685 3344
rect 9641 3318 9685 3324
rect 9735 3348 9784 3360
rect 9735 3328 9753 3348
rect 9773 3328 9784 3348
rect 9735 3318 9784 3328
rect 9849 3344 9893 3360
rect 9849 3324 9858 3344
rect 9878 3324 9893 3344
rect 9849 3318 9893 3324
rect 9943 3348 9992 3360
rect 9943 3328 9961 3348
rect 9981 3328 9992 3348
rect 9943 3318 9992 3328
rect 10062 3344 10106 3360
rect 10062 3324 10071 3344
rect 10091 3324 10106 3344
rect 10062 3318 10106 3324
rect 10156 3348 10205 3360
rect 10156 3328 10174 3348
rect 10194 3328 10205 3348
rect 10156 3318 10205 3328
rect 14808 3377 14857 3389
rect 6661 3255 6710 3265
rect 6661 3235 6672 3255
rect 6692 3235 6710 3255
rect 6661 3223 6710 3235
rect 6760 3259 6804 3265
rect 6760 3239 6775 3259
rect 6795 3239 6804 3259
rect 6760 3223 6804 3239
rect 6874 3255 6923 3265
rect 6874 3235 6885 3255
rect 6905 3235 6923 3255
rect 6874 3223 6923 3235
rect 6973 3259 7017 3265
rect 6973 3239 6988 3259
rect 7008 3239 7017 3259
rect 6973 3223 7017 3239
rect 7082 3255 7131 3265
rect 7082 3235 7093 3255
rect 7113 3235 7131 3255
rect 7082 3223 7131 3235
rect 7181 3259 7225 3265
rect 7181 3239 7196 3259
rect 7216 3239 7225 3259
rect 7181 3223 7225 3239
rect 7295 3259 7339 3265
rect 7295 3239 7304 3259
rect 7324 3239 7339 3259
rect 7295 3223 7339 3239
rect 7389 3255 7438 3265
rect 7389 3235 7407 3255
rect 7427 3235 7438 3255
rect 14808 3357 14819 3377
rect 14839 3357 14857 3377
rect 14808 3347 14857 3357
rect 14907 3373 14951 3389
rect 14907 3353 14922 3373
rect 14942 3353 14951 3373
rect 14907 3347 14951 3353
rect 15021 3373 15065 3389
rect 15021 3353 15030 3373
rect 15050 3353 15065 3373
rect 15021 3347 15065 3353
rect 15115 3377 15164 3389
rect 15115 3357 15133 3377
rect 15153 3357 15164 3377
rect 15115 3347 15164 3357
rect 15229 3373 15273 3389
rect 15229 3353 15238 3373
rect 15258 3353 15273 3373
rect 15229 3347 15273 3353
rect 15323 3377 15372 3389
rect 15323 3357 15341 3377
rect 15361 3357 15372 3377
rect 15323 3347 15372 3357
rect 15442 3373 15486 3389
rect 15442 3353 15451 3373
rect 15471 3353 15486 3373
rect 15442 3347 15486 3353
rect 15536 3377 15585 3389
rect 15536 3357 15554 3377
rect 15574 3357 15585 3377
rect 15536 3347 15585 3357
rect 12041 3284 12090 3294
rect 12041 3264 12052 3284
rect 12072 3264 12090 3284
rect 12041 3252 12090 3264
rect 12140 3288 12184 3294
rect 12140 3268 12155 3288
rect 12175 3268 12184 3288
rect 12140 3252 12184 3268
rect 12254 3284 12303 3294
rect 12254 3264 12265 3284
rect 12285 3264 12303 3284
rect 12254 3252 12303 3264
rect 12353 3288 12397 3294
rect 12353 3268 12368 3288
rect 12388 3268 12397 3288
rect 12353 3252 12397 3268
rect 12462 3284 12511 3294
rect 12462 3264 12473 3284
rect 12493 3264 12511 3284
rect 12462 3252 12511 3264
rect 12561 3288 12605 3294
rect 12561 3268 12576 3288
rect 12596 3268 12605 3288
rect 12561 3252 12605 3268
rect 12675 3288 12719 3294
rect 12675 3268 12684 3288
rect 12704 3268 12719 3288
rect 12675 3252 12719 3268
rect 12769 3284 12818 3294
rect 12769 3264 12787 3284
rect 12807 3264 12818 3284
rect 20089 3356 20138 3368
rect 12769 3252 12818 3264
rect 7389 3223 7438 3235
rect 3134 3135 3183 3147
rect 3134 3115 3145 3135
rect 3165 3115 3183 3135
rect 3134 3105 3183 3115
rect 3233 3131 3277 3147
rect 3233 3111 3248 3131
rect 3268 3111 3277 3131
rect 3233 3105 3277 3111
rect 3347 3131 3391 3147
rect 3347 3111 3356 3131
rect 3376 3111 3391 3131
rect 3347 3105 3391 3111
rect 3441 3135 3490 3147
rect 3441 3115 3459 3135
rect 3479 3115 3490 3135
rect 3441 3105 3490 3115
rect 3555 3131 3599 3147
rect 3555 3111 3564 3131
rect 3584 3111 3599 3131
rect 3555 3105 3599 3111
rect 3649 3135 3698 3147
rect 3649 3115 3667 3135
rect 3687 3115 3698 3135
rect 3649 3105 3698 3115
rect 3768 3131 3812 3147
rect 3768 3111 3777 3131
rect 3797 3111 3812 3131
rect 3768 3105 3812 3111
rect 3862 3135 3911 3147
rect 3862 3115 3880 3135
rect 3900 3115 3911 3135
rect 3862 3105 3911 3115
rect 318 3037 367 3047
rect 318 3017 329 3037
rect 349 3017 367 3037
rect 318 3005 367 3017
rect 417 3041 461 3047
rect 417 3021 432 3041
rect 452 3021 461 3041
rect 417 3005 461 3021
rect 531 3037 580 3047
rect 531 3017 542 3037
rect 562 3017 580 3037
rect 531 3005 580 3017
rect 630 3041 674 3047
rect 630 3021 645 3041
rect 665 3021 674 3041
rect 630 3005 674 3021
rect 739 3037 788 3047
rect 739 3017 750 3037
rect 770 3017 788 3037
rect 739 3005 788 3017
rect 838 3041 882 3047
rect 838 3021 853 3041
rect 873 3021 882 3041
rect 838 3005 882 3021
rect 952 3041 996 3047
rect 952 3021 961 3041
rect 981 3021 996 3041
rect 952 3005 996 3021
rect 1046 3037 1095 3047
rect 1046 3017 1064 3037
rect 1084 3017 1095 3037
rect 1046 3005 1095 3017
rect 8415 3114 8464 3126
rect 8415 3094 8426 3114
rect 8446 3094 8464 3114
rect 8415 3084 8464 3094
rect 8514 3110 8558 3126
rect 8514 3090 8529 3110
rect 8549 3090 8558 3110
rect 8514 3084 8558 3090
rect 8628 3110 8672 3126
rect 8628 3090 8637 3110
rect 8657 3090 8672 3110
rect 8628 3084 8672 3090
rect 8722 3114 8771 3126
rect 8722 3094 8740 3114
rect 8760 3094 8771 3114
rect 8722 3084 8771 3094
rect 8836 3110 8880 3126
rect 8836 3090 8845 3110
rect 8865 3090 8880 3110
rect 8836 3084 8880 3090
rect 8930 3114 8979 3126
rect 8930 3094 8948 3114
rect 8968 3094 8979 3114
rect 8930 3084 8979 3094
rect 9049 3110 9093 3126
rect 9049 3090 9058 3110
rect 9078 3090 9093 3110
rect 9049 3084 9093 3090
rect 9143 3114 9192 3126
rect 9143 3094 9161 3114
rect 9181 3094 9192 3114
rect 20089 3336 20100 3356
rect 20120 3336 20138 3356
rect 20089 3326 20138 3336
rect 20188 3352 20232 3368
rect 20188 3332 20203 3352
rect 20223 3332 20232 3352
rect 20188 3326 20232 3332
rect 20302 3352 20346 3368
rect 20302 3332 20311 3352
rect 20331 3332 20346 3352
rect 20302 3326 20346 3332
rect 20396 3356 20445 3368
rect 20396 3336 20414 3356
rect 20434 3336 20445 3356
rect 20396 3326 20445 3336
rect 20510 3352 20554 3368
rect 20510 3332 20519 3352
rect 20539 3332 20554 3352
rect 20510 3326 20554 3332
rect 20604 3356 20653 3368
rect 20604 3336 20622 3356
rect 20642 3336 20653 3356
rect 20604 3326 20653 3336
rect 20723 3352 20767 3368
rect 20723 3332 20732 3352
rect 20752 3332 20767 3352
rect 20723 3326 20767 3332
rect 20817 3356 20866 3368
rect 20817 3336 20835 3356
rect 20855 3336 20866 3356
rect 20817 3326 20866 3336
rect 17322 3263 17371 3273
rect 17322 3243 17333 3263
rect 17353 3243 17371 3263
rect 17322 3231 17371 3243
rect 17421 3267 17465 3273
rect 17421 3247 17436 3267
rect 17456 3247 17465 3267
rect 17421 3231 17465 3247
rect 17535 3263 17584 3273
rect 17535 3243 17546 3263
rect 17566 3243 17584 3263
rect 17535 3231 17584 3243
rect 17634 3267 17678 3273
rect 17634 3247 17649 3267
rect 17669 3247 17678 3267
rect 17634 3231 17678 3247
rect 17743 3263 17792 3273
rect 17743 3243 17754 3263
rect 17774 3243 17792 3263
rect 17743 3231 17792 3243
rect 17842 3267 17886 3273
rect 17842 3247 17857 3267
rect 17877 3247 17886 3267
rect 17842 3231 17886 3247
rect 17956 3267 18000 3273
rect 17956 3247 17965 3267
rect 17985 3247 18000 3267
rect 17956 3231 18000 3247
rect 18050 3263 18099 3273
rect 18050 3243 18068 3263
rect 18088 3243 18099 3263
rect 18050 3231 18099 3243
rect 13795 3143 13844 3155
rect 9143 3084 9192 3094
rect 5599 3016 5648 3026
rect 5599 2996 5610 3016
rect 5630 2996 5648 3016
rect 5599 2984 5648 2996
rect 5698 3020 5742 3026
rect 5698 3000 5713 3020
rect 5733 3000 5742 3020
rect 5698 2984 5742 3000
rect 5812 3016 5861 3026
rect 5812 2996 5823 3016
rect 5843 2996 5861 3016
rect 5812 2984 5861 2996
rect 5911 3020 5955 3026
rect 5911 3000 5926 3020
rect 5946 3000 5955 3020
rect 5911 2984 5955 3000
rect 6020 3016 6069 3026
rect 6020 2996 6031 3016
rect 6051 2996 6069 3016
rect 6020 2984 6069 2996
rect 6119 3020 6163 3026
rect 6119 3000 6134 3020
rect 6154 3000 6163 3020
rect 6119 2984 6163 3000
rect 6233 3020 6277 3026
rect 6233 3000 6242 3020
rect 6262 3000 6277 3020
rect 6233 2984 6277 3000
rect 6327 3016 6376 3026
rect 6327 2996 6345 3016
rect 6365 2996 6376 3016
rect 6327 2984 6376 2996
rect 4146 2954 4195 2966
rect 4146 2934 4157 2954
rect 4177 2934 4195 2954
rect 4146 2924 4195 2934
rect 4245 2950 4289 2966
rect 4245 2930 4260 2950
rect 4280 2930 4289 2950
rect 4245 2924 4289 2930
rect 4359 2950 4403 2966
rect 4359 2930 4368 2950
rect 4388 2930 4403 2950
rect 4359 2924 4403 2930
rect 4453 2954 4502 2966
rect 4453 2934 4471 2954
rect 4491 2934 4502 2954
rect 4453 2924 4502 2934
rect 4567 2950 4611 2966
rect 4567 2930 4576 2950
rect 4596 2930 4611 2950
rect 4567 2924 4611 2930
rect 4661 2954 4710 2966
rect 4661 2934 4679 2954
rect 4699 2934 4710 2954
rect 4661 2924 4710 2934
rect 4780 2950 4824 2966
rect 4780 2930 4789 2950
rect 4809 2930 4824 2950
rect 4780 2924 4824 2930
rect 4874 2954 4923 2966
rect 4874 2934 4892 2954
rect 4912 2934 4923 2954
rect 4874 2924 4923 2934
rect 1330 2856 1379 2866
rect 1330 2836 1341 2856
rect 1361 2836 1379 2856
rect 1330 2824 1379 2836
rect 1429 2860 1473 2866
rect 1429 2840 1444 2860
rect 1464 2840 1473 2860
rect 1429 2824 1473 2840
rect 1543 2856 1592 2866
rect 1543 2836 1554 2856
rect 1574 2836 1592 2856
rect 1543 2824 1592 2836
rect 1642 2860 1686 2866
rect 1642 2840 1657 2860
rect 1677 2840 1686 2860
rect 1642 2824 1686 2840
rect 1751 2856 1800 2866
rect 1751 2836 1762 2856
rect 1782 2836 1800 2856
rect 1751 2824 1800 2836
rect 1850 2860 1894 2866
rect 1850 2840 1865 2860
rect 1885 2840 1894 2860
rect 1850 2824 1894 2840
rect 1964 2860 2008 2866
rect 1964 2840 1973 2860
rect 1993 2840 2008 2860
rect 1964 2824 2008 2840
rect 2058 2856 2107 2866
rect 2058 2836 2076 2856
rect 2096 2836 2107 2856
rect 13795 3123 13806 3143
rect 13826 3123 13844 3143
rect 13795 3113 13844 3123
rect 13894 3139 13938 3155
rect 13894 3119 13909 3139
rect 13929 3119 13938 3139
rect 13894 3113 13938 3119
rect 14008 3139 14052 3155
rect 14008 3119 14017 3139
rect 14037 3119 14052 3139
rect 14008 3113 14052 3119
rect 14102 3143 14151 3155
rect 14102 3123 14120 3143
rect 14140 3123 14151 3143
rect 14102 3113 14151 3123
rect 14216 3139 14260 3155
rect 14216 3119 14225 3139
rect 14245 3119 14260 3139
rect 14216 3113 14260 3119
rect 14310 3143 14359 3155
rect 14310 3123 14328 3143
rect 14348 3123 14359 3143
rect 14310 3113 14359 3123
rect 14429 3139 14473 3155
rect 14429 3119 14438 3139
rect 14458 3119 14473 3139
rect 14429 3113 14473 3119
rect 14523 3143 14572 3155
rect 14523 3123 14541 3143
rect 14561 3123 14572 3143
rect 14523 3113 14572 3123
rect 10979 3045 11028 3055
rect 10979 3025 10990 3045
rect 11010 3025 11028 3045
rect 10979 3013 11028 3025
rect 11078 3049 11122 3055
rect 11078 3029 11093 3049
rect 11113 3029 11122 3049
rect 11078 3013 11122 3029
rect 11192 3045 11241 3055
rect 11192 3025 11203 3045
rect 11223 3025 11241 3045
rect 11192 3013 11241 3025
rect 11291 3049 11335 3055
rect 11291 3029 11306 3049
rect 11326 3029 11335 3049
rect 11291 3013 11335 3029
rect 11400 3045 11449 3055
rect 11400 3025 11411 3045
rect 11431 3025 11449 3045
rect 11400 3013 11449 3025
rect 11499 3049 11543 3055
rect 11499 3029 11514 3049
rect 11534 3029 11543 3049
rect 11499 3013 11543 3029
rect 11613 3049 11657 3055
rect 11613 3029 11622 3049
rect 11642 3029 11657 3049
rect 11613 3013 11657 3029
rect 11707 3045 11756 3055
rect 11707 3025 11725 3045
rect 11745 3025 11756 3045
rect 11707 3013 11756 3025
rect 2058 2824 2107 2836
rect 19076 3122 19125 3134
rect 9427 2933 9476 2945
rect 9427 2913 9438 2933
rect 9458 2913 9476 2933
rect 9427 2903 9476 2913
rect 9526 2929 9570 2945
rect 9526 2909 9541 2929
rect 9561 2909 9570 2929
rect 9526 2903 9570 2909
rect 9640 2929 9684 2945
rect 9640 2909 9649 2929
rect 9669 2909 9684 2929
rect 9640 2903 9684 2909
rect 9734 2933 9783 2945
rect 9734 2913 9752 2933
rect 9772 2913 9783 2933
rect 9734 2903 9783 2913
rect 9848 2929 9892 2945
rect 9848 2909 9857 2929
rect 9877 2909 9892 2929
rect 9848 2903 9892 2909
rect 9942 2933 9991 2945
rect 9942 2913 9960 2933
rect 9980 2913 9991 2933
rect 9942 2903 9991 2913
rect 10061 2929 10105 2945
rect 10061 2909 10070 2929
rect 10090 2909 10105 2929
rect 10061 2903 10105 2909
rect 10155 2933 10204 2945
rect 10155 2913 10173 2933
rect 10193 2913 10204 2933
rect 10155 2903 10204 2913
rect 6611 2835 6660 2845
rect 6611 2815 6622 2835
rect 6642 2815 6660 2835
rect 6611 2803 6660 2815
rect 6710 2839 6754 2845
rect 6710 2819 6725 2839
rect 6745 2819 6754 2839
rect 6710 2803 6754 2819
rect 6824 2835 6873 2845
rect 6824 2815 6835 2835
rect 6855 2815 6873 2835
rect 6824 2803 6873 2815
rect 6923 2839 6967 2845
rect 6923 2819 6938 2839
rect 6958 2819 6967 2839
rect 6923 2803 6967 2819
rect 7032 2835 7081 2845
rect 7032 2815 7043 2835
rect 7063 2815 7081 2835
rect 7032 2803 7081 2815
rect 7131 2839 7175 2845
rect 7131 2819 7146 2839
rect 7166 2819 7175 2839
rect 7131 2803 7175 2819
rect 7245 2839 7289 2845
rect 7245 2819 7254 2839
rect 7274 2819 7289 2839
rect 7245 2803 7289 2819
rect 7339 2835 7388 2845
rect 7339 2815 7357 2835
rect 7377 2815 7388 2835
rect 19076 3102 19087 3122
rect 19107 3102 19125 3122
rect 19076 3092 19125 3102
rect 19175 3118 19219 3134
rect 19175 3098 19190 3118
rect 19210 3098 19219 3118
rect 19175 3092 19219 3098
rect 19289 3118 19333 3134
rect 19289 3098 19298 3118
rect 19318 3098 19333 3118
rect 19289 3092 19333 3098
rect 19383 3122 19432 3134
rect 19383 3102 19401 3122
rect 19421 3102 19432 3122
rect 19383 3092 19432 3102
rect 19497 3118 19541 3134
rect 19497 3098 19506 3118
rect 19526 3098 19541 3118
rect 19497 3092 19541 3098
rect 19591 3122 19640 3134
rect 19591 3102 19609 3122
rect 19629 3102 19640 3122
rect 19591 3092 19640 3102
rect 19710 3118 19754 3134
rect 19710 3098 19719 3118
rect 19739 3098 19754 3118
rect 19710 3092 19754 3098
rect 19804 3122 19853 3134
rect 19804 3102 19822 3122
rect 19842 3102 19853 3122
rect 19804 3092 19853 3102
rect 16260 3024 16309 3034
rect 16260 3004 16271 3024
rect 16291 3004 16309 3024
rect 16260 2992 16309 3004
rect 16359 3028 16403 3034
rect 16359 3008 16374 3028
rect 16394 3008 16403 3028
rect 16359 2992 16403 3008
rect 16473 3024 16522 3034
rect 16473 3004 16484 3024
rect 16504 3004 16522 3024
rect 16473 2992 16522 3004
rect 16572 3028 16616 3034
rect 16572 3008 16587 3028
rect 16607 3008 16616 3028
rect 16572 2992 16616 3008
rect 16681 3024 16730 3034
rect 16681 3004 16692 3024
rect 16712 3004 16730 3024
rect 16681 2992 16730 3004
rect 16780 3028 16824 3034
rect 16780 3008 16795 3028
rect 16815 3008 16824 3028
rect 16780 2992 16824 3008
rect 16894 3028 16938 3034
rect 16894 3008 16903 3028
rect 16923 3008 16938 3028
rect 16894 2992 16938 3008
rect 16988 3024 17037 3034
rect 16988 3004 17006 3024
rect 17026 3004 17037 3024
rect 16988 2992 17037 3004
rect 14807 2962 14856 2974
rect 14807 2942 14818 2962
rect 14838 2942 14856 2962
rect 14807 2932 14856 2942
rect 14906 2958 14950 2974
rect 14906 2938 14921 2958
rect 14941 2938 14950 2958
rect 14906 2932 14950 2938
rect 15020 2958 15064 2974
rect 15020 2938 15029 2958
rect 15049 2938 15064 2958
rect 15020 2932 15064 2938
rect 15114 2962 15163 2974
rect 15114 2942 15132 2962
rect 15152 2942 15163 2962
rect 15114 2932 15163 2942
rect 15228 2958 15272 2974
rect 15228 2938 15237 2958
rect 15257 2938 15272 2958
rect 15228 2932 15272 2938
rect 15322 2962 15371 2974
rect 15322 2942 15340 2962
rect 15360 2942 15371 2962
rect 15322 2932 15371 2942
rect 15441 2958 15485 2974
rect 15441 2938 15450 2958
rect 15470 2938 15485 2958
rect 15441 2932 15485 2938
rect 15535 2962 15584 2974
rect 15535 2942 15553 2962
rect 15573 2942 15584 2962
rect 15535 2932 15584 2942
rect 11991 2864 12040 2874
rect 7339 2803 7388 2815
rect 2926 2668 2975 2680
rect 2926 2648 2937 2668
rect 2957 2648 2975 2668
rect 2926 2638 2975 2648
rect 3025 2664 3069 2680
rect 3025 2644 3040 2664
rect 3060 2644 3069 2664
rect 3025 2638 3069 2644
rect 3139 2664 3183 2680
rect 3139 2644 3148 2664
rect 3168 2644 3183 2664
rect 3139 2638 3183 2644
rect 3233 2668 3282 2680
rect 3233 2648 3251 2668
rect 3271 2648 3282 2668
rect 3233 2638 3282 2648
rect 3347 2664 3391 2680
rect 3347 2644 3356 2664
rect 3376 2644 3391 2664
rect 3347 2638 3391 2644
rect 3441 2668 3490 2680
rect 3441 2648 3459 2668
rect 3479 2648 3490 2668
rect 3441 2638 3490 2648
rect 3560 2664 3604 2680
rect 3560 2644 3569 2664
rect 3589 2644 3604 2664
rect 3560 2638 3604 2644
rect 3654 2668 3703 2680
rect 3654 2648 3672 2668
rect 3692 2648 3703 2668
rect 3654 2638 3703 2648
rect 11991 2844 12002 2864
rect 12022 2844 12040 2864
rect 11991 2832 12040 2844
rect 12090 2868 12134 2874
rect 12090 2848 12105 2868
rect 12125 2848 12134 2868
rect 12090 2832 12134 2848
rect 12204 2864 12253 2874
rect 12204 2844 12215 2864
rect 12235 2844 12253 2864
rect 12204 2832 12253 2844
rect 12303 2868 12347 2874
rect 12303 2848 12318 2868
rect 12338 2848 12347 2868
rect 12303 2832 12347 2848
rect 12412 2864 12461 2874
rect 12412 2844 12423 2864
rect 12443 2844 12461 2864
rect 12412 2832 12461 2844
rect 12511 2868 12555 2874
rect 12511 2848 12526 2868
rect 12546 2848 12555 2868
rect 12511 2832 12555 2848
rect 12625 2868 12669 2874
rect 12625 2848 12634 2868
rect 12654 2848 12669 2868
rect 12625 2832 12669 2848
rect 12719 2864 12768 2874
rect 12719 2844 12737 2864
rect 12757 2844 12768 2864
rect 12719 2832 12768 2844
rect 20088 2941 20137 2953
rect 20088 2921 20099 2941
rect 20119 2921 20137 2941
rect 20088 2911 20137 2921
rect 20187 2937 20231 2953
rect 20187 2917 20202 2937
rect 20222 2917 20231 2937
rect 20187 2911 20231 2917
rect 20301 2937 20345 2953
rect 20301 2917 20310 2937
rect 20330 2917 20345 2937
rect 20301 2911 20345 2917
rect 20395 2941 20444 2953
rect 20395 2921 20413 2941
rect 20433 2921 20444 2941
rect 20395 2911 20444 2921
rect 20509 2937 20553 2953
rect 20509 2917 20518 2937
rect 20538 2917 20553 2937
rect 20509 2911 20553 2917
rect 20603 2941 20652 2953
rect 20603 2921 20621 2941
rect 20641 2921 20652 2941
rect 20603 2911 20652 2921
rect 20722 2937 20766 2953
rect 20722 2917 20731 2937
rect 20751 2917 20766 2937
rect 20722 2911 20766 2917
rect 20816 2941 20865 2953
rect 20816 2921 20834 2941
rect 20854 2921 20865 2941
rect 20816 2911 20865 2921
rect 17272 2843 17321 2853
rect 17272 2823 17283 2843
rect 17303 2823 17321 2843
rect 17272 2811 17321 2823
rect 17371 2847 17415 2853
rect 17371 2827 17386 2847
rect 17406 2827 17415 2847
rect 17371 2811 17415 2827
rect 17485 2843 17534 2853
rect 17485 2823 17496 2843
rect 17516 2823 17534 2843
rect 17485 2811 17534 2823
rect 17584 2847 17628 2853
rect 17584 2827 17599 2847
rect 17619 2827 17628 2847
rect 17584 2811 17628 2827
rect 17693 2843 17742 2853
rect 17693 2823 17704 2843
rect 17724 2823 17742 2843
rect 17693 2811 17742 2823
rect 17792 2847 17836 2853
rect 17792 2827 17807 2847
rect 17827 2827 17836 2847
rect 17792 2811 17836 2827
rect 17906 2847 17950 2853
rect 17906 2827 17915 2847
rect 17935 2827 17950 2847
rect 17906 2811 17950 2827
rect 18000 2843 18049 2853
rect 18000 2823 18018 2843
rect 18038 2823 18049 2843
rect 18000 2811 18049 2823
rect 317 2622 366 2632
rect 317 2602 328 2622
rect 348 2602 366 2622
rect 317 2590 366 2602
rect 416 2626 460 2632
rect 416 2606 431 2626
rect 451 2606 460 2626
rect 416 2590 460 2606
rect 530 2622 579 2632
rect 530 2602 541 2622
rect 561 2602 579 2622
rect 530 2590 579 2602
rect 629 2626 673 2632
rect 629 2606 644 2626
rect 664 2606 673 2626
rect 629 2590 673 2606
rect 738 2622 787 2632
rect 738 2602 749 2622
rect 769 2602 787 2622
rect 738 2590 787 2602
rect 837 2626 881 2632
rect 837 2606 852 2626
rect 872 2606 881 2626
rect 837 2590 881 2606
rect 951 2626 995 2632
rect 951 2606 960 2626
rect 980 2606 995 2626
rect 951 2590 995 2606
rect 1045 2622 1094 2632
rect 1045 2602 1063 2622
rect 1083 2602 1094 2622
rect 1045 2590 1094 2602
rect 8207 2647 8256 2659
rect 8207 2627 8218 2647
rect 8238 2627 8256 2647
rect 8207 2617 8256 2627
rect 8306 2643 8350 2659
rect 8306 2623 8321 2643
rect 8341 2623 8350 2643
rect 8306 2617 8350 2623
rect 8420 2643 8464 2659
rect 8420 2623 8429 2643
rect 8449 2623 8464 2643
rect 8420 2617 8464 2623
rect 8514 2647 8563 2659
rect 8514 2627 8532 2647
rect 8552 2627 8563 2647
rect 8514 2617 8563 2627
rect 8628 2643 8672 2659
rect 8628 2623 8637 2643
rect 8657 2623 8672 2643
rect 8628 2617 8672 2623
rect 8722 2647 8771 2659
rect 8722 2627 8740 2647
rect 8760 2627 8771 2647
rect 8722 2617 8771 2627
rect 8841 2643 8885 2659
rect 8841 2623 8850 2643
rect 8870 2623 8885 2643
rect 8841 2617 8885 2623
rect 8935 2647 8984 2659
rect 8935 2627 8953 2647
rect 8973 2627 8984 2647
rect 8935 2617 8984 2627
rect 5598 2601 5647 2611
rect 5598 2581 5609 2601
rect 5629 2581 5647 2601
rect 5598 2569 5647 2581
rect 5697 2605 5741 2611
rect 5697 2585 5712 2605
rect 5732 2585 5741 2605
rect 5697 2569 5741 2585
rect 5811 2601 5860 2611
rect 5811 2581 5822 2601
rect 5842 2581 5860 2601
rect 5811 2569 5860 2581
rect 5910 2605 5954 2611
rect 5910 2585 5925 2605
rect 5945 2585 5954 2605
rect 5910 2569 5954 2585
rect 6019 2601 6068 2611
rect 6019 2581 6030 2601
rect 6050 2581 6068 2601
rect 6019 2569 6068 2581
rect 6118 2605 6162 2611
rect 6118 2585 6133 2605
rect 6153 2585 6162 2605
rect 6118 2569 6162 2585
rect 6232 2605 6276 2611
rect 6232 2585 6241 2605
rect 6261 2585 6276 2605
rect 6232 2569 6276 2585
rect 6326 2601 6375 2611
rect 6326 2581 6344 2601
rect 6364 2581 6375 2601
rect 6326 2569 6375 2581
rect 13587 2676 13636 2688
rect 13587 2656 13598 2676
rect 13618 2656 13636 2676
rect 13587 2646 13636 2656
rect 13686 2672 13730 2688
rect 13686 2652 13701 2672
rect 13721 2652 13730 2672
rect 13686 2646 13730 2652
rect 13800 2672 13844 2688
rect 13800 2652 13809 2672
rect 13829 2652 13844 2672
rect 13800 2646 13844 2652
rect 13894 2676 13943 2688
rect 13894 2656 13912 2676
rect 13932 2656 13943 2676
rect 13894 2646 13943 2656
rect 14008 2672 14052 2688
rect 14008 2652 14017 2672
rect 14037 2652 14052 2672
rect 14008 2646 14052 2652
rect 14102 2676 14151 2688
rect 14102 2656 14120 2676
rect 14140 2656 14151 2676
rect 14102 2646 14151 2656
rect 14221 2672 14265 2688
rect 14221 2652 14230 2672
rect 14250 2652 14265 2672
rect 14221 2646 14265 2652
rect 14315 2676 14364 2688
rect 14315 2656 14333 2676
rect 14353 2656 14364 2676
rect 14315 2646 14364 2656
rect 10978 2630 11027 2640
rect 10978 2610 10989 2630
rect 11009 2610 11027 2630
rect 10978 2598 11027 2610
rect 11077 2634 11121 2640
rect 11077 2614 11092 2634
rect 11112 2614 11121 2634
rect 11077 2598 11121 2614
rect 11191 2630 11240 2640
rect 11191 2610 11202 2630
rect 11222 2610 11240 2630
rect 11191 2598 11240 2610
rect 11290 2634 11334 2640
rect 11290 2614 11305 2634
rect 11325 2614 11334 2634
rect 11290 2598 11334 2614
rect 11399 2630 11448 2640
rect 11399 2610 11410 2630
rect 11430 2610 11448 2630
rect 11399 2598 11448 2610
rect 11498 2634 11542 2640
rect 11498 2614 11513 2634
rect 11533 2614 11542 2634
rect 11498 2598 11542 2614
rect 11612 2634 11656 2640
rect 11612 2614 11621 2634
rect 11641 2614 11656 2634
rect 11612 2598 11656 2614
rect 11706 2630 11755 2640
rect 11706 2610 11724 2630
rect 11744 2610 11755 2630
rect 11706 2598 11755 2610
rect 18868 2655 18917 2667
rect 18868 2635 18879 2655
rect 18899 2635 18917 2655
rect 18868 2625 18917 2635
rect 18967 2651 19011 2667
rect 18967 2631 18982 2651
rect 19002 2631 19011 2651
rect 18967 2625 19011 2631
rect 19081 2651 19125 2667
rect 19081 2631 19090 2651
rect 19110 2631 19125 2651
rect 19081 2625 19125 2631
rect 19175 2655 19224 2667
rect 19175 2635 19193 2655
rect 19213 2635 19224 2655
rect 19175 2625 19224 2635
rect 19289 2651 19333 2667
rect 19289 2631 19298 2651
rect 19318 2631 19333 2651
rect 19289 2625 19333 2631
rect 19383 2655 19432 2667
rect 19383 2635 19401 2655
rect 19421 2635 19432 2655
rect 19383 2625 19432 2635
rect 19502 2651 19546 2667
rect 19502 2631 19511 2651
rect 19531 2631 19546 2651
rect 19502 2625 19546 2631
rect 19596 2655 19645 2667
rect 19596 2635 19614 2655
rect 19634 2635 19645 2655
rect 19596 2625 19645 2635
rect 4154 2390 4203 2402
rect 4154 2370 4165 2390
rect 4185 2370 4203 2390
rect 4154 2360 4203 2370
rect 4253 2386 4297 2402
rect 4253 2366 4268 2386
rect 4288 2366 4297 2386
rect 4253 2360 4297 2366
rect 4367 2386 4411 2402
rect 4367 2366 4376 2386
rect 4396 2366 4411 2386
rect 4367 2360 4411 2366
rect 4461 2390 4510 2402
rect 4461 2370 4479 2390
rect 4499 2370 4510 2390
rect 4461 2360 4510 2370
rect 4575 2386 4619 2402
rect 4575 2366 4584 2386
rect 4604 2366 4619 2386
rect 4575 2360 4619 2366
rect 4669 2390 4718 2402
rect 4669 2370 4687 2390
rect 4707 2370 4718 2390
rect 4669 2360 4718 2370
rect 4788 2386 4832 2402
rect 4788 2366 4797 2386
rect 4817 2366 4832 2386
rect 4788 2360 4832 2366
rect 4882 2390 4931 2402
rect 4882 2370 4900 2390
rect 4920 2370 4931 2390
rect 4882 2360 4931 2370
rect 16259 2609 16308 2619
rect 16259 2589 16270 2609
rect 16290 2589 16308 2609
rect 16259 2577 16308 2589
rect 16358 2613 16402 2619
rect 16358 2593 16373 2613
rect 16393 2593 16402 2613
rect 16358 2577 16402 2593
rect 16472 2609 16521 2619
rect 16472 2589 16483 2609
rect 16503 2589 16521 2609
rect 16472 2577 16521 2589
rect 16571 2613 16615 2619
rect 16571 2593 16586 2613
rect 16606 2593 16615 2613
rect 16571 2577 16615 2593
rect 16680 2609 16729 2619
rect 16680 2589 16691 2609
rect 16711 2589 16729 2609
rect 16680 2577 16729 2589
rect 16779 2613 16823 2619
rect 16779 2593 16794 2613
rect 16814 2593 16823 2613
rect 16779 2577 16823 2593
rect 16893 2613 16937 2619
rect 16893 2593 16902 2613
rect 16922 2593 16937 2613
rect 16893 2577 16937 2593
rect 16987 2609 17036 2619
rect 16987 2589 17005 2609
rect 17025 2589 17036 2609
rect 16987 2577 17036 2589
rect 1545 2344 1594 2354
rect 1545 2324 1556 2344
rect 1576 2324 1594 2344
rect 1545 2312 1594 2324
rect 1644 2348 1688 2354
rect 1644 2328 1659 2348
rect 1679 2328 1688 2348
rect 1644 2312 1688 2328
rect 1758 2344 1807 2354
rect 1758 2324 1769 2344
rect 1789 2324 1807 2344
rect 1758 2312 1807 2324
rect 1857 2348 1901 2354
rect 1857 2328 1872 2348
rect 1892 2328 1901 2348
rect 1857 2312 1901 2328
rect 1966 2344 2015 2354
rect 1966 2324 1977 2344
rect 1997 2324 2015 2344
rect 1966 2312 2015 2324
rect 2065 2348 2109 2354
rect 2065 2328 2080 2348
rect 2100 2328 2109 2348
rect 2065 2312 2109 2328
rect 2179 2348 2223 2354
rect 2179 2328 2188 2348
rect 2208 2328 2223 2348
rect 2179 2312 2223 2328
rect 2273 2344 2322 2354
rect 2273 2324 2291 2344
rect 2311 2324 2322 2344
rect 2273 2312 2322 2324
rect 9435 2369 9484 2381
rect 9435 2349 9446 2369
rect 9466 2349 9484 2369
rect 9435 2339 9484 2349
rect 9534 2365 9578 2381
rect 9534 2345 9549 2365
rect 9569 2345 9578 2365
rect 9534 2339 9578 2345
rect 9648 2365 9692 2381
rect 9648 2345 9657 2365
rect 9677 2345 9692 2365
rect 9648 2339 9692 2345
rect 9742 2369 9791 2381
rect 9742 2349 9760 2369
rect 9780 2349 9791 2369
rect 9742 2339 9791 2349
rect 9856 2365 9900 2381
rect 9856 2345 9865 2365
rect 9885 2345 9900 2365
rect 9856 2339 9900 2345
rect 9950 2369 9999 2381
rect 9950 2349 9968 2369
rect 9988 2349 9999 2369
rect 9950 2339 9999 2349
rect 10069 2365 10113 2381
rect 10069 2345 10078 2365
rect 10098 2345 10113 2365
rect 10069 2339 10113 2345
rect 10163 2369 10212 2381
rect 10163 2349 10181 2369
rect 10201 2349 10212 2369
rect 10163 2339 10212 2349
rect 6826 2323 6875 2333
rect 6826 2303 6837 2323
rect 6857 2303 6875 2323
rect 6826 2291 6875 2303
rect 6925 2327 6969 2333
rect 6925 2307 6940 2327
rect 6960 2307 6969 2327
rect 6925 2291 6969 2307
rect 7039 2323 7088 2333
rect 7039 2303 7050 2323
rect 7070 2303 7088 2323
rect 7039 2291 7088 2303
rect 7138 2327 7182 2333
rect 7138 2307 7153 2327
rect 7173 2307 7182 2327
rect 7138 2291 7182 2307
rect 7247 2323 7296 2333
rect 7247 2303 7258 2323
rect 7278 2303 7296 2323
rect 7247 2291 7296 2303
rect 7346 2327 7390 2333
rect 7346 2307 7361 2327
rect 7381 2307 7390 2327
rect 7346 2291 7390 2307
rect 7460 2327 7504 2333
rect 7460 2307 7469 2327
rect 7489 2307 7504 2327
rect 7460 2291 7504 2307
rect 7554 2323 7603 2333
rect 7554 2303 7572 2323
rect 7592 2303 7603 2323
rect 7554 2291 7603 2303
rect 14815 2398 14864 2410
rect 14815 2378 14826 2398
rect 14846 2378 14864 2398
rect 14815 2368 14864 2378
rect 14914 2394 14958 2410
rect 14914 2374 14929 2394
rect 14949 2374 14958 2394
rect 14914 2368 14958 2374
rect 15028 2394 15072 2410
rect 15028 2374 15037 2394
rect 15057 2374 15072 2394
rect 15028 2368 15072 2374
rect 15122 2398 15171 2410
rect 15122 2378 15140 2398
rect 15160 2378 15171 2398
rect 15122 2368 15171 2378
rect 15236 2394 15280 2410
rect 15236 2374 15245 2394
rect 15265 2374 15280 2394
rect 15236 2368 15280 2374
rect 15330 2398 15379 2410
rect 15330 2378 15348 2398
rect 15368 2378 15379 2398
rect 15330 2368 15379 2378
rect 15449 2394 15493 2410
rect 15449 2374 15458 2394
rect 15478 2374 15493 2394
rect 15449 2368 15493 2374
rect 15543 2398 15592 2410
rect 15543 2378 15561 2398
rect 15581 2378 15592 2398
rect 15543 2368 15592 2378
rect 12206 2352 12255 2362
rect 12206 2332 12217 2352
rect 12237 2332 12255 2352
rect 12206 2320 12255 2332
rect 12305 2356 12349 2362
rect 12305 2336 12320 2356
rect 12340 2336 12349 2356
rect 12305 2320 12349 2336
rect 12419 2352 12468 2362
rect 12419 2332 12430 2352
rect 12450 2332 12468 2352
rect 12419 2320 12468 2332
rect 12518 2356 12562 2362
rect 12518 2336 12533 2356
rect 12553 2336 12562 2356
rect 12518 2320 12562 2336
rect 12627 2352 12676 2362
rect 12627 2332 12638 2352
rect 12658 2332 12676 2352
rect 12627 2320 12676 2332
rect 12726 2356 12770 2362
rect 12726 2336 12741 2356
rect 12761 2336 12770 2356
rect 12726 2320 12770 2336
rect 12840 2356 12884 2362
rect 12840 2336 12849 2356
rect 12869 2336 12884 2356
rect 12840 2320 12884 2336
rect 12934 2352 12983 2362
rect 12934 2332 12952 2352
rect 12972 2332 12983 2352
rect 12934 2320 12983 2332
rect 20096 2377 20145 2389
rect 20096 2357 20107 2377
rect 20127 2357 20145 2377
rect 20096 2347 20145 2357
rect 20195 2373 20239 2389
rect 20195 2353 20210 2373
rect 20230 2353 20239 2373
rect 20195 2347 20239 2353
rect 20309 2373 20353 2389
rect 20309 2353 20318 2373
rect 20338 2353 20353 2373
rect 20309 2347 20353 2353
rect 20403 2377 20452 2389
rect 20403 2357 20421 2377
rect 20441 2357 20452 2377
rect 20403 2347 20452 2357
rect 20517 2373 20561 2389
rect 20517 2353 20526 2373
rect 20546 2353 20561 2373
rect 20517 2347 20561 2353
rect 20611 2377 20660 2389
rect 20611 2357 20629 2377
rect 20649 2357 20660 2377
rect 20611 2347 20660 2357
rect 20730 2373 20774 2389
rect 20730 2353 20739 2373
rect 20759 2353 20774 2373
rect 20730 2347 20774 2353
rect 20824 2377 20873 2389
rect 20824 2357 20842 2377
rect 20862 2357 20873 2377
rect 20824 2347 20873 2357
rect 3141 2156 3190 2168
rect 3141 2136 3152 2156
rect 3172 2136 3190 2156
rect 3141 2126 3190 2136
rect 3240 2152 3284 2168
rect 3240 2132 3255 2152
rect 3275 2132 3284 2152
rect 3240 2126 3284 2132
rect 3354 2152 3398 2168
rect 3354 2132 3363 2152
rect 3383 2132 3398 2152
rect 3354 2126 3398 2132
rect 3448 2156 3497 2168
rect 3448 2136 3466 2156
rect 3486 2136 3497 2156
rect 3448 2126 3497 2136
rect 3562 2152 3606 2168
rect 3562 2132 3571 2152
rect 3591 2132 3606 2152
rect 3562 2126 3606 2132
rect 3656 2156 3705 2168
rect 3656 2136 3674 2156
rect 3694 2136 3705 2156
rect 3656 2126 3705 2136
rect 3775 2152 3819 2168
rect 3775 2132 3784 2152
rect 3804 2132 3819 2152
rect 3775 2126 3819 2132
rect 3869 2156 3918 2168
rect 3869 2136 3887 2156
rect 3907 2136 3918 2156
rect 3869 2126 3918 2136
rect 325 2058 374 2068
rect 325 2038 336 2058
rect 356 2038 374 2058
rect 325 2026 374 2038
rect 424 2062 468 2068
rect 424 2042 439 2062
rect 459 2042 468 2062
rect 424 2026 468 2042
rect 538 2058 587 2068
rect 538 2038 549 2058
rect 569 2038 587 2058
rect 538 2026 587 2038
rect 637 2062 681 2068
rect 637 2042 652 2062
rect 672 2042 681 2062
rect 637 2026 681 2042
rect 746 2058 795 2068
rect 746 2038 757 2058
rect 777 2038 795 2058
rect 746 2026 795 2038
rect 845 2062 889 2068
rect 845 2042 860 2062
rect 880 2042 889 2062
rect 845 2026 889 2042
rect 959 2062 1003 2068
rect 959 2042 968 2062
rect 988 2042 1003 2062
rect 959 2026 1003 2042
rect 1053 2058 1102 2068
rect 1053 2038 1071 2058
rect 1091 2038 1102 2058
rect 1053 2026 1102 2038
rect 8422 2135 8471 2147
rect 8422 2115 8433 2135
rect 8453 2115 8471 2135
rect 8422 2105 8471 2115
rect 8521 2131 8565 2147
rect 8521 2111 8536 2131
rect 8556 2111 8565 2131
rect 8521 2105 8565 2111
rect 8635 2131 8679 2147
rect 8635 2111 8644 2131
rect 8664 2111 8679 2131
rect 8635 2105 8679 2111
rect 8729 2135 8778 2147
rect 8729 2115 8747 2135
rect 8767 2115 8778 2135
rect 8729 2105 8778 2115
rect 8843 2131 8887 2147
rect 8843 2111 8852 2131
rect 8872 2111 8887 2131
rect 8843 2105 8887 2111
rect 8937 2135 8986 2147
rect 8937 2115 8955 2135
rect 8975 2115 8986 2135
rect 8937 2105 8986 2115
rect 9056 2131 9100 2147
rect 9056 2111 9065 2131
rect 9085 2111 9100 2131
rect 9056 2105 9100 2111
rect 9150 2135 9199 2147
rect 9150 2115 9168 2135
rect 9188 2115 9199 2135
rect 17487 2331 17536 2341
rect 17487 2311 17498 2331
rect 17518 2311 17536 2331
rect 17487 2299 17536 2311
rect 17586 2335 17630 2341
rect 17586 2315 17601 2335
rect 17621 2315 17630 2335
rect 17586 2299 17630 2315
rect 17700 2331 17749 2341
rect 17700 2311 17711 2331
rect 17731 2311 17749 2331
rect 17700 2299 17749 2311
rect 17799 2335 17843 2341
rect 17799 2315 17814 2335
rect 17834 2315 17843 2335
rect 17799 2299 17843 2315
rect 17908 2331 17957 2341
rect 17908 2311 17919 2331
rect 17939 2311 17957 2331
rect 17908 2299 17957 2311
rect 18007 2335 18051 2341
rect 18007 2315 18022 2335
rect 18042 2315 18051 2335
rect 18007 2299 18051 2315
rect 18121 2335 18165 2341
rect 18121 2315 18130 2335
rect 18150 2315 18165 2335
rect 18121 2299 18165 2315
rect 18215 2331 18264 2341
rect 18215 2311 18233 2331
rect 18253 2311 18264 2331
rect 18215 2299 18264 2311
rect 13802 2164 13851 2176
rect 9150 2105 9199 2115
rect 5606 2037 5655 2047
rect 5606 2017 5617 2037
rect 5637 2017 5655 2037
rect 5606 2005 5655 2017
rect 5705 2041 5749 2047
rect 5705 2021 5720 2041
rect 5740 2021 5749 2041
rect 5705 2005 5749 2021
rect 5819 2037 5868 2047
rect 5819 2017 5830 2037
rect 5850 2017 5868 2037
rect 5819 2005 5868 2017
rect 5918 2041 5962 2047
rect 5918 2021 5933 2041
rect 5953 2021 5962 2041
rect 5918 2005 5962 2021
rect 6027 2037 6076 2047
rect 6027 2017 6038 2037
rect 6058 2017 6076 2037
rect 6027 2005 6076 2017
rect 6126 2041 6170 2047
rect 6126 2021 6141 2041
rect 6161 2021 6170 2041
rect 6126 2005 6170 2021
rect 6240 2041 6284 2047
rect 6240 2021 6249 2041
rect 6269 2021 6284 2041
rect 6240 2005 6284 2021
rect 6334 2037 6383 2047
rect 6334 2017 6352 2037
rect 6372 2017 6383 2037
rect 6334 2005 6383 2017
rect 4153 1975 4202 1987
rect 4153 1955 4164 1975
rect 4184 1955 4202 1975
rect 4153 1945 4202 1955
rect 4252 1971 4296 1987
rect 4252 1951 4267 1971
rect 4287 1951 4296 1971
rect 4252 1945 4296 1951
rect 4366 1971 4410 1987
rect 4366 1951 4375 1971
rect 4395 1951 4410 1971
rect 4366 1945 4410 1951
rect 4460 1975 4509 1987
rect 4460 1955 4478 1975
rect 4498 1955 4509 1975
rect 4460 1945 4509 1955
rect 4574 1971 4618 1987
rect 4574 1951 4583 1971
rect 4603 1951 4618 1971
rect 4574 1945 4618 1951
rect 4668 1975 4717 1987
rect 4668 1955 4686 1975
rect 4706 1955 4717 1975
rect 4668 1945 4717 1955
rect 4787 1971 4831 1987
rect 4787 1951 4796 1971
rect 4816 1951 4831 1971
rect 4787 1945 4831 1951
rect 4881 1975 4930 1987
rect 4881 1955 4899 1975
rect 4919 1955 4930 1975
rect 4881 1945 4930 1955
rect 1337 1877 1386 1887
rect 1337 1857 1348 1877
rect 1368 1857 1386 1877
rect 1337 1845 1386 1857
rect 1436 1881 1480 1887
rect 1436 1861 1451 1881
rect 1471 1861 1480 1881
rect 1436 1845 1480 1861
rect 1550 1877 1599 1887
rect 1550 1857 1561 1877
rect 1581 1857 1599 1877
rect 1550 1845 1599 1857
rect 1649 1881 1693 1887
rect 1649 1861 1664 1881
rect 1684 1861 1693 1881
rect 1649 1845 1693 1861
rect 1758 1877 1807 1887
rect 1758 1857 1769 1877
rect 1789 1857 1807 1877
rect 1758 1845 1807 1857
rect 1857 1881 1901 1887
rect 1857 1861 1872 1881
rect 1892 1861 1901 1881
rect 1857 1845 1901 1861
rect 1971 1881 2015 1887
rect 1971 1861 1980 1881
rect 2000 1861 2015 1881
rect 1971 1845 2015 1861
rect 2065 1877 2114 1887
rect 2065 1857 2083 1877
rect 2103 1857 2114 1877
rect 13802 2144 13813 2164
rect 13833 2144 13851 2164
rect 13802 2134 13851 2144
rect 13901 2160 13945 2176
rect 13901 2140 13916 2160
rect 13936 2140 13945 2160
rect 13901 2134 13945 2140
rect 14015 2160 14059 2176
rect 14015 2140 14024 2160
rect 14044 2140 14059 2160
rect 14015 2134 14059 2140
rect 14109 2164 14158 2176
rect 14109 2144 14127 2164
rect 14147 2144 14158 2164
rect 14109 2134 14158 2144
rect 14223 2160 14267 2176
rect 14223 2140 14232 2160
rect 14252 2140 14267 2160
rect 14223 2134 14267 2140
rect 14317 2164 14366 2176
rect 14317 2144 14335 2164
rect 14355 2144 14366 2164
rect 14317 2134 14366 2144
rect 14436 2160 14480 2176
rect 14436 2140 14445 2160
rect 14465 2140 14480 2160
rect 14436 2134 14480 2140
rect 14530 2164 14579 2176
rect 14530 2144 14548 2164
rect 14568 2144 14579 2164
rect 14530 2134 14579 2144
rect 10986 2066 11035 2076
rect 10986 2046 10997 2066
rect 11017 2046 11035 2066
rect 10986 2034 11035 2046
rect 11085 2070 11129 2076
rect 11085 2050 11100 2070
rect 11120 2050 11129 2070
rect 11085 2034 11129 2050
rect 11199 2066 11248 2076
rect 11199 2046 11210 2066
rect 11230 2046 11248 2066
rect 11199 2034 11248 2046
rect 11298 2070 11342 2076
rect 11298 2050 11313 2070
rect 11333 2050 11342 2070
rect 11298 2034 11342 2050
rect 11407 2066 11456 2076
rect 11407 2046 11418 2066
rect 11438 2046 11456 2066
rect 11407 2034 11456 2046
rect 11506 2070 11550 2076
rect 11506 2050 11521 2070
rect 11541 2050 11550 2070
rect 11506 2034 11550 2050
rect 11620 2070 11664 2076
rect 11620 2050 11629 2070
rect 11649 2050 11664 2070
rect 11620 2034 11664 2050
rect 11714 2066 11763 2076
rect 11714 2046 11732 2066
rect 11752 2046 11763 2066
rect 11714 2034 11763 2046
rect 2065 1845 2114 1857
rect 19083 2143 19132 2155
rect 9434 1954 9483 1966
rect 9434 1934 9445 1954
rect 9465 1934 9483 1954
rect 9434 1924 9483 1934
rect 9533 1950 9577 1966
rect 9533 1930 9548 1950
rect 9568 1930 9577 1950
rect 9533 1924 9577 1930
rect 9647 1950 9691 1966
rect 9647 1930 9656 1950
rect 9676 1930 9691 1950
rect 9647 1924 9691 1930
rect 9741 1954 9790 1966
rect 9741 1934 9759 1954
rect 9779 1934 9790 1954
rect 9741 1924 9790 1934
rect 9855 1950 9899 1966
rect 9855 1930 9864 1950
rect 9884 1930 9899 1950
rect 9855 1924 9899 1930
rect 9949 1954 9998 1966
rect 9949 1934 9967 1954
rect 9987 1934 9998 1954
rect 9949 1924 9998 1934
rect 10068 1950 10112 1966
rect 10068 1930 10077 1950
rect 10097 1930 10112 1950
rect 10068 1924 10112 1930
rect 10162 1954 10211 1966
rect 10162 1934 10180 1954
rect 10200 1934 10211 1954
rect 10162 1924 10211 1934
rect 6618 1856 6667 1866
rect 6618 1836 6629 1856
rect 6649 1836 6667 1856
rect 6618 1824 6667 1836
rect 6717 1860 6761 1866
rect 6717 1840 6732 1860
rect 6752 1840 6761 1860
rect 6717 1824 6761 1840
rect 6831 1856 6880 1866
rect 6831 1836 6842 1856
rect 6862 1836 6880 1856
rect 6831 1824 6880 1836
rect 6930 1860 6974 1866
rect 6930 1840 6945 1860
rect 6965 1840 6974 1860
rect 6930 1824 6974 1840
rect 7039 1856 7088 1866
rect 7039 1836 7050 1856
rect 7070 1836 7088 1856
rect 7039 1824 7088 1836
rect 7138 1860 7182 1866
rect 7138 1840 7153 1860
rect 7173 1840 7182 1860
rect 7138 1824 7182 1840
rect 7252 1860 7296 1866
rect 7252 1840 7261 1860
rect 7281 1840 7296 1860
rect 7252 1824 7296 1840
rect 7346 1856 7395 1866
rect 7346 1836 7364 1856
rect 7384 1836 7395 1856
rect 19083 2123 19094 2143
rect 19114 2123 19132 2143
rect 19083 2113 19132 2123
rect 19182 2139 19226 2155
rect 19182 2119 19197 2139
rect 19217 2119 19226 2139
rect 19182 2113 19226 2119
rect 19296 2139 19340 2155
rect 19296 2119 19305 2139
rect 19325 2119 19340 2139
rect 19296 2113 19340 2119
rect 19390 2143 19439 2155
rect 19390 2123 19408 2143
rect 19428 2123 19439 2143
rect 19390 2113 19439 2123
rect 19504 2139 19548 2155
rect 19504 2119 19513 2139
rect 19533 2119 19548 2139
rect 19504 2113 19548 2119
rect 19598 2143 19647 2155
rect 19598 2123 19616 2143
rect 19636 2123 19647 2143
rect 19598 2113 19647 2123
rect 19717 2139 19761 2155
rect 19717 2119 19726 2139
rect 19746 2119 19761 2139
rect 19717 2113 19761 2119
rect 19811 2143 19860 2155
rect 19811 2123 19829 2143
rect 19849 2123 19860 2143
rect 19811 2113 19860 2123
rect 16267 2045 16316 2055
rect 16267 2025 16278 2045
rect 16298 2025 16316 2045
rect 16267 2013 16316 2025
rect 16366 2049 16410 2055
rect 16366 2029 16381 2049
rect 16401 2029 16410 2049
rect 16366 2013 16410 2029
rect 16480 2045 16529 2055
rect 16480 2025 16491 2045
rect 16511 2025 16529 2045
rect 16480 2013 16529 2025
rect 16579 2049 16623 2055
rect 16579 2029 16594 2049
rect 16614 2029 16623 2049
rect 16579 2013 16623 2029
rect 16688 2045 16737 2055
rect 16688 2025 16699 2045
rect 16719 2025 16737 2045
rect 16688 2013 16737 2025
rect 16787 2049 16831 2055
rect 16787 2029 16802 2049
rect 16822 2029 16831 2049
rect 16787 2013 16831 2029
rect 16901 2049 16945 2055
rect 16901 2029 16910 2049
rect 16930 2029 16945 2049
rect 16901 2013 16945 2029
rect 16995 2045 17044 2055
rect 16995 2025 17013 2045
rect 17033 2025 17044 2045
rect 16995 2013 17044 2025
rect 14814 1983 14863 1995
rect 14814 1963 14825 1983
rect 14845 1963 14863 1983
rect 14814 1953 14863 1963
rect 14913 1979 14957 1995
rect 14913 1959 14928 1979
rect 14948 1959 14957 1979
rect 14913 1953 14957 1959
rect 15027 1979 15071 1995
rect 15027 1959 15036 1979
rect 15056 1959 15071 1979
rect 15027 1953 15071 1959
rect 15121 1983 15170 1995
rect 15121 1963 15139 1983
rect 15159 1963 15170 1983
rect 15121 1953 15170 1963
rect 15235 1979 15279 1995
rect 15235 1959 15244 1979
rect 15264 1959 15279 1979
rect 15235 1953 15279 1959
rect 15329 1983 15378 1995
rect 15329 1963 15347 1983
rect 15367 1963 15378 1983
rect 15329 1953 15378 1963
rect 15448 1979 15492 1995
rect 15448 1959 15457 1979
rect 15477 1959 15492 1979
rect 15448 1953 15492 1959
rect 15542 1983 15591 1995
rect 15542 1963 15560 1983
rect 15580 1963 15591 1983
rect 15542 1953 15591 1963
rect 11998 1885 12047 1895
rect 7346 1824 7395 1836
rect 3091 1736 3140 1748
rect 3091 1716 3102 1736
rect 3122 1716 3140 1736
rect 3091 1706 3140 1716
rect 3190 1732 3234 1748
rect 3190 1712 3205 1732
rect 3225 1712 3234 1732
rect 3190 1706 3234 1712
rect 3304 1732 3348 1748
rect 3304 1712 3313 1732
rect 3333 1712 3348 1732
rect 3304 1706 3348 1712
rect 3398 1736 3447 1748
rect 3398 1716 3416 1736
rect 3436 1716 3447 1736
rect 3398 1706 3447 1716
rect 3512 1732 3556 1748
rect 3512 1712 3521 1732
rect 3541 1712 3556 1732
rect 3512 1706 3556 1712
rect 3606 1736 3655 1748
rect 3606 1716 3624 1736
rect 3644 1716 3655 1736
rect 3606 1706 3655 1716
rect 3725 1732 3769 1748
rect 3725 1712 3734 1732
rect 3754 1712 3769 1732
rect 3725 1706 3769 1712
rect 3819 1736 3868 1748
rect 3819 1716 3837 1736
rect 3857 1716 3868 1736
rect 3819 1706 3868 1716
rect 324 1643 373 1653
rect 324 1623 335 1643
rect 355 1623 373 1643
rect 324 1611 373 1623
rect 423 1647 467 1653
rect 423 1627 438 1647
rect 458 1627 467 1647
rect 423 1611 467 1627
rect 537 1643 586 1653
rect 537 1623 548 1643
rect 568 1623 586 1643
rect 537 1611 586 1623
rect 636 1647 680 1653
rect 636 1627 651 1647
rect 671 1627 680 1647
rect 636 1611 680 1627
rect 745 1643 794 1653
rect 745 1623 756 1643
rect 776 1623 794 1643
rect 745 1611 794 1623
rect 844 1647 888 1653
rect 844 1627 859 1647
rect 879 1627 888 1647
rect 844 1611 888 1627
rect 958 1647 1002 1653
rect 958 1627 967 1647
rect 987 1627 1002 1647
rect 958 1611 1002 1627
rect 1052 1643 1101 1653
rect 1052 1623 1070 1643
rect 1090 1623 1101 1643
rect 11998 1865 12009 1885
rect 12029 1865 12047 1885
rect 11998 1853 12047 1865
rect 12097 1889 12141 1895
rect 12097 1869 12112 1889
rect 12132 1869 12141 1889
rect 12097 1853 12141 1869
rect 12211 1885 12260 1895
rect 12211 1865 12222 1885
rect 12242 1865 12260 1885
rect 12211 1853 12260 1865
rect 12310 1889 12354 1895
rect 12310 1869 12325 1889
rect 12345 1869 12354 1889
rect 12310 1853 12354 1869
rect 12419 1885 12468 1895
rect 12419 1865 12430 1885
rect 12450 1865 12468 1885
rect 12419 1853 12468 1865
rect 12518 1889 12562 1895
rect 12518 1869 12533 1889
rect 12553 1869 12562 1889
rect 12518 1853 12562 1869
rect 12632 1889 12676 1895
rect 12632 1869 12641 1889
rect 12661 1869 12676 1889
rect 12632 1853 12676 1869
rect 12726 1885 12775 1895
rect 12726 1865 12744 1885
rect 12764 1865 12775 1885
rect 12726 1853 12775 1865
rect 20095 1962 20144 1974
rect 20095 1942 20106 1962
rect 20126 1942 20144 1962
rect 20095 1932 20144 1942
rect 20194 1958 20238 1974
rect 20194 1938 20209 1958
rect 20229 1938 20238 1958
rect 20194 1932 20238 1938
rect 20308 1958 20352 1974
rect 20308 1938 20317 1958
rect 20337 1938 20352 1958
rect 20308 1932 20352 1938
rect 20402 1962 20451 1974
rect 20402 1942 20420 1962
rect 20440 1942 20451 1962
rect 20402 1932 20451 1942
rect 20516 1958 20560 1974
rect 20516 1938 20525 1958
rect 20545 1938 20560 1958
rect 20516 1932 20560 1938
rect 20610 1962 20659 1974
rect 20610 1942 20628 1962
rect 20648 1942 20659 1962
rect 20610 1932 20659 1942
rect 20729 1958 20773 1974
rect 20729 1938 20738 1958
rect 20758 1938 20773 1958
rect 20729 1932 20773 1938
rect 20823 1962 20872 1974
rect 20823 1942 20841 1962
rect 20861 1942 20872 1962
rect 20823 1932 20872 1942
rect 17279 1864 17328 1874
rect 17279 1844 17290 1864
rect 17310 1844 17328 1864
rect 17279 1832 17328 1844
rect 17378 1868 17422 1874
rect 17378 1848 17393 1868
rect 17413 1848 17422 1868
rect 17378 1832 17422 1848
rect 17492 1864 17541 1874
rect 17492 1844 17503 1864
rect 17523 1844 17541 1864
rect 17492 1832 17541 1844
rect 17591 1868 17635 1874
rect 17591 1848 17606 1868
rect 17626 1848 17635 1868
rect 17591 1832 17635 1848
rect 17700 1864 17749 1874
rect 17700 1844 17711 1864
rect 17731 1844 17749 1864
rect 17700 1832 17749 1844
rect 17799 1868 17843 1874
rect 17799 1848 17814 1868
rect 17834 1848 17843 1868
rect 17799 1832 17843 1848
rect 17913 1868 17957 1874
rect 17913 1848 17922 1868
rect 17942 1848 17957 1868
rect 17913 1832 17957 1848
rect 18007 1864 18056 1874
rect 18007 1844 18025 1864
rect 18045 1844 18056 1864
rect 18007 1832 18056 1844
rect 13752 1744 13801 1756
rect 8372 1715 8421 1727
rect 1052 1611 1101 1623
rect 8372 1695 8383 1715
rect 8403 1695 8421 1715
rect 8372 1685 8421 1695
rect 8471 1711 8515 1727
rect 8471 1691 8486 1711
rect 8506 1691 8515 1711
rect 8471 1685 8515 1691
rect 8585 1711 8629 1727
rect 8585 1691 8594 1711
rect 8614 1691 8629 1711
rect 8585 1685 8629 1691
rect 8679 1715 8728 1727
rect 8679 1695 8697 1715
rect 8717 1695 8728 1715
rect 8679 1685 8728 1695
rect 8793 1711 8837 1727
rect 8793 1691 8802 1711
rect 8822 1691 8837 1711
rect 8793 1685 8837 1691
rect 8887 1715 8936 1727
rect 8887 1695 8905 1715
rect 8925 1695 8936 1715
rect 8887 1685 8936 1695
rect 9006 1711 9050 1727
rect 9006 1691 9015 1711
rect 9035 1691 9050 1711
rect 9006 1685 9050 1691
rect 9100 1715 9149 1727
rect 9100 1695 9118 1715
rect 9138 1695 9149 1715
rect 9100 1685 9149 1695
rect 5605 1622 5654 1632
rect 5605 1602 5616 1622
rect 5636 1602 5654 1622
rect 5605 1590 5654 1602
rect 5704 1626 5748 1632
rect 5704 1606 5719 1626
rect 5739 1606 5748 1626
rect 5704 1590 5748 1606
rect 5818 1622 5867 1632
rect 5818 1602 5829 1622
rect 5849 1602 5867 1622
rect 5818 1590 5867 1602
rect 5917 1626 5961 1632
rect 5917 1606 5932 1626
rect 5952 1606 5961 1626
rect 5917 1590 5961 1606
rect 6026 1622 6075 1632
rect 6026 1602 6037 1622
rect 6057 1602 6075 1622
rect 6026 1590 6075 1602
rect 6125 1626 6169 1632
rect 6125 1606 6140 1626
rect 6160 1606 6169 1626
rect 6125 1590 6169 1606
rect 6239 1626 6283 1632
rect 6239 1606 6248 1626
rect 6268 1606 6283 1626
rect 6239 1590 6283 1606
rect 6333 1622 6382 1632
rect 6333 1602 6351 1622
rect 6371 1602 6382 1622
rect 13752 1724 13763 1744
rect 13783 1724 13801 1744
rect 13752 1714 13801 1724
rect 13851 1740 13895 1756
rect 13851 1720 13866 1740
rect 13886 1720 13895 1740
rect 13851 1714 13895 1720
rect 13965 1740 14009 1756
rect 13965 1720 13974 1740
rect 13994 1720 14009 1740
rect 13965 1714 14009 1720
rect 14059 1744 14108 1756
rect 14059 1724 14077 1744
rect 14097 1724 14108 1744
rect 14059 1714 14108 1724
rect 14173 1740 14217 1756
rect 14173 1720 14182 1740
rect 14202 1720 14217 1740
rect 14173 1714 14217 1720
rect 14267 1744 14316 1756
rect 14267 1724 14285 1744
rect 14305 1724 14316 1744
rect 14267 1714 14316 1724
rect 14386 1740 14430 1756
rect 14386 1720 14395 1740
rect 14415 1720 14430 1740
rect 14386 1714 14430 1720
rect 14480 1744 14529 1756
rect 14480 1724 14498 1744
rect 14518 1724 14529 1744
rect 14480 1714 14529 1724
rect 6333 1590 6382 1602
rect 10985 1651 11034 1661
rect 10985 1631 10996 1651
rect 11016 1631 11034 1651
rect 10985 1619 11034 1631
rect 11084 1655 11128 1661
rect 11084 1635 11099 1655
rect 11119 1635 11128 1655
rect 11084 1619 11128 1635
rect 11198 1651 11247 1661
rect 11198 1631 11209 1651
rect 11229 1631 11247 1651
rect 11198 1619 11247 1631
rect 11297 1655 11341 1661
rect 11297 1635 11312 1655
rect 11332 1635 11341 1655
rect 11297 1619 11341 1635
rect 11406 1651 11455 1661
rect 11406 1631 11417 1651
rect 11437 1631 11455 1651
rect 11406 1619 11455 1631
rect 11505 1655 11549 1661
rect 11505 1635 11520 1655
rect 11540 1635 11549 1655
rect 11505 1619 11549 1635
rect 11619 1655 11663 1661
rect 11619 1635 11628 1655
rect 11648 1635 11663 1655
rect 11619 1619 11663 1635
rect 11713 1651 11762 1661
rect 11713 1631 11731 1651
rect 11751 1631 11762 1651
rect 19033 1723 19082 1735
rect 11713 1619 11762 1631
rect 19033 1703 19044 1723
rect 19064 1703 19082 1723
rect 19033 1693 19082 1703
rect 19132 1719 19176 1735
rect 19132 1699 19147 1719
rect 19167 1699 19176 1719
rect 19132 1693 19176 1699
rect 19246 1719 19290 1735
rect 19246 1699 19255 1719
rect 19275 1699 19290 1719
rect 19246 1693 19290 1699
rect 19340 1723 19389 1735
rect 19340 1703 19358 1723
rect 19378 1703 19389 1723
rect 19340 1693 19389 1703
rect 19454 1719 19498 1735
rect 19454 1699 19463 1719
rect 19483 1699 19498 1719
rect 19454 1693 19498 1699
rect 19548 1723 19597 1735
rect 19548 1703 19566 1723
rect 19586 1703 19597 1723
rect 19548 1693 19597 1703
rect 19667 1719 19711 1735
rect 19667 1699 19676 1719
rect 19696 1699 19711 1719
rect 19667 1693 19711 1699
rect 19761 1723 19810 1735
rect 19761 1703 19779 1723
rect 19799 1703 19810 1723
rect 19761 1693 19810 1703
rect 16266 1630 16315 1640
rect 16266 1610 16277 1630
rect 16297 1610 16315 1630
rect 16266 1598 16315 1610
rect 16365 1634 16409 1640
rect 16365 1614 16380 1634
rect 16400 1614 16409 1634
rect 16365 1598 16409 1614
rect 16479 1630 16528 1640
rect 16479 1610 16490 1630
rect 16510 1610 16528 1630
rect 16479 1598 16528 1610
rect 16578 1634 16622 1640
rect 16578 1614 16593 1634
rect 16613 1614 16622 1634
rect 16578 1598 16622 1614
rect 16687 1630 16736 1640
rect 16687 1610 16698 1630
rect 16718 1610 16736 1630
rect 16687 1598 16736 1610
rect 16786 1634 16830 1640
rect 16786 1614 16801 1634
rect 16821 1614 16830 1634
rect 16786 1598 16830 1614
rect 16900 1634 16944 1640
rect 16900 1614 16909 1634
rect 16929 1614 16944 1634
rect 16900 1598 16944 1614
rect 16994 1630 17043 1640
rect 16994 1610 17012 1630
rect 17032 1610 17043 1630
rect 16994 1598 17043 1610
rect 4159 1409 4208 1421
rect 4159 1389 4170 1409
rect 4190 1389 4208 1409
rect 4159 1379 4208 1389
rect 4258 1405 4302 1421
rect 4258 1385 4273 1405
rect 4293 1385 4302 1405
rect 4258 1379 4302 1385
rect 4372 1405 4416 1421
rect 4372 1385 4381 1405
rect 4401 1385 4416 1405
rect 4372 1379 4416 1385
rect 4466 1409 4515 1421
rect 4466 1389 4484 1409
rect 4504 1389 4515 1409
rect 4466 1379 4515 1389
rect 4580 1405 4624 1421
rect 4580 1385 4589 1405
rect 4609 1385 4624 1405
rect 4580 1379 4624 1385
rect 4674 1409 4723 1421
rect 4674 1389 4692 1409
rect 4712 1389 4723 1409
rect 4674 1379 4723 1389
rect 4793 1405 4837 1421
rect 4793 1385 4802 1405
rect 4822 1385 4837 1405
rect 4793 1379 4837 1385
rect 4887 1409 4936 1421
rect 4887 1389 4905 1409
rect 4925 1389 4936 1409
rect 4887 1379 4936 1389
rect 1392 1316 1441 1326
rect 1392 1296 1403 1316
rect 1423 1296 1441 1316
rect 1392 1284 1441 1296
rect 1491 1320 1535 1326
rect 1491 1300 1506 1320
rect 1526 1300 1535 1320
rect 1491 1284 1535 1300
rect 1605 1316 1654 1326
rect 1605 1296 1616 1316
rect 1636 1296 1654 1316
rect 1605 1284 1654 1296
rect 1704 1320 1748 1326
rect 1704 1300 1719 1320
rect 1739 1300 1748 1320
rect 1704 1284 1748 1300
rect 1813 1316 1862 1326
rect 1813 1296 1824 1316
rect 1844 1296 1862 1316
rect 1813 1284 1862 1296
rect 1912 1320 1956 1326
rect 1912 1300 1927 1320
rect 1947 1300 1956 1320
rect 1912 1284 1956 1300
rect 2026 1320 2070 1326
rect 2026 1300 2035 1320
rect 2055 1300 2070 1320
rect 2026 1284 2070 1300
rect 2120 1316 2169 1326
rect 2120 1296 2138 1316
rect 2158 1296 2169 1316
rect 9440 1388 9489 1400
rect 2120 1284 2169 1296
rect 9440 1368 9451 1388
rect 9471 1368 9489 1388
rect 9440 1358 9489 1368
rect 9539 1384 9583 1400
rect 9539 1364 9554 1384
rect 9574 1364 9583 1384
rect 9539 1358 9583 1364
rect 9653 1384 9697 1400
rect 9653 1364 9662 1384
rect 9682 1364 9697 1384
rect 9653 1358 9697 1364
rect 9747 1388 9796 1400
rect 9747 1368 9765 1388
rect 9785 1368 9796 1388
rect 9747 1358 9796 1368
rect 9861 1384 9905 1400
rect 9861 1364 9870 1384
rect 9890 1364 9905 1384
rect 9861 1358 9905 1364
rect 9955 1388 10004 1400
rect 9955 1368 9973 1388
rect 9993 1368 10004 1388
rect 9955 1358 10004 1368
rect 10074 1384 10118 1400
rect 10074 1364 10083 1384
rect 10103 1364 10118 1384
rect 10074 1358 10118 1364
rect 10168 1388 10217 1400
rect 10168 1368 10186 1388
rect 10206 1368 10217 1388
rect 10168 1358 10217 1368
rect 14820 1417 14869 1429
rect 6673 1295 6722 1305
rect 6673 1275 6684 1295
rect 6704 1275 6722 1295
rect 6673 1263 6722 1275
rect 6772 1299 6816 1305
rect 6772 1279 6787 1299
rect 6807 1279 6816 1299
rect 6772 1263 6816 1279
rect 6886 1295 6935 1305
rect 6886 1275 6897 1295
rect 6917 1275 6935 1295
rect 6886 1263 6935 1275
rect 6985 1299 7029 1305
rect 6985 1279 7000 1299
rect 7020 1279 7029 1299
rect 6985 1263 7029 1279
rect 7094 1295 7143 1305
rect 7094 1275 7105 1295
rect 7125 1275 7143 1295
rect 7094 1263 7143 1275
rect 7193 1299 7237 1305
rect 7193 1279 7208 1299
rect 7228 1279 7237 1299
rect 7193 1263 7237 1279
rect 7307 1299 7351 1305
rect 7307 1279 7316 1299
rect 7336 1279 7351 1299
rect 7307 1263 7351 1279
rect 7401 1295 7450 1305
rect 7401 1275 7419 1295
rect 7439 1275 7450 1295
rect 14820 1397 14831 1417
rect 14851 1397 14869 1417
rect 14820 1387 14869 1397
rect 14919 1413 14963 1429
rect 14919 1393 14934 1413
rect 14954 1393 14963 1413
rect 14919 1387 14963 1393
rect 15033 1413 15077 1429
rect 15033 1393 15042 1413
rect 15062 1393 15077 1413
rect 15033 1387 15077 1393
rect 15127 1417 15176 1429
rect 15127 1397 15145 1417
rect 15165 1397 15176 1417
rect 15127 1387 15176 1397
rect 15241 1413 15285 1429
rect 15241 1393 15250 1413
rect 15270 1393 15285 1413
rect 15241 1387 15285 1393
rect 15335 1417 15384 1429
rect 15335 1397 15353 1417
rect 15373 1397 15384 1417
rect 15335 1387 15384 1397
rect 15454 1413 15498 1429
rect 15454 1393 15463 1413
rect 15483 1393 15498 1413
rect 15454 1387 15498 1393
rect 15548 1417 15597 1429
rect 15548 1397 15566 1417
rect 15586 1397 15597 1417
rect 15548 1387 15597 1397
rect 12053 1324 12102 1334
rect 12053 1304 12064 1324
rect 12084 1304 12102 1324
rect 12053 1292 12102 1304
rect 12152 1328 12196 1334
rect 12152 1308 12167 1328
rect 12187 1308 12196 1328
rect 12152 1292 12196 1308
rect 12266 1324 12315 1334
rect 12266 1304 12277 1324
rect 12297 1304 12315 1324
rect 12266 1292 12315 1304
rect 12365 1328 12409 1334
rect 12365 1308 12380 1328
rect 12400 1308 12409 1328
rect 12365 1292 12409 1308
rect 12474 1324 12523 1334
rect 12474 1304 12485 1324
rect 12505 1304 12523 1324
rect 12474 1292 12523 1304
rect 12573 1328 12617 1334
rect 12573 1308 12588 1328
rect 12608 1308 12617 1328
rect 12573 1292 12617 1308
rect 12687 1328 12731 1334
rect 12687 1308 12696 1328
rect 12716 1308 12731 1328
rect 12687 1292 12731 1308
rect 12781 1324 12830 1334
rect 12781 1304 12799 1324
rect 12819 1304 12830 1324
rect 20101 1396 20150 1408
rect 12781 1292 12830 1304
rect 7401 1263 7450 1275
rect 3146 1175 3195 1187
rect 3146 1155 3157 1175
rect 3177 1155 3195 1175
rect 3146 1145 3195 1155
rect 3245 1171 3289 1187
rect 3245 1151 3260 1171
rect 3280 1151 3289 1171
rect 3245 1145 3289 1151
rect 3359 1171 3403 1187
rect 3359 1151 3368 1171
rect 3388 1151 3403 1171
rect 3359 1145 3403 1151
rect 3453 1175 3502 1187
rect 3453 1155 3471 1175
rect 3491 1155 3502 1175
rect 3453 1145 3502 1155
rect 3567 1171 3611 1187
rect 3567 1151 3576 1171
rect 3596 1151 3611 1171
rect 3567 1145 3611 1151
rect 3661 1175 3710 1187
rect 3661 1155 3679 1175
rect 3699 1155 3710 1175
rect 3661 1145 3710 1155
rect 3780 1171 3824 1187
rect 3780 1151 3789 1171
rect 3809 1151 3824 1171
rect 3780 1145 3824 1151
rect 3874 1175 3923 1187
rect 3874 1155 3892 1175
rect 3912 1155 3923 1175
rect 3874 1145 3923 1155
rect 330 1077 379 1087
rect 330 1057 341 1077
rect 361 1057 379 1077
rect 330 1045 379 1057
rect 429 1081 473 1087
rect 429 1061 444 1081
rect 464 1061 473 1081
rect 429 1045 473 1061
rect 543 1077 592 1087
rect 543 1057 554 1077
rect 574 1057 592 1077
rect 543 1045 592 1057
rect 642 1081 686 1087
rect 642 1061 657 1081
rect 677 1061 686 1081
rect 642 1045 686 1061
rect 751 1077 800 1087
rect 751 1057 762 1077
rect 782 1057 800 1077
rect 751 1045 800 1057
rect 850 1081 894 1087
rect 850 1061 865 1081
rect 885 1061 894 1081
rect 850 1045 894 1061
rect 964 1081 1008 1087
rect 964 1061 973 1081
rect 993 1061 1008 1081
rect 964 1045 1008 1061
rect 1058 1077 1107 1087
rect 1058 1057 1076 1077
rect 1096 1057 1107 1077
rect 1058 1045 1107 1057
rect 8427 1154 8476 1166
rect 8427 1134 8438 1154
rect 8458 1134 8476 1154
rect 8427 1124 8476 1134
rect 8526 1150 8570 1166
rect 8526 1130 8541 1150
rect 8561 1130 8570 1150
rect 8526 1124 8570 1130
rect 8640 1150 8684 1166
rect 8640 1130 8649 1150
rect 8669 1130 8684 1150
rect 8640 1124 8684 1130
rect 8734 1154 8783 1166
rect 8734 1134 8752 1154
rect 8772 1134 8783 1154
rect 8734 1124 8783 1134
rect 8848 1150 8892 1166
rect 8848 1130 8857 1150
rect 8877 1130 8892 1150
rect 8848 1124 8892 1130
rect 8942 1154 8991 1166
rect 8942 1134 8960 1154
rect 8980 1134 8991 1154
rect 8942 1124 8991 1134
rect 9061 1150 9105 1166
rect 9061 1130 9070 1150
rect 9090 1130 9105 1150
rect 9061 1124 9105 1130
rect 9155 1154 9204 1166
rect 9155 1134 9173 1154
rect 9193 1134 9204 1154
rect 20101 1376 20112 1396
rect 20132 1376 20150 1396
rect 20101 1366 20150 1376
rect 20200 1392 20244 1408
rect 20200 1372 20215 1392
rect 20235 1372 20244 1392
rect 20200 1366 20244 1372
rect 20314 1392 20358 1408
rect 20314 1372 20323 1392
rect 20343 1372 20358 1392
rect 20314 1366 20358 1372
rect 20408 1396 20457 1408
rect 20408 1376 20426 1396
rect 20446 1376 20457 1396
rect 20408 1366 20457 1376
rect 20522 1392 20566 1408
rect 20522 1372 20531 1392
rect 20551 1372 20566 1392
rect 20522 1366 20566 1372
rect 20616 1396 20665 1408
rect 20616 1376 20634 1396
rect 20654 1376 20665 1396
rect 20616 1366 20665 1376
rect 20735 1392 20779 1408
rect 20735 1372 20744 1392
rect 20764 1372 20779 1392
rect 20735 1366 20779 1372
rect 20829 1396 20878 1408
rect 20829 1376 20847 1396
rect 20867 1376 20878 1396
rect 20829 1366 20878 1376
rect 17334 1303 17383 1313
rect 17334 1283 17345 1303
rect 17365 1283 17383 1303
rect 17334 1271 17383 1283
rect 17433 1307 17477 1313
rect 17433 1287 17448 1307
rect 17468 1287 17477 1307
rect 17433 1271 17477 1287
rect 17547 1303 17596 1313
rect 17547 1283 17558 1303
rect 17578 1283 17596 1303
rect 17547 1271 17596 1283
rect 17646 1307 17690 1313
rect 17646 1287 17661 1307
rect 17681 1287 17690 1307
rect 17646 1271 17690 1287
rect 17755 1303 17804 1313
rect 17755 1283 17766 1303
rect 17786 1283 17804 1303
rect 17755 1271 17804 1283
rect 17854 1307 17898 1313
rect 17854 1287 17869 1307
rect 17889 1287 17898 1307
rect 17854 1271 17898 1287
rect 17968 1307 18012 1313
rect 17968 1287 17977 1307
rect 17997 1287 18012 1307
rect 17968 1271 18012 1287
rect 18062 1303 18111 1313
rect 18062 1283 18080 1303
rect 18100 1283 18111 1303
rect 18062 1271 18111 1283
rect 13807 1183 13856 1195
rect 9155 1124 9204 1134
rect 5611 1056 5660 1066
rect 5611 1036 5622 1056
rect 5642 1036 5660 1056
rect 5611 1024 5660 1036
rect 5710 1060 5754 1066
rect 5710 1040 5725 1060
rect 5745 1040 5754 1060
rect 5710 1024 5754 1040
rect 5824 1056 5873 1066
rect 5824 1036 5835 1056
rect 5855 1036 5873 1056
rect 5824 1024 5873 1036
rect 5923 1060 5967 1066
rect 5923 1040 5938 1060
rect 5958 1040 5967 1060
rect 5923 1024 5967 1040
rect 6032 1056 6081 1066
rect 6032 1036 6043 1056
rect 6063 1036 6081 1056
rect 6032 1024 6081 1036
rect 6131 1060 6175 1066
rect 6131 1040 6146 1060
rect 6166 1040 6175 1060
rect 6131 1024 6175 1040
rect 6245 1060 6289 1066
rect 6245 1040 6254 1060
rect 6274 1040 6289 1060
rect 6245 1024 6289 1040
rect 6339 1056 6388 1066
rect 6339 1036 6357 1056
rect 6377 1036 6388 1056
rect 6339 1024 6388 1036
rect 4158 994 4207 1006
rect 4158 974 4169 994
rect 4189 974 4207 994
rect 4158 964 4207 974
rect 4257 990 4301 1006
rect 4257 970 4272 990
rect 4292 970 4301 990
rect 4257 964 4301 970
rect 4371 990 4415 1006
rect 4371 970 4380 990
rect 4400 970 4415 990
rect 4371 964 4415 970
rect 4465 994 4514 1006
rect 4465 974 4483 994
rect 4503 974 4514 994
rect 4465 964 4514 974
rect 4579 990 4623 1006
rect 4579 970 4588 990
rect 4608 970 4623 990
rect 4579 964 4623 970
rect 4673 994 4722 1006
rect 4673 974 4691 994
rect 4711 974 4722 994
rect 4673 964 4722 974
rect 4792 990 4836 1006
rect 4792 970 4801 990
rect 4821 970 4836 990
rect 4792 964 4836 970
rect 4886 994 4935 1006
rect 4886 974 4904 994
rect 4924 974 4935 994
rect 4886 964 4935 974
rect 1342 896 1391 906
rect 1342 876 1353 896
rect 1373 876 1391 896
rect 1342 864 1391 876
rect 1441 900 1485 906
rect 1441 880 1456 900
rect 1476 880 1485 900
rect 1441 864 1485 880
rect 1555 896 1604 906
rect 1555 876 1566 896
rect 1586 876 1604 896
rect 1555 864 1604 876
rect 1654 900 1698 906
rect 1654 880 1669 900
rect 1689 880 1698 900
rect 1654 864 1698 880
rect 1763 896 1812 906
rect 1763 876 1774 896
rect 1794 876 1812 896
rect 1763 864 1812 876
rect 1862 900 1906 906
rect 1862 880 1877 900
rect 1897 880 1906 900
rect 1862 864 1906 880
rect 1976 900 2020 906
rect 1976 880 1985 900
rect 2005 880 2020 900
rect 1976 864 2020 880
rect 2070 896 2119 906
rect 2070 876 2088 896
rect 2108 876 2119 896
rect 13807 1163 13818 1183
rect 13838 1163 13856 1183
rect 13807 1153 13856 1163
rect 13906 1179 13950 1195
rect 13906 1159 13921 1179
rect 13941 1159 13950 1179
rect 13906 1153 13950 1159
rect 14020 1179 14064 1195
rect 14020 1159 14029 1179
rect 14049 1159 14064 1179
rect 14020 1153 14064 1159
rect 14114 1183 14163 1195
rect 14114 1163 14132 1183
rect 14152 1163 14163 1183
rect 14114 1153 14163 1163
rect 14228 1179 14272 1195
rect 14228 1159 14237 1179
rect 14257 1159 14272 1179
rect 14228 1153 14272 1159
rect 14322 1183 14371 1195
rect 14322 1163 14340 1183
rect 14360 1163 14371 1183
rect 14322 1153 14371 1163
rect 14441 1179 14485 1195
rect 14441 1159 14450 1179
rect 14470 1159 14485 1179
rect 14441 1153 14485 1159
rect 14535 1183 14584 1195
rect 14535 1163 14553 1183
rect 14573 1163 14584 1183
rect 14535 1153 14584 1163
rect 10991 1085 11040 1095
rect 10991 1065 11002 1085
rect 11022 1065 11040 1085
rect 10991 1053 11040 1065
rect 11090 1089 11134 1095
rect 11090 1069 11105 1089
rect 11125 1069 11134 1089
rect 11090 1053 11134 1069
rect 11204 1085 11253 1095
rect 11204 1065 11215 1085
rect 11235 1065 11253 1085
rect 11204 1053 11253 1065
rect 11303 1089 11347 1095
rect 11303 1069 11318 1089
rect 11338 1069 11347 1089
rect 11303 1053 11347 1069
rect 11412 1085 11461 1095
rect 11412 1065 11423 1085
rect 11443 1065 11461 1085
rect 11412 1053 11461 1065
rect 11511 1089 11555 1095
rect 11511 1069 11526 1089
rect 11546 1069 11555 1089
rect 11511 1053 11555 1069
rect 11625 1089 11669 1095
rect 11625 1069 11634 1089
rect 11654 1069 11669 1089
rect 11625 1053 11669 1069
rect 11719 1085 11768 1095
rect 11719 1065 11737 1085
rect 11757 1065 11768 1085
rect 11719 1053 11768 1065
rect 2070 864 2119 876
rect 19088 1162 19137 1174
rect 9439 973 9488 985
rect 9439 953 9450 973
rect 9470 953 9488 973
rect 9439 943 9488 953
rect 9538 969 9582 985
rect 9538 949 9553 969
rect 9573 949 9582 969
rect 9538 943 9582 949
rect 9652 969 9696 985
rect 9652 949 9661 969
rect 9681 949 9696 969
rect 9652 943 9696 949
rect 9746 973 9795 985
rect 9746 953 9764 973
rect 9784 953 9795 973
rect 9746 943 9795 953
rect 9860 969 9904 985
rect 9860 949 9869 969
rect 9889 949 9904 969
rect 9860 943 9904 949
rect 9954 973 10003 985
rect 9954 953 9972 973
rect 9992 953 10003 973
rect 9954 943 10003 953
rect 10073 969 10117 985
rect 10073 949 10082 969
rect 10102 949 10117 969
rect 10073 943 10117 949
rect 10167 973 10216 985
rect 10167 953 10185 973
rect 10205 953 10216 973
rect 10167 943 10216 953
rect 6623 875 6672 885
rect 6623 855 6634 875
rect 6654 855 6672 875
rect 6623 843 6672 855
rect 6722 879 6766 885
rect 6722 859 6737 879
rect 6757 859 6766 879
rect 6722 843 6766 859
rect 6836 875 6885 885
rect 6836 855 6847 875
rect 6867 855 6885 875
rect 6836 843 6885 855
rect 6935 879 6979 885
rect 6935 859 6950 879
rect 6970 859 6979 879
rect 6935 843 6979 859
rect 7044 875 7093 885
rect 7044 855 7055 875
rect 7075 855 7093 875
rect 7044 843 7093 855
rect 7143 879 7187 885
rect 7143 859 7158 879
rect 7178 859 7187 879
rect 7143 843 7187 859
rect 7257 879 7301 885
rect 7257 859 7266 879
rect 7286 859 7301 879
rect 7257 843 7301 859
rect 7351 875 7400 885
rect 7351 855 7369 875
rect 7389 855 7400 875
rect 19088 1142 19099 1162
rect 19119 1142 19137 1162
rect 19088 1132 19137 1142
rect 19187 1158 19231 1174
rect 19187 1138 19202 1158
rect 19222 1138 19231 1158
rect 19187 1132 19231 1138
rect 19301 1158 19345 1174
rect 19301 1138 19310 1158
rect 19330 1138 19345 1158
rect 19301 1132 19345 1138
rect 19395 1162 19444 1174
rect 19395 1142 19413 1162
rect 19433 1142 19444 1162
rect 19395 1132 19444 1142
rect 19509 1158 19553 1174
rect 19509 1138 19518 1158
rect 19538 1138 19553 1158
rect 19509 1132 19553 1138
rect 19603 1162 19652 1174
rect 19603 1142 19621 1162
rect 19641 1142 19652 1162
rect 19603 1132 19652 1142
rect 19722 1158 19766 1174
rect 19722 1138 19731 1158
rect 19751 1138 19766 1158
rect 19722 1132 19766 1138
rect 19816 1162 19865 1174
rect 19816 1142 19834 1162
rect 19854 1142 19865 1162
rect 19816 1132 19865 1142
rect 16272 1064 16321 1074
rect 16272 1044 16283 1064
rect 16303 1044 16321 1064
rect 16272 1032 16321 1044
rect 16371 1068 16415 1074
rect 16371 1048 16386 1068
rect 16406 1048 16415 1068
rect 16371 1032 16415 1048
rect 16485 1064 16534 1074
rect 16485 1044 16496 1064
rect 16516 1044 16534 1064
rect 16485 1032 16534 1044
rect 16584 1068 16628 1074
rect 16584 1048 16599 1068
rect 16619 1048 16628 1068
rect 16584 1032 16628 1048
rect 16693 1064 16742 1074
rect 16693 1044 16704 1064
rect 16724 1044 16742 1064
rect 16693 1032 16742 1044
rect 16792 1068 16836 1074
rect 16792 1048 16807 1068
rect 16827 1048 16836 1068
rect 16792 1032 16836 1048
rect 16906 1068 16950 1074
rect 16906 1048 16915 1068
rect 16935 1048 16950 1068
rect 16906 1032 16950 1048
rect 17000 1064 17049 1074
rect 17000 1044 17018 1064
rect 17038 1044 17049 1064
rect 17000 1032 17049 1044
rect 14819 1002 14868 1014
rect 14819 982 14830 1002
rect 14850 982 14868 1002
rect 14819 972 14868 982
rect 14918 998 14962 1014
rect 14918 978 14933 998
rect 14953 978 14962 998
rect 14918 972 14962 978
rect 15032 998 15076 1014
rect 15032 978 15041 998
rect 15061 978 15076 998
rect 15032 972 15076 978
rect 15126 1002 15175 1014
rect 15126 982 15144 1002
rect 15164 982 15175 1002
rect 15126 972 15175 982
rect 15240 998 15284 1014
rect 15240 978 15249 998
rect 15269 978 15284 998
rect 15240 972 15284 978
rect 15334 1002 15383 1014
rect 15334 982 15352 1002
rect 15372 982 15383 1002
rect 15334 972 15383 982
rect 15453 998 15497 1014
rect 15453 978 15462 998
rect 15482 978 15497 998
rect 15453 972 15497 978
rect 15547 1002 15596 1014
rect 15547 982 15565 1002
rect 15585 982 15596 1002
rect 15547 972 15596 982
rect 12003 904 12052 914
rect 7351 843 7400 855
rect 12003 884 12014 904
rect 12034 884 12052 904
rect 12003 872 12052 884
rect 12102 908 12146 914
rect 12102 888 12117 908
rect 12137 888 12146 908
rect 12102 872 12146 888
rect 12216 904 12265 914
rect 12216 884 12227 904
rect 12247 884 12265 904
rect 12216 872 12265 884
rect 12315 908 12359 914
rect 12315 888 12330 908
rect 12350 888 12359 908
rect 12315 872 12359 888
rect 12424 904 12473 914
rect 12424 884 12435 904
rect 12455 884 12473 904
rect 12424 872 12473 884
rect 12523 908 12567 914
rect 12523 888 12538 908
rect 12558 888 12567 908
rect 12523 872 12567 888
rect 12637 908 12681 914
rect 12637 888 12646 908
rect 12666 888 12681 908
rect 12637 872 12681 888
rect 12731 904 12780 914
rect 12731 884 12749 904
rect 12769 884 12780 904
rect 12731 872 12780 884
rect 20100 981 20149 993
rect 20100 961 20111 981
rect 20131 961 20149 981
rect 20100 951 20149 961
rect 20199 977 20243 993
rect 20199 957 20214 977
rect 20234 957 20243 977
rect 20199 951 20243 957
rect 20313 977 20357 993
rect 20313 957 20322 977
rect 20342 957 20357 977
rect 20313 951 20357 957
rect 20407 981 20456 993
rect 20407 961 20425 981
rect 20445 961 20456 981
rect 20407 951 20456 961
rect 20521 977 20565 993
rect 20521 957 20530 977
rect 20550 957 20565 977
rect 20521 951 20565 957
rect 20615 981 20664 993
rect 20615 961 20633 981
rect 20653 961 20664 981
rect 20615 951 20664 961
rect 20734 977 20778 993
rect 20734 957 20743 977
rect 20763 957 20778 977
rect 20734 951 20778 957
rect 20828 981 20877 993
rect 20828 961 20846 981
rect 20866 961 20877 981
rect 20828 951 20877 961
rect 17284 883 17333 893
rect 17284 863 17295 883
rect 17315 863 17333 883
rect 17284 851 17333 863
rect 17383 887 17427 893
rect 17383 867 17398 887
rect 17418 867 17427 887
rect 17383 851 17427 867
rect 17497 883 17546 893
rect 17497 863 17508 883
rect 17528 863 17546 883
rect 17497 851 17546 863
rect 17596 887 17640 893
rect 17596 867 17611 887
rect 17631 867 17640 887
rect 17596 851 17640 867
rect 17705 883 17754 893
rect 17705 863 17716 883
rect 17736 863 17754 883
rect 17705 851 17754 863
rect 17804 887 17848 893
rect 17804 867 17819 887
rect 17839 867 17848 887
rect 17804 851 17848 867
rect 17918 887 17962 893
rect 17918 867 17927 887
rect 17947 867 17962 887
rect 17918 851 17962 867
rect 18012 883 18061 893
rect 18012 863 18030 883
rect 18050 863 18061 883
rect 18012 851 18061 863
rect 329 662 378 672
rect 329 642 340 662
rect 360 642 378 662
rect 329 630 378 642
rect 428 666 472 672
rect 428 646 443 666
rect 463 646 472 666
rect 428 630 472 646
rect 542 662 591 672
rect 542 642 553 662
rect 573 642 591 662
rect 542 630 591 642
rect 641 666 685 672
rect 641 646 656 666
rect 676 646 685 666
rect 641 630 685 646
rect 750 662 799 672
rect 750 642 761 662
rect 781 642 799 662
rect 750 630 799 642
rect 849 666 893 672
rect 849 646 864 666
rect 884 646 893 666
rect 849 630 893 646
rect 963 666 1007 672
rect 963 646 972 666
rect 992 646 1007 666
rect 963 630 1007 646
rect 1057 662 1106 672
rect 1057 642 1075 662
rect 1095 642 1106 662
rect 1057 630 1106 642
rect 5610 641 5659 651
rect 5610 621 5621 641
rect 5641 621 5659 641
rect 5610 609 5659 621
rect 5709 645 5753 651
rect 5709 625 5724 645
rect 5744 625 5753 645
rect 5709 609 5753 625
rect 5823 641 5872 651
rect 5823 621 5834 641
rect 5854 621 5872 641
rect 5823 609 5872 621
rect 5922 645 5966 651
rect 5922 625 5937 645
rect 5957 625 5966 645
rect 5922 609 5966 625
rect 6031 641 6080 651
rect 6031 621 6042 641
rect 6062 621 6080 641
rect 6031 609 6080 621
rect 6130 645 6174 651
rect 6130 625 6145 645
rect 6165 625 6174 645
rect 6130 609 6174 625
rect 6244 645 6288 651
rect 6244 625 6253 645
rect 6273 625 6288 645
rect 6244 609 6288 625
rect 6338 641 6387 651
rect 6338 621 6356 641
rect 6376 621 6387 641
rect 6338 609 6387 621
rect 10990 670 11039 680
rect 10990 650 11001 670
rect 11021 650 11039 670
rect 10990 638 11039 650
rect 11089 674 11133 680
rect 11089 654 11104 674
rect 11124 654 11133 674
rect 11089 638 11133 654
rect 11203 670 11252 680
rect 11203 650 11214 670
rect 11234 650 11252 670
rect 11203 638 11252 650
rect 11302 674 11346 680
rect 11302 654 11317 674
rect 11337 654 11346 674
rect 11302 638 11346 654
rect 11411 670 11460 680
rect 11411 650 11422 670
rect 11442 650 11460 670
rect 11411 638 11460 650
rect 11510 674 11554 680
rect 11510 654 11525 674
rect 11545 654 11554 674
rect 11510 638 11554 654
rect 11624 674 11668 680
rect 11624 654 11633 674
rect 11653 654 11668 674
rect 11624 638 11668 654
rect 11718 670 11767 680
rect 11718 650 11736 670
rect 11756 650 11767 670
rect 11718 638 11767 650
rect 16271 649 16320 659
rect 16271 629 16282 649
rect 16302 629 16320 649
rect 16271 617 16320 629
rect 16370 653 16414 659
rect 16370 633 16385 653
rect 16405 633 16414 653
rect 16370 617 16414 633
rect 16484 649 16533 659
rect 16484 629 16495 649
rect 16515 629 16533 649
rect 16484 617 16533 629
rect 16583 653 16627 659
rect 16583 633 16598 653
rect 16618 633 16627 653
rect 16583 617 16627 633
rect 16692 649 16741 659
rect 16692 629 16703 649
rect 16723 629 16741 649
rect 16692 617 16741 629
rect 16791 653 16835 659
rect 16791 633 16806 653
rect 16826 633 16835 653
rect 16791 617 16835 633
rect 16905 653 16949 659
rect 16905 633 16914 653
rect 16934 633 16949 653
rect 16905 617 16949 633
rect 16999 649 17048 659
rect 16999 629 17017 649
rect 17037 629 17048 649
rect 16999 617 17048 629
rect 1732 181 1781 191
rect 1732 161 1743 181
rect 1763 161 1781 181
rect 1732 149 1781 161
rect 1831 185 1875 191
rect 1831 165 1846 185
rect 1866 165 1875 185
rect 1831 149 1875 165
rect 1945 181 1994 191
rect 1945 161 1956 181
rect 1976 161 1994 181
rect 1945 149 1994 161
rect 2044 185 2088 191
rect 2044 165 2059 185
rect 2079 165 2088 185
rect 2044 149 2088 165
rect 2153 181 2202 191
rect 2153 161 2164 181
rect 2184 161 2202 181
rect 2153 149 2202 161
rect 2252 185 2296 191
rect 2252 165 2267 185
rect 2287 165 2296 185
rect 2252 149 2296 165
rect 2366 185 2410 191
rect 2366 165 2375 185
rect 2395 165 2410 185
rect 2366 149 2410 165
rect 2460 181 2509 191
rect 2460 161 2478 181
rect 2498 161 2509 181
rect 2460 149 2509 161
rect 12393 189 12442 199
rect 7013 160 7062 170
rect 7013 140 7024 160
rect 7044 140 7062 160
rect 7013 128 7062 140
rect 7112 164 7156 170
rect 7112 144 7127 164
rect 7147 144 7156 164
rect 7112 128 7156 144
rect 7226 160 7275 170
rect 7226 140 7237 160
rect 7257 140 7275 160
rect 7226 128 7275 140
rect 7325 164 7369 170
rect 7325 144 7340 164
rect 7360 144 7369 164
rect 7325 128 7369 144
rect 7434 160 7483 170
rect 7434 140 7445 160
rect 7465 140 7483 160
rect 7434 128 7483 140
rect 7533 164 7577 170
rect 7533 144 7548 164
rect 7568 144 7577 164
rect 7533 128 7577 144
rect 7647 164 7691 170
rect 7647 144 7656 164
rect 7676 144 7691 164
rect 7647 128 7691 144
rect 7741 160 7790 170
rect 7741 140 7759 160
rect 7779 140 7790 160
rect 7741 128 7790 140
rect 4822 93 4871 103
rect 4822 73 4833 93
rect 4853 73 4871 93
rect 4822 61 4871 73
rect 4921 97 4965 103
rect 4921 77 4936 97
rect 4956 77 4965 97
rect 4921 61 4965 77
rect 5035 93 5084 103
rect 5035 73 5046 93
rect 5066 73 5084 93
rect 5035 61 5084 73
rect 5134 97 5178 103
rect 5134 77 5149 97
rect 5169 77 5178 97
rect 5134 61 5178 77
rect 5243 93 5292 103
rect 5243 73 5254 93
rect 5274 73 5292 93
rect 5243 61 5292 73
rect 5342 97 5386 103
rect 5342 77 5357 97
rect 5377 77 5386 97
rect 5342 61 5386 77
rect 5456 97 5500 103
rect 5456 77 5465 97
rect 5485 77 5500 97
rect 5456 61 5500 77
rect 5550 93 5599 103
rect 12393 169 12404 189
rect 12424 169 12442 189
rect 12393 157 12442 169
rect 12492 193 12536 199
rect 12492 173 12507 193
rect 12527 173 12536 193
rect 12492 157 12536 173
rect 12606 189 12655 199
rect 12606 169 12617 189
rect 12637 169 12655 189
rect 12606 157 12655 169
rect 12705 193 12749 199
rect 12705 173 12720 193
rect 12740 173 12749 193
rect 12705 157 12749 173
rect 12814 189 12863 199
rect 12814 169 12825 189
rect 12845 169 12863 189
rect 12814 157 12863 169
rect 12913 193 12957 199
rect 12913 173 12928 193
rect 12948 173 12957 193
rect 12913 157 12957 173
rect 13027 193 13071 199
rect 13027 173 13036 193
rect 13056 173 13071 193
rect 13027 157 13071 173
rect 13121 189 13170 199
rect 13121 169 13139 189
rect 13159 169 13170 189
rect 13121 157 13170 169
rect 17674 168 17723 178
rect 17674 148 17685 168
rect 17705 148 17723 168
rect 17674 136 17723 148
rect 17773 172 17817 178
rect 17773 152 17788 172
rect 17808 152 17817 172
rect 17773 136 17817 152
rect 17887 168 17936 178
rect 17887 148 17898 168
rect 17918 148 17936 168
rect 17887 136 17936 148
rect 17986 172 18030 178
rect 17986 152 18001 172
rect 18021 152 18030 172
rect 17986 136 18030 152
rect 18095 168 18144 178
rect 18095 148 18106 168
rect 18126 148 18144 168
rect 18095 136 18144 148
rect 18194 172 18238 178
rect 18194 152 18209 172
rect 18229 152 18238 172
rect 18194 136 18238 152
rect 18308 172 18352 178
rect 18308 152 18317 172
rect 18337 152 18352 172
rect 18308 136 18352 152
rect 18402 168 18451 178
rect 18402 148 18420 168
rect 18440 148 18451 168
rect 18402 136 18451 148
rect 15483 101 15532 111
rect 5550 73 5568 93
rect 5588 73 5599 93
rect 5550 61 5599 73
rect 10083 86 10132 96
rect 10083 66 10094 86
rect 10114 66 10132 86
rect 10083 54 10132 66
rect 10182 90 10226 96
rect 10182 70 10197 90
rect 10217 70 10226 90
rect 10182 54 10226 70
rect 10296 86 10345 96
rect 10296 66 10307 86
rect 10327 66 10345 86
rect 10296 54 10345 66
rect 10395 90 10439 96
rect 10395 70 10410 90
rect 10430 70 10439 90
rect 10395 54 10439 70
rect 10504 86 10553 96
rect 10504 66 10515 86
rect 10535 66 10553 86
rect 10504 54 10553 66
rect 10603 90 10647 96
rect 10603 70 10618 90
rect 10638 70 10647 90
rect 10603 54 10647 70
rect 10717 90 10761 96
rect 10717 70 10726 90
rect 10746 70 10761 90
rect 10717 54 10761 70
rect 10811 86 10860 96
rect 10811 66 10829 86
rect 10849 66 10860 86
rect 15483 81 15494 101
rect 15514 81 15532 101
rect 15483 69 15532 81
rect 15582 105 15626 111
rect 15582 85 15597 105
rect 15617 85 15626 105
rect 15582 69 15626 85
rect 15696 101 15745 111
rect 15696 81 15707 101
rect 15727 81 15745 101
rect 15696 69 15745 81
rect 15795 105 15839 111
rect 15795 85 15810 105
rect 15830 85 15839 105
rect 15795 69 15839 85
rect 15904 101 15953 111
rect 15904 81 15915 101
rect 15935 81 15953 101
rect 15904 69 15953 81
rect 16003 105 16047 111
rect 16003 85 16018 105
rect 16038 85 16047 105
rect 16003 69 16047 85
rect 16117 105 16161 111
rect 16117 85 16126 105
rect 16146 85 16161 105
rect 16117 69 16161 85
rect 16211 101 16260 111
rect 16211 81 16229 101
rect 16249 81 16260 101
rect 16211 69 16260 81
rect 10811 54 10860 66
<< pdiff >>
rect 298 8084 342 8122
rect 298 8064 310 8084
rect 330 8064 342 8084
rect 298 8022 342 8064
rect 392 8084 434 8122
rect 392 8064 406 8084
rect 426 8064 434 8084
rect 392 8022 434 8064
rect 511 8084 555 8122
rect 511 8064 523 8084
rect 543 8064 555 8084
rect 511 8022 555 8064
rect 605 8084 647 8122
rect 605 8064 619 8084
rect 639 8064 647 8084
rect 605 8022 647 8064
rect 719 8084 763 8122
rect 719 8064 731 8084
rect 751 8064 763 8084
rect 719 8022 763 8064
rect 813 8084 855 8122
rect 813 8064 827 8084
rect 847 8064 855 8084
rect 813 8022 855 8064
rect 929 8084 971 8122
rect 929 8064 937 8084
rect 957 8064 971 8084
rect 929 8022 971 8064
rect 1021 8091 1066 8122
rect 4127 8118 4171 8160
rect 4127 8098 4139 8118
rect 4159 8098 4171 8118
rect 4127 8091 4171 8098
rect 1021 8084 1065 8091
rect 1021 8064 1033 8084
rect 1053 8064 1065 8084
rect 1021 8022 1065 8064
rect 4126 8060 4171 8091
rect 4221 8118 4263 8160
rect 4221 8098 4235 8118
rect 4255 8098 4263 8118
rect 4221 8060 4263 8098
rect 4337 8118 4379 8160
rect 4337 8098 4345 8118
rect 4365 8098 4379 8118
rect 4337 8060 4379 8098
rect 4429 8118 4473 8160
rect 4429 8098 4441 8118
rect 4461 8098 4473 8118
rect 4429 8060 4473 8098
rect 4545 8118 4587 8160
rect 4545 8098 4553 8118
rect 4573 8098 4587 8118
rect 4545 8060 4587 8098
rect 4637 8118 4681 8160
rect 4637 8098 4649 8118
rect 4669 8098 4681 8118
rect 4637 8060 4681 8098
rect 4758 8118 4800 8160
rect 4758 8098 4766 8118
rect 4786 8098 4800 8118
rect 4758 8060 4800 8098
rect 4850 8118 4894 8160
rect 4850 8098 4862 8118
rect 4882 8098 4894 8118
rect 4850 8060 4894 8098
rect 5579 8063 5623 8101
rect 5579 8043 5591 8063
rect 5611 8043 5623 8063
rect 1310 7903 1354 7941
rect 1310 7883 1322 7903
rect 1342 7883 1354 7903
rect 1310 7841 1354 7883
rect 1404 7903 1446 7941
rect 1404 7883 1418 7903
rect 1438 7883 1446 7903
rect 1404 7841 1446 7883
rect 1523 7903 1567 7941
rect 1523 7883 1535 7903
rect 1555 7883 1567 7903
rect 1523 7841 1567 7883
rect 1617 7903 1659 7941
rect 1617 7883 1631 7903
rect 1651 7883 1659 7903
rect 1617 7841 1659 7883
rect 1731 7903 1775 7941
rect 1731 7883 1743 7903
rect 1763 7883 1775 7903
rect 1731 7841 1775 7883
rect 1825 7903 1867 7941
rect 1825 7883 1839 7903
rect 1859 7883 1867 7903
rect 1825 7841 1867 7883
rect 1941 7903 1983 7941
rect 1941 7883 1949 7903
rect 1969 7883 1983 7903
rect 1941 7841 1983 7883
rect 2033 7910 2078 7941
rect 5579 8001 5623 8043
rect 5673 8063 5715 8101
rect 5673 8043 5687 8063
rect 5707 8043 5715 8063
rect 5673 8001 5715 8043
rect 5792 8063 5836 8101
rect 5792 8043 5804 8063
rect 5824 8043 5836 8063
rect 5792 8001 5836 8043
rect 5886 8063 5928 8101
rect 5886 8043 5900 8063
rect 5920 8043 5928 8063
rect 5886 8001 5928 8043
rect 6000 8063 6044 8101
rect 6000 8043 6012 8063
rect 6032 8043 6044 8063
rect 6000 8001 6044 8043
rect 6094 8063 6136 8101
rect 6094 8043 6108 8063
rect 6128 8043 6136 8063
rect 6094 8001 6136 8043
rect 6210 8063 6252 8101
rect 6210 8043 6218 8063
rect 6238 8043 6252 8063
rect 6210 8001 6252 8043
rect 6302 8070 6347 8101
rect 9408 8097 9452 8139
rect 9408 8077 9420 8097
rect 9440 8077 9452 8097
rect 9408 8070 9452 8077
rect 6302 8063 6346 8070
rect 6302 8043 6314 8063
rect 6334 8043 6346 8063
rect 6302 8001 6346 8043
rect 9407 8039 9452 8070
rect 9502 8097 9544 8139
rect 9502 8077 9516 8097
rect 9536 8077 9544 8097
rect 9502 8039 9544 8077
rect 9618 8097 9660 8139
rect 9618 8077 9626 8097
rect 9646 8077 9660 8097
rect 9618 8039 9660 8077
rect 9710 8097 9754 8139
rect 9710 8077 9722 8097
rect 9742 8077 9754 8097
rect 9710 8039 9754 8077
rect 9826 8097 9868 8139
rect 9826 8077 9834 8097
rect 9854 8077 9868 8097
rect 9826 8039 9868 8077
rect 9918 8097 9962 8139
rect 9918 8077 9930 8097
rect 9950 8077 9962 8097
rect 9918 8039 9962 8077
rect 10039 8097 10081 8139
rect 10039 8077 10047 8097
rect 10067 8077 10081 8097
rect 10039 8039 10081 8077
rect 10131 8097 10175 8139
rect 10131 8077 10143 8097
rect 10163 8077 10175 8097
rect 10131 8039 10175 8077
rect 10959 8092 11003 8130
rect 10959 8072 10971 8092
rect 10991 8072 11003 8092
rect 2033 7903 2077 7910
rect 2033 7883 2045 7903
rect 2065 7883 2077 7903
rect 2033 7841 2077 7883
rect 3114 7884 3158 7926
rect 3114 7864 3126 7884
rect 3146 7864 3158 7884
rect 3114 7857 3158 7864
rect 3113 7826 3158 7857
rect 3208 7884 3250 7926
rect 3208 7864 3222 7884
rect 3242 7864 3250 7884
rect 3208 7826 3250 7864
rect 3324 7884 3366 7926
rect 3324 7864 3332 7884
rect 3352 7864 3366 7884
rect 3324 7826 3366 7864
rect 3416 7884 3460 7926
rect 3416 7864 3428 7884
rect 3448 7864 3460 7884
rect 3416 7826 3460 7864
rect 3532 7884 3574 7926
rect 3532 7864 3540 7884
rect 3560 7864 3574 7884
rect 3532 7826 3574 7864
rect 3624 7884 3668 7926
rect 3624 7864 3636 7884
rect 3656 7864 3668 7884
rect 3624 7826 3668 7864
rect 3745 7884 3787 7926
rect 3745 7864 3753 7884
rect 3773 7864 3787 7884
rect 3745 7826 3787 7864
rect 3837 7884 3881 7926
rect 10959 8030 11003 8072
rect 11053 8092 11095 8130
rect 11053 8072 11067 8092
rect 11087 8072 11095 8092
rect 11053 8030 11095 8072
rect 11172 8092 11216 8130
rect 11172 8072 11184 8092
rect 11204 8072 11216 8092
rect 11172 8030 11216 8072
rect 11266 8092 11308 8130
rect 11266 8072 11280 8092
rect 11300 8072 11308 8092
rect 11266 8030 11308 8072
rect 11380 8092 11424 8130
rect 11380 8072 11392 8092
rect 11412 8072 11424 8092
rect 11380 8030 11424 8072
rect 11474 8092 11516 8130
rect 11474 8072 11488 8092
rect 11508 8072 11516 8092
rect 11474 8030 11516 8072
rect 11590 8092 11632 8130
rect 11590 8072 11598 8092
rect 11618 8072 11632 8092
rect 11590 8030 11632 8072
rect 11682 8099 11727 8130
rect 14788 8126 14832 8168
rect 14788 8106 14800 8126
rect 14820 8106 14832 8126
rect 14788 8099 14832 8106
rect 11682 8092 11726 8099
rect 11682 8072 11694 8092
rect 11714 8072 11726 8092
rect 11682 8030 11726 8072
rect 14787 8068 14832 8099
rect 14882 8126 14924 8168
rect 14882 8106 14896 8126
rect 14916 8106 14924 8126
rect 14882 8068 14924 8106
rect 14998 8126 15040 8168
rect 14998 8106 15006 8126
rect 15026 8106 15040 8126
rect 14998 8068 15040 8106
rect 15090 8126 15134 8168
rect 15090 8106 15102 8126
rect 15122 8106 15134 8126
rect 15090 8068 15134 8106
rect 15206 8126 15248 8168
rect 15206 8106 15214 8126
rect 15234 8106 15248 8126
rect 15206 8068 15248 8106
rect 15298 8126 15342 8168
rect 15298 8106 15310 8126
rect 15330 8106 15342 8126
rect 15298 8068 15342 8106
rect 15419 8126 15461 8168
rect 15419 8106 15427 8126
rect 15447 8106 15461 8126
rect 15419 8068 15461 8106
rect 15511 8126 15555 8168
rect 15511 8106 15523 8126
rect 15543 8106 15555 8126
rect 15511 8068 15555 8106
rect 3837 7864 3849 7884
rect 3869 7864 3881 7884
rect 6591 7882 6635 7920
rect 3837 7826 3881 7864
rect 6591 7862 6603 7882
rect 6623 7862 6635 7882
rect 6591 7820 6635 7862
rect 6685 7882 6727 7920
rect 6685 7862 6699 7882
rect 6719 7862 6727 7882
rect 6685 7820 6727 7862
rect 6804 7882 6848 7920
rect 6804 7862 6816 7882
rect 6836 7862 6848 7882
rect 6804 7820 6848 7862
rect 6898 7882 6940 7920
rect 6898 7862 6912 7882
rect 6932 7862 6940 7882
rect 6898 7820 6940 7862
rect 7012 7882 7056 7920
rect 7012 7862 7024 7882
rect 7044 7862 7056 7882
rect 7012 7820 7056 7862
rect 7106 7882 7148 7920
rect 7106 7862 7120 7882
rect 7140 7862 7148 7882
rect 7106 7820 7148 7862
rect 7222 7882 7264 7920
rect 7222 7862 7230 7882
rect 7250 7862 7264 7882
rect 7222 7820 7264 7862
rect 7314 7889 7359 7920
rect 16240 8071 16284 8109
rect 16240 8051 16252 8071
rect 16272 8051 16284 8071
rect 11971 7911 12015 7949
rect 7314 7882 7358 7889
rect 7314 7862 7326 7882
rect 7346 7862 7358 7882
rect 7314 7820 7358 7862
rect 8395 7863 8439 7905
rect 8395 7843 8407 7863
rect 8427 7843 8439 7863
rect 8395 7836 8439 7843
rect 297 7669 341 7707
rect 297 7649 309 7669
rect 329 7649 341 7669
rect 297 7607 341 7649
rect 391 7669 433 7707
rect 391 7649 405 7669
rect 425 7649 433 7669
rect 391 7607 433 7649
rect 510 7669 554 7707
rect 510 7649 522 7669
rect 542 7649 554 7669
rect 510 7607 554 7649
rect 604 7669 646 7707
rect 604 7649 618 7669
rect 638 7649 646 7669
rect 604 7607 646 7649
rect 718 7669 762 7707
rect 718 7649 730 7669
rect 750 7649 762 7669
rect 718 7607 762 7649
rect 812 7669 854 7707
rect 812 7649 826 7669
rect 846 7649 854 7669
rect 812 7607 854 7649
rect 928 7669 970 7707
rect 928 7649 936 7669
rect 956 7649 970 7669
rect 928 7607 970 7649
rect 1020 7676 1065 7707
rect 4126 7703 4170 7745
rect 4126 7683 4138 7703
rect 4158 7683 4170 7703
rect 4126 7676 4170 7683
rect 1020 7669 1064 7676
rect 1020 7649 1032 7669
rect 1052 7649 1064 7669
rect 1020 7607 1064 7649
rect 4125 7645 4170 7676
rect 4220 7703 4262 7745
rect 4220 7683 4234 7703
rect 4254 7683 4262 7703
rect 4220 7645 4262 7683
rect 4336 7703 4378 7745
rect 4336 7683 4344 7703
rect 4364 7683 4378 7703
rect 4336 7645 4378 7683
rect 4428 7703 4472 7745
rect 4428 7683 4440 7703
rect 4460 7683 4472 7703
rect 4428 7645 4472 7683
rect 4544 7703 4586 7745
rect 4544 7683 4552 7703
rect 4572 7683 4586 7703
rect 4544 7645 4586 7683
rect 4636 7703 4680 7745
rect 4636 7683 4648 7703
rect 4668 7683 4680 7703
rect 4636 7645 4680 7683
rect 4757 7703 4799 7745
rect 4757 7683 4765 7703
rect 4785 7683 4799 7703
rect 4757 7645 4799 7683
rect 4849 7703 4893 7745
rect 8394 7805 8439 7836
rect 8489 7863 8531 7905
rect 8489 7843 8503 7863
rect 8523 7843 8531 7863
rect 8489 7805 8531 7843
rect 8605 7863 8647 7905
rect 8605 7843 8613 7863
rect 8633 7843 8647 7863
rect 8605 7805 8647 7843
rect 8697 7863 8741 7905
rect 8697 7843 8709 7863
rect 8729 7843 8741 7863
rect 8697 7805 8741 7843
rect 8813 7863 8855 7905
rect 8813 7843 8821 7863
rect 8841 7843 8855 7863
rect 8813 7805 8855 7843
rect 8905 7863 8949 7905
rect 8905 7843 8917 7863
rect 8937 7843 8949 7863
rect 8905 7805 8949 7843
rect 9026 7863 9068 7905
rect 9026 7843 9034 7863
rect 9054 7843 9068 7863
rect 9026 7805 9068 7843
rect 9118 7863 9162 7905
rect 9118 7843 9130 7863
rect 9150 7843 9162 7863
rect 11971 7891 11983 7911
rect 12003 7891 12015 7911
rect 11971 7849 12015 7891
rect 12065 7911 12107 7949
rect 12065 7891 12079 7911
rect 12099 7891 12107 7911
rect 12065 7849 12107 7891
rect 12184 7911 12228 7949
rect 12184 7891 12196 7911
rect 12216 7891 12228 7911
rect 12184 7849 12228 7891
rect 12278 7911 12320 7949
rect 12278 7891 12292 7911
rect 12312 7891 12320 7911
rect 12278 7849 12320 7891
rect 12392 7911 12436 7949
rect 12392 7891 12404 7911
rect 12424 7891 12436 7911
rect 12392 7849 12436 7891
rect 12486 7911 12528 7949
rect 12486 7891 12500 7911
rect 12520 7891 12528 7911
rect 12486 7849 12528 7891
rect 12602 7911 12644 7949
rect 12602 7891 12610 7911
rect 12630 7891 12644 7911
rect 12602 7849 12644 7891
rect 12694 7918 12739 7949
rect 16240 8009 16284 8051
rect 16334 8071 16376 8109
rect 16334 8051 16348 8071
rect 16368 8051 16376 8071
rect 16334 8009 16376 8051
rect 16453 8071 16497 8109
rect 16453 8051 16465 8071
rect 16485 8051 16497 8071
rect 16453 8009 16497 8051
rect 16547 8071 16589 8109
rect 16547 8051 16561 8071
rect 16581 8051 16589 8071
rect 16547 8009 16589 8051
rect 16661 8071 16705 8109
rect 16661 8051 16673 8071
rect 16693 8051 16705 8071
rect 16661 8009 16705 8051
rect 16755 8071 16797 8109
rect 16755 8051 16769 8071
rect 16789 8051 16797 8071
rect 16755 8009 16797 8051
rect 16871 8071 16913 8109
rect 16871 8051 16879 8071
rect 16899 8051 16913 8071
rect 16871 8009 16913 8051
rect 16963 8078 17008 8109
rect 20069 8105 20113 8147
rect 20069 8085 20081 8105
rect 20101 8085 20113 8105
rect 20069 8078 20113 8085
rect 16963 8071 17007 8078
rect 16963 8051 16975 8071
rect 16995 8051 17007 8071
rect 16963 8009 17007 8051
rect 20068 8047 20113 8078
rect 20163 8105 20205 8147
rect 20163 8085 20177 8105
rect 20197 8085 20205 8105
rect 20163 8047 20205 8085
rect 20279 8105 20321 8147
rect 20279 8085 20287 8105
rect 20307 8085 20321 8105
rect 20279 8047 20321 8085
rect 20371 8105 20415 8147
rect 20371 8085 20383 8105
rect 20403 8085 20415 8105
rect 20371 8047 20415 8085
rect 20487 8105 20529 8147
rect 20487 8085 20495 8105
rect 20515 8085 20529 8105
rect 20487 8047 20529 8085
rect 20579 8105 20623 8147
rect 20579 8085 20591 8105
rect 20611 8085 20623 8105
rect 20579 8047 20623 8085
rect 20700 8105 20742 8147
rect 20700 8085 20708 8105
rect 20728 8085 20742 8105
rect 20700 8047 20742 8085
rect 20792 8105 20836 8147
rect 20792 8085 20804 8105
rect 20824 8085 20836 8105
rect 20792 8047 20836 8085
rect 12694 7911 12738 7918
rect 12694 7891 12706 7911
rect 12726 7891 12738 7911
rect 12694 7849 12738 7891
rect 13775 7892 13819 7934
rect 13775 7872 13787 7892
rect 13807 7872 13819 7892
rect 13775 7865 13819 7872
rect 9118 7805 9162 7843
rect 4849 7683 4861 7703
rect 4881 7683 4893 7703
rect 4849 7645 4893 7683
rect 13774 7834 13819 7865
rect 13869 7892 13911 7934
rect 13869 7872 13883 7892
rect 13903 7872 13911 7892
rect 13869 7834 13911 7872
rect 13985 7892 14027 7934
rect 13985 7872 13993 7892
rect 14013 7872 14027 7892
rect 13985 7834 14027 7872
rect 14077 7892 14121 7934
rect 14077 7872 14089 7892
rect 14109 7872 14121 7892
rect 14077 7834 14121 7872
rect 14193 7892 14235 7934
rect 14193 7872 14201 7892
rect 14221 7872 14235 7892
rect 14193 7834 14235 7872
rect 14285 7892 14329 7934
rect 14285 7872 14297 7892
rect 14317 7872 14329 7892
rect 14285 7834 14329 7872
rect 14406 7892 14448 7934
rect 14406 7872 14414 7892
rect 14434 7872 14448 7892
rect 14406 7834 14448 7872
rect 14498 7892 14542 7934
rect 14498 7872 14510 7892
rect 14530 7872 14542 7892
rect 17252 7890 17296 7928
rect 14498 7834 14542 7872
rect 17252 7870 17264 7890
rect 17284 7870 17296 7890
rect 5578 7648 5622 7686
rect 5578 7628 5590 7648
rect 5610 7628 5622 7648
rect 5578 7586 5622 7628
rect 5672 7648 5714 7686
rect 5672 7628 5686 7648
rect 5706 7628 5714 7648
rect 5672 7586 5714 7628
rect 5791 7648 5835 7686
rect 5791 7628 5803 7648
rect 5823 7628 5835 7648
rect 5791 7586 5835 7628
rect 5885 7648 5927 7686
rect 5885 7628 5899 7648
rect 5919 7628 5927 7648
rect 5885 7586 5927 7628
rect 5999 7648 6043 7686
rect 5999 7628 6011 7648
rect 6031 7628 6043 7648
rect 5999 7586 6043 7628
rect 6093 7648 6135 7686
rect 6093 7628 6107 7648
rect 6127 7628 6135 7648
rect 6093 7586 6135 7628
rect 6209 7648 6251 7686
rect 6209 7628 6217 7648
rect 6237 7628 6251 7648
rect 6209 7586 6251 7628
rect 6301 7655 6346 7686
rect 9407 7682 9451 7724
rect 9407 7662 9419 7682
rect 9439 7662 9451 7682
rect 9407 7655 9451 7662
rect 6301 7648 6345 7655
rect 6301 7628 6313 7648
rect 6333 7628 6345 7648
rect 6301 7586 6345 7628
rect 9406 7624 9451 7655
rect 9501 7682 9543 7724
rect 9501 7662 9515 7682
rect 9535 7662 9543 7682
rect 9501 7624 9543 7662
rect 9617 7682 9659 7724
rect 9617 7662 9625 7682
rect 9645 7662 9659 7682
rect 9617 7624 9659 7662
rect 9709 7682 9753 7724
rect 9709 7662 9721 7682
rect 9741 7662 9753 7682
rect 9709 7624 9753 7662
rect 9825 7682 9867 7724
rect 9825 7662 9833 7682
rect 9853 7662 9867 7682
rect 9825 7624 9867 7662
rect 9917 7682 9961 7724
rect 9917 7662 9929 7682
rect 9949 7662 9961 7682
rect 9917 7624 9961 7662
rect 10038 7682 10080 7724
rect 10038 7662 10046 7682
rect 10066 7662 10080 7682
rect 10038 7624 10080 7662
rect 10130 7682 10174 7724
rect 17252 7828 17296 7870
rect 17346 7890 17388 7928
rect 17346 7870 17360 7890
rect 17380 7870 17388 7890
rect 17346 7828 17388 7870
rect 17465 7890 17509 7928
rect 17465 7870 17477 7890
rect 17497 7870 17509 7890
rect 17465 7828 17509 7870
rect 17559 7890 17601 7928
rect 17559 7870 17573 7890
rect 17593 7870 17601 7890
rect 17559 7828 17601 7870
rect 17673 7890 17717 7928
rect 17673 7870 17685 7890
rect 17705 7870 17717 7890
rect 17673 7828 17717 7870
rect 17767 7890 17809 7928
rect 17767 7870 17781 7890
rect 17801 7870 17809 7890
rect 17767 7828 17809 7870
rect 17883 7890 17925 7928
rect 17883 7870 17891 7890
rect 17911 7870 17925 7890
rect 17883 7828 17925 7870
rect 17975 7897 18020 7928
rect 17975 7890 18019 7897
rect 17975 7870 17987 7890
rect 18007 7870 18019 7890
rect 17975 7828 18019 7870
rect 19056 7871 19100 7913
rect 19056 7851 19068 7871
rect 19088 7851 19100 7871
rect 19056 7844 19100 7851
rect 10130 7662 10142 7682
rect 10162 7662 10174 7682
rect 10130 7624 10174 7662
rect 10958 7677 11002 7715
rect 10958 7657 10970 7677
rect 10990 7657 11002 7677
rect 10958 7615 11002 7657
rect 11052 7677 11094 7715
rect 11052 7657 11066 7677
rect 11086 7657 11094 7677
rect 11052 7615 11094 7657
rect 11171 7677 11215 7715
rect 11171 7657 11183 7677
rect 11203 7657 11215 7677
rect 11171 7615 11215 7657
rect 11265 7677 11307 7715
rect 11265 7657 11279 7677
rect 11299 7657 11307 7677
rect 11265 7615 11307 7657
rect 11379 7677 11423 7715
rect 11379 7657 11391 7677
rect 11411 7657 11423 7677
rect 11379 7615 11423 7657
rect 11473 7677 11515 7715
rect 11473 7657 11487 7677
rect 11507 7657 11515 7677
rect 11473 7615 11515 7657
rect 11589 7677 11631 7715
rect 11589 7657 11597 7677
rect 11617 7657 11631 7677
rect 11589 7615 11631 7657
rect 11681 7684 11726 7715
rect 14787 7711 14831 7753
rect 14787 7691 14799 7711
rect 14819 7691 14831 7711
rect 14787 7684 14831 7691
rect 11681 7677 11725 7684
rect 11681 7657 11693 7677
rect 11713 7657 11725 7677
rect 11681 7615 11725 7657
rect 14786 7653 14831 7684
rect 14881 7711 14923 7753
rect 14881 7691 14895 7711
rect 14915 7691 14923 7711
rect 14881 7653 14923 7691
rect 14997 7711 15039 7753
rect 14997 7691 15005 7711
rect 15025 7691 15039 7711
rect 14997 7653 15039 7691
rect 15089 7711 15133 7753
rect 15089 7691 15101 7711
rect 15121 7691 15133 7711
rect 15089 7653 15133 7691
rect 15205 7711 15247 7753
rect 15205 7691 15213 7711
rect 15233 7691 15247 7711
rect 15205 7653 15247 7691
rect 15297 7711 15341 7753
rect 15297 7691 15309 7711
rect 15329 7691 15341 7711
rect 15297 7653 15341 7691
rect 15418 7711 15460 7753
rect 15418 7691 15426 7711
rect 15446 7691 15460 7711
rect 15418 7653 15460 7691
rect 15510 7711 15554 7753
rect 19055 7813 19100 7844
rect 19150 7871 19192 7913
rect 19150 7851 19164 7871
rect 19184 7851 19192 7871
rect 19150 7813 19192 7851
rect 19266 7871 19308 7913
rect 19266 7851 19274 7871
rect 19294 7851 19308 7871
rect 19266 7813 19308 7851
rect 19358 7871 19402 7913
rect 19358 7851 19370 7871
rect 19390 7851 19402 7871
rect 19358 7813 19402 7851
rect 19474 7871 19516 7913
rect 19474 7851 19482 7871
rect 19502 7851 19516 7871
rect 19474 7813 19516 7851
rect 19566 7871 19610 7913
rect 19566 7851 19578 7871
rect 19598 7851 19610 7871
rect 19566 7813 19610 7851
rect 19687 7871 19729 7913
rect 19687 7851 19695 7871
rect 19715 7851 19729 7871
rect 19687 7813 19729 7851
rect 19779 7871 19823 7913
rect 19779 7851 19791 7871
rect 19811 7851 19823 7871
rect 19779 7813 19823 7851
rect 15510 7691 15522 7711
rect 15542 7691 15554 7711
rect 15510 7653 15554 7691
rect 16239 7656 16283 7694
rect 16239 7636 16251 7656
rect 16271 7636 16283 7656
rect 3064 7464 3108 7506
rect 3064 7444 3076 7464
rect 3096 7444 3108 7464
rect 3064 7437 3108 7444
rect 3063 7406 3108 7437
rect 3158 7464 3200 7506
rect 3158 7444 3172 7464
rect 3192 7444 3200 7464
rect 3158 7406 3200 7444
rect 3274 7464 3316 7506
rect 3274 7444 3282 7464
rect 3302 7444 3316 7464
rect 3274 7406 3316 7444
rect 3366 7464 3410 7506
rect 3366 7444 3378 7464
rect 3398 7444 3410 7464
rect 3366 7406 3410 7444
rect 3482 7464 3524 7506
rect 3482 7444 3490 7464
rect 3510 7444 3524 7464
rect 3482 7406 3524 7444
rect 3574 7464 3618 7506
rect 3574 7444 3586 7464
rect 3606 7444 3618 7464
rect 3574 7406 3618 7444
rect 3695 7464 3737 7506
rect 3695 7444 3703 7464
rect 3723 7444 3737 7464
rect 3695 7406 3737 7444
rect 3787 7464 3831 7506
rect 3787 7444 3799 7464
rect 3819 7444 3831 7464
rect 3787 7406 3831 7444
rect 8345 7443 8389 7485
rect 8345 7423 8357 7443
rect 8377 7423 8389 7443
rect 8345 7416 8389 7423
rect 8344 7385 8389 7416
rect 8439 7443 8481 7485
rect 8439 7423 8453 7443
rect 8473 7423 8481 7443
rect 8439 7385 8481 7423
rect 8555 7443 8597 7485
rect 8555 7423 8563 7443
rect 8583 7423 8597 7443
rect 8555 7385 8597 7423
rect 8647 7443 8691 7485
rect 8647 7423 8659 7443
rect 8679 7423 8691 7443
rect 8647 7385 8691 7423
rect 8763 7443 8805 7485
rect 8763 7423 8771 7443
rect 8791 7423 8805 7443
rect 8763 7385 8805 7423
rect 8855 7443 8899 7485
rect 8855 7423 8867 7443
rect 8887 7423 8899 7443
rect 8855 7385 8899 7423
rect 8976 7443 9018 7485
rect 8976 7423 8984 7443
rect 9004 7423 9018 7443
rect 8976 7385 9018 7423
rect 9068 7443 9112 7485
rect 16239 7594 16283 7636
rect 16333 7656 16375 7694
rect 16333 7636 16347 7656
rect 16367 7636 16375 7656
rect 16333 7594 16375 7636
rect 16452 7656 16496 7694
rect 16452 7636 16464 7656
rect 16484 7636 16496 7656
rect 16452 7594 16496 7636
rect 16546 7656 16588 7694
rect 16546 7636 16560 7656
rect 16580 7636 16588 7656
rect 16546 7594 16588 7636
rect 16660 7656 16704 7694
rect 16660 7636 16672 7656
rect 16692 7636 16704 7656
rect 16660 7594 16704 7636
rect 16754 7656 16796 7694
rect 16754 7636 16768 7656
rect 16788 7636 16796 7656
rect 16754 7594 16796 7636
rect 16870 7656 16912 7694
rect 16870 7636 16878 7656
rect 16898 7636 16912 7656
rect 16870 7594 16912 7636
rect 16962 7663 17007 7694
rect 20068 7690 20112 7732
rect 20068 7670 20080 7690
rect 20100 7670 20112 7690
rect 20068 7663 20112 7670
rect 16962 7656 17006 7663
rect 16962 7636 16974 7656
rect 16994 7636 17006 7656
rect 16962 7594 17006 7636
rect 20067 7632 20112 7663
rect 20162 7690 20204 7732
rect 20162 7670 20176 7690
rect 20196 7670 20204 7690
rect 20162 7632 20204 7670
rect 20278 7690 20320 7732
rect 20278 7670 20286 7690
rect 20306 7670 20320 7690
rect 20278 7632 20320 7670
rect 20370 7690 20414 7732
rect 20370 7670 20382 7690
rect 20402 7670 20414 7690
rect 20370 7632 20414 7670
rect 20486 7690 20528 7732
rect 20486 7670 20494 7690
rect 20514 7670 20528 7690
rect 20486 7632 20528 7670
rect 20578 7690 20622 7732
rect 20578 7670 20590 7690
rect 20610 7670 20622 7690
rect 20578 7632 20622 7670
rect 20699 7690 20741 7732
rect 20699 7670 20707 7690
rect 20727 7670 20741 7690
rect 20699 7632 20741 7670
rect 20791 7690 20835 7732
rect 20791 7670 20803 7690
rect 20823 7670 20835 7690
rect 20791 7632 20835 7670
rect 9068 7423 9080 7443
rect 9100 7423 9112 7443
rect 9068 7385 9112 7423
rect 13725 7472 13769 7514
rect 13725 7452 13737 7472
rect 13757 7452 13769 7472
rect 13725 7445 13769 7452
rect 13724 7414 13769 7445
rect 13819 7472 13861 7514
rect 13819 7452 13833 7472
rect 13853 7452 13861 7472
rect 13819 7414 13861 7452
rect 13935 7472 13977 7514
rect 13935 7452 13943 7472
rect 13963 7452 13977 7472
rect 13935 7414 13977 7452
rect 14027 7472 14071 7514
rect 14027 7452 14039 7472
rect 14059 7452 14071 7472
rect 14027 7414 14071 7452
rect 14143 7472 14185 7514
rect 14143 7452 14151 7472
rect 14171 7452 14185 7472
rect 14143 7414 14185 7452
rect 14235 7472 14279 7514
rect 14235 7452 14247 7472
rect 14267 7452 14279 7472
rect 14235 7414 14279 7452
rect 14356 7472 14398 7514
rect 14356 7452 14364 7472
rect 14384 7452 14398 7472
rect 14356 7414 14398 7452
rect 14448 7472 14492 7514
rect 14448 7452 14460 7472
rect 14480 7452 14492 7472
rect 14448 7414 14492 7452
rect 19006 7451 19050 7493
rect 19006 7431 19018 7451
rect 19038 7431 19050 7451
rect 19006 7424 19050 7431
rect 19005 7393 19050 7424
rect 19100 7451 19142 7493
rect 19100 7431 19114 7451
rect 19134 7431 19142 7451
rect 19100 7393 19142 7431
rect 19216 7451 19258 7493
rect 19216 7431 19224 7451
rect 19244 7431 19258 7451
rect 19216 7393 19258 7431
rect 19308 7451 19352 7493
rect 19308 7431 19320 7451
rect 19340 7431 19352 7451
rect 19308 7393 19352 7431
rect 19424 7451 19466 7493
rect 19424 7431 19432 7451
rect 19452 7431 19466 7451
rect 19424 7393 19466 7431
rect 19516 7451 19560 7493
rect 19516 7431 19528 7451
rect 19548 7431 19560 7451
rect 19516 7393 19560 7431
rect 19637 7451 19679 7493
rect 19637 7431 19645 7451
rect 19665 7431 19679 7451
rect 19637 7393 19679 7431
rect 19729 7451 19773 7493
rect 19729 7431 19741 7451
rect 19761 7431 19773 7451
rect 19729 7393 19773 7431
rect 1365 7342 1409 7380
rect 1365 7322 1377 7342
rect 1397 7322 1409 7342
rect 1365 7280 1409 7322
rect 1459 7342 1501 7380
rect 1459 7322 1473 7342
rect 1493 7322 1501 7342
rect 1459 7280 1501 7322
rect 1578 7342 1622 7380
rect 1578 7322 1590 7342
rect 1610 7322 1622 7342
rect 1578 7280 1622 7322
rect 1672 7342 1714 7380
rect 1672 7322 1686 7342
rect 1706 7322 1714 7342
rect 1672 7280 1714 7322
rect 1786 7342 1830 7380
rect 1786 7322 1798 7342
rect 1818 7322 1830 7342
rect 1786 7280 1830 7322
rect 1880 7342 1922 7380
rect 1880 7322 1894 7342
rect 1914 7322 1922 7342
rect 1880 7280 1922 7322
rect 1996 7342 2038 7380
rect 1996 7322 2004 7342
rect 2024 7322 2038 7342
rect 1996 7280 2038 7322
rect 2088 7349 2133 7380
rect 2088 7342 2132 7349
rect 2088 7322 2100 7342
rect 2120 7322 2132 7342
rect 2088 7280 2132 7322
rect 6646 7321 6690 7359
rect 6646 7301 6658 7321
rect 6678 7301 6690 7321
rect 6646 7259 6690 7301
rect 6740 7321 6782 7359
rect 6740 7301 6754 7321
rect 6774 7301 6782 7321
rect 6740 7259 6782 7301
rect 6859 7321 6903 7359
rect 6859 7301 6871 7321
rect 6891 7301 6903 7321
rect 6859 7259 6903 7301
rect 6953 7321 6995 7359
rect 6953 7301 6967 7321
rect 6987 7301 6995 7321
rect 6953 7259 6995 7301
rect 7067 7321 7111 7359
rect 7067 7301 7079 7321
rect 7099 7301 7111 7321
rect 7067 7259 7111 7301
rect 7161 7321 7203 7359
rect 7161 7301 7175 7321
rect 7195 7301 7203 7321
rect 7161 7259 7203 7301
rect 7277 7321 7319 7359
rect 7277 7301 7285 7321
rect 7305 7301 7319 7321
rect 7277 7259 7319 7301
rect 7369 7328 7414 7359
rect 7369 7321 7413 7328
rect 7369 7301 7381 7321
rect 7401 7301 7413 7321
rect 7369 7259 7413 7301
rect 12026 7350 12070 7388
rect 12026 7330 12038 7350
rect 12058 7330 12070 7350
rect 303 7103 347 7141
rect 303 7083 315 7103
rect 335 7083 347 7103
rect 303 7041 347 7083
rect 397 7103 439 7141
rect 397 7083 411 7103
rect 431 7083 439 7103
rect 397 7041 439 7083
rect 516 7103 560 7141
rect 516 7083 528 7103
rect 548 7083 560 7103
rect 516 7041 560 7083
rect 610 7103 652 7141
rect 610 7083 624 7103
rect 644 7083 652 7103
rect 610 7041 652 7083
rect 724 7103 768 7141
rect 724 7083 736 7103
rect 756 7083 768 7103
rect 724 7041 768 7083
rect 818 7103 860 7141
rect 818 7083 832 7103
rect 852 7083 860 7103
rect 818 7041 860 7083
rect 934 7103 976 7141
rect 934 7083 942 7103
rect 962 7083 976 7103
rect 934 7041 976 7083
rect 1026 7110 1071 7141
rect 4132 7137 4176 7179
rect 4132 7117 4144 7137
rect 4164 7117 4176 7137
rect 4132 7110 4176 7117
rect 1026 7103 1070 7110
rect 1026 7083 1038 7103
rect 1058 7083 1070 7103
rect 1026 7041 1070 7083
rect 4131 7079 4176 7110
rect 4226 7137 4268 7179
rect 4226 7117 4240 7137
rect 4260 7117 4268 7137
rect 4226 7079 4268 7117
rect 4342 7137 4384 7179
rect 4342 7117 4350 7137
rect 4370 7117 4384 7137
rect 4342 7079 4384 7117
rect 4434 7137 4478 7179
rect 4434 7117 4446 7137
rect 4466 7117 4478 7137
rect 4434 7079 4478 7117
rect 4550 7137 4592 7179
rect 4550 7117 4558 7137
rect 4578 7117 4592 7137
rect 4550 7079 4592 7117
rect 4642 7137 4686 7179
rect 4642 7117 4654 7137
rect 4674 7117 4686 7137
rect 4642 7079 4686 7117
rect 4763 7137 4805 7179
rect 4763 7117 4771 7137
rect 4791 7117 4805 7137
rect 4763 7079 4805 7117
rect 4855 7137 4899 7179
rect 12026 7288 12070 7330
rect 12120 7350 12162 7388
rect 12120 7330 12134 7350
rect 12154 7330 12162 7350
rect 12120 7288 12162 7330
rect 12239 7350 12283 7388
rect 12239 7330 12251 7350
rect 12271 7330 12283 7350
rect 12239 7288 12283 7330
rect 12333 7350 12375 7388
rect 12333 7330 12347 7350
rect 12367 7330 12375 7350
rect 12333 7288 12375 7330
rect 12447 7350 12491 7388
rect 12447 7330 12459 7350
rect 12479 7330 12491 7350
rect 12447 7288 12491 7330
rect 12541 7350 12583 7388
rect 12541 7330 12555 7350
rect 12575 7330 12583 7350
rect 12541 7288 12583 7330
rect 12657 7350 12699 7388
rect 12657 7330 12665 7350
rect 12685 7330 12699 7350
rect 12657 7288 12699 7330
rect 12749 7357 12794 7388
rect 12749 7350 12793 7357
rect 12749 7330 12761 7350
rect 12781 7330 12793 7350
rect 12749 7288 12793 7330
rect 17307 7329 17351 7367
rect 17307 7309 17319 7329
rect 17339 7309 17351 7329
rect 17307 7267 17351 7309
rect 17401 7329 17443 7367
rect 17401 7309 17415 7329
rect 17435 7309 17443 7329
rect 17401 7267 17443 7309
rect 17520 7329 17564 7367
rect 17520 7309 17532 7329
rect 17552 7309 17564 7329
rect 17520 7267 17564 7309
rect 17614 7329 17656 7367
rect 17614 7309 17628 7329
rect 17648 7309 17656 7329
rect 17614 7267 17656 7309
rect 17728 7329 17772 7367
rect 17728 7309 17740 7329
rect 17760 7309 17772 7329
rect 17728 7267 17772 7309
rect 17822 7329 17864 7367
rect 17822 7309 17836 7329
rect 17856 7309 17864 7329
rect 17822 7267 17864 7309
rect 17938 7329 17980 7367
rect 17938 7309 17946 7329
rect 17966 7309 17980 7329
rect 17938 7267 17980 7309
rect 18030 7336 18075 7367
rect 18030 7329 18074 7336
rect 18030 7309 18042 7329
rect 18062 7309 18074 7329
rect 18030 7267 18074 7309
rect 4855 7117 4867 7137
rect 4887 7117 4899 7137
rect 4855 7079 4899 7117
rect 5584 7082 5628 7120
rect 5584 7062 5596 7082
rect 5616 7062 5628 7082
rect 1315 6922 1359 6960
rect 1315 6902 1327 6922
rect 1347 6902 1359 6922
rect 1315 6860 1359 6902
rect 1409 6922 1451 6960
rect 1409 6902 1423 6922
rect 1443 6902 1451 6922
rect 1409 6860 1451 6902
rect 1528 6922 1572 6960
rect 1528 6902 1540 6922
rect 1560 6902 1572 6922
rect 1528 6860 1572 6902
rect 1622 6922 1664 6960
rect 1622 6902 1636 6922
rect 1656 6902 1664 6922
rect 1622 6860 1664 6902
rect 1736 6922 1780 6960
rect 1736 6902 1748 6922
rect 1768 6902 1780 6922
rect 1736 6860 1780 6902
rect 1830 6922 1872 6960
rect 1830 6902 1844 6922
rect 1864 6902 1872 6922
rect 1830 6860 1872 6902
rect 1946 6922 1988 6960
rect 1946 6902 1954 6922
rect 1974 6902 1988 6922
rect 1946 6860 1988 6902
rect 2038 6929 2083 6960
rect 5584 7020 5628 7062
rect 5678 7082 5720 7120
rect 5678 7062 5692 7082
rect 5712 7062 5720 7082
rect 5678 7020 5720 7062
rect 5797 7082 5841 7120
rect 5797 7062 5809 7082
rect 5829 7062 5841 7082
rect 5797 7020 5841 7062
rect 5891 7082 5933 7120
rect 5891 7062 5905 7082
rect 5925 7062 5933 7082
rect 5891 7020 5933 7062
rect 6005 7082 6049 7120
rect 6005 7062 6017 7082
rect 6037 7062 6049 7082
rect 6005 7020 6049 7062
rect 6099 7082 6141 7120
rect 6099 7062 6113 7082
rect 6133 7062 6141 7082
rect 6099 7020 6141 7062
rect 6215 7082 6257 7120
rect 6215 7062 6223 7082
rect 6243 7062 6257 7082
rect 6215 7020 6257 7062
rect 6307 7089 6352 7120
rect 9413 7116 9457 7158
rect 9413 7096 9425 7116
rect 9445 7096 9457 7116
rect 9413 7089 9457 7096
rect 6307 7082 6351 7089
rect 6307 7062 6319 7082
rect 6339 7062 6351 7082
rect 6307 7020 6351 7062
rect 9412 7058 9457 7089
rect 9507 7116 9549 7158
rect 9507 7096 9521 7116
rect 9541 7096 9549 7116
rect 9507 7058 9549 7096
rect 9623 7116 9665 7158
rect 9623 7096 9631 7116
rect 9651 7096 9665 7116
rect 9623 7058 9665 7096
rect 9715 7116 9759 7158
rect 9715 7096 9727 7116
rect 9747 7096 9759 7116
rect 9715 7058 9759 7096
rect 9831 7116 9873 7158
rect 9831 7096 9839 7116
rect 9859 7096 9873 7116
rect 9831 7058 9873 7096
rect 9923 7116 9967 7158
rect 9923 7096 9935 7116
rect 9955 7096 9967 7116
rect 9923 7058 9967 7096
rect 10044 7116 10086 7158
rect 10044 7096 10052 7116
rect 10072 7096 10086 7116
rect 10044 7058 10086 7096
rect 10136 7116 10180 7158
rect 10136 7096 10148 7116
rect 10168 7096 10180 7116
rect 10136 7058 10180 7096
rect 10964 7111 11008 7149
rect 10964 7091 10976 7111
rect 10996 7091 11008 7111
rect 2038 6922 2082 6929
rect 2038 6902 2050 6922
rect 2070 6902 2082 6922
rect 2038 6860 2082 6902
rect 3119 6903 3163 6945
rect 3119 6883 3131 6903
rect 3151 6883 3163 6903
rect 3119 6876 3163 6883
rect 3118 6845 3163 6876
rect 3213 6903 3255 6945
rect 3213 6883 3227 6903
rect 3247 6883 3255 6903
rect 3213 6845 3255 6883
rect 3329 6903 3371 6945
rect 3329 6883 3337 6903
rect 3357 6883 3371 6903
rect 3329 6845 3371 6883
rect 3421 6903 3465 6945
rect 3421 6883 3433 6903
rect 3453 6883 3465 6903
rect 3421 6845 3465 6883
rect 3537 6903 3579 6945
rect 3537 6883 3545 6903
rect 3565 6883 3579 6903
rect 3537 6845 3579 6883
rect 3629 6903 3673 6945
rect 3629 6883 3641 6903
rect 3661 6883 3673 6903
rect 3629 6845 3673 6883
rect 3750 6903 3792 6945
rect 3750 6883 3758 6903
rect 3778 6883 3792 6903
rect 3750 6845 3792 6883
rect 3842 6903 3886 6945
rect 10964 7049 11008 7091
rect 11058 7111 11100 7149
rect 11058 7091 11072 7111
rect 11092 7091 11100 7111
rect 11058 7049 11100 7091
rect 11177 7111 11221 7149
rect 11177 7091 11189 7111
rect 11209 7091 11221 7111
rect 11177 7049 11221 7091
rect 11271 7111 11313 7149
rect 11271 7091 11285 7111
rect 11305 7091 11313 7111
rect 11271 7049 11313 7091
rect 11385 7111 11429 7149
rect 11385 7091 11397 7111
rect 11417 7091 11429 7111
rect 11385 7049 11429 7091
rect 11479 7111 11521 7149
rect 11479 7091 11493 7111
rect 11513 7091 11521 7111
rect 11479 7049 11521 7091
rect 11595 7111 11637 7149
rect 11595 7091 11603 7111
rect 11623 7091 11637 7111
rect 11595 7049 11637 7091
rect 11687 7118 11732 7149
rect 14793 7145 14837 7187
rect 14793 7125 14805 7145
rect 14825 7125 14837 7145
rect 14793 7118 14837 7125
rect 11687 7111 11731 7118
rect 11687 7091 11699 7111
rect 11719 7091 11731 7111
rect 11687 7049 11731 7091
rect 14792 7087 14837 7118
rect 14887 7145 14929 7187
rect 14887 7125 14901 7145
rect 14921 7125 14929 7145
rect 14887 7087 14929 7125
rect 15003 7145 15045 7187
rect 15003 7125 15011 7145
rect 15031 7125 15045 7145
rect 15003 7087 15045 7125
rect 15095 7145 15139 7187
rect 15095 7125 15107 7145
rect 15127 7125 15139 7145
rect 15095 7087 15139 7125
rect 15211 7145 15253 7187
rect 15211 7125 15219 7145
rect 15239 7125 15253 7145
rect 15211 7087 15253 7125
rect 15303 7145 15347 7187
rect 15303 7125 15315 7145
rect 15335 7125 15347 7145
rect 15303 7087 15347 7125
rect 15424 7145 15466 7187
rect 15424 7125 15432 7145
rect 15452 7125 15466 7145
rect 15424 7087 15466 7125
rect 15516 7145 15560 7187
rect 15516 7125 15528 7145
rect 15548 7125 15560 7145
rect 15516 7087 15560 7125
rect 3842 6883 3854 6903
rect 3874 6883 3886 6903
rect 6596 6901 6640 6939
rect 3842 6845 3886 6883
rect 6596 6881 6608 6901
rect 6628 6881 6640 6901
rect 6596 6839 6640 6881
rect 6690 6901 6732 6939
rect 6690 6881 6704 6901
rect 6724 6881 6732 6901
rect 6690 6839 6732 6881
rect 6809 6901 6853 6939
rect 6809 6881 6821 6901
rect 6841 6881 6853 6901
rect 6809 6839 6853 6881
rect 6903 6901 6945 6939
rect 6903 6881 6917 6901
rect 6937 6881 6945 6901
rect 6903 6839 6945 6881
rect 7017 6901 7061 6939
rect 7017 6881 7029 6901
rect 7049 6881 7061 6901
rect 7017 6839 7061 6881
rect 7111 6901 7153 6939
rect 7111 6881 7125 6901
rect 7145 6881 7153 6901
rect 7111 6839 7153 6881
rect 7227 6901 7269 6939
rect 7227 6881 7235 6901
rect 7255 6881 7269 6901
rect 7227 6839 7269 6881
rect 7319 6908 7364 6939
rect 16245 7090 16289 7128
rect 16245 7070 16257 7090
rect 16277 7070 16289 7090
rect 11976 6930 12020 6968
rect 7319 6901 7363 6908
rect 7319 6881 7331 6901
rect 7351 6881 7363 6901
rect 7319 6839 7363 6881
rect 8400 6882 8444 6924
rect 8400 6862 8412 6882
rect 8432 6862 8444 6882
rect 8400 6855 8444 6862
rect 302 6688 346 6726
rect 302 6668 314 6688
rect 334 6668 346 6688
rect 302 6626 346 6668
rect 396 6688 438 6726
rect 396 6668 410 6688
rect 430 6668 438 6688
rect 396 6626 438 6668
rect 515 6688 559 6726
rect 515 6668 527 6688
rect 547 6668 559 6688
rect 515 6626 559 6668
rect 609 6688 651 6726
rect 609 6668 623 6688
rect 643 6668 651 6688
rect 609 6626 651 6668
rect 723 6688 767 6726
rect 723 6668 735 6688
rect 755 6668 767 6688
rect 723 6626 767 6668
rect 817 6688 859 6726
rect 817 6668 831 6688
rect 851 6668 859 6688
rect 817 6626 859 6668
rect 933 6688 975 6726
rect 933 6668 941 6688
rect 961 6668 975 6688
rect 933 6626 975 6668
rect 1025 6695 1070 6726
rect 4131 6722 4175 6764
rect 4131 6702 4143 6722
rect 4163 6702 4175 6722
rect 4131 6695 4175 6702
rect 1025 6688 1069 6695
rect 1025 6668 1037 6688
rect 1057 6668 1069 6688
rect 1025 6626 1069 6668
rect 4130 6664 4175 6695
rect 4225 6722 4267 6764
rect 4225 6702 4239 6722
rect 4259 6702 4267 6722
rect 4225 6664 4267 6702
rect 4341 6722 4383 6764
rect 4341 6702 4349 6722
rect 4369 6702 4383 6722
rect 4341 6664 4383 6702
rect 4433 6722 4477 6764
rect 4433 6702 4445 6722
rect 4465 6702 4477 6722
rect 4433 6664 4477 6702
rect 4549 6722 4591 6764
rect 4549 6702 4557 6722
rect 4577 6702 4591 6722
rect 4549 6664 4591 6702
rect 4641 6722 4685 6764
rect 4641 6702 4653 6722
rect 4673 6702 4685 6722
rect 4641 6664 4685 6702
rect 4762 6722 4804 6764
rect 4762 6702 4770 6722
rect 4790 6702 4804 6722
rect 4762 6664 4804 6702
rect 4854 6722 4898 6764
rect 8399 6824 8444 6855
rect 8494 6882 8536 6924
rect 8494 6862 8508 6882
rect 8528 6862 8536 6882
rect 8494 6824 8536 6862
rect 8610 6882 8652 6924
rect 8610 6862 8618 6882
rect 8638 6862 8652 6882
rect 8610 6824 8652 6862
rect 8702 6882 8746 6924
rect 8702 6862 8714 6882
rect 8734 6862 8746 6882
rect 8702 6824 8746 6862
rect 8818 6882 8860 6924
rect 8818 6862 8826 6882
rect 8846 6862 8860 6882
rect 8818 6824 8860 6862
rect 8910 6882 8954 6924
rect 8910 6862 8922 6882
rect 8942 6862 8954 6882
rect 8910 6824 8954 6862
rect 9031 6882 9073 6924
rect 9031 6862 9039 6882
rect 9059 6862 9073 6882
rect 9031 6824 9073 6862
rect 9123 6882 9167 6924
rect 9123 6862 9135 6882
rect 9155 6862 9167 6882
rect 11976 6910 11988 6930
rect 12008 6910 12020 6930
rect 11976 6868 12020 6910
rect 12070 6930 12112 6968
rect 12070 6910 12084 6930
rect 12104 6910 12112 6930
rect 12070 6868 12112 6910
rect 12189 6930 12233 6968
rect 12189 6910 12201 6930
rect 12221 6910 12233 6930
rect 12189 6868 12233 6910
rect 12283 6930 12325 6968
rect 12283 6910 12297 6930
rect 12317 6910 12325 6930
rect 12283 6868 12325 6910
rect 12397 6930 12441 6968
rect 12397 6910 12409 6930
rect 12429 6910 12441 6930
rect 12397 6868 12441 6910
rect 12491 6930 12533 6968
rect 12491 6910 12505 6930
rect 12525 6910 12533 6930
rect 12491 6868 12533 6910
rect 12607 6930 12649 6968
rect 12607 6910 12615 6930
rect 12635 6910 12649 6930
rect 12607 6868 12649 6910
rect 12699 6937 12744 6968
rect 16245 7028 16289 7070
rect 16339 7090 16381 7128
rect 16339 7070 16353 7090
rect 16373 7070 16381 7090
rect 16339 7028 16381 7070
rect 16458 7090 16502 7128
rect 16458 7070 16470 7090
rect 16490 7070 16502 7090
rect 16458 7028 16502 7070
rect 16552 7090 16594 7128
rect 16552 7070 16566 7090
rect 16586 7070 16594 7090
rect 16552 7028 16594 7070
rect 16666 7090 16710 7128
rect 16666 7070 16678 7090
rect 16698 7070 16710 7090
rect 16666 7028 16710 7070
rect 16760 7090 16802 7128
rect 16760 7070 16774 7090
rect 16794 7070 16802 7090
rect 16760 7028 16802 7070
rect 16876 7090 16918 7128
rect 16876 7070 16884 7090
rect 16904 7070 16918 7090
rect 16876 7028 16918 7070
rect 16968 7097 17013 7128
rect 20074 7124 20118 7166
rect 20074 7104 20086 7124
rect 20106 7104 20118 7124
rect 20074 7097 20118 7104
rect 16968 7090 17012 7097
rect 16968 7070 16980 7090
rect 17000 7070 17012 7090
rect 16968 7028 17012 7070
rect 20073 7066 20118 7097
rect 20168 7124 20210 7166
rect 20168 7104 20182 7124
rect 20202 7104 20210 7124
rect 20168 7066 20210 7104
rect 20284 7124 20326 7166
rect 20284 7104 20292 7124
rect 20312 7104 20326 7124
rect 20284 7066 20326 7104
rect 20376 7124 20420 7166
rect 20376 7104 20388 7124
rect 20408 7104 20420 7124
rect 20376 7066 20420 7104
rect 20492 7124 20534 7166
rect 20492 7104 20500 7124
rect 20520 7104 20534 7124
rect 20492 7066 20534 7104
rect 20584 7124 20628 7166
rect 20584 7104 20596 7124
rect 20616 7104 20628 7124
rect 20584 7066 20628 7104
rect 20705 7124 20747 7166
rect 20705 7104 20713 7124
rect 20733 7104 20747 7124
rect 20705 7066 20747 7104
rect 20797 7124 20841 7166
rect 20797 7104 20809 7124
rect 20829 7104 20841 7124
rect 20797 7066 20841 7104
rect 12699 6930 12743 6937
rect 12699 6910 12711 6930
rect 12731 6910 12743 6930
rect 12699 6868 12743 6910
rect 13780 6911 13824 6953
rect 13780 6891 13792 6911
rect 13812 6891 13824 6911
rect 13780 6884 13824 6891
rect 9123 6824 9167 6862
rect 4854 6702 4866 6722
rect 4886 6702 4898 6722
rect 4854 6664 4898 6702
rect 13779 6853 13824 6884
rect 13874 6911 13916 6953
rect 13874 6891 13888 6911
rect 13908 6891 13916 6911
rect 13874 6853 13916 6891
rect 13990 6911 14032 6953
rect 13990 6891 13998 6911
rect 14018 6891 14032 6911
rect 13990 6853 14032 6891
rect 14082 6911 14126 6953
rect 14082 6891 14094 6911
rect 14114 6891 14126 6911
rect 14082 6853 14126 6891
rect 14198 6911 14240 6953
rect 14198 6891 14206 6911
rect 14226 6891 14240 6911
rect 14198 6853 14240 6891
rect 14290 6911 14334 6953
rect 14290 6891 14302 6911
rect 14322 6891 14334 6911
rect 14290 6853 14334 6891
rect 14411 6911 14453 6953
rect 14411 6891 14419 6911
rect 14439 6891 14453 6911
rect 14411 6853 14453 6891
rect 14503 6911 14547 6953
rect 14503 6891 14515 6911
rect 14535 6891 14547 6911
rect 17257 6909 17301 6947
rect 14503 6853 14547 6891
rect 17257 6889 17269 6909
rect 17289 6889 17301 6909
rect 5583 6667 5627 6705
rect 5583 6647 5595 6667
rect 5615 6647 5627 6667
rect 5583 6605 5627 6647
rect 5677 6667 5719 6705
rect 5677 6647 5691 6667
rect 5711 6647 5719 6667
rect 5677 6605 5719 6647
rect 5796 6667 5840 6705
rect 5796 6647 5808 6667
rect 5828 6647 5840 6667
rect 5796 6605 5840 6647
rect 5890 6667 5932 6705
rect 5890 6647 5904 6667
rect 5924 6647 5932 6667
rect 5890 6605 5932 6647
rect 6004 6667 6048 6705
rect 6004 6647 6016 6667
rect 6036 6647 6048 6667
rect 6004 6605 6048 6647
rect 6098 6667 6140 6705
rect 6098 6647 6112 6667
rect 6132 6647 6140 6667
rect 6098 6605 6140 6647
rect 6214 6667 6256 6705
rect 6214 6647 6222 6667
rect 6242 6647 6256 6667
rect 6214 6605 6256 6647
rect 6306 6674 6351 6705
rect 9412 6701 9456 6743
rect 9412 6681 9424 6701
rect 9444 6681 9456 6701
rect 9412 6674 9456 6681
rect 6306 6667 6350 6674
rect 6306 6647 6318 6667
rect 6338 6647 6350 6667
rect 6306 6605 6350 6647
rect 9411 6643 9456 6674
rect 9506 6701 9548 6743
rect 9506 6681 9520 6701
rect 9540 6681 9548 6701
rect 9506 6643 9548 6681
rect 9622 6701 9664 6743
rect 9622 6681 9630 6701
rect 9650 6681 9664 6701
rect 9622 6643 9664 6681
rect 9714 6701 9758 6743
rect 9714 6681 9726 6701
rect 9746 6681 9758 6701
rect 9714 6643 9758 6681
rect 9830 6701 9872 6743
rect 9830 6681 9838 6701
rect 9858 6681 9872 6701
rect 9830 6643 9872 6681
rect 9922 6701 9966 6743
rect 9922 6681 9934 6701
rect 9954 6681 9966 6701
rect 9922 6643 9966 6681
rect 10043 6701 10085 6743
rect 10043 6681 10051 6701
rect 10071 6681 10085 6701
rect 10043 6643 10085 6681
rect 10135 6701 10179 6743
rect 17257 6847 17301 6889
rect 17351 6909 17393 6947
rect 17351 6889 17365 6909
rect 17385 6889 17393 6909
rect 17351 6847 17393 6889
rect 17470 6909 17514 6947
rect 17470 6889 17482 6909
rect 17502 6889 17514 6909
rect 17470 6847 17514 6889
rect 17564 6909 17606 6947
rect 17564 6889 17578 6909
rect 17598 6889 17606 6909
rect 17564 6847 17606 6889
rect 17678 6909 17722 6947
rect 17678 6889 17690 6909
rect 17710 6889 17722 6909
rect 17678 6847 17722 6889
rect 17772 6909 17814 6947
rect 17772 6889 17786 6909
rect 17806 6889 17814 6909
rect 17772 6847 17814 6889
rect 17888 6909 17930 6947
rect 17888 6889 17896 6909
rect 17916 6889 17930 6909
rect 17888 6847 17930 6889
rect 17980 6916 18025 6947
rect 17980 6909 18024 6916
rect 17980 6889 17992 6909
rect 18012 6889 18024 6909
rect 17980 6847 18024 6889
rect 19061 6890 19105 6932
rect 19061 6870 19073 6890
rect 19093 6870 19105 6890
rect 19061 6863 19105 6870
rect 10135 6681 10147 6701
rect 10167 6681 10179 6701
rect 10135 6643 10179 6681
rect 10963 6696 11007 6734
rect 10963 6676 10975 6696
rect 10995 6676 11007 6696
rect 10963 6634 11007 6676
rect 11057 6696 11099 6734
rect 11057 6676 11071 6696
rect 11091 6676 11099 6696
rect 11057 6634 11099 6676
rect 11176 6696 11220 6734
rect 11176 6676 11188 6696
rect 11208 6676 11220 6696
rect 11176 6634 11220 6676
rect 11270 6696 11312 6734
rect 11270 6676 11284 6696
rect 11304 6676 11312 6696
rect 11270 6634 11312 6676
rect 11384 6696 11428 6734
rect 11384 6676 11396 6696
rect 11416 6676 11428 6696
rect 11384 6634 11428 6676
rect 11478 6696 11520 6734
rect 11478 6676 11492 6696
rect 11512 6676 11520 6696
rect 11478 6634 11520 6676
rect 11594 6696 11636 6734
rect 11594 6676 11602 6696
rect 11622 6676 11636 6696
rect 11594 6634 11636 6676
rect 11686 6703 11731 6734
rect 14792 6730 14836 6772
rect 14792 6710 14804 6730
rect 14824 6710 14836 6730
rect 14792 6703 14836 6710
rect 11686 6696 11730 6703
rect 11686 6676 11698 6696
rect 11718 6676 11730 6696
rect 11686 6634 11730 6676
rect 14791 6672 14836 6703
rect 14886 6730 14928 6772
rect 14886 6710 14900 6730
rect 14920 6710 14928 6730
rect 14886 6672 14928 6710
rect 15002 6730 15044 6772
rect 15002 6710 15010 6730
rect 15030 6710 15044 6730
rect 15002 6672 15044 6710
rect 15094 6730 15138 6772
rect 15094 6710 15106 6730
rect 15126 6710 15138 6730
rect 15094 6672 15138 6710
rect 15210 6730 15252 6772
rect 15210 6710 15218 6730
rect 15238 6710 15252 6730
rect 15210 6672 15252 6710
rect 15302 6730 15346 6772
rect 15302 6710 15314 6730
rect 15334 6710 15346 6730
rect 15302 6672 15346 6710
rect 15423 6730 15465 6772
rect 15423 6710 15431 6730
rect 15451 6710 15465 6730
rect 15423 6672 15465 6710
rect 15515 6730 15559 6772
rect 19060 6832 19105 6863
rect 19155 6890 19197 6932
rect 19155 6870 19169 6890
rect 19189 6870 19197 6890
rect 19155 6832 19197 6870
rect 19271 6890 19313 6932
rect 19271 6870 19279 6890
rect 19299 6870 19313 6890
rect 19271 6832 19313 6870
rect 19363 6890 19407 6932
rect 19363 6870 19375 6890
rect 19395 6870 19407 6890
rect 19363 6832 19407 6870
rect 19479 6890 19521 6932
rect 19479 6870 19487 6890
rect 19507 6870 19521 6890
rect 19479 6832 19521 6870
rect 19571 6890 19615 6932
rect 19571 6870 19583 6890
rect 19603 6870 19615 6890
rect 19571 6832 19615 6870
rect 19692 6890 19734 6932
rect 19692 6870 19700 6890
rect 19720 6870 19734 6890
rect 19692 6832 19734 6870
rect 19784 6890 19828 6932
rect 19784 6870 19796 6890
rect 19816 6870 19828 6890
rect 19784 6832 19828 6870
rect 15515 6710 15527 6730
rect 15547 6710 15559 6730
rect 15515 6672 15559 6710
rect 16244 6675 16288 6713
rect 16244 6655 16256 6675
rect 16276 6655 16288 6675
rect 1530 6410 1574 6448
rect 1530 6390 1542 6410
rect 1562 6390 1574 6410
rect 1530 6348 1574 6390
rect 1624 6410 1666 6448
rect 1624 6390 1638 6410
rect 1658 6390 1666 6410
rect 1624 6348 1666 6390
rect 1743 6410 1787 6448
rect 1743 6390 1755 6410
rect 1775 6390 1787 6410
rect 1743 6348 1787 6390
rect 1837 6410 1879 6448
rect 1837 6390 1851 6410
rect 1871 6390 1879 6410
rect 1837 6348 1879 6390
rect 1951 6410 1995 6448
rect 1951 6390 1963 6410
rect 1983 6390 1995 6410
rect 1951 6348 1995 6390
rect 2045 6410 2087 6448
rect 2045 6390 2059 6410
rect 2079 6390 2087 6410
rect 2045 6348 2087 6390
rect 2161 6410 2203 6448
rect 2161 6390 2169 6410
rect 2189 6390 2203 6410
rect 2161 6348 2203 6390
rect 2253 6417 2298 6448
rect 2911 6436 2955 6478
rect 2253 6410 2297 6417
rect 2253 6390 2265 6410
rect 2285 6390 2297 6410
rect 2911 6416 2923 6436
rect 2943 6416 2955 6436
rect 2911 6409 2955 6416
rect 2253 6348 2297 6390
rect 2910 6378 2955 6409
rect 3005 6436 3047 6478
rect 3005 6416 3019 6436
rect 3039 6416 3047 6436
rect 3005 6378 3047 6416
rect 3121 6436 3163 6478
rect 3121 6416 3129 6436
rect 3149 6416 3163 6436
rect 3121 6378 3163 6416
rect 3213 6436 3257 6478
rect 3213 6416 3225 6436
rect 3245 6416 3257 6436
rect 3213 6378 3257 6416
rect 3329 6436 3371 6478
rect 3329 6416 3337 6436
rect 3357 6416 3371 6436
rect 3329 6378 3371 6416
rect 3421 6436 3465 6478
rect 3421 6416 3433 6436
rect 3453 6416 3465 6436
rect 3421 6378 3465 6416
rect 3542 6436 3584 6478
rect 3542 6416 3550 6436
rect 3570 6416 3584 6436
rect 3542 6378 3584 6416
rect 3634 6436 3678 6478
rect 16244 6613 16288 6655
rect 16338 6675 16380 6713
rect 16338 6655 16352 6675
rect 16372 6655 16380 6675
rect 16338 6613 16380 6655
rect 16457 6675 16501 6713
rect 16457 6655 16469 6675
rect 16489 6655 16501 6675
rect 16457 6613 16501 6655
rect 16551 6675 16593 6713
rect 16551 6655 16565 6675
rect 16585 6655 16593 6675
rect 16551 6613 16593 6655
rect 16665 6675 16709 6713
rect 16665 6655 16677 6675
rect 16697 6655 16709 6675
rect 16665 6613 16709 6655
rect 16759 6675 16801 6713
rect 16759 6655 16773 6675
rect 16793 6655 16801 6675
rect 16759 6613 16801 6655
rect 16875 6675 16917 6713
rect 16875 6655 16883 6675
rect 16903 6655 16917 6675
rect 16875 6613 16917 6655
rect 16967 6682 17012 6713
rect 20073 6709 20117 6751
rect 20073 6689 20085 6709
rect 20105 6689 20117 6709
rect 20073 6682 20117 6689
rect 16967 6675 17011 6682
rect 16967 6655 16979 6675
rect 16999 6655 17011 6675
rect 16967 6613 17011 6655
rect 20072 6651 20117 6682
rect 20167 6709 20209 6751
rect 20167 6689 20181 6709
rect 20201 6689 20209 6709
rect 20167 6651 20209 6689
rect 20283 6709 20325 6751
rect 20283 6689 20291 6709
rect 20311 6689 20325 6709
rect 20283 6651 20325 6689
rect 20375 6709 20419 6751
rect 20375 6689 20387 6709
rect 20407 6689 20419 6709
rect 20375 6651 20419 6689
rect 20491 6709 20533 6751
rect 20491 6689 20499 6709
rect 20519 6689 20533 6709
rect 20491 6651 20533 6689
rect 20583 6709 20627 6751
rect 20583 6689 20595 6709
rect 20615 6689 20627 6709
rect 20583 6651 20627 6689
rect 20704 6709 20746 6751
rect 20704 6689 20712 6709
rect 20732 6689 20746 6709
rect 20704 6651 20746 6689
rect 20796 6709 20840 6751
rect 20796 6689 20808 6709
rect 20828 6689 20840 6709
rect 20796 6651 20840 6689
rect 3634 6416 3646 6436
rect 3666 6416 3678 6436
rect 3634 6378 3678 6416
rect 6811 6389 6855 6427
rect 6811 6369 6823 6389
rect 6843 6369 6855 6389
rect 6811 6327 6855 6369
rect 6905 6389 6947 6427
rect 6905 6369 6919 6389
rect 6939 6369 6947 6389
rect 6905 6327 6947 6369
rect 7024 6389 7068 6427
rect 7024 6369 7036 6389
rect 7056 6369 7068 6389
rect 7024 6327 7068 6369
rect 7118 6389 7160 6427
rect 7118 6369 7132 6389
rect 7152 6369 7160 6389
rect 7118 6327 7160 6369
rect 7232 6389 7276 6427
rect 7232 6369 7244 6389
rect 7264 6369 7276 6389
rect 7232 6327 7276 6369
rect 7326 6389 7368 6427
rect 7326 6369 7340 6389
rect 7360 6369 7368 6389
rect 7326 6327 7368 6369
rect 7442 6389 7484 6427
rect 7442 6369 7450 6389
rect 7470 6369 7484 6389
rect 7442 6327 7484 6369
rect 7534 6396 7579 6427
rect 8192 6415 8236 6457
rect 7534 6389 7578 6396
rect 7534 6369 7546 6389
rect 7566 6369 7578 6389
rect 8192 6395 8204 6415
rect 8224 6395 8236 6415
rect 8192 6388 8236 6395
rect 7534 6327 7578 6369
rect 8191 6357 8236 6388
rect 8286 6415 8328 6457
rect 8286 6395 8300 6415
rect 8320 6395 8328 6415
rect 8286 6357 8328 6395
rect 8402 6415 8444 6457
rect 8402 6395 8410 6415
rect 8430 6395 8444 6415
rect 8402 6357 8444 6395
rect 8494 6415 8538 6457
rect 8494 6395 8506 6415
rect 8526 6395 8538 6415
rect 8494 6357 8538 6395
rect 8610 6415 8652 6457
rect 8610 6395 8618 6415
rect 8638 6395 8652 6415
rect 8610 6357 8652 6395
rect 8702 6415 8746 6457
rect 8702 6395 8714 6415
rect 8734 6395 8746 6415
rect 8702 6357 8746 6395
rect 8823 6415 8865 6457
rect 8823 6395 8831 6415
rect 8851 6395 8865 6415
rect 8823 6357 8865 6395
rect 8915 6415 8959 6457
rect 8915 6395 8927 6415
rect 8947 6395 8959 6415
rect 8915 6357 8959 6395
rect 12191 6418 12235 6456
rect 12191 6398 12203 6418
rect 12223 6398 12235 6418
rect 12191 6356 12235 6398
rect 12285 6418 12327 6456
rect 12285 6398 12299 6418
rect 12319 6398 12327 6418
rect 12285 6356 12327 6398
rect 12404 6418 12448 6456
rect 12404 6398 12416 6418
rect 12436 6398 12448 6418
rect 12404 6356 12448 6398
rect 12498 6418 12540 6456
rect 12498 6398 12512 6418
rect 12532 6398 12540 6418
rect 12498 6356 12540 6398
rect 12612 6418 12656 6456
rect 12612 6398 12624 6418
rect 12644 6398 12656 6418
rect 12612 6356 12656 6398
rect 12706 6418 12748 6456
rect 12706 6398 12720 6418
rect 12740 6398 12748 6418
rect 12706 6356 12748 6398
rect 12822 6418 12864 6456
rect 12822 6398 12830 6418
rect 12850 6398 12864 6418
rect 12822 6356 12864 6398
rect 12914 6425 12959 6456
rect 13572 6444 13616 6486
rect 12914 6418 12958 6425
rect 12914 6398 12926 6418
rect 12946 6398 12958 6418
rect 13572 6424 13584 6444
rect 13604 6424 13616 6444
rect 13572 6417 13616 6424
rect 12914 6356 12958 6398
rect 13571 6386 13616 6417
rect 13666 6444 13708 6486
rect 13666 6424 13680 6444
rect 13700 6424 13708 6444
rect 13666 6386 13708 6424
rect 13782 6444 13824 6486
rect 13782 6424 13790 6444
rect 13810 6424 13824 6444
rect 13782 6386 13824 6424
rect 13874 6444 13918 6486
rect 13874 6424 13886 6444
rect 13906 6424 13918 6444
rect 13874 6386 13918 6424
rect 13990 6444 14032 6486
rect 13990 6424 13998 6444
rect 14018 6424 14032 6444
rect 13990 6386 14032 6424
rect 14082 6444 14126 6486
rect 14082 6424 14094 6444
rect 14114 6424 14126 6444
rect 14082 6386 14126 6424
rect 14203 6444 14245 6486
rect 14203 6424 14211 6444
rect 14231 6424 14245 6444
rect 14203 6386 14245 6424
rect 14295 6444 14339 6486
rect 14295 6424 14307 6444
rect 14327 6424 14339 6444
rect 14295 6386 14339 6424
rect 17472 6397 17516 6435
rect 17472 6377 17484 6397
rect 17504 6377 17516 6397
rect 310 6124 354 6162
rect 310 6104 322 6124
rect 342 6104 354 6124
rect 310 6062 354 6104
rect 404 6124 446 6162
rect 404 6104 418 6124
rect 438 6104 446 6124
rect 404 6062 446 6104
rect 523 6124 567 6162
rect 523 6104 535 6124
rect 555 6104 567 6124
rect 523 6062 567 6104
rect 617 6124 659 6162
rect 617 6104 631 6124
rect 651 6104 659 6124
rect 617 6062 659 6104
rect 731 6124 775 6162
rect 731 6104 743 6124
rect 763 6104 775 6124
rect 731 6062 775 6104
rect 825 6124 867 6162
rect 825 6104 839 6124
rect 859 6104 867 6124
rect 825 6062 867 6104
rect 941 6124 983 6162
rect 941 6104 949 6124
rect 969 6104 983 6124
rect 941 6062 983 6104
rect 1033 6131 1078 6162
rect 4139 6158 4183 6200
rect 4139 6138 4151 6158
rect 4171 6138 4183 6158
rect 4139 6131 4183 6138
rect 1033 6124 1077 6131
rect 1033 6104 1045 6124
rect 1065 6104 1077 6124
rect 1033 6062 1077 6104
rect 4138 6100 4183 6131
rect 4233 6158 4275 6200
rect 4233 6138 4247 6158
rect 4267 6138 4275 6158
rect 4233 6100 4275 6138
rect 4349 6158 4391 6200
rect 4349 6138 4357 6158
rect 4377 6138 4391 6158
rect 4349 6100 4391 6138
rect 4441 6158 4485 6200
rect 4441 6138 4453 6158
rect 4473 6138 4485 6158
rect 4441 6100 4485 6138
rect 4557 6158 4599 6200
rect 4557 6138 4565 6158
rect 4585 6138 4599 6158
rect 4557 6100 4599 6138
rect 4649 6158 4693 6200
rect 4649 6138 4661 6158
rect 4681 6138 4693 6158
rect 4649 6100 4693 6138
rect 4770 6158 4812 6200
rect 4770 6138 4778 6158
rect 4798 6138 4812 6158
rect 4770 6100 4812 6138
rect 4862 6158 4906 6200
rect 17472 6335 17516 6377
rect 17566 6397 17608 6435
rect 17566 6377 17580 6397
rect 17600 6377 17608 6397
rect 17566 6335 17608 6377
rect 17685 6397 17729 6435
rect 17685 6377 17697 6397
rect 17717 6377 17729 6397
rect 17685 6335 17729 6377
rect 17779 6397 17821 6435
rect 17779 6377 17793 6397
rect 17813 6377 17821 6397
rect 17779 6335 17821 6377
rect 17893 6397 17937 6435
rect 17893 6377 17905 6397
rect 17925 6377 17937 6397
rect 17893 6335 17937 6377
rect 17987 6397 18029 6435
rect 17987 6377 18001 6397
rect 18021 6377 18029 6397
rect 17987 6335 18029 6377
rect 18103 6397 18145 6435
rect 18103 6377 18111 6397
rect 18131 6377 18145 6397
rect 18103 6335 18145 6377
rect 18195 6404 18240 6435
rect 18853 6423 18897 6465
rect 18195 6397 18239 6404
rect 18195 6377 18207 6397
rect 18227 6377 18239 6397
rect 18853 6403 18865 6423
rect 18885 6403 18897 6423
rect 18853 6396 18897 6403
rect 18195 6335 18239 6377
rect 18852 6365 18897 6396
rect 18947 6423 18989 6465
rect 18947 6403 18961 6423
rect 18981 6403 18989 6423
rect 18947 6365 18989 6403
rect 19063 6423 19105 6465
rect 19063 6403 19071 6423
rect 19091 6403 19105 6423
rect 19063 6365 19105 6403
rect 19155 6423 19199 6465
rect 19155 6403 19167 6423
rect 19187 6403 19199 6423
rect 19155 6365 19199 6403
rect 19271 6423 19313 6465
rect 19271 6403 19279 6423
rect 19299 6403 19313 6423
rect 19271 6365 19313 6403
rect 19363 6423 19407 6465
rect 19363 6403 19375 6423
rect 19395 6403 19407 6423
rect 19363 6365 19407 6403
rect 19484 6423 19526 6465
rect 19484 6403 19492 6423
rect 19512 6403 19526 6423
rect 19484 6365 19526 6403
rect 19576 6423 19620 6465
rect 19576 6403 19588 6423
rect 19608 6403 19620 6423
rect 19576 6365 19620 6403
rect 4862 6138 4874 6158
rect 4894 6138 4906 6158
rect 4862 6100 4906 6138
rect 5591 6103 5635 6141
rect 5591 6083 5603 6103
rect 5623 6083 5635 6103
rect 1322 5943 1366 5981
rect 1322 5923 1334 5943
rect 1354 5923 1366 5943
rect 1322 5881 1366 5923
rect 1416 5943 1458 5981
rect 1416 5923 1430 5943
rect 1450 5923 1458 5943
rect 1416 5881 1458 5923
rect 1535 5943 1579 5981
rect 1535 5923 1547 5943
rect 1567 5923 1579 5943
rect 1535 5881 1579 5923
rect 1629 5943 1671 5981
rect 1629 5923 1643 5943
rect 1663 5923 1671 5943
rect 1629 5881 1671 5923
rect 1743 5943 1787 5981
rect 1743 5923 1755 5943
rect 1775 5923 1787 5943
rect 1743 5881 1787 5923
rect 1837 5943 1879 5981
rect 1837 5923 1851 5943
rect 1871 5923 1879 5943
rect 1837 5881 1879 5923
rect 1953 5943 1995 5981
rect 1953 5923 1961 5943
rect 1981 5923 1995 5943
rect 1953 5881 1995 5923
rect 2045 5950 2090 5981
rect 5591 6041 5635 6083
rect 5685 6103 5727 6141
rect 5685 6083 5699 6103
rect 5719 6083 5727 6103
rect 5685 6041 5727 6083
rect 5804 6103 5848 6141
rect 5804 6083 5816 6103
rect 5836 6083 5848 6103
rect 5804 6041 5848 6083
rect 5898 6103 5940 6141
rect 5898 6083 5912 6103
rect 5932 6083 5940 6103
rect 5898 6041 5940 6083
rect 6012 6103 6056 6141
rect 6012 6083 6024 6103
rect 6044 6083 6056 6103
rect 6012 6041 6056 6083
rect 6106 6103 6148 6141
rect 6106 6083 6120 6103
rect 6140 6083 6148 6103
rect 6106 6041 6148 6083
rect 6222 6103 6264 6141
rect 6222 6083 6230 6103
rect 6250 6083 6264 6103
rect 6222 6041 6264 6083
rect 6314 6110 6359 6141
rect 9420 6137 9464 6179
rect 9420 6117 9432 6137
rect 9452 6117 9464 6137
rect 9420 6110 9464 6117
rect 6314 6103 6358 6110
rect 6314 6083 6326 6103
rect 6346 6083 6358 6103
rect 6314 6041 6358 6083
rect 9419 6079 9464 6110
rect 9514 6137 9556 6179
rect 9514 6117 9528 6137
rect 9548 6117 9556 6137
rect 9514 6079 9556 6117
rect 9630 6137 9672 6179
rect 9630 6117 9638 6137
rect 9658 6117 9672 6137
rect 9630 6079 9672 6117
rect 9722 6137 9766 6179
rect 9722 6117 9734 6137
rect 9754 6117 9766 6137
rect 9722 6079 9766 6117
rect 9838 6137 9880 6179
rect 9838 6117 9846 6137
rect 9866 6117 9880 6137
rect 9838 6079 9880 6117
rect 9930 6137 9974 6179
rect 9930 6117 9942 6137
rect 9962 6117 9974 6137
rect 9930 6079 9974 6117
rect 10051 6137 10093 6179
rect 10051 6117 10059 6137
rect 10079 6117 10093 6137
rect 10051 6079 10093 6117
rect 10143 6137 10187 6179
rect 10143 6117 10155 6137
rect 10175 6117 10187 6137
rect 10143 6079 10187 6117
rect 10971 6132 11015 6170
rect 10971 6112 10983 6132
rect 11003 6112 11015 6132
rect 2045 5943 2089 5950
rect 2045 5923 2057 5943
rect 2077 5923 2089 5943
rect 2045 5881 2089 5923
rect 3126 5924 3170 5966
rect 3126 5904 3138 5924
rect 3158 5904 3170 5924
rect 3126 5897 3170 5904
rect 3125 5866 3170 5897
rect 3220 5924 3262 5966
rect 3220 5904 3234 5924
rect 3254 5904 3262 5924
rect 3220 5866 3262 5904
rect 3336 5924 3378 5966
rect 3336 5904 3344 5924
rect 3364 5904 3378 5924
rect 3336 5866 3378 5904
rect 3428 5924 3472 5966
rect 3428 5904 3440 5924
rect 3460 5904 3472 5924
rect 3428 5866 3472 5904
rect 3544 5924 3586 5966
rect 3544 5904 3552 5924
rect 3572 5904 3586 5924
rect 3544 5866 3586 5904
rect 3636 5924 3680 5966
rect 3636 5904 3648 5924
rect 3668 5904 3680 5924
rect 3636 5866 3680 5904
rect 3757 5924 3799 5966
rect 3757 5904 3765 5924
rect 3785 5904 3799 5924
rect 3757 5866 3799 5904
rect 3849 5924 3893 5966
rect 10971 6070 11015 6112
rect 11065 6132 11107 6170
rect 11065 6112 11079 6132
rect 11099 6112 11107 6132
rect 11065 6070 11107 6112
rect 11184 6132 11228 6170
rect 11184 6112 11196 6132
rect 11216 6112 11228 6132
rect 11184 6070 11228 6112
rect 11278 6132 11320 6170
rect 11278 6112 11292 6132
rect 11312 6112 11320 6132
rect 11278 6070 11320 6112
rect 11392 6132 11436 6170
rect 11392 6112 11404 6132
rect 11424 6112 11436 6132
rect 11392 6070 11436 6112
rect 11486 6132 11528 6170
rect 11486 6112 11500 6132
rect 11520 6112 11528 6132
rect 11486 6070 11528 6112
rect 11602 6132 11644 6170
rect 11602 6112 11610 6132
rect 11630 6112 11644 6132
rect 11602 6070 11644 6112
rect 11694 6139 11739 6170
rect 14800 6166 14844 6208
rect 14800 6146 14812 6166
rect 14832 6146 14844 6166
rect 14800 6139 14844 6146
rect 11694 6132 11738 6139
rect 11694 6112 11706 6132
rect 11726 6112 11738 6132
rect 11694 6070 11738 6112
rect 14799 6108 14844 6139
rect 14894 6166 14936 6208
rect 14894 6146 14908 6166
rect 14928 6146 14936 6166
rect 14894 6108 14936 6146
rect 15010 6166 15052 6208
rect 15010 6146 15018 6166
rect 15038 6146 15052 6166
rect 15010 6108 15052 6146
rect 15102 6166 15146 6208
rect 15102 6146 15114 6166
rect 15134 6146 15146 6166
rect 15102 6108 15146 6146
rect 15218 6166 15260 6208
rect 15218 6146 15226 6166
rect 15246 6146 15260 6166
rect 15218 6108 15260 6146
rect 15310 6166 15354 6208
rect 15310 6146 15322 6166
rect 15342 6146 15354 6166
rect 15310 6108 15354 6146
rect 15431 6166 15473 6208
rect 15431 6146 15439 6166
rect 15459 6146 15473 6166
rect 15431 6108 15473 6146
rect 15523 6166 15567 6208
rect 15523 6146 15535 6166
rect 15555 6146 15567 6166
rect 15523 6108 15567 6146
rect 3849 5904 3861 5924
rect 3881 5904 3893 5924
rect 6603 5922 6647 5960
rect 3849 5866 3893 5904
rect 6603 5902 6615 5922
rect 6635 5902 6647 5922
rect 6603 5860 6647 5902
rect 6697 5922 6739 5960
rect 6697 5902 6711 5922
rect 6731 5902 6739 5922
rect 6697 5860 6739 5902
rect 6816 5922 6860 5960
rect 6816 5902 6828 5922
rect 6848 5902 6860 5922
rect 6816 5860 6860 5902
rect 6910 5922 6952 5960
rect 6910 5902 6924 5922
rect 6944 5902 6952 5922
rect 6910 5860 6952 5902
rect 7024 5922 7068 5960
rect 7024 5902 7036 5922
rect 7056 5902 7068 5922
rect 7024 5860 7068 5902
rect 7118 5922 7160 5960
rect 7118 5902 7132 5922
rect 7152 5902 7160 5922
rect 7118 5860 7160 5902
rect 7234 5922 7276 5960
rect 7234 5902 7242 5922
rect 7262 5902 7276 5922
rect 7234 5860 7276 5902
rect 7326 5929 7371 5960
rect 16252 6111 16296 6149
rect 16252 6091 16264 6111
rect 16284 6091 16296 6111
rect 11983 5951 12027 5989
rect 7326 5922 7370 5929
rect 7326 5902 7338 5922
rect 7358 5902 7370 5922
rect 7326 5860 7370 5902
rect 8407 5903 8451 5945
rect 8407 5883 8419 5903
rect 8439 5883 8451 5903
rect 8407 5876 8451 5883
rect 309 5709 353 5747
rect 309 5689 321 5709
rect 341 5689 353 5709
rect 309 5647 353 5689
rect 403 5709 445 5747
rect 403 5689 417 5709
rect 437 5689 445 5709
rect 403 5647 445 5689
rect 522 5709 566 5747
rect 522 5689 534 5709
rect 554 5689 566 5709
rect 522 5647 566 5689
rect 616 5709 658 5747
rect 616 5689 630 5709
rect 650 5689 658 5709
rect 616 5647 658 5689
rect 730 5709 774 5747
rect 730 5689 742 5709
rect 762 5689 774 5709
rect 730 5647 774 5689
rect 824 5709 866 5747
rect 824 5689 838 5709
rect 858 5689 866 5709
rect 824 5647 866 5689
rect 940 5709 982 5747
rect 940 5689 948 5709
rect 968 5689 982 5709
rect 940 5647 982 5689
rect 1032 5716 1077 5747
rect 4138 5743 4182 5785
rect 4138 5723 4150 5743
rect 4170 5723 4182 5743
rect 4138 5716 4182 5723
rect 1032 5709 1076 5716
rect 1032 5689 1044 5709
rect 1064 5689 1076 5709
rect 1032 5647 1076 5689
rect 4137 5685 4182 5716
rect 4232 5743 4274 5785
rect 4232 5723 4246 5743
rect 4266 5723 4274 5743
rect 4232 5685 4274 5723
rect 4348 5743 4390 5785
rect 4348 5723 4356 5743
rect 4376 5723 4390 5743
rect 4348 5685 4390 5723
rect 4440 5743 4484 5785
rect 4440 5723 4452 5743
rect 4472 5723 4484 5743
rect 4440 5685 4484 5723
rect 4556 5743 4598 5785
rect 4556 5723 4564 5743
rect 4584 5723 4598 5743
rect 4556 5685 4598 5723
rect 4648 5743 4692 5785
rect 4648 5723 4660 5743
rect 4680 5723 4692 5743
rect 4648 5685 4692 5723
rect 4769 5743 4811 5785
rect 4769 5723 4777 5743
rect 4797 5723 4811 5743
rect 4769 5685 4811 5723
rect 4861 5743 4905 5785
rect 8406 5845 8451 5876
rect 8501 5903 8543 5945
rect 8501 5883 8515 5903
rect 8535 5883 8543 5903
rect 8501 5845 8543 5883
rect 8617 5903 8659 5945
rect 8617 5883 8625 5903
rect 8645 5883 8659 5903
rect 8617 5845 8659 5883
rect 8709 5903 8753 5945
rect 8709 5883 8721 5903
rect 8741 5883 8753 5903
rect 8709 5845 8753 5883
rect 8825 5903 8867 5945
rect 8825 5883 8833 5903
rect 8853 5883 8867 5903
rect 8825 5845 8867 5883
rect 8917 5903 8961 5945
rect 8917 5883 8929 5903
rect 8949 5883 8961 5903
rect 8917 5845 8961 5883
rect 9038 5903 9080 5945
rect 9038 5883 9046 5903
rect 9066 5883 9080 5903
rect 9038 5845 9080 5883
rect 9130 5903 9174 5945
rect 9130 5883 9142 5903
rect 9162 5883 9174 5903
rect 11983 5931 11995 5951
rect 12015 5931 12027 5951
rect 11983 5889 12027 5931
rect 12077 5951 12119 5989
rect 12077 5931 12091 5951
rect 12111 5931 12119 5951
rect 12077 5889 12119 5931
rect 12196 5951 12240 5989
rect 12196 5931 12208 5951
rect 12228 5931 12240 5951
rect 12196 5889 12240 5931
rect 12290 5951 12332 5989
rect 12290 5931 12304 5951
rect 12324 5931 12332 5951
rect 12290 5889 12332 5931
rect 12404 5951 12448 5989
rect 12404 5931 12416 5951
rect 12436 5931 12448 5951
rect 12404 5889 12448 5931
rect 12498 5951 12540 5989
rect 12498 5931 12512 5951
rect 12532 5931 12540 5951
rect 12498 5889 12540 5931
rect 12614 5951 12656 5989
rect 12614 5931 12622 5951
rect 12642 5931 12656 5951
rect 12614 5889 12656 5931
rect 12706 5958 12751 5989
rect 16252 6049 16296 6091
rect 16346 6111 16388 6149
rect 16346 6091 16360 6111
rect 16380 6091 16388 6111
rect 16346 6049 16388 6091
rect 16465 6111 16509 6149
rect 16465 6091 16477 6111
rect 16497 6091 16509 6111
rect 16465 6049 16509 6091
rect 16559 6111 16601 6149
rect 16559 6091 16573 6111
rect 16593 6091 16601 6111
rect 16559 6049 16601 6091
rect 16673 6111 16717 6149
rect 16673 6091 16685 6111
rect 16705 6091 16717 6111
rect 16673 6049 16717 6091
rect 16767 6111 16809 6149
rect 16767 6091 16781 6111
rect 16801 6091 16809 6111
rect 16767 6049 16809 6091
rect 16883 6111 16925 6149
rect 16883 6091 16891 6111
rect 16911 6091 16925 6111
rect 16883 6049 16925 6091
rect 16975 6118 17020 6149
rect 20081 6145 20125 6187
rect 20081 6125 20093 6145
rect 20113 6125 20125 6145
rect 20081 6118 20125 6125
rect 16975 6111 17019 6118
rect 16975 6091 16987 6111
rect 17007 6091 17019 6111
rect 16975 6049 17019 6091
rect 20080 6087 20125 6118
rect 20175 6145 20217 6187
rect 20175 6125 20189 6145
rect 20209 6125 20217 6145
rect 20175 6087 20217 6125
rect 20291 6145 20333 6187
rect 20291 6125 20299 6145
rect 20319 6125 20333 6145
rect 20291 6087 20333 6125
rect 20383 6145 20427 6187
rect 20383 6125 20395 6145
rect 20415 6125 20427 6145
rect 20383 6087 20427 6125
rect 20499 6145 20541 6187
rect 20499 6125 20507 6145
rect 20527 6125 20541 6145
rect 20499 6087 20541 6125
rect 20591 6145 20635 6187
rect 20591 6125 20603 6145
rect 20623 6125 20635 6145
rect 20591 6087 20635 6125
rect 20712 6145 20754 6187
rect 20712 6125 20720 6145
rect 20740 6125 20754 6145
rect 20712 6087 20754 6125
rect 20804 6145 20848 6187
rect 20804 6125 20816 6145
rect 20836 6125 20848 6145
rect 20804 6087 20848 6125
rect 12706 5951 12750 5958
rect 12706 5931 12718 5951
rect 12738 5931 12750 5951
rect 12706 5889 12750 5931
rect 13787 5932 13831 5974
rect 13787 5912 13799 5932
rect 13819 5912 13831 5932
rect 13787 5905 13831 5912
rect 9130 5845 9174 5883
rect 4861 5723 4873 5743
rect 4893 5723 4905 5743
rect 4861 5685 4905 5723
rect 13786 5874 13831 5905
rect 13881 5932 13923 5974
rect 13881 5912 13895 5932
rect 13915 5912 13923 5932
rect 13881 5874 13923 5912
rect 13997 5932 14039 5974
rect 13997 5912 14005 5932
rect 14025 5912 14039 5932
rect 13997 5874 14039 5912
rect 14089 5932 14133 5974
rect 14089 5912 14101 5932
rect 14121 5912 14133 5932
rect 14089 5874 14133 5912
rect 14205 5932 14247 5974
rect 14205 5912 14213 5932
rect 14233 5912 14247 5932
rect 14205 5874 14247 5912
rect 14297 5932 14341 5974
rect 14297 5912 14309 5932
rect 14329 5912 14341 5932
rect 14297 5874 14341 5912
rect 14418 5932 14460 5974
rect 14418 5912 14426 5932
rect 14446 5912 14460 5932
rect 14418 5874 14460 5912
rect 14510 5932 14554 5974
rect 14510 5912 14522 5932
rect 14542 5912 14554 5932
rect 17264 5930 17308 5968
rect 14510 5874 14554 5912
rect 17264 5910 17276 5930
rect 17296 5910 17308 5930
rect 5590 5688 5634 5726
rect 5590 5668 5602 5688
rect 5622 5668 5634 5688
rect 5590 5626 5634 5668
rect 5684 5688 5726 5726
rect 5684 5668 5698 5688
rect 5718 5668 5726 5688
rect 5684 5626 5726 5668
rect 5803 5688 5847 5726
rect 5803 5668 5815 5688
rect 5835 5668 5847 5688
rect 5803 5626 5847 5668
rect 5897 5688 5939 5726
rect 5897 5668 5911 5688
rect 5931 5668 5939 5688
rect 5897 5626 5939 5668
rect 6011 5688 6055 5726
rect 6011 5668 6023 5688
rect 6043 5668 6055 5688
rect 6011 5626 6055 5668
rect 6105 5688 6147 5726
rect 6105 5668 6119 5688
rect 6139 5668 6147 5688
rect 6105 5626 6147 5668
rect 6221 5688 6263 5726
rect 6221 5668 6229 5688
rect 6249 5668 6263 5688
rect 6221 5626 6263 5668
rect 6313 5695 6358 5726
rect 9419 5722 9463 5764
rect 9419 5702 9431 5722
rect 9451 5702 9463 5722
rect 9419 5695 9463 5702
rect 6313 5688 6357 5695
rect 6313 5668 6325 5688
rect 6345 5668 6357 5688
rect 6313 5626 6357 5668
rect 9418 5664 9463 5695
rect 9513 5722 9555 5764
rect 9513 5702 9527 5722
rect 9547 5702 9555 5722
rect 9513 5664 9555 5702
rect 9629 5722 9671 5764
rect 9629 5702 9637 5722
rect 9657 5702 9671 5722
rect 9629 5664 9671 5702
rect 9721 5722 9765 5764
rect 9721 5702 9733 5722
rect 9753 5702 9765 5722
rect 9721 5664 9765 5702
rect 9837 5722 9879 5764
rect 9837 5702 9845 5722
rect 9865 5702 9879 5722
rect 9837 5664 9879 5702
rect 9929 5722 9973 5764
rect 9929 5702 9941 5722
rect 9961 5702 9973 5722
rect 9929 5664 9973 5702
rect 10050 5722 10092 5764
rect 10050 5702 10058 5722
rect 10078 5702 10092 5722
rect 10050 5664 10092 5702
rect 10142 5722 10186 5764
rect 17264 5868 17308 5910
rect 17358 5930 17400 5968
rect 17358 5910 17372 5930
rect 17392 5910 17400 5930
rect 17358 5868 17400 5910
rect 17477 5930 17521 5968
rect 17477 5910 17489 5930
rect 17509 5910 17521 5930
rect 17477 5868 17521 5910
rect 17571 5930 17613 5968
rect 17571 5910 17585 5930
rect 17605 5910 17613 5930
rect 17571 5868 17613 5910
rect 17685 5930 17729 5968
rect 17685 5910 17697 5930
rect 17717 5910 17729 5930
rect 17685 5868 17729 5910
rect 17779 5930 17821 5968
rect 17779 5910 17793 5930
rect 17813 5910 17821 5930
rect 17779 5868 17821 5910
rect 17895 5930 17937 5968
rect 17895 5910 17903 5930
rect 17923 5910 17937 5930
rect 17895 5868 17937 5910
rect 17987 5937 18032 5968
rect 17987 5930 18031 5937
rect 17987 5910 17999 5930
rect 18019 5910 18031 5930
rect 17987 5868 18031 5910
rect 19068 5911 19112 5953
rect 19068 5891 19080 5911
rect 19100 5891 19112 5911
rect 19068 5884 19112 5891
rect 10142 5702 10154 5722
rect 10174 5702 10186 5722
rect 10142 5664 10186 5702
rect 10970 5717 11014 5755
rect 10970 5697 10982 5717
rect 11002 5697 11014 5717
rect 10970 5655 11014 5697
rect 11064 5717 11106 5755
rect 11064 5697 11078 5717
rect 11098 5697 11106 5717
rect 11064 5655 11106 5697
rect 11183 5717 11227 5755
rect 11183 5697 11195 5717
rect 11215 5697 11227 5717
rect 11183 5655 11227 5697
rect 11277 5717 11319 5755
rect 11277 5697 11291 5717
rect 11311 5697 11319 5717
rect 11277 5655 11319 5697
rect 11391 5717 11435 5755
rect 11391 5697 11403 5717
rect 11423 5697 11435 5717
rect 11391 5655 11435 5697
rect 11485 5717 11527 5755
rect 11485 5697 11499 5717
rect 11519 5697 11527 5717
rect 11485 5655 11527 5697
rect 11601 5717 11643 5755
rect 11601 5697 11609 5717
rect 11629 5697 11643 5717
rect 11601 5655 11643 5697
rect 11693 5724 11738 5755
rect 14799 5751 14843 5793
rect 14799 5731 14811 5751
rect 14831 5731 14843 5751
rect 14799 5724 14843 5731
rect 11693 5717 11737 5724
rect 11693 5697 11705 5717
rect 11725 5697 11737 5717
rect 11693 5655 11737 5697
rect 14798 5693 14843 5724
rect 14893 5751 14935 5793
rect 14893 5731 14907 5751
rect 14927 5731 14935 5751
rect 14893 5693 14935 5731
rect 15009 5751 15051 5793
rect 15009 5731 15017 5751
rect 15037 5731 15051 5751
rect 15009 5693 15051 5731
rect 15101 5751 15145 5793
rect 15101 5731 15113 5751
rect 15133 5731 15145 5751
rect 15101 5693 15145 5731
rect 15217 5751 15259 5793
rect 15217 5731 15225 5751
rect 15245 5731 15259 5751
rect 15217 5693 15259 5731
rect 15309 5751 15353 5793
rect 15309 5731 15321 5751
rect 15341 5731 15353 5751
rect 15309 5693 15353 5731
rect 15430 5751 15472 5793
rect 15430 5731 15438 5751
rect 15458 5731 15472 5751
rect 15430 5693 15472 5731
rect 15522 5751 15566 5793
rect 19067 5853 19112 5884
rect 19162 5911 19204 5953
rect 19162 5891 19176 5911
rect 19196 5891 19204 5911
rect 19162 5853 19204 5891
rect 19278 5911 19320 5953
rect 19278 5891 19286 5911
rect 19306 5891 19320 5911
rect 19278 5853 19320 5891
rect 19370 5911 19414 5953
rect 19370 5891 19382 5911
rect 19402 5891 19414 5911
rect 19370 5853 19414 5891
rect 19486 5911 19528 5953
rect 19486 5891 19494 5911
rect 19514 5891 19528 5911
rect 19486 5853 19528 5891
rect 19578 5911 19622 5953
rect 19578 5891 19590 5911
rect 19610 5891 19622 5911
rect 19578 5853 19622 5891
rect 19699 5911 19741 5953
rect 19699 5891 19707 5911
rect 19727 5891 19741 5911
rect 19699 5853 19741 5891
rect 19791 5911 19835 5953
rect 19791 5891 19803 5911
rect 19823 5891 19835 5911
rect 19791 5853 19835 5891
rect 15522 5731 15534 5751
rect 15554 5731 15566 5751
rect 15522 5693 15566 5731
rect 16251 5696 16295 5734
rect 16251 5676 16263 5696
rect 16283 5676 16295 5696
rect 3076 5504 3120 5546
rect 3076 5484 3088 5504
rect 3108 5484 3120 5504
rect 3076 5477 3120 5484
rect 3075 5446 3120 5477
rect 3170 5504 3212 5546
rect 3170 5484 3184 5504
rect 3204 5484 3212 5504
rect 3170 5446 3212 5484
rect 3286 5504 3328 5546
rect 3286 5484 3294 5504
rect 3314 5484 3328 5504
rect 3286 5446 3328 5484
rect 3378 5504 3422 5546
rect 3378 5484 3390 5504
rect 3410 5484 3422 5504
rect 3378 5446 3422 5484
rect 3494 5504 3536 5546
rect 3494 5484 3502 5504
rect 3522 5484 3536 5504
rect 3494 5446 3536 5484
rect 3586 5504 3630 5546
rect 3586 5484 3598 5504
rect 3618 5484 3630 5504
rect 3586 5446 3630 5484
rect 3707 5504 3749 5546
rect 3707 5484 3715 5504
rect 3735 5484 3749 5504
rect 3707 5446 3749 5484
rect 3799 5504 3843 5546
rect 3799 5484 3811 5504
rect 3831 5484 3843 5504
rect 3799 5446 3843 5484
rect 8357 5483 8401 5525
rect 8357 5463 8369 5483
rect 8389 5463 8401 5483
rect 8357 5456 8401 5463
rect 8356 5425 8401 5456
rect 8451 5483 8493 5525
rect 8451 5463 8465 5483
rect 8485 5463 8493 5483
rect 8451 5425 8493 5463
rect 8567 5483 8609 5525
rect 8567 5463 8575 5483
rect 8595 5463 8609 5483
rect 8567 5425 8609 5463
rect 8659 5483 8703 5525
rect 8659 5463 8671 5483
rect 8691 5463 8703 5483
rect 8659 5425 8703 5463
rect 8775 5483 8817 5525
rect 8775 5463 8783 5483
rect 8803 5463 8817 5483
rect 8775 5425 8817 5463
rect 8867 5483 8911 5525
rect 8867 5463 8879 5483
rect 8899 5463 8911 5483
rect 8867 5425 8911 5463
rect 8988 5483 9030 5525
rect 8988 5463 8996 5483
rect 9016 5463 9030 5483
rect 8988 5425 9030 5463
rect 9080 5483 9124 5525
rect 16251 5634 16295 5676
rect 16345 5696 16387 5734
rect 16345 5676 16359 5696
rect 16379 5676 16387 5696
rect 16345 5634 16387 5676
rect 16464 5696 16508 5734
rect 16464 5676 16476 5696
rect 16496 5676 16508 5696
rect 16464 5634 16508 5676
rect 16558 5696 16600 5734
rect 16558 5676 16572 5696
rect 16592 5676 16600 5696
rect 16558 5634 16600 5676
rect 16672 5696 16716 5734
rect 16672 5676 16684 5696
rect 16704 5676 16716 5696
rect 16672 5634 16716 5676
rect 16766 5696 16808 5734
rect 16766 5676 16780 5696
rect 16800 5676 16808 5696
rect 16766 5634 16808 5676
rect 16882 5696 16924 5734
rect 16882 5676 16890 5696
rect 16910 5676 16924 5696
rect 16882 5634 16924 5676
rect 16974 5703 17019 5734
rect 20080 5730 20124 5772
rect 20080 5710 20092 5730
rect 20112 5710 20124 5730
rect 20080 5703 20124 5710
rect 16974 5696 17018 5703
rect 16974 5676 16986 5696
rect 17006 5676 17018 5696
rect 16974 5634 17018 5676
rect 20079 5672 20124 5703
rect 20174 5730 20216 5772
rect 20174 5710 20188 5730
rect 20208 5710 20216 5730
rect 20174 5672 20216 5710
rect 20290 5730 20332 5772
rect 20290 5710 20298 5730
rect 20318 5710 20332 5730
rect 20290 5672 20332 5710
rect 20382 5730 20426 5772
rect 20382 5710 20394 5730
rect 20414 5710 20426 5730
rect 20382 5672 20426 5710
rect 20498 5730 20540 5772
rect 20498 5710 20506 5730
rect 20526 5710 20540 5730
rect 20498 5672 20540 5710
rect 20590 5730 20634 5772
rect 20590 5710 20602 5730
rect 20622 5710 20634 5730
rect 20590 5672 20634 5710
rect 20711 5730 20753 5772
rect 20711 5710 20719 5730
rect 20739 5710 20753 5730
rect 20711 5672 20753 5710
rect 20803 5730 20847 5772
rect 20803 5710 20815 5730
rect 20835 5710 20847 5730
rect 20803 5672 20847 5710
rect 9080 5463 9092 5483
rect 9112 5463 9124 5483
rect 9080 5425 9124 5463
rect 13737 5512 13781 5554
rect 13737 5492 13749 5512
rect 13769 5492 13781 5512
rect 13737 5485 13781 5492
rect 13736 5454 13781 5485
rect 13831 5512 13873 5554
rect 13831 5492 13845 5512
rect 13865 5492 13873 5512
rect 13831 5454 13873 5492
rect 13947 5512 13989 5554
rect 13947 5492 13955 5512
rect 13975 5492 13989 5512
rect 13947 5454 13989 5492
rect 14039 5512 14083 5554
rect 14039 5492 14051 5512
rect 14071 5492 14083 5512
rect 14039 5454 14083 5492
rect 14155 5512 14197 5554
rect 14155 5492 14163 5512
rect 14183 5492 14197 5512
rect 14155 5454 14197 5492
rect 14247 5512 14291 5554
rect 14247 5492 14259 5512
rect 14279 5492 14291 5512
rect 14247 5454 14291 5492
rect 14368 5512 14410 5554
rect 14368 5492 14376 5512
rect 14396 5492 14410 5512
rect 14368 5454 14410 5492
rect 14460 5512 14504 5554
rect 14460 5492 14472 5512
rect 14492 5492 14504 5512
rect 14460 5454 14504 5492
rect 19018 5491 19062 5533
rect 19018 5471 19030 5491
rect 19050 5471 19062 5491
rect 19018 5464 19062 5471
rect 19017 5433 19062 5464
rect 19112 5491 19154 5533
rect 19112 5471 19126 5491
rect 19146 5471 19154 5491
rect 19112 5433 19154 5471
rect 19228 5491 19270 5533
rect 19228 5471 19236 5491
rect 19256 5471 19270 5491
rect 19228 5433 19270 5471
rect 19320 5491 19364 5533
rect 19320 5471 19332 5491
rect 19352 5471 19364 5491
rect 19320 5433 19364 5471
rect 19436 5491 19478 5533
rect 19436 5471 19444 5491
rect 19464 5471 19478 5491
rect 19436 5433 19478 5471
rect 19528 5491 19572 5533
rect 19528 5471 19540 5491
rect 19560 5471 19572 5491
rect 19528 5433 19572 5471
rect 19649 5491 19691 5533
rect 19649 5471 19657 5491
rect 19677 5471 19691 5491
rect 19649 5433 19691 5471
rect 19741 5491 19785 5533
rect 19741 5471 19753 5491
rect 19773 5471 19785 5491
rect 19741 5433 19785 5471
rect 1377 5382 1421 5420
rect 1377 5362 1389 5382
rect 1409 5362 1421 5382
rect 1377 5320 1421 5362
rect 1471 5382 1513 5420
rect 1471 5362 1485 5382
rect 1505 5362 1513 5382
rect 1471 5320 1513 5362
rect 1590 5382 1634 5420
rect 1590 5362 1602 5382
rect 1622 5362 1634 5382
rect 1590 5320 1634 5362
rect 1684 5382 1726 5420
rect 1684 5362 1698 5382
rect 1718 5362 1726 5382
rect 1684 5320 1726 5362
rect 1798 5382 1842 5420
rect 1798 5362 1810 5382
rect 1830 5362 1842 5382
rect 1798 5320 1842 5362
rect 1892 5382 1934 5420
rect 1892 5362 1906 5382
rect 1926 5362 1934 5382
rect 1892 5320 1934 5362
rect 2008 5382 2050 5420
rect 2008 5362 2016 5382
rect 2036 5362 2050 5382
rect 2008 5320 2050 5362
rect 2100 5389 2145 5420
rect 2100 5382 2144 5389
rect 2100 5362 2112 5382
rect 2132 5362 2144 5382
rect 2100 5320 2144 5362
rect 6658 5361 6702 5399
rect 6658 5341 6670 5361
rect 6690 5341 6702 5361
rect 6658 5299 6702 5341
rect 6752 5361 6794 5399
rect 6752 5341 6766 5361
rect 6786 5341 6794 5361
rect 6752 5299 6794 5341
rect 6871 5361 6915 5399
rect 6871 5341 6883 5361
rect 6903 5341 6915 5361
rect 6871 5299 6915 5341
rect 6965 5361 7007 5399
rect 6965 5341 6979 5361
rect 6999 5341 7007 5361
rect 6965 5299 7007 5341
rect 7079 5361 7123 5399
rect 7079 5341 7091 5361
rect 7111 5341 7123 5361
rect 7079 5299 7123 5341
rect 7173 5361 7215 5399
rect 7173 5341 7187 5361
rect 7207 5341 7215 5361
rect 7173 5299 7215 5341
rect 7289 5361 7331 5399
rect 7289 5341 7297 5361
rect 7317 5341 7331 5361
rect 7289 5299 7331 5341
rect 7381 5368 7426 5399
rect 7381 5361 7425 5368
rect 7381 5341 7393 5361
rect 7413 5341 7425 5361
rect 7381 5299 7425 5341
rect 12038 5390 12082 5428
rect 12038 5370 12050 5390
rect 12070 5370 12082 5390
rect 315 5143 359 5181
rect 315 5123 327 5143
rect 347 5123 359 5143
rect 315 5081 359 5123
rect 409 5143 451 5181
rect 409 5123 423 5143
rect 443 5123 451 5143
rect 409 5081 451 5123
rect 528 5143 572 5181
rect 528 5123 540 5143
rect 560 5123 572 5143
rect 528 5081 572 5123
rect 622 5143 664 5181
rect 622 5123 636 5143
rect 656 5123 664 5143
rect 622 5081 664 5123
rect 736 5143 780 5181
rect 736 5123 748 5143
rect 768 5123 780 5143
rect 736 5081 780 5123
rect 830 5143 872 5181
rect 830 5123 844 5143
rect 864 5123 872 5143
rect 830 5081 872 5123
rect 946 5143 988 5181
rect 946 5123 954 5143
rect 974 5123 988 5143
rect 946 5081 988 5123
rect 1038 5150 1083 5181
rect 4144 5177 4188 5219
rect 4144 5157 4156 5177
rect 4176 5157 4188 5177
rect 4144 5150 4188 5157
rect 1038 5143 1082 5150
rect 1038 5123 1050 5143
rect 1070 5123 1082 5143
rect 1038 5081 1082 5123
rect 4143 5119 4188 5150
rect 4238 5177 4280 5219
rect 4238 5157 4252 5177
rect 4272 5157 4280 5177
rect 4238 5119 4280 5157
rect 4354 5177 4396 5219
rect 4354 5157 4362 5177
rect 4382 5157 4396 5177
rect 4354 5119 4396 5157
rect 4446 5177 4490 5219
rect 4446 5157 4458 5177
rect 4478 5157 4490 5177
rect 4446 5119 4490 5157
rect 4562 5177 4604 5219
rect 4562 5157 4570 5177
rect 4590 5157 4604 5177
rect 4562 5119 4604 5157
rect 4654 5177 4698 5219
rect 4654 5157 4666 5177
rect 4686 5157 4698 5177
rect 4654 5119 4698 5157
rect 4775 5177 4817 5219
rect 4775 5157 4783 5177
rect 4803 5157 4817 5177
rect 4775 5119 4817 5157
rect 4867 5177 4911 5219
rect 12038 5328 12082 5370
rect 12132 5390 12174 5428
rect 12132 5370 12146 5390
rect 12166 5370 12174 5390
rect 12132 5328 12174 5370
rect 12251 5390 12295 5428
rect 12251 5370 12263 5390
rect 12283 5370 12295 5390
rect 12251 5328 12295 5370
rect 12345 5390 12387 5428
rect 12345 5370 12359 5390
rect 12379 5370 12387 5390
rect 12345 5328 12387 5370
rect 12459 5390 12503 5428
rect 12459 5370 12471 5390
rect 12491 5370 12503 5390
rect 12459 5328 12503 5370
rect 12553 5390 12595 5428
rect 12553 5370 12567 5390
rect 12587 5370 12595 5390
rect 12553 5328 12595 5370
rect 12669 5390 12711 5428
rect 12669 5370 12677 5390
rect 12697 5370 12711 5390
rect 12669 5328 12711 5370
rect 12761 5397 12806 5428
rect 12761 5390 12805 5397
rect 12761 5370 12773 5390
rect 12793 5370 12805 5390
rect 12761 5328 12805 5370
rect 17319 5369 17363 5407
rect 17319 5349 17331 5369
rect 17351 5349 17363 5369
rect 17319 5307 17363 5349
rect 17413 5369 17455 5407
rect 17413 5349 17427 5369
rect 17447 5349 17455 5369
rect 17413 5307 17455 5349
rect 17532 5369 17576 5407
rect 17532 5349 17544 5369
rect 17564 5349 17576 5369
rect 17532 5307 17576 5349
rect 17626 5369 17668 5407
rect 17626 5349 17640 5369
rect 17660 5349 17668 5369
rect 17626 5307 17668 5349
rect 17740 5369 17784 5407
rect 17740 5349 17752 5369
rect 17772 5349 17784 5369
rect 17740 5307 17784 5349
rect 17834 5369 17876 5407
rect 17834 5349 17848 5369
rect 17868 5349 17876 5369
rect 17834 5307 17876 5349
rect 17950 5369 17992 5407
rect 17950 5349 17958 5369
rect 17978 5349 17992 5369
rect 17950 5307 17992 5349
rect 18042 5376 18087 5407
rect 18042 5369 18086 5376
rect 18042 5349 18054 5369
rect 18074 5349 18086 5369
rect 18042 5307 18086 5349
rect 4867 5157 4879 5177
rect 4899 5157 4911 5177
rect 4867 5119 4911 5157
rect 5596 5122 5640 5160
rect 5596 5102 5608 5122
rect 5628 5102 5640 5122
rect 1327 4962 1371 5000
rect 1327 4942 1339 4962
rect 1359 4942 1371 4962
rect 1327 4900 1371 4942
rect 1421 4962 1463 5000
rect 1421 4942 1435 4962
rect 1455 4942 1463 4962
rect 1421 4900 1463 4942
rect 1540 4962 1584 5000
rect 1540 4942 1552 4962
rect 1572 4942 1584 4962
rect 1540 4900 1584 4942
rect 1634 4962 1676 5000
rect 1634 4942 1648 4962
rect 1668 4942 1676 4962
rect 1634 4900 1676 4942
rect 1748 4962 1792 5000
rect 1748 4942 1760 4962
rect 1780 4942 1792 4962
rect 1748 4900 1792 4942
rect 1842 4962 1884 5000
rect 1842 4942 1856 4962
rect 1876 4942 1884 4962
rect 1842 4900 1884 4942
rect 1958 4962 2000 5000
rect 1958 4942 1966 4962
rect 1986 4942 2000 4962
rect 1958 4900 2000 4942
rect 2050 4969 2095 5000
rect 5596 5060 5640 5102
rect 5690 5122 5732 5160
rect 5690 5102 5704 5122
rect 5724 5102 5732 5122
rect 5690 5060 5732 5102
rect 5809 5122 5853 5160
rect 5809 5102 5821 5122
rect 5841 5102 5853 5122
rect 5809 5060 5853 5102
rect 5903 5122 5945 5160
rect 5903 5102 5917 5122
rect 5937 5102 5945 5122
rect 5903 5060 5945 5102
rect 6017 5122 6061 5160
rect 6017 5102 6029 5122
rect 6049 5102 6061 5122
rect 6017 5060 6061 5102
rect 6111 5122 6153 5160
rect 6111 5102 6125 5122
rect 6145 5102 6153 5122
rect 6111 5060 6153 5102
rect 6227 5122 6269 5160
rect 6227 5102 6235 5122
rect 6255 5102 6269 5122
rect 6227 5060 6269 5102
rect 6319 5129 6364 5160
rect 9425 5156 9469 5198
rect 9425 5136 9437 5156
rect 9457 5136 9469 5156
rect 9425 5129 9469 5136
rect 6319 5122 6363 5129
rect 6319 5102 6331 5122
rect 6351 5102 6363 5122
rect 6319 5060 6363 5102
rect 9424 5098 9469 5129
rect 9519 5156 9561 5198
rect 9519 5136 9533 5156
rect 9553 5136 9561 5156
rect 9519 5098 9561 5136
rect 9635 5156 9677 5198
rect 9635 5136 9643 5156
rect 9663 5136 9677 5156
rect 9635 5098 9677 5136
rect 9727 5156 9771 5198
rect 9727 5136 9739 5156
rect 9759 5136 9771 5156
rect 9727 5098 9771 5136
rect 9843 5156 9885 5198
rect 9843 5136 9851 5156
rect 9871 5136 9885 5156
rect 9843 5098 9885 5136
rect 9935 5156 9979 5198
rect 9935 5136 9947 5156
rect 9967 5136 9979 5156
rect 9935 5098 9979 5136
rect 10056 5156 10098 5198
rect 10056 5136 10064 5156
rect 10084 5136 10098 5156
rect 10056 5098 10098 5136
rect 10148 5156 10192 5198
rect 10148 5136 10160 5156
rect 10180 5136 10192 5156
rect 10148 5098 10192 5136
rect 10976 5151 11020 5189
rect 10976 5131 10988 5151
rect 11008 5131 11020 5151
rect 2050 4962 2094 4969
rect 2050 4942 2062 4962
rect 2082 4942 2094 4962
rect 2050 4900 2094 4942
rect 3131 4943 3175 4985
rect 3131 4923 3143 4943
rect 3163 4923 3175 4943
rect 3131 4916 3175 4923
rect 3130 4885 3175 4916
rect 3225 4943 3267 4985
rect 3225 4923 3239 4943
rect 3259 4923 3267 4943
rect 3225 4885 3267 4923
rect 3341 4943 3383 4985
rect 3341 4923 3349 4943
rect 3369 4923 3383 4943
rect 3341 4885 3383 4923
rect 3433 4943 3477 4985
rect 3433 4923 3445 4943
rect 3465 4923 3477 4943
rect 3433 4885 3477 4923
rect 3549 4943 3591 4985
rect 3549 4923 3557 4943
rect 3577 4923 3591 4943
rect 3549 4885 3591 4923
rect 3641 4943 3685 4985
rect 3641 4923 3653 4943
rect 3673 4923 3685 4943
rect 3641 4885 3685 4923
rect 3762 4943 3804 4985
rect 3762 4923 3770 4943
rect 3790 4923 3804 4943
rect 3762 4885 3804 4923
rect 3854 4943 3898 4985
rect 10976 5089 11020 5131
rect 11070 5151 11112 5189
rect 11070 5131 11084 5151
rect 11104 5131 11112 5151
rect 11070 5089 11112 5131
rect 11189 5151 11233 5189
rect 11189 5131 11201 5151
rect 11221 5131 11233 5151
rect 11189 5089 11233 5131
rect 11283 5151 11325 5189
rect 11283 5131 11297 5151
rect 11317 5131 11325 5151
rect 11283 5089 11325 5131
rect 11397 5151 11441 5189
rect 11397 5131 11409 5151
rect 11429 5131 11441 5151
rect 11397 5089 11441 5131
rect 11491 5151 11533 5189
rect 11491 5131 11505 5151
rect 11525 5131 11533 5151
rect 11491 5089 11533 5131
rect 11607 5151 11649 5189
rect 11607 5131 11615 5151
rect 11635 5131 11649 5151
rect 11607 5089 11649 5131
rect 11699 5158 11744 5189
rect 14805 5185 14849 5227
rect 14805 5165 14817 5185
rect 14837 5165 14849 5185
rect 14805 5158 14849 5165
rect 11699 5151 11743 5158
rect 11699 5131 11711 5151
rect 11731 5131 11743 5151
rect 11699 5089 11743 5131
rect 14804 5127 14849 5158
rect 14899 5185 14941 5227
rect 14899 5165 14913 5185
rect 14933 5165 14941 5185
rect 14899 5127 14941 5165
rect 15015 5185 15057 5227
rect 15015 5165 15023 5185
rect 15043 5165 15057 5185
rect 15015 5127 15057 5165
rect 15107 5185 15151 5227
rect 15107 5165 15119 5185
rect 15139 5165 15151 5185
rect 15107 5127 15151 5165
rect 15223 5185 15265 5227
rect 15223 5165 15231 5185
rect 15251 5165 15265 5185
rect 15223 5127 15265 5165
rect 15315 5185 15359 5227
rect 15315 5165 15327 5185
rect 15347 5165 15359 5185
rect 15315 5127 15359 5165
rect 15436 5185 15478 5227
rect 15436 5165 15444 5185
rect 15464 5165 15478 5185
rect 15436 5127 15478 5165
rect 15528 5185 15572 5227
rect 15528 5165 15540 5185
rect 15560 5165 15572 5185
rect 15528 5127 15572 5165
rect 3854 4923 3866 4943
rect 3886 4923 3898 4943
rect 6608 4941 6652 4979
rect 3854 4885 3898 4923
rect 6608 4921 6620 4941
rect 6640 4921 6652 4941
rect 6608 4879 6652 4921
rect 6702 4941 6744 4979
rect 6702 4921 6716 4941
rect 6736 4921 6744 4941
rect 6702 4879 6744 4921
rect 6821 4941 6865 4979
rect 6821 4921 6833 4941
rect 6853 4921 6865 4941
rect 6821 4879 6865 4921
rect 6915 4941 6957 4979
rect 6915 4921 6929 4941
rect 6949 4921 6957 4941
rect 6915 4879 6957 4921
rect 7029 4941 7073 4979
rect 7029 4921 7041 4941
rect 7061 4921 7073 4941
rect 7029 4879 7073 4921
rect 7123 4941 7165 4979
rect 7123 4921 7137 4941
rect 7157 4921 7165 4941
rect 7123 4879 7165 4921
rect 7239 4941 7281 4979
rect 7239 4921 7247 4941
rect 7267 4921 7281 4941
rect 7239 4879 7281 4921
rect 7331 4948 7376 4979
rect 16257 5130 16301 5168
rect 16257 5110 16269 5130
rect 16289 5110 16301 5130
rect 11988 4970 12032 5008
rect 7331 4941 7375 4948
rect 7331 4921 7343 4941
rect 7363 4921 7375 4941
rect 7331 4879 7375 4921
rect 8412 4922 8456 4964
rect 8412 4902 8424 4922
rect 8444 4902 8456 4922
rect 8412 4895 8456 4902
rect 314 4728 358 4766
rect 314 4708 326 4728
rect 346 4708 358 4728
rect 314 4666 358 4708
rect 408 4728 450 4766
rect 408 4708 422 4728
rect 442 4708 450 4728
rect 408 4666 450 4708
rect 527 4728 571 4766
rect 527 4708 539 4728
rect 559 4708 571 4728
rect 527 4666 571 4708
rect 621 4728 663 4766
rect 621 4708 635 4728
rect 655 4708 663 4728
rect 621 4666 663 4708
rect 735 4728 779 4766
rect 735 4708 747 4728
rect 767 4708 779 4728
rect 735 4666 779 4708
rect 829 4728 871 4766
rect 829 4708 843 4728
rect 863 4708 871 4728
rect 829 4666 871 4708
rect 945 4728 987 4766
rect 945 4708 953 4728
rect 973 4708 987 4728
rect 945 4666 987 4708
rect 1037 4735 1082 4766
rect 4143 4762 4187 4804
rect 4143 4742 4155 4762
rect 4175 4742 4187 4762
rect 4143 4735 4187 4742
rect 1037 4728 1081 4735
rect 1037 4708 1049 4728
rect 1069 4708 1081 4728
rect 1037 4666 1081 4708
rect 4142 4704 4187 4735
rect 4237 4762 4279 4804
rect 4237 4742 4251 4762
rect 4271 4742 4279 4762
rect 4237 4704 4279 4742
rect 4353 4762 4395 4804
rect 4353 4742 4361 4762
rect 4381 4742 4395 4762
rect 4353 4704 4395 4742
rect 4445 4762 4489 4804
rect 4445 4742 4457 4762
rect 4477 4742 4489 4762
rect 4445 4704 4489 4742
rect 4561 4762 4603 4804
rect 4561 4742 4569 4762
rect 4589 4742 4603 4762
rect 4561 4704 4603 4742
rect 4653 4762 4697 4804
rect 4653 4742 4665 4762
rect 4685 4742 4697 4762
rect 4653 4704 4697 4742
rect 4774 4762 4816 4804
rect 4774 4742 4782 4762
rect 4802 4742 4816 4762
rect 4774 4704 4816 4742
rect 4866 4762 4910 4804
rect 8411 4864 8456 4895
rect 8506 4922 8548 4964
rect 8506 4902 8520 4922
rect 8540 4902 8548 4922
rect 8506 4864 8548 4902
rect 8622 4922 8664 4964
rect 8622 4902 8630 4922
rect 8650 4902 8664 4922
rect 8622 4864 8664 4902
rect 8714 4922 8758 4964
rect 8714 4902 8726 4922
rect 8746 4902 8758 4922
rect 8714 4864 8758 4902
rect 8830 4922 8872 4964
rect 8830 4902 8838 4922
rect 8858 4902 8872 4922
rect 8830 4864 8872 4902
rect 8922 4922 8966 4964
rect 8922 4902 8934 4922
rect 8954 4902 8966 4922
rect 8922 4864 8966 4902
rect 9043 4922 9085 4964
rect 9043 4902 9051 4922
rect 9071 4902 9085 4922
rect 9043 4864 9085 4902
rect 9135 4922 9179 4964
rect 9135 4902 9147 4922
rect 9167 4902 9179 4922
rect 11988 4950 12000 4970
rect 12020 4950 12032 4970
rect 11988 4908 12032 4950
rect 12082 4970 12124 5008
rect 12082 4950 12096 4970
rect 12116 4950 12124 4970
rect 12082 4908 12124 4950
rect 12201 4970 12245 5008
rect 12201 4950 12213 4970
rect 12233 4950 12245 4970
rect 12201 4908 12245 4950
rect 12295 4970 12337 5008
rect 12295 4950 12309 4970
rect 12329 4950 12337 4970
rect 12295 4908 12337 4950
rect 12409 4970 12453 5008
rect 12409 4950 12421 4970
rect 12441 4950 12453 4970
rect 12409 4908 12453 4950
rect 12503 4970 12545 5008
rect 12503 4950 12517 4970
rect 12537 4950 12545 4970
rect 12503 4908 12545 4950
rect 12619 4970 12661 5008
rect 12619 4950 12627 4970
rect 12647 4950 12661 4970
rect 12619 4908 12661 4950
rect 12711 4977 12756 5008
rect 16257 5068 16301 5110
rect 16351 5130 16393 5168
rect 16351 5110 16365 5130
rect 16385 5110 16393 5130
rect 16351 5068 16393 5110
rect 16470 5130 16514 5168
rect 16470 5110 16482 5130
rect 16502 5110 16514 5130
rect 16470 5068 16514 5110
rect 16564 5130 16606 5168
rect 16564 5110 16578 5130
rect 16598 5110 16606 5130
rect 16564 5068 16606 5110
rect 16678 5130 16722 5168
rect 16678 5110 16690 5130
rect 16710 5110 16722 5130
rect 16678 5068 16722 5110
rect 16772 5130 16814 5168
rect 16772 5110 16786 5130
rect 16806 5110 16814 5130
rect 16772 5068 16814 5110
rect 16888 5130 16930 5168
rect 16888 5110 16896 5130
rect 16916 5110 16930 5130
rect 16888 5068 16930 5110
rect 16980 5137 17025 5168
rect 20086 5164 20130 5206
rect 20086 5144 20098 5164
rect 20118 5144 20130 5164
rect 20086 5137 20130 5144
rect 16980 5130 17024 5137
rect 16980 5110 16992 5130
rect 17012 5110 17024 5130
rect 16980 5068 17024 5110
rect 20085 5106 20130 5137
rect 20180 5164 20222 5206
rect 20180 5144 20194 5164
rect 20214 5144 20222 5164
rect 20180 5106 20222 5144
rect 20296 5164 20338 5206
rect 20296 5144 20304 5164
rect 20324 5144 20338 5164
rect 20296 5106 20338 5144
rect 20388 5164 20432 5206
rect 20388 5144 20400 5164
rect 20420 5144 20432 5164
rect 20388 5106 20432 5144
rect 20504 5164 20546 5206
rect 20504 5144 20512 5164
rect 20532 5144 20546 5164
rect 20504 5106 20546 5144
rect 20596 5164 20640 5206
rect 20596 5144 20608 5164
rect 20628 5144 20640 5164
rect 20596 5106 20640 5144
rect 20717 5164 20759 5206
rect 20717 5144 20725 5164
rect 20745 5144 20759 5164
rect 20717 5106 20759 5144
rect 20809 5164 20853 5206
rect 20809 5144 20821 5164
rect 20841 5144 20853 5164
rect 20809 5106 20853 5144
rect 12711 4970 12755 4977
rect 12711 4950 12723 4970
rect 12743 4950 12755 4970
rect 12711 4908 12755 4950
rect 13792 4951 13836 4993
rect 13792 4931 13804 4951
rect 13824 4931 13836 4951
rect 13792 4924 13836 4931
rect 9135 4864 9179 4902
rect 4866 4742 4878 4762
rect 4898 4742 4910 4762
rect 4866 4704 4910 4742
rect 13791 4893 13836 4924
rect 13886 4951 13928 4993
rect 13886 4931 13900 4951
rect 13920 4931 13928 4951
rect 13886 4893 13928 4931
rect 14002 4951 14044 4993
rect 14002 4931 14010 4951
rect 14030 4931 14044 4951
rect 14002 4893 14044 4931
rect 14094 4951 14138 4993
rect 14094 4931 14106 4951
rect 14126 4931 14138 4951
rect 14094 4893 14138 4931
rect 14210 4951 14252 4993
rect 14210 4931 14218 4951
rect 14238 4931 14252 4951
rect 14210 4893 14252 4931
rect 14302 4951 14346 4993
rect 14302 4931 14314 4951
rect 14334 4931 14346 4951
rect 14302 4893 14346 4931
rect 14423 4951 14465 4993
rect 14423 4931 14431 4951
rect 14451 4931 14465 4951
rect 14423 4893 14465 4931
rect 14515 4951 14559 4993
rect 14515 4931 14527 4951
rect 14547 4931 14559 4951
rect 17269 4949 17313 4987
rect 14515 4893 14559 4931
rect 17269 4929 17281 4949
rect 17301 4929 17313 4949
rect 5595 4707 5639 4745
rect 5595 4687 5607 4707
rect 5627 4687 5639 4707
rect 5595 4645 5639 4687
rect 5689 4707 5731 4745
rect 5689 4687 5703 4707
rect 5723 4687 5731 4707
rect 5689 4645 5731 4687
rect 5808 4707 5852 4745
rect 5808 4687 5820 4707
rect 5840 4687 5852 4707
rect 5808 4645 5852 4687
rect 5902 4707 5944 4745
rect 5902 4687 5916 4707
rect 5936 4687 5944 4707
rect 5902 4645 5944 4687
rect 6016 4707 6060 4745
rect 6016 4687 6028 4707
rect 6048 4687 6060 4707
rect 6016 4645 6060 4687
rect 6110 4707 6152 4745
rect 6110 4687 6124 4707
rect 6144 4687 6152 4707
rect 6110 4645 6152 4687
rect 6226 4707 6268 4745
rect 6226 4687 6234 4707
rect 6254 4687 6268 4707
rect 6226 4645 6268 4687
rect 6318 4714 6363 4745
rect 9424 4741 9468 4783
rect 9424 4721 9436 4741
rect 9456 4721 9468 4741
rect 9424 4714 9468 4721
rect 6318 4707 6362 4714
rect 6318 4687 6330 4707
rect 6350 4687 6362 4707
rect 6318 4645 6362 4687
rect 9423 4683 9468 4714
rect 9518 4741 9560 4783
rect 9518 4721 9532 4741
rect 9552 4721 9560 4741
rect 9518 4683 9560 4721
rect 9634 4741 9676 4783
rect 9634 4721 9642 4741
rect 9662 4721 9676 4741
rect 9634 4683 9676 4721
rect 9726 4741 9770 4783
rect 9726 4721 9738 4741
rect 9758 4721 9770 4741
rect 9726 4683 9770 4721
rect 9842 4741 9884 4783
rect 9842 4721 9850 4741
rect 9870 4721 9884 4741
rect 9842 4683 9884 4721
rect 9934 4741 9978 4783
rect 9934 4721 9946 4741
rect 9966 4721 9978 4741
rect 9934 4683 9978 4721
rect 10055 4741 10097 4783
rect 10055 4721 10063 4741
rect 10083 4721 10097 4741
rect 10055 4683 10097 4721
rect 10147 4741 10191 4783
rect 17269 4887 17313 4929
rect 17363 4949 17405 4987
rect 17363 4929 17377 4949
rect 17397 4929 17405 4949
rect 17363 4887 17405 4929
rect 17482 4949 17526 4987
rect 17482 4929 17494 4949
rect 17514 4929 17526 4949
rect 17482 4887 17526 4929
rect 17576 4949 17618 4987
rect 17576 4929 17590 4949
rect 17610 4929 17618 4949
rect 17576 4887 17618 4929
rect 17690 4949 17734 4987
rect 17690 4929 17702 4949
rect 17722 4929 17734 4949
rect 17690 4887 17734 4929
rect 17784 4949 17826 4987
rect 17784 4929 17798 4949
rect 17818 4929 17826 4949
rect 17784 4887 17826 4929
rect 17900 4949 17942 4987
rect 17900 4929 17908 4949
rect 17928 4929 17942 4949
rect 17900 4887 17942 4929
rect 17992 4956 18037 4987
rect 17992 4949 18036 4956
rect 17992 4929 18004 4949
rect 18024 4929 18036 4949
rect 17992 4887 18036 4929
rect 19073 4930 19117 4972
rect 19073 4910 19085 4930
rect 19105 4910 19117 4930
rect 19073 4903 19117 4910
rect 10147 4721 10159 4741
rect 10179 4721 10191 4741
rect 10147 4683 10191 4721
rect 10975 4736 11019 4774
rect 10975 4716 10987 4736
rect 11007 4716 11019 4736
rect 10975 4674 11019 4716
rect 11069 4736 11111 4774
rect 11069 4716 11083 4736
rect 11103 4716 11111 4736
rect 11069 4674 11111 4716
rect 11188 4736 11232 4774
rect 11188 4716 11200 4736
rect 11220 4716 11232 4736
rect 11188 4674 11232 4716
rect 11282 4736 11324 4774
rect 11282 4716 11296 4736
rect 11316 4716 11324 4736
rect 11282 4674 11324 4716
rect 11396 4736 11440 4774
rect 11396 4716 11408 4736
rect 11428 4716 11440 4736
rect 11396 4674 11440 4716
rect 11490 4736 11532 4774
rect 11490 4716 11504 4736
rect 11524 4716 11532 4736
rect 11490 4674 11532 4716
rect 11606 4736 11648 4774
rect 11606 4716 11614 4736
rect 11634 4716 11648 4736
rect 11606 4674 11648 4716
rect 11698 4743 11743 4774
rect 14804 4770 14848 4812
rect 14804 4750 14816 4770
rect 14836 4750 14848 4770
rect 14804 4743 14848 4750
rect 11698 4736 11742 4743
rect 11698 4716 11710 4736
rect 11730 4716 11742 4736
rect 11698 4674 11742 4716
rect 14803 4712 14848 4743
rect 14898 4770 14940 4812
rect 14898 4750 14912 4770
rect 14932 4750 14940 4770
rect 14898 4712 14940 4750
rect 15014 4770 15056 4812
rect 15014 4750 15022 4770
rect 15042 4750 15056 4770
rect 15014 4712 15056 4750
rect 15106 4770 15150 4812
rect 15106 4750 15118 4770
rect 15138 4750 15150 4770
rect 15106 4712 15150 4750
rect 15222 4770 15264 4812
rect 15222 4750 15230 4770
rect 15250 4750 15264 4770
rect 15222 4712 15264 4750
rect 15314 4770 15358 4812
rect 15314 4750 15326 4770
rect 15346 4750 15358 4770
rect 15314 4712 15358 4750
rect 15435 4770 15477 4812
rect 15435 4750 15443 4770
rect 15463 4750 15477 4770
rect 15435 4712 15477 4750
rect 15527 4770 15571 4812
rect 19072 4872 19117 4903
rect 19167 4930 19209 4972
rect 19167 4910 19181 4930
rect 19201 4910 19209 4930
rect 19167 4872 19209 4910
rect 19283 4930 19325 4972
rect 19283 4910 19291 4930
rect 19311 4910 19325 4930
rect 19283 4872 19325 4910
rect 19375 4930 19419 4972
rect 19375 4910 19387 4930
rect 19407 4910 19419 4930
rect 19375 4872 19419 4910
rect 19491 4930 19533 4972
rect 19491 4910 19499 4930
rect 19519 4910 19533 4930
rect 19491 4872 19533 4910
rect 19583 4930 19627 4972
rect 19583 4910 19595 4930
rect 19615 4910 19627 4930
rect 19583 4872 19627 4910
rect 19704 4930 19746 4972
rect 19704 4910 19712 4930
rect 19732 4910 19746 4930
rect 19704 4872 19746 4910
rect 19796 4930 19840 4972
rect 19796 4910 19808 4930
rect 19828 4910 19840 4930
rect 19796 4872 19840 4910
rect 15527 4750 15539 4770
rect 15559 4750 15571 4770
rect 15527 4712 15571 4750
rect 16256 4715 16300 4753
rect 16256 4695 16268 4715
rect 16288 4695 16300 4715
rect 2836 4511 2880 4553
rect 2836 4491 2848 4511
rect 2868 4491 2880 4511
rect 2836 4484 2880 4491
rect 1625 4418 1669 4456
rect 1625 4398 1637 4418
rect 1657 4398 1669 4418
rect 1625 4356 1669 4398
rect 1719 4418 1761 4456
rect 1719 4398 1733 4418
rect 1753 4398 1761 4418
rect 1719 4356 1761 4398
rect 1838 4418 1882 4456
rect 1838 4398 1850 4418
rect 1870 4398 1882 4418
rect 1838 4356 1882 4398
rect 1932 4418 1974 4456
rect 1932 4398 1946 4418
rect 1966 4398 1974 4418
rect 1932 4356 1974 4398
rect 2046 4418 2090 4456
rect 2046 4398 2058 4418
rect 2078 4398 2090 4418
rect 2046 4356 2090 4398
rect 2140 4418 2182 4456
rect 2140 4398 2154 4418
rect 2174 4398 2182 4418
rect 2140 4356 2182 4398
rect 2256 4418 2298 4456
rect 2256 4398 2264 4418
rect 2284 4398 2298 4418
rect 2256 4356 2298 4398
rect 2348 4425 2393 4456
rect 2835 4453 2880 4484
rect 2930 4511 2972 4553
rect 2930 4491 2944 4511
rect 2964 4491 2972 4511
rect 2930 4453 2972 4491
rect 3046 4511 3088 4553
rect 3046 4491 3054 4511
rect 3074 4491 3088 4511
rect 3046 4453 3088 4491
rect 3138 4511 3182 4553
rect 3138 4491 3150 4511
rect 3170 4491 3182 4511
rect 3138 4453 3182 4491
rect 3254 4511 3296 4553
rect 3254 4491 3262 4511
rect 3282 4491 3296 4511
rect 3254 4453 3296 4491
rect 3346 4511 3390 4553
rect 3346 4491 3358 4511
rect 3378 4491 3390 4511
rect 3346 4453 3390 4491
rect 3467 4511 3509 4553
rect 3467 4491 3475 4511
rect 3495 4491 3509 4511
rect 3467 4453 3509 4491
rect 3559 4511 3603 4553
rect 3559 4491 3571 4511
rect 3591 4491 3603 4511
rect 3559 4453 3603 4491
rect 16256 4653 16300 4695
rect 16350 4715 16392 4753
rect 16350 4695 16364 4715
rect 16384 4695 16392 4715
rect 16350 4653 16392 4695
rect 16469 4715 16513 4753
rect 16469 4695 16481 4715
rect 16501 4695 16513 4715
rect 16469 4653 16513 4695
rect 16563 4715 16605 4753
rect 16563 4695 16577 4715
rect 16597 4695 16605 4715
rect 16563 4653 16605 4695
rect 16677 4715 16721 4753
rect 16677 4695 16689 4715
rect 16709 4695 16721 4715
rect 16677 4653 16721 4695
rect 16771 4715 16813 4753
rect 16771 4695 16785 4715
rect 16805 4695 16813 4715
rect 16771 4653 16813 4695
rect 16887 4715 16929 4753
rect 16887 4695 16895 4715
rect 16915 4695 16929 4715
rect 16887 4653 16929 4695
rect 16979 4722 17024 4753
rect 20085 4749 20129 4791
rect 20085 4729 20097 4749
rect 20117 4729 20129 4749
rect 20085 4722 20129 4729
rect 16979 4715 17023 4722
rect 16979 4695 16991 4715
rect 17011 4695 17023 4715
rect 16979 4653 17023 4695
rect 20084 4691 20129 4722
rect 20179 4749 20221 4791
rect 20179 4729 20193 4749
rect 20213 4729 20221 4749
rect 20179 4691 20221 4729
rect 20295 4749 20337 4791
rect 20295 4729 20303 4749
rect 20323 4729 20337 4749
rect 20295 4691 20337 4729
rect 20387 4749 20431 4791
rect 20387 4729 20399 4749
rect 20419 4729 20431 4749
rect 20387 4691 20431 4729
rect 20503 4749 20545 4791
rect 20503 4729 20511 4749
rect 20531 4729 20545 4749
rect 20503 4691 20545 4729
rect 20595 4749 20639 4791
rect 20595 4729 20607 4749
rect 20627 4729 20639 4749
rect 20595 4691 20639 4729
rect 20716 4749 20758 4791
rect 20716 4729 20724 4749
rect 20744 4729 20758 4749
rect 20716 4691 20758 4729
rect 20808 4749 20852 4791
rect 20808 4729 20820 4749
rect 20840 4729 20852 4749
rect 20808 4691 20852 4729
rect 8117 4490 8161 4532
rect 8117 4470 8129 4490
rect 8149 4470 8161 4490
rect 8117 4463 8161 4470
rect 2348 4418 2392 4425
rect 2348 4398 2360 4418
rect 2380 4398 2392 4418
rect 2348 4356 2392 4398
rect 6906 4397 6950 4435
rect 6906 4377 6918 4397
rect 6938 4377 6950 4397
rect 6906 4335 6950 4377
rect 7000 4397 7042 4435
rect 7000 4377 7014 4397
rect 7034 4377 7042 4397
rect 7000 4335 7042 4377
rect 7119 4397 7163 4435
rect 7119 4377 7131 4397
rect 7151 4377 7163 4397
rect 7119 4335 7163 4377
rect 7213 4397 7255 4435
rect 7213 4377 7227 4397
rect 7247 4377 7255 4397
rect 7213 4335 7255 4377
rect 7327 4397 7371 4435
rect 7327 4377 7339 4397
rect 7359 4377 7371 4397
rect 7327 4335 7371 4377
rect 7421 4397 7463 4435
rect 7421 4377 7435 4397
rect 7455 4377 7463 4397
rect 7421 4335 7463 4377
rect 7537 4397 7579 4435
rect 7537 4377 7545 4397
rect 7565 4377 7579 4397
rect 7537 4335 7579 4377
rect 7629 4404 7674 4435
rect 8116 4432 8161 4463
rect 8211 4490 8253 4532
rect 8211 4470 8225 4490
rect 8245 4470 8253 4490
rect 8211 4432 8253 4470
rect 8327 4490 8369 4532
rect 8327 4470 8335 4490
rect 8355 4470 8369 4490
rect 8327 4432 8369 4470
rect 8419 4490 8463 4532
rect 8419 4470 8431 4490
rect 8451 4470 8463 4490
rect 8419 4432 8463 4470
rect 8535 4490 8577 4532
rect 8535 4470 8543 4490
rect 8563 4470 8577 4490
rect 8535 4432 8577 4470
rect 8627 4490 8671 4532
rect 8627 4470 8639 4490
rect 8659 4470 8671 4490
rect 8627 4432 8671 4470
rect 8748 4490 8790 4532
rect 8748 4470 8756 4490
rect 8776 4470 8790 4490
rect 8748 4432 8790 4470
rect 8840 4490 8884 4532
rect 8840 4470 8852 4490
rect 8872 4470 8884 4490
rect 8840 4432 8884 4470
rect 13497 4519 13541 4561
rect 13497 4499 13509 4519
rect 13529 4499 13541 4519
rect 13497 4492 13541 4499
rect 7629 4397 7673 4404
rect 7629 4377 7641 4397
rect 7661 4377 7673 4397
rect 7629 4335 7673 4377
rect 12286 4426 12330 4464
rect 12286 4406 12298 4426
rect 12318 4406 12330 4426
rect 12286 4364 12330 4406
rect 12380 4426 12422 4464
rect 12380 4406 12394 4426
rect 12414 4406 12422 4426
rect 12380 4364 12422 4406
rect 12499 4426 12543 4464
rect 12499 4406 12511 4426
rect 12531 4406 12543 4426
rect 12499 4364 12543 4406
rect 12593 4426 12635 4464
rect 12593 4406 12607 4426
rect 12627 4406 12635 4426
rect 12593 4364 12635 4406
rect 12707 4426 12751 4464
rect 12707 4406 12719 4426
rect 12739 4406 12751 4426
rect 12707 4364 12751 4406
rect 12801 4426 12843 4464
rect 12801 4406 12815 4426
rect 12835 4406 12843 4426
rect 12801 4364 12843 4406
rect 12917 4426 12959 4464
rect 12917 4406 12925 4426
rect 12945 4406 12959 4426
rect 12917 4364 12959 4406
rect 13009 4433 13054 4464
rect 13496 4461 13541 4492
rect 13591 4519 13633 4561
rect 13591 4499 13605 4519
rect 13625 4499 13633 4519
rect 13591 4461 13633 4499
rect 13707 4519 13749 4561
rect 13707 4499 13715 4519
rect 13735 4499 13749 4519
rect 13707 4461 13749 4499
rect 13799 4519 13843 4561
rect 13799 4499 13811 4519
rect 13831 4499 13843 4519
rect 13799 4461 13843 4499
rect 13915 4519 13957 4561
rect 13915 4499 13923 4519
rect 13943 4499 13957 4519
rect 13915 4461 13957 4499
rect 14007 4519 14051 4561
rect 14007 4499 14019 4519
rect 14039 4499 14051 4519
rect 14007 4461 14051 4499
rect 14128 4519 14170 4561
rect 14128 4499 14136 4519
rect 14156 4499 14170 4519
rect 14128 4461 14170 4499
rect 14220 4519 14264 4561
rect 14220 4499 14232 4519
rect 14252 4499 14264 4519
rect 14220 4461 14264 4499
rect 18778 4498 18822 4540
rect 18778 4478 18790 4498
rect 18810 4478 18822 4498
rect 18778 4471 18822 4478
rect 13009 4426 13053 4433
rect 13009 4406 13021 4426
rect 13041 4406 13053 4426
rect 13009 4364 13053 4406
rect 318 4167 362 4205
rect 318 4147 330 4167
rect 350 4147 362 4167
rect 318 4105 362 4147
rect 412 4167 454 4205
rect 412 4147 426 4167
rect 446 4147 454 4167
rect 412 4105 454 4147
rect 531 4167 575 4205
rect 531 4147 543 4167
rect 563 4147 575 4167
rect 531 4105 575 4147
rect 625 4167 667 4205
rect 625 4147 639 4167
rect 659 4147 667 4167
rect 625 4105 667 4147
rect 739 4167 783 4205
rect 739 4147 751 4167
rect 771 4147 783 4167
rect 739 4105 783 4147
rect 833 4167 875 4205
rect 833 4147 847 4167
rect 867 4147 875 4167
rect 833 4105 875 4147
rect 949 4167 991 4205
rect 949 4147 957 4167
rect 977 4147 991 4167
rect 949 4105 991 4147
rect 1041 4174 1086 4205
rect 4147 4201 4191 4243
rect 4147 4181 4159 4201
rect 4179 4181 4191 4201
rect 4147 4174 4191 4181
rect 1041 4167 1085 4174
rect 1041 4147 1053 4167
rect 1073 4147 1085 4167
rect 1041 4105 1085 4147
rect 4146 4143 4191 4174
rect 4241 4201 4283 4243
rect 4241 4181 4255 4201
rect 4275 4181 4283 4201
rect 4241 4143 4283 4181
rect 4357 4201 4399 4243
rect 4357 4181 4365 4201
rect 4385 4181 4399 4201
rect 4357 4143 4399 4181
rect 4449 4201 4493 4243
rect 4449 4181 4461 4201
rect 4481 4181 4493 4201
rect 4449 4143 4493 4181
rect 4565 4201 4607 4243
rect 4565 4181 4573 4201
rect 4593 4181 4607 4201
rect 4565 4143 4607 4181
rect 4657 4201 4701 4243
rect 4657 4181 4669 4201
rect 4689 4181 4701 4201
rect 4657 4143 4701 4181
rect 4778 4201 4820 4243
rect 4778 4181 4786 4201
rect 4806 4181 4820 4201
rect 4778 4143 4820 4181
rect 4870 4201 4914 4243
rect 17567 4405 17611 4443
rect 17567 4385 17579 4405
rect 17599 4385 17611 4405
rect 17567 4343 17611 4385
rect 17661 4405 17703 4443
rect 17661 4385 17675 4405
rect 17695 4385 17703 4405
rect 17661 4343 17703 4385
rect 17780 4405 17824 4443
rect 17780 4385 17792 4405
rect 17812 4385 17824 4405
rect 17780 4343 17824 4385
rect 17874 4405 17916 4443
rect 17874 4385 17888 4405
rect 17908 4385 17916 4405
rect 17874 4343 17916 4385
rect 17988 4405 18032 4443
rect 17988 4385 18000 4405
rect 18020 4385 18032 4405
rect 17988 4343 18032 4385
rect 18082 4405 18124 4443
rect 18082 4385 18096 4405
rect 18116 4385 18124 4405
rect 18082 4343 18124 4385
rect 18198 4405 18240 4443
rect 18198 4385 18206 4405
rect 18226 4385 18240 4405
rect 18198 4343 18240 4385
rect 18290 4412 18335 4443
rect 18777 4440 18822 4471
rect 18872 4498 18914 4540
rect 18872 4478 18886 4498
rect 18906 4478 18914 4498
rect 18872 4440 18914 4478
rect 18988 4498 19030 4540
rect 18988 4478 18996 4498
rect 19016 4478 19030 4498
rect 18988 4440 19030 4478
rect 19080 4498 19124 4540
rect 19080 4478 19092 4498
rect 19112 4478 19124 4498
rect 19080 4440 19124 4478
rect 19196 4498 19238 4540
rect 19196 4478 19204 4498
rect 19224 4478 19238 4498
rect 19196 4440 19238 4478
rect 19288 4498 19332 4540
rect 19288 4478 19300 4498
rect 19320 4478 19332 4498
rect 19288 4440 19332 4478
rect 19409 4498 19451 4540
rect 19409 4478 19417 4498
rect 19437 4478 19451 4498
rect 19409 4440 19451 4478
rect 19501 4498 19545 4540
rect 19501 4478 19513 4498
rect 19533 4478 19545 4498
rect 19501 4440 19545 4478
rect 18290 4405 18334 4412
rect 18290 4385 18302 4405
rect 18322 4385 18334 4405
rect 18290 4343 18334 4385
rect 4870 4181 4882 4201
rect 4902 4181 4914 4201
rect 4870 4143 4914 4181
rect 5599 4146 5643 4184
rect 5599 4126 5611 4146
rect 5631 4126 5643 4146
rect 1330 3986 1374 4024
rect 1330 3966 1342 3986
rect 1362 3966 1374 3986
rect 1330 3924 1374 3966
rect 1424 3986 1466 4024
rect 1424 3966 1438 3986
rect 1458 3966 1466 3986
rect 1424 3924 1466 3966
rect 1543 3986 1587 4024
rect 1543 3966 1555 3986
rect 1575 3966 1587 3986
rect 1543 3924 1587 3966
rect 1637 3986 1679 4024
rect 1637 3966 1651 3986
rect 1671 3966 1679 3986
rect 1637 3924 1679 3966
rect 1751 3986 1795 4024
rect 1751 3966 1763 3986
rect 1783 3966 1795 3986
rect 1751 3924 1795 3966
rect 1845 3986 1887 4024
rect 1845 3966 1859 3986
rect 1879 3966 1887 3986
rect 1845 3924 1887 3966
rect 1961 3986 2003 4024
rect 1961 3966 1969 3986
rect 1989 3966 2003 3986
rect 1961 3924 2003 3966
rect 2053 3993 2098 4024
rect 5599 4084 5643 4126
rect 5693 4146 5735 4184
rect 5693 4126 5707 4146
rect 5727 4126 5735 4146
rect 5693 4084 5735 4126
rect 5812 4146 5856 4184
rect 5812 4126 5824 4146
rect 5844 4126 5856 4146
rect 5812 4084 5856 4126
rect 5906 4146 5948 4184
rect 5906 4126 5920 4146
rect 5940 4126 5948 4146
rect 5906 4084 5948 4126
rect 6020 4146 6064 4184
rect 6020 4126 6032 4146
rect 6052 4126 6064 4146
rect 6020 4084 6064 4126
rect 6114 4146 6156 4184
rect 6114 4126 6128 4146
rect 6148 4126 6156 4146
rect 6114 4084 6156 4126
rect 6230 4146 6272 4184
rect 6230 4126 6238 4146
rect 6258 4126 6272 4146
rect 6230 4084 6272 4126
rect 6322 4153 6367 4184
rect 9428 4180 9472 4222
rect 9428 4160 9440 4180
rect 9460 4160 9472 4180
rect 9428 4153 9472 4160
rect 6322 4146 6366 4153
rect 6322 4126 6334 4146
rect 6354 4126 6366 4146
rect 6322 4084 6366 4126
rect 9427 4122 9472 4153
rect 9522 4180 9564 4222
rect 9522 4160 9536 4180
rect 9556 4160 9564 4180
rect 9522 4122 9564 4160
rect 9638 4180 9680 4222
rect 9638 4160 9646 4180
rect 9666 4160 9680 4180
rect 9638 4122 9680 4160
rect 9730 4180 9774 4222
rect 9730 4160 9742 4180
rect 9762 4160 9774 4180
rect 9730 4122 9774 4160
rect 9846 4180 9888 4222
rect 9846 4160 9854 4180
rect 9874 4160 9888 4180
rect 9846 4122 9888 4160
rect 9938 4180 9982 4222
rect 9938 4160 9950 4180
rect 9970 4160 9982 4180
rect 9938 4122 9982 4160
rect 10059 4180 10101 4222
rect 10059 4160 10067 4180
rect 10087 4160 10101 4180
rect 10059 4122 10101 4160
rect 10151 4180 10195 4222
rect 10151 4160 10163 4180
rect 10183 4160 10195 4180
rect 10151 4122 10195 4160
rect 10979 4175 11023 4213
rect 10979 4155 10991 4175
rect 11011 4155 11023 4175
rect 2053 3986 2097 3993
rect 2053 3966 2065 3986
rect 2085 3966 2097 3986
rect 2053 3924 2097 3966
rect 3134 3967 3178 4009
rect 3134 3947 3146 3967
rect 3166 3947 3178 3967
rect 3134 3940 3178 3947
rect 3133 3909 3178 3940
rect 3228 3967 3270 4009
rect 3228 3947 3242 3967
rect 3262 3947 3270 3967
rect 3228 3909 3270 3947
rect 3344 3967 3386 4009
rect 3344 3947 3352 3967
rect 3372 3947 3386 3967
rect 3344 3909 3386 3947
rect 3436 3967 3480 4009
rect 3436 3947 3448 3967
rect 3468 3947 3480 3967
rect 3436 3909 3480 3947
rect 3552 3967 3594 4009
rect 3552 3947 3560 3967
rect 3580 3947 3594 3967
rect 3552 3909 3594 3947
rect 3644 3967 3688 4009
rect 3644 3947 3656 3967
rect 3676 3947 3688 3967
rect 3644 3909 3688 3947
rect 3765 3967 3807 4009
rect 3765 3947 3773 3967
rect 3793 3947 3807 3967
rect 3765 3909 3807 3947
rect 3857 3967 3901 4009
rect 10979 4113 11023 4155
rect 11073 4175 11115 4213
rect 11073 4155 11087 4175
rect 11107 4155 11115 4175
rect 11073 4113 11115 4155
rect 11192 4175 11236 4213
rect 11192 4155 11204 4175
rect 11224 4155 11236 4175
rect 11192 4113 11236 4155
rect 11286 4175 11328 4213
rect 11286 4155 11300 4175
rect 11320 4155 11328 4175
rect 11286 4113 11328 4155
rect 11400 4175 11444 4213
rect 11400 4155 11412 4175
rect 11432 4155 11444 4175
rect 11400 4113 11444 4155
rect 11494 4175 11536 4213
rect 11494 4155 11508 4175
rect 11528 4155 11536 4175
rect 11494 4113 11536 4155
rect 11610 4175 11652 4213
rect 11610 4155 11618 4175
rect 11638 4155 11652 4175
rect 11610 4113 11652 4155
rect 11702 4182 11747 4213
rect 14808 4209 14852 4251
rect 14808 4189 14820 4209
rect 14840 4189 14852 4209
rect 14808 4182 14852 4189
rect 11702 4175 11746 4182
rect 11702 4155 11714 4175
rect 11734 4155 11746 4175
rect 11702 4113 11746 4155
rect 14807 4151 14852 4182
rect 14902 4209 14944 4251
rect 14902 4189 14916 4209
rect 14936 4189 14944 4209
rect 14902 4151 14944 4189
rect 15018 4209 15060 4251
rect 15018 4189 15026 4209
rect 15046 4189 15060 4209
rect 15018 4151 15060 4189
rect 15110 4209 15154 4251
rect 15110 4189 15122 4209
rect 15142 4189 15154 4209
rect 15110 4151 15154 4189
rect 15226 4209 15268 4251
rect 15226 4189 15234 4209
rect 15254 4189 15268 4209
rect 15226 4151 15268 4189
rect 15318 4209 15362 4251
rect 15318 4189 15330 4209
rect 15350 4189 15362 4209
rect 15318 4151 15362 4189
rect 15439 4209 15481 4251
rect 15439 4189 15447 4209
rect 15467 4189 15481 4209
rect 15439 4151 15481 4189
rect 15531 4209 15575 4251
rect 15531 4189 15543 4209
rect 15563 4189 15575 4209
rect 15531 4151 15575 4189
rect 3857 3947 3869 3967
rect 3889 3947 3901 3967
rect 6611 3965 6655 4003
rect 3857 3909 3901 3947
rect 6611 3945 6623 3965
rect 6643 3945 6655 3965
rect 6611 3903 6655 3945
rect 6705 3965 6747 4003
rect 6705 3945 6719 3965
rect 6739 3945 6747 3965
rect 6705 3903 6747 3945
rect 6824 3965 6868 4003
rect 6824 3945 6836 3965
rect 6856 3945 6868 3965
rect 6824 3903 6868 3945
rect 6918 3965 6960 4003
rect 6918 3945 6932 3965
rect 6952 3945 6960 3965
rect 6918 3903 6960 3945
rect 7032 3965 7076 4003
rect 7032 3945 7044 3965
rect 7064 3945 7076 3965
rect 7032 3903 7076 3945
rect 7126 3965 7168 4003
rect 7126 3945 7140 3965
rect 7160 3945 7168 3965
rect 7126 3903 7168 3945
rect 7242 3965 7284 4003
rect 7242 3945 7250 3965
rect 7270 3945 7284 3965
rect 7242 3903 7284 3945
rect 7334 3972 7379 4003
rect 16260 4154 16304 4192
rect 16260 4134 16272 4154
rect 16292 4134 16304 4154
rect 11991 3994 12035 4032
rect 7334 3965 7378 3972
rect 7334 3945 7346 3965
rect 7366 3945 7378 3965
rect 7334 3903 7378 3945
rect 8415 3946 8459 3988
rect 8415 3926 8427 3946
rect 8447 3926 8459 3946
rect 8415 3919 8459 3926
rect 317 3752 361 3790
rect 317 3732 329 3752
rect 349 3732 361 3752
rect 317 3690 361 3732
rect 411 3752 453 3790
rect 411 3732 425 3752
rect 445 3732 453 3752
rect 411 3690 453 3732
rect 530 3752 574 3790
rect 530 3732 542 3752
rect 562 3732 574 3752
rect 530 3690 574 3732
rect 624 3752 666 3790
rect 624 3732 638 3752
rect 658 3732 666 3752
rect 624 3690 666 3732
rect 738 3752 782 3790
rect 738 3732 750 3752
rect 770 3732 782 3752
rect 738 3690 782 3732
rect 832 3752 874 3790
rect 832 3732 846 3752
rect 866 3732 874 3752
rect 832 3690 874 3732
rect 948 3752 990 3790
rect 948 3732 956 3752
rect 976 3732 990 3752
rect 948 3690 990 3732
rect 1040 3759 1085 3790
rect 4146 3786 4190 3828
rect 4146 3766 4158 3786
rect 4178 3766 4190 3786
rect 4146 3759 4190 3766
rect 1040 3752 1084 3759
rect 1040 3732 1052 3752
rect 1072 3732 1084 3752
rect 1040 3690 1084 3732
rect 4145 3728 4190 3759
rect 4240 3786 4282 3828
rect 4240 3766 4254 3786
rect 4274 3766 4282 3786
rect 4240 3728 4282 3766
rect 4356 3786 4398 3828
rect 4356 3766 4364 3786
rect 4384 3766 4398 3786
rect 4356 3728 4398 3766
rect 4448 3786 4492 3828
rect 4448 3766 4460 3786
rect 4480 3766 4492 3786
rect 4448 3728 4492 3766
rect 4564 3786 4606 3828
rect 4564 3766 4572 3786
rect 4592 3766 4606 3786
rect 4564 3728 4606 3766
rect 4656 3786 4700 3828
rect 4656 3766 4668 3786
rect 4688 3766 4700 3786
rect 4656 3728 4700 3766
rect 4777 3786 4819 3828
rect 4777 3766 4785 3786
rect 4805 3766 4819 3786
rect 4777 3728 4819 3766
rect 4869 3786 4913 3828
rect 8414 3888 8459 3919
rect 8509 3946 8551 3988
rect 8509 3926 8523 3946
rect 8543 3926 8551 3946
rect 8509 3888 8551 3926
rect 8625 3946 8667 3988
rect 8625 3926 8633 3946
rect 8653 3926 8667 3946
rect 8625 3888 8667 3926
rect 8717 3946 8761 3988
rect 8717 3926 8729 3946
rect 8749 3926 8761 3946
rect 8717 3888 8761 3926
rect 8833 3946 8875 3988
rect 8833 3926 8841 3946
rect 8861 3926 8875 3946
rect 8833 3888 8875 3926
rect 8925 3946 8969 3988
rect 8925 3926 8937 3946
rect 8957 3926 8969 3946
rect 8925 3888 8969 3926
rect 9046 3946 9088 3988
rect 9046 3926 9054 3946
rect 9074 3926 9088 3946
rect 9046 3888 9088 3926
rect 9138 3946 9182 3988
rect 9138 3926 9150 3946
rect 9170 3926 9182 3946
rect 11991 3974 12003 3994
rect 12023 3974 12035 3994
rect 11991 3932 12035 3974
rect 12085 3994 12127 4032
rect 12085 3974 12099 3994
rect 12119 3974 12127 3994
rect 12085 3932 12127 3974
rect 12204 3994 12248 4032
rect 12204 3974 12216 3994
rect 12236 3974 12248 3994
rect 12204 3932 12248 3974
rect 12298 3994 12340 4032
rect 12298 3974 12312 3994
rect 12332 3974 12340 3994
rect 12298 3932 12340 3974
rect 12412 3994 12456 4032
rect 12412 3974 12424 3994
rect 12444 3974 12456 3994
rect 12412 3932 12456 3974
rect 12506 3994 12548 4032
rect 12506 3974 12520 3994
rect 12540 3974 12548 3994
rect 12506 3932 12548 3974
rect 12622 3994 12664 4032
rect 12622 3974 12630 3994
rect 12650 3974 12664 3994
rect 12622 3932 12664 3974
rect 12714 4001 12759 4032
rect 16260 4092 16304 4134
rect 16354 4154 16396 4192
rect 16354 4134 16368 4154
rect 16388 4134 16396 4154
rect 16354 4092 16396 4134
rect 16473 4154 16517 4192
rect 16473 4134 16485 4154
rect 16505 4134 16517 4154
rect 16473 4092 16517 4134
rect 16567 4154 16609 4192
rect 16567 4134 16581 4154
rect 16601 4134 16609 4154
rect 16567 4092 16609 4134
rect 16681 4154 16725 4192
rect 16681 4134 16693 4154
rect 16713 4134 16725 4154
rect 16681 4092 16725 4134
rect 16775 4154 16817 4192
rect 16775 4134 16789 4154
rect 16809 4134 16817 4154
rect 16775 4092 16817 4134
rect 16891 4154 16933 4192
rect 16891 4134 16899 4154
rect 16919 4134 16933 4154
rect 16891 4092 16933 4134
rect 16983 4161 17028 4192
rect 20089 4188 20133 4230
rect 20089 4168 20101 4188
rect 20121 4168 20133 4188
rect 20089 4161 20133 4168
rect 16983 4154 17027 4161
rect 16983 4134 16995 4154
rect 17015 4134 17027 4154
rect 16983 4092 17027 4134
rect 20088 4130 20133 4161
rect 20183 4188 20225 4230
rect 20183 4168 20197 4188
rect 20217 4168 20225 4188
rect 20183 4130 20225 4168
rect 20299 4188 20341 4230
rect 20299 4168 20307 4188
rect 20327 4168 20341 4188
rect 20299 4130 20341 4168
rect 20391 4188 20435 4230
rect 20391 4168 20403 4188
rect 20423 4168 20435 4188
rect 20391 4130 20435 4168
rect 20507 4188 20549 4230
rect 20507 4168 20515 4188
rect 20535 4168 20549 4188
rect 20507 4130 20549 4168
rect 20599 4188 20643 4230
rect 20599 4168 20611 4188
rect 20631 4168 20643 4188
rect 20599 4130 20643 4168
rect 20720 4188 20762 4230
rect 20720 4168 20728 4188
rect 20748 4168 20762 4188
rect 20720 4130 20762 4168
rect 20812 4188 20856 4230
rect 20812 4168 20824 4188
rect 20844 4168 20856 4188
rect 20812 4130 20856 4168
rect 12714 3994 12758 4001
rect 12714 3974 12726 3994
rect 12746 3974 12758 3994
rect 12714 3932 12758 3974
rect 13795 3975 13839 4017
rect 13795 3955 13807 3975
rect 13827 3955 13839 3975
rect 13795 3948 13839 3955
rect 9138 3888 9182 3926
rect 4869 3766 4881 3786
rect 4901 3766 4913 3786
rect 4869 3728 4913 3766
rect 13794 3917 13839 3948
rect 13889 3975 13931 4017
rect 13889 3955 13903 3975
rect 13923 3955 13931 3975
rect 13889 3917 13931 3955
rect 14005 3975 14047 4017
rect 14005 3955 14013 3975
rect 14033 3955 14047 3975
rect 14005 3917 14047 3955
rect 14097 3975 14141 4017
rect 14097 3955 14109 3975
rect 14129 3955 14141 3975
rect 14097 3917 14141 3955
rect 14213 3975 14255 4017
rect 14213 3955 14221 3975
rect 14241 3955 14255 3975
rect 14213 3917 14255 3955
rect 14305 3975 14349 4017
rect 14305 3955 14317 3975
rect 14337 3955 14349 3975
rect 14305 3917 14349 3955
rect 14426 3975 14468 4017
rect 14426 3955 14434 3975
rect 14454 3955 14468 3975
rect 14426 3917 14468 3955
rect 14518 3975 14562 4017
rect 14518 3955 14530 3975
rect 14550 3955 14562 3975
rect 17272 3973 17316 4011
rect 14518 3917 14562 3955
rect 17272 3953 17284 3973
rect 17304 3953 17316 3973
rect 5598 3731 5642 3769
rect 5598 3711 5610 3731
rect 5630 3711 5642 3731
rect 5598 3669 5642 3711
rect 5692 3731 5734 3769
rect 5692 3711 5706 3731
rect 5726 3711 5734 3731
rect 5692 3669 5734 3711
rect 5811 3731 5855 3769
rect 5811 3711 5823 3731
rect 5843 3711 5855 3731
rect 5811 3669 5855 3711
rect 5905 3731 5947 3769
rect 5905 3711 5919 3731
rect 5939 3711 5947 3731
rect 5905 3669 5947 3711
rect 6019 3731 6063 3769
rect 6019 3711 6031 3731
rect 6051 3711 6063 3731
rect 6019 3669 6063 3711
rect 6113 3731 6155 3769
rect 6113 3711 6127 3731
rect 6147 3711 6155 3731
rect 6113 3669 6155 3711
rect 6229 3731 6271 3769
rect 6229 3711 6237 3731
rect 6257 3711 6271 3731
rect 6229 3669 6271 3711
rect 6321 3738 6366 3769
rect 9427 3765 9471 3807
rect 9427 3745 9439 3765
rect 9459 3745 9471 3765
rect 9427 3738 9471 3745
rect 6321 3731 6365 3738
rect 6321 3711 6333 3731
rect 6353 3711 6365 3731
rect 6321 3669 6365 3711
rect 9426 3707 9471 3738
rect 9521 3765 9563 3807
rect 9521 3745 9535 3765
rect 9555 3745 9563 3765
rect 9521 3707 9563 3745
rect 9637 3765 9679 3807
rect 9637 3745 9645 3765
rect 9665 3745 9679 3765
rect 9637 3707 9679 3745
rect 9729 3765 9773 3807
rect 9729 3745 9741 3765
rect 9761 3745 9773 3765
rect 9729 3707 9773 3745
rect 9845 3765 9887 3807
rect 9845 3745 9853 3765
rect 9873 3745 9887 3765
rect 9845 3707 9887 3745
rect 9937 3765 9981 3807
rect 9937 3745 9949 3765
rect 9969 3745 9981 3765
rect 9937 3707 9981 3745
rect 10058 3765 10100 3807
rect 10058 3745 10066 3765
rect 10086 3745 10100 3765
rect 10058 3707 10100 3745
rect 10150 3765 10194 3807
rect 17272 3911 17316 3953
rect 17366 3973 17408 4011
rect 17366 3953 17380 3973
rect 17400 3953 17408 3973
rect 17366 3911 17408 3953
rect 17485 3973 17529 4011
rect 17485 3953 17497 3973
rect 17517 3953 17529 3973
rect 17485 3911 17529 3953
rect 17579 3973 17621 4011
rect 17579 3953 17593 3973
rect 17613 3953 17621 3973
rect 17579 3911 17621 3953
rect 17693 3973 17737 4011
rect 17693 3953 17705 3973
rect 17725 3953 17737 3973
rect 17693 3911 17737 3953
rect 17787 3973 17829 4011
rect 17787 3953 17801 3973
rect 17821 3953 17829 3973
rect 17787 3911 17829 3953
rect 17903 3973 17945 4011
rect 17903 3953 17911 3973
rect 17931 3953 17945 3973
rect 17903 3911 17945 3953
rect 17995 3980 18040 4011
rect 17995 3973 18039 3980
rect 17995 3953 18007 3973
rect 18027 3953 18039 3973
rect 17995 3911 18039 3953
rect 19076 3954 19120 3996
rect 19076 3934 19088 3954
rect 19108 3934 19120 3954
rect 19076 3927 19120 3934
rect 10150 3745 10162 3765
rect 10182 3745 10194 3765
rect 10150 3707 10194 3745
rect 10978 3760 11022 3798
rect 10978 3740 10990 3760
rect 11010 3740 11022 3760
rect 10978 3698 11022 3740
rect 11072 3760 11114 3798
rect 11072 3740 11086 3760
rect 11106 3740 11114 3760
rect 11072 3698 11114 3740
rect 11191 3760 11235 3798
rect 11191 3740 11203 3760
rect 11223 3740 11235 3760
rect 11191 3698 11235 3740
rect 11285 3760 11327 3798
rect 11285 3740 11299 3760
rect 11319 3740 11327 3760
rect 11285 3698 11327 3740
rect 11399 3760 11443 3798
rect 11399 3740 11411 3760
rect 11431 3740 11443 3760
rect 11399 3698 11443 3740
rect 11493 3760 11535 3798
rect 11493 3740 11507 3760
rect 11527 3740 11535 3760
rect 11493 3698 11535 3740
rect 11609 3760 11651 3798
rect 11609 3740 11617 3760
rect 11637 3740 11651 3760
rect 11609 3698 11651 3740
rect 11701 3767 11746 3798
rect 14807 3794 14851 3836
rect 14807 3774 14819 3794
rect 14839 3774 14851 3794
rect 14807 3767 14851 3774
rect 11701 3760 11745 3767
rect 11701 3740 11713 3760
rect 11733 3740 11745 3760
rect 11701 3698 11745 3740
rect 14806 3736 14851 3767
rect 14901 3794 14943 3836
rect 14901 3774 14915 3794
rect 14935 3774 14943 3794
rect 14901 3736 14943 3774
rect 15017 3794 15059 3836
rect 15017 3774 15025 3794
rect 15045 3774 15059 3794
rect 15017 3736 15059 3774
rect 15109 3794 15153 3836
rect 15109 3774 15121 3794
rect 15141 3774 15153 3794
rect 15109 3736 15153 3774
rect 15225 3794 15267 3836
rect 15225 3774 15233 3794
rect 15253 3774 15267 3794
rect 15225 3736 15267 3774
rect 15317 3794 15361 3836
rect 15317 3774 15329 3794
rect 15349 3774 15361 3794
rect 15317 3736 15361 3774
rect 15438 3794 15480 3836
rect 15438 3774 15446 3794
rect 15466 3774 15480 3794
rect 15438 3736 15480 3774
rect 15530 3794 15574 3836
rect 19075 3896 19120 3927
rect 19170 3954 19212 3996
rect 19170 3934 19184 3954
rect 19204 3934 19212 3954
rect 19170 3896 19212 3934
rect 19286 3954 19328 3996
rect 19286 3934 19294 3954
rect 19314 3934 19328 3954
rect 19286 3896 19328 3934
rect 19378 3954 19422 3996
rect 19378 3934 19390 3954
rect 19410 3934 19422 3954
rect 19378 3896 19422 3934
rect 19494 3954 19536 3996
rect 19494 3934 19502 3954
rect 19522 3934 19536 3954
rect 19494 3896 19536 3934
rect 19586 3954 19630 3996
rect 19586 3934 19598 3954
rect 19618 3934 19630 3954
rect 19586 3896 19630 3934
rect 19707 3954 19749 3996
rect 19707 3934 19715 3954
rect 19735 3934 19749 3954
rect 19707 3896 19749 3934
rect 19799 3954 19843 3996
rect 19799 3934 19811 3954
rect 19831 3934 19843 3954
rect 19799 3896 19843 3934
rect 15530 3774 15542 3794
rect 15562 3774 15574 3794
rect 15530 3736 15574 3774
rect 16259 3739 16303 3777
rect 16259 3719 16271 3739
rect 16291 3719 16303 3739
rect 3084 3547 3128 3589
rect 3084 3527 3096 3547
rect 3116 3527 3128 3547
rect 3084 3520 3128 3527
rect 3083 3489 3128 3520
rect 3178 3547 3220 3589
rect 3178 3527 3192 3547
rect 3212 3527 3220 3547
rect 3178 3489 3220 3527
rect 3294 3547 3336 3589
rect 3294 3527 3302 3547
rect 3322 3527 3336 3547
rect 3294 3489 3336 3527
rect 3386 3547 3430 3589
rect 3386 3527 3398 3547
rect 3418 3527 3430 3547
rect 3386 3489 3430 3527
rect 3502 3547 3544 3589
rect 3502 3527 3510 3547
rect 3530 3527 3544 3547
rect 3502 3489 3544 3527
rect 3594 3547 3638 3589
rect 3594 3527 3606 3547
rect 3626 3527 3638 3547
rect 3594 3489 3638 3527
rect 3715 3547 3757 3589
rect 3715 3527 3723 3547
rect 3743 3527 3757 3547
rect 3715 3489 3757 3527
rect 3807 3547 3851 3589
rect 3807 3527 3819 3547
rect 3839 3527 3851 3547
rect 3807 3489 3851 3527
rect 8365 3526 8409 3568
rect 8365 3506 8377 3526
rect 8397 3506 8409 3526
rect 8365 3499 8409 3506
rect 8364 3468 8409 3499
rect 8459 3526 8501 3568
rect 8459 3506 8473 3526
rect 8493 3506 8501 3526
rect 8459 3468 8501 3506
rect 8575 3526 8617 3568
rect 8575 3506 8583 3526
rect 8603 3506 8617 3526
rect 8575 3468 8617 3506
rect 8667 3526 8711 3568
rect 8667 3506 8679 3526
rect 8699 3506 8711 3526
rect 8667 3468 8711 3506
rect 8783 3526 8825 3568
rect 8783 3506 8791 3526
rect 8811 3506 8825 3526
rect 8783 3468 8825 3506
rect 8875 3526 8919 3568
rect 8875 3506 8887 3526
rect 8907 3506 8919 3526
rect 8875 3468 8919 3506
rect 8996 3526 9038 3568
rect 8996 3506 9004 3526
rect 9024 3506 9038 3526
rect 8996 3468 9038 3506
rect 9088 3526 9132 3568
rect 16259 3677 16303 3719
rect 16353 3739 16395 3777
rect 16353 3719 16367 3739
rect 16387 3719 16395 3739
rect 16353 3677 16395 3719
rect 16472 3739 16516 3777
rect 16472 3719 16484 3739
rect 16504 3719 16516 3739
rect 16472 3677 16516 3719
rect 16566 3739 16608 3777
rect 16566 3719 16580 3739
rect 16600 3719 16608 3739
rect 16566 3677 16608 3719
rect 16680 3739 16724 3777
rect 16680 3719 16692 3739
rect 16712 3719 16724 3739
rect 16680 3677 16724 3719
rect 16774 3739 16816 3777
rect 16774 3719 16788 3739
rect 16808 3719 16816 3739
rect 16774 3677 16816 3719
rect 16890 3739 16932 3777
rect 16890 3719 16898 3739
rect 16918 3719 16932 3739
rect 16890 3677 16932 3719
rect 16982 3746 17027 3777
rect 20088 3773 20132 3815
rect 20088 3753 20100 3773
rect 20120 3753 20132 3773
rect 20088 3746 20132 3753
rect 16982 3739 17026 3746
rect 16982 3719 16994 3739
rect 17014 3719 17026 3739
rect 16982 3677 17026 3719
rect 20087 3715 20132 3746
rect 20182 3773 20224 3815
rect 20182 3753 20196 3773
rect 20216 3753 20224 3773
rect 20182 3715 20224 3753
rect 20298 3773 20340 3815
rect 20298 3753 20306 3773
rect 20326 3753 20340 3773
rect 20298 3715 20340 3753
rect 20390 3773 20434 3815
rect 20390 3753 20402 3773
rect 20422 3753 20434 3773
rect 20390 3715 20434 3753
rect 20506 3773 20548 3815
rect 20506 3753 20514 3773
rect 20534 3753 20548 3773
rect 20506 3715 20548 3753
rect 20598 3773 20642 3815
rect 20598 3753 20610 3773
rect 20630 3753 20642 3773
rect 20598 3715 20642 3753
rect 20719 3773 20761 3815
rect 20719 3753 20727 3773
rect 20747 3753 20761 3773
rect 20719 3715 20761 3753
rect 20811 3773 20855 3815
rect 20811 3753 20823 3773
rect 20843 3753 20855 3773
rect 20811 3715 20855 3753
rect 9088 3506 9100 3526
rect 9120 3506 9132 3526
rect 9088 3468 9132 3506
rect 13745 3555 13789 3597
rect 13745 3535 13757 3555
rect 13777 3535 13789 3555
rect 13745 3528 13789 3535
rect 13744 3497 13789 3528
rect 13839 3555 13881 3597
rect 13839 3535 13853 3555
rect 13873 3535 13881 3555
rect 13839 3497 13881 3535
rect 13955 3555 13997 3597
rect 13955 3535 13963 3555
rect 13983 3535 13997 3555
rect 13955 3497 13997 3535
rect 14047 3555 14091 3597
rect 14047 3535 14059 3555
rect 14079 3535 14091 3555
rect 14047 3497 14091 3535
rect 14163 3555 14205 3597
rect 14163 3535 14171 3555
rect 14191 3535 14205 3555
rect 14163 3497 14205 3535
rect 14255 3555 14299 3597
rect 14255 3535 14267 3555
rect 14287 3535 14299 3555
rect 14255 3497 14299 3535
rect 14376 3555 14418 3597
rect 14376 3535 14384 3555
rect 14404 3535 14418 3555
rect 14376 3497 14418 3535
rect 14468 3555 14512 3597
rect 14468 3535 14480 3555
rect 14500 3535 14512 3555
rect 14468 3497 14512 3535
rect 19026 3534 19070 3576
rect 19026 3514 19038 3534
rect 19058 3514 19070 3534
rect 19026 3507 19070 3514
rect 19025 3476 19070 3507
rect 19120 3534 19162 3576
rect 19120 3514 19134 3534
rect 19154 3514 19162 3534
rect 19120 3476 19162 3514
rect 19236 3534 19278 3576
rect 19236 3514 19244 3534
rect 19264 3514 19278 3534
rect 19236 3476 19278 3514
rect 19328 3534 19372 3576
rect 19328 3514 19340 3534
rect 19360 3514 19372 3534
rect 19328 3476 19372 3514
rect 19444 3534 19486 3576
rect 19444 3514 19452 3534
rect 19472 3514 19486 3534
rect 19444 3476 19486 3514
rect 19536 3534 19580 3576
rect 19536 3514 19548 3534
rect 19568 3514 19580 3534
rect 19536 3476 19580 3514
rect 19657 3534 19699 3576
rect 19657 3514 19665 3534
rect 19685 3514 19699 3534
rect 19657 3476 19699 3514
rect 19749 3534 19793 3576
rect 19749 3514 19761 3534
rect 19781 3514 19793 3534
rect 19749 3476 19793 3514
rect 1385 3425 1429 3463
rect 1385 3405 1397 3425
rect 1417 3405 1429 3425
rect 1385 3363 1429 3405
rect 1479 3425 1521 3463
rect 1479 3405 1493 3425
rect 1513 3405 1521 3425
rect 1479 3363 1521 3405
rect 1598 3425 1642 3463
rect 1598 3405 1610 3425
rect 1630 3405 1642 3425
rect 1598 3363 1642 3405
rect 1692 3425 1734 3463
rect 1692 3405 1706 3425
rect 1726 3405 1734 3425
rect 1692 3363 1734 3405
rect 1806 3425 1850 3463
rect 1806 3405 1818 3425
rect 1838 3405 1850 3425
rect 1806 3363 1850 3405
rect 1900 3425 1942 3463
rect 1900 3405 1914 3425
rect 1934 3405 1942 3425
rect 1900 3363 1942 3405
rect 2016 3425 2058 3463
rect 2016 3405 2024 3425
rect 2044 3405 2058 3425
rect 2016 3363 2058 3405
rect 2108 3432 2153 3463
rect 2108 3425 2152 3432
rect 2108 3405 2120 3425
rect 2140 3405 2152 3425
rect 2108 3363 2152 3405
rect 6666 3404 6710 3442
rect 6666 3384 6678 3404
rect 6698 3384 6710 3404
rect 6666 3342 6710 3384
rect 6760 3404 6802 3442
rect 6760 3384 6774 3404
rect 6794 3384 6802 3404
rect 6760 3342 6802 3384
rect 6879 3404 6923 3442
rect 6879 3384 6891 3404
rect 6911 3384 6923 3404
rect 6879 3342 6923 3384
rect 6973 3404 7015 3442
rect 6973 3384 6987 3404
rect 7007 3384 7015 3404
rect 6973 3342 7015 3384
rect 7087 3404 7131 3442
rect 7087 3384 7099 3404
rect 7119 3384 7131 3404
rect 7087 3342 7131 3384
rect 7181 3404 7223 3442
rect 7181 3384 7195 3404
rect 7215 3384 7223 3404
rect 7181 3342 7223 3384
rect 7297 3404 7339 3442
rect 7297 3384 7305 3404
rect 7325 3384 7339 3404
rect 7297 3342 7339 3384
rect 7389 3411 7434 3442
rect 7389 3404 7433 3411
rect 7389 3384 7401 3404
rect 7421 3384 7433 3404
rect 7389 3342 7433 3384
rect 12046 3433 12090 3471
rect 12046 3413 12058 3433
rect 12078 3413 12090 3433
rect 323 3186 367 3224
rect 323 3166 335 3186
rect 355 3166 367 3186
rect 323 3124 367 3166
rect 417 3186 459 3224
rect 417 3166 431 3186
rect 451 3166 459 3186
rect 417 3124 459 3166
rect 536 3186 580 3224
rect 536 3166 548 3186
rect 568 3166 580 3186
rect 536 3124 580 3166
rect 630 3186 672 3224
rect 630 3166 644 3186
rect 664 3166 672 3186
rect 630 3124 672 3166
rect 744 3186 788 3224
rect 744 3166 756 3186
rect 776 3166 788 3186
rect 744 3124 788 3166
rect 838 3186 880 3224
rect 838 3166 852 3186
rect 872 3166 880 3186
rect 838 3124 880 3166
rect 954 3186 996 3224
rect 954 3166 962 3186
rect 982 3166 996 3186
rect 954 3124 996 3166
rect 1046 3193 1091 3224
rect 4152 3220 4196 3262
rect 4152 3200 4164 3220
rect 4184 3200 4196 3220
rect 4152 3193 4196 3200
rect 1046 3186 1090 3193
rect 1046 3166 1058 3186
rect 1078 3166 1090 3186
rect 1046 3124 1090 3166
rect 4151 3162 4196 3193
rect 4246 3220 4288 3262
rect 4246 3200 4260 3220
rect 4280 3200 4288 3220
rect 4246 3162 4288 3200
rect 4362 3220 4404 3262
rect 4362 3200 4370 3220
rect 4390 3200 4404 3220
rect 4362 3162 4404 3200
rect 4454 3220 4498 3262
rect 4454 3200 4466 3220
rect 4486 3200 4498 3220
rect 4454 3162 4498 3200
rect 4570 3220 4612 3262
rect 4570 3200 4578 3220
rect 4598 3200 4612 3220
rect 4570 3162 4612 3200
rect 4662 3220 4706 3262
rect 4662 3200 4674 3220
rect 4694 3200 4706 3220
rect 4662 3162 4706 3200
rect 4783 3220 4825 3262
rect 4783 3200 4791 3220
rect 4811 3200 4825 3220
rect 4783 3162 4825 3200
rect 4875 3220 4919 3262
rect 12046 3371 12090 3413
rect 12140 3433 12182 3471
rect 12140 3413 12154 3433
rect 12174 3413 12182 3433
rect 12140 3371 12182 3413
rect 12259 3433 12303 3471
rect 12259 3413 12271 3433
rect 12291 3413 12303 3433
rect 12259 3371 12303 3413
rect 12353 3433 12395 3471
rect 12353 3413 12367 3433
rect 12387 3413 12395 3433
rect 12353 3371 12395 3413
rect 12467 3433 12511 3471
rect 12467 3413 12479 3433
rect 12499 3413 12511 3433
rect 12467 3371 12511 3413
rect 12561 3433 12603 3471
rect 12561 3413 12575 3433
rect 12595 3413 12603 3433
rect 12561 3371 12603 3413
rect 12677 3433 12719 3471
rect 12677 3413 12685 3433
rect 12705 3413 12719 3433
rect 12677 3371 12719 3413
rect 12769 3440 12814 3471
rect 12769 3433 12813 3440
rect 12769 3413 12781 3433
rect 12801 3413 12813 3433
rect 12769 3371 12813 3413
rect 17327 3412 17371 3450
rect 17327 3392 17339 3412
rect 17359 3392 17371 3412
rect 17327 3350 17371 3392
rect 17421 3412 17463 3450
rect 17421 3392 17435 3412
rect 17455 3392 17463 3412
rect 17421 3350 17463 3392
rect 17540 3412 17584 3450
rect 17540 3392 17552 3412
rect 17572 3392 17584 3412
rect 17540 3350 17584 3392
rect 17634 3412 17676 3450
rect 17634 3392 17648 3412
rect 17668 3392 17676 3412
rect 17634 3350 17676 3392
rect 17748 3412 17792 3450
rect 17748 3392 17760 3412
rect 17780 3392 17792 3412
rect 17748 3350 17792 3392
rect 17842 3412 17884 3450
rect 17842 3392 17856 3412
rect 17876 3392 17884 3412
rect 17842 3350 17884 3392
rect 17958 3412 18000 3450
rect 17958 3392 17966 3412
rect 17986 3392 18000 3412
rect 17958 3350 18000 3392
rect 18050 3419 18095 3450
rect 18050 3412 18094 3419
rect 18050 3392 18062 3412
rect 18082 3392 18094 3412
rect 18050 3350 18094 3392
rect 4875 3200 4887 3220
rect 4907 3200 4919 3220
rect 4875 3162 4919 3200
rect 5604 3165 5648 3203
rect 5604 3145 5616 3165
rect 5636 3145 5648 3165
rect 1335 3005 1379 3043
rect 1335 2985 1347 3005
rect 1367 2985 1379 3005
rect 1335 2943 1379 2985
rect 1429 3005 1471 3043
rect 1429 2985 1443 3005
rect 1463 2985 1471 3005
rect 1429 2943 1471 2985
rect 1548 3005 1592 3043
rect 1548 2985 1560 3005
rect 1580 2985 1592 3005
rect 1548 2943 1592 2985
rect 1642 3005 1684 3043
rect 1642 2985 1656 3005
rect 1676 2985 1684 3005
rect 1642 2943 1684 2985
rect 1756 3005 1800 3043
rect 1756 2985 1768 3005
rect 1788 2985 1800 3005
rect 1756 2943 1800 2985
rect 1850 3005 1892 3043
rect 1850 2985 1864 3005
rect 1884 2985 1892 3005
rect 1850 2943 1892 2985
rect 1966 3005 2008 3043
rect 1966 2985 1974 3005
rect 1994 2985 2008 3005
rect 1966 2943 2008 2985
rect 2058 3012 2103 3043
rect 5604 3103 5648 3145
rect 5698 3165 5740 3203
rect 5698 3145 5712 3165
rect 5732 3145 5740 3165
rect 5698 3103 5740 3145
rect 5817 3165 5861 3203
rect 5817 3145 5829 3165
rect 5849 3145 5861 3165
rect 5817 3103 5861 3145
rect 5911 3165 5953 3203
rect 5911 3145 5925 3165
rect 5945 3145 5953 3165
rect 5911 3103 5953 3145
rect 6025 3165 6069 3203
rect 6025 3145 6037 3165
rect 6057 3145 6069 3165
rect 6025 3103 6069 3145
rect 6119 3165 6161 3203
rect 6119 3145 6133 3165
rect 6153 3145 6161 3165
rect 6119 3103 6161 3145
rect 6235 3165 6277 3203
rect 6235 3145 6243 3165
rect 6263 3145 6277 3165
rect 6235 3103 6277 3145
rect 6327 3172 6372 3203
rect 9433 3199 9477 3241
rect 9433 3179 9445 3199
rect 9465 3179 9477 3199
rect 9433 3172 9477 3179
rect 6327 3165 6371 3172
rect 6327 3145 6339 3165
rect 6359 3145 6371 3165
rect 6327 3103 6371 3145
rect 9432 3141 9477 3172
rect 9527 3199 9569 3241
rect 9527 3179 9541 3199
rect 9561 3179 9569 3199
rect 9527 3141 9569 3179
rect 9643 3199 9685 3241
rect 9643 3179 9651 3199
rect 9671 3179 9685 3199
rect 9643 3141 9685 3179
rect 9735 3199 9779 3241
rect 9735 3179 9747 3199
rect 9767 3179 9779 3199
rect 9735 3141 9779 3179
rect 9851 3199 9893 3241
rect 9851 3179 9859 3199
rect 9879 3179 9893 3199
rect 9851 3141 9893 3179
rect 9943 3199 9987 3241
rect 9943 3179 9955 3199
rect 9975 3179 9987 3199
rect 9943 3141 9987 3179
rect 10064 3199 10106 3241
rect 10064 3179 10072 3199
rect 10092 3179 10106 3199
rect 10064 3141 10106 3179
rect 10156 3199 10200 3241
rect 10156 3179 10168 3199
rect 10188 3179 10200 3199
rect 10156 3141 10200 3179
rect 10984 3194 11028 3232
rect 10984 3174 10996 3194
rect 11016 3174 11028 3194
rect 2058 3005 2102 3012
rect 2058 2985 2070 3005
rect 2090 2985 2102 3005
rect 2058 2943 2102 2985
rect 3139 2986 3183 3028
rect 3139 2966 3151 2986
rect 3171 2966 3183 2986
rect 3139 2959 3183 2966
rect 3138 2928 3183 2959
rect 3233 2986 3275 3028
rect 3233 2966 3247 2986
rect 3267 2966 3275 2986
rect 3233 2928 3275 2966
rect 3349 2986 3391 3028
rect 3349 2966 3357 2986
rect 3377 2966 3391 2986
rect 3349 2928 3391 2966
rect 3441 2986 3485 3028
rect 3441 2966 3453 2986
rect 3473 2966 3485 2986
rect 3441 2928 3485 2966
rect 3557 2986 3599 3028
rect 3557 2966 3565 2986
rect 3585 2966 3599 2986
rect 3557 2928 3599 2966
rect 3649 2986 3693 3028
rect 3649 2966 3661 2986
rect 3681 2966 3693 2986
rect 3649 2928 3693 2966
rect 3770 2986 3812 3028
rect 3770 2966 3778 2986
rect 3798 2966 3812 2986
rect 3770 2928 3812 2966
rect 3862 2986 3906 3028
rect 10984 3132 11028 3174
rect 11078 3194 11120 3232
rect 11078 3174 11092 3194
rect 11112 3174 11120 3194
rect 11078 3132 11120 3174
rect 11197 3194 11241 3232
rect 11197 3174 11209 3194
rect 11229 3174 11241 3194
rect 11197 3132 11241 3174
rect 11291 3194 11333 3232
rect 11291 3174 11305 3194
rect 11325 3174 11333 3194
rect 11291 3132 11333 3174
rect 11405 3194 11449 3232
rect 11405 3174 11417 3194
rect 11437 3174 11449 3194
rect 11405 3132 11449 3174
rect 11499 3194 11541 3232
rect 11499 3174 11513 3194
rect 11533 3174 11541 3194
rect 11499 3132 11541 3174
rect 11615 3194 11657 3232
rect 11615 3174 11623 3194
rect 11643 3174 11657 3194
rect 11615 3132 11657 3174
rect 11707 3201 11752 3232
rect 14813 3228 14857 3270
rect 14813 3208 14825 3228
rect 14845 3208 14857 3228
rect 14813 3201 14857 3208
rect 11707 3194 11751 3201
rect 11707 3174 11719 3194
rect 11739 3174 11751 3194
rect 11707 3132 11751 3174
rect 14812 3170 14857 3201
rect 14907 3228 14949 3270
rect 14907 3208 14921 3228
rect 14941 3208 14949 3228
rect 14907 3170 14949 3208
rect 15023 3228 15065 3270
rect 15023 3208 15031 3228
rect 15051 3208 15065 3228
rect 15023 3170 15065 3208
rect 15115 3228 15159 3270
rect 15115 3208 15127 3228
rect 15147 3208 15159 3228
rect 15115 3170 15159 3208
rect 15231 3228 15273 3270
rect 15231 3208 15239 3228
rect 15259 3208 15273 3228
rect 15231 3170 15273 3208
rect 15323 3228 15367 3270
rect 15323 3208 15335 3228
rect 15355 3208 15367 3228
rect 15323 3170 15367 3208
rect 15444 3228 15486 3270
rect 15444 3208 15452 3228
rect 15472 3208 15486 3228
rect 15444 3170 15486 3208
rect 15536 3228 15580 3270
rect 15536 3208 15548 3228
rect 15568 3208 15580 3228
rect 15536 3170 15580 3208
rect 3862 2966 3874 2986
rect 3894 2966 3906 2986
rect 6616 2984 6660 3022
rect 3862 2928 3906 2966
rect 6616 2964 6628 2984
rect 6648 2964 6660 2984
rect 6616 2922 6660 2964
rect 6710 2984 6752 3022
rect 6710 2964 6724 2984
rect 6744 2964 6752 2984
rect 6710 2922 6752 2964
rect 6829 2984 6873 3022
rect 6829 2964 6841 2984
rect 6861 2964 6873 2984
rect 6829 2922 6873 2964
rect 6923 2984 6965 3022
rect 6923 2964 6937 2984
rect 6957 2964 6965 2984
rect 6923 2922 6965 2964
rect 7037 2984 7081 3022
rect 7037 2964 7049 2984
rect 7069 2964 7081 2984
rect 7037 2922 7081 2964
rect 7131 2984 7173 3022
rect 7131 2964 7145 2984
rect 7165 2964 7173 2984
rect 7131 2922 7173 2964
rect 7247 2984 7289 3022
rect 7247 2964 7255 2984
rect 7275 2964 7289 2984
rect 7247 2922 7289 2964
rect 7339 2991 7384 3022
rect 16265 3173 16309 3211
rect 16265 3153 16277 3173
rect 16297 3153 16309 3173
rect 11996 3013 12040 3051
rect 7339 2984 7383 2991
rect 7339 2964 7351 2984
rect 7371 2964 7383 2984
rect 7339 2922 7383 2964
rect 8420 2965 8464 3007
rect 8420 2945 8432 2965
rect 8452 2945 8464 2965
rect 8420 2938 8464 2945
rect 322 2771 366 2809
rect 322 2751 334 2771
rect 354 2751 366 2771
rect 322 2709 366 2751
rect 416 2771 458 2809
rect 416 2751 430 2771
rect 450 2751 458 2771
rect 416 2709 458 2751
rect 535 2771 579 2809
rect 535 2751 547 2771
rect 567 2751 579 2771
rect 535 2709 579 2751
rect 629 2771 671 2809
rect 629 2751 643 2771
rect 663 2751 671 2771
rect 629 2709 671 2751
rect 743 2771 787 2809
rect 743 2751 755 2771
rect 775 2751 787 2771
rect 743 2709 787 2751
rect 837 2771 879 2809
rect 837 2751 851 2771
rect 871 2751 879 2771
rect 837 2709 879 2751
rect 953 2771 995 2809
rect 953 2751 961 2771
rect 981 2751 995 2771
rect 953 2709 995 2751
rect 1045 2778 1090 2809
rect 4151 2805 4195 2847
rect 4151 2785 4163 2805
rect 4183 2785 4195 2805
rect 4151 2778 4195 2785
rect 1045 2771 1089 2778
rect 1045 2751 1057 2771
rect 1077 2751 1089 2771
rect 1045 2709 1089 2751
rect 4150 2747 4195 2778
rect 4245 2805 4287 2847
rect 4245 2785 4259 2805
rect 4279 2785 4287 2805
rect 4245 2747 4287 2785
rect 4361 2805 4403 2847
rect 4361 2785 4369 2805
rect 4389 2785 4403 2805
rect 4361 2747 4403 2785
rect 4453 2805 4497 2847
rect 4453 2785 4465 2805
rect 4485 2785 4497 2805
rect 4453 2747 4497 2785
rect 4569 2805 4611 2847
rect 4569 2785 4577 2805
rect 4597 2785 4611 2805
rect 4569 2747 4611 2785
rect 4661 2805 4705 2847
rect 4661 2785 4673 2805
rect 4693 2785 4705 2805
rect 4661 2747 4705 2785
rect 4782 2805 4824 2847
rect 4782 2785 4790 2805
rect 4810 2785 4824 2805
rect 4782 2747 4824 2785
rect 4874 2805 4918 2847
rect 8419 2907 8464 2938
rect 8514 2965 8556 3007
rect 8514 2945 8528 2965
rect 8548 2945 8556 2965
rect 8514 2907 8556 2945
rect 8630 2965 8672 3007
rect 8630 2945 8638 2965
rect 8658 2945 8672 2965
rect 8630 2907 8672 2945
rect 8722 2965 8766 3007
rect 8722 2945 8734 2965
rect 8754 2945 8766 2965
rect 8722 2907 8766 2945
rect 8838 2965 8880 3007
rect 8838 2945 8846 2965
rect 8866 2945 8880 2965
rect 8838 2907 8880 2945
rect 8930 2965 8974 3007
rect 8930 2945 8942 2965
rect 8962 2945 8974 2965
rect 8930 2907 8974 2945
rect 9051 2965 9093 3007
rect 9051 2945 9059 2965
rect 9079 2945 9093 2965
rect 9051 2907 9093 2945
rect 9143 2965 9187 3007
rect 9143 2945 9155 2965
rect 9175 2945 9187 2965
rect 11996 2993 12008 3013
rect 12028 2993 12040 3013
rect 11996 2951 12040 2993
rect 12090 3013 12132 3051
rect 12090 2993 12104 3013
rect 12124 2993 12132 3013
rect 12090 2951 12132 2993
rect 12209 3013 12253 3051
rect 12209 2993 12221 3013
rect 12241 2993 12253 3013
rect 12209 2951 12253 2993
rect 12303 3013 12345 3051
rect 12303 2993 12317 3013
rect 12337 2993 12345 3013
rect 12303 2951 12345 2993
rect 12417 3013 12461 3051
rect 12417 2993 12429 3013
rect 12449 2993 12461 3013
rect 12417 2951 12461 2993
rect 12511 3013 12553 3051
rect 12511 2993 12525 3013
rect 12545 2993 12553 3013
rect 12511 2951 12553 2993
rect 12627 3013 12669 3051
rect 12627 2993 12635 3013
rect 12655 2993 12669 3013
rect 12627 2951 12669 2993
rect 12719 3020 12764 3051
rect 16265 3111 16309 3153
rect 16359 3173 16401 3211
rect 16359 3153 16373 3173
rect 16393 3153 16401 3173
rect 16359 3111 16401 3153
rect 16478 3173 16522 3211
rect 16478 3153 16490 3173
rect 16510 3153 16522 3173
rect 16478 3111 16522 3153
rect 16572 3173 16614 3211
rect 16572 3153 16586 3173
rect 16606 3153 16614 3173
rect 16572 3111 16614 3153
rect 16686 3173 16730 3211
rect 16686 3153 16698 3173
rect 16718 3153 16730 3173
rect 16686 3111 16730 3153
rect 16780 3173 16822 3211
rect 16780 3153 16794 3173
rect 16814 3153 16822 3173
rect 16780 3111 16822 3153
rect 16896 3173 16938 3211
rect 16896 3153 16904 3173
rect 16924 3153 16938 3173
rect 16896 3111 16938 3153
rect 16988 3180 17033 3211
rect 20094 3207 20138 3249
rect 20094 3187 20106 3207
rect 20126 3187 20138 3207
rect 20094 3180 20138 3187
rect 16988 3173 17032 3180
rect 16988 3153 17000 3173
rect 17020 3153 17032 3173
rect 16988 3111 17032 3153
rect 20093 3149 20138 3180
rect 20188 3207 20230 3249
rect 20188 3187 20202 3207
rect 20222 3187 20230 3207
rect 20188 3149 20230 3187
rect 20304 3207 20346 3249
rect 20304 3187 20312 3207
rect 20332 3187 20346 3207
rect 20304 3149 20346 3187
rect 20396 3207 20440 3249
rect 20396 3187 20408 3207
rect 20428 3187 20440 3207
rect 20396 3149 20440 3187
rect 20512 3207 20554 3249
rect 20512 3187 20520 3207
rect 20540 3187 20554 3207
rect 20512 3149 20554 3187
rect 20604 3207 20648 3249
rect 20604 3187 20616 3207
rect 20636 3187 20648 3207
rect 20604 3149 20648 3187
rect 20725 3207 20767 3249
rect 20725 3187 20733 3207
rect 20753 3187 20767 3207
rect 20725 3149 20767 3187
rect 20817 3207 20861 3249
rect 20817 3187 20829 3207
rect 20849 3187 20861 3207
rect 20817 3149 20861 3187
rect 12719 3013 12763 3020
rect 12719 2993 12731 3013
rect 12751 2993 12763 3013
rect 12719 2951 12763 2993
rect 13800 2994 13844 3036
rect 13800 2974 13812 2994
rect 13832 2974 13844 2994
rect 13800 2967 13844 2974
rect 9143 2907 9187 2945
rect 4874 2785 4886 2805
rect 4906 2785 4918 2805
rect 4874 2747 4918 2785
rect 13799 2936 13844 2967
rect 13894 2994 13936 3036
rect 13894 2974 13908 2994
rect 13928 2974 13936 2994
rect 13894 2936 13936 2974
rect 14010 2994 14052 3036
rect 14010 2974 14018 2994
rect 14038 2974 14052 2994
rect 14010 2936 14052 2974
rect 14102 2994 14146 3036
rect 14102 2974 14114 2994
rect 14134 2974 14146 2994
rect 14102 2936 14146 2974
rect 14218 2994 14260 3036
rect 14218 2974 14226 2994
rect 14246 2974 14260 2994
rect 14218 2936 14260 2974
rect 14310 2994 14354 3036
rect 14310 2974 14322 2994
rect 14342 2974 14354 2994
rect 14310 2936 14354 2974
rect 14431 2994 14473 3036
rect 14431 2974 14439 2994
rect 14459 2974 14473 2994
rect 14431 2936 14473 2974
rect 14523 2994 14567 3036
rect 14523 2974 14535 2994
rect 14555 2974 14567 2994
rect 17277 2992 17321 3030
rect 14523 2936 14567 2974
rect 17277 2972 17289 2992
rect 17309 2972 17321 2992
rect 5603 2750 5647 2788
rect 5603 2730 5615 2750
rect 5635 2730 5647 2750
rect 5603 2688 5647 2730
rect 5697 2750 5739 2788
rect 5697 2730 5711 2750
rect 5731 2730 5739 2750
rect 5697 2688 5739 2730
rect 5816 2750 5860 2788
rect 5816 2730 5828 2750
rect 5848 2730 5860 2750
rect 5816 2688 5860 2730
rect 5910 2750 5952 2788
rect 5910 2730 5924 2750
rect 5944 2730 5952 2750
rect 5910 2688 5952 2730
rect 6024 2750 6068 2788
rect 6024 2730 6036 2750
rect 6056 2730 6068 2750
rect 6024 2688 6068 2730
rect 6118 2750 6160 2788
rect 6118 2730 6132 2750
rect 6152 2730 6160 2750
rect 6118 2688 6160 2730
rect 6234 2750 6276 2788
rect 6234 2730 6242 2750
rect 6262 2730 6276 2750
rect 6234 2688 6276 2730
rect 6326 2757 6371 2788
rect 9432 2784 9476 2826
rect 9432 2764 9444 2784
rect 9464 2764 9476 2784
rect 9432 2757 9476 2764
rect 6326 2750 6370 2757
rect 6326 2730 6338 2750
rect 6358 2730 6370 2750
rect 6326 2688 6370 2730
rect 9431 2726 9476 2757
rect 9526 2784 9568 2826
rect 9526 2764 9540 2784
rect 9560 2764 9568 2784
rect 9526 2726 9568 2764
rect 9642 2784 9684 2826
rect 9642 2764 9650 2784
rect 9670 2764 9684 2784
rect 9642 2726 9684 2764
rect 9734 2784 9778 2826
rect 9734 2764 9746 2784
rect 9766 2764 9778 2784
rect 9734 2726 9778 2764
rect 9850 2784 9892 2826
rect 9850 2764 9858 2784
rect 9878 2764 9892 2784
rect 9850 2726 9892 2764
rect 9942 2784 9986 2826
rect 9942 2764 9954 2784
rect 9974 2764 9986 2784
rect 9942 2726 9986 2764
rect 10063 2784 10105 2826
rect 10063 2764 10071 2784
rect 10091 2764 10105 2784
rect 10063 2726 10105 2764
rect 10155 2784 10199 2826
rect 17277 2930 17321 2972
rect 17371 2992 17413 3030
rect 17371 2972 17385 2992
rect 17405 2972 17413 2992
rect 17371 2930 17413 2972
rect 17490 2992 17534 3030
rect 17490 2972 17502 2992
rect 17522 2972 17534 2992
rect 17490 2930 17534 2972
rect 17584 2992 17626 3030
rect 17584 2972 17598 2992
rect 17618 2972 17626 2992
rect 17584 2930 17626 2972
rect 17698 2992 17742 3030
rect 17698 2972 17710 2992
rect 17730 2972 17742 2992
rect 17698 2930 17742 2972
rect 17792 2992 17834 3030
rect 17792 2972 17806 2992
rect 17826 2972 17834 2992
rect 17792 2930 17834 2972
rect 17908 2992 17950 3030
rect 17908 2972 17916 2992
rect 17936 2972 17950 2992
rect 17908 2930 17950 2972
rect 18000 2999 18045 3030
rect 18000 2992 18044 2999
rect 18000 2972 18012 2992
rect 18032 2972 18044 2992
rect 18000 2930 18044 2972
rect 19081 2973 19125 3015
rect 19081 2953 19093 2973
rect 19113 2953 19125 2973
rect 19081 2946 19125 2953
rect 10155 2764 10167 2784
rect 10187 2764 10199 2784
rect 10155 2726 10199 2764
rect 10983 2779 11027 2817
rect 10983 2759 10995 2779
rect 11015 2759 11027 2779
rect 10983 2717 11027 2759
rect 11077 2779 11119 2817
rect 11077 2759 11091 2779
rect 11111 2759 11119 2779
rect 11077 2717 11119 2759
rect 11196 2779 11240 2817
rect 11196 2759 11208 2779
rect 11228 2759 11240 2779
rect 11196 2717 11240 2759
rect 11290 2779 11332 2817
rect 11290 2759 11304 2779
rect 11324 2759 11332 2779
rect 11290 2717 11332 2759
rect 11404 2779 11448 2817
rect 11404 2759 11416 2779
rect 11436 2759 11448 2779
rect 11404 2717 11448 2759
rect 11498 2779 11540 2817
rect 11498 2759 11512 2779
rect 11532 2759 11540 2779
rect 11498 2717 11540 2759
rect 11614 2779 11656 2817
rect 11614 2759 11622 2779
rect 11642 2759 11656 2779
rect 11614 2717 11656 2759
rect 11706 2786 11751 2817
rect 14812 2813 14856 2855
rect 14812 2793 14824 2813
rect 14844 2793 14856 2813
rect 14812 2786 14856 2793
rect 11706 2779 11750 2786
rect 11706 2759 11718 2779
rect 11738 2759 11750 2779
rect 11706 2717 11750 2759
rect 14811 2755 14856 2786
rect 14906 2813 14948 2855
rect 14906 2793 14920 2813
rect 14940 2793 14948 2813
rect 14906 2755 14948 2793
rect 15022 2813 15064 2855
rect 15022 2793 15030 2813
rect 15050 2793 15064 2813
rect 15022 2755 15064 2793
rect 15114 2813 15158 2855
rect 15114 2793 15126 2813
rect 15146 2793 15158 2813
rect 15114 2755 15158 2793
rect 15230 2813 15272 2855
rect 15230 2793 15238 2813
rect 15258 2793 15272 2813
rect 15230 2755 15272 2793
rect 15322 2813 15366 2855
rect 15322 2793 15334 2813
rect 15354 2793 15366 2813
rect 15322 2755 15366 2793
rect 15443 2813 15485 2855
rect 15443 2793 15451 2813
rect 15471 2793 15485 2813
rect 15443 2755 15485 2793
rect 15535 2813 15579 2855
rect 19080 2915 19125 2946
rect 19175 2973 19217 3015
rect 19175 2953 19189 2973
rect 19209 2953 19217 2973
rect 19175 2915 19217 2953
rect 19291 2973 19333 3015
rect 19291 2953 19299 2973
rect 19319 2953 19333 2973
rect 19291 2915 19333 2953
rect 19383 2973 19427 3015
rect 19383 2953 19395 2973
rect 19415 2953 19427 2973
rect 19383 2915 19427 2953
rect 19499 2973 19541 3015
rect 19499 2953 19507 2973
rect 19527 2953 19541 2973
rect 19499 2915 19541 2953
rect 19591 2973 19635 3015
rect 19591 2953 19603 2973
rect 19623 2953 19635 2973
rect 19591 2915 19635 2953
rect 19712 2973 19754 3015
rect 19712 2953 19720 2973
rect 19740 2953 19754 2973
rect 19712 2915 19754 2953
rect 19804 2973 19848 3015
rect 19804 2953 19816 2973
rect 19836 2953 19848 2973
rect 19804 2915 19848 2953
rect 15535 2793 15547 2813
rect 15567 2793 15579 2813
rect 15535 2755 15579 2793
rect 16264 2758 16308 2796
rect 16264 2738 16276 2758
rect 16296 2738 16308 2758
rect 1550 2493 1594 2531
rect 1550 2473 1562 2493
rect 1582 2473 1594 2493
rect 1550 2431 1594 2473
rect 1644 2493 1686 2531
rect 1644 2473 1658 2493
rect 1678 2473 1686 2493
rect 1644 2431 1686 2473
rect 1763 2493 1807 2531
rect 1763 2473 1775 2493
rect 1795 2473 1807 2493
rect 1763 2431 1807 2473
rect 1857 2493 1899 2531
rect 1857 2473 1871 2493
rect 1891 2473 1899 2493
rect 1857 2431 1899 2473
rect 1971 2493 2015 2531
rect 1971 2473 1983 2493
rect 2003 2473 2015 2493
rect 1971 2431 2015 2473
rect 2065 2493 2107 2531
rect 2065 2473 2079 2493
rect 2099 2473 2107 2493
rect 2065 2431 2107 2473
rect 2181 2493 2223 2531
rect 2181 2473 2189 2493
rect 2209 2473 2223 2493
rect 2181 2431 2223 2473
rect 2273 2500 2318 2531
rect 2931 2519 2975 2561
rect 2273 2493 2317 2500
rect 2273 2473 2285 2493
rect 2305 2473 2317 2493
rect 2931 2499 2943 2519
rect 2963 2499 2975 2519
rect 2931 2492 2975 2499
rect 2273 2431 2317 2473
rect 2930 2461 2975 2492
rect 3025 2519 3067 2561
rect 3025 2499 3039 2519
rect 3059 2499 3067 2519
rect 3025 2461 3067 2499
rect 3141 2519 3183 2561
rect 3141 2499 3149 2519
rect 3169 2499 3183 2519
rect 3141 2461 3183 2499
rect 3233 2519 3277 2561
rect 3233 2499 3245 2519
rect 3265 2499 3277 2519
rect 3233 2461 3277 2499
rect 3349 2519 3391 2561
rect 3349 2499 3357 2519
rect 3377 2499 3391 2519
rect 3349 2461 3391 2499
rect 3441 2519 3485 2561
rect 3441 2499 3453 2519
rect 3473 2499 3485 2519
rect 3441 2461 3485 2499
rect 3562 2519 3604 2561
rect 3562 2499 3570 2519
rect 3590 2499 3604 2519
rect 3562 2461 3604 2499
rect 3654 2519 3698 2561
rect 16264 2696 16308 2738
rect 16358 2758 16400 2796
rect 16358 2738 16372 2758
rect 16392 2738 16400 2758
rect 16358 2696 16400 2738
rect 16477 2758 16521 2796
rect 16477 2738 16489 2758
rect 16509 2738 16521 2758
rect 16477 2696 16521 2738
rect 16571 2758 16613 2796
rect 16571 2738 16585 2758
rect 16605 2738 16613 2758
rect 16571 2696 16613 2738
rect 16685 2758 16729 2796
rect 16685 2738 16697 2758
rect 16717 2738 16729 2758
rect 16685 2696 16729 2738
rect 16779 2758 16821 2796
rect 16779 2738 16793 2758
rect 16813 2738 16821 2758
rect 16779 2696 16821 2738
rect 16895 2758 16937 2796
rect 16895 2738 16903 2758
rect 16923 2738 16937 2758
rect 16895 2696 16937 2738
rect 16987 2765 17032 2796
rect 20093 2792 20137 2834
rect 20093 2772 20105 2792
rect 20125 2772 20137 2792
rect 20093 2765 20137 2772
rect 16987 2758 17031 2765
rect 16987 2738 16999 2758
rect 17019 2738 17031 2758
rect 16987 2696 17031 2738
rect 20092 2734 20137 2765
rect 20187 2792 20229 2834
rect 20187 2772 20201 2792
rect 20221 2772 20229 2792
rect 20187 2734 20229 2772
rect 20303 2792 20345 2834
rect 20303 2772 20311 2792
rect 20331 2772 20345 2792
rect 20303 2734 20345 2772
rect 20395 2792 20439 2834
rect 20395 2772 20407 2792
rect 20427 2772 20439 2792
rect 20395 2734 20439 2772
rect 20511 2792 20553 2834
rect 20511 2772 20519 2792
rect 20539 2772 20553 2792
rect 20511 2734 20553 2772
rect 20603 2792 20647 2834
rect 20603 2772 20615 2792
rect 20635 2772 20647 2792
rect 20603 2734 20647 2772
rect 20724 2792 20766 2834
rect 20724 2772 20732 2792
rect 20752 2772 20766 2792
rect 20724 2734 20766 2772
rect 20816 2792 20860 2834
rect 20816 2772 20828 2792
rect 20848 2772 20860 2792
rect 20816 2734 20860 2772
rect 3654 2499 3666 2519
rect 3686 2499 3698 2519
rect 3654 2461 3698 2499
rect 6831 2472 6875 2510
rect 6831 2452 6843 2472
rect 6863 2452 6875 2472
rect 6831 2410 6875 2452
rect 6925 2472 6967 2510
rect 6925 2452 6939 2472
rect 6959 2452 6967 2472
rect 6925 2410 6967 2452
rect 7044 2472 7088 2510
rect 7044 2452 7056 2472
rect 7076 2452 7088 2472
rect 7044 2410 7088 2452
rect 7138 2472 7180 2510
rect 7138 2452 7152 2472
rect 7172 2452 7180 2472
rect 7138 2410 7180 2452
rect 7252 2472 7296 2510
rect 7252 2452 7264 2472
rect 7284 2452 7296 2472
rect 7252 2410 7296 2452
rect 7346 2472 7388 2510
rect 7346 2452 7360 2472
rect 7380 2452 7388 2472
rect 7346 2410 7388 2452
rect 7462 2472 7504 2510
rect 7462 2452 7470 2472
rect 7490 2452 7504 2472
rect 7462 2410 7504 2452
rect 7554 2479 7599 2510
rect 8212 2498 8256 2540
rect 7554 2472 7598 2479
rect 7554 2452 7566 2472
rect 7586 2452 7598 2472
rect 8212 2478 8224 2498
rect 8244 2478 8256 2498
rect 8212 2471 8256 2478
rect 7554 2410 7598 2452
rect 8211 2440 8256 2471
rect 8306 2498 8348 2540
rect 8306 2478 8320 2498
rect 8340 2478 8348 2498
rect 8306 2440 8348 2478
rect 8422 2498 8464 2540
rect 8422 2478 8430 2498
rect 8450 2478 8464 2498
rect 8422 2440 8464 2478
rect 8514 2498 8558 2540
rect 8514 2478 8526 2498
rect 8546 2478 8558 2498
rect 8514 2440 8558 2478
rect 8630 2498 8672 2540
rect 8630 2478 8638 2498
rect 8658 2478 8672 2498
rect 8630 2440 8672 2478
rect 8722 2498 8766 2540
rect 8722 2478 8734 2498
rect 8754 2478 8766 2498
rect 8722 2440 8766 2478
rect 8843 2498 8885 2540
rect 8843 2478 8851 2498
rect 8871 2478 8885 2498
rect 8843 2440 8885 2478
rect 8935 2498 8979 2540
rect 8935 2478 8947 2498
rect 8967 2478 8979 2498
rect 8935 2440 8979 2478
rect 12211 2501 12255 2539
rect 12211 2481 12223 2501
rect 12243 2481 12255 2501
rect 12211 2439 12255 2481
rect 12305 2501 12347 2539
rect 12305 2481 12319 2501
rect 12339 2481 12347 2501
rect 12305 2439 12347 2481
rect 12424 2501 12468 2539
rect 12424 2481 12436 2501
rect 12456 2481 12468 2501
rect 12424 2439 12468 2481
rect 12518 2501 12560 2539
rect 12518 2481 12532 2501
rect 12552 2481 12560 2501
rect 12518 2439 12560 2481
rect 12632 2501 12676 2539
rect 12632 2481 12644 2501
rect 12664 2481 12676 2501
rect 12632 2439 12676 2481
rect 12726 2501 12768 2539
rect 12726 2481 12740 2501
rect 12760 2481 12768 2501
rect 12726 2439 12768 2481
rect 12842 2501 12884 2539
rect 12842 2481 12850 2501
rect 12870 2481 12884 2501
rect 12842 2439 12884 2481
rect 12934 2508 12979 2539
rect 13592 2527 13636 2569
rect 12934 2501 12978 2508
rect 12934 2481 12946 2501
rect 12966 2481 12978 2501
rect 13592 2507 13604 2527
rect 13624 2507 13636 2527
rect 13592 2500 13636 2507
rect 12934 2439 12978 2481
rect 13591 2469 13636 2500
rect 13686 2527 13728 2569
rect 13686 2507 13700 2527
rect 13720 2507 13728 2527
rect 13686 2469 13728 2507
rect 13802 2527 13844 2569
rect 13802 2507 13810 2527
rect 13830 2507 13844 2527
rect 13802 2469 13844 2507
rect 13894 2527 13938 2569
rect 13894 2507 13906 2527
rect 13926 2507 13938 2527
rect 13894 2469 13938 2507
rect 14010 2527 14052 2569
rect 14010 2507 14018 2527
rect 14038 2507 14052 2527
rect 14010 2469 14052 2507
rect 14102 2527 14146 2569
rect 14102 2507 14114 2527
rect 14134 2507 14146 2527
rect 14102 2469 14146 2507
rect 14223 2527 14265 2569
rect 14223 2507 14231 2527
rect 14251 2507 14265 2527
rect 14223 2469 14265 2507
rect 14315 2527 14359 2569
rect 14315 2507 14327 2527
rect 14347 2507 14359 2527
rect 14315 2469 14359 2507
rect 17492 2480 17536 2518
rect 17492 2460 17504 2480
rect 17524 2460 17536 2480
rect 330 2207 374 2245
rect 330 2187 342 2207
rect 362 2187 374 2207
rect 330 2145 374 2187
rect 424 2207 466 2245
rect 424 2187 438 2207
rect 458 2187 466 2207
rect 424 2145 466 2187
rect 543 2207 587 2245
rect 543 2187 555 2207
rect 575 2187 587 2207
rect 543 2145 587 2187
rect 637 2207 679 2245
rect 637 2187 651 2207
rect 671 2187 679 2207
rect 637 2145 679 2187
rect 751 2207 795 2245
rect 751 2187 763 2207
rect 783 2187 795 2207
rect 751 2145 795 2187
rect 845 2207 887 2245
rect 845 2187 859 2207
rect 879 2187 887 2207
rect 845 2145 887 2187
rect 961 2207 1003 2245
rect 961 2187 969 2207
rect 989 2187 1003 2207
rect 961 2145 1003 2187
rect 1053 2214 1098 2245
rect 4159 2241 4203 2283
rect 4159 2221 4171 2241
rect 4191 2221 4203 2241
rect 4159 2214 4203 2221
rect 1053 2207 1097 2214
rect 1053 2187 1065 2207
rect 1085 2187 1097 2207
rect 1053 2145 1097 2187
rect 4158 2183 4203 2214
rect 4253 2241 4295 2283
rect 4253 2221 4267 2241
rect 4287 2221 4295 2241
rect 4253 2183 4295 2221
rect 4369 2241 4411 2283
rect 4369 2221 4377 2241
rect 4397 2221 4411 2241
rect 4369 2183 4411 2221
rect 4461 2241 4505 2283
rect 4461 2221 4473 2241
rect 4493 2221 4505 2241
rect 4461 2183 4505 2221
rect 4577 2241 4619 2283
rect 4577 2221 4585 2241
rect 4605 2221 4619 2241
rect 4577 2183 4619 2221
rect 4669 2241 4713 2283
rect 4669 2221 4681 2241
rect 4701 2221 4713 2241
rect 4669 2183 4713 2221
rect 4790 2241 4832 2283
rect 4790 2221 4798 2241
rect 4818 2221 4832 2241
rect 4790 2183 4832 2221
rect 4882 2241 4926 2283
rect 17492 2418 17536 2460
rect 17586 2480 17628 2518
rect 17586 2460 17600 2480
rect 17620 2460 17628 2480
rect 17586 2418 17628 2460
rect 17705 2480 17749 2518
rect 17705 2460 17717 2480
rect 17737 2460 17749 2480
rect 17705 2418 17749 2460
rect 17799 2480 17841 2518
rect 17799 2460 17813 2480
rect 17833 2460 17841 2480
rect 17799 2418 17841 2460
rect 17913 2480 17957 2518
rect 17913 2460 17925 2480
rect 17945 2460 17957 2480
rect 17913 2418 17957 2460
rect 18007 2480 18049 2518
rect 18007 2460 18021 2480
rect 18041 2460 18049 2480
rect 18007 2418 18049 2460
rect 18123 2480 18165 2518
rect 18123 2460 18131 2480
rect 18151 2460 18165 2480
rect 18123 2418 18165 2460
rect 18215 2487 18260 2518
rect 18873 2506 18917 2548
rect 18215 2480 18259 2487
rect 18215 2460 18227 2480
rect 18247 2460 18259 2480
rect 18873 2486 18885 2506
rect 18905 2486 18917 2506
rect 18873 2479 18917 2486
rect 18215 2418 18259 2460
rect 18872 2448 18917 2479
rect 18967 2506 19009 2548
rect 18967 2486 18981 2506
rect 19001 2486 19009 2506
rect 18967 2448 19009 2486
rect 19083 2506 19125 2548
rect 19083 2486 19091 2506
rect 19111 2486 19125 2506
rect 19083 2448 19125 2486
rect 19175 2506 19219 2548
rect 19175 2486 19187 2506
rect 19207 2486 19219 2506
rect 19175 2448 19219 2486
rect 19291 2506 19333 2548
rect 19291 2486 19299 2506
rect 19319 2486 19333 2506
rect 19291 2448 19333 2486
rect 19383 2506 19427 2548
rect 19383 2486 19395 2506
rect 19415 2486 19427 2506
rect 19383 2448 19427 2486
rect 19504 2506 19546 2548
rect 19504 2486 19512 2506
rect 19532 2486 19546 2506
rect 19504 2448 19546 2486
rect 19596 2506 19640 2548
rect 19596 2486 19608 2506
rect 19628 2486 19640 2506
rect 19596 2448 19640 2486
rect 4882 2221 4894 2241
rect 4914 2221 4926 2241
rect 4882 2183 4926 2221
rect 5611 2186 5655 2224
rect 5611 2166 5623 2186
rect 5643 2166 5655 2186
rect 1342 2026 1386 2064
rect 1342 2006 1354 2026
rect 1374 2006 1386 2026
rect 1342 1964 1386 2006
rect 1436 2026 1478 2064
rect 1436 2006 1450 2026
rect 1470 2006 1478 2026
rect 1436 1964 1478 2006
rect 1555 2026 1599 2064
rect 1555 2006 1567 2026
rect 1587 2006 1599 2026
rect 1555 1964 1599 2006
rect 1649 2026 1691 2064
rect 1649 2006 1663 2026
rect 1683 2006 1691 2026
rect 1649 1964 1691 2006
rect 1763 2026 1807 2064
rect 1763 2006 1775 2026
rect 1795 2006 1807 2026
rect 1763 1964 1807 2006
rect 1857 2026 1899 2064
rect 1857 2006 1871 2026
rect 1891 2006 1899 2026
rect 1857 1964 1899 2006
rect 1973 2026 2015 2064
rect 1973 2006 1981 2026
rect 2001 2006 2015 2026
rect 1973 1964 2015 2006
rect 2065 2033 2110 2064
rect 5611 2124 5655 2166
rect 5705 2186 5747 2224
rect 5705 2166 5719 2186
rect 5739 2166 5747 2186
rect 5705 2124 5747 2166
rect 5824 2186 5868 2224
rect 5824 2166 5836 2186
rect 5856 2166 5868 2186
rect 5824 2124 5868 2166
rect 5918 2186 5960 2224
rect 5918 2166 5932 2186
rect 5952 2166 5960 2186
rect 5918 2124 5960 2166
rect 6032 2186 6076 2224
rect 6032 2166 6044 2186
rect 6064 2166 6076 2186
rect 6032 2124 6076 2166
rect 6126 2186 6168 2224
rect 6126 2166 6140 2186
rect 6160 2166 6168 2186
rect 6126 2124 6168 2166
rect 6242 2186 6284 2224
rect 6242 2166 6250 2186
rect 6270 2166 6284 2186
rect 6242 2124 6284 2166
rect 6334 2193 6379 2224
rect 9440 2220 9484 2262
rect 9440 2200 9452 2220
rect 9472 2200 9484 2220
rect 9440 2193 9484 2200
rect 6334 2186 6378 2193
rect 6334 2166 6346 2186
rect 6366 2166 6378 2186
rect 6334 2124 6378 2166
rect 9439 2162 9484 2193
rect 9534 2220 9576 2262
rect 9534 2200 9548 2220
rect 9568 2200 9576 2220
rect 9534 2162 9576 2200
rect 9650 2220 9692 2262
rect 9650 2200 9658 2220
rect 9678 2200 9692 2220
rect 9650 2162 9692 2200
rect 9742 2220 9786 2262
rect 9742 2200 9754 2220
rect 9774 2200 9786 2220
rect 9742 2162 9786 2200
rect 9858 2220 9900 2262
rect 9858 2200 9866 2220
rect 9886 2200 9900 2220
rect 9858 2162 9900 2200
rect 9950 2220 9994 2262
rect 9950 2200 9962 2220
rect 9982 2200 9994 2220
rect 9950 2162 9994 2200
rect 10071 2220 10113 2262
rect 10071 2200 10079 2220
rect 10099 2200 10113 2220
rect 10071 2162 10113 2200
rect 10163 2220 10207 2262
rect 10163 2200 10175 2220
rect 10195 2200 10207 2220
rect 10163 2162 10207 2200
rect 10991 2215 11035 2253
rect 10991 2195 11003 2215
rect 11023 2195 11035 2215
rect 2065 2026 2109 2033
rect 2065 2006 2077 2026
rect 2097 2006 2109 2026
rect 2065 1964 2109 2006
rect 3146 2007 3190 2049
rect 3146 1987 3158 2007
rect 3178 1987 3190 2007
rect 3146 1980 3190 1987
rect 3145 1949 3190 1980
rect 3240 2007 3282 2049
rect 3240 1987 3254 2007
rect 3274 1987 3282 2007
rect 3240 1949 3282 1987
rect 3356 2007 3398 2049
rect 3356 1987 3364 2007
rect 3384 1987 3398 2007
rect 3356 1949 3398 1987
rect 3448 2007 3492 2049
rect 3448 1987 3460 2007
rect 3480 1987 3492 2007
rect 3448 1949 3492 1987
rect 3564 2007 3606 2049
rect 3564 1987 3572 2007
rect 3592 1987 3606 2007
rect 3564 1949 3606 1987
rect 3656 2007 3700 2049
rect 3656 1987 3668 2007
rect 3688 1987 3700 2007
rect 3656 1949 3700 1987
rect 3777 2007 3819 2049
rect 3777 1987 3785 2007
rect 3805 1987 3819 2007
rect 3777 1949 3819 1987
rect 3869 2007 3913 2049
rect 10991 2153 11035 2195
rect 11085 2215 11127 2253
rect 11085 2195 11099 2215
rect 11119 2195 11127 2215
rect 11085 2153 11127 2195
rect 11204 2215 11248 2253
rect 11204 2195 11216 2215
rect 11236 2195 11248 2215
rect 11204 2153 11248 2195
rect 11298 2215 11340 2253
rect 11298 2195 11312 2215
rect 11332 2195 11340 2215
rect 11298 2153 11340 2195
rect 11412 2215 11456 2253
rect 11412 2195 11424 2215
rect 11444 2195 11456 2215
rect 11412 2153 11456 2195
rect 11506 2215 11548 2253
rect 11506 2195 11520 2215
rect 11540 2195 11548 2215
rect 11506 2153 11548 2195
rect 11622 2215 11664 2253
rect 11622 2195 11630 2215
rect 11650 2195 11664 2215
rect 11622 2153 11664 2195
rect 11714 2222 11759 2253
rect 14820 2249 14864 2291
rect 14820 2229 14832 2249
rect 14852 2229 14864 2249
rect 14820 2222 14864 2229
rect 11714 2215 11758 2222
rect 11714 2195 11726 2215
rect 11746 2195 11758 2215
rect 11714 2153 11758 2195
rect 14819 2191 14864 2222
rect 14914 2249 14956 2291
rect 14914 2229 14928 2249
rect 14948 2229 14956 2249
rect 14914 2191 14956 2229
rect 15030 2249 15072 2291
rect 15030 2229 15038 2249
rect 15058 2229 15072 2249
rect 15030 2191 15072 2229
rect 15122 2249 15166 2291
rect 15122 2229 15134 2249
rect 15154 2229 15166 2249
rect 15122 2191 15166 2229
rect 15238 2249 15280 2291
rect 15238 2229 15246 2249
rect 15266 2229 15280 2249
rect 15238 2191 15280 2229
rect 15330 2249 15374 2291
rect 15330 2229 15342 2249
rect 15362 2229 15374 2249
rect 15330 2191 15374 2229
rect 15451 2249 15493 2291
rect 15451 2229 15459 2249
rect 15479 2229 15493 2249
rect 15451 2191 15493 2229
rect 15543 2249 15587 2291
rect 15543 2229 15555 2249
rect 15575 2229 15587 2249
rect 15543 2191 15587 2229
rect 3869 1987 3881 2007
rect 3901 1987 3913 2007
rect 6623 2005 6667 2043
rect 3869 1949 3913 1987
rect 6623 1985 6635 2005
rect 6655 1985 6667 2005
rect 6623 1943 6667 1985
rect 6717 2005 6759 2043
rect 6717 1985 6731 2005
rect 6751 1985 6759 2005
rect 6717 1943 6759 1985
rect 6836 2005 6880 2043
rect 6836 1985 6848 2005
rect 6868 1985 6880 2005
rect 6836 1943 6880 1985
rect 6930 2005 6972 2043
rect 6930 1985 6944 2005
rect 6964 1985 6972 2005
rect 6930 1943 6972 1985
rect 7044 2005 7088 2043
rect 7044 1985 7056 2005
rect 7076 1985 7088 2005
rect 7044 1943 7088 1985
rect 7138 2005 7180 2043
rect 7138 1985 7152 2005
rect 7172 1985 7180 2005
rect 7138 1943 7180 1985
rect 7254 2005 7296 2043
rect 7254 1985 7262 2005
rect 7282 1985 7296 2005
rect 7254 1943 7296 1985
rect 7346 2012 7391 2043
rect 16272 2194 16316 2232
rect 16272 2174 16284 2194
rect 16304 2174 16316 2194
rect 12003 2034 12047 2072
rect 7346 2005 7390 2012
rect 7346 1985 7358 2005
rect 7378 1985 7390 2005
rect 7346 1943 7390 1985
rect 8427 1986 8471 2028
rect 8427 1966 8439 1986
rect 8459 1966 8471 1986
rect 8427 1959 8471 1966
rect 329 1792 373 1830
rect 329 1772 341 1792
rect 361 1772 373 1792
rect 329 1730 373 1772
rect 423 1792 465 1830
rect 423 1772 437 1792
rect 457 1772 465 1792
rect 423 1730 465 1772
rect 542 1792 586 1830
rect 542 1772 554 1792
rect 574 1772 586 1792
rect 542 1730 586 1772
rect 636 1792 678 1830
rect 636 1772 650 1792
rect 670 1772 678 1792
rect 636 1730 678 1772
rect 750 1792 794 1830
rect 750 1772 762 1792
rect 782 1772 794 1792
rect 750 1730 794 1772
rect 844 1792 886 1830
rect 844 1772 858 1792
rect 878 1772 886 1792
rect 844 1730 886 1772
rect 960 1792 1002 1830
rect 960 1772 968 1792
rect 988 1772 1002 1792
rect 960 1730 1002 1772
rect 1052 1799 1097 1830
rect 4158 1826 4202 1868
rect 4158 1806 4170 1826
rect 4190 1806 4202 1826
rect 4158 1799 4202 1806
rect 1052 1792 1096 1799
rect 1052 1772 1064 1792
rect 1084 1772 1096 1792
rect 1052 1730 1096 1772
rect 4157 1768 4202 1799
rect 4252 1826 4294 1868
rect 4252 1806 4266 1826
rect 4286 1806 4294 1826
rect 4252 1768 4294 1806
rect 4368 1826 4410 1868
rect 4368 1806 4376 1826
rect 4396 1806 4410 1826
rect 4368 1768 4410 1806
rect 4460 1826 4504 1868
rect 4460 1806 4472 1826
rect 4492 1806 4504 1826
rect 4460 1768 4504 1806
rect 4576 1826 4618 1868
rect 4576 1806 4584 1826
rect 4604 1806 4618 1826
rect 4576 1768 4618 1806
rect 4668 1826 4712 1868
rect 4668 1806 4680 1826
rect 4700 1806 4712 1826
rect 4668 1768 4712 1806
rect 4789 1826 4831 1868
rect 4789 1806 4797 1826
rect 4817 1806 4831 1826
rect 4789 1768 4831 1806
rect 4881 1826 4925 1868
rect 8426 1928 8471 1959
rect 8521 1986 8563 2028
rect 8521 1966 8535 1986
rect 8555 1966 8563 1986
rect 8521 1928 8563 1966
rect 8637 1986 8679 2028
rect 8637 1966 8645 1986
rect 8665 1966 8679 1986
rect 8637 1928 8679 1966
rect 8729 1986 8773 2028
rect 8729 1966 8741 1986
rect 8761 1966 8773 1986
rect 8729 1928 8773 1966
rect 8845 1986 8887 2028
rect 8845 1966 8853 1986
rect 8873 1966 8887 1986
rect 8845 1928 8887 1966
rect 8937 1986 8981 2028
rect 8937 1966 8949 1986
rect 8969 1966 8981 1986
rect 8937 1928 8981 1966
rect 9058 1986 9100 2028
rect 9058 1966 9066 1986
rect 9086 1966 9100 1986
rect 9058 1928 9100 1966
rect 9150 1986 9194 2028
rect 9150 1966 9162 1986
rect 9182 1966 9194 1986
rect 12003 2014 12015 2034
rect 12035 2014 12047 2034
rect 12003 1972 12047 2014
rect 12097 2034 12139 2072
rect 12097 2014 12111 2034
rect 12131 2014 12139 2034
rect 12097 1972 12139 2014
rect 12216 2034 12260 2072
rect 12216 2014 12228 2034
rect 12248 2014 12260 2034
rect 12216 1972 12260 2014
rect 12310 2034 12352 2072
rect 12310 2014 12324 2034
rect 12344 2014 12352 2034
rect 12310 1972 12352 2014
rect 12424 2034 12468 2072
rect 12424 2014 12436 2034
rect 12456 2014 12468 2034
rect 12424 1972 12468 2014
rect 12518 2034 12560 2072
rect 12518 2014 12532 2034
rect 12552 2014 12560 2034
rect 12518 1972 12560 2014
rect 12634 2034 12676 2072
rect 12634 2014 12642 2034
rect 12662 2014 12676 2034
rect 12634 1972 12676 2014
rect 12726 2041 12771 2072
rect 16272 2132 16316 2174
rect 16366 2194 16408 2232
rect 16366 2174 16380 2194
rect 16400 2174 16408 2194
rect 16366 2132 16408 2174
rect 16485 2194 16529 2232
rect 16485 2174 16497 2194
rect 16517 2174 16529 2194
rect 16485 2132 16529 2174
rect 16579 2194 16621 2232
rect 16579 2174 16593 2194
rect 16613 2174 16621 2194
rect 16579 2132 16621 2174
rect 16693 2194 16737 2232
rect 16693 2174 16705 2194
rect 16725 2174 16737 2194
rect 16693 2132 16737 2174
rect 16787 2194 16829 2232
rect 16787 2174 16801 2194
rect 16821 2174 16829 2194
rect 16787 2132 16829 2174
rect 16903 2194 16945 2232
rect 16903 2174 16911 2194
rect 16931 2174 16945 2194
rect 16903 2132 16945 2174
rect 16995 2201 17040 2232
rect 20101 2228 20145 2270
rect 20101 2208 20113 2228
rect 20133 2208 20145 2228
rect 20101 2201 20145 2208
rect 16995 2194 17039 2201
rect 16995 2174 17007 2194
rect 17027 2174 17039 2194
rect 16995 2132 17039 2174
rect 20100 2170 20145 2201
rect 20195 2228 20237 2270
rect 20195 2208 20209 2228
rect 20229 2208 20237 2228
rect 20195 2170 20237 2208
rect 20311 2228 20353 2270
rect 20311 2208 20319 2228
rect 20339 2208 20353 2228
rect 20311 2170 20353 2208
rect 20403 2228 20447 2270
rect 20403 2208 20415 2228
rect 20435 2208 20447 2228
rect 20403 2170 20447 2208
rect 20519 2228 20561 2270
rect 20519 2208 20527 2228
rect 20547 2208 20561 2228
rect 20519 2170 20561 2208
rect 20611 2228 20655 2270
rect 20611 2208 20623 2228
rect 20643 2208 20655 2228
rect 20611 2170 20655 2208
rect 20732 2228 20774 2270
rect 20732 2208 20740 2228
rect 20760 2208 20774 2228
rect 20732 2170 20774 2208
rect 20824 2228 20868 2270
rect 20824 2208 20836 2228
rect 20856 2208 20868 2228
rect 20824 2170 20868 2208
rect 12726 2034 12770 2041
rect 12726 2014 12738 2034
rect 12758 2014 12770 2034
rect 12726 1972 12770 2014
rect 13807 2015 13851 2057
rect 13807 1995 13819 2015
rect 13839 1995 13851 2015
rect 13807 1988 13851 1995
rect 9150 1928 9194 1966
rect 4881 1806 4893 1826
rect 4913 1806 4925 1826
rect 4881 1768 4925 1806
rect 13806 1957 13851 1988
rect 13901 2015 13943 2057
rect 13901 1995 13915 2015
rect 13935 1995 13943 2015
rect 13901 1957 13943 1995
rect 14017 2015 14059 2057
rect 14017 1995 14025 2015
rect 14045 1995 14059 2015
rect 14017 1957 14059 1995
rect 14109 2015 14153 2057
rect 14109 1995 14121 2015
rect 14141 1995 14153 2015
rect 14109 1957 14153 1995
rect 14225 2015 14267 2057
rect 14225 1995 14233 2015
rect 14253 1995 14267 2015
rect 14225 1957 14267 1995
rect 14317 2015 14361 2057
rect 14317 1995 14329 2015
rect 14349 1995 14361 2015
rect 14317 1957 14361 1995
rect 14438 2015 14480 2057
rect 14438 1995 14446 2015
rect 14466 1995 14480 2015
rect 14438 1957 14480 1995
rect 14530 2015 14574 2057
rect 14530 1995 14542 2015
rect 14562 1995 14574 2015
rect 17284 2013 17328 2051
rect 14530 1957 14574 1995
rect 17284 1993 17296 2013
rect 17316 1993 17328 2013
rect 5610 1771 5654 1809
rect 5610 1751 5622 1771
rect 5642 1751 5654 1771
rect 5610 1709 5654 1751
rect 5704 1771 5746 1809
rect 5704 1751 5718 1771
rect 5738 1751 5746 1771
rect 5704 1709 5746 1751
rect 5823 1771 5867 1809
rect 5823 1751 5835 1771
rect 5855 1751 5867 1771
rect 5823 1709 5867 1751
rect 5917 1771 5959 1809
rect 5917 1751 5931 1771
rect 5951 1751 5959 1771
rect 5917 1709 5959 1751
rect 6031 1771 6075 1809
rect 6031 1751 6043 1771
rect 6063 1751 6075 1771
rect 6031 1709 6075 1751
rect 6125 1771 6167 1809
rect 6125 1751 6139 1771
rect 6159 1751 6167 1771
rect 6125 1709 6167 1751
rect 6241 1771 6283 1809
rect 6241 1751 6249 1771
rect 6269 1751 6283 1771
rect 6241 1709 6283 1751
rect 6333 1778 6378 1809
rect 9439 1805 9483 1847
rect 9439 1785 9451 1805
rect 9471 1785 9483 1805
rect 9439 1778 9483 1785
rect 6333 1771 6377 1778
rect 6333 1751 6345 1771
rect 6365 1751 6377 1771
rect 6333 1709 6377 1751
rect 9438 1747 9483 1778
rect 9533 1805 9575 1847
rect 9533 1785 9547 1805
rect 9567 1785 9575 1805
rect 9533 1747 9575 1785
rect 9649 1805 9691 1847
rect 9649 1785 9657 1805
rect 9677 1785 9691 1805
rect 9649 1747 9691 1785
rect 9741 1805 9785 1847
rect 9741 1785 9753 1805
rect 9773 1785 9785 1805
rect 9741 1747 9785 1785
rect 9857 1805 9899 1847
rect 9857 1785 9865 1805
rect 9885 1785 9899 1805
rect 9857 1747 9899 1785
rect 9949 1805 9993 1847
rect 9949 1785 9961 1805
rect 9981 1785 9993 1805
rect 9949 1747 9993 1785
rect 10070 1805 10112 1847
rect 10070 1785 10078 1805
rect 10098 1785 10112 1805
rect 10070 1747 10112 1785
rect 10162 1805 10206 1847
rect 17284 1951 17328 1993
rect 17378 2013 17420 2051
rect 17378 1993 17392 2013
rect 17412 1993 17420 2013
rect 17378 1951 17420 1993
rect 17497 2013 17541 2051
rect 17497 1993 17509 2013
rect 17529 1993 17541 2013
rect 17497 1951 17541 1993
rect 17591 2013 17633 2051
rect 17591 1993 17605 2013
rect 17625 1993 17633 2013
rect 17591 1951 17633 1993
rect 17705 2013 17749 2051
rect 17705 1993 17717 2013
rect 17737 1993 17749 2013
rect 17705 1951 17749 1993
rect 17799 2013 17841 2051
rect 17799 1993 17813 2013
rect 17833 1993 17841 2013
rect 17799 1951 17841 1993
rect 17915 2013 17957 2051
rect 17915 1993 17923 2013
rect 17943 1993 17957 2013
rect 17915 1951 17957 1993
rect 18007 2020 18052 2051
rect 18007 2013 18051 2020
rect 18007 1993 18019 2013
rect 18039 1993 18051 2013
rect 18007 1951 18051 1993
rect 19088 1994 19132 2036
rect 19088 1974 19100 1994
rect 19120 1974 19132 1994
rect 19088 1967 19132 1974
rect 10162 1785 10174 1805
rect 10194 1785 10206 1805
rect 10162 1747 10206 1785
rect 10990 1800 11034 1838
rect 10990 1780 11002 1800
rect 11022 1780 11034 1800
rect 10990 1738 11034 1780
rect 11084 1800 11126 1838
rect 11084 1780 11098 1800
rect 11118 1780 11126 1800
rect 11084 1738 11126 1780
rect 11203 1800 11247 1838
rect 11203 1780 11215 1800
rect 11235 1780 11247 1800
rect 11203 1738 11247 1780
rect 11297 1800 11339 1838
rect 11297 1780 11311 1800
rect 11331 1780 11339 1800
rect 11297 1738 11339 1780
rect 11411 1800 11455 1838
rect 11411 1780 11423 1800
rect 11443 1780 11455 1800
rect 11411 1738 11455 1780
rect 11505 1800 11547 1838
rect 11505 1780 11519 1800
rect 11539 1780 11547 1800
rect 11505 1738 11547 1780
rect 11621 1800 11663 1838
rect 11621 1780 11629 1800
rect 11649 1780 11663 1800
rect 11621 1738 11663 1780
rect 11713 1807 11758 1838
rect 14819 1834 14863 1876
rect 14819 1814 14831 1834
rect 14851 1814 14863 1834
rect 14819 1807 14863 1814
rect 11713 1800 11757 1807
rect 11713 1780 11725 1800
rect 11745 1780 11757 1800
rect 11713 1738 11757 1780
rect 14818 1776 14863 1807
rect 14913 1834 14955 1876
rect 14913 1814 14927 1834
rect 14947 1814 14955 1834
rect 14913 1776 14955 1814
rect 15029 1834 15071 1876
rect 15029 1814 15037 1834
rect 15057 1814 15071 1834
rect 15029 1776 15071 1814
rect 15121 1834 15165 1876
rect 15121 1814 15133 1834
rect 15153 1814 15165 1834
rect 15121 1776 15165 1814
rect 15237 1834 15279 1876
rect 15237 1814 15245 1834
rect 15265 1814 15279 1834
rect 15237 1776 15279 1814
rect 15329 1834 15373 1876
rect 15329 1814 15341 1834
rect 15361 1814 15373 1834
rect 15329 1776 15373 1814
rect 15450 1834 15492 1876
rect 15450 1814 15458 1834
rect 15478 1814 15492 1834
rect 15450 1776 15492 1814
rect 15542 1834 15586 1876
rect 19087 1936 19132 1967
rect 19182 1994 19224 2036
rect 19182 1974 19196 1994
rect 19216 1974 19224 1994
rect 19182 1936 19224 1974
rect 19298 1994 19340 2036
rect 19298 1974 19306 1994
rect 19326 1974 19340 1994
rect 19298 1936 19340 1974
rect 19390 1994 19434 2036
rect 19390 1974 19402 1994
rect 19422 1974 19434 1994
rect 19390 1936 19434 1974
rect 19506 1994 19548 2036
rect 19506 1974 19514 1994
rect 19534 1974 19548 1994
rect 19506 1936 19548 1974
rect 19598 1994 19642 2036
rect 19598 1974 19610 1994
rect 19630 1974 19642 1994
rect 19598 1936 19642 1974
rect 19719 1994 19761 2036
rect 19719 1974 19727 1994
rect 19747 1974 19761 1994
rect 19719 1936 19761 1974
rect 19811 1994 19855 2036
rect 19811 1974 19823 1994
rect 19843 1974 19855 1994
rect 19811 1936 19855 1974
rect 15542 1814 15554 1834
rect 15574 1814 15586 1834
rect 15542 1776 15586 1814
rect 16271 1779 16315 1817
rect 16271 1759 16283 1779
rect 16303 1759 16315 1779
rect 3096 1587 3140 1629
rect 3096 1567 3108 1587
rect 3128 1567 3140 1587
rect 3096 1560 3140 1567
rect 3095 1529 3140 1560
rect 3190 1587 3232 1629
rect 3190 1567 3204 1587
rect 3224 1567 3232 1587
rect 3190 1529 3232 1567
rect 3306 1587 3348 1629
rect 3306 1567 3314 1587
rect 3334 1567 3348 1587
rect 3306 1529 3348 1567
rect 3398 1587 3442 1629
rect 3398 1567 3410 1587
rect 3430 1567 3442 1587
rect 3398 1529 3442 1567
rect 3514 1587 3556 1629
rect 3514 1567 3522 1587
rect 3542 1567 3556 1587
rect 3514 1529 3556 1567
rect 3606 1587 3650 1629
rect 3606 1567 3618 1587
rect 3638 1567 3650 1587
rect 3606 1529 3650 1567
rect 3727 1587 3769 1629
rect 3727 1567 3735 1587
rect 3755 1567 3769 1587
rect 3727 1529 3769 1567
rect 3819 1587 3863 1629
rect 3819 1567 3831 1587
rect 3851 1567 3863 1587
rect 3819 1529 3863 1567
rect 8377 1566 8421 1608
rect 8377 1546 8389 1566
rect 8409 1546 8421 1566
rect 8377 1539 8421 1546
rect 8376 1508 8421 1539
rect 8471 1566 8513 1608
rect 8471 1546 8485 1566
rect 8505 1546 8513 1566
rect 8471 1508 8513 1546
rect 8587 1566 8629 1608
rect 8587 1546 8595 1566
rect 8615 1546 8629 1566
rect 8587 1508 8629 1546
rect 8679 1566 8723 1608
rect 8679 1546 8691 1566
rect 8711 1546 8723 1566
rect 8679 1508 8723 1546
rect 8795 1566 8837 1608
rect 8795 1546 8803 1566
rect 8823 1546 8837 1566
rect 8795 1508 8837 1546
rect 8887 1566 8931 1608
rect 8887 1546 8899 1566
rect 8919 1546 8931 1566
rect 8887 1508 8931 1546
rect 9008 1566 9050 1608
rect 9008 1546 9016 1566
rect 9036 1546 9050 1566
rect 9008 1508 9050 1546
rect 9100 1566 9144 1608
rect 16271 1717 16315 1759
rect 16365 1779 16407 1817
rect 16365 1759 16379 1779
rect 16399 1759 16407 1779
rect 16365 1717 16407 1759
rect 16484 1779 16528 1817
rect 16484 1759 16496 1779
rect 16516 1759 16528 1779
rect 16484 1717 16528 1759
rect 16578 1779 16620 1817
rect 16578 1759 16592 1779
rect 16612 1759 16620 1779
rect 16578 1717 16620 1759
rect 16692 1779 16736 1817
rect 16692 1759 16704 1779
rect 16724 1759 16736 1779
rect 16692 1717 16736 1759
rect 16786 1779 16828 1817
rect 16786 1759 16800 1779
rect 16820 1759 16828 1779
rect 16786 1717 16828 1759
rect 16902 1779 16944 1817
rect 16902 1759 16910 1779
rect 16930 1759 16944 1779
rect 16902 1717 16944 1759
rect 16994 1786 17039 1817
rect 20100 1813 20144 1855
rect 20100 1793 20112 1813
rect 20132 1793 20144 1813
rect 20100 1786 20144 1793
rect 16994 1779 17038 1786
rect 16994 1759 17006 1779
rect 17026 1759 17038 1779
rect 16994 1717 17038 1759
rect 20099 1755 20144 1786
rect 20194 1813 20236 1855
rect 20194 1793 20208 1813
rect 20228 1793 20236 1813
rect 20194 1755 20236 1793
rect 20310 1813 20352 1855
rect 20310 1793 20318 1813
rect 20338 1793 20352 1813
rect 20310 1755 20352 1793
rect 20402 1813 20446 1855
rect 20402 1793 20414 1813
rect 20434 1793 20446 1813
rect 20402 1755 20446 1793
rect 20518 1813 20560 1855
rect 20518 1793 20526 1813
rect 20546 1793 20560 1813
rect 20518 1755 20560 1793
rect 20610 1813 20654 1855
rect 20610 1793 20622 1813
rect 20642 1793 20654 1813
rect 20610 1755 20654 1793
rect 20731 1813 20773 1855
rect 20731 1793 20739 1813
rect 20759 1793 20773 1813
rect 20731 1755 20773 1793
rect 20823 1813 20867 1855
rect 20823 1793 20835 1813
rect 20855 1793 20867 1813
rect 20823 1755 20867 1793
rect 9100 1546 9112 1566
rect 9132 1546 9144 1566
rect 9100 1508 9144 1546
rect 13757 1595 13801 1637
rect 13757 1575 13769 1595
rect 13789 1575 13801 1595
rect 13757 1568 13801 1575
rect 13756 1537 13801 1568
rect 13851 1595 13893 1637
rect 13851 1575 13865 1595
rect 13885 1575 13893 1595
rect 13851 1537 13893 1575
rect 13967 1595 14009 1637
rect 13967 1575 13975 1595
rect 13995 1575 14009 1595
rect 13967 1537 14009 1575
rect 14059 1595 14103 1637
rect 14059 1575 14071 1595
rect 14091 1575 14103 1595
rect 14059 1537 14103 1575
rect 14175 1595 14217 1637
rect 14175 1575 14183 1595
rect 14203 1575 14217 1595
rect 14175 1537 14217 1575
rect 14267 1595 14311 1637
rect 14267 1575 14279 1595
rect 14299 1575 14311 1595
rect 14267 1537 14311 1575
rect 14388 1595 14430 1637
rect 14388 1575 14396 1595
rect 14416 1575 14430 1595
rect 14388 1537 14430 1575
rect 14480 1595 14524 1637
rect 14480 1575 14492 1595
rect 14512 1575 14524 1595
rect 14480 1537 14524 1575
rect 19038 1574 19082 1616
rect 19038 1554 19050 1574
rect 19070 1554 19082 1574
rect 19038 1547 19082 1554
rect 19037 1516 19082 1547
rect 19132 1574 19174 1616
rect 19132 1554 19146 1574
rect 19166 1554 19174 1574
rect 19132 1516 19174 1554
rect 19248 1574 19290 1616
rect 19248 1554 19256 1574
rect 19276 1554 19290 1574
rect 19248 1516 19290 1554
rect 19340 1574 19384 1616
rect 19340 1554 19352 1574
rect 19372 1554 19384 1574
rect 19340 1516 19384 1554
rect 19456 1574 19498 1616
rect 19456 1554 19464 1574
rect 19484 1554 19498 1574
rect 19456 1516 19498 1554
rect 19548 1574 19592 1616
rect 19548 1554 19560 1574
rect 19580 1554 19592 1574
rect 19548 1516 19592 1554
rect 19669 1574 19711 1616
rect 19669 1554 19677 1574
rect 19697 1554 19711 1574
rect 19669 1516 19711 1554
rect 19761 1574 19805 1616
rect 19761 1554 19773 1574
rect 19793 1554 19805 1574
rect 19761 1516 19805 1554
rect 1397 1465 1441 1503
rect 1397 1445 1409 1465
rect 1429 1445 1441 1465
rect 1397 1403 1441 1445
rect 1491 1465 1533 1503
rect 1491 1445 1505 1465
rect 1525 1445 1533 1465
rect 1491 1403 1533 1445
rect 1610 1465 1654 1503
rect 1610 1445 1622 1465
rect 1642 1445 1654 1465
rect 1610 1403 1654 1445
rect 1704 1465 1746 1503
rect 1704 1445 1718 1465
rect 1738 1445 1746 1465
rect 1704 1403 1746 1445
rect 1818 1465 1862 1503
rect 1818 1445 1830 1465
rect 1850 1445 1862 1465
rect 1818 1403 1862 1445
rect 1912 1465 1954 1503
rect 1912 1445 1926 1465
rect 1946 1445 1954 1465
rect 1912 1403 1954 1445
rect 2028 1465 2070 1503
rect 2028 1445 2036 1465
rect 2056 1445 2070 1465
rect 2028 1403 2070 1445
rect 2120 1472 2165 1503
rect 2120 1465 2164 1472
rect 2120 1445 2132 1465
rect 2152 1445 2164 1465
rect 2120 1403 2164 1445
rect 6678 1444 6722 1482
rect 6678 1424 6690 1444
rect 6710 1424 6722 1444
rect 6678 1382 6722 1424
rect 6772 1444 6814 1482
rect 6772 1424 6786 1444
rect 6806 1424 6814 1444
rect 6772 1382 6814 1424
rect 6891 1444 6935 1482
rect 6891 1424 6903 1444
rect 6923 1424 6935 1444
rect 6891 1382 6935 1424
rect 6985 1444 7027 1482
rect 6985 1424 6999 1444
rect 7019 1424 7027 1444
rect 6985 1382 7027 1424
rect 7099 1444 7143 1482
rect 7099 1424 7111 1444
rect 7131 1424 7143 1444
rect 7099 1382 7143 1424
rect 7193 1444 7235 1482
rect 7193 1424 7207 1444
rect 7227 1424 7235 1444
rect 7193 1382 7235 1424
rect 7309 1444 7351 1482
rect 7309 1424 7317 1444
rect 7337 1424 7351 1444
rect 7309 1382 7351 1424
rect 7401 1451 7446 1482
rect 7401 1444 7445 1451
rect 7401 1424 7413 1444
rect 7433 1424 7445 1444
rect 7401 1382 7445 1424
rect 12058 1473 12102 1511
rect 12058 1453 12070 1473
rect 12090 1453 12102 1473
rect 335 1226 379 1264
rect 335 1206 347 1226
rect 367 1206 379 1226
rect 335 1164 379 1206
rect 429 1226 471 1264
rect 429 1206 443 1226
rect 463 1206 471 1226
rect 429 1164 471 1206
rect 548 1226 592 1264
rect 548 1206 560 1226
rect 580 1206 592 1226
rect 548 1164 592 1206
rect 642 1226 684 1264
rect 642 1206 656 1226
rect 676 1206 684 1226
rect 642 1164 684 1206
rect 756 1226 800 1264
rect 756 1206 768 1226
rect 788 1206 800 1226
rect 756 1164 800 1206
rect 850 1226 892 1264
rect 850 1206 864 1226
rect 884 1206 892 1226
rect 850 1164 892 1206
rect 966 1226 1008 1264
rect 966 1206 974 1226
rect 994 1206 1008 1226
rect 966 1164 1008 1206
rect 1058 1233 1103 1264
rect 4164 1260 4208 1302
rect 4164 1240 4176 1260
rect 4196 1240 4208 1260
rect 4164 1233 4208 1240
rect 1058 1226 1102 1233
rect 1058 1206 1070 1226
rect 1090 1206 1102 1226
rect 1058 1164 1102 1206
rect 4163 1202 4208 1233
rect 4258 1260 4300 1302
rect 4258 1240 4272 1260
rect 4292 1240 4300 1260
rect 4258 1202 4300 1240
rect 4374 1260 4416 1302
rect 4374 1240 4382 1260
rect 4402 1240 4416 1260
rect 4374 1202 4416 1240
rect 4466 1260 4510 1302
rect 4466 1240 4478 1260
rect 4498 1240 4510 1260
rect 4466 1202 4510 1240
rect 4582 1260 4624 1302
rect 4582 1240 4590 1260
rect 4610 1240 4624 1260
rect 4582 1202 4624 1240
rect 4674 1260 4718 1302
rect 4674 1240 4686 1260
rect 4706 1240 4718 1260
rect 4674 1202 4718 1240
rect 4795 1260 4837 1302
rect 4795 1240 4803 1260
rect 4823 1240 4837 1260
rect 4795 1202 4837 1240
rect 4887 1260 4931 1302
rect 12058 1411 12102 1453
rect 12152 1473 12194 1511
rect 12152 1453 12166 1473
rect 12186 1453 12194 1473
rect 12152 1411 12194 1453
rect 12271 1473 12315 1511
rect 12271 1453 12283 1473
rect 12303 1453 12315 1473
rect 12271 1411 12315 1453
rect 12365 1473 12407 1511
rect 12365 1453 12379 1473
rect 12399 1453 12407 1473
rect 12365 1411 12407 1453
rect 12479 1473 12523 1511
rect 12479 1453 12491 1473
rect 12511 1453 12523 1473
rect 12479 1411 12523 1453
rect 12573 1473 12615 1511
rect 12573 1453 12587 1473
rect 12607 1453 12615 1473
rect 12573 1411 12615 1453
rect 12689 1473 12731 1511
rect 12689 1453 12697 1473
rect 12717 1453 12731 1473
rect 12689 1411 12731 1453
rect 12781 1480 12826 1511
rect 12781 1473 12825 1480
rect 12781 1453 12793 1473
rect 12813 1453 12825 1473
rect 12781 1411 12825 1453
rect 17339 1452 17383 1490
rect 17339 1432 17351 1452
rect 17371 1432 17383 1452
rect 17339 1390 17383 1432
rect 17433 1452 17475 1490
rect 17433 1432 17447 1452
rect 17467 1432 17475 1452
rect 17433 1390 17475 1432
rect 17552 1452 17596 1490
rect 17552 1432 17564 1452
rect 17584 1432 17596 1452
rect 17552 1390 17596 1432
rect 17646 1452 17688 1490
rect 17646 1432 17660 1452
rect 17680 1432 17688 1452
rect 17646 1390 17688 1432
rect 17760 1452 17804 1490
rect 17760 1432 17772 1452
rect 17792 1432 17804 1452
rect 17760 1390 17804 1432
rect 17854 1452 17896 1490
rect 17854 1432 17868 1452
rect 17888 1432 17896 1452
rect 17854 1390 17896 1432
rect 17970 1452 18012 1490
rect 17970 1432 17978 1452
rect 17998 1432 18012 1452
rect 17970 1390 18012 1432
rect 18062 1459 18107 1490
rect 18062 1452 18106 1459
rect 18062 1432 18074 1452
rect 18094 1432 18106 1452
rect 18062 1390 18106 1432
rect 4887 1240 4899 1260
rect 4919 1240 4931 1260
rect 4887 1202 4931 1240
rect 5616 1205 5660 1243
rect 5616 1185 5628 1205
rect 5648 1185 5660 1205
rect 1347 1045 1391 1083
rect 1347 1025 1359 1045
rect 1379 1025 1391 1045
rect 1347 983 1391 1025
rect 1441 1045 1483 1083
rect 1441 1025 1455 1045
rect 1475 1025 1483 1045
rect 1441 983 1483 1025
rect 1560 1045 1604 1083
rect 1560 1025 1572 1045
rect 1592 1025 1604 1045
rect 1560 983 1604 1025
rect 1654 1045 1696 1083
rect 1654 1025 1668 1045
rect 1688 1025 1696 1045
rect 1654 983 1696 1025
rect 1768 1045 1812 1083
rect 1768 1025 1780 1045
rect 1800 1025 1812 1045
rect 1768 983 1812 1025
rect 1862 1045 1904 1083
rect 1862 1025 1876 1045
rect 1896 1025 1904 1045
rect 1862 983 1904 1025
rect 1978 1045 2020 1083
rect 1978 1025 1986 1045
rect 2006 1025 2020 1045
rect 1978 983 2020 1025
rect 2070 1052 2115 1083
rect 5616 1143 5660 1185
rect 5710 1205 5752 1243
rect 5710 1185 5724 1205
rect 5744 1185 5752 1205
rect 5710 1143 5752 1185
rect 5829 1205 5873 1243
rect 5829 1185 5841 1205
rect 5861 1185 5873 1205
rect 5829 1143 5873 1185
rect 5923 1205 5965 1243
rect 5923 1185 5937 1205
rect 5957 1185 5965 1205
rect 5923 1143 5965 1185
rect 6037 1205 6081 1243
rect 6037 1185 6049 1205
rect 6069 1185 6081 1205
rect 6037 1143 6081 1185
rect 6131 1205 6173 1243
rect 6131 1185 6145 1205
rect 6165 1185 6173 1205
rect 6131 1143 6173 1185
rect 6247 1205 6289 1243
rect 6247 1185 6255 1205
rect 6275 1185 6289 1205
rect 6247 1143 6289 1185
rect 6339 1212 6384 1243
rect 9445 1239 9489 1281
rect 9445 1219 9457 1239
rect 9477 1219 9489 1239
rect 9445 1212 9489 1219
rect 6339 1205 6383 1212
rect 6339 1185 6351 1205
rect 6371 1185 6383 1205
rect 6339 1143 6383 1185
rect 9444 1181 9489 1212
rect 9539 1239 9581 1281
rect 9539 1219 9553 1239
rect 9573 1219 9581 1239
rect 9539 1181 9581 1219
rect 9655 1239 9697 1281
rect 9655 1219 9663 1239
rect 9683 1219 9697 1239
rect 9655 1181 9697 1219
rect 9747 1239 9791 1281
rect 9747 1219 9759 1239
rect 9779 1219 9791 1239
rect 9747 1181 9791 1219
rect 9863 1239 9905 1281
rect 9863 1219 9871 1239
rect 9891 1219 9905 1239
rect 9863 1181 9905 1219
rect 9955 1239 9999 1281
rect 9955 1219 9967 1239
rect 9987 1219 9999 1239
rect 9955 1181 9999 1219
rect 10076 1239 10118 1281
rect 10076 1219 10084 1239
rect 10104 1219 10118 1239
rect 10076 1181 10118 1219
rect 10168 1239 10212 1281
rect 10168 1219 10180 1239
rect 10200 1219 10212 1239
rect 10168 1181 10212 1219
rect 10996 1234 11040 1272
rect 10996 1214 11008 1234
rect 11028 1214 11040 1234
rect 2070 1045 2114 1052
rect 2070 1025 2082 1045
rect 2102 1025 2114 1045
rect 2070 983 2114 1025
rect 3151 1026 3195 1068
rect 3151 1006 3163 1026
rect 3183 1006 3195 1026
rect 3151 999 3195 1006
rect 3150 968 3195 999
rect 3245 1026 3287 1068
rect 3245 1006 3259 1026
rect 3279 1006 3287 1026
rect 3245 968 3287 1006
rect 3361 1026 3403 1068
rect 3361 1006 3369 1026
rect 3389 1006 3403 1026
rect 3361 968 3403 1006
rect 3453 1026 3497 1068
rect 3453 1006 3465 1026
rect 3485 1006 3497 1026
rect 3453 968 3497 1006
rect 3569 1026 3611 1068
rect 3569 1006 3577 1026
rect 3597 1006 3611 1026
rect 3569 968 3611 1006
rect 3661 1026 3705 1068
rect 3661 1006 3673 1026
rect 3693 1006 3705 1026
rect 3661 968 3705 1006
rect 3782 1026 3824 1068
rect 3782 1006 3790 1026
rect 3810 1006 3824 1026
rect 3782 968 3824 1006
rect 3874 1026 3918 1068
rect 10996 1172 11040 1214
rect 11090 1234 11132 1272
rect 11090 1214 11104 1234
rect 11124 1214 11132 1234
rect 11090 1172 11132 1214
rect 11209 1234 11253 1272
rect 11209 1214 11221 1234
rect 11241 1214 11253 1234
rect 11209 1172 11253 1214
rect 11303 1234 11345 1272
rect 11303 1214 11317 1234
rect 11337 1214 11345 1234
rect 11303 1172 11345 1214
rect 11417 1234 11461 1272
rect 11417 1214 11429 1234
rect 11449 1214 11461 1234
rect 11417 1172 11461 1214
rect 11511 1234 11553 1272
rect 11511 1214 11525 1234
rect 11545 1214 11553 1234
rect 11511 1172 11553 1214
rect 11627 1234 11669 1272
rect 11627 1214 11635 1234
rect 11655 1214 11669 1234
rect 11627 1172 11669 1214
rect 11719 1241 11764 1272
rect 14825 1268 14869 1310
rect 14825 1248 14837 1268
rect 14857 1248 14869 1268
rect 14825 1241 14869 1248
rect 11719 1234 11763 1241
rect 11719 1214 11731 1234
rect 11751 1214 11763 1234
rect 11719 1172 11763 1214
rect 14824 1210 14869 1241
rect 14919 1268 14961 1310
rect 14919 1248 14933 1268
rect 14953 1248 14961 1268
rect 14919 1210 14961 1248
rect 15035 1268 15077 1310
rect 15035 1248 15043 1268
rect 15063 1248 15077 1268
rect 15035 1210 15077 1248
rect 15127 1268 15171 1310
rect 15127 1248 15139 1268
rect 15159 1248 15171 1268
rect 15127 1210 15171 1248
rect 15243 1268 15285 1310
rect 15243 1248 15251 1268
rect 15271 1248 15285 1268
rect 15243 1210 15285 1248
rect 15335 1268 15379 1310
rect 15335 1248 15347 1268
rect 15367 1248 15379 1268
rect 15335 1210 15379 1248
rect 15456 1268 15498 1310
rect 15456 1248 15464 1268
rect 15484 1248 15498 1268
rect 15456 1210 15498 1248
rect 15548 1268 15592 1310
rect 15548 1248 15560 1268
rect 15580 1248 15592 1268
rect 15548 1210 15592 1248
rect 3874 1006 3886 1026
rect 3906 1006 3918 1026
rect 6628 1024 6672 1062
rect 3874 968 3918 1006
rect 6628 1004 6640 1024
rect 6660 1004 6672 1024
rect 6628 962 6672 1004
rect 6722 1024 6764 1062
rect 6722 1004 6736 1024
rect 6756 1004 6764 1024
rect 6722 962 6764 1004
rect 6841 1024 6885 1062
rect 6841 1004 6853 1024
rect 6873 1004 6885 1024
rect 6841 962 6885 1004
rect 6935 1024 6977 1062
rect 6935 1004 6949 1024
rect 6969 1004 6977 1024
rect 6935 962 6977 1004
rect 7049 1024 7093 1062
rect 7049 1004 7061 1024
rect 7081 1004 7093 1024
rect 7049 962 7093 1004
rect 7143 1024 7185 1062
rect 7143 1004 7157 1024
rect 7177 1004 7185 1024
rect 7143 962 7185 1004
rect 7259 1024 7301 1062
rect 7259 1004 7267 1024
rect 7287 1004 7301 1024
rect 7259 962 7301 1004
rect 7351 1031 7396 1062
rect 16277 1213 16321 1251
rect 16277 1193 16289 1213
rect 16309 1193 16321 1213
rect 12008 1053 12052 1091
rect 7351 1024 7395 1031
rect 7351 1004 7363 1024
rect 7383 1004 7395 1024
rect 7351 962 7395 1004
rect 8432 1005 8476 1047
rect 8432 985 8444 1005
rect 8464 985 8476 1005
rect 8432 978 8476 985
rect 334 811 378 849
rect 334 791 346 811
rect 366 791 378 811
rect 334 749 378 791
rect 428 811 470 849
rect 428 791 442 811
rect 462 791 470 811
rect 428 749 470 791
rect 547 811 591 849
rect 547 791 559 811
rect 579 791 591 811
rect 547 749 591 791
rect 641 811 683 849
rect 641 791 655 811
rect 675 791 683 811
rect 641 749 683 791
rect 755 811 799 849
rect 755 791 767 811
rect 787 791 799 811
rect 755 749 799 791
rect 849 811 891 849
rect 849 791 863 811
rect 883 791 891 811
rect 849 749 891 791
rect 965 811 1007 849
rect 965 791 973 811
rect 993 791 1007 811
rect 965 749 1007 791
rect 1057 818 1102 849
rect 4163 845 4207 887
rect 4163 825 4175 845
rect 4195 825 4207 845
rect 4163 818 4207 825
rect 1057 811 1101 818
rect 1057 791 1069 811
rect 1089 791 1101 811
rect 1057 749 1101 791
rect 4162 787 4207 818
rect 4257 845 4299 887
rect 4257 825 4271 845
rect 4291 825 4299 845
rect 4257 787 4299 825
rect 4373 845 4415 887
rect 4373 825 4381 845
rect 4401 825 4415 845
rect 4373 787 4415 825
rect 4465 845 4509 887
rect 4465 825 4477 845
rect 4497 825 4509 845
rect 4465 787 4509 825
rect 4581 845 4623 887
rect 4581 825 4589 845
rect 4609 825 4623 845
rect 4581 787 4623 825
rect 4673 845 4717 887
rect 4673 825 4685 845
rect 4705 825 4717 845
rect 4673 787 4717 825
rect 4794 845 4836 887
rect 4794 825 4802 845
rect 4822 825 4836 845
rect 4794 787 4836 825
rect 4886 845 4930 887
rect 8431 947 8476 978
rect 8526 1005 8568 1047
rect 8526 985 8540 1005
rect 8560 985 8568 1005
rect 8526 947 8568 985
rect 8642 1005 8684 1047
rect 8642 985 8650 1005
rect 8670 985 8684 1005
rect 8642 947 8684 985
rect 8734 1005 8778 1047
rect 8734 985 8746 1005
rect 8766 985 8778 1005
rect 8734 947 8778 985
rect 8850 1005 8892 1047
rect 8850 985 8858 1005
rect 8878 985 8892 1005
rect 8850 947 8892 985
rect 8942 1005 8986 1047
rect 8942 985 8954 1005
rect 8974 985 8986 1005
rect 8942 947 8986 985
rect 9063 1005 9105 1047
rect 9063 985 9071 1005
rect 9091 985 9105 1005
rect 9063 947 9105 985
rect 9155 1005 9199 1047
rect 9155 985 9167 1005
rect 9187 985 9199 1005
rect 12008 1033 12020 1053
rect 12040 1033 12052 1053
rect 12008 991 12052 1033
rect 12102 1053 12144 1091
rect 12102 1033 12116 1053
rect 12136 1033 12144 1053
rect 12102 991 12144 1033
rect 12221 1053 12265 1091
rect 12221 1033 12233 1053
rect 12253 1033 12265 1053
rect 12221 991 12265 1033
rect 12315 1053 12357 1091
rect 12315 1033 12329 1053
rect 12349 1033 12357 1053
rect 12315 991 12357 1033
rect 12429 1053 12473 1091
rect 12429 1033 12441 1053
rect 12461 1033 12473 1053
rect 12429 991 12473 1033
rect 12523 1053 12565 1091
rect 12523 1033 12537 1053
rect 12557 1033 12565 1053
rect 12523 991 12565 1033
rect 12639 1053 12681 1091
rect 12639 1033 12647 1053
rect 12667 1033 12681 1053
rect 12639 991 12681 1033
rect 12731 1060 12776 1091
rect 16277 1151 16321 1193
rect 16371 1213 16413 1251
rect 16371 1193 16385 1213
rect 16405 1193 16413 1213
rect 16371 1151 16413 1193
rect 16490 1213 16534 1251
rect 16490 1193 16502 1213
rect 16522 1193 16534 1213
rect 16490 1151 16534 1193
rect 16584 1213 16626 1251
rect 16584 1193 16598 1213
rect 16618 1193 16626 1213
rect 16584 1151 16626 1193
rect 16698 1213 16742 1251
rect 16698 1193 16710 1213
rect 16730 1193 16742 1213
rect 16698 1151 16742 1193
rect 16792 1213 16834 1251
rect 16792 1193 16806 1213
rect 16826 1193 16834 1213
rect 16792 1151 16834 1193
rect 16908 1213 16950 1251
rect 16908 1193 16916 1213
rect 16936 1193 16950 1213
rect 16908 1151 16950 1193
rect 17000 1220 17045 1251
rect 20106 1247 20150 1289
rect 20106 1227 20118 1247
rect 20138 1227 20150 1247
rect 20106 1220 20150 1227
rect 17000 1213 17044 1220
rect 17000 1193 17012 1213
rect 17032 1193 17044 1213
rect 17000 1151 17044 1193
rect 20105 1189 20150 1220
rect 20200 1247 20242 1289
rect 20200 1227 20214 1247
rect 20234 1227 20242 1247
rect 20200 1189 20242 1227
rect 20316 1247 20358 1289
rect 20316 1227 20324 1247
rect 20344 1227 20358 1247
rect 20316 1189 20358 1227
rect 20408 1247 20452 1289
rect 20408 1227 20420 1247
rect 20440 1227 20452 1247
rect 20408 1189 20452 1227
rect 20524 1247 20566 1289
rect 20524 1227 20532 1247
rect 20552 1227 20566 1247
rect 20524 1189 20566 1227
rect 20616 1247 20660 1289
rect 20616 1227 20628 1247
rect 20648 1227 20660 1247
rect 20616 1189 20660 1227
rect 20737 1247 20779 1289
rect 20737 1227 20745 1247
rect 20765 1227 20779 1247
rect 20737 1189 20779 1227
rect 20829 1247 20873 1289
rect 20829 1227 20841 1247
rect 20861 1227 20873 1247
rect 20829 1189 20873 1227
rect 12731 1053 12775 1060
rect 12731 1033 12743 1053
rect 12763 1033 12775 1053
rect 12731 991 12775 1033
rect 13812 1034 13856 1076
rect 13812 1014 13824 1034
rect 13844 1014 13856 1034
rect 13812 1007 13856 1014
rect 9155 947 9199 985
rect 4886 825 4898 845
rect 4918 825 4930 845
rect 4886 787 4930 825
rect 13811 976 13856 1007
rect 13906 1034 13948 1076
rect 13906 1014 13920 1034
rect 13940 1014 13948 1034
rect 13906 976 13948 1014
rect 14022 1034 14064 1076
rect 14022 1014 14030 1034
rect 14050 1014 14064 1034
rect 14022 976 14064 1014
rect 14114 1034 14158 1076
rect 14114 1014 14126 1034
rect 14146 1014 14158 1034
rect 14114 976 14158 1014
rect 14230 1034 14272 1076
rect 14230 1014 14238 1034
rect 14258 1014 14272 1034
rect 14230 976 14272 1014
rect 14322 1034 14366 1076
rect 14322 1014 14334 1034
rect 14354 1014 14366 1034
rect 14322 976 14366 1014
rect 14443 1034 14485 1076
rect 14443 1014 14451 1034
rect 14471 1014 14485 1034
rect 14443 976 14485 1014
rect 14535 1034 14579 1076
rect 14535 1014 14547 1034
rect 14567 1014 14579 1034
rect 17289 1032 17333 1070
rect 14535 976 14579 1014
rect 17289 1012 17301 1032
rect 17321 1012 17333 1032
rect 5615 790 5659 828
rect 5615 770 5627 790
rect 5647 770 5659 790
rect 5615 728 5659 770
rect 5709 790 5751 828
rect 5709 770 5723 790
rect 5743 770 5751 790
rect 5709 728 5751 770
rect 5828 790 5872 828
rect 5828 770 5840 790
rect 5860 770 5872 790
rect 5828 728 5872 770
rect 5922 790 5964 828
rect 5922 770 5936 790
rect 5956 770 5964 790
rect 5922 728 5964 770
rect 6036 790 6080 828
rect 6036 770 6048 790
rect 6068 770 6080 790
rect 6036 728 6080 770
rect 6130 790 6172 828
rect 6130 770 6144 790
rect 6164 770 6172 790
rect 6130 728 6172 770
rect 6246 790 6288 828
rect 6246 770 6254 790
rect 6274 770 6288 790
rect 6246 728 6288 770
rect 6338 797 6383 828
rect 9444 824 9488 866
rect 9444 804 9456 824
rect 9476 804 9488 824
rect 9444 797 9488 804
rect 6338 790 6382 797
rect 6338 770 6350 790
rect 6370 770 6382 790
rect 6338 728 6382 770
rect 9443 766 9488 797
rect 9538 824 9580 866
rect 9538 804 9552 824
rect 9572 804 9580 824
rect 9538 766 9580 804
rect 9654 824 9696 866
rect 9654 804 9662 824
rect 9682 804 9696 824
rect 9654 766 9696 804
rect 9746 824 9790 866
rect 9746 804 9758 824
rect 9778 804 9790 824
rect 9746 766 9790 804
rect 9862 824 9904 866
rect 9862 804 9870 824
rect 9890 804 9904 824
rect 9862 766 9904 804
rect 9954 824 9998 866
rect 9954 804 9966 824
rect 9986 804 9998 824
rect 9954 766 9998 804
rect 10075 824 10117 866
rect 10075 804 10083 824
rect 10103 804 10117 824
rect 10075 766 10117 804
rect 10167 824 10211 866
rect 17289 970 17333 1012
rect 17383 1032 17425 1070
rect 17383 1012 17397 1032
rect 17417 1012 17425 1032
rect 17383 970 17425 1012
rect 17502 1032 17546 1070
rect 17502 1012 17514 1032
rect 17534 1012 17546 1032
rect 17502 970 17546 1012
rect 17596 1032 17638 1070
rect 17596 1012 17610 1032
rect 17630 1012 17638 1032
rect 17596 970 17638 1012
rect 17710 1032 17754 1070
rect 17710 1012 17722 1032
rect 17742 1012 17754 1032
rect 17710 970 17754 1012
rect 17804 1032 17846 1070
rect 17804 1012 17818 1032
rect 17838 1012 17846 1032
rect 17804 970 17846 1012
rect 17920 1032 17962 1070
rect 17920 1012 17928 1032
rect 17948 1012 17962 1032
rect 17920 970 17962 1012
rect 18012 1039 18057 1070
rect 18012 1032 18056 1039
rect 18012 1012 18024 1032
rect 18044 1012 18056 1032
rect 18012 970 18056 1012
rect 19093 1013 19137 1055
rect 19093 993 19105 1013
rect 19125 993 19137 1013
rect 19093 986 19137 993
rect 10167 804 10179 824
rect 10199 804 10211 824
rect 10167 766 10211 804
rect 10995 819 11039 857
rect 10995 799 11007 819
rect 11027 799 11039 819
rect 10995 757 11039 799
rect 11089 819 11131 857
rect 11089 799 11103 819
rect 11123 799 11131 819
rect 11089 757 11131 799
rect 11208 819 11252 857
rect 11208 799 11220 819
rect 11240 799 11252 819
rect 11208 757 11252 799
rect 11302 819 11344 857
rect 11302 799 11316 819
rect 11336 799 11344 819
rect 11302 757 11344 799
rect 11416 819 11460 857
rect 11416 799 11428 819
rect 11448 799 11460 819
rect 11416 757 11460 799
rect 11510 819 11552 857
rect 11510 799 11524 819
rect 11544 799 11552 819
rect 11510 757 11552 799
rect 11626 819 11668 857
rect 11626 799 11634 819
rect 11654 799 11668 819
rect 11626 757 11668 799
rect 11718 826 11763 857
rect 14824 853 14868 895
rect 14824 833 14836 853
rect 14856 833 14868 853
rect 14824 826 14868 833
rect 11718 819 11762 826
rect 11718 799 11730 819
rect 11750 799 11762 819
rect 11718 757 11762 799
rect 14823 795 14868 826
rect 14918 853 14960 895
rect 14918 833 14932 853
rect 14952 833 14960 853
rect 14918 795 14960 833
rect 15034 853 15076 895
rect 15034 833 15042 853
rect 15062 833 15076 853
rect 15034 795 15076 833
rect 15126 853 15170 895
rect 15126 833 15138 853
rect 15158 833 15170 853
rect 15126 795 15170 833
rect 15242 853 15284 895
rect 15242 833 15250 853
rect 15270 833 15284 853
rect 15242 795 15284 833
rect 15334 853 15378 895
rect 15334 833 15346 853
rect 15366 833 15378 853
rect 15334 795 15378 833
rect 15455 853 15497 895
rect 15455 833 15463 853
rect 15483 833 15497 853
rect 15455 795 15497 833
rect 15547 853 15591 895
rect 19092 955 19137 986
rect 19187 1013 19229 1055
rect 19187 993 19201 1013
rect 19221 993 19229 1013
rect 19187 955 19229 993
rect 19303 1013 19345 1055
rect 19303 993 19311 1013
rect 19331 993 19345 1013
rect 19303 955 19345 993
rect 19395 1013 19439 1055
rect 19395 993 19407 1013
rect 19427 993 19439 1013
rect 19395 955 19439 993
rect 19511 1013 19553 1055
rect 19511 993 19519 1013
rect 19539 993 19553 1013
rect 19511 955 19553 993
rect 19603 1013 19647 1055
rect 19603 993 19615 1013
rect 19635 993 19647 1013
rect 19603 955 19647 993
rect 19724 1013 19766 1055
rect 19724 993 19732 1013
rect 19752 993 19766 1013
rect 19724 955 19766 993
rect 19816 1013 19860 1055
rect 19816 993 19828 1013
rect 19848 993 19860 1013
rect 19816 955 19860 993
rect 15547 833 15559 853
rect 15579 833 15591 853
rect 15547 795 15591 833
rect 16276 798 16320 836
rect 16276 778 16288 798
rect 16308 778 16320 798
rect 16276 736 16320 778
rect 16370 798 16412 836
rect 16370 778 16384 798
rect 16404 778 16412 798
rect 16370 736 16412 778
rect 16489 798 16533 836
rect 16489 778 16501 798
rect 16521 778 16533 798
rect 16489 736 16533 778
rect 16583 798 16625 836
rect 16583 778 16597 798
rect 16617 778 16625 798
rect 16583 736 16625 778
rect 16697 798 16741 836
rect 16697 778 16709 798
rect 16729 778 16741 798
rect 16697 736 16741 778
rect 16791 798 16833 836
rect 16791 778 16805 798
rect 16825 778 16833 798
rect 16791 736 16833 778
rect 16907 798 16949 836
rect 16907 778 16915 798
rect 16935 778 16949 798
rect 16907 736 16949 778
rect 16999 805 17044 836
rect 20105 832 20149 874
rect 20105 812 20117 832
rect 20137 812 20149 832
rect 20105 805 20149 812
rect 16999 798 17043 805
rect 16999 778 17011 798
rect 17031 778 17043 798
rect 16999 736 17043 778
rect 20104 774 20149 805
rect 20199 832 20241 874
rect 20199 812 20213 832
rect 20233 812 20241 832
rect 20199 774 20241 812
rect 20315 832 20357 874
rect 20315 812 20323 832
rect 20343 812 20357 832
rect 20315 774 20357 812
rect 20407 832 20451 874
rect 20407 812 20419 832
rect 20439 812 20451 832
rect 20407 774 20451 812
rect 20523 832 20565 874
rect 20523 812 20531 832
rect 20551 812 20565 832
rect 20523 774 20565 812
rect 20615 832 20659 874
rect 20615 812 20627 832
rect 20647 812 20659 832
rect 20615 774 20659 812
rect 20736 832 20778 874
rect 20736 812 20744 832
rect 20764 812 20778 832
rect 20736 774 20778 812
rect 20828 832 20872 874
rect 20828 812 20840 832
rect 20860 812 20872 832
rect 20828 774 20872 812
rect 1737 330 1781 368
rect 1737 310 1749 330
rect 1769 310 1781 330
rect 1737 268 1781 310
rect 1831 330 1873 368
rect 1831 310 1845 330
rect 1865 310 1873 330
rect 1831 268 1873 310
rect 1950 330 1994 368
rect 1950 310 1962 330
rect 1982 310 1994 330
rect 1950 268 1994 310
rect 2044 330 2086 368
rect 2044 310 2058 330
rect 2078 310 2086 330
rect 2044 268 2086 310
rect 2158 330 2202 368
rect 2158 310 2170 330
rect 2190 310 2202 330
rect 2158 268 2202 310
rect 2252 330 2294 368
rect 2252 310 2266 330
rect 2286 310 2294 330
rect 2252 268 2294 310
rect 2368 330 2410 368
rect 2368 310 2376 330
rect 2396 310 2410 330
rect 2368 268 2410 310
rect 2460 337 2505 368
rect 2460 330 2504 337
rect 2460 310 2472 330
rect 2492 310 2504 330
rect 2460 268 2504 310
rect 7018 309 7062 347
rect 7018 289 7030 309
rect 7050 289 7062 309
rect 4827 242 4871 280
rect 4827 222 4839 242
rect 4859 222 4871 242
rect 4827 180 4871 222
rect 4921 242 4963 280
rect 4921 222 4935 242
rect 4955 222 4963 242
rect 4921 180 4963 222
rect 5040 242 5084 280
rect 5040 222 5052 242
rect 5072 222 5084 242
rect 5040 180 5084 222
rect 5134 242 5176 280
rect 5134 222 5148 242
rect 5168 222 5176 242
rect 5134 180 5176 222
rect 5248 242 5292 280
rect 5248 222 5260 242
rect 5280 222 5292 242
rect 5248 180 5292 222
rect 5342 242 5384 280
rect 5342 222 5356 242
rect 5376 222 5384 242
rect 5342 180 5384 222
rect 5458 242 5500 280
rect 5458 222 5466 242
rect 5486 222 5500 242
rect 5458 180 5500 222
rect 5550 249 5595 280
rect 5550 242 5594 249
rect 7018 247 7062 289
rect 7112 309 7154 347
rect 7112 289 7126 309
rect 7146 289 7154 309
rect 7112 247 7154 289
rect 7231 309 7275 347
rect 7231 289 7243 309
rect 7263 289 7275 309
rect 7231 247 7275 289
rect 7325 309 7367 347
rect 7325 289 7339 309
rect 7359 289 7367 309
rect 7325 247 7367 289
rect 7439 309 7483 347
rect 7439 289 7451 309
rect 7471 289 7483 309
rect 7439 247 7483 289
rect 7533 309 7575 347
rect 7533 289 7547 309
rect 7567 289 7575 309
rect 7533 247 7575 289
rect 7649 309 7691 347
rect 7649 289 7657 309
rect 7677 289 7691 309
rect 7649 247 7691 289
rect 7741 316 7786 347
rect 12398 338 12442 376
rect 12398 318 12410 338
rect 12430 318 12442 338
rect 7741 309 7785 316
rect 7741 289 7753 309
rect 7773 289 7785 309
rect 7741 247 7785 289
rect 12398 276 12442 318
rect 12492 338 12534 376
rect 12492 318 12506 338
rect 12526 318 12534 338
rect 12492 276 12534 318
rect 12611 338 12655 376
rect 12611 318 12623 338
rect 12643 318 12655 338
rect 12611 276 12655 318
rect 12705 338 12747 376
rect 12705 318 12719 338
rect 12739 318 12747 338
rect 12705 276 12747 318
rect 12819 338 12863 376
rect 12819 318 12831 338
rect 12851 318 12863 338
rect 12819 276 12863 318
rect 12913 338 12955 376
rect 12913 318 12927 338
rect 12947 318 12955 338
rect 12913 276 12955 318
rect 13029 338 13071 376
rect 13029 318 13037 338
rect 13057 318 13071 338
rect 13029 276 13071 318
rect 13121 345 13166 376
rect 13121 338 13165 345
rect 13121 318 13133 338
rect 13153 318 13165 338
rect 13121 276 13165 318
rect 17679 317 17723 355
rect 17679 297 17691 317
rect 17711 297 17723 317
rect 5550 222 5562 242
rect 5582 222 5594 242
rect 5550 180 5594 222
rect 10088 235 10132 273
rect 10088 215 10100 235
rect 10120 215 10132 235
rect 10088 173 10132 215
rect 10182 235 10224 273
rect 10182 215 10196 235
rect 10216 215 10224 235
rect 10182 173 10224 215
rect 10301 235 10345 273
rect 10301 215 10313 235
rect 10333 215 10345 235
rect 10301 173 10345 215
rect 10395 235 10437 273
rect 10395 215 10409 235
rect 10429 215 10437 235
rect 10395 173 10437 215
rect 10509 235 10553 273
rect 10509 215 10521 235
rect 10541 215 10553 235
rect 10509 173 10553 215
rect 10603 235 10645 273
rect 10603 215 10617 235
rect 10637 215 10645 235
rect 10603 173 10645 215
rect 10719 235 10761 273
rect 10719 215 10727 235
rect 10747 215 10761 235
rect 10719 173 10761 215
rect 10811 242 10856 273
rect 10811 235 10855 242
rect 10811 215 10823 235
rect 10843 215 10855 235
rect 10811 173 10855 215
rect 15488 250 15532 288
rect 15488 230 15500 250
rect 15520 230 15532 250
rect 15488 188 15532 230
rect 15582 250 15624 288
rect 15582 230 15596 250
rect 15616 230 15624 250
rect 15582 188 15624 230
rect 15701 250 15745 288
rect 15701 230 15713 250
rect 15733 230 15745 250
rect 15701 188 15745 230
rect 15795 250 15837 288
rect 15795 230 15809 250
rect 15829 230 15837 250
rect 15795 188 15837 230
rect 15909 250 15953 288
rect 15909 230 15921 250
rect 15941 230 15953 250
rect 15909 188 15953 230
rect 16003 250 16045 288
rect 16003 230 16017 250
rect 16037 230 16045 250
rect 16003 188 16045 230
rect 16119 250 16161 288
rect 16119 230 16127 250
rect 16147 230 16161 250
rect 16119 188 16161 230
rect 16211 257 16256 288
rect 16211 250 16255 257
rect 17679 255 17723 297
rect 17773 317 17815 355
rect 17773 297 17787 317
rect 17807 297 17815 317
rect 17773 255 17815 297
rect 17892 317 17936 355
rect 17892 297 17904 317
rect 17924 297 17936 317
rect 17892 255 17936 297
rect 17986 317 18028 355
rect 17986 297 18000 317
rect 18020 297 18028 317
rect 17986 255 18028 297
rect 18100 317 18144 355
rect 18100 297 18112 317
rect 18132 297 18144 317
rect 18100 255 18144 297
rect 18194 317 18236 355
rect 18194 297 18208 317
rect 18228 297 18236 317
rect 18194 255 18236 297
rect 18310 317 18352 355
rect 18310 297 18318 317
rect 18338 297 18352 317
rect 18310 255 18352 297
rect 18402 324 18447 355
rect 18402 317 18446 324
rect 18402 297 18414 317
rect 18434 297 18446 317
rect 18402 255 18446 297
rect 16211 230 16223 250
rect 16243 230 16255 250
rect 16211 188 16255 230
<< ndiffc >>
rect 118 8299 136 8317
rect 4133 8247 4153 8267
rect 4236 8243 4256 8263
rect 4344 8243 4364 8263
rect 4447 8247 4467 8267
rect 4552 8243 4572 8263
rect 4655 8247 4675 8267
rect 4765 8243 4785 8263
rect 4868 8247 4888 8267
rect 5399 8278 5417 8296
rect 5048 8246 5066 8264
rect 120 8200 138 8218
rect 10779 8307 10797 8325
rect 9414 8226 9434 8246
rect 9517 8222 9537 8242
rect 9625 8222 9645 8242
rect 9728 8226 9748 8246
rect 9833 8222 9853 8242
rect 9936 8226 9956 8246
rect 10046 8222 10066 8242
rect 10149 8226 10169 8246
rect 14794 8255 14814 8275
rect 10329 8225 10347 8243
rect 5401 8179 5419 8197
rect 116 8085 134 8103
rect 5050 8147 5068 8165
rect 14897 8251 14917 8271
rect 15005 8251 15025 8271
rect 15108 8255 15128 8275
rect 15213 8251 15233 8271
rect 15316 8255 15336 8275
rect 15426 8251 15446 8271
rect 15529 8255 15549 8275
rect 16060 8286 16078 8304
rect 15709 8254 15727 8272
rect 10781 8208 10799 8226
rect 20075 8234 20095 8254
rect 20178 8230 20198 8250
rect 20286 8230 20306 8250
rect 20389 8234 20409 8254
rect 20494 8230 20514 8250
rect 20597 8234 20617 8254
rect 20707 8230 20727 8250
rect 20810 8234 20830 8254
rect 20990 8233 21008 8251
rect 16062 8187 16080 8205
rect 5055 8045 5073 8063
rect 118 7986 136 8004
rect 3120 8013 3140 8033
rect 3223 8009 3243 8029
rect 3331 8009 3351 8029
rect 3434 8013 3454 8033
rect 3539 8009 3559 8029
rect 3642 8013 3662 8033
rect 3752 8009 3772 8029
rect 3855 8013 3875 8033
rect 5397 8064 5415 8082
rect 304 7915 324 7935
rect 407 7919 427 7939
rect 517 7915 537 7935
rect 620 7919 640 7939
rect 725 7915 745 7935
rect 828 7919 848 7939
rect 936 7919 956 7939
rect 1039 7915 1059 7935
rect 5057 7946 5075 7964
rect 10331 8126 10349 8144
rect 10777 8093 10795 8111
rect 10336 8024 10354 8042
rect 5399 7965 5417 7983
rect 116 7803 134 7821
rect 8401 7992 8421 8012
rect 8504 7988 8524 8008
rect 8612 7988 8632 8008
rect 8715 7992 8735 8012
rect 8820 7988 8840 8008
rect 8923 7992 8943 8012
rect 9033 7988 9053 8008
rect 9136 7992 9156 8012
rect 15711 8155 15729 8173
rect 15716 8053 15734 8071
rect 5585 7894 5605 7914
rect 5688 7898 5708 7918
rect 5798 7894 5818 7914
rect 5901 7898 5921 7918
rect 6006 7894 6026 7914
rect 6109 7898 6129 7918
rect 6217 7898 6237 7918
rect 6320 7894 6340 7914
rect 4132 7832 4152 7852
rect 4235 7828 4255 7848
rect 4343 7828 4363 7848
rect 4446 7832 4466 7852
rect 4551 7828 4571 7848
rect 4654 7832 4674 7852
rect 4764 7828 4784 7848
rect 4867 7832 4887 7852
rect 1316 7734 1336 7754
rect 1419 7738 1439 7758
rect 1529 7734 1549 7754
rect 1632 7738 1652 7758
rect 1737 7734 1757 7754
rect 1840 7738 1860 7758
rect 1948 7738 1968 7758
rect 2051 7734 2071 7754
rect 10779 7994 10797 8012
rect 13781 8021 13801 8041
rect 13884 8017 13904 8037
rect 13992 8017 14012 8037
rect 14095 8021 14115 8041
rect 14200 8017 14220 8037
rect 14303 8021 14323 8041
rect 14413 8017 14433 8037
rect 14516 8021 14536 8041
rect 16058 8072 16076 8090
rect 10338 7925 10356 7943
rect 10965 7923 10985 7943
rect 11068 7927 11088 7947
rect 11178 7923 11198 7943
rect 11281 7927 11301 7947
rect 11386 7923 11406 7943
rect 11489 7927 11509 7947
rect 11597 7927 11617 7947
rect 11700 7923 11720 7943
rect 5055 7763 5073 7781
rect 118 7704 136 7722
rect 123 7602 141 7620
rect 5397 7782 5415 7800
rect 15718 7954 15736 7972
rect 20992 8134 21010 8152
rect 20997 8032 21015 8050
rect 16060 7973 16078 7991
rect 9413 7811 9433 7831
rect 9516 7807 9536 7827
rect 9624 7807 9644 7827
rect 9727 7811 9747 7831
rect 9832 7807 9852 7827
rect 9935 7811 9955 7831
rect 10045 7807 10065 7827
rect 10148 7811 10168 7831
rect 10777 7811 10795 7829
rect 5057 7664 5075 7682
rect 6597 7713 6617 7733
rect 6700 7717 6720 7737
rect 6810 7713 6830 7733
rect 6913 7717 6933 7737
rect 7018 7713 7038 7733
rect 7121 7717 7141 7737
rect 7229 7717 7249 7737
rect 7332 7713 7352 7733
rect 10336 7742 10354 7760
rect 19062 8000 19082 8020
rect 19165 7996 19185 8016
rect 19273 7996 19293 8016
rect 19376 8000 19396 8020
rect 19481 7996 19501 8016
rect 19584 8000 19604 8020
rect 19694 7996 19714 8016
rect 19797 8000 19817 8020
rect 16246 7902 16266 7922
rect 16349 7906 16369 7926
rect 16459 7902 16479 7922
rect 16562 7906 16582 7926
rect 16667 7902 16687 7922
rect 16770 7906 16790 7926
rect 16878 7906 16898 7926
rect 16981 7902 17001 7922
rect 14793 7840 14813 7860
rect 14896 7836 14916 7856
rect 15004 7836 15024 7856
rect 15107 7840 15127 7860
rect 15212 7836 15232 7856
rect 15315 7840 15335 7860
rect 15425 7836 15445 7856
rect 15528 7840 15548 7860
rect 5399 7683 5417 7701
rect 3070 7593 3090 7613
rect 3173 7589 3193 7609
rect 3281 7589 3301 7609
rect 3384 7593 3404 7613
rect 3489 7589 3509 7609
rect 3592 7593 3612 7613
rect 3702 7589 3722 7609
rect 3805 7593 3825 7613
rect 125 7503 143 7521
rect 303 7500 323 7520
rect 406 7504 426 7524
rect 516 7500 536 7520
rect 619 7504 639 7524
rect 724 7500 744 7520
rect 827 7504 847 7524
rect 935 7504 955 7524
rect 1038 7500 1058 7520
rect 5404 7581 5422 7599
rect 11977 7742 11997 7762
rect 12080 7746 12100 7766
rect 12190 7742 12210 7762
rect 12293 7746 12313 7766
rect 12398 7742 12418 7762
rect 12501 7746 12521 7766
rect 12609 7746 12629 7766
rect 12712 7742 12732 7762
rect 20999 7933 21017 7951
rect 15716 7771 15734 7789
rect 10779 7712 10797 7730
rect 10338 7643 10356 7661
rect 10784 7610 10802 7628
rect 16058 7790 16076 7808
rect 20074 7819 20094 7839
rect 20177 7815 20197 7835
rect 20285 7815 20305 7835
rect 20388 7819 20408 7839
rect 20493 7815 20513 7835
rect 20596 7819 20616 7839
rect 20706 7815 20726 7835
rect 20809 7819 20829 7839
rect 15718 7672 15736 7690
rect 17258 7721 17278 7741
rect 17361 7725 17381 7745
rect 17471 7721 17491 7741
rect 17574 7725 17594 7745
rect 17679 7721 17699 7741
rect 17782 7725 17802 7745
rect 17890 7725 17910 7745
rect 17993 7721 18013 7741
rect 20997 7750 21015 7768
rect 16060 7691 16078 7709
rect 5053 7549 5071 7567
rect 8351 7572 8371 7592
rect 8454 7568 8474 7588
rect 8562 7568 8582 7588
rect 8665 7572 8685 7592
rect 8770 7568 8790 7588
rect 8873 7572 8893 7592
rect 8983 7568 9003 7588
rect 9086 7572 9106 7592
rect 5406 7482 5424 7500
rect 5055 7450 5073 7468
rect 5584 7479 5604 7499
rect 5687 7483 5707 7503
rect 5797 7479 5817 7499
rect 5900 7483 5920 7503
rect 6005 7479 6025 7499
rect 6108 7483 6128 7503
rect 6216 7483 6236 7503
rect 6319 7479 6339 7499
rect 10334 7528 10352 7546
rect 13731 7601 13751 7621
rect 13834 7597 13854 7617
rect 13942 7597 13962 7617
rect 14045 7601 14065 7621
rect 14150 7597 14170 7617
rect 14253 7601 14273 7621
rect 14363 7597 14383 7617
rect 14466 7601 14486 7621
rect 10786 7511 10804 7529
rect 10964 7508 10984 7528
rect 11067 7512 11087 7532
rect 11177 7508 11197 7528
rect 11280 7512 11300 7532
rect 11385 7508 11405 7528
rect 11488 7512 11508 7532
rect 11596 7512 11616 7532
rect 11699 7508 11719 7528
rect 16065 7589 16083 7607
rect 20999 7651 21017 7669
rect 15714 7557 15732 7575
rect 10336 7429 10354 7447
rect 19012 7580 19032 7600
rect 19115 7576 19135 7596
rect 19223 7576 19243 7596
rect 19326 7580 19346 7600
rect 19431 7576 19451 7596
rect 19534 7580 19554 7600
rect 19644 7576 19664 7596
rect 19747 7580 19767 7600
rect 16067 7490 16085 7508
rect 15716 7458 15734 7476
rect 16245 7487 16265 7507
rect 16348 7491 16368 7511
rect 16458 7487 16478 7507
rect 16561 7491 16581 7511
rect 16666 7487 16686 7507
rect 16769 7491 16789 7511
rect 16877 7491 16897 7511
rect 16980 7487 17000 7507
rect 20995 7536 21013 7554
rect 20997 7437 21015 7455
rect 123 7318 141 7336
rect 125 7219 143 7237
rect 4138 7266 4158 7286
rect 4241 7262 4261 7282
rect 4349 7262 4369 7282
rect 4452 7266 4472 7286
rect 4557 7262 4577 7282
rect 4660 7266 4680 7286
rect 4770 7262 4790 7282
rect 4873 7266 4893 7286
rect 5404 7297 5422 7315
rect 5053 7265 5071 7283
rect 1371 7173 1391 7193
rect 1474 7177 1494 7197
rect 1584 7173 1604 7193
rect 1687 7177 1707 7197
rect 1792 7173 1812 7193
rect 1895 7177 1915 7197
rect 2003 7177 2023 7197
rect 2106 7173 2126 7193
rect 10784 7326 10802 7344
rect 5406 7198 5424 7216
rect 121 7104 139 7122
rect 5055 7166 5073 7184
rect 9419 7245 9439 7265
rect 9522 7241 9542 7261
rect 9630 7241 9650 7261
rect 9733 7245 9753 7265
rect 9838 7241 9858 7261
rect 9941 7245 9961 7265
rect 10051 7241 10071 7261
rect 10154 7245 10174 7265
rect 10334 7244 10352 7262
rect 6652 7152 6672 7172
rect 6755 7156 6775 7176
rect 6865 7152 6885 7172
rect 6968 7156 6988 7176
rect 7073 7152 7093 7172
rect 7176 7156 7196 7176
rect 7284 7156 7304 7176
rect 7387 7152 7407 7172
rect 10786 7227 10804 7245
rect 14799 7274 14819 7294
rect 14902 7270 14922 7290
rect 15010 7270 15030 7290
rect 15113 7274 15133 7294
rect 15218 7270 15238 7290
rect 15321 7274 15341 7294
rect 15431 7270 15451 7290
rect 15534 7274 15554 7294
rect 16065 7305 16083 7323
rect 15714 7273 15732 7291
rect 12032 7181 12052 7201
rect 12135 7185 12155 7205
rect 12245 7181 12265 7201
rect 12348 7185 12368 7205
rect 12453 7181 12473 7201
rect 12556 7185 12576 7205
rect 12664 7185 12684 7205
rect 12767 7181 12787 7201
rect 16067 7206 16085 7224
rect 5060 7064 5078 7082
rect 123 7005 141 7023
rect 3125 7032 3145 7052
rect 3228 7028 3248 7048
rect 3336 7028 3356 7048
rect 3439 7032 3459 7052
rect 3544 7028 3564 7048
rect 3647 7032 3667 7052
rect 3757 7028 3777 7048
rect 3860 7032 3880 7052
rect 5402 7083 5420 7101
rect 309 6934 329 6954
rect 412 6938 432 6958
rect 522 6934 542 6954
rect 625 6938 645 6958
rect 730 6934 750 6954
rect 833 6938 853 6958
rect 941 6938 961 6958
rect 1044 6934 1064 6954
rect 5062 6965 5080 6983
rect 10336 7145 10354 7163
rect 10782 7112 10800 7130
rect 10341 7043 10359 7061
rect 5404 6984 5422 7002
rect 121 6822 139 6840
rect 8406 7011 8426 7031
rect 8509 7007 8529 7027
rect 8617 7007 8637 7027
rect 8720 7011 8740 7031
rect 8825 7007 8845 7027
rect 8928 7011 8948 7031
rect 9038 7007 9058 7027
rect 9141 7011 9161 7031
rect 15716 7174 15734 7192
rect 20080 7253 20100 7273
rect 20183 7249 20203 7269
rect 20291 7249 20311 7269
rect 20394 7253 20414 7273
rect 20499 7249 20519 7269
rect 20602 7253 20622 7273
rect 20712 7249 20732 7269
rect 20815 7253 20835 7273
rect 20995 7252 21013 7270
rect 17313 7160 17333 7180
rect 17416 7164 17436 7184
rect 17526 7160 17546 7180
rect 17629 7164 17649 7184
rect 17734 7160 17754 7180
rect 17837 7164 17857 7184
rect 17945 7164 17965 7184
rect 18048 7160 18068 7180
rect 15721 7072 15739 7090
rect 5590 6913 5610 6933
rect 5693 6917 5713 6937
rect 5803 6913 5823 6933
rect 5906 6917 5926 6937
rect 6011 6913 6031 6933
rect 6114 6917 6134 6937
rect 6222 6917 6242 6937
rect 6325 6913 6345 6933
rect 4137 6851 4157 6871
rect 4240 6847 4260 6867
rect 4348 6847 4368 6867
rect 4451 6851 4471 6871
rect 4556 6847 4576 6867
rect 4659 6851 4679 6871
rect 4769 6847 4789 6867
rect 4872 6851 4892 6871
rect 1321 6753 1341 6773
rect 1424 6757 1444 6777
rect 1534 6753 1554 6773
rect 1637 6757 1657 6777
rect 1742 6753 1762 6773
rect 1845 6757 1865 6777
rect 1953 6757 1973 6777
rect 2056 6753 2076 6773
rect 10784 7013 10802 7031
rect 13786 7040 13806 7060
rect 13889 7036 13909 7056
rect 13997 7036 14017 7056
rect 14100 7040 14120 7060
rect 14205 7036 14225 7056
rect 14308 7040 14328 7060
rect 14418 7036 14438 7056
rect 14521 7040 14541 7060
rect 16063 7091 16081 7109
rect 10343 6944 10361 6962
rect 10970 6942 10990 6962
rect 11073 6946 11093 6966
rect 11183 6942 11203 6962
rect 11286 6946 11306 6966
rect 11391 6942 11411 6962
rect 11494 6946 11514 6966
rect 11602 6946 11622 6966
rect 11705 6942 11725 6962
rect 5060 6782 5078 6800
rect 123 6723 141 6741
rect 128 6621 146 6639
rect 5402 6801 5420 6819
rect 15723 6973 15741 6991
rect 20997 7153 21015 7171
rect 21002 7051 21020 7069
rect 16065 6992 16083 7010
rect 9418 6830 9438 6850
rect 9521 6826 9541 6846
rect 9629 6826 9649 6846
rect 9732 6830 9752 6850
rect 9837 6826 9857 6846
rect 9940 6830 9960 6850
rect 10050 6826 10070 6846
rect 10153 6830 10173 6850
rect 10782 6830 10800 6848
rect 5062 6683 5080 6701
rect 6602 6732 6622 6752
rect 6705 6736 6725 6756
rect 6815 6732 6835 6752
rect 6918 6736 6938 6756
rect 7023 6732 7043 6752
rect 7126 6736 7146 6756
rect 7234 6736 7254 6756
rect 7337 6732 7357 6752
rect 10341 6761 10359 6779
rect 19067 7019 19087 7039
rect 19170 7015 19190 7035
rect 19278 7015 19298 7035
rect 19381 7019 19401 7039
rect 19486 7015 19506 7035
rect 19589 7019 19609 7039
rect 19699 7015 19719 7035
rect 19802 7019 19822 7039
rect 16251 6921 16271 6941
rect 16354 6925 16374 6945
rect 16464 6921 16484 6941
rect 16567 6925 16587 6945
rect 16672 6921 16692 6941
rect 16775 6925 16795 6945
rect 16883 6925 16903 6945
rect 16986 6921 17006 6941
rect 14798 6859 14818 6879
rect 14901 6855 14921 6875
rect 15009 6855 15029 6875
rect 15112 6859 15132 6879
rect 15217 6855 15237 6875
rect 15320 6859 15340 6879
rect 15430 6855 15450 6875
rect 15533 6859 15553 6879
rect 5404 6702 5422 6720
rect 2917 6565 2937 6585
rect 3020 6561 3040 6581
rect 3128 6561 3148 6581
rect 3231 6565 3251 6585
rect 3336 6561 3356 6581
rect 3439 6565 3459 6585
rect 3549 6561 3569 6581
rect 3652 6565 3672 6585
rect 5409 6600 5427 6618
rect 11982 6761 12002 6781
rect 12085 6765 12105 6785
rect 12195 6761 12215 6781
rect 12298 6765 12318 6785
rect 12403 6761 12423 6781
rect 12506 6765 12526 6785
rect 12614 6765 12634 6785
rect 12717 6761 12737 6781
rect 21004 6952 21022 6970
rect 15721 6790 15739 6808
rect 10784 6731 10802 6749
rect 10343 6662 10361 6680
rect 10789 6629 10807 6647
rect 16063 6809 16081 6827
rect 20079 6838 20099 6858
rect 20182 6834 20202 6854
rect 20290 6834 20310 6854
rect 20393 6838 20413 6858
rect 20498 6834 20518 6854
rect 20601 6838 20621 6858
rect 20711 6834 20731 6854
rect 20814 6838 20834 6858
rect 15723 6691 15741 6709
rect 17263 6740 17283 6760
rect 17366 6744 17386 6764
rect 17476 6740 17496 6760
rect 17579 6744 17599 6764
rect 17684 6740 17704 6760
rect 17787 6744 17807 6764
rect 17895 6744 17915 6764
rect 17998 6740 18018 6760
rect 21002 6769 21020 6787
rect 16065 6710 16083 6728
rect 5058 6568 5076 6586
rect 130 6522 148 6540
rect 308 6519 328 6539
rect 411 6523 431 6543
rect 521 6519 541 6539
rect 624 6523 644 6543
rect 729 6519 749 6539
rect 832 6523 852 6543
rect 940 6523 960 6543
rect 1043 6519 1063 6539
rect 8198 6544 8218 6564
rect 8301 6540 8321 6560
rect 8409 6540 8429 6560
rect 8512 6544 8532 6564
rect 8617 6540 8637 6560
rect 8720 6544 8740 6564
rect 8830 6540 8850 6560
rect 8933 6544 8953 6564
rect 10339 6547 10357 6565
rect 5411 6501 5429 6519
rect 130 6339 148 6357
rect 5060 6469 5078 6487
rect 5589 6498 5609 6518
rect 5692 6502 5712 6522
rect 5802 6498 5822 6518
rect 5905 6502 5925 6522
rect 6010 6498 6030 6518
rect 6113 6502 6133 6522
rect 6221 6502 6241 6522
rect 6324 6498 6344 6518
rect 13578 6573 13598 6593
rect 13681 6569 13701 6589
rect 13789 6569 13809 6589
rect 13892 6573 13912 6593
rect 13997 6569 14017 6589
rect 14100 6573 14120 6593
rect 14210 6569 14230 6589
rect 14313 6573 14333 6593
rect 16070 6608 16088 6626
rect 21004 6670 21022 6688
rect 15719 6576 15737 6594
rect 10791 6530 10809 6548
rect 10969 6527 10989 6547
rect 11072 6531 11092 6551
rect 11182 6527 11202 6547
rect 11285 6531 11305 6551
rect 11390 6527 11410 6547
rect 11493 6531 11513 6551
rect 11601 6531 11621 6551
rect 11704 6527 11724 6547
rect 18859 6552 18879 6572
rect 18962 6548 18982 6568
rect 19070 6548 19090 6568
rect 19173 6552 19193 6572
rect 19278 6548 19298 6568
rect 19381 6552 19401 6572
rect 19491 6548 19511 6568
rect 19594 6552 19614 6572
rect 21000 6555 21018 6573
rect 16072 6509 16090 6527
rect 4145 6287 4165 6307
rect 4248 6283 4268 6303
rect 4356 6283 4376 6303
rect 4459 6287 4479 6307
rect 4564 6283 4584 6303
rect 4667 6287 4687 6307
rect 4777 6283 4797 6303
rect 4880 6287 4900 6307
rect 5411 6318 5429 6336
rect 10341 6448 10359 6466
rect 10791 6347 10809 6365
rect 15721 6477 15739 6495
rect 16250 6506 16270 6526
rect 16353 6510 16373 6530
rect 16463 6506 16483 6526
rect 16566 6510 16586 6530
rect 16671 6506 16691 6526
rect 16774 6510 16794 6530
rect 16882 6510 16902 6530
rect 16985 6506 17005 6526
rect 5060 6286 5078 6304
rect 132 6240 150 6258
rect 1536 6241 1556 6261
rect 1639 6245 1659 6265
rect 1749 6241 1769 6261
rect 1852 6245 1872 6265
rect 1957 6241 1977 6261
rect 2060 6245 2080 6265
rect 2168 6245 2188 6265
rect 2271 6241 2291 6261
rect 9426 6266 9446 6286
rect 9529 6262 9549 6282
rect 9637 6262 9657 6282
rect 9740 6266 9760 6286
rect 9845 6262 9865 6282
rect 9948 6266 9968 6286
rect 10058 6262 10078 6282
rect 10161 6266 10181 6286
rect 10341 6265 10359 6283
rect 5413 6219 5431 6237
rect 128 6125 146 6143
rect 5062 6187 5080 6205
rect 6817 6220 6837 6240
rect 6920 6224 6940 6244
rect 7030 6220 7050 6240
rect 7133 6224 7153 6244
rect 7238 6220 7258 6240
rect 7341 6224 7361 6244
rect 7449 6224 7469 6244
rect 7552 6220 7572 6240
rect 14806 6295 14826 6315
rect 14909 6291 14929 6311
rect 15017 6291 15037 6311
rect 15120 6295 15140 6315
rect 15225 6291 15245 6311
rect 15328 6295 15348 6315
rect 15438 6291 15458 6311
rect 15541 6295 15561 6315
rect 16072 6326 16090 6344
rect 21002 6456 21020 6474
rect 15721 6294 15739 6312
rect 10793 6248 10811 6266
rect 12197 6249 12217 6269
rect 12300 6253 12320 6273
rect 12410 6249 12430 6269
rect 12513 6253 12533 6273
rect 12618 6249 12638 6269
rect 12721 6253 12741 6273
rect 12829 6253 12849 6273
rect 12932 6249 12952 6269
rect 20087 6274 20107 6294
rect 20190 6270 20210 6290
rect 20298 6270 20318 6290
rect 20401 6274 20421 6294
rect 20506 6270 20526 6290
rect 20609 6274 20629 6294
rect 20719 6270 20739 6290
rect 20822 6274 20842 6294
rect 21002 6273 21020 6291
rect 16074 6227 16092 6245
rect 5067 6085 5085 6103
rect 130 6026 148 6044
rect 3132 6053 3152 6073
rect 3235 6049 3255 6069
rect 3343 6049 3363 6069
rect 3446 6053 3466 6073
rect 3551 6049 3571 6069
rect 3654 6053 3674 6073
rect 3764 6049 3784 6069
rect 3867 6053 3887 6073
rect 5409 6104 5427 6122
rect 316 5955 336 5975
rect 419 5959 439 5979
rect 529 5955 549 5975
rect 632 5959 652 5979
rect 737 5955 757 5975
rect 840 5959 860 5979
rect 948 5959 968 5979
rect 1051 5955 1071 5975
rect 5069 5986 5087 6004
rect 10343 6166 10361 6184
rect 10789 6133 10807 6151
rect 10348 6064 10366 6082
rect 5411 6005 5429 6023
rect 128 5843 146 5861
rect 8413 6032 8433 6052
rect 8516 6028 8536 6048
rect 8624 6028 8644 6048
rect 8727 6032 8747 6052
rect 8832 6028 8852 6048
rect 8935 6032 8955 6052
rect 9045 6028 9065 6048
rect 9148 6032 9168 6052
rect 15723 6195 15741 6213
rect 17478 6228 17498 6248
rect 17581 6232 17601 6252
rect 17691 6228 17711 6248
rect 17794 6232 17814 6252
rect 17899 6228 17919 6248
rect 18002 6232 18022 6252
rect 18110 6232 18130 6252
rect 18213 6228 18233 6248
rect 15728 6093 15746 6111
rect 5597 5934 5617 5954
rect 5700 5938 5720 5958
rect 5810 5934 5830 5954
rect 5913 5938 5933 5958
rect 6018 5934 6038 5954
rect 6121 5938 6141 5958
rect 6229 5938 6249 5958
rect 6332 5934 6352 5954
rect 4144 5872 4164 5892
rect 4247 5868 4267 5888
rect 4355 5868 4375 5888
rect 4458 5872 4478 5892
rect 4563 5868 4583 5888
rect 4666 5872 4686 5892
rect 4776 5868 4796 5888
rect 4879 5872 4899 5892
rect 1328 5774 1348 5794
rect 1431 5778 1451 5798
rect 1541 5774 1561 5794
rect 1644 5778 1664 5798
rect 1749 5774 1769 5794
rect 1852 5778 1872 5798
rect 1960 5778 1980 5798
rect 2063 5774 2083 5794
rect 10791 6034 10809 6052
rect 13793 6061 13813 6081
rect 13896 6057 13916 6077
rect 14004 6057 14024 6077
rect 14107 6061 14127 6081
rect 14212 6057 14232 6077
rect 14315 6061 14335 6081
rect 14425 6057 14445 6077
rect 14528 6061 14548 6081
rect 16070 6112 16088 6130
rect 10350 5965 10368 5983
rect 10977 5963 10997 5983
rect 11080 5967 11100 5987
rect 11190 5963 11210 5983
rect 11293 5967 11313 5987
rect 11398 5963 11418 5983
rect 11501 5967 11521 5987
rect 11609 5967 11629 5987
rect 11712 5963 11732 5983
rect 5067 5803 5085 5821
rect 130 5744 148 5762
rect 135 5642 153 5660
rect 5409 5822 5427 5840
rect 15730 5994 15748 6012
rect 21004 6174 21022 6192
rect 21009 6072 21027 6090
rect 16072 6013 16090 6031
rect 9425 5851 9445 5871
rect 9528 5847 9548 5867
rect 9636 5847 9656 5867
rect 9739 5851 9759 5871
rect 9844 5847 9864 5867
rect 9947 5851 9967 5871
rect 10057 5847 10077 5867
rect 10160 5851 10180 5871
rect 10789 5851 10807 5869
rect 5069 5704 5087 5722
rect 6609 5753 6629 5773
rect 6712 5757 6732 5777
rect 6822 5753 6842 5773
rect 6925 5757 6945 5777
rect 7030 5753 7050 5773
rect 7133 5757 7153 5777
rect 7241 5757 7261 5777
rect 7344 5753 7364 5773
rect 10348 5782 10366 5800
rect 19074 6040 19094 6060
rect 19177 6036 19197 6056
rect 19285 6036 19305 6056
rect 19388 6040 19408 6060
rect 19493 6036 19513 6056
rect 19596 6040 19616 6060
rect 19706 6036 19726 6056
rect 19809 6040 19829 6060
rect 16258 5942 16278 5962
rect 16361 5946 16381 5966
rect 16471 5942 16491 5962
rect 16574 5946 16594 5966
rect 16679 5942 16699 5962
rect 16782 5946 16802 5966
rect 16890 5946 16910 5966
rect 16993 5942 17013 5962
rect 14805 5880 14825 5900
rect 14908 5876 14928 5896
rect 15016 5876 15036 5896
rect 15119 5880 15139 5900
rect 15224 5876 15244 5896
rect 15327 5880 15347 5900
rect 15437 5876 15457 5896
rect 15540 5880 15560 5900
rect 5411 5723 5429 5741
rect 3082 5633 3102 5653
rect 3185 5629 3205 5649
rect 3293 5629 3313 5649
rect 3396 5633 3416 5653
rect 3501 5629 3521 5649
rect 3604 5633 3624 5653
rect 3714 5629 3734 5649
rect 3817 5633 3837 5653
rect 137 5543 155 5561
rect 315 5540 335 5560
rect 418 5544 438 5564
rect 528 5540 548 5560
rect 631 5544 651 5564
rect 736 5540 756 5560
rect 839 5544 859 5564
rect 947 5544 967 5564
rect 1050 5540 1070 5560
rect 5416 5621 5434 5639
rect 11989 5782 12009 5802
rect 12092 5786 12112 5806
rect 12202 5782 12222 5802
rect 12305 5786 12325 5806
rect 12410 5782 12430 5802
rect 12513 5786 12533 5806
rect 12621 5786 12641 5806
rect 12724 5782 12744 5802
rect 21011 5973 21029 5991
rect 15728 5811 15746 5829
rect 10791 5752 10809 5770
rect 10350 5683 10368 5701
rect 10796 5650 10814 5668
rect 16070 5830 16088 5848
rect 20086 5859 20106 5879
rect 20189 5855 20209 5875
rect 20297 5855 20317 5875
rect 20400 5859 20420 5879
rect 20505 5855 20525 5875
rect 20608 5859 20628 5879
rect 20718 5855 20738 5875
rect 20821 5859 20841 5879
rect 15730 5712 15748 5730
rect 17270 5761 17290 5781
rect 17373 5765 17393 5785
rect 17483 5761 17503 5781
rect 17586 5765 17606 5785
rect 17691 5761 17711 5781
rect 17794 5765 17814 5785
rect 17902 5765 17922 5785
rect 18005 5761 18025 5781
rect 21009 5790 21027 5808
rect 16072 5731 16090 5749
rect 5065 5589 5083 5607
rect 8363 5612 8383 5632
rect 8466 5608 8486 5628
rect 8574 5608 8594 5628
rect 8677 5612 8697 5632
rect 8782 5608 8802 5628
rect 8885 5612 8905 5632
rect 8995 5608 9015 5628
rect 9098 5612 9118 5632
rect 5418 5522 5436 5540
rect 5067 5490 5085 5508
rect 5596 5519 5616 5539
rect 5699 5523 5719 5543
rect 5809 5519 5829 5539
rect 5912 5523 5932 5543
rect 6017 5519 6037 5539
rect 6120 5523 6140 5543
rect 6228 5523 6248 5543
rect 6331 5519 6351 5539
rect 10346 5568 10364 5586
rect 13743 5641 13763 5661
rect 13846 5637 13866 5657
rect 13954 5637 13974 5657
rect 14057 5641 14077 5661
rect 14162 5637 14182 5657
rect 14265 5641 14285 5661
rect 14375 5637 14395 5657
rect 14478 5641 14498 5661
rect 10798 5551 10816 5569
rect 10976 5548 10996 5568
rect 11079 5552 11099 5572
rect 11189 5548 11209 5568
rect 11292 5552 11312 5572
rect 11397 5548 11417 5568
rect 11500 5552 11520 5572
rect 11608 5552 11628 5572
rect 11711 5548 11731 5568
rect 16077 5629 16095 5647
rect 21011 5691 21029 5709
rect 15726 5597 15744 5615
rect 10348 5469 10366 5487
rect 19024 5620 19044 5640
rect 19127 5616 19147 5636
rect 19235 5616 19255 5636
rect 19338 5620 19358 5640
rect 19443 5616 19463 5636
rect 19546 5620 19566 5640
rect 19656 5616 19676 5636
rect 19759 5620 19779 5640
rect 16079 5530 16097 5548
rect 15728 5498 15746 5516
rect 16257 5527 16277 5547
rect 16360 5531 16380 5551
rect 16470 5527 16490 5547
rect 16573 5531 16593 5551
rect 16678 5527 16698 5547
rect 16781 5531 16801 5551
rect 16889 5531 16909 5551
rect 16992 5527 17012 5547
rect 21007 5576 21025 5594
rect 21009 5477 21027 5495
rect 135 5358 153 5376
rect 137 5259 155 5277
rect 4150 5306 4170 5326
rect 4253 5302 4273 5322
rect 4361 5302 4381 5322
rect 4464 5306 4484 5326
rect 4569 5302 4589 5322
rect 4672 5306 4692 5326
rect 4782 5302 4802 5322
rect 4885 5306 4905 5326
rect 5416 5337 5434 5355
rect 5065 5305 5083 5323
rect 1383 5213 1403 5233
rect 1486 5217 1506 5237
rect 1596 5213 1616 5233
rect 1699 5217 1719 5237
rect 1804 5213 1824 5233
rect 1907 5217 1927 5237
rect 2015 5217 2035 5237
rect 2118 5213 2138 5233
rect 10796 5366 10814 5384
rect 5418 5238 5436 5256
rect 133 5144 151 5162
rect 5067 5206 5085 5224
rect 9431 5285 9451 5305
rect 9534 5281 9554 5301
rect 9642 5281 9662 5301
rect 9745 5285 9765 5305
rect 9850 5281 9870 5301
rect 9953 5285 9973 5305
rect 10063 5281 10083 5301
rect 10166 5285 10186 5305
rect 10346 5284 10364 5302
rect 6664 5192 6684 5212
rect 6767 5196 6787 5216
rect 6877 5192 6897 5212
rect 6980 5196 7000 5216
rect 7085 5192 7105 5212
rect 7188 5196 7208 5216
rect 7296 5196 7316 5216
rect 7399 5192 7419 5212
rect 10798 5267 10816 5285
rect 14811 5314 14831 5334
rect 14914 5310 14934 5330
rect 15022 5310 15042 5330
rect 15125 5314 15145 5334
rect 15230 5310 15250 5330
rect 15333 5314 15353 5334
rect 15443 5310 15463 5330
rect 15546 5314 15566 5334
rect 16077 5345 16095 5363
rect 15726 5313 15744 5331
rect 12044 5221 12064 5241
rect 12147 5225 12167 5245
rect 12257 5221 12277 5241
rect 12360 5225 12380 5245
rect 12465 5221 12485 5241
rect 12568 5225 12588 5245
rect 12676 5225 12696 5245
rect 12779 5221 12799 5241
rect 16079 5246 16097 5264
rect 5072 5104 5090 5122
rect 135 5045 153 5063
rect 3137 5072 3157 5092
rect 3240 5068 3260 5088
rect 3348 5068 3368 5088
rect 3451 5072 3471 5092
rect 3556 5068 3576 5088
rect 3659 5072 3679 5092
rect 3769 5068 3789 5088
rect 3872 5072 3892 5092
rect 5414 5123 5432 5141
rect 321 4974 341 4994
rect 424 4978 444 4998
rect 534 4974 554 4994
rect 637 4978 657 4998
rect 742 4974 762 4994
rect 845 4978 865 4998
rect 953 4978 973 4998
rect 1056 4974 1076 4994
rect 5074 5005 5092 5023
rect 10348 5185 10366 5203
rect 10794 5152 10812 5170
rect 10353 5083 10371 5101
rect 5416 5024 5434 5042
rect 133 4862 151 4880
rect 8418 5051 8438 5071
rect 8521 5047 8541 5067
rect 8629 5047 8649 5067
rect 8732 5051 8752 5071
rect 8837 5047 8857 5067
rect 8940 5051 8960 5071
rect 9050 5047 9070 5067
rect 9153 5051 9173 5071
rect 15728 5214 15746 5232
rect 20092 5293 20112 5313
rect 20195 5289 20215 5309
rect 20303 5289 20323 5309
rect 20406 5293 20426 5313
rect 20511 5289 20531 5309
rect 20614 5293 20634 5313
rect 20724 5289 20744 5309
rect 20827 5293 20847 5313
rect 21007 5292 21025 5310
rect 17325 5200 17345 5220
rect 17428 5204 17448 5224
rect 17538 5200 17558 5220
rect 17641 5204 17661 5224
rect 17746 5200 17766 5220
rect 17849 5204 17869 5224
rect 17957 5204 17977 5224
rect 18060 5200 18080 5220
rect 15733 5112 15751 5130
rect 5602 4953 5622 4973
rect 5705 4957 5725 4977
rect 5815 4953 5835 4973
rect 5918 4957 5938 4977
rect 6023 4953 6043 4973
rect 6126 4957 6146 4977
rect 6234 4957 6254 4977
rect 6337 4953 6357 4973
rect 4149 4891 4169 4911
rect 4252 4887 4272 4907
rect 4360 4887 4380 4907
rect 4463 4891 4483 4911
rect 4568 4887 4588 4907
rect 4671 4891 4691 4911
rect 4781 4887 4801 4907
rect 4884 4891 4904 4911
rect 1333 4793 1353 4813
rect 1436 4797 1456 4817
rect 1546 4793 1566 4813
rect 1649 4797 1669 4817
rect 1754 4793 1774 4813
rect 1857 4797 1877 4817
rect 1965 4797 1985 4817
rect 2068 4793 2088 4813
rect 10796 5053 10814 5071
rect 13798 5080 13818 5100
rect 13901 5076 13921 5096
rect 14009 5076 14029 5096
rect 14112 5080 14132 5100
rect 14217 5076 14237 5096
rect 14320 5080 14340 5100
rect 14430 5076 14450 5096
rect 14533 5080 14553 5100
rect 16075 5131 16093 5149
rect 10355 4984 10373 5002
rect 10982 4982 11002 5002
rect 11085 4986 11105 5006
rect 11195 4982 11215 5002
rect 11298 4986 11318 5006
rect 11403 4982 11423 5002
rect 11506 4986 11526 5006
rect 11614 4986 11634 5006
rect 11717 4982 11737 5002
rect 5072 4822 5090 4840
rect 135 4763 153 4781
rect 140 4661 158 4679
rect 5414 4841 5432 4859
rect 15735 5013 15753 5031
rect 21009 5193 21027 5211
rect 21014 5091 21032 5109
rect 16077 5032 16095 5050
rect 9430 4870 9450 4890
rect 9533 4866 9553 4886
rect 9641 4866 9661 4886
rect 9744 4870 9764 4890
rect 9849 4866 9869 4886
rect 9952 4870 9972 4890
rect 10062 4866 10082 4886
rect 10165 4870 10185 4890
rect 10794 4870 10812 4888
rect 5074 4723 5092 4741
rect 6614 4772 6634 4792
rect 6717 4776 6737 4796
rect 6827 4772 6847 4792
rect 6930 4776 6950 4796
rect 7035 4772 7055 4792
rect 7138 4776 7158 4796
rect 7246 4776 7266 4796
rect 7349 4772 7369 4792
rect 10353 4801 10371 4819
rect 19079 5059 19099 5079
rect 19182 5055 19202 5075
rect 19290 5055 19310 5075
rect 19393 5059 19413 5079
rect 19498 5055 19518 5075
rect 19601 5059 19621 5079
rect 19711 5055 19731 5075
rect 19814 5059 19834 5079
rect 16263 4961 16283 4981
rect 16366 4965 16386 4985
rect 16476 4961 16496 4981
rect 16579 4965 16599 4985
rect 16684 4961 16704 4981
rect 16787 4965 16807 4985
rect 16895 4965 16915 4985
rect 16998 4961 17018 4981
rect 14810 4899 14830 4919
rect 14913 4895 14933 4915
rect 15021 4895 15041 4915
rect 15124 4899 15144 4919
rect 15229 4895 15249 4915
rect 15332 4899 15352 4919
rect 15442 4895 15462 4915
rect 15545 4899 15565 4919
rect 5416 4742 5434 4760
rect 2842 4640 2862 4660
rect 2945 4636 2965 4656
rect 3053 4636 3073 4656
rect 3156 4640 3176 4660
rect 3261 4636 3281 4656
rect 3364 4640 3384 4660
rect 3474 4636 3494 4656
rect 3577 4640 3597 4660
rect 5421 4640 5439 4658
rect 11994 4801 12014 4821
rect 12097 4805 12117 4825
rect 12207 4801 12227 4821
rect 12310 4805 12330 4825
rect 12415 4801 12435 4821
rect 12518 4805 12538 4825
rect 12626 4805 12646 4825
rect 12729 4801 12749 4821
rect 21016 4992 21034 5010
rect 15733 4830 15751 4848
rect 10796 4771 10814 4789
rect 10355 4702 10373 4720
rect 10801 4669 10819 4687
rect 16075 4849 16093 4867
rect 20091 4878 20111 4898
rect 20194 4874 20214 4894
rect 20302 4874 20322 4894
rect 20405 4878 20425 4898
rect 20510 4874 20530 4894
rect 20613 4878 20633 4898
rect 20723 4874 20743 4894
rect 20826 4878 20846 4898
rect 15735 4731 15753 4749
rect 17275 4780 17295 4800
rect 17378 4784 17398 4804
rect 17488 4780 17508 4800
rect 17591 4784 17611 4804
rect 17696 4780 17716 4800
rect 17799 4784 17819 4804
rect 17907 4784 17927 4804
rect 18010 4780 18030 4800
rect 21014 4809 21032 4827
rect 16077 4750 16095 4768
rect 142 4562 160 4580
rect 320 4559 340 4579
rect 423 4563 443 4583
rect 533 4559 553 4579
rect 636 4563 656 4583
rect 741 4559 761 4579
rect 844 4563 864 4583
rect 952 4563 972 4583
rect 1055 4559 1075 4579
rect 5070 4608 5088 4626
rect 138 4382 156 4400
rect 8123 4619 8143 4639
rect 8226 4615 8246 4635
rect 8334 4615 8354 4635
rect 8437 4619 8457 4639
rect 8542 4615 8562 4635
rect 8645 4619 8665 4639
rect 8755 4615 8775 4635
rect 8858 4619 8878 4639
rect 5423 4541 5441 4559
rect 5072 4509 5090 4527
rect 5601 4538 5621 4558
rect 5704 4542 5724 4562
rect 5814 4538 5834 4558
rect 5917 4542 5937 4562
rect 6022 4538 6042 4558
rect 6125 4542 6145 4562
rect 6233 4542 6253 4562
rect 6336 4538 6356 4558
rect 10351 4587 10369 4605
rect 13503 4648 13523 4668
rect 13606 4644 13626 4664
rect 13714 4644 13734 4664
rect 13817 4648 13837 4668
rect 13922 4644 13942 4664
rect 14025 4648 14045 4668
rect 14135 4644 14155 4664
rect 14238 4648 14258 4668
rect 16082 4648 16100 4666
rect 21016 4710 21034 4728
rect 10803 4570 10821 4588
rect 140 4283 158 4301
rect 4153 4330 4173 4350
rect 4256 4326 4276 4346
rect 4364 4326 4384 4346
rect 4467 4330 4487 4350
rect 4572 4326 4592 4346
rect 4675 4330 4695 4350
rect 4785 4326 4805 4346
rect 4888 4330 4908 4350
rect 5419 4361 5437 4379
rect 5068 4329 5086 4347
rect 1631 4249 1651 4269
rect 1734 4253 1754 4273
rect 1844 4249 1864 4269
rect 1947 4253 1967 4273
rect 2052 4249 2072 4269
rect 2155 4253 2175 4273
rect 2263 4253 2283 4273
rect 2366 4249 2386 4269
rect 10981 4567 11001 4587
rect 11084 4571 11104 4591
rect 11194 4567 11214 4587
rect 11297 4571 11317 4591
rect 11402 4567 11422 4587
rect 11505 4571 11525 4591
rect 11613 4571 11633 4591
rect 11716 4567 11736 4587
rect 15731 4616 15749 4634
rect 10353 4488 10371 4506
rect 10799 4390 10817 4408
rect 5421 4262 5439 4280
rect 9434 4309 9454 4329
rect 9537 4305 9557 4325
rect 9645 4305 9665 4325
rect 9748 4309 9768 4329
rect 9853 4305 9873 4325
rect 9956 4309 9976 4329
rect 10066 4305 10086 4325
rect 10169 4309 10189 4329
rect 18784 4627 18804 4647
rect 18887 4623 18907 4643
rect 18995 4623 19015 4643
rect 19098 4627 19118 4647
rect 19203 4623 19223 4643
rect 19306 4627 19326 4647
rect 19416 4623 19436 4643
rect 19519 4627 19539 4647
rect 16084 4549 16102 4567
rect 15733 4517 15751 4535
rect 16262 4546 16282 4566
rect 16365 4550 16385 4570
rect 16475 4546 16495 4566
rect 16578 4550 16598 4570
rect 16683 4546 16703 4566
rect 16786 4550 16806 4570
rect 16894 4550 16914 4570
rect 16997 4546 17017 4566
rect 21012 4595 21030 4613
rect 10349 4308 10367 4326
rect 136 4168 154 4186
rect 5070 4230 5088 4248
rect 6912 4228 6932 4248
rect 7015 4232 7035 4252
rect 7125 4228 7145 4248
rect 7228 4232 7248 4252
rect 7333 4228 7353 4248
rect 7436 4232 7456 4252
rect 7544 4232 7564 4252
rect 7647 4228 7667 4248
rect 10801 4291 10819 4309
rect 14814 4338 14834 4358
rect 14917 4334 14937 4354
rect 15025 4334 15045 4354
rect 15128 4338 15148 4358
rect 15233 4334 15253 4354
rect 15336 4338 15356 4358
rect 15446 4334 15466 4354
rect 15549 4338 15569 4358
rect 16080 4369 16098 4387
rect 15729 4337 15747 4355
rect 12292 4257 12312 4277
rect 12395 4261 12415 4281
rect 12505 4257 12525 4277
rect 12608 4261 12628 4281
rect 12713 4257 12733 4277
rect 12816 4261 12836 4281
rect 12924 4261 12944 4281
rect 13027 4257 13047 4277
rect 21014 4496 21032 4514
rect 16082 4270 16100 4288
rect 20095 4317 20115 4337
rect 20198 4313 20218 4333
rect 20306 4313 20326 4333
rect 20409 4317 20429 4337
rect 20514 4313 20534 4333
rect 20617 4317 20637 4337
rect 20727 4313 20747 4333
rect 20830 4317 20850 4337
rect 21010 4316 21028 4334
rect 5075 4128 5093 4146
rect 138 4069 156 4087
rect 3140 4096 3160 4116
rect 3243 4092 3263 4112
rect 3351 4092 3371 4112
rect 3454 4096 3474 4116
rect 3559 4092 3579 4112
rect 3662 4096 3682 4116
rect 3772 4092 3792 4112
rect 3875 4096 3895 4116
rect 5417 4147 5435 4165
rect 324 3998 344 4018
rect 427 4002 447 4022
rect 537 3998 557 4018
rect 640 4002 660 4022
rect 745 3998 765 4018
rect 848 4002 868 4022
rect 956 4002 976 4022
rect 1059 3998 1079 4018
rect 5077 4029 5095 4047
rect 10351 4209 10369 4227
rect 10797 4176 10815 4194
rect 10356 4107 10374 4125
rect 5419 4048 5437 4066
rect 136 3886 154 3904
rect 8421 4075 8441 4095
rect 8524 4071 8544 4091
rect 8632 4071 8652 4091
rect 8735 4075 8755 4095
rect 8840 4071 8860 4091
rect 8943 4075 8963 4095
rect 9053 4071 9073 4091
rect 9156 4075 9176 4095
rect 15731 4238 15749 4256
rect 17573 4236 17593 4256
rect 17676 4240 17696 4260
rect 17786 4236 17806 4256
rect 17889 4240 17909 4260
rect 17994 4236 18014 4256
rect 18097 4240 18117 4260
rect 18205 4240 18225 4260
rect 18308 4236 18328 4256
rect 15736 4136 15754 4154
rect 5605 3977 5625 3997
rect 5708 3981 5728 4001
rect 5818 3977 5838 3997
rect 5921 3981 5941 4001
rect 6026 3977 6046 3997
rect 6129 3981 6149 4001
rect 6237 3981 6257 4001
rect 6340 3977 6360 3997
rect 4152 3915 4172 3935
rect 4255 3911 4275 3931
rect 4363 3911 4383 3931
rect 4466 3915 4486 3935
rect 4571 3911 4591 3931
rect 4674 3915 4694 3935
rect 4784 3911 4804 3931
rect 4887 3915 4907 3935
rect 1336 3817 1356 3837
rect 1439 3821 1459 3841
rect 1549 3817 1569 3837
rect 1652 3821 1672 3841
rect 1757 3817 1777 3837
rect 1860 3821 1880 3841
rect 1968 3821 1988 3841
rect 2071 3817 2091 3837
rect 10799 4077 10817 4095
rect 13801 4104 13821 4124
rect 13904 4100 13924 4120
rect 14012 4100 14032 4120
rect 14115 4104 14135 4124
rect 14220 4100 14240 4120
rect 14323 4104 14343 4124
rect 14433 4100 14453 4120
rect 14536 4104 14556 4124
rect 16078 4155 16096 4173
rect 10358 4008 10376 4026
rect 10985 4006 11005 4026
rect 11088 4010 11108 4030
rect 11198 4006 11218 4026
rect 11301 4010 11321 4030
rect 11406 4006 11426 4026
rect 11509 4010 11529 4030
rect 11617 4010 11637 4030
rect 11720 4006 11740 4026
rect 5075 3846 5093 3864
rect 138 3787 156 3805
rect 143 3685 161 3703
rect 5417 3865 5435 3883
rect 15738 4037 15756 4055
rect 21012 4217 21030 4235
rect 21017 4115 21035 4133
rect 16080 4056 16098 4074
rect 9433 3894 9453 3914
rect 9536 3890 9556 3910
rect 9644 3890 9664 3910
rect 9747 3894 9767 3914
rect 9852 3890 9872 3910
rect 9955 3894 9975 3914
rect 10065 3890 10085 3910
rect 10168 3894 10188 3914
rect 10797 3894 10815 3912
rect 5077 3747 5095 3765
rect 6617 3796 6637 3816
rect 6720 3800 6740 3820
rect 6830 3796 6850 3816
rect 6933 3800 6953 3820
rect 7038 3796 7058 3816
rect 7141 3800 7161 3820
rect 7249 3800 7269 3820
rect 7352 3796 7372 3816
rect 10356 3825 10374 3843
rect 19082 4083 19102 4103
rect 19185 4079 19205 4099
rect 19293 4079 19313 4099
rect 19396 4083 19416 4103
rect 19501 4079 19521 4099
rect 19604 4083 19624 4103
rect 19714 4079 19734 4099
rect 19817 4083 19837 4103
rect 16266 3985 16286 4005
rect 16369 3989 16389 4009
rect 16479 3985 16499 4005
rect 16582 3989 16602 4009
rect 16687 3985 16707 4005
rect 16790 3989 16810 4009
rect 16898 3989 16918 4009
rect 17001 3985 17021 4005
rect 14813 3923 14833 3943
rect 14916 3919 14936 3939
rect 15024 3919 15044 3939
rect 15127 3923 15147 3943
rect 15232 3919 15252 3939
rect 15335 3923 15355 3943
rect 15445 3919 15465 3939
rect 15548 3923 15568 3943
rect 5419 3766 5437 3784
rect 3090 3676 3110 3696
rect 3193 3672 3213 3692
rect 3301 3672 3321 3692
rect 3404 3676 3424 3696
rect 3509 3672 3529 3692
rect 3612 3676 3632 3696
rect 3722 3672 3742 3692
rect 3825 3676 3845 3696
rect 145 3586 163 3604
rect 323 3583 343 3603
rect 426 3587 446 3607
rect 536 3583 556 3603
rect 639 3587 659 3607
rect 744 3583 764 3603
rect 847 3587 867 3607
rect 955 3587 975 3607
rect 1058 3583 1078 3603
rect 5424 3664 5442 3682
rect 11997 3825 12017 3845
rect 12100 3829 12120 3849
rect 12210 3825 12230 3845
rect 12313 3829 12333 3849
rect 12418 3825 12438 3845
rect 12521 3829 12541 3849
rect 12629 3829 12649 3849
rect 12732 3825 12752 3845
rect 21019 4016 21037 4034
rect 15736 3854 15754 3872
rect 10799 3795 10817 3813
rect 10358 3726 10376 3744
rect 10804 3693 10822 3711
rect 16078 3873 16096 3891
rect 20094 3902 20114 3922
rect 20197 3898 20217 3918
rect 20305 3898 20325 3918
rect 20408 3902 20428 3922
rect 20513 3898 20533 3918
rect 20616 3902 20636 3922
rect 20726 3898 20746 3918
rect 20829 3902 20849 3922
rect 15738 3755 15756 3773
rect 17278 3804 17298 3824
rect 17381 3808 17401 3828
rect 17491 3804 17511 3824
rect 17594 3808 17614 3828
rect 17699 3804 17719 3824
rect 17802 3808 17822 3828
rect 17910 3808 17930 3828
rect 18013 3804 18033 3824
rect 21017 3833 21035 3851
rect 16080 3774 16098 3792
rect 5073 3632 5091 3650
rect 8371 3655 8391 3675
rect 8474 3651 8494 3671
rect 8582 3651 8602 3671
rect 8685 3655 8705 3675
rect 8790 3651 8810 3671
rect 8893 3655 8913 3675
rect 9003 3651 9023 3671
rect 9106 3655 9126 3675
rect 5426 3565 5444 3583
rect 5075 3533 5093 3551
rect 5604 3562 5624 3582
rect 5707 3566 5727 3586
rect 5817 3562 5837 3582
rect 5920 3566 5940 3586
rect 6025 3562 6045 3582
rect 6128 3566 6148 3586
rect 6236 3566 6256 3586
rect 6339 3562 6359 3582
rect 10354 3611 10372 3629
rect 13751 3684 13771 3704
rect 13854 3680 13874 3700
rect 13962 3680 13982 3700
rect 14065 3684 14085 3704
rect 14170 3680 14190 3700
rect 14273 3684 14293 3704
rect 14383 3680 14403 3700
rect 14486 3684 14506 3704
rect 10806 3594 10824 3612
rect 10984 3591 11004 3611
rect 11087 3595 11107 3615
rect 11197 3591 11217 3611
rect 11300 3595 11320 3615
rect 11405 3591 11425 3611
rect 11508 3595 11528 3615
rect 11616 3595 11636 3615
rect 11719 3591 11739 3611
rect 16085 3672 16103 3690
rect 21019 3734 21037 3752
rect 15734 3640 15752 3658
rect 10356 3512 10374 3530
rect 19032 3663 19052 3683
rect 19135 3659 19155 3679
rect 19243 3659 19263 3679
rect 19346 3663 19366 3683
rect 19451 3659 19471 3679
rect 19554 3663 19574 3683
rect 19664 3659 19684 3679
rect 19767 3663 19787 3683
rect 16087 3573 16105 3591
rect 15736 3541 15754 3559
rect 16265 3570 16285 3590
rect 16368 3574 16388 3594
rect 16478 3570 16498 3590
rect 16581 3574 16601 3594
rect 16686 3570 16706 3590
rect 16789 3574 16809 3594
rect 16897 3574 16917 3594
rect 17000 3570 17020 3590
rect 21015 3619 21033 3637
rect 21017 3520 21035 3538
rect 143 3401 161 3419
rect 145 3302 163 3320
rect 4158 3349 4178 3369
rect 4261 3345 4281 3365
rect 4369 3345 4389 3365
rect 4472 3349 4492 3369
rect 4577 3345 4597 3365
rect 4680 3349 4700 3369
rect 4790 3345 4810 3365
rect 4893 3349 4913 3369
rect 5424 3380 5442 3398
rect 5073 3348 5091 3366
rect 1391 3256 1411 3276
rect 1494 3260 1514 3280
rect 1604 3256 1624 3276
rect 1707 3260 1727 3280
rect 1812 3256 1832 3276
rect 1915 3260 1935 3280
rect 2023 3260 2043 3280
rect 2126 3256 2146 3276
rect 10804 3409 10822 3427
rect 5426 3281 5444 3299
rect 141 3187 159 3205
rect 5075 3249 5093 3267
rect 9439 3328 9459 3348
rect 9542 3324 9562 3344
rect 9650 3324 9670 3344
rect 9753 3328 9773 3348
rect 9858 3324 9878 3344
rect 9961 3328 9981 3348
rect 10071 3324 10091 3344
rect 10174 3328 10194 3348
rect 10354 3327 10372 3345
rect 6672 3235 6692 3255
rect 6775 3239 6795 3259
rect 6885 3235 6905 3255
rect 6988 3239 7008 3259
rect 7093 3235 7113 3255
rect 7196 3239 7216 3259
rect 7304 3239 7324 3259
rect 7407 3235 7427 3255
rect 10806 3310 10824 3328
rect 14819 3357 14839 3377
rect 14922 3353 14942 3373
rect 15030 3353 15050 3373
rect 15133 3357 15153 3377
rect 15238 3353 15258 3373
rect 15341 3357 15361 3377
rect 15451 3353 15471 3373
rect 15554 3357 15574 3377
rect 16085 3388 16103 3406
rect 15734 3356 15752 3374
rect 12052 3264 12072 3284
rect 12155 3268 12175 3288
rect 12265 3264 12285 3284
rect 12368 3268 12388 3288
rect 12473 3264 12493 3284
rect 12576 3268 12596 3288
rect 12684 3268 12704 3288
rect 12787 3264 12807 3284
rect 16087 3289 16105 3307
rect 5080 3147 5098 3165
rect 143 3088 161 3106
rect 3145 3115 3165 3135
rect 3248 3111 3268 3131
rect 3356 3111 3376 3131
rect 3459 3115 3479 3135
rect 3564 3111 3584 3131
rect 3667 3115 3687 3135
rect 3777 3111 3797 3131
rect 3880 3115 3900 3135
rect 5422 3166 5440 3184
rect 329 3017 349 3037
rect 432 3021 452 3041
rect 542 3017 562 3037
rect 645 3021 665 3041
rect 750 3017 770 3037
rect 853 3021 873 3041
rect 961 3021 981 3041
rect 1064 3017 1084 3037
rect 5082 3048 5100 3066
rect 10356 3228 10374 3246
rect 10802 3195 10820 3213
rect 10361 3126 10379 3144
rect 5424 3067 5442 3085
rect 141 2905 159 2923
rect 8426 3094 8446 3114
rect 8529 3090 8549 3110
rect 8637 3090 8657 3110
rect 8740 3094 8760 3114
rect 8845 3090 8865 3110
rect 8948 3094 8968 3114
rect 9058 3090 9078 3110
rect 9161 3094 9181 3114
rect 15736 3257 15754 3275
rect 20100 3336 20120 3356
rect 20203 3332 20223 3352
rect 20311 3332 20331 3352
rect 20414 3336 20434 3356
rect 20519 3332 20539 3352
rect 20622 3336 20642 3356
rect 20732 3332 20752 3352
rect 20835 3336 20855 3356
rect 21015 3335 21033 3353
rect 17333 3243 17353 3263
rect 17436 3247 17456 3267
rect 17546 3243 17566 3263
rect 17649 3247 17669 3267
rect 17754 3243 17774 3263
rect 17857 3247 17877 3267
rect 17965 3247 17985 3267
rect 18068 3243 18088 3263
rect 15741 3155 15759 3173
rect 5610 2996 5630 3016
rect 5713 3000 5733 3020
rect 5823 2996 5843 3016
rect 5926 3000 5946 3020
rect 6031 2996 6051 3016
rect 6134 3000 6154 3020
rect 6242 3000 6262 3020
rect 6345 2996 6365 3016
rect 4157 2934 4177 2954
rect 4260 2930 4280 2950
rect 4368 2930 4388 2950
rect 4471 2934 4491 2954
rect 4576 2930 4596 2950
rect 4679 2934 4699 2954
rect 4789 2930 4809 2950
rect 4892 2934 4912 2954
rect 1341 2836 1361 2856
rect 1444 2840 1464 2860
rect 1554 2836 1574 2856
rect 1657 2840 1677 2860
rect 1762 2836 1782 2856
rect 1865 2840 1885 2860
rect 1973 2840 1993 2860
rect 2076 2836 2096 2856
rect 10804 3096 10822 3114
rect 13806 3123 13826 3143
rect 13909 3119 13929 3139
rect 14017 3119 14037 3139
rect 14120 3123 14140 3143
rect 14225 3119 14245 3139
rect 14328 3123 14348 3143
rect 14438 3119 14458 3139
rect 14541 3123 14561 3143
rect 16083 3174 16101 3192
rect 10363 3027 10381 3045
rect 10990 3025 11010 3045
rect 11093 3029 11113 3049
rect 11203 3025 11223 3045
rect 11306 3029 11326 3049
rect 11411 3025 11431 3045
rect 11514 3029 11534 3049
rect 11622 3029 11642 3049
rect 11725 3025 11745 3045
rect 5080 2865 5098 2883
rect 143 2806 161 2824
rect 148 2704 166 2722
rect 5422 2884 5440 2902
rect 15743 3056 15761 3074
rect 21017 3236 21035 3254
rect 21022 3134 21040 3152
rect 16085 3075 16103 3093
rect 9438 2913 9458 2933
rect 9541 2909 9561 2929
rect 9649 2909 9669 2929
rect 9752 2913 9772 2933
rect 9857 2909 9877 2929
rect 9960 2913 9980 2933
rect 10070 2909 10090 2929
rect 10173 2913 10193 2933
rect 10802 2913 10820 2931
rect 5082 2766 5100 2784
rect 6622 2815 6642 2835
rect 6725 2819 6745 2839
rect 6835 2815 6855 2835
rect 6938 2819 6958 2839
rect 7043 2815 7063 2835
rect 7146 2819 7166 2839
rect 7254 2819 7274 2839
rect 7357 2815 7377 2835
rect 10361 2844 10379 2862
rect 19087 3102 19107 3122
rect 19190 3098 19210 3118
rect 19298 3098 19318 3118
rect 19401 3102 19421 3122
rect 19506 3098 19526 3118
rect 19609 3102 19629 3122
rect 19719 3098 19739 3118
rect 19822 3102 19842 3122
rect 16271 3004 16291 3024
rect 16374 3008 16394 3028
rect 16484 3004 16504 3024
rect 16587 3008 16607 3028
rect 16692 3004 16712 3024
rect 16795 3008 16815 3028
rect 16903 3008 16923 3028
rect 17006 3004 17026 3024
rect 14818 2942 14838 2962
rect 14921 2938 14941 2958
rect 15029 2938 15049 2958
rect 15132 2942 15152 2962
rect 15237 2938 15257 2958
rect 15340 2942 15360 2962
rect 15450 2938 15470 2958
rect 15553 2942 15573 2962
rect 5424 2785 5442 2803
rect 2937 2648 2957 2668
rect 3040 2644 3060 2664
rect 3148 2644 3168 2664
rect 3251 2648 3271 2668
rect 3356 2644 3376 2664
rect 3459 2648 3479 2668
rect 3569 2644 3589 2664
rect 3672 2648 3692 2668
rect 5429 2683 5447 2701
rect 12002 2844 12022 2864
rect 12105 2848 12125 2868
rect 12215 2844 12235 2864
rect 12318 2848 12338 2868
rect 12423 2844 12443 2864
rect 12526 2848 12546 2868
rect 12634 2848 12654 2868
rect 12737 2844 12757 2864
rect 21024 3035 21042 3053
rect 15741 2873 15759 2891
rect 10804 2814 10822 2832
rect 10363 2745 10381 2763
rect 10809 2712 10827 2730
rect 16083 2892 16101 2910
rect 20099 2921 20119 2941
rect 20202 2917 20222 2937
rect 20310 2917 20330 2937
rect 20413 2921 20433 2941
rect 20518 2917 20538 2937
rect 20621 2921 20641 2941
rect 20731 2917 20751 2937
rect 20834 2921 20854 2941
rect 15743 2774 15761 2792
rect 17283 2823 17303 2843
rect 17386 2827 17406 2847
rect 17496 2823 17516 2843
rect 17599 2827 17619 2847
rect 17704 2823 17724 2843
rect 17807 2827 17827 2847
rect 17915 2827 17935 2847
rect 18018 2823 18038 2843
rect 21022 2852 21040 2870
rect 16085 2793 16103 2811
rect 5078 2651 5096 2669
rect 150 2605 168 2623
rect 328 2602 348 2622
rect 431 2606 451 2626
rect 541 2602 561 2622
rect 644 2606 664 2626
rect 749 2602 769 2622
rect 852 2606 872 2626
rect 960 2606 980 2626
rect 1063 2602 1083 2622
rect 8218 2627 8238 2647
rect 8321 2623 8341 2643
rect 8429 2623 8449 2643
rect 8532 2627 8552 2647
rect 8637 2623 8657 2643
rect 8740 2627 8760 2647
rect 8850 2623 8870 2643
rect 8953 2627 8973 2647
rect 10359 2630 10377 2648
rect 5431 2584 5449 2602
rect 150 2422 168 2440
rect 5080 2552 5098 2570
rect 5609 2581 5629 2601
rect 5712 2585 5732 2605
rect 5822 2581 5842 2601
rect 5925 2585 5945 2605
rect 6030 2581 6050 2601
rect 6133 2585 6153 2605
rect 6241 2585 6261 2605
rect 6344 2581 6364 2601
rect 13598 2656 13618 2676
rect 13701 2652 13721 2672
rect 13809 2652 13829 2672
rect 13912 2656 13932 2676
rect 14017 2652 14037 2672
rect 14120 2656 14140 2676
rect 14230 2652 14250 2672
rect 14333 2656 14353 2676
rect 16090 2691 16108 2709
rect 21024 2753 21042 2771
rect 15739 2659 15757 2677
rect 10811 2613 10829 2631
rect 10989 2610 11009 2630
rect 11092 2614 11112 2634
rect 11202 2610 11222 2630
rect 11305 2614 11325 2634
rect 11410 2610 11430 2630
rect 11513 2614 11533 2634
rect 11621 2614 11641 2634
rect 11724 2610 11744 2630
rect 18879 2635 18899 2655
rect 18982 2631 19002 2651
rect 19090 2631 19110 2651
rect 19193 2635 19213 2655
rect 19298 2631 19318 2651
rect 19401 2635 19421 2655
rect 19511 2631 19531 2651
rect 19614 2635 19634 2655
rect 21020 2638 21038 2656
rect 16092 2592 16110 2610
rect 4165 2370 4185 2390
rect 4268 2366 4288 2386
rect 4376 2366 4396 2386
rect 4479 2370 4499 2390
rect 4584 2366 4604 2386
rect 4687 2370 4707 2390
rect 4797 2366 4817 2386
rect 4900 2370 4920 2390
rect 5431 2401 5449 2419
rect 10361 2531 10379 2549
rect 10811 2430 10829 2448
rect 15741 2560 15759 2578
rect 16270 2589 16290 2609
rect 16373 2593 16393 2613
rect 16483 2589 16503 2609
rect 16586 2593 16606 2613
rect 16691 2589 16711 2609
rect 16794 2593 16814 2613
rect 16902 2593 16922 2613
rect 17005 2589 17025 2609
rect 5080 2369 5098 2387
rect 152 2323 170 2341
rect 1556 2324 1576 2344
rect 1659 2328 1679 2348
rect 1769 2324 1789 2344
rect 1872 2328 1892 2348
rect 1977 2324 1997 2344
rect 2080 2328 2100 2348
rect 2188 2328 2208 2348
rect 2291 2324 2311 2344
rect 9446 2349 9466 2369
rect 9549 2345 9569 2365
rect 9657 2345 9677 2365
rect 9760 2349 9780 2369
rect 9865 2345 9885 2365
rect 9968 2349 9988 2369
rect 10078 2345 10098 2365
rect 10181 2349 10201 2369
rect 10361 2348 10379 2366
rect 5433 2302 5451 2320
rect 148 2208 166 2226
rect 5082 2270 5100 2288
rect 6837 2303 6857 2323
rect 6940 2307 6960 2327
rect 7050 2303 7070 2323
rect 7153 2307 7173 2327
rect 7258 2303 7278 2323
rect 7361 2307 7381 2327
rect 7469 2307 7489 2327
rect 7572 2303 7592 2323
rect 14826 2378 14846 2398
rect 14929 2374 14949 2394
rect 15037 2374 15057 2394
rect 15140 2378 15160 2398
rect 15245 2374 15265 2394
rect 15348 2378 15368 2398
rect 15458 2374 15478 2394
rect 15561 2378 15581 2398
rect 16092 2409 16110 2427
rect 21022 2539 21040 2557
rect 15741 2377 15759 2395
rect 10813 2331 10831 2349
rect 12217 2332 12237 2352
rect 12320 2336 12340 2356
rect 12430 2332 12450 2352
rect 12533 2336 12553 2356
rect 12638 2332 12658 2352
rect 12741 2336 12761 2356
rect 12849 2336 12869 2356
rect 12952 2332 12972 2352
rect 20107 2357 20127 2377
rect 20210 2353 20230 2373
rect 20318 2353 20338 2373
rect 20421 2357 20441 2377
rect 20526 2353 20546 2373
rect 20629 2357 20649 2377
rect 20739 2353 20759 2373
rect 20842 2357 20862 2377
rect 21022 2356 21040 2374
rect 16094 2310 16112 2328
rect 5087 2168 5105 2186
rect 150 2109 168 2127
rect 3152 2136 3172 2156
rect 3255 2132 3275 2152
rect 3363 2132 3383 2152
rect 3466 2136 3486 2156
rect 3571 2132 3591 2152
rect 3674 2136 3694 2156
rect 3784 2132 3804 2152
rect 3887 2136 3907 2156
rect 5429 2187 5447 2205
rect 336 2038 356 2058
rect 439 2042 459 2062
rect 549 2038 569 2058
rect 652 2042 672 2062
rect 757 2038 777 2058
rect 860 2042 880 2062
rect 968 2042 988 2062
rect 1071 2038 1091 2058
rect 5089 2069 5107 2087
rect 10363 2249 10381 2267
rect 10809 2216 10827 2234
rect 10368 2147 10386 2165
rect 5431 2088 5449 2106
rect 148 1926 166 1944
rect 8433 2115 8453 2135
rect 8536 2111 8556 2131
rect 8644 2111 8664 2131
rect 8747 2115 8767 2135
rect 8852 2111 8872 2131
rect 8955 2115 8975 2135
rect 9065 2111 9085 2131
rect 9168 2115 9188 2135
rect 15743 2278 15761 2296
rect 17498 2311 17518 2331
rect 17601 2315 17621 2335
rect 17711 2311 17731 2331
rect 17814 2315 17834 2335
rect 17919 2311 17939 2331
rect 18022 2315 18042 2335
rect 18130 2315 18150 2335
rect 18233 2311 18253 2331
rect 15748 2176 15766 2194
rect 5617 2017 5637 2037
rect 5720 2021 5740 2041
rect 5830 2017 5850 2037
rect 5933 2021 5953 2041
rect 6038 2017 6058 2037
rect 6141 2021 6161 2041
rect 6249 2021 6269 2041
rect 6352 2017 6372 2037
rect 4164 1955 4184 1975
rect 4267 1951 4287 1971
rect 4375 1951 4395 1971
rect 4478 1955 4498 1975
rect 4583 1951 4603 1971
rect 4686 1955 4706 1975
rect 4796 1951 4816 1971
rect 4899 1955 4919 1975
rect 1348 1857 1368 1877
rect 1451 1861 1471 1881
rect 1561 1857 1581 1877
rect 1664 1861 1684 1881
rect 1769 1857 1789 1877
rect 1872 1861 1892 1881
rect 1980 1861 2000 1881
rect 2083 1857 2103 1877
rect 10811 2117 10829 2135
rect 13813 2144 13833 2164
rect 13916 2140 13936 2160
rect 14024 2140 14044 2160
rect 14127 2144 14147 2164
rect 14232 2140 14252 2160
rect 14335 2144 14355 2164
rect 14445 2140 14465 2160
rect 14548 2144 14568 2164
rect 16090 2195 16108 2213
rect 10370 2048 10388 2066
rect 10997 2046 11017 2066
rect 11100 2050 11120 2070
rect 11210 2046 11230 2066
rect 11313 2050 11333 2070
rect 11418 2046 11438 2066
rect 11521 2050 11541 2070
rect 11629 2050 11649 2070
rect 11732 2046 11752 2066
rect 5087 1886 5105 1904
rect 150 1827 168 1845
rect 155 1725 173 1743
rect 5429 1905 5447 1923
rect 15750 2077 15768 2095
rect 21024 2257 21042 2275
rect 21029 2155 21047 2173
rect 16092 2096 16110 2114
rect 9445 1934 9465 1954
rect 9548 1930 9568 1950
rect 9656 1930 9676 1950
rect 9759 1934 9779 1954
rect 9864 1930 9884 1950
rect 9967 1934 9987 1954
rect 10077 1930 10097 1950
rect 10180 1934 10200 1954
rect 10809 1934 10827 1952
rect 5089 1787 5107 1805
rect 6629 1836 6649 1856
rect 6732 1840 6752 1860
rect 6842 1836 6862 1856
rect 6945 1840 6965 1860
rect 7050 1836 7070 1856
rect 7153 1840 7173 1860
rect 7261 1840 7281 1860
rect 7364 1836 7384 1856
rect 10368 1865 10386 1883
rect 19094 2123 19114 2143
rect 19197 2119 19217 2139
rect 19305 2119 19325 2139
rect 19408 2123 19428 2143
rect 19513 2119 19533 2139
rect 19616 2123 19636 2143
rect 19726 2119 19746 2139
rect 19829 2123 19849 2143
rect 16278 2025 16298 2045
rect 16381 2029 16401 2049
rect 16491 2025 16511 2045
rect 16594 2029 16614 2049
rect 16699 2025 16719 2045
rect 16802 2029 16822 2049
rect 16910 2029 16930 2049
rect 17013 2025 17033 2045
rect 14825 1963 14845 1983
rect 14928 1959 14948 1979
rect 15036 1959 15056 1979
rect 15139 1963 15159 1983
rect 15244 1959 15264 1979
rect 15347 1963 15367 1983
rect 15457 1959 15477 1979
rect 15560 1963 15580 1983
rect 5431 1806 5449 1824
rect 3102 1716 3122 1736
rect 3205 1712 3225 1732
rect 3313 1712 3333 1732
rect 3416 1716 3436 1736
rect 3521 1712 3541 1732
rect 3624 1716 3644 1736
rect 3734 1712 3754 1732
rect 3837 1716 3857 1736
rect 157 1626 175 1644
rect 335 1623 355 1643
rect 438 1627 458 1647
rect 548 1623 568 1643
rect 651 1627 671 1647
rect 756 1623 776 1643
rect 859 1627 879 1647
rect 967 1627 987 1647
rect 1070 1623 1090 1643
rect 5436 1704 5454 1722
rect 12009 1865 12029 1885
rect 12112 1869 12132 1889
rect 12222 1865 12242 1885
rect 12325 1869 12345 1889
rect 12430 1865 12450 1885
rect 12533 1869 12553 1889
rect 12641 1869 12661 1889
rect 12744 1865 12764 1885
rect 21031 2056 21049 2074
rect 15748 1894 15766 1912
rect 10811 1835 10829 1853
rect 10370 1766 10388 1784
rect 10816 1733 10834 1751
rect 16090 1913 16108 1931
rect 20106 1942 20126 1962
rect 20209 1938 20229 1958
rect 20317 1938 20337 1958
rect 20420 1942 20440 1962
rect 20525 1938 20545 1958
rect 20628 1942 20648 1962
rect 20738 1938 20758 1958
rect 20841 1942 20861 1962
rect 15750 1795 15768 1813
rect 17290 1844 17310 1864
rect 17393 1848 17413 1868
rect 17503 1844 17523 1864
rect 17606 1848 17626 1868
rect 17711 1844 17731 1864
rect 17814 1848 17834 1868
rect 17922 1848 17942 1868
rect 18025 1844 18045 1864
rect 21029 1873 21047 1891
rect 16092 1814 16110 1832
rect 5085 1672 5103 1690
rect 8383 1695 8403 1715
rect 8486 1691 8506 1711
rect 8594 1691 8614 1711
rect 8697 1695 8717 1715
rect 8802 1691 8822 1711
rect 8905 1695 8925 1715
rect 9015 1691 9035 1711
rect 9118 1695 9138 1715
rect 5438 1605 5456 1623
rect 5087 1573 5105 1591
rect 5616 1602 5636 1622
rect 5719 1606 5739 1626
rect 5829 1602 5849 1622
rect 5932 1606 5952 1626
rect 6037 1602 6057 1622
rect 6140 1606 6160 1626
rect 6248 1606 6268 1626
rect 6351 1602 6371 1622
rect 10366 1651 10384 1669
rect 13763 1724 13783 1744
rect 13866 1720 13886 1740
rect 13974 1720 13994 1740
rect 14077 1724 14097 1744
rect 14182 1720 14202 1740
rect 14285 1724 14305 1744
rect 14395 1720 14415 1740
rect 14498 1724 14518 1744
rect 10818 1634 10836 1652
rect 10996 1631 11016 1651
rect 11099 1635 11119 1655
rect 11209 1631 11229 1651
rect 11312 1635 11332 1655
rect 11417 1631 11437 1651
rect 11520 1635 11540 1655
rect 11628 1635 11648 1655
rect 11731 1631 11751 1651
rect 16097 1712 16115 1730
rect 21031 1774 21049 1792
rect 15746 1680 15764 1698
rect 10368 1552 10386 1570
rect 19044 1703 19064 1723
rect 19147 1699 19167 1719
rect 19255 1699 19275 1719
rect 19358 1703 19378 1723
rect 19463 1699 19483 1719
rect 19566 1703 19586 1723
rect 19676 1699 19696 1719
rect 19779 1703 19799 1723
rect 16099 1613 16117 1631
rect 15748 1581 15766 1599
rect 16277 1610 16297 1630
rect 16380 1614 16400 1634
rect 16490 1610 16510 1630
rect 16593 1614 16613 1634
rect 16698 1610 16718 1630
rect 16801 1614 16821 1634
rect 16909 1614 16929 1634
rect 17012 1610 17032 1630
rect 21027 1659 21045 1677
rect 21029 1560 21047 1578
rect 155 1441 173 1459
rect 157 1342 175 1360
rect 4170 1389 4190 1409
rect 4273 1385 4293 1405
rect 4381 1385 4401 1405
rect 4484 1389 4504 1409
rect 4589 1385 4609 1405
rect 4692 1389 4712 1409
rect 4802 1385 4822 1405
rect 4905 1389 4925 1409
rect 5436 1420 5454 1438
rect 5085 1388 5103 1406
rect 1403 1296 1423 1316
rect 1506 1300 1526 1320
rect 1616 1296 1636 1316
rect 1719 1300 1739 1320
rect 1824 1296 1844 1316
rect 1927 1300 1947 1320
rect 2035 1300 2055 1320
rect 2138 1296 2158 1316
rect 10816 1449 10834 1467
rect 5438 1321 5456 1339
rect 153 1227 171 1245
rect 5087 1289 5105 1307
rect 9451 1368 9471 1388
rect 9554 1364 9574 1384
rect 9662 1364 9682 1384
rect 9765 1368 9785 1388
rect 9870 1364 9890 1384
rect 9973 1368 9993 1388
rect 10083 1364 10103 1384
rect 10186 1368 10206 1388
rect 10366 1367 10384 1385
rect 6684 1275 6704 1295
rect 6787 1279 6807 1299
rect 6897 1275 6917 1295
rect 7000 1279 7020 1299
rect 7105 1275 7125 1295
rect 7208 1279 7228 1299
rect 7316 1279 7336 1299
rect 7419 1275 7439 1295
rect 10818 1350 10836 1368
rect 14831 1397 14851 1417
rect 14934 1393 14954 1413
rect 15042 1393 15062 1413
rect 15145 1397 15165 1417
rect 15250 1393 15270 1413
rect 15353 1397 15373 1417
rect 15463 1393 15483 1413
rect 15566 1397 15586 1417
rect 16097 1428 16115 1446
rect 15746 1396 15764 1414
rect 12064 1304 12084 1324
rect 12167 1308 12187 1328
rect 12277 1304 12297 1324
rect 12380 1308 12400 1328
rect 12485 1304 12505 1324
rect 12588 1308 12608 1328
rect 12696 1308 12716 1328
rect 12799 1304 12819 1324
rect 16099 1329 16117 1347
rect 5092 1187 5110 1205
rect 155 1128 173 1146
rect 3157 1155 3177 1175
rect 3260 1151 3280 1171
rect 3368 1151 3388 1171
rect 3471 1155 3491 1175
rect 3576 1151 3596 1171
rect 3679 1155 3699 1175
rect 3789 1151 3809 1171
rect 3892 1155 3912 1175
rect 5434 1206 5452 1224
rect 341 1057 361 1077
rect 444 1061 464 1081
rect 554 1057 574 1077
rect 657 1061 677 1081
rect 762 1057 782 1077
rect 865 1061 885 1081
rect 973 1061 993 1081
rect 1076 1057 1096 1077
rect 5094 1088 5112 1106
rect 10368 1268 10386 1286
rect 10814 1235 10832 1253
rect 10373 1166 10391 1184
rect 5436 1107 5454 1125
rect 153 945 171 963
rect 8438 1134 8458 1154
rect 8541 1130 8561 1150
rect 8649 1130 8669 1150
rect 8752 1134 8772 1154
rect 8857 1130 8877 1150
rect 8960 1134 8980 1154
rect 9070 1130 9090 1150
rect 9173 1134 9193 1154
rect 15748 1297 15766 1315
rect 20112 1376 20132 1396
rect 20215 1372 20235 1392
rect 20323 1372 20343 1392
rect 20426 1376 20446 1396
rect 20531 1372 20551 1392
rect 20634 1376 20654 1396
rect 20744 1372 20764 1392
rect 20847 1376 20867 1396
rect 21027 1375 21045 1393
rect 17345 1283 17365 1303
rect 17448 1287 17468 1307
rect 17558 1283 17578 1303
rect 17661 1287 17681 1307
rect 17766 1283 17786 1303
rect 17869 1287 17889 1307
rect 17977 1287 17997 1307
rect 18080 1283 18100 1303
rect 15753 1195 15771 1213
rect 5622 1036 5642 1056
rect 5725 1040 5745 1060
rect 5835 1036 5855 1056
rect 5938 1040 5958 1060
rect 6043 1036 6063 1056
rect 6146 1040 6166 1060
rect 6254 1040 6274 1060
rect 6357 1036 6377 1056
rect 4169 974 4189 994
rect 4272 970 4292 990
rect 4380 970 4400 990
rect 4483 974 4503 994
rect 4588 970 4608 990
rect 4691 974 4711 994
rect 4801 970 4821 990
rect 4904 974 4924 994
rect 1353 876 1373 896
rect 1456 880 1476 900
rect 1566 876 1586 896
rect 1669 880 1689 900
rect 1774 876 1794 896
rect 1877 880 1897 900
rect 1985 880 2005 900
rect 2088 876 2108 896
rect 10816 1136 10834 1154
rect 13818 1163 13838 1183
rect 13921 1159 13941 1179
rect 14029 1159 14049 1179
rect 14132 1163 14152 1183
rect 14237 1159 14257 1179
rect 14340 1163 14360 1183
rect 14450 1159 14470 1179
rect 14553 1163 14573 1183
rect 16095 1214 16113 1232
rect 10375 1067 10393 1085
rect 11002 1065 11022 1085
rect 11105 1069 11125 1089
rect 11215 1065 11235 1085
rect 11318 1069 11338 1089
rect 11423 1065 11443 1085
rect 11526 1069 11546 1089
rect 11634 1069 11654 1089
rect 11737 1065 11757 1085
rect 5092 905 5110 923
rect 155 846 173 864
rect 160 744 178 762
rect 5434 924 5452 942
rect 15755 1096 15773 1114
rect 21029 1276 21047 1294
rect 21034 1174 21052 1192
rect 16097 1115 16115 1133
rect 9450 953 9470 973
rect 9553 949 9573 969
rect 9661 949 9681 969
rect 9764 953 9784 973
rect 9869 949 9889 969
rect 9972 953 9992 973
rect 10082 949 10102 969
rect 10185 953 10205 973
rect 10814 953 10832 971
rect 5094 806 5112 824
rect 6634 855 6654 875
rect 6737 859 6757 879
rect 6847 855 6867 875
rect 6950 859 6970 879
rect 7055 855 7075 875
rect 7158 859 7178 879
rect 7266 859 7286 879
rect 7369 855 7389 875
rect 10373 884 10391 902
rect 19099 1142 19119 1162
rect 19202 1138 19222 1158
rect 19310 1138 19330 1158
rect 19413 1142 19433 1162
rect 19518 1138 19538 1158
rect 19621 1142 19641 1162
rect 19731 1138 19751 1158
rect 19834 1142 19854 1162
rect 16283 1044 16303 1064
rect 16386 1048 16406 1068
rect 16496 1044 16516 1064
rect 16599 1048 16619 1068
rect 16704 1044 16724 1064
rect 16807 1048 16827 1068
rect 16915 1048 16935 1068
rect 17018 1044 17038 1064
rect 14830 982 14850 1002
rect 14933 978 14953 998
rect 15041 978 15061 998
rect 15144 982 15164 1002
rect 15249 978 15269 998
rect 15352 982 15372 1002
rect 15462 978 15482 998
rect 15565 982 15585 1002
rect 5436 825 5454 843
rect 5441 723 5459 741
rect 12014 884 12034 904
rect 12117 888 12137 908
rect 12227 884 12247 904
rect 12330 888 12350 908
rect 12435 884 12455 904
rect 12538 888 12558 908
rect 12646 888 12666 908
rect 12749 884 12769 904
rect 21036 1075 21054 1093
rect 15753 913 15771 931
rect 10816 854 10834 872
rect 10375 785 10393 803
rect 10821 752 10839 770
rect 16095 932 16113 950
rect 20111 961 20131 981
rect 20214 957 20234 977
rect 20322 957 20342 977
rect 20425 961 20445 981
rect 20530 957 20550 977
rect 20633 961 20653 981
rect 20743 957 20763 977
rect 20846 961 20866 981
rect 15755 814 15773 832
rect 17295 863 17315 883
rect 17398 867 17418 887
rect 17508 863 17528 883
rect 17611 867 17631 887
rect 17716 863 17736 883
rect 17819 867 17839 887
rect 17927 867 17947 887
rect 18030 863 18050 883
rect 21034 892 21052 910
rect 16097 833 16115 851
rect 5090 691 5108 709
rect 162 645 180 663
rect 340 642 360 662
rect 443 646 463 666
rect 553 642 573 662
rect 656 646 676 666
rect 761 642 781 662
rect 864 646 884 666
rect 972 646 992 666
rect 1075 642 1095 662
rect 10371 670 10389 688
rect 5443 624 5461 642
rect 5092 592 5110 610
rect 5621 621 5641 641
rect 5724 625 5744 645
rect 5834 621 5854 641
rect 5937 625 5957 645
rect 6042 621 6062 641
rect 6145 625 6165 645
rect 6253 625 6273 645
rect 16102 731 16120 749
rect 21036 793 21054 811
rect 15751 699 15769 717
rect 10823 653 10841 671
rect 6356 621 6376 641
rect 11001 650 11021 670
rect 11104 654 11124 674
rect 11214 650 11234 670
rect 11317 654 11337 674
rect 11422 650 11442 670
rect 11525 654 11545 674
rect 11633 654 11653 674
rect 11736 650 11756 670
rect 10373 571 10391 589
rect 21032 678 21050 696
rect 16104 632 16122 650
rect 15753 600 15771 618
rect 16282 629 16302 649
rect 16385 633 16405 653
rect 16495 629 16515 649
rect 16598 633 16618 653
rect 16703 629 16723 649
rect 16806 633 16826 653
rect 16914 633 16934 653
rect 17017 629 17037 649
rect 21034 579 21052 597
rect 1743 161 1763 181
rect 1846 165 1866 185
rect 1956 161 1976 181
rect 2059 165 2079 185
rect 2164 161 2184 181
rect 2267 165 2287 185
rect 2375 165 2395 185
rect 2478 161 2498 181
rect 7024 140 7044 160
rect 7127 144 7147 164
rect 7237 140 7257 160
rect 7340 144 7360 164
rect 7445 140 7465 160
rect 7548 144 7568 164
rect 7656 144 7676 164
rect 7759 140 7779 160
rect 4833 73 4853 93
rect 4936 77 4956 97
rect 5046 73 5066 93
rect 5149 77 5169 97
rect 5254 73 5274 93
rect 5357 77 5377 97
rect 5465 77 5485 97
rect 12404 169 12424 189
rect 12507 173 12527 193
rect 12617 169 12637 189
rect 12720 173 12740 193
rect 12825 169 12845 189
rect 12928 173 12948 193
rect 13036 173 13056 193
rect 13139 169 13159 189
rect 17685 148 17705 168
rect 17788 152 17808 172
rect 17898 148 17918 168
rect 18001 152 18021 172
rect 18106 148 18126 168
rect 18209 152 18229 172
rect 18317 152 18337 172
rect 18420 148 18440 168
rect 5568 73 5588 93
rect 10094 66 10114 86
rect 10197 70 10217 90
rect 10307 66 10327 86
rect 10410 70 10430 90
rect 10515 66 10535 86
rect 10618 70 10638 90
rect 10726 70 10746 90
rect 10829 66 10849 86
rect 15494 81 15514 101
rect 15597 85 15617 105
rect 15707 81 15727 101
rect 15810 85 15830 105
rect 15915 81 15935 101
rect 16018 85 16038 105
rect 16126 85 16146 105
rect 16229 81 16249 101
<< pdiffc >>
rect 310 8064 330 8084
rect 406 8064 426 8084
rect 523 8064 543 8084
rect 619 8064 639 8084
rect 731 8064 751 8084
rect 827 8064 847 8084
rect 937 8064 957 8084
rect 4139 8098 4159 8118
rect 1033 8064 1053 8084
rect 4235 8098 4255 8118
rect 4345 8098 4365 8118
rect 4441 8098 4461 8118
rect 4553 8098 4573 8118
rect 4649 8098 4669 8118
rect 4766 8098 4786 8118
rect 4862 8098 4882 8118
rect 5591 8043 5611 8063
rect 1322 7883 1342 7903
rect 1418 7883 1438 7903
rect 1535 7883 1555 7903
rect 1631 7883 1651 7903
rect 1743 7883 1763 7903
rect 1839 7883 1859 7903
rect 1949 7883 1969 7903
rect 5687 8043 5707 8063
rect 5804 8043 5824 8063
rect 5900 8043 5920 8063
rect 6012 8043 6032 8063
rect 6108 8043 6128 8063
rect 6218 8043 6238 8063
rect 9420 8077 9440 8097
rect 6314 8043 6334 8063
rect 9516 8077 9536 8097
rect 9626 8077 9646 8097
rect 9722 8077 9742 8097
rect 9834 8077 9854 8097
rect 9930 8077 9950 8097
rect 10047 8077 10067 8097
rect 10143 8077 10163 8097
rect 10971 8072 10991 8092
rect 2045 7883 2065 7903
rect 3126 7864 3146 7884
rect 3222 7864 3242 7884
rect 3332 7864 3352 7884
rect 3428 7864 3448 7884
rect 3540 7864 3560 7884
rect 3636 7864 3656 7884
rect 3753 7864 3773 7884
rect 11067 8072 11087 8092
rect 11184 8072 11204 8092
rect 11280 8072 11300 8092
rect 11392 8072 11412 8092
rect 11488 8072 11508 8092
rect 11598 8072 11618 8092
rect 14800 8106 14820 8126
rect 11694 8072 11714 8092
rect 14896 8106 14916 8126
rect 15006 8106 15026 8126
rect 15102 8106 15122 8126
rect 15214 8106 15234 8126
rect 15310 8106 15330 8126
rect 15427 8106 15447 8126
rect 15523 8106 15543 8126
rect 3849 7864 3869 7884
rect 6603 7862 6623 7882
rect 6699 7862 6719 7882
rect 6816 7862 6836 7882
rect 6912 7862 6932 7882
rect 7024 7862 7044 7882
rect 7120 7862 7140 7882
rect 7230 7862 7250 7882
rect 16252 8051 16272 8071
rect 7326 7862 7346 7882
rect 8407 7843 8427 7863
rect 309 7649 329 7669
rect 405 7649 425 7669
rect 522 7649 542 7669
rect 618 7649 638 7669
rect 730 7649 750 7669
rect 826 7649 846 7669
rect 936 7649 956 7669
rect 4138 7683 4158 7703
rect 1032 7649 1052 7669
rect 4234 7683 4254 7703
rect 4344 7683 4364 7703
rect 4440 7683 4460 7703
rect 4552 7683 4572 7703
rect 4648 7683 4668 7703
rect 4765 7683 4785 7703
rect 8503 7843 8523 7863
rect 8613 7843 8633 7863
rect 8709 7843 8729 7863
rect 8821 7843 8841 7863
rect 8917 7843 8937 7863
rect 9034 7843 9054 7863
rect 9130 7843 9150 7863
rect 11983 7891 12003 7911
rect 12079 7891 12099 7911
rect 12196 7891 12216 7911
rect 12292 7891 12312 7911
rect 12404 7891 12424 7911
rect 12500 7891 12520 7911
rect 12610 7891 12630 7911
rect 16348 8051 16368 8071
rect 16465 8051 16485 8071
rect 16561 8051 16581 8071
rect 16673 8051 16693 8071
rect 16769 8051 16789 8071
rect 16879 8051 16899 8071
rect 20081 8085 20101 8105
rect 16975 8051 16995 8071
rect 20177 8085 20197 8105
rect 20287 8085 20307 8105
rect 20383 8085 20403 8105
rect 20495 8085 20515 8105
rect 20591 8085 20611 8105
rect 20708 8085 20728 8105
rect 20804 8085 20824 8105
rect 12706 7891 12726 7911
rect 13787 7872 13807 7892
rect 4861 7683 4881 7703
rect 13883 7872 13903 7892
rect 13993 7872 14013 7892
rect 14089 7872 14109 7892
rect 14201 7872 14221 7892
rect 14297 7872 14317 7892
rect 14414 7872 14434 7892
rect 14510 7872 14530 7892
rect 17264 7870 17284 7890
rect 5590 7628 5610 7648
rect 5686 7628 5706 7648
rect 5803 7628 5823 7648
rect 5899 7628 5919 7648
rect 6011 7628 6031 7648
rect 6107 7628 6127 7648
rect 6217 7628 6237 7648
rect 9419 7662 9439 7682
rect 6313 7628 6333 7648
rect 9515 7662 9535 7682
rect 9625 7662 9645 7682
rect 9721 7662 9741 7682
rect 9833 7662 9853 7682
rect 9929 7662 9949 7682
rect 10046 7662 10066 7682
rect 17360 7870 17380 7890
rect 17477 7870 17497 7890
rect 17573 7870 17593 7890
rect 17685 7870 17705 7890
rect 17781 7870 17801 7890
rect 17891 7870 17911 7890
rect 17987 7870 18007 7890
rect 19068 7851 19088 7871
rect 10142 7662 10162 7682
rect 10970 7657 10990 7677
rect 11066 7657 11086 7677
rect 11183 7657 11203 7677
rect 11279 7657 11299 7677
rect 11391 7657 11411 7677
rect 11487 7657 11507 7677
rect 11597 7657 11617 7677
rect 14799 7691 14819 7711
rect 11693 7657 11713 7677
rect 14895 7691 14915 7711
rect 15005 7691 15025 7711
rect 15101 7691 15121 7711
rect 15213 7691 15233 7711
rect 15309 7691 15329 7711
rect 15426 7691 15446 7711
rect 19164 7851 19184 7871
rect 19274 7851 19294 7871
rect 19370 7851 19390 7871
rect 19482 7851 19502 7871
rect 19578 7851 19598 7871
rect 19695 7851 19715 7871
rect 19791 7851 19811 7871
rect 15522 7691 15542 7711
rect 16251 7636 16271 7656
rect 3076 7444 3096 7464
rect 3172 7444 3192 7464
rect 3282 7444 3302 7464
rect 3378 7444 3398 7464
rect 3490 7444 3510 7464
rect 3586 7444 3606 7464
rect 3703 7444 3723 7464
rect 3799 7444 3819 7464
rect 8357 7423 8377 7443
rect 8453 7423 8473 7443
rect 8563 7423 8583 7443
rect 8659 7423 8679 7443
rect 8771 7423 8791 7443
rect 8867 7423 8887 7443
rect 8984 7423 9004 7443
rect 16347 7636 16367 7656
rect 16464 7636 16484 7656
rect 16560 7636 16580 7656
rect 16672 7636 16692 7656
rect 16768 7636 16788 7656
rect 16878 7636 16898 7656
rect 20080 7670 20100 7690
rect 16974 7636 16994 7656
rect 20176 7670 20196 7690
rect 20286 7670 20306 7690
rect 20382 7670 20402 7690
rect 20494 7670 20514 7690
rect 20590 7670 20610 7690
rect 20707 7670 20727 7690
rect 20803 7670 20823 7690
rect 9080 7423 9100 7443
rect 13737 7452 13757 7472
rect 13833 7452 13853 7472
rect 13943 7452 13963 7472
rect 14039 7452 14059 7472
rect 14151 7452 14171 7472
rect 14247 7452 14267 7472
rect 14364 7452 14384 7472
rect 14460 7452 14480 7472
rect 19018 7431 19038 7451
rect 19114 7431 19134 7451
rect 19224 7431 19244 7451
rect 19320 7431 19340 7451
rect 19432 7431 19452 7451
rect 19528 7431 19548 7451
rect 19645 7431 19665 7451
rect 19741 7431 19761 7451
rect 1377 7322 1397 7342
rect 1473 7322 1493 7342
rect 1590 7322 1610 7342
rect 1686 7322 1706 7342
rect 1798 7322 1818 7342
rect 1894 7322 1914 7342
rect 2004 7322 2024 7342
rect 2100 7322 2120 7342
rect 6658 7301 6678 7321
rect 6754 7301 6774 7321
rect 6871 7301 6891 7321
rect 6967 7301 6987 7321
rect 7079 7301 7099 7321
rect 7175 7301 7195 7321
rect 7285 7301 7305 7321
rect 7381 7301 7401 7321
rect 12038 7330 12058 7350
rect 315 7083 335 7103
rect 411 7083 431 7103
rect 528 7083 548 7103
rect 624 7083 644 7103
rect 736 7083 756 7103
rect 832 7083 852 7103
rect 942 7083 962 7103
rect 4144 7117 4164 7137
rect 1038 7083 1058 7103
rect 4240 7117 4260 7137
rect 4350 7117 4370 7137
rect 4446 7117 4466 7137
rect 4558 7117 4578 7137
rect 4654 7117 4674 7137
rect 4771 7117 4791 7137
rect 12134 7330 12154 7350
rect 12251 7330 12271 7350
rect 12347 7330 12367 7350
rect 12459 7330 12479 7350
rect 12555 7330 12575 7350
rect 12665 7330 12685 7350
rect 12761 7330 12781 7350
rect 17319 7309 17339 7329
rect 17415 7309 17435 7329
rect 17532 7309 17552 7329
rect 17628 7309 17648 7329
rect 17740 7309 17760 7329
rect 17836 7309 17856 7329
rect 17946 7309 17966 7329
rect 18042 7309 18062 7329
rect 4867 7117 4887 7137
rect 5596 7062 5616 7082
rect 1327 6902 1347 6922
rect 1423 6902 1443 6922
rect 1540 6902 1560 6922
rect 1636 6902 1656 6922
rect 1748 6902 1768 6922
rect 1844 6902 1864 6922
rect 1954 6902 1974 6922
rect 5692 7062 5712 7082
rect 5809 7062 5829 7082
rect 5905 7062 5925 7082
rect 6017 7062 6037 7082
rect 6113 7062 6133 7082
rect 6223 7062 6243 7082
rect 9425 7096 9445 7116
rect 6319 7062 6339 7082
rect 9521 7096 9541 7116
rect 9631 7096 9651 7116
rect 9727 7096 9747 7116
rect 9839 7096 9859 7116
rect 9935 7096 9955 7116
rect 10052 7096 10072 7116
rect 10148 7096 10168 7116
rect 10976 7091 10996 7111
rect 2050 6902 2070 6922
rect 3131 6883 3151 6903
rect 3227 6883 3247 6903
rect 3337 6883 3357 6903
rect 3433 6883 3453 6903
rect 3545 6883 3565 6903
rect 3641 6883 3661 6903
rect 3758 6883 3778 6903
rect 11072 7091 11092 7111
rect 11189 7091 11209 7111
rect 11285 7091 11305 7111
rect 11397 7091 11417 7111
rect 11493 7091 11513 7111
rect 11603 7091 11623 7111
rect 14805 7125 14825 7145
rect 11699 7091 11719 7111
rect 14901 7125 14921 7145
rect 15011 7125 15031 7145
rect 15107 7125 15127 7145
rect 15219 7125 15239 7145
rect 15315 7125 15335 7145
rect 15432 7125 15452 7145
rect 15528 7125 15548 7145
rect 3854 6883 3874 6903
rect 6608 6881 6628 6901
rect 6704 6881 6724 6901
rect 6821 6881 6841 6901
rect 6917 6881 6937 6901
rect 7029 6881 7049 6901
rect 7125 6881 7145 6901
rect 7235 6881 7255 6901
rect 16257 7070 16277 7090
rect 7331 6881 7351 6901
rect 8412 6862 8432 6882
rect 314 6668 334 6688
rect 410 6668 430 6688
rect 527 6668 547 6688
rect 623 6668 643 6688
rect 735 6668 755 6688
rect 831 6668 851 6688
rect 941 6668 961 6688
rect 4143 6702 4163 6722
rect 1037 6668 1057 6688
rect 4239 6702 4259 6722
rect 4349 6702 4369 6722
rect 4445 6702 4465 6722
rect 4557 6702 4577 6722
rect 4653 6702 4673 6722
rect 4770 6702 4790 6722
rect 8508 6862 8528 6882
rect 8618 6862 8638 6882
rect 8714 6862 8734 6882
rect 8826 6862 8846 6882
rect 8922 6862 8942 6882
rect 9039 6862 9059 6882
rect 9135 6862 9155 6882
rect 11988 6910 12008 6930
rect 12084 6910 12104 6930
rect 12201 6910 12221 6930
rect 12297 6910 12317 6930
rect 12409 6910 12429 6930
rect 12505 6910 12525 6930
rect 12615 6910 12635 6930
rect 16353 7070 16373 7090
rect 16470 7070 16490 7090
rect 16566 7070 16586 7090
rect 16678 7070 16698 7090
rect 16774 7070 16794 7090
rect 16884 7070 16904 7090
rect 20086 7104 20106 7124
rect 16980 7070 17000 7090
rect 20182 7104 20202 7124
rect 20292 7104 20312 7124
rect 20388 7104 20408 7124
rect 20500 7104 20520 7124
rect 20596 7104 20616 7124
rect 20713 7104 20733 7124
rect 20809 7104 20829 7124
rect 12711 6910 12731 6930
rect 13792 6891 13812 6911
rect 4866 6702 4886 6722
rect 13888 6891 13908 6911
rect 13998 6891 14018 6911
rect 14094 6891 14114 6911
rect 14206 6891 14226 6911
rect 14302 6891 14322 6911
rect 14419 6891 14439 6911
rect 14515 6891 14535 6911
rect 17269 6889 17289 6909
rect 5595 6647 5615 6667
rect 5691 6647 5711 6667
rect 5808 6647 5828 6667
rect 5904 6647 5924 6667
rect 6016 6647 6036 6667
rect 6112 6647 6132 6667
rect 6222 6647 6242 6667
rect 9424 6681 9444 6701
rect 6318 6647 6338 6667
rect 9520 6681 9540 6701
rect 9630 6681 9650 6701
rect 9726 6681 9746 6701
rect 9838 6681 9858 6701
rect 9934 6681 9954 6701
rect 10051 6681 10071 6701
rect 17365 6889 17385 6909
rect 17482 6889 17502 6909
rect 17578 6889 17598 6909
rect 17690 6889 17710 6909
rect 17786 6889 17806 6909
rect 17896 6889 17916 6909
rect 17992 6889 18012 6909
rect 19073 6870 19093 6890
rect 10147 6681 10167 6701
rect 10975 6676 10995 6696
rect 11071 6676 11091 6696
rect 11188 6676 11208 6696
rect 11284 6676 11304 6696
rect 11396 6676 11416 6696
rect 11492 6676 11512 6696
rect 11602 6676 11622 6696
rect 14804 6710 14824 6730
rect 11698 6676 11718 6696
rect 14900 6710 14920 6730
rect 15010 6710 15030 6730
rect 15106 6710 15126 6730
rect 15218 6710 15238 6730
rect 15314 6710 15334 6730
rect 15431 6710 15451 6730
rect 19169 6870 19189 6890
rect 19279 6870 19299 6890
rect 19375 6870 19395 6890
rect 19487 6870 19507 6890
rect 19583 6870 19603 6890
rect 19700 6870 19720 6890
rect 19796 6870 19816 6890
rect 15527 6710 15547 6730
rect 16256 6655 16276 6675
rect 1542 6390 1562 6410
rect 1638 6390 1658 6410
rect 1755 6390 1775 6410
rect 1851 6390 1871 6410
rect 1963 6390 1983 6410
rect 2059 6390 2079 6410
rect 2169 6390 2189 6410
rect 2265 6390 2285 6410
rect 2923 6416 2943 6436
rect 3019 6416 3039 6436
rect 3129 6416 3149 6436
rect 3225 6416 3245 6436
rect 3337 6416 3357 6436
rect 3433 6416 3453 6436
rect 3550 6416 3570 6436
rect 16352 6655 16372 6675
rect 16469 6655 16489 6675
rect 16565 6655 16585 6675
rect 16677 6655 16697 6675
rect 16773 6655 16793 6675
rect 16883 6655 16903 6675
rect 20085 6689 20105 6709
rect 16979 6655 16999 6675
rect 20181 6689 20201 6709
rect 20291 6689 20311 6709
rect 20387 6689 20407 6709
rect 20499 6689 20519 6709
rect 20595 6689 20615 6709
rect 20712 6689 20732 6709
rect 20808 6689 20828 6709
rect 3646 6416 3666 6436
rect 6823 6369 6843 6389
rect 6919 6369 6939 6389
rect 7036 6369 7056 6389
rect 7132 6369 7152 6389
rect 7244 6369 7264 6389
rect 7340 6369 7360 6389
rect 7450 6369 7470 6389
rect 7546 6369 7566 6389
rect 8204 6395 8224 6415
rect 8300 6395 8320 6415
rect 8410 6395 8430 6415
rect 8506 6395 8526 6415
rect 8618 6395 8638 6415
rect 8714 6395 8734 6415
rect 8831 6395 8851 6415
rect 8927 6395 8947 6415
rect 12203 6398 12223 6418
rect 12299 6398 12319 6418
rect 12416 6398 12436 6418
rect 12512 6398 12532 6418
rect 12624 6398 12644 6418
rect 12720 6398 12740 6418
rect 12830 6398 12850 6418
rect 12926 6398 12946 6418
rect 13584 6424 13604 6444
rect 13680 6424 13700 6444
rect 13790 6424 13810 6444
rect 13886 6424 13906 6444
rect 13998 6424 14018 6444
rect 14094 6424 14114 6444
rect 14211 6424 14231 6444
rect 14307 6424 14327 6444
rect 17484 6377 17504 6397
rect 322 6104 342 6124
rect 418 6104 438 6124
rect 535 6104 555 6124
rect 631 6104 651 6124
rect 743 6104 763 6124
rect 839 6104 859 6124
rect 949 6104 969 6124
rect 4151 6138 4171 6158
rect 1045 6104 1065 6124
rect 4247 6138 4267 6158
rect 4357 6138 4377 6158
rect 4453 6138 4473 6158
rect 4565 6138 4585 6158
rect 4661 6138 4681 6158
rect 4778 6138 4798 6158
rect 17580 6377 17600 6397
rect 17697 6377 17717 6397
rect 17793 6377 17813 6397
rect 17905 6377 17925 6397
rect 18001 6377 18021 6397
rect 18111 6377 18131 6397
rect 18207 6377 18227 6397
rect 18865 6403 18885 6423
rect 18961 6403 18981 6423
rect 19071 6403 19091 6423
rect 19167 6403 19187 6423
rect 19279 6403 19299 6423
rect 19375 6403 19395 6423
rect 19492 6403 19512 6423
rect 19588 6403 19608 6423
rect 4874 6138 4894 6158
rect 5603 6083 5623 6103
rect 1334 5923 1354 5943
rect 1430 5923 1450 5943
rect 1547 5923 1567 5943
rect 1643 5923 1663 5943
rect 1755 5923 1775 5943
rect 1851 5923 1871 5943
rect 1961 5923 1981 5943
rect 5699 6083 5719 6103
rect 5816 6083 5836 6103
rect 5912 6083 5932 6103
rect 6024 6083 6044 6103
rect 6120 6083 6140 6103
rect 6230 6083 6250 6103
rect 9432 6117 9452 6137
rect 6326 6083 6346 6103
rect 9528 6117 9548 6137
rect 9638 6117 9658 6137
rect 9734 6117 9754 6137
rect 9846 6117 9866 6137
rect 9942 6117 9962 6137
rect 10059 6117 10079 6137
rect 10155 6117 10175 6137
rect 10983 6112 11003 6132
rect 2057 5923 2077 5943
rect 3138 5904 3158 5924
rect 3234 5904 3254 5924
rect 3344 5904 3364 5924
rect 3440 5904 3460 5924
rect 3552 5904 3572 5924
rect 3648 5904 3668 5924
rect 3765 5904 3785 5924
rect 11079 6112 11099 6132
rect 11196 6112 11216 6132
rect 11292 6112 11312 6132
rect 11404 6112 11424 6132
rect 11500 6112 11520 6132
rect 11610 6112 11630 6132
rect 14812 6146 14832 6166
rect 11706 6112 11726 6132
rect 14908 6146 14928 6166
rect 15018 6146 15038 6166
rect 15114 6146 15134 6166
rect 15226 6146 15246 6166
rect 15322 6146 15342 6166
rect 15439 6146 15459 6166
rect 15535 6146 15555 6166
rect 3861 5904 3881 5924
rect 6615 5902 6635 5922
rect 6711 5902 6731 5922
rect 6828 5902 6848 5922
rect 6924 5902 6944 5922
rect 7036 5902 7056 5922
rect 7132 5902 7152 5922
rect 7242 5902 7262 5922
rect 16264 6091 16284 6111
rect 7338 5902 7358 5922
rect 8419 5883 8439 5903
rect 321 5689 341 5709
rect 417 5689 437 5709
rect 534 5689 554 5709
rect 630 5689 650 5709
rect 742 5689 762 5709
rect 838 5689 858 5709
rect 948 5689 968 5709
rect 4150 5723 4170 5743
rect 1044 5689 1064 5709
rect 4246 5723 4266 5743
rect 4356 5723 4376 5743
rect 4452 5723 4472 5743
rect 4564 5723 4584 5743
rect 4660 5723 4680 5743
rect 4777 5723 4797 5743
rect 8515 5883 8535 5903
rect 8625 5883 8645 5903
rect 8721 5883 8741 5903
rect 8833 5883 8853 5903
rect 8929 5883 8949 5903
rect 9046 5883 9066 5903
rect 9142 5883 9162 5903
rect 11995 5931 12015 5951
rect 12091 5931 12111 5951
rect 12208 5931 12228 5951
rect 12304 5931 12324 5951
rect 12416 5931 12436 5951
rect 12512 5931 12532 5951
rect 12622 5931 12642 5951
rect 16360 6091 16380 6111
rect 16477 6091 16497 6111
rect 16573 6091 16593 6111
rect 16685 6091 16705 6111
rect 16781 6091 16801 6111
rect 16891 6091 16911 6111
rect 20093 6125 20113 6145
rect 16987 6091 17007 6111
rect 20189 6125 20209 6145
rect 20299 6125 20319 6145
rect 20395 6125 20415 6145
rect 20507 6125 20527 6145
rect 20603 6125 20623 6145
rect 20720 6125 20740 6145
rect 20816 6125 20836 6145
rect 12718 5931 12738 5951
rect 13799 5912 13819 5932
rect 4873 5723 4893 5743
rect 13895 5912 13915 5932
rect 14005 5912 14025 5932
rect 14101 5912 14121 5932
rect 14213 5912 14233 5932
rect 14309 5912 14329 5932
rect 14426 5912 14446 5932
rect 14522 5912 14542 5932
rect 17276 5910 17296 5930
rect 5602 5668 5622 5688
rect 5698 5668 5718 5688
rect 5815 5668 5835 5688
rect 5911 5668 5931 5688
rect 6023 5668 6043 5688
rect 6119 5668 6139 5688
rect 6229 5668 6249 5688
rect 9431 5702 9451 5722
rect 6325 5668 6345 5688
rect 9527 5702 9547 5722
rect 9637 5702 9657 5722
rect 9733 5702 9753 5722
rect 9845 5702 9865 5722
rect 9941 5702 9961 5722
rect 10058 5702 10078 5722
rect 17372 5910 17392 5930
rect 17489 5910 17509 5930
rect 17585 5910 17605 5930
rect 17697 5910 17717 5930
rect 17793 5910 17813 5930
rect 17903 5910 17923 5930
rect 17999 5910 18019 5930
rect 19080 5891 19100 5911
rect 10154 5702 10174 5722
rect 10982 5697 11002 5717
rect 11078 5697 11098 5717
rect 11195 5697 11215 5717
rect 11291 5697 11311 5717
rect 11403 5697 11423 5717
rect 11499 5697 11519 5717
rect 11609 5697 11629 5717
rect 14811 5731 14831 5751
rect 11705 5697 11725 5717
rect 14907 5731 14927 5751
rect 15017 5731 15037 5751
rect 15113 5731 15133 5751
rect 15225 5731 15245 5751
rect 15321 5731 15341 5751
rect 15438 5731 15458 5751
rect 19176 5891 19196 5911
rect 19286 5891 19306 5911
rect 19382 5891 19402 5911
rect 19494 5891 19514 5911
rect 19590 5891 19610 5911
rect 19707 5891 19727 5911
rect 19803 5891 19823 5911
rect 15534 5731 15554 5751
rect 16263 5676 16283 5696
rect 3088 5484 3108 5504
rect 3184 5484 3204 5504
rect 3294 5484 3314 5504
rect 3390 5484 3410 5504
rect 3502 5484 3522 5504
rect 3598 5484 3618 5504
rect 3715 5484 3735 5504
rect 3811 5484 3831 5504
rect 8369 5463 8389 5483
rect 8465 5463 8485 5483
rect 8575 5463 8595 5483
rect 8671 5463 8691 5483
rect 8783 5463 8803 5483
rect 8879 5463 8899 5483
rect 8996 5463 9016 5483
rect 16359 5676 16379 5696
rect 16476 5676 16496 5696
rect 16572 5676 16592 5696
rect 16684 5676 16704 5696
rect 16780 5676 16800 5696
rect 16890 5676 16910 5696
rect 20092 5710 20112 5730
rect 16986 5676 17006 5696
rect 20188 5710 20208 5730
rect 20298 5710 20318 5730
rect 20394 5710 20414 5730
rect 20506 5710 20526 5730
rect 20602 5710 20622 5730
rect 20719 5710 20739 5730
rect 20815 5710 20835 5730
rect 9092 5463 9112 5483
rect 13749 5492 13769 5512
rect 13845 5492 13865 5512
rect 13955 5492 13975 5512
rect 14051 5492 14071 5512
rect 14163 5492 14183 5512
rect 14259 5492 14279 5512
rect 14376 5492 14396 5512
rect 14472 5492 14492 5512
rect 19030 5471 19050 5491
rect 19126 5471 19146 5491
rect 19236 5471 19256 5491
rect 19332 5471 19352 5491
rect 19444 5471 19464 5491
rect 19540 5471 19560 5491
rect 19657 5471 19677 5491
rect 19753 5471 19773 5491
rect 1389 5362 1409 5382
rect 1485 5362 1505 5382
rect 1602 5362 1622 5382
rect 1698 5362 1718 5382
rect 1810 5362 1830 5382
rect 1906 5362 1926 5382
rect 2016 5362 2036 5382
rect 2112 5362 2132 5382
rect 6670 5341 6690 5361
rect 6766 5341 6786 5361
rect 6883 5341 6903 5361
rect 6979 5341 6999 5361
rect 7091 5341 7111 5361
rect 7187 5341 7207 5361
rect 7297 5341 7317 5361
rect 7393 5341 7413 5361
rect 12050 5370 12070 5390
rect 327 5123 347 5143
rect 423 5123 443 5143
rect 540 5123 560 5143
rect 636 5123 656 5143
rect 748 5123 768 5143
rect 844 5123 864 5143
rect 954 5123 974 5143
rect 4156 5157 4176 5177
rect 1050 5123 1070 5143
rect 4252 5157 4272 5177
rect 4362 5157 4382 5177
rect 4458 5157 4478 5177
rect 4570 5157 4590 5177
rect 4666 5157 4686 5177
rect 4783 5157 4803 5177
rect 12146 5370 12166 5390
rect 12263 5370 12283 5390
rect 12359 5370 12379 5390
rect 12471 5370 12491 5390
rect 12567 5370 12587 5390
rect 12677 5370 12697 5390
rect 12773 5370 12793 5390
rect 17331 5349 17351 5369
rect 17427 5349 17447 5369
rect 17544 5349 17564 5369
rect 17640 5349 17660 5369
rect 17752 5349 17772 5369
rect 17848 5349 17868 5369
rect 17958 5349 17978 5369
rect 18054 5349 18074 5369
rect 4879 5157 4899 5177
rect 5608 5102 5628 5122
rect 1339 4942 1359 4962
rect 1435 4942 1455 4962
rect 1552 4942 1572 4962
rect 1648 4942 1668 4962
rect 1760 4942 1780 4962
rect 1856 4942 1876 4962
rect 1966 4942 1986 4962
rect 5704 5102 5724 5122
rect 5821 5102 5841 5122
rect 5917 5102 5937 5122
rect 6029 5102 6049 5122
rect 6125 5102 6145 5122
rect 6235 5102 6255 5122
rect 9437 5136 9457 5156
rect 6331 5102 6351 5122
rect 9533 5136 9553 5156
rect 9643 5136 9663 5156
rect 9739 5136 9759 5156
rect 9851 5136 9871 5156
rect 9947 5136 9967 5156
rect 10064 5136 10084 5156
rect 10160 5136 10180 5156
rect 10988 5131 11008 5151
rect 2062 4942 2082 4962
rect 3143 4923 3163 4943
rect 3239 4923 3259 4943
rect 3349 4923 3369 4943
rect 3445 4923 3465 4943
rect 3557 4923 3577 4943
rect 3653 4923 3673 4943
rect 3770 4923 3790 4943
rect 11084 5131 11104 5151
rect 11201 5131 11221 5151
rect 11297 5131 11317 5151
rect 11409 5131 11429 5151
rect 11505 5131 11525 5151
rect 11615 5131 11635 5151
rect 14817 5165 14837 5185
rect 11711 5131 11731 5151
rect 14913 5165 14933 5185
rect 15023 5165 15043 5185
rect 15119 5165 15139 5185
rect 15231 5165 15251 5185
rect 15327 5165 15347 5185
rect 15444 5165 15464 5185
rect 15540 5165 15560 5185
rect 3866 4923 3886 4943
rect 6620 4921 6640 4941
rect 6716 4921 6736 4941
rect 6833 4921 6853 4941
rect 6929 4921 6949 4941
rect 7041 4921 7061 4941
rect 7137 4921 7157 4941
rect 7247 4921 7267 4941
rect 16269 5110 16289 5130
rect 7343 4921 7363 4941
rect 8424 4902 8444 4922
rect 326 4708 346 4728
rect 422 4708 442 4728
rect 539 4708 559 4728
rect 635 4708 655 4728
rect 747 4708 767 4728
rect 843 4708 863 4728
rect 953 4708 973 4728
rect 4155 4742 4175 4762
rect 1049 4708 1069 4728
rect 4251 4742 4271 4762
rect 4361 4742 4381 4762
rect 4457 4742 4477 4762
rect 4569 4742 4589 4762
rect 4665 4742 4685 4762
rect 4782 4742 4802 4762
rect 8520 4902 8540 4922
rect 8630 4902 8650 4922
rect 8726 4902 8746 4922
rect 8838 4902 8858 4922
rect 8934 4902 8954 4922
rect 9051 4902 9071 4922
rect 9147 4902 9167 4922
rect 12000 4950 12020 4970
rect 12096 4950 12116 4970
rect 12213 4950 12233 4970
rect 12309 4950 12329 4970
rect 12421 4950 12441 4970
rect 12517 4950 12537 4970
rect 12627 4950 12647 4970
rect 16365 5110 16385 5130
rect 16482 5110 16502 5130
rect 16578 5110 16598 5130
rect 16690 5110 16710 5130
rect 16786 5110 16806 5130
rect 16896 5110 16916 5130
rect 20098 5144 20118 5164
rect 16992 5110 17012 5130
rect 20194 5144 20214 5164
rect 20304 5144 20324 5164
rect 20400 5144 20420 5164
rect 20512 5144 20532 5164
rect 20608 5144 20628 5164
rect 20725 5144 20745 5164
rect 20821 5144 20841 5164
rect 12723 4950 12743 4970
rect 13804 4931 13824 4951
rect 4878 4742 4898 4762
rect 13900 4931 13920 4951
rect 14010 4931 14030 4951
rect 14106 4931 14126 4951
rect 14218 4931 14238 4951
rect 14314 4931 14334 4951
rect 14431 4931 14451 4951
rect 14527 4931 14547 4951
rect 17281 4929 17301 4949
rect 5607 4687 5627 4707
rect 5703 4687 5723 4707
rect 5820 4687 5840 4707
rect 5916 4687 5936 4707
rect 6028 4687 6048 4707
rect 6124 4687 6144 4707
rect 6234 4687 6254 4707
rect 9436 4721 9456 4741
rect 6330 4687 6350 4707
rect 9532 4721 9552 4741
rect 9642 4721 9662 4741
rect 9738 4721 9758 4741
rect 9850 4721 9870 4741
rect 9946 4721 9966 4741
rect 10063 4721 10083 4741
rect 17377 4929 17397 4949
rect 17494 4929 17514 4949
rect 17590 4929 17610 4949
rect 17702 4929 17722 4949
rect 17798 4929 17818 4949
rect 17908 4929 17928 4949
rect 18004 4929 18024 4949
rect 19085 4910 19105 4930
rect 10159 4721 10179 4741
rect 10987 4716 11007 4736
rect 11083 4716 11103 4736
rect 11200 4716 11220 4736
rect 11296 4716 11316 4736
rect 11408 4716 11428 4736
rect 11504 4716 11524 4736
rect 11614 4716 11634 4736
rect 14816 4750 14836 4770
rect 11710 4716 11730 4736
rect 14912 4750 14932 4770
rect 15022 4750 15042 4770
rect 15118 4750 15138 4770
rect 15230 4750 15250 4770
rect 15326 4750 15346 4770
rect 15443 4750 15463 4770
rect 19181 4910 19201 4930
rect 19291 4910 19311 4930
rect 19387 4910 19407 4930
rect 19499 4910 19519 4930
rect 19595 4910 19615 4930
rect 19712 4910 19732 4930
rect 19808 4910 19828 4930
rect 15539 4750 15559 4770
rect 16268 4695 16288 4715
rect 2848 4491 2868 4511
rect 1637 4398 1657 4418
rect 1733 4398 1753 4418
rect 1850 4398 1870 4418
rect 1946 4398 1966 4418
rect 2058 4398 2078 4418
rect 2154 4398 2174 4418
rect 2264 4398 2284 4418
rect 2944 4491 2964 4511
rect 3054 4491 3074 4511
rect 3150 4491 3170 4511
rect 3262 4491 3282 4511
rect 3358 4491 3378 4511
rect 3475 4491 3495 4511
rect 3571 4491 3591 4511
rect 16364 4695 16384 4715
rect 16481 4695 16501 4715
rect 16577 4695 16597 4715
rect 16689 4695 16709 4715
rect 16785 4695 16805 4715
rect 16895 4695 16915 4715
rect 20097 4729 20117 4749
rect 16991 4695 17011 4715
rect 20193 4729 20213 4749
rect 20303 4729 20323 4749
rect 20399 4729 20419 4749
rect 20511 4729 20531 4749
rect 20607 4729 20627 4749
rect 20724 4729 20744 4749
rect 20820 4729 20840 4749
rect 8129 4470 8149 4490
rect 2360 4398 2380 4418
rect 6918 4377 6938 4397
rect 7014 4377 7034 4397
rect 7131 4377 7151 4397
rect 7227 4377 7247 4397
rect 7339 4377 7359 4397
rect 7435 4377 7455 4397
rect 7545 4377 7565 4397
rect 8225 4470 8245 4490
rect 8335 4470 8355 4490
rect 8431 4470 8451 4490
rect 8543 4470 8563 4490
rect 8639 4470 8659 4490
rect 8756 4470 8776 4490
rect 8852 4470 8872 4490
rect 13509 4499 13529 4519
rect 7641 4377 7661 4397
rect 12298 4406 12318 4426
rect 12394 4406 12414 4426
rect 12511 4406 12531 4426
rect 12607 4406 12627 4426
rect 12719 4406 12739 4426
rect 12815 4406 12835 4426
rect 12925 4406 12945 4426
rect 13605 4499 13625 4519
rect 13715 4499 13735 4519
rect 13811 4499 13831 4519
rect 13923 4499 13943 4519
rect 14019 4499 14039 4519
rect 14136 4499 14156 4519
rect 14232 4499 14252 4519
rect 18790 4478 18810 4498
rect 13021 4406 13041 4426
rect 330 4147 350 4167
rect 426 4147 446 4167
rect 543 4147 563 4167
rect 639 4147 659 4167
rect 751 4147 771 4167
rect 847 4147 867 4167
rect 957 4147 977 4167
rect 4159 4181 4179 4201
rect 1053 4147 1073 4167
rect 4255 4181 4275 4201
rect 4365 4181 4385 4201
rect 4461 4181 4481 4201
rect 4573 4181 4593 4201
rect 4669 4181 4689 4201
rect 4786 4181 4806 4201
rect 17579 4385 17599 4405
rect 17675 4385 17695 4405
rect 17792 4385 17812 4405
rect 17888 4385 17908 4405
rect 18000 4385 18020 4405
rect 18096 4385 18116 4405
rect 18206 4385 18226 4405
rect 18886 4478 18906 4498
rect 18996 4478 19016 4498
rect 19092 4478 19112 4498
rect 19204 4478 19224 4498
rect 19300 4478 19320 4498
rect 19417 4478 19437 4498
rect 19513 4478 19533 4498
rect 18302 4385 18322 4405
rect 4882 4181 4902 4201
rect 5611 4126 5631 4146
rect 1342 3966 1362 3986
rect 1438 3966 1458 3986
rect 1555 3966 1575 3986
rect 1651 3966 1671 3986
rect 1763 3966 1783 3986
rect 1859 3966 1879 3986
rect 1969 3966 1989 3986
rect 5707 4126 5727 4146
rect 5824 4126 5844 4146
rect 5920 4126 5940 4146
rect 6032 4126 6052 4146
rect 6128 4126 6148 4146
rect 6238 4126 6258 4146
rect 9440 4160 9460 4180
rect 6334 4126 6354 4146
rect 9536 4160 9556 4180
rect 9646 4160 9666 4180
rect 9742 4160 9762 4180
rect 9854 4160 9874 4180
rect 9950 4160 9970 4180
rect 10067 4160 10087 4180
rect 10163 4160 10183 4180
rect 10991 4155 11011 4175
rect 2065 3966 2085 3986
rect 3146 3947 3166 3967
rect 3242 3947 3262 3967
rect 3352 3947 3372 3967
rect 3448 3947 3468 3967
rect 3560 3947 3580 3967
rect 3656 3947 3676 3967
rect 3773 3947 3793 3967
rect 11087 4155 11107 4175
rect 11204 4155 11224 4175
rect 11300 4155 11320 4175
rect 11412 4155 11432 4175
rect 11508 4155 11528 4175
rect 11618 4155 11638 4175
rect 14820 4189 14840 4209
rect 11714 4155 11734 4175
rect 14916 4189 14936 4209
rect 15026 4189 15046 4209
rect 15122 4189 15142 4209
rect 15234 4189 15254 4209
rect 15330 4189 15350 4209
rect 15447 4189 15467 4209
rect 15543 4189 15563 4209
rect 3869 3947 3889 3967
rect 6623 3945 6643 3965
rect 6719 3945 6739 3965
rect 6836 3945 6856 3965
rect 6932 3945 6952 3965
rect 7044 3945 7064 3965
rect 7140 3945 7160 3965
rect 7250 3945 7270 3965
rect 16272 4134 16292 4154
rect 7346 3945 7366 3965
rect 8427 3926 8447 3946
rect 329 3732 349 3752
rect 425 3732 445 3752
rect 542 3732 562 3752
rect 638 3732 658 3752
rect 750 3732 770 3752
rect 846 3732 866 3752
rect 956 3732 976 3752
rect 4158 3766 4178 3786
rect 1052 3732 1072 3752
rect 4254 3766 4274 3786
rect 4364 3766 4384 3786
rect 4460 3766 4480 3786
rect 4572 3766 4592 3786
rect 4668 3766 4688 3786
rect 4785 3766 4805 3786
rect 8523 3926 8543 3946
rect 8633 3926 8653 3946
rect 8729 3926 8749 3946
rect 8841 3926 8861 3946
rect 8937 3926 8957 3946
rect 9054 3926 9074 3946
rect 9150 3926 9170 3946
rect 12003 3974 12023 3994
rect 12099 3974 12119 3994
rect 12216 3974 12236 3994
rect 12312 3974 12332 3994
rect 12424 3974 12444 3994
rect 12520 3974 12540 3994
rect 12630 3974 12650 3994
rect 16368 4134 16388 4154
rect 16485 4134 16505 4154
rect 16581 4134 16601 4154
rect 16693 4134 16713 4154
rect 16789 4134 16809 4154
rect 16899 4134 16919 4154
rect 20101 4168 20121 4188
rect 16995 4134 17015 4154
rect 20197 4168 20217 4188
rect 20307 4168 20327 4188
rect 20403 4168 20423 4188
rect 20515 4168 20535 4188
rect 20611 4168 20631 4188
rect 20728 4168 20748 4188
rect 20824 4168 20844 4188
rect 12726 3974 12746 3994
rect 13807 3955 13827 3975
rect 4881 3766 4901 3786
rect 13903 3955 13923 3975
rect 14013 3955 14033 3975
rect 14109 3955 14129 3975
rect 14221 3955 14241 3975
rect 14317 3955 14337 3975
rect 14434 3955 14454 3975
rect 14530 3955 14550 3975
rect 17284 3953 17304 3973
rect 5610 3711 5630 3731
rect 5706 3711 5726 3731
rect 5823 3711 5843 3731
rect 5919 3711 5939 3731
rect 6031 3711 6051 3731
rect 6127 3711 6147 3731
rect 6237 3711 6257 3731
rect 9439 3745 9459 3765
rect 6333 3711 6353 3731
rect 9535 3745 9555 3765
rect 9645 3745 9665 3765
rect 9741 3745 9761 3765
rect 9853 3745 9873 3765
rect 9949 3745 9969 3765
rect 10066 3745 10086 3765
rect 17380 3953 17400 3973
rect 17497 3953 17517 3973
rect 17593 3953 17613 3973
rect 17705 3953 17725 3973
rect 17801 3953 17821 3973
rect 17911 3953 17931 3973
rect 18007 3953 18027 3973
rect 19088 3934 19108 3954
rect 10162 3745 10182 3765
rect 10990 3740 11010 3760
rect 11086 3740 11106 3760
rect 11203 3740 11223 3760
rect 11299 3740 11319 3760
rect 11411 3740 11431 3760
rect 11507 3740 11527 3760
rect 11617 3740 11637 3760
rect 14819 3774 14839 3794
rect 11713 3740 11733 3760
rect 14915 3774 14935 3794
rect 15025 3774 15045 3794
rect 15121 3774 15141 3794
rect 15233 3774 15253 3794
rect 15329 3774 15349 3794
rect 15446 3774 15466 3794
rect 19184 3934 19204 3954
rect 19294 3934 19314 3954
rect 19390 3934 19410 3954
rect 19502 3934 19522 3954
rect 19598 3934 19618 3954
rect 19715 3934 19735 3954
rect 19811 3934 19831 3954
rect 15542 3774 15562 3794
rect 16271 3719 16291 3739
rect 3096 3527 3116 3547
rect 3192 3527 3212 3547
rect 3302 3527 3322 3547
rect 3398 3527 3418 3547
rect 3510 3527 3530 3547
rect 3606 3527 3626 3547
rect 3723 3527 3743 3547
rect 3819 3527 3839 3547
rect 8377 3506 8397 3526
rect 8473 3506 8493 3526
rect 8583 3506 8603 3526
rect 8679 3506 8699 3526
rect 8791 3506 8811 3526
rect 8887 3506 8907 3526
rect 9004 3506 9024 3526
rect 16367 3719 16387 3739
rect 16484 3719 16504 3739
rect 16580 3719 16600 3739
rect 16692 3719 16712 3739
rect 16788 3719 16808 3739
rect 16898 3719 16918 3739
rect 20100 3753 20120 3773
rect 16994 3719 17014 3739
rect 20196 3753 20216 3773
rect 20306 3753 20326 3773
rect 20402 3753 20422 3773
rect 20514 3753 20534 3773
rect 20610 3753 20630 3773
rect 20727 3753 20747 3773
rect 20823 3753 20843 3773
rect 9100 3506 9120 3526
rect 13757 3535 13777 3555
rect 13853 3535 13873 3555
rect 13963 3535 13983 3555
rect 14059 3535 14079 3555
rect 14171 3535 14191 3555
rect 14267 3535 14287 3555
rect 14384 3535 14404 3555
rect 14480 3535 14500 3555
rect 19038 3514 19058 3534
rect 19134 3514 19154 3534
rect 19244 3514 19264 3534
rect 19340 3514 19360 3534
rect 19452 3514 19472 3534
rect 19548 3514 19568 3534
rect 19665 3514 19685 3534
rect 19761 3514 19781 3534
rect 1397 3405 1417 3425
rect 1493 3405 1513 3425
rect 1610 3405 1630 3425
rect 1706 3405 1726 3425
rect 1818 3405 1838 3425
rect 1914 3405 1934 3425
rect 2024 3405 2044 3425
rect 2120 3405 2140 3425
rect 6678 3384 6698 3404
rect 6774 3384 6794 3404
rect 6891 3384 6911 3404
rect 6987 3384 7007 3404
rect 7099 3384 7119 3404
rect 7195 3384 7215 3404
rect 7305 3384 7325 3404
rect 7401 3384 7421 3404
rect 12058 3413 12078 3433
rect 335 3166 355 3186
rect 431 3166 451 3186
rect 548 3166 568 3186
rect 644 3166 664 3186
rect 756 3166 776 3186
rect 852 3166 872 3186
rect 962 3166 982 3186
rect 4164 3200 4184 3220
rect 1058 3166 1078 3186
rect 4260 3200 4280 3220
rect 4370 3200 4390 3220
rect 4466 3200 4486 3220
rect 4578 3200 4598 3220
rect 4674 3200 4694 3220
rect 4791 3200 4811 3220
rect 12154 3413 12174 3433
rect 12271 3413 12291 3433
rect 12367 3413 12387 3433
rect 12479 3413 12499 3433
rect 12575 3413 12595 3433
rect 12685 3413 12705 3433
rect 12781 3413 12801 3433
rect 17339 3392 17359 3412
rect 17435 3392 17455 3412
rect 17552 3392 17572 3412
rect 17648 3392 17668 3412
rect 17760 3392 17780 3412
rect 17856 3392 17876 3412
rect 17966 3392 17986 3412
rect 18062 3392 18082 3412
rect 4887 3200 4907 3220
rect 5616 3145 5636 3165
rect 1347 2985 1367 3005
rect 1443 2985 1463 3005
rect 1560 2985 1580 3005
rect 1656 2985 1676 3005
rect 1768 2985 1788 3005
rect 1864 2985 1884 3005
rect 1974 2985 1994 3005
rect 5712 3145 5732 3165
rect 5829 3145 5849 3165
rect 5925 3145 5945 3165
rect 6037 3145 6057 3165
rect 6133 3145 6153 3165
rect 6243 3145 6263 3165
rect 9445 3179 9465 3199
rect 6339 3145 6359 3165
rect 9541 3179 9561 3199
rect 9651 3179 9671 3199
rect 9747 3179 9767 3199
rect 9859 3179 9879 3199
rect 9955 3179 9975 3199
rect 10072 3179 10092 3199
rect 10168 3179 10188 3199
rect 10996 3174 11016 3194
rect 2070 2985 2090 3005
rect 3151 2966 3171 2986
rect 3247 2966 3267 2986
rect 3357 2966 3377 2986
rect 3453 2966 3473 2986
rect 3565 2966 3585 2986
rect 3661 2966 3681 2986
rect 3778 2966 3798 2986
rect 11092 3174 11112 3194
rect 11209 3174 11229 3194
rect 11305 3174 11325 3194
rect 11417 3174 11437 3194
rect 11513 3174 11533 3194
rect 11623 3174 11643 3194
rect 14825 3208 14845 3228
rect 11719 3174 11739 3194
rect 14921 3208 14941 3228
rect 15031 3208 15051 3228
rect 15127 3208 15147 3228
rect 15239 3208 15259 3228
rect 15335 3208 15355 3228
rect 15452 3208 15472 3228
rect 15548 3208 15568 3228
rect 3874 2966 3894 2986
rect 6628 2964 6648 2984
rect 6724 2964 6744 2984
rect 6841 2964 6861 2984
rect 6937 2964 6957 2984
rect 7049 2964 7069 2984
rect 7145 2964 7165 2984
rect 7255 2964 7275 2984
rect 16277 3153 16297 3173
rect 7351 2964 7371 2984
rect 8432 2945 8452 2965
rect 334 2751 354 2771
rect 430 2751 450 2771
rect 547 2751 567 2771
rect 643 2751 663 2771
rect 755 2751 775 2771
rect 851 2751 871 2771
rect 961 2751 981 2771
rect 4163 2785 4183 2805
rect 1057 2751 1077 2771
rect 4259 2785 4279 2805
rect 4369 2785 4389 2805
rect 4465 2785 4485 2805
rect 4577 2785 4597 2805
rect 4673 2785 4693 2805
rect 4790 2785 4810 2805
rect 8528 2945 8548 2965
rect 8638 2945 8658 2965
rect 8734 2945 8754 2965
rect 8846 2945 8866 2965
rect 8942 2945 8962 2965
rect 9059 2945 9079 2965
rect 9155 2945 9175 2965
rect 12008 2993 12028 3013
rect 12104 2993 12124 3013
rect 12221 2993 12241 3013
rect 12317 2993 12337 3013
rect 12429 2993 12449 3013
rect 12525 2993 12545 3013
rect 12635 2993 12655 3013
rect 16373 3153 16393 3173
rect 16490 3153 16510 3173
rect 16586 3153 16606 3173
rect 16698 3153 16718 3173
rect 16794 3153 16814 3173
rect 16904 3153 16924 3173
rect 20106 3187 20126 3207
rect 17000 3153 17020 3173
rect 20202 3187 20222 3207
rect 20312 3187 20332 3207
rect 20408 3187 20428 3207
rect 20520 3187 20540 3207
rect 20616 3187 20636 3207
rect 20733 3187 20753 3207
rect 20829 3187 20849 3207
rect 12731 2993 12751 3013
rect 13812 2974 13832 2994
rect 4886 2785 4906 2805
rect 13908 2974 13928 2994
rect 14018 2974 14038 2994
rect 14114 2974 14134 2994
rect 14226 2974 14246 2994
rect 14322 2974 14342 2994
rect 14439 2974 14459 2994
rect 14535 2974 14555 2994
rect 17289 2972 17309 2992
rect 5615 2730 5635 2750
rect 5711 2730 5731 2750
rect 5828 2730 5848 2750
rect 5924 2730 5944 2750
rect 6036 2730 6056 2750
rect 6132 2730 6152 2750
rect 6242 2730 6262 2750
rect 9444 2764 9464 2784
rect 6338 2730 6358 2750
rect 9540 2764 9560 2784
rect 9650 2764 9670 2784
rect 9746 2764 9766 2784
rect 9858 2764 9878 2784
rect 9954 2764 9974 2784
rect 10071 2764 10091 2784
rect 17385 2972 17405 2992
rect 17502 2972 17522 2992
rect 17598 2972 17618 2992
rect 17710 2972 17730 2992
rect 17806 2972 17826 2992
rect 17916 2972 17936 2992
rect 18012 2972 18032 2992
rect 19093 2953 19113 2973
rect 10167 2764 10187 2784
rect 10995 2759 11015 2779
rect 11091 2759 11111 2779
rect 11208 2759 11228 2779
rect 11304 2759 11324 2779
rect 11416 2759 11436 2779
rect 11512 2759 11532 2779
rect 11622 2759 11642 2779
rect 14824 2793 14844 2813
rect 11718 2759 11738 2779
rect 14920 2793 14940 2813
rect 15030 2793 15050 2813
rect 15126 2793 15146 2813
rect 15238 2793 15258 2813
rect 15334 2793 15354 2813
rect 15451 2793 15471 2813
rect 19189 2953 19209 2973
rect 19299 2953 19319 2973
rect 19395 2953 19415 2973
rect 19507 2953 19527 2973
rect 19603 2953 19623 2973
rect 19720 2953 19740 2973
rect 19816 2953 19836 2973
rect 15547 2793 15567 2813
rect 16276 2738 16296 2758
rect 1562 2473 1582 2493
rect 1658 2473 1678 2493
rect 1775 2473 1795 2493
rect 1871 2473 1891 2493
rect 1983 2473 2003 2493
rect 2079 2473 2099 2493
rect 2189 2473 2209 2493
rect 2285 2473 2305 2493
rect 2943 2499 2963 2519
rect 3039 2499 3059 2519
rect 3149 2499 3169 2519
rect 3245 2499 3265 2519
rect 3357 2499 3377 2519
rect 3453 2499 3473 2519
rect 3570 2499 3590 2519
rect 16372 2738 16392 2758
rect 16489 2738 16509 2758
rect 16585 2738 16605 2758
rect 16697 2738 16717 2758
rect 16793 2738 16813 2758
rect 16903 2738 16923 2758
rect 20105 2772 20125 2792
rect 16999 2738 17019 2758
rect 20201 2772 20221 2792
rect 20311 2772 20331 2792
rect 20407 2772 20427 2792
rect 20519 2772 20539 2792
rect 20615 2772 20635 2792
rect 20732 2772 20752 2792
rect 20828 2772 20848 2792
rect 3666 2499 3686 2519
rect 6843 2452 6863 2472
rect 6939 2452 6959 2472
rect 7056 2452 7076 2472
rect 7152 2452 7172 2472
rect 7264 2452 7284 2472
rect 7360 2452 7380 2472
rect 7470 2452 7490 2472
rect 7566 2452 7586 2472
rect 8224 2478 8244 2498
rect 8320 2478 8340 2498
rect 8430 2478 8450 2498
rect 8526 2478 8546 2498
rect 8638 2478 8658 2498
rect 8734 2478 8754 2498
rect 8851 2478 8871 2498
rect 8947 2478 8967 2498
rect 12223 2481 12243 2501
rect 12319 2481 12339 2501
rect 12436 2481 12456 2501
rect 12532 2481 12552 2501
rect 12644 2481 12664 2501
rect 12740 2481 12760 2501
rect 12850 2481 12870 2501
rect 12946 2481 12966 2501
rect 13604 2507 13624 2527
rect 13700 2507 13720 2527
rect 13810 2507 13830 2527
rect 13906 2507 13926 2527
rect 14018 2507 14038 2527
rect 14114 2507 14134 2527
rect 14231 2507 14251 2527
rect 14327 2507 14347 2527
rect 17504 2460 17524 2480
rect 342 2187 362 2207
rect 438 2187 458 2207
rect 555 2187 575 2207
rect 651 2187 671 2207
rect 763 2187 783 2207
rect 859 2187 879 2207
rect 969 2187 989 2207
rect 4171 2221 4191 2241
rect 1065 2187 1085 2207
rect 4267 2221 4287 2241
rect 4377 2221 4397 2241
rect 4473 2221 4493 2241
rect 4585 2221 4605 2241
rect 4681 2221 4701 2241
rect 4798 2221 4818 2241
rect 17600 2460 17620 2480
rect 17717 2460 17737 2480
rect 17813 2460 17833 2480
rect 17925 2460 17945 2480
rect 18021 2460 18041 2480
rect 18131 2460 18151 2480
rect 18227 2460 18247 2480
rect 18885 2486 18905 2506
rect 18981 2486 19001 2506
rect 19091 2486 19111 2506
rect 19187 2486 19207 2506
rect 19299 2486 19319 2506
rect 19395 2486 19415 2506
rect 19512 2486 19532 2506
rect 19608 2486 19628 2506
rect 4894 2221 4914 2241
rect 5623 2166 5643 2186
rect 1354 2006 1374 2026
rect 1450 2006 1470 2026
rect 1567 2006 1587 2026
rect 1663 2006 1683 2026
rect 1775 2006 1795 2026
rect 1871 2006 1891 2026
rect 1981 2006 2001 2026
rect 5719 2166 5739 2186
rect 5836 2166 5856 2186
rect 5932 2166 5952 2186
rect 6044 2166 6064 2186
rect 6140 2166 6160 2186
rect 6250 2166 6270 2186
rect 9452 2200 9472 2220
rect 6346 2166 6366 2186
rect 9548 2200 9568 2220
rect 9658 2200 9678 2220
rect 9754 2200 9774 2220
rect 9866 2200 9886 2220
rect 9962 2200 9982 2220
rect 10079 2200 10099 2220
rect 10175 2200 10195 2220
rect 11003 2195 11023 2215
rect 2077 2006 2097 2026
rect 3158 1987 3178 2007
rect 3254 1987 3274 2007
rect 3364 1987 3384 2007
rect 3460 1987 3480 2007
rect 3572 1987 3592 2007
rect 3668 1987 3688 2007
rect 3785 1987 3805 2007
rect 11099 2195 11119 2215
rect 11216 2195 11236 2215
rect 11312 2195 11332 2215
rect 11424 2195 11444 2215
rect 11520 2195 11540 2215
rect 11630 2195 11650 2215
rect 14832 2229 14852 2249
rect 11726 2195 11746 2215
rect 14928 2229 14948 2249
rect 15038 2229 15058 2249
rect 15134 2229 15154 2249
rect 15246 2229 15266 2249
rect 15342 2229 15362 2249
rect 15459 2229 15479 2249
rect 15555 2229 15575 2249
rect 3881 1987 3901 2007
rect 6635 1985 6655 2005
rect 6731 1985 6751 2005
rect 6848 1985 6868 2005
rect 6944 1985 6964 2005
rect 7056 1985 7076 2005
rect 7152 1985 7172 2005
rect 7262 1985 7282 2005
rect 16284 2174 16304 2194
rect 7358 1985 7378 2005
rect 8439 1966 8459 1986
rect 341 1772 361 1792
rect 437 1772 457 1792
rect 554 1772 574 1792
rect 650 1772 670 1792
rect 762 1772 782 1792
rect 858 1772 878 1792
rect 968 1772 988 1792
rect 4170 1806 4190 1826
rect 1064 1772 1084 1792
rect 4266 1806 4286 1826
rect 4376 1806 4396 1826
rect 4472 1806 4492 1826
rect 4584 1806 4604 1826
rect 4680 1806 4700 1826
rect 4797 1806 4817 1826
rect 8535 1966 8555 1986
rect 8645 1966 8665 1986
rect 8741 1966 8761 1986
rect 8853 1966 8873 1986
rect 8949 1966 8969 1986
rect 9066 1966 9086 1986
rect 9162 1966 9182 1986
rect 12015 2014 12035 2034
rect 12111 2014 12131 2034
rect 12228 2014 12248 2034
rect 12324 2014 12344 2034
rect 12436 2014 12456 2034
rect 12532 2014 12552 2034
rect 12642 2014 12662 2034
rect 16380 2174 16400 2194
rect 16497 2174 16517 2194
rect 16593 2174 16613 2194
rect 16705 2174 16725 2194
rect 16801 2174 16821 2194
rect 16911 2174 16931 2194
rect 20113 2208 20133 2228
rect 17007 2174 17027 2194
rect 20209 2208 20229 2228
rect 20319 2208 20339 2228
rect 20415 2208 20435 2228
rect 20527 2208 20547 2228
rect 20623 2208 20643 2228
rect 20740 2208 20760 2228
rect 20836 2208 20856 2228
rect 12738 2014 12758 2034
rect 13819 1995 13839 2015
rect 4893 1806 4913 1826
rect 13915 1995 13935 2015
rect 14025 1995 14045 2015
rect 14121 1995 14141 2015
rect 14233 1995 14253 2015
rect 14329 1995 14349 2015
rect 14446 1995 14466 2015
rect 14542 1995 14562 2015
rect 17296 1993 17316 2013
rect 5622 1751 5642 1771
rect 5718 1751 5738 1771
rect 5835 1751 5855 1771
rect 5931 1751 5951 1771
rect 6043 1751 6063 1771
rect 6139 1751 6159 1771
rect 6249 1751 6269 1771
rect 9451 1785 9471 1805
rect 6345 1751 6365 1771
rect 9547 1785 9567 1805
rect 9657 1785 9677 1805
rect 9753 1785 9773 1805
rect 9865 1785 9885 1805
rect 9961 1785 9981 1805
rect 10078 1785 10098 1805
rect 17392 1993 17412 2013
rect 17509 1993 17529 2013
rect 17605 1993 17625 2013
rect 17717 1993 17737 2013
rect 17813 1993 17833 2013
rect 17923 1993 17943 2013
rect 18019 1993 18039 2013
rect 19100 1974 19120 1994
rect 10174 1785 10194 1805
rect 11002 1780 11022 1800
rect 11098 1780 11118 1800
rect 11215 1780 11235 1800
rect 11311 1780 11331 1800
rect 11423 1780 11443 1800
rect 11519 1780 11539 1800
rect 11629 1780 11649 1800
rect 14831 1814 14851 1834
rect 11725 1780 11745 1800
rect 14927 1814 14947 1834
rect 15037 1814 15057 1834
rect 15133 1814 15153 1834
rect 15245 1814 15265 1834
rect 15341 1814 15361 1834
rect 15458 1814 15478 1834
rect 19196 1974 19216 1994
rect 19306 1974 19326 1994
rect 19402 1974 19422 1994
rect 19514 1974 19534 1994
rect 19610 1974 19630 1994
rect 19727 1974 19747 1994
rect 19823 1974 19843 1994
rect 15554 1814 15574 1834
rect 16283 1759 16303 1779
rect 3108 1567 3128 1587
rect 3204 1567 3224 1587
rect 3314 1567 3334 1587
rect 3410 1567 3430 1587
rect 3522 1567 3542 1587
rect 3618 1567 3638 1587
rect 3735 1567 3755 1587
rect 3831 1567 3851 1587
rect 8389 1546 8409 1566
rect 8485 1546 8505 1566
rect 8595 1546 8615 1566
rect 8691 1546 8711 1566
rect 8803 1546 8823 1566
rect 8899 1546 8919 1566
rect 9016 1546 9036 1566
rect 16379 1759 16399 1779
rect 16496 1759 16516 1779
rect 16592 1759 16612 1779
rect 16704 1759 16724 1779
rect 16800 1759 16820 1779
rect 16910 1759 16930 1779
rect 20112 1793 20132 1813
rect 17006 1759 17026 1779
rect 20208 1793 20228 1813
rect 20318 1793 20338 1813
rect 20414 1793 20434 1813
rect 20526 1793 20546 1813
rect 20622 1793 20642 1813
rect 20739 1793 20759 1813
rect 20835 1793 20855 1813
rect 9112 1546 9132 1566
rect 13769 1575 13789 1595
rect 13865 1575 13885 1595
rect 13975 1575 13995 1595
rect 14071 1575 14091 1595
rect 14183 1575 14203 1595
rect 14279 1575 14299 1595
rect 14396 1575 14416 1595
rect 14492 1575 14512 1595
rect 19050 1554 19070 1574
rect 19146 1554 19166 1574
rect 19256 1554 19276 1574
rect 19352 1554 19372 1574
rect 19464 1554 19484 1574
rect 19560 1554 19580 1574
rect 19677 1554 19697 1574
rect 19773 1554 19793 1574
rect 1409 1445 1429 1465
rect 1505 1445 1525 1465
rect 1622 1445 1642 1465
rect 1718 1445 1738 1465
rect 1830 1445 1850 1465
rect 1926 1445 1946 1465
rect 2036 1445 2056 1465
rect 2132 1445 2152 1465
rect 6690 1424 6710 1444
rect 6786 1424 6806 1444
rect 6903 1424 6923 1444
rect 6999 1424 7019 1444
rect 7111 1424 7131 1444
rect 7207 1424 7227 1444
rect 7317 1424 7337 1444
rect 7413 1424 7433 1444
rect 12070 1453 12090 1473
rect 347 1206 367 1226
rect 443 1206 463 1226
rect 560 1206 580 1226
rect 656 1206 676 1226
rect 768 1206 788 1226
rect 864 1206 884 1226
rect 974 1206 994 1226
rect 4176 1240 4196 1260
rect 1070 1206 1090 1226
rect 4272 1240 4292 1260
rect 4382 1240 4402 1260
rect 4478 1240 4498 1260
rect 4590 1240 4610 1260
rect 4686 1240 4706 1260
rect 4803 1240 4823 1260
rect 12166 1453 12186 1473
rect 12283 1453 12303 1473
rect 12379 1453 12399 1473
rect 12491 1453 12511 1473
rect 12587 1453 12607 1473
rect 12697 1453 12717 1473
rect 12793 1453 12813 1473
rect 17351 1432 17371 1452
rect 17447 1432 17467 1452
rect 17564 1432 17584 1452
rect 17660 1432 17680 1452
rect 17772 1432 17792 1452
rect 17868 1432 17888 1452
rect 17978 1432 17998 1452
rect 18074 1432 18094 1452
rect 4899 1240 4919 1260
rect 5628 1185 5648 1205
rect 1359 1025 1379 1045
rect 1455 1025 1475 1045
rect 1572 1025 1592 1045
rect 1668 1025 1688 1045
rect 1780 1025 1800 1045
rect 1876 1025 1896 1045
rect 1986 1025 2006 1045
rect 5724 1185 5744 1205
rect 5841 1185 5861 1205
rect 5937 1185 5957 1205
rect 6049 1185 6069 1205
rect 6145 1185 6165 1205
rect 6255 1185 6275 1205
rect 9457 1219 9477 1239
rect 6351 1185 6371 1205
rect 9553 1219 9573 1239
rect 9663 1219 9683 1239
rect 9759 1219 9779 1239
rect 9871 1219 9891 1239
rect 9967 1219 9987 1239
rect 10084 1219 10104 1239
rect 10180 1219 10200 1239
rect 11008 1214 11028 1234
rect 2082 1025 2102 1045
rect 3163 1006 3183 1026
rect 3259 1006 3279 1026
rect 3369 1006 3389 1026
rect 3465 1006 3485 1026
rect 3577 1006 3597 1026
rect 3673 1006 3693 1026
rect 3790 1006 3810 1026
rect 11104 1214 11124 1234
rect 11221 1214 11241 1234
rect 11317 1214 11337 1234
rect 11429 1214 11449 1234
rect 11525 1214 11545 1234
rect 11635 1214 11655 1234
rect 14837 1248 14857 1268
rect 11731 1214 11751 1234
rect 14933 1248 14953 1268
rect 15043 1248 15063 1268
rect 15139 1248 15159 1268
rect 15251 1248 15271 1268
rect 15347 1248 15367 1268
rect 15464 1248 15484 1268
rect 15560 1248 15580 1268
rect 3886 1006 3906 1026
rect 6640 1004 6660 1024
rect 6736 1004 6756 1024
rect 6853 1004 6873 1024
rect 6949 1004 6969 1024
rect 7061 1004 7081 1024
rect 7157 1004 7177 1024
rect 7267 1004 7287 1024
rect 16289 1193 16309 1213
rect 7363 1004 7383 1024
rect 8444 985 8464 1005
rect 346 791 366 811
rect 442 791 462 811
rect 559 791 579 811
rect 655 791 675 811
rect 767 791 787 811
rect 863 791 883 811
rect 973 791 993 811
rect 4175 825 4195 845
rect 1069 791 1089 811
rect 4271 825 4291 845
rect 4381 825 4401 845
rect 4477 825 4497 845
rect 4589 825 4609 845
rect 4685 825 4705 845
rect 4802 825 4822 845
rect 8540 985 8560 1005
rect 8650 985 8670 1005
rect 8746 985 8766 1005
rect 8858 985 8878 1005
rect 8954 985 8974 1005
rect 9071 985 9091 1005
rect 9167 985 9187 1005
rect 12020 1033 12040 1053
rect 12116 1033 12136 1053
rect 12233 1033 12253 1053
rect 12329 1033 12349 1053
rect 12441 1033 12461 1053
rect 12537 1033 12557 1053
rect 12647 1033 12667 1053
rect 16385 1193 16405 1213
rect 16502 1193 16522 1213
rect 16598 1193 16618 1213
rect 16710 1193 16730 1213
rect 16806 1193 16826 1213
rect 16916 1193 16936 1213
rect 20118 1227 20138 1247
rect 17012 1193 17032 1213
rect 20214 1227 20234 1247
rect 20324 1227 20344 1247
rect 20420 1227 20440 1247
rect 20532 1227 20552 1247
rect 20628 1227 20648 1247
rect 20745 1227 20765 1247
rect 20841 1227 20861 1247
rect 12743 1033 12763 1053
rect 13824 1014 13844 1034
rect 4898 825 4918 845
rect 13920 1014 13940 1034
rect 14030 1014 14050 1034
rect 14126 1014 14146 1034
rect 14238 1014 14258 1034
rect 14334 1014 14354 1034
rect 14451 1014 14471 1034
rect 14547 1014 14567 1034
rect 17301 1012 17321 1032
rect 5627 770 5647 790
rect 5723 770 5743 790
rect 5840 770 5860 790
rect 5936 770 5956 790
rect 6048 770 6068 790
rect 6144 770 6164 790
rect 6254 770 6274 790
rect 9456 804 9476 824
rect 6350 770 6370 790
rect 9552 804 9572 824
rect 9662 804 9682 824
rect 9758 804 9778 824
rect 9870 804 9890 824
rect 9966 804 9986 824
rect 10083 804 10103 824
rect 17397 1012 17417 1032
rect 17514 1012 17534 1032
rect 17610 1012 17630 1032
rect 17722 1012 17742 1032
rect 17818 1012 17838 1032
rect 17928 1012 17948 1032
rect 18024 1012 18044 1032
rect 19105 993 19125 1013
rect 10179 804 10199 824
rect 11007 799 11027 819
rect 11103 799 11123 819
rect 11220 799 11240 819
rect 11316 799 11336 819
rect 11428 799 11448 819
rect 11524 799 11544 819
rect 11634 799 11654 819
rect 14836 833 14856 853
rect 11730 799 11750 819
rect 14932 833 14952 853
rect 15042 833 15062 853
rect 15138 833 15158 853
rect 15250 833 15270 853
rect 15346 833 15366 853
rect 15463 833 15483 853
rect 19201 993 19221 1013
rect 19311 993 19331 1013
rect 19407 993 19427 1013
rect 19519 993 19539 1013
rect 19615 993 19635 1013
rect 19732 993 19752 1013
rect 19828 993 19848 1013
rect 15559 833 15579 853
rect 16288 778 16308 798
rect 16384 778 16404 798
rect 16501 778 16521 798
rect 16597 778 16617 798
rect 16709 778 16729 798
rect 16805 778 16825 798
rect 16915 778 16935 798
rect 20117 812 20137 832
rect 17011 778 17031 798
rect 20213 812 20233 832
rect 20323 812 20343 832
rect 20419 812 20439 832
rect 20531 812 20551 832
rect 20627 812 20647 832
rect 20744 812 20764 832
rect 20840 812 20860 832
rect 1749 310 1769 330
rect 1845 310 1865 330
rect 1962 310 1982 330
rect 2058 310 2078 330
rect 2170 310 2190 330
rect 2266 310 2286 330
rect 2376 310 2396 330
rect 2472 310 2492 330
rect 7030 289 7050 309
rect 4839 222 4859 242
rect 4935 222 4955 242
rect 5052 222 5072 242
rect 5148 222 5168 242
rect 5260 222 5280 242
rect 5356 222 5376 242
rect 5466 222 5486 242
rect 7126 289 7146 309
rect 7243 289 7263 309
rect 7339 289 7359 309
rect 7451 289 7471 309
rect 7547 289 7567 309
rect 7657 289 7677 309
rect 12410 318 12430 338
rect 7753 289 7773 309
rect 12506 318 12526 338
rect 12623 318 12643 338
rect 12719 318 12739 338
rect 12831 318 12851 338
rect 12927 318 12947 338
rect 13037 318 13057 338
rect 13133 318 13153 338
rect 17691 297 17711 317
rect 5562 222 5582 242
rect 10100 215 10120 235
rect 10196 215 10216 235
rect 10313 215 10333 235
rect 10409 215 10429 235
rect 10521 215 10541 235
rect 10617 215 10637 235
rect 10727 215 10747 235
rect 10823 215 10843 235
rect 15500 230 15520 250
rect 15596 230 15616 250
rect 15713 230 15733 250
rect 15809 230 15829 250
rect 15921 230 15941 250
rect 16017 230 16037 250
rect 16127 230 16147 250
rect 17787 297 17807 317
rect 17904 297 17924 317
rect 18000 297 18020 317
rect 18112 297 18132 317
rect 18208 297 18228 317
rect 18318 297 18338 317
rect 18414 297 18434 317
rect 16223 230 16243 250
<< poly >>
rect 4171 8279 4221 8295
rect 4379 8279 4429 8295
rect 4587 8279 4637 8295
rect 4800 8279 4850 8295
rect 4171 8212 4221 8237
rect 4171 8186 4177 8212
rect 4203 8186 4221 8212
rect 4171 8160 4221 8186
rect 4379 8208 4429 8237
rect 4379 8184 4393 8208
rect 4417 8184 4429 8208
rect 4379 8160 4429 8184
rect 4587 8213 4637 8237
rect 4587 8189 4602 8213
rect 4626 8189 4637 8213
rect 4587 8160 4637 8189
rect 4800 8208 4850 8237
rect 14832 8287 14882 8303
rect 15040 8287 15090 8303
rect 15248 8287 15298 8303
rect 15461 8287 15511 8303
rect 9452 8258 9502 8274
rect 9660 8258 9710 8274
rect 9868 8258 9918 8274
rect 10081 8258 10131 8274
rect 4800 8188 4817 8208
rect 4837 8188 4850 8208
rect 4800 8160 4850 8188
rect 342 8122 392 8135
rect 555 8122 605 8135
rect 763 8122 813 8135
rect 971 8122 1021 8135
rect 3158 8045 3208 8061
rect 3366 8045 3416 8061
rect 3574 8045 3624 8061
rect 3787 8045 3837 8061
rect 9452 8191 9502 8216
rect 9452 8165 9458 8191
rect 9484 8165 9502 8191
rect 9452 8139 9502 8165
rect 9660 8187 9710 8216
rect 9660 8163 9674 8187
rect 9698 8163 9710 8187
rect 9660 8139 9710 8163
rect 9868 8192 9918 8216
rect 9868 8168 9883 8192
rect 9907 8168 9918 8192
rect 9868 8139 9918 8168
rect 10081 8187 10131 8216
rect 10081 8167 10098 8187
rect 10118 8167 10131 8187
rect 14832 8220 14882 8245
rect 14832 8194 14838 8220
rect 14864 8194 14882 8220
rect 14832 8168 14882 8194
rect 15040 8216 15090 8245
rect 15040 8192 15054 8216
rect 15078 8192 15090 8216
rect 15040 8168 15090 8192
rect 15248 8221 15298 8245
rect 15248 8197 15263 8221
rect 15287 8197 15298 8221
rect 15248 8168 15298 8197
rect 15461 8216 15511 8245
rect 20113 8266 20163 8282
rect 20321 8266 20371 8282
rect 20529 8266 20579 8282
rect 20742 8266 20792 8282
rect 15461 8196 15478 8216
rect 15498 8196 15511 8216
rect 15461 8168 15511 8196
rect 10081 8139 10131 8167
rect 5623 8101 5673 8114
rect 5836 8101 5886 8114
rect 6044 8101 6094 8114
rect 6252 8101 6302 8114
rect 4171 8047 4221 8060
rect 4379 8047 4429 8060
rect 4587 8047 4637 8060
rect 4800 8047 4850 8060
rect 342 7994 392 8022
rect 342 7974 355 7994
rect 375 7974 392 7994
rect 342 7945 392 7974
rect 555 7993 605 8022
rect 555 7969 566 7993
rect 590 7969 605 7993
rect 555 7945 605 7969
rect 763 7998 813 8022
rect 763 7974 775 7998
rect 799 7974 813 7998
rect 763 7945 813 7974
rect 971 7996 1021 8022
rect 971 7970 989 7996
rect 1015 7970 1021 7996
rect 971 7945 1021 7970
rect 3158 7978 3208 8003
rect 1354 7941 1404 7954
rect 1567 7941 1617 7954
rect 1775 7941 1825 7954
rect 1983 7941 2033 7954
rect 3158 7952 3164 7978
rect 3190 7952 3208 7978
rect 342 7887 392 7903
rect 555 7887 605 7903
rect 763 7887 813 7903
rect 971 7887 1021 7903
rect 3158 7926 3208 7952
rect 3366 7974 3416 8003
rect 3366 7950 3380 7974
rect 3404 7950 3416 7974
rect 3366 7926 3416 7950
rect 3574 7979 3624 8003
rect 3574 7955 3589 7979
rect 3613 7955 3624 7979
rect 3574 7926 3624 7955
rect 3787 7974 3837 8003
rect 3787 7954 3804 7974
rect 3824 7954 3837 7974
rect 3787 7926 3837 7954
rect 8439 8024 8489 8040
rect 8647 8024 8697 8040
rect 8855 8024 8905 8040
rect 9068 8024 9118 8040
rect 11003 8130 11053 8143
rect 11216 8130 11266 8143
rect 11424 8130 11474 8143
rect 11632 8130 11682 8143
rect 9452 8026 9502 8039
rect 9660 8026 9710 8039
rect 9868 8026 9918 8039
rect 10081 8026 10131 8039
rect 5623 7973 5673 8001
rect 5623 7953 5636 7973
rect 5656 7953 5673 7973
rect 1354 7813 1404 7841
rect 1354 7793 1367 7813
rect 1387 7793 1404 7813
rect 1354 7764 1404 7793
rect 1567 7812 1617 7841
rect 1567 7788 1578 7812
rect 1602 7788 1617 7812
rect 1567 7764 1617 7788
rect 1775 7817 1825 7841
rect 1775 7793 1787 7817
rect 1811 7793 1825 7817
rect 1775 7764 1825 7793
rect 1983 7815 2033 7841
rect 5623 7924 5673 7953
rect 5836 7972 5886 8001
rect 5836 7948 5847 7972
rect 5871 7948 5886 7972
rect 5836 7924 5886 7948
rect 6044 7977 6094 8001
rect 6044 7953 6056 7977
rect 6080 7953 6094 7977
rect 6044 7924 6094 7953
rect 6252 7975 6302 8001
rect 13819 8053 13869 8069
rect 14027 8053 14077 8069
rect 14235 8053 14285 8069
rect 14448 8053 14498 8069
rect 20113 8199 20163 8224
rect 20113 8173 20119 8199
rect 20145 8173 20163 8199
rect 20113 8147 20163 8173
rect 20321 8195 20371 8224
rect 20321 8171 20335 8195
rect 20359 8171 20371 8195
rect 20321 8147 20371 8171
rect 20529 8200 20579 8224
rect 20529 8176 20544 8200
rect 20568 8176 20579 8200
rect 20529 8147 20579 8176
rect 20742 8195 20792 8224
rect 20742 8175 20759 8195
rect 20779 8175 20792 8195
rect 20742 8147 20792 8175
rect 16284 8109 16334 8122
rect 16497 8109 16547 8122
rect 16705 8109 16755 8122
rect 16913 8109 16963 8122
rect 14832 8055 14882 8068
rect 15040 8055 15090 8068
rect 15248 8055 15298 8068
rect 15461 8055 15511 8068
rect 6252 7949 6270 7975
rect 6296 7949 6302 7975
rect 6252 7924 6302 7949
rect 8439 7957 8489 7982
rect 6635 7920 6685 7933
rect 6848 7920 6898 7933
rect 7056 7920 7106 7933
rect 7264 7920 7314 7933
rect 8439 7931 8445 7957
rect 8471 7931 8489 7957
rect 4170 7864 4220 7880
rect 4378 7864 4428 7880
rect 4586 7864 4636 7880
rect 4799 7864 4849 7880
rect 5623 7866 5673 7882
rect 5836 7866 5886 7882
rect 6044 7866 6094 7882
rect 6252 7866 6302 7882
rect 1983 7789 2001 7815
rect 2027 7789 2033 7815
rect 3158 7813 3208 7826
rect 3366 7813 3416 7826
rect 3574 7813 3624 7826
rect 3787 7813 3837 7826
rect 1983 7764 2033 7789
rect 4170 7797 4220 7822
rect 4170 7771 4176 7797
rect 4202 7771 4220 7797
rect 4170 7745 4220 7771
rect 4378 7793 4428 7822
rect 4378 7769 4392 7793
rect 4416 7769 4428 7793
rect 4378 7745 4428 7769
rect 4586 7798 4636 7822
rect 4586 7774 4601 7798
rect 4625 7774 4636 7798
rect 4586 7745 4636 7774
rect 4799 7793 4849 7822
rect 8439 7905 8489 7931
rect 8647 7953 8697 7982
rect 8647 7929 8661 7953
rect 8685 7929 8697 7953
rect 8647 7905 8697 7929
rect 8855 7958 8905 7982
rect 8855 7934 8870 7958
rect 8894 7934 8905 7958
rect 8855 7905 8905 7934
rect 9068 7953 9118 7982
rect 11003 8002 11053 8030
rect 11003 7982 11016 8002
rect 11036 7982 11053 8002
rect 9068 7933 9085 7953
rect 9105 7933 9118 7953
rect 9068 7905 9118 7933
rect 11003 7953 11053 7982
rect 11216 8001 11266 8030
rect 11216 7977 11227 8001
rect 11251 7977 11266 8001
rect 11216 7953 11266 7977
rect 11424 8006 11474 8030
rect 11424 7982 11436 8006
rect 11460 7982 11474 8006
rect 11424 7953 11474 7982
rect 11632 8004 11682 8030
rect 11632 7978 11650 8004
rect 11676 7978 11682 8004
rect 11632 7953 11682 7978
rect 13819 7986 13869 8011
rect 12015 7949 12065 7962
rect 12228 7949 12278 7962
rect 12436 7949 12486 7962
rect 12644 7949 12694 7962
rect 13819 7960 13825 7986
rect 13851 7960 13869 7986
rect 4799 7773 4816 7793
rect 4836 7773 4849 7793
rect 4799 7745 4849 7773
rect 341 7707 391 7720
rect 554 7707 604 7720
rect 762 7707 812 7720
rect 970 7707 1020 7720
rect 1354 7706 1404 7722
rect 1567 7706 1617 7722
rect 1775 7706 1825 7722
rect 1983 7706 2033 7722
rect 6635 7792 6685 7820
rect 6635 7772 6648 7792
rect 6668 7772 6685 7792
rect 6635 7743 6685 7772
rect 6848 7791 6898 7820
rect 6848 7767 6859 7791
rect 6883 7767 6898 7791
rect 6848 7743 6898 7767
rect 7056 7796 7106 7820
rect 7056 7772 7068 7796
rect 7092 7772 7106 7796
rect 7056 7743 7106 7772
rect 7264 7794 7314 7820
rect 11003 7895 11053 7911
rect 11216 7895 11266 7911
rect 11424 7895 11474 7911
rect 11632 7895 11682 7911
rect 9451 7843 9501 7859
rect 9659 7843 9709 7859
rect 9867 7843 9917 7859
rect 10080 7843 10130 7859
rect 13819 7934 13869 7960
rect 14027 7982 14077 8011
rect 14027 7958 14041 7982
rect 14065 7958 14077 7982
rect 14027 7934 14077 7958
rect 14235 7987 14285 8011
rect 14235 7963 14250 7987
rect 14274 7963 14285 7987
rect 14235 7934 14285 7963
rect 14448 7982 14498 8011
rect 14448 7962 14465 7982
rect 14485 7962 14498 7982
rect 14448 7934 14498 7962
rect 19100 8032 19150 8048
rect 19308 8032 19358 8048
rect 19516 8032 19566 8048
rect 19729 8032 19779 8048
rect 20113 8034 20163 8047
rect 20321 8034 20371 8047
rect 20529 8034 20579 8047
rect 20742 8034 20792 8047
rect 16284 7981 16334 8009
rect 16284 7961 16297 7981
rect 16317 7961 16334 7981
rect 7264 7768 7282 7794
rect 7308 7768 7314 7794
rect 8439 7792 8489 7805
rect 8647 7792 8697 7805
rect 8855 7792 8905 7805
rect 9068 7792 9118 7805
rect 7264 7743 7314 7768
rect 9451 7776 9501 7801
rect 9451 7750 9457 7776
rect 9483 7750 9501 7776
rect 9451 7724 9501 7750
rect 9659 7772 9709 7801
rect 9659 7748 9673 7772
rect 9697 7748 9709 7772
rect 9659 7724 9709 7748
rect 9867 7777 9917 7801
rect 9867 7753 9882 7777
rect 9906 7753 9917 7777
rect 9867 7724 9917 7753
rect 10080 7772 10130 7801
rect 12015 7821 12065 7849
rect 12015 7801 12028 7821
rect 12048 7801 12065 7821
rect 10080 7752 10097 7772
rect 10117 7752 10130 7772
rect 10080 7724 10130 7752
rect 12015 7772 12065 7801
rect 12228 7820 12278 7849
rect 12228 7796 12239 7820
rect 12263 7796 12278 7820
rect 12228 7772 12278 7796
rect 12436 7825 12486 7849
rect 12436 7801 12448 7825
rect 12472 7801 12486 7825
rect 12436 7772 12486 7801
rect 12644 7823 12694 7849
rect 16284 7932 16334 7961
rect 16497 7980 16547 8009
rect 16497 7956 16508 7980
rect 16532 7956 16547 7980
rect 16497 7932 16547 7956
rect 16705 7985 16755 8009
rect 16705 7961 16717 7985
rect 16741 7961 16755 7985
rect 16705 7932 16755 7961
rect 16913 7983 16963 8009
rect 16913 7957 16931 7983
rect 16957 7957 16963 7983
rect 16913 7932 16963 7957
rect 19100 7965 19150 7990
rect 17296 7928 17346 7941
rect 17509 7928 17559 7941
rect 17717 7928 17767 7941
rect 17925 7928 17975 7941
rect 19100 7939 19106 7965
rect 19132 7939 19150 7965
rect 14831 7872 14881 7888
rect 15039 7872 15089 7888
rect 15247 7872 15297 7888
rect 15460 7872 15510 7888
rect 16284 7874 16334 7890
rect 16497 7874 16547 7890
rect 16705 7874 16755 7890
rect 16913 7874 16963 7890
rect 12644 7797 12662 7823
rect 12688 7797 12694 7823
rect 13819 7821 13869 7834
rect 14027 7821 14077 7834
rect 14235 7821 14285 7834
rect 14448 7821 14498 7834
rect 12644 7772 12694 7797
rect 14831 7805 14881 7830
rect 14831 7779 14837 7805
rect 14863 7779 14881 7805
rect 5622 7686 5672 7699
rect 5835 7686 5885 7699
rect 6043 7686 6093 7699
rect 6251 7686 6301 7699
rect 3108 7625 3158 7641
rect 3316 7625 3366 7641
rect 3524 7625 3574 7641
rect 3737 7625 3787 7641
rect 4170 7632 4220 7645
rect 4378 7632 4428 7645
rect 4586 7632 4636 7645
rect 4799 7632 4849 7645
rect 341 7579 391 7607
rect 341 7559 354 7579
rect 374 7559 391 7579
rect 341 7530 391 7559
rect 554 7578 604 7607
rect 554 7554 565 7578
rect 589 7554 604 7578
rect 554 7530 604 7554
rect 762 7583 812 7607
rect 762 7559 774 7583
rect 798 7559 812 7583
rect 762 7530 812 7559
rect 970 7581 1020 7607
rect 970 7555 988 7581
rect 1014 7555 1020 7581
rect 970 7530 1020 7555
rect 3108 7558 3158 7583
rect 3108 7532 3114 7558
rect 3140 7532 3158 7558
rect 3108 7506 3158 7532
rect 3316 7554 3366 7583
rect 3316 7530 3330 7554
rect 3354 7530 3366 7554
rect 3316 7506 3366 7530
rect 3524 7559 3574 7583
rect 3524 7535 3539 7559
rect 3563 7535 3574 7559
rect 3524 7506 3574 7535
rect 3737 7554 3787 7583
rect 3737 7534 3754 7554
rect 3774 7534 3787 7554
rect 3737 7506 3787 7534
rect 6635 7685 6685 7701
rect 6848 7685 6898 7701
rect 7056 7685 7106 7701
rect 7264 7685 7314 7701
rect 14831 7753 14881 7779
rect 15039 7801 15089 7830
rect 15039 7777 15053 7801
rect 15077 7777 15089 7801
rect 15039 7753 15089 7777
rect 15247 7806 15297 7830
rect 15247 7782 15262 7806
rect 15286 7782 15297 7806
rect 15247 7753 15297 7782
rect 15460 7801 15510 7830
rect 19100 7913 19150 7939
rect 19308 7961 19358 7990
rect 19308 7937 19322 7961
rect 19346 7937 19358 7961
rect 19308 7913 19358 7937
rect 19516 7966 19566 7990
rect 19516 7942 19531 7966
rect 19555 7942 19566 7966
rect 19516 7913 19566 7942
rect 19729 7961 19779 7990
rect 19729 7941 19746 7961
rect 19766 7941 19779 7961
rect 19729 7913 19779 7941
rect 15460 7781 15477 7801
rect 15497 7781 15510 7801
rect 15460 7753 15510 7781
rect 11002 7715 11052 7728
rect 11215 7715 11265 7728
rect 11423 7715 11473 7728
rect 11631 7715 11681 7728
rect 8389 7604 8439 7620
rect 8597 7604 8647 7620
rect 8805 7604 8855 7620
rect 9018 7604 9068 7620
rect 9451 7611 9501 7624
rect 9659 7611 9709 7624
rect 9867 7611 9917 7624
rect 10080 7611 10130 7624
rect 12015 7714 12065 7730
rect 12228 7714 12278 7730
rect 12436 7714 12486 7730
rect 12644 7714 12694 7730
rect 17296 7800 17346 7828
rect 17296 7780 17309 7800
rect 17329 7780 17346 7800
rect 17296 7751 17346 7780
rect 17509 7799 17559 7828
rect 17509 7775 17520 7799
rect 17544 7775 17559 7799
rect 17509 7751 17559 7775
rect 17717 7804 17767 7828
rect 17717 7780 17729 7804
rect 17753 7780 17767 7804
rect 17717 7751 17767 7780
rect 17925 7802 17975 7828
rect 20112 7851 20162 7867
rect 20320 7851 20370 7867
rect 20528 7851 20578 7867
rect 20741 7851 20791 7867
rect 17925 7776 17943 7802
rect 17969 7776 17975 7802
rect 19100 7800 19150 7813
rect 19308 7800 19358 7813
rect 19516 7800 19566 7813
rect 19729 7800 19779 7813
rect 17925 7751 17975 7776
rect 20112 7784 20162 7809
rect 20112 7758 20118 7784
rect 20144 7758 20162 7784
rect 20112 7732 20162 7758
rect 20320 7780 20370 7809
rect 20320 7756 20334 7780
rect 20358 7756 20370 7780
rect 20320 7732 20370 7756
rect 20528 7785 20578 7809
rect 20528 7761 20543 7785
rect 20567 7761 20578 7785
rect 20528 7732 20578 7761
rect 20741 7780 20791 7809
rect 20741 7760 20758 7780
rect 20778 7760 20791 7780
rect 20741 7732 20791 7760
rect 16283 7694 16333 7707
rect 16496 7694 16546 7707
rect 16704 7694 16754 7707
rect 16912 7694 16962 7707
rect 13769 7633 13819 7649
rect 13977 7633 14027 7649
rect 14185 7633 14235 7649
rect 14398 7633 14448 7649
rect 14831 7640 14881 7653
rect 15039 7640 15089 7653
rect 15247 7640 15297 7653
rect 15460 7640 15510 7653
rect 5622 7558 5672 7586
rect 341 7472 391 7488
rect 554 7472 604 7488
rect 762 7472 812 7488
rect 970 7472 1020 7488
rect 5622 7538 5635 7558
rect 5655 7538 5672 7558
rect 5622 7509 5672 7538
rect 5835 7557 5885 7586
rect 5835 7533 5846 7557
rect 5870 7533 5885 7557
rect 5835 7509 5885 7533
rect 6043 7562 6093 7586
rect 6043 7538 6055 7562
rect 6079 7538 6093 7562
rect 6043 7509 6093 7538
rect 6251 7560 6301 7586
rect 11002 7587 11052 7615
rect 6251 7534 6269 7560
rect 6295 7534 6301 7560
rect 6251 7509 6301 7534
rect 8389 7537 8439 7562
rect 8389 7511 8395 7537
rect 8421 7511 8439 7537
rect 8389 7485 8439 7511
rect 8597 7533 8647 7562
rect 8597 7509 8611 7533
rect 8635 7509 8647 7533
rect 8597 7485 8647 7509
rect 8805 7538 8855 7562
rect 8805 7514 8820 7538
rect 8844 7514 8855 7538
rect 8805 7485 8855 7514
rect 9018 7533 9068 7562
rect 9018 7513 9035 7533
rect 9055 7513 9068 7533
rect 9018 7485 9068 7513
rect 11002 7567 11015 7587
rect 11035 7567 11052 7587
rect 11002 7538 11052 7567
rect 11215 7586 11265 7615
rect 11215 7562 11226 7586
rect 11250 7562 11265 7586
rect 11215 7538 11265 7562
rect 11423 7591 11473 7615
rect 11423 7567 11435 7591
rect 11459 7567 11473 7591
rect 11423 7538 11473 7567
rect 11631 7589 11681 7615
rect 11631 7563 11649 7589
rect 11675 7563 11681 7589
rect 11631 7538 11681 7563
rect 13769 7566 13819 7591
rect 13769 7540 13775 7566
rect 13801 7540 13819 7566
rect 5622 7451 5672 7467
rect 5835 7451 5885 7467
rect 6043 7451 6093 7467
rect 6251 7451 6301 7467
rect 3108 7393 3158 7406
rect 3316 7393 3366 7406
rect 3524 7393 3574 7406
rect 3737 7393 3787 7406
rect 1409 7380 1459 7393
rect 1622 7380 1672 7393
rect 1830 7380 1880 7393
rect 2038 7380 2088 7393
rect 13769 7514 13819 7540
rect 13977 7562 14027 7591
rect 13977 7538 13991 7562
rect 14015 7538 14027 7562
rect 13977 7514 14027 7538
rect 14185 7567 14235 7591
rect 14185 7543 14200 7567
rect 14224 7543 14235 7567
rect 14185 7514 14235 7543
rect 14398 7562 14448 7591
rect 14398 7542 14415 7562
rect 14435 7542 14448 7562
rect 14398 7514 14448 7542
rect 17296 7693 17346 7709
rect 17509 7693 17559 7709
rect 17717 7693 17767 7709
rect 17925 7693 17975 7709
rect 19050 7612 19100 7628
rect 19258 7612 19308 7628
rect 19466 7612 19516 7628
rect 19679 7612 19729 7628
rect 20112 7619 20162 7632
rect 20320 7619 20370 7632
rect 20528 7619 20578 7632
rect 20741 7619 20791 7632
rect 16283 7566 16333 7594
rect 11002 7480 11052 7496
rect 11215 7480 11265 7496
rect 11423 7480 11473 7496
rect 11631 7480 11681 7496
rect 16283 7546 16296 7566
rect 16316 7546 16333 7566
rect 16283 7517 16333 7546
rect 16496 7565 16546 7594
rect 16496 7541 16507 7565
rect 16531 7541 16546 7565
rect 16496 7517 16546 7541
rect 16704 7570 16754 7594
rect 16704 7546 16716 7570
rect 16740 7546 16754 7570
rect 16704 7517 16754 7546
rect 16912 7568 16962 7594
rect 16912 7542 16930 7568
rect 16956 7542 16962 7568
rect 16912 7517 16962 7542
rect 19050 7545 19100 7570
rect 19050 7519 19056 7545
rect 19082 7519 19100 7545
rect 19050 7493 19100 7519
rect 19258 7541 19308 7570
rect 19258 7517 19272 7541
rect 19296 7517 19308 7541
rect 19258 7493 19308 7517
rect 19466 7546 19516 7570
rect 19466 7522 19481 7546
rect 19505 7522 19516 7546
rect 19466 7493 19516 7522
rect 19679 7541 19729 7570
rect 19679 7521 19696 7541
rect 19716 7521 19729 7541
rect 19679 7493 19729 7521
rect 16283 7459 16333 7475
rect 16496 7459 16546 7475
rect 16704 7459 16754 7475
rect 16912 7459 16962 7475
rect 13769 7401 13819 7414
rect 13977 7401 14027 7414
rect 14185 7401 14235 7414
rect 14398 7401 14448 7414
rect 12070 7388 12120 7401
rect 12283 7388 12333 7401
rect 12491 7388 12541 7401
rect 12699 7388 12749 7401
rect 8389 7372 8439 7385
rect 8597 7372 8647 7385
rect 8805 7372 8855 7385
rect 9018 7372 9068 7385
rect 6690 7359 6740 7372
rect 6903 7359 6953 7372
rect 7111 7359 7161 7372
rect 7319 7359 7369 7372
rect 4176 7298 4226 7314
rect 4384 7298 4434 7314
rect 4592 7298 4642 7314
rect 4805 7298 4855 7314
rect 1409 7252 1459 7280
rect 1409 7232 1422 7252
rect 1442 7232 1459 7252
rect 1409 7203 1459 7232
rect 1622 7251 1672 7280
rect 1622 7227 1633 7251
rect 1657 7227 1672 7251
rect 1622 7203 1672 7227
rect 1830 7256 1880 7280
rect 1830 7232 1842 7256
rect 1866 7232 1880 7256
rect 1830 7203 1880 7232
rect 2038 7254 2088 7280
rect 2038 7228 2056 7254
rect 2082 7228 2088 7254
rect 2038 7203 2088 7228
rect 4176 7231 4226 7256
rect 4176 7205 4182 7231
rect 4208 7205 4226 7231
rect 4176 7179 4226 7205
rect 4384 7227 4434 7256
rect 4384 7203 4398 7227
rect 4422 7203 4434 7227
rect 4384 7179 4434 7203
rect 4592 7232 4642 7256
rect 4592 7208 4607 7232
rect 4631 7208 4642 7232
rect 4592 7179 4642 7208
rect 4805 7227 4855 7256
rect 4805 7207 4822 7227
rect 4842 7207 4855 7227
rect 9457 7277 9507 7293
rect 9665 7277 9715 7293
rect 9873 7277 9923 7293
rect 10086 7277 10136 7293
rect 4805 7179 4855 7207
rect 347 7141 397 7154
rect 560 7141 610 7154
rect 768 7141 818 7154
rect 976 7141 1026 7154
rect 1409 7145 1459 7161
rect 1622 7145 1672 7161
rect 1830 7145 1880 7161
rect 2038 7145 2088 7161
rect 3163 7064 3213 7080
rect 3371 7064 3421 7080
rect 3579 7064 3629 7080
rect 3792 7064 3842 7080
rect 6690 7231 6740 7259
rect 6690 7211 6703 7231
rect 6723 7211 6740 7231
rect 6690 7182 6740 7211
rect 6903 7230 6953 7259
rect 6903 7206 6914 7230
rect 6938 7206 6953 7230
rect 6903 7182 6953 7206
rect 7111 7235 7161 7259
rect 7111 7211 7123 7235
rect 7147 7211 7161 7235
rect 7111 7182 7161 7211
rect 7319 7233 7369 7259
rect 19050 7380 19100 7393
rect 19258 7380 19308 7393
rect 19466 7380 19516 7393
rect 19679 7380 19729 7393
rect 17351 7367 17401 7380
rect 17564 7367 17614 7380
rect 17772 7367 17822 7380
rect 17980 7367 18030 7380
rect 14837 7306 14887 7322
rect 15045 7306 15095 7322
rect 15253 7306 15303 7322
rect 15466 7306 15516 7322
rect 7319 7207 7337 7233
rect 7363 7207 7369 7233
rect 7319 7182 7369 7207
rect 9457 7210 9507 7235
rect 9457 7184 9463 7210
rect 9489 7184 9507 7210
rect 9457 7158 9507 7184
rect 9665 7206 9715 7235
rect 9665 7182 9679 7206
rect 9703 7182 9715 7206
rect 9665 7158 9715 7182
rect 9873 7211 9923 7235
rect 9873 7187 9888 7211
rect 9912 7187 9923 7211
rect 9873 7158 9923 7187
rect 10086 7206 10136 7235
rect 10086 7186 10103 7206
rect 10123 7186 10136 7206
rect 12070 7260 12120 7288
rect 12070 7240 12083 7260
rect 12103 7240 12120 7260
rect 12070 7211 12120 7240
rect 12283 7259 12333 7288
rect 12283 7235 12294 7259
rect 12318 7235 12333 7259
rect 12283 7211 12333 7235
rect 12491 7264 12541 7288
rect 12491 7240 12503 7264
rect 12527 7240 12541 7264
rect 12491 7211 12541 7240
rect 12699 7262 12749 7288
rect 12699 7236 12717 7262
rect 12743 7236 12749 7262
rect 12699 7211 12749 7236
rect 14837 7239 14887 7264
rect 14837 7213 14843 7239
rect 14869 7213 14887 7239
rect 10086 7158 10136 7186
rect 14837 7187 14887 7213
rect 15045 7235 15095 7264
rect 15045 7211 15059 7235
rect 15083 7211 15095 7235
rect 15045 7187 15095 7211
rect 15253 7240 15303 7264
rect 15253 7216 15268 7240
rect 15292 7216 15303 7240
rect 15253 7187 15303 7216
rect 15466 7235 15516 7264
rect 15466 7215 15483 7235
rect 15503 7215 15516 7235
rect 20118 7285 20168 7301
rect 20326 7285 20376 7301
rect 20534 7285 20584 7301
rect 20747 7285 20797 7301
rect 15466 7187 15516 7215
rect 5628 7120 5678 7133
rect 5841 7120 5891 7133
rect 6049 7120 6099 7133
rect 6257 7120 6307 7133
rect 6690 7124 6740 7140
rect 6903 7124 6953 7140
rect 7111 7124 7161 7140
rect 7319 7124 7369 7140
rect 4176 7066 4226 7079
rect 4384 7066 4434 7079
rect 4592 7066 4642 7079
rect 4805 7066 4855 7079
rect 347 7013 397 7041
rect 347 6993 360 7013
rect 380 6993 397 7013
rect 347 6964 397 6993
rect 560 7012 610 7041
rect 560 6988 571 7012
rect 595 6988 610 7012
rect 560 6964 610 6988
rect 768 7017 818 7041
rect 768 6993 780 7017
rect 804 6993 818 7017
rect 768 6964 818 6993
rect 976 7015 1026 7041
rect 976 6989 994 7015
rect 1020 6989 1026 7015
rect 976 6964 1026 6989
rect 3163 6997 3213 7022
rect 1359 6960 1409 6973
rect 1572 6960 1622 6973
rect 1780 6960 1830 6973
rect 1988 6960 2038 6973
rect 3163 6971 3169 6997
rect 3195 6971 3213 6997
rect 347 6906 397 6922
rect 560 6906 610 6922
rect 768 6906 818 6922
rect 976 6906 1026 6922
rect 3163 6945 3213 6971
rect 3371 6993 3421 7022
rect 3371 6969 3385 6993
rect 3409 6969 3421 6993
rect 3371 6945 3421 6969
rect 3579 6998 3629 7022
rect 3579 6974 3594 6998
rect 3618 6974 3629 6998
rect 3579 6945 3629 6974
rect 3792 6993 3842 7022
rect 3792 6973 3809 6993
rect 3829 6973 3842 6993
rect 3792 6945 3842 6973
rect 8444 7043 8494 7059
rect 8652 7043 8702 7059
rect 8860 7043 8910 7059
rect 9073 7043 9123 7059
rect 11008 7149 11058 7162
rect 11221 7149 11271 7162
rect 11429 7149 11479 7162
rect 11637 7149 11687 7162
rect 12070 7153 12120 7169
rect 12283 7153 12333 7169
rect 12491 7153 12541 7169
rect 12699 7153 12749 7169
rect 9457 7045 9507 7058
rect 9665 7045 9715 7058
rect 9873 7045 9923 7058
rect 10086 7045 10136 7058
rect 5628 6992 5678 7020
rect 5628 6972 5641 6992
rect 5661 6972 5678 6992
rect 1359 6832 1409 6860
rect 1359 6812 1372 6832
rect 1392 6812 1409 6832
rect 1359 6783 1409 6812
rect 1572 6831 1622 6860
rect 1572 6807 1583 6831
rect 1607 6807 1622 6831
rect 1572 6783 1622 6807
rect 1780 6836 1830 6860
rect 1780 6812 1792 6836
rect 1816 6812 1830 6836
rect 1780 6783 1830 6812
rect 1988 6834 2038 6860
rect 5628 6943 5678 6972
rect 5841 6991 5891 7020
rect 5841 6967 5852 6991
rect 5876 6967 5891 6991
rect 5841 6943 5891 6967
rect 6049 6996 6099 7020
rect 6049 6972 6061 6996
rect 6085 6972 6099 6996
rect 6049 6943 6099 6972
rect 6257 6994 6307 7020
rect 13824 7072 13874 7088
rect 14032 7072 14082 7088
rect 14240 7072 14290 7088
rect 14453 7072 14503 7088
rect 17351 7239 17401 7267
rect 17351 7219 17364 7239
rect 17384 7219 17401 7239
rect 17351 7190 17401 7219
rect 17564 7238 17614 7267
rect 17564 7214 17575 7238
rect 17599 7214 17614 7238
rect 17564 7190 17614 7214
rect 17772 7243 17822 7267
rect 17772 7219 17784 7243
rect 17808 7219 17822 7243
rect 17772 7190 17822 7219
rect 17980 7241 18030 7267
rect 17980 7215 17998 7241
rect 18024 7215 18030 7241
rect 17980 7190 18030 7215
rect 20118 7218 20168 7243
rect 20118 7192 20124 7218
rect 20150 7192 20168 7218
rect 20118 7166 20168 7192
rect 20326 7214 20376 7243
rect 20326 7190 20340 7214
rect 20364 7190 20376 7214
rect 20326 7166 20376 7190
rect 20534 7219 20584 7243
rect 20534 7195 20549 7219
rect 20573 7195 20584 7219
rect 20534 7166 20584 7195
rect 20747 7214 20797 7243
rect 20747 7194 20764 7214
rect 20784 7194 20797 7214
rect 20747 7166 20797 7194
rect 16289 7128 16339 7141
rect 16502 7128 16552 7141
rect 16710 7128 16760 7141
rect 16918 7128 16968 7141
rect 17351 7132 17401 7148
rect 17564 7132 17614 7148
rect 17772 7132 17822 7148
rect 17980 7132 18030 7148
rect 14837 7074 14887 7087
rect 15045 7074 15095 7087
rect 15253 7074 15303 7087
rect 15466 7074 15516 7087
rect 6257 6968 6275 6994
rect 6301 6968 6307 6994
rect 6257 6943 6307 6968
rect 8444 6976 8494 7001
rect 6640 6939 6690 6952
rect 6853 6939 6903 6952
rect 7061 6939 7111 6952
rect 7269 6939 7319 6952
rect 8444 6950 8450 6976
rect 8476 6950 8494 6976
rect 4175 6883 4225 6899
rect 4383 6883 4433 6899
rect 4591 6883 4641 6899
rect 4804 6883 4854 6899
rect 5628 6885 5678 6901
rect 5841 6885 5891 6901
rect 6049 6885 6099 6901
rect 6257 6885 6307 6901
rect 1988 6808 2006 6834
rect 2032 6808 2038 6834
rect 3163 6832 3213 6845
rect 3371 6832 3421 6845
rect 3579 6832 3629 6845
rect 3792 6832 3842 6845
rect 1988 6783 2038 6808
rect 4175 6816 4225 6841
rect 4175 6790 4181 6816
rect 4207 6790 4225 6816
rect 4175 6764 4225 6790
rect 4383 6812 4433 6841
rect 4383 6788 4397 6812
rect 4421 6788 4433 6812
rect 4383 6764 4433 6788
rect 4591 6817 4641 6841
rect 4591 6793 4606 6817
rect 4630 6793 4641 6817
rect 4591 6764 4641 6793
rect 4804 6812 4854 6841
rect 8444 6924 8494 6950
rect 8652 6972 8702 7001
rect 8652 6948 8666 6972
rect 8690 6948 8702 6972
rect 8652 6924 8702 6948
rect 8860 6977 8910 7001
rect 8860 6953 8875 6977
rect 8899 6953 8910 6977
rect 8860 6924 8910 6953
rect 9073 6972 9123 7001
rect 11008 7021 11058 7049
rect 11008 7001 11021 7021
rect 11041 7001 11058 7021
rect 9073 6952 9090 6972
rect 9110 6952 9123 6972
rect 9073 6924 9123 6952
rect 11008 6972 11058 7001
rect 11221 7020 11271 7049
rect 11221 6996 11232 7020
rect 11256 6996 11271 7020
rect 11221 6972 11271 6996
rect 11429 7025 11479 7049
rect 11429 7001 11441 7025
rect 11465 7001 11479 7025
rect 11429 6972 11479 7001
rect 11637 7023 11687 7049
rect 11637 6997 11655 7023
rect 11681 6997 11687 7023
rect 11637 6972 11687 6997
rect 13824 7005 13874 7030
rect 12020 6968 12070 6981
rect 12233 6968 12283 6981
rect 12441 6968 12491 6981
rect 12649 6968 12699 6981
rect 13824 6979 13830 7005
rect 13856 6979 13874 7005
rect 4804 6792 4821 6812
rect 4841 6792 4854 6812
rect 4804 6764 4854 6792
rect 346 6726 396 6739
rect 559 6726 609 6739
rect 767 6726 817 6739
rect 975 6726 1025 6739
rect 1359 6725 1409 6741
rect 1572 6725 1622 6741
rect 1780 6725 1830 6741
rect 1988 6725 2038 6741
rect 6640 6811 6690 6839
rect 6640 6791 6653 6811
rect 6673 6791 6690 6811
rect 6640 6762 6690 6791
rect 6853 6810 6903 6839
rect 6853 6786 6864 6810
rect 6888 6786 6903 6810
rect 6853 6762 6903 6786
rect 7061 6815 7111 6839
rect 7061 6791 7073 6815
rect 7097 6791 7111 6815
rect 7061 6762 7111 6791
rect 7269 6813 7319 6839
rect 11008 6914 11058 6930
rect 11221 6914 11271 6930
rect 11429 6914 11479 6930
rect 11637 6914 11687 6930
rect 9456 6862 9506 6878
rect 9664 6862 9714 6878
rect 9872 6862 9922 6878
rect 10085 6862 10135 6878
rect 13824 6953 13874 6979
rect 14032 7001 14082 7030
rect 14032 6977 14046 7001
rect 14070 6977 14082 7001
rect 14032 6953 14082 6977
rect 14240 7006 14290 7030
rect 14240 6982 14255 7006
rect 14279 6982 14290 7006
rect 14240 6953 14290 6982
rect 14453 7001 14503 7030
rect 14453 6981 14470 7001
rect 14490 6981 14503 7001
rect 14453 6953 14503 6981
rect 19105 7051 19155 7067
rect 19313 7051 19363 7067
rect 19521 7051 19571 7067
rect 19734 7051 19784 7067
rect 20118 7053 20168 7066
rect 20326 7053 20376 7066
rect 20534 7053 20584 7066
rect 20747 7053 20797 7066
rect 16289 7000 16339 7028
rect 16289 6980 16302 7000
rect 16322 6980 16339 7000
rect 7269 6787 7287 6813
rect 7313 6787 7319 6813
rect 8444 6811 8494 6824
rect 8652 6811 8702 6824
rect 8860 6811 8910 6824
rect 9073 6811 9123 6824
rect 7269 6762 7319 6787
rect 9456 6795 9506 6820
rect 9456 6769 9462 6795
rect 9488 6769 9506 6795
rect 9456 6743 9506 6769
rect 9664 6791 9714 6820
rect 9664 6767 9678 6791
rect 9702 6767 9714 6791
rect 9664 6743 9714 6767
rect 9872 6796 9922 6820
rect 9872 6772 9887 6796
rect 9911 6772 9922 6796
rect 9872 6743 9922 6772
rect 10085 6791 10135 6820
rect 12020 6840 12070 6868
rect 12020 6820 12033 6840
rect 12053 6820 12070 6840
rect 10085 6771 10102 6791
rect 10122 6771 10135 6791
rect 10085 6743 10135 6771
rect 12020 6791 12070 6820
rect 12233 6839 12283 6868
rect 12233 6815 12244 6839
rect 12268 6815 12283 6839
rect 12233 6791 12283 6815
rect 12441 6844 12491 6868
rect 12441 6820 12453 6844
rect 12477 6820 12491 6844
rect 12441 6791 12491 6820
rect 12649 6842 12699 6868
rect 16289 6951 16339 6980
rect 16502 6999 16552 7028
rect 16502 6975 16513 6999
rect 16537 6975 16552 6999
rect 16502 6951 16552 6975
rect 16710 7004 16760 7028
rect 16710 6980 16722 7004
rect 16746 6980 16760 7004
rect 16710 6951 16760 6980
rect 16918 7002 16968 7028
rect 16918 6976 16936 7002
rect 16962 6976 16968 7002
rect 16918 6951 16968 6976
rect 19105 6984 19155 7009
rect 17301 6947 17351 6960
rect 17514 6947 17564 6960
rect 17722 6947 17772 6960
rect 17930 6947 17980 6960
rect 19105 6958 19111 6984
rect 19137 6958 19155 6984
rect 14836 6891 14886 6907
rect 15044 6891 15094 6907
rect 15252 6891 15302 6907
rect 15465 6891 15515 6907
rect 16289 6893 16339 6909
rect 16502 6893 16552 6909
rect 16710 6893 16760 6909
rect 16918 6893 16968 6909
rect 12649 6816 12667 6842
rect 12693 6816 12699 6842
rect 13824 6840 13874 6853
rect 14032 6840 14082 6853
rect 14240 6840 14290 6853
rect 14453 6840 14503 6853
rect 12649 6791 12699 6816
rect 14836 6824 14886 6849
rect 14836 6798 14842 6824
rect 14868 6798 14886 6824
rect 5627 6705 5677 6718
rect 5840 6705 5890 6718
rect 6048 6705 6098 6718
rect 6256 6705 6306 6718
rect 4175 6651 4225 6664
rect 4383 6651 4433 6664
rect 4591 6651 4641 6664
rect 4804 6651 4854 6664
rect 346 6598 396 6626
rect 346 6578 359 6598
rect 379 6578 396 6598
rect 346 6549 396 6578
rect 559 6597 609 6626
rect 559 6573 570 6597
rect 594 6573 609 6597
rect 559 6549 609 6573
rect 767 6602 817 6626
rect 767 6578 779 6602
rect 803 6578 817 6602
rect 767 6549 817 6578
rect 975 6600 1025 6626
rect 975 6574 993 6600
rect 1019 6574 1025 6600
rect 2955 6597 3005 6613
rect 3163 6597 3213 6613
rect 3371 6597 3421 6613
rect 3584 6597 3634 6613
rect 975 6549 1025 6574
rect 6640 6704 6690 6720
rect 6853 6704 6903 6720
rect 7061 6704 7111 6720
rect 7269 6704 7319 6720
rect 14836 6772 14886 6798
rect 15044 6820 15094 6849
rect 15044 6796 15058 6820
rect 15082 6796 15094 6820
rect 15044 6772 15094 6796
rect 15252 6825 15302 6849
rect 15252 6801 15267 6825
rect 15291 6801 15302 6825
rect 15252 6772 15302 6801
rect 15465 6820 15515 6849
rect 19105 6932 19155 6958
rect 19313 6980 19363 7009
rect 19313 6956 19327 6980
rect 19351 6956 19363 6980
rect 19313 6932 19363 6956
rect 19521 6985 19571 7009
rect 19521 6961 19536 6985
rect 19560 6961 19571 6985
rect 19521 6932 19571 6961
rect 19734 6980 19784 7009
rect 19734 6960 19751 6980
rect 19771 6960 19784 6980
rect 19734 6932 19784 6960
rect 15465 6800 15482 6820
rect 15502 6800 15515 6820
rect 15465 6772 15515 6800
rect 11007 6734 11057 6747
rect 11220 6734 11270 6747
rect 11428 6734 11478 6747
rect 11636 6734 11686 6747
rect 9456 6630 9506 6643
rect 9664 6630 9714 6643
rect 9872 6630 9922 6643
rect 10085 6630 10135 6643
rect 12020 6733 12070 6749
rect 12233 6733 12283 6749
rect 12441 6733 12491 6749
rect 12649 6733 12699 6749
rect 17301 6819 17351 6847
rect 17301 6799 17314 6819
rect 17334 6799 17351 6819
rect 17301 6770 17351 6799
rect 17514 6818 17564 6847
rect 17514 6794 17525 6818
rect 17549 6794 17564 6818
rect 17514 6770 17564 6794
rect 17722 6823 17772 6847
rect 17722 6799 17734 6823
rect 17758 6799 17772 6823
rect 17722 6770 17772 6799
rect 17930 6821 17980 6847
rect 20117 6870 20167 6886
rect 20325 6870 20375 6886
rect 20533 6870 20583 6886
rect 20746 6870 20796 6886
rect 17930 6795 17948 6821
rect 17974 6795 17980 6821
rect 19105 6819 19155 6832
rect 19313 6819 19363 6832
rect 19521 6819 19571 6832
rect 19734 6819 19784 6832
rect 17930 6770 17980 6795
rect 20117 6803 20167 6828
rect 20117 6777 20123 6803
rect 20149 6777 20167 6803
rect 20117 6751 20167 6777
rect 20325 6799 20375 6828
rect 20325 6775 20339 6799
rect 20363 6775 20375 6799
rect 20325 6751 20375 6775
rect 20533 6804 20583 6828
rect 20533 6780 20548 6804
rect 20572 6780 20583 6804
rect 20533 6751 20583 6780
rect 20746 6799 20796 6828
rect 20746 6779 20763 6799
rect 20783 6779 20796 6799
rect 20746 6751 20796 6779
rect 16288 6713 16338 6726
rect 16501 6713 16551 6726
rect 16709 6713 16759 6726
rect 16917 6713 16967 6726
rect 14836 6659 14886 6672
rect 15044 6659 15094 6672
rect 15252 6659 15302 6672
rect 15465 6659 15515 6672
rect 11007 6606 11057 6634
rect 2955 6530 3005 6555
rect 346 6491 396 6507
rect 559 6491 609 6507
rect 767 6491 817 6507
rect 975 6491 1025 6507
rect 2955 6504 2961 6530
rect 2987 6504 3005 6530
rect 2955 6478 3005 6504
rect 3163 6526 3213 6555
rect 3163 6502 3177 6526
rect 3201 6502 3213 6526
rect 3163 6478 3213 6502
rect 3371 6531 3421 6555
rect 3371 6507 3386 6531
rect 3410 6507 3421 6531
rect 3371 6478 3421 6507
rect 3584 6526 3634 6555
rect 5627 6577 5677 6605
rect 3584 6506 3601 6526
rect 3621 6506 3634 6526
rect 5627 6557 5640 6577
rect 5660 6557 5677 6577
rect 3584 6478 3634 6506
rect 5627 6528 5677 6557
rect 5840 6576 5890 6605
rect 5840 6552 5851 6576
rect 5875 6552 5890 6576
rect 5840 6528 5890 6552
rect 6048 6581 6098 6605
rect 6048 6557 6060 6581
rect 6084 6557 6098 6581
rect 6048 6528 6098 6557
rect 6256 6579 6306 6605
rect 6256 6553 6274 6579
rect 6300 6553 6306 6579
rect 8236 6576 8286 6592
rect 8444 6576 8494 6592
rect 8652 6576 8702 6592
rect 8865 6576 8915 6592
rect 6256 6528 6306 6553
rect 11007 6586 11020 6606
rect 11040 6586 11057 6606
rect 1574 6448 1624 6461
rect 1787 6448 1837 6461
rect 1995 6448 2045 6461
rect 2203 6448 2253 6461
rect 8236 6509 8286 6534
rect 5627 6470 5677 6486
rect 5840 6470 5890 6486
rect 6048 6470 6098 6486
rect 6256 6470 6306 6486
rect 8236 6483 8242 6509
rect 8268 6483 8286 6509
rect 8236 6457 8286 6483
rect 8444 6505 8494 6534
rect 8444 6481 8458 6505
rect 8482 6481 8494 6505
rect 8444 6457 8494 6481
rect 8652 6510 8702 6534
rect 8652 6486 8667 6510
rect 8691 6486 8702 6510
rect 8652 6457 8702 6486
rect 8865 6505 8915 6534
rect 11007 6557 11057 6586
rect 11220 6605 11270 6634
rect 11220 6581 11231 6605
rect 11255 6581 11270 6605
rect 11220 6557 11270 6581
rect 11428 6610 11478 6634
rect 11428 6586 11440 6610
rect 11464 6586 11478 6610
rect 11428 6557 11478 6586
rect 11636 6608 11686 6634
rect 11636 6582 11654 6608
rect 11680 6582 11686 6608
rect 13616 6605 13666 6621
rect 13824 6605 13874 6621
rect 14032 6605 14082 6621
rect 14245 6605 14295 6621
rect 11636 6557 11686 6582
rect 17301 6712 17351 6728
rect 17514 6712 17564 6728
rect 17722 6712 17772 6728
rect 17930 6712 17980 6728
rect 20117 6638 20167 6651
rect 20325 6638 20375 6651
rect 20533 6638 20583 6651
rect 20746 6638 20796 6651
rect 8865 6485 8882 6505
rect 8902 6485 8915 6505
rect 13616 6538 13666 6563
rect 11007 6499 11057 6515
rect 11220 6499 11270 6515
rect 11428 6499 11478 6515
rect 11636 6499 11686 6515
rect 13616 6512 13622 6538
rect 13648 6512 13666 6538
rect 8865 6457 8915 6485
rect 13616 6486 13666 6512
rect 13824 6534 13874 6563
rect 13824 6510 13838 6534
rect 13862 6510 13874 6534
rect 13824 6486 13874 6510
rect 14032 6539 14082 6563
rect 14032 6515 14047 6539
rect 14071 6515 14082 6539
rect 14032 6486 14082 6515
rect 14245 6534 14295 6563
rect 16288 6585 16338 6613
rect 14245 6514 14262 6534
rect 14282 6514 14295 6534
rect 16288 6565 16301 6585
rect 16321 6565 16338 6585
rect 14245 6486 14295 6514
rect 16288 6536 16338 6565
rect 16501 6584 16551 6613
rect 16501 6560 16512 6584
rect 16536 6560 16551 6584
rect 16501 6536 16551 6560
rect 16709 6589 16759 6613
rect 16709 6565 16721 6589
rect 16745 6565 16759 6589
rect 16709 6536 16759 6565
rect 16917 6587 16967 6613
rect 16917 6561 16935 6587
rect 16961 6561 16967 6587
rect 18897 6584 18947 6600
rect 19105 6584 19155 6600
rect 19313 6584 19363 6600
rect 19526 6584 19576 6600
rect 16917 6536 16967 6561
rect 6855 6427 6905 6440
rect 7068 6427 7118 6440
rect 7276 6427 7326 6440
rect 7484 6427 7534 6440
rect 2955 6365 3005 6378
rect 3163 6365 3213 6378
rect 3371 6365 3421 6378
rect 3584 6365 3634 6378
rect 1574 6320 1624 6348
rect 1574 6300 1587 6320
rect 1607 6300 1624 6320
rect 1574 6271 1624 6300
rect 1787 6319 1837 6348
rect 1787 6295 1798 6319
rect 1822 6295 1837 6319
rect 1787 6271 1837 6295
rect 1995 6324 2045 6348
rect 1995 6300 2007 6324
rect 2031 6300 2045 6324
rect 1995 6271 2045 6300
rect 2203 6322 2253 6348
rect 2203 6296 2221 6322
rect 2247 6296 2253 6322
rect 4183 6319 4233 6335
rect 4391 6319 4441 6335
rect 4599 6319 4649 6335
rect 4812 6319 4862 6335
rect 2203 6271 2253 6296
rect 12235 6456 12285 6469
rect 12448 6456 12498 6469
rect 12656 6456 12706 6469
rect 12864 6456 12914 6469
rect 8236 6344 8286 6357
rect 8444 6344 8494 6357
rect 8652 6344 8702 6357
rect 8865 6344 8915 6357
rect 18897 6517 18947 6542
rect 16288 6478 16338 6494
rect 16501 6478 16551 6494
rect 16709 6478 16759 6494
rect 16917 6478 16967 6494
rect 18897 6491 18903 6517
rect 18929 6491 18947 6517
rect 18897 6465 18947 6491
rect 19105 6513 19155 6542
rect 19105 6489 19119 6513
rect 19143 6489 19155 6513
rect 19105 6465 19155 6489
rect 19313 6518 19363 6542
rect 19313 6494 19328 6518
rect 19352 6494 19363 6518
rect 19313 6465 19363 6494
rect 19526 6513 19576 6542
rect 19526 6493 19543 6513
rect 19563 6493 19576 6513
rect 19526 6465 19576 6493
rect 17516 6435 17566 6448
rect 17729 6435 17779 6448
rect 17937 6435 17987 6448
rect 18145 6435 18195 6448
rect 13616 6373 13666 6386
rect 13824 6373 13874 6386
rect 14032 6373 14082 6386
rect 14245 6373 14295 6386
rect 4183 6252 4233 6277
rect 1574 6213 1624 6229
rect 1787 6213 1837 6229
rect 1995 6213 2045 6229
rect 2203 6213 2253 6229
rect 4183 6226 4189 6252
rect 4215 6226 4233 6252
rect 4183 6200 4233 6226
rect 4391 6248 4441 6277
rect 4391 6224 4405 6248
rect 4429 6224 4441 6248
rect 4391 6200 4441 6224
rect 4599 6253 4649 6277
rect 4599 6229 4614 6253
rect 4638 6229 4649 6253
rect 4599 6200 4649 6229
rect 4812 6248 4862 6277
rect 6855 6299 6905 6327
rect 4812 6228 4829 6248
rect 4849 6228 4862 6248
rect 6855 6279 6868 6299
rect 6888 6279 6905 6299
rect 4812 6200 4862 6228
rect 6855 6250 6905 6279
rect 7068 6298 7118 6327
rect 7068 6274 7079 6298
rect 7103 6274 7118 6298
rect 7068 6250 7118 6274
rect 7276 6303 7326 6327
rect 7276 6279 7288 6303
rect 7312 6279 7326 6303
rect 7276 6250 7326 6279
rect 7484 6301 7534 6327
rect 12235 6328 12285 6356
rect 7484 6275 7502 6301
rect 7528 6275 7534 6301
rect 9464 6298 9514 6314
rect 9672 6298 9722 6314
rect 9880 6298 9930 6314
rect 10093 6298 10143 6314
rect 7484 6250 7534 6275
rect 12235 6308 12248 6328
rect 12268 6308 12285 6328
rect 354 6162 404 6175
rect 567 6162 617 6175
rect 775 6162 825 6175
rect 983 6162 1033 6175
rect 3170 6085 3220 6101
rect 3378 6085 3428 6101
rect 3586 6085 3636 6101
rect 3799 6085 3849 6101
rect 9464 6231 9514 6256
rect 6855 6192 6905 6208
rect 7068 6192 7118 6208
rect 7276 6192 7326 6208
rect 7484 6192 7534 6208
rect 9464 6205 9470 6231
rect 9496 6205 9514 6231
rect 9464 6179 9514 6205
rect 9672 6227 9722 6256
rect 9672 6203 9686 6227
rect 9710 6203 9722 6227
rect 9672 6179 9722 6203
rect 9880 6232 9930 6256
rect 9880 6208 9895 6232
rect 9919 6208 9930 6232
rect 9880 6179 9930 6208
rect 10093 6227 10143 6256
rect 12235 6279 12285 6308
rect 12448 6327 12498 6356
rect 12448 6303 12459 6327
rect 12483 6303 12498 6327
rect 12448 6279 12498 6303
rect 12656 6332 12706 6356
rect 12656 6308 12668 6332
rect 12692 6308 12706 6332
rect 12656 6279 12706 6308
rect 12864 6330 12914 6356
rect 12864 6304 12882 6330
rect 12908 6304 12914 6330
rect 14844 6327 14894 6343
rect 15052 6327 15102 6343
rect 15260 6327 15310 6343
rect 15473 6327 15523 6343
rect 12864 6279 12914 6304
rect 18897 6352 18947 6365
rect 19105 6352 19155 6365
rect 19313 6352 19363 6365
rect 19526 6352 19576 6365
rect 10093 6207 10110 6227
rect 10130 6207 10143 6227
rect 14844 6260 14894 6285
rect 12235 6221 12285 6237
rect 12448 6221 12498 6237
rect 12656 6221 12706 6237
rect 12864 6221 12914 6237
rect 14844 6234 14850 6260
rect 14876 6234 14894 6260
rect 14844 6208 14894 6234
rect 15052 6256 15102 6285
rect 15052 6232 15066 6256
rect 15090 6232 15102 6256
rect 15052 6208 15102 6232
rect 15260 6261 15310 6285
rect 15260 6237 15275 6261
rect 15299 6237 15310 6261
rect 15260 6208 15310 6237
rect 15473 6256 15523 6285
rect 17516 6307 17566 6335
rect 15473 6236 15490 6256
rect 15510 6236 15523 6256
rect 17516 6287 17529 6307
rect 17549 6287 17566 6307
rect 15473 6208 15523 6236
rect 17516 6258 17566 6287
rect 17729 6306 17779 6335
rect 17729 6282 17740 6306
rect 17764 6282 17779 6306
rect 17729 6258 17779 6282
rect 17937 6311 17987 6335
rect 17937 6287 17949 6311
rect 17973 6287 17987 6311
rect 17937 6258 17987 6287
rect 18145 6309 18195 6335
rect 18145 6283 18163 6309
rect 18189 6283 18195 6309
rect 20125 6306 20175 6322
rect 20333 6306 20383 6322
rect 20541 6306 20591 6322
rect 20754 6306 20804 6322
rect 18145 6258 18195 6283
rect 10093 6179 10143 6207
rect 5635 6141 5685 6154
rect 5848 6141 5898 6154
rect 6056 6141 6106 6154
rect 6264 6141 6314 6154
rect 4183 6087 4233 6100
rect 4391 6087 4441 6100
rect 4599 6087 4649 6100
rect 4812 6087 4862 6100
rect 354 6034 404 6062
rect 354 6014 367 6034
rect 387 6014 404 6034
rect 354 5985 404 6014
rect 567 6033 617 6062
rect 567 6009 578 6033
rect 602 6009 617 6033
rect 567 5985 617 6009
rect 775 6038 825 6062
rect 775 6014 787 6038
rect 811 6014 825 6038
rect 775 5985 825 6014
rect 983 6036 1033 6062
rect 983 6010 1001 6036
rect 1027 6010 1033 6036
rect 983 5985 1033 6010
rect 3170 6018 3220 6043
rect 1366 5981 1416 5994
rect 1579 5981 1629 5994
rect 1787 5981 1837 5994
rect 1995 5981 2045 5994
rect 3170 5992 3176 6018
rect 3202 5992 3220 6018
rect 354 5927 404 5943
rect 567 5927 617 5943
rect 775 5927 825 5943
rect 983 5927 1033 5943
rect 3170 5966 3220 5992
rect 3378 6014 3428 6043
rect 3378 5990 3392 6014
rect 3416 5990 3428 6014
rect 3378 5966 3428 5990
rect 3586 6019 3636 6043
rect 3586 5995 3601 6019
rect 3625 5995 3636 6019
rect 3586 5966 3636 5995
rect 3799 6014 3849 6043
rect 3799 5994 3816 6014
rect 3836 5994 3849 6014
rect 3799 5966 3849 5994
rect 8451 6064 8501 6080
rect 8659 6064 8709 6080
rect 8867 6064 8917 6080
rect 9080 6064 9130 6080
rect 11015 6170 11065 6183
rect 11228 6170 11278 6183
rect 11436 6170 11486 6183
rect 11644 6170 11694 6183
rect 9464 6066 9514 6079
rect 9672 6066 9722 6079
rect 9880 6066 9930 6079
rect 10093 6066 10143 6079
rect 5635 6013 5685 6041
rect 5635 5993 5648 6013
rect 5668 5993 5685 6013
rect 1366 5853 1416 5881
rect 1366 5833 1379 5853
rect 1399 5833 1416 5853
rect 1366 5804 1416 5833
rect 1579 5852 1629 5881
rect 1579 5828 1590 5852
rect 1614 5828 1629 5852
rect 1579 5804 1629 5828
rect 1787 5857 1837 5881
rect 1787 5833 1799 5857
rect 1823 5833 1837 5857
rect 1787 5804 1837 5833
rect 1995 5855 2045 5881
rect 5635 5964 5685 5993
rect 5848 6012 5898 6041
rect 5848 5988 5859 6012
rect 5883 5988 5898 6012
rect 5848 5964 5898 5988
rect 6056 6017 6106 6041
rect 6056 5993 6068 6017
rect 6092 5993 6106 6017
rect 6056 5964 6106 5993
rect 6264 6015 6314 6041
rect 13831 6093 13881 6109
rect 14039 6093 14089 6109
rect 14247 6093 14297 6109
rect 14460 6093 14510 6109
rect 20125 6239 20175 6264
rect 17516 6200 17566 6216
rect 17729 6200 17779 6216
rect 17937 6200 17987 6216
rect 18145 6200 18195 6216
rect 20125 6213 20131 6239
rect 20157 6213 20175 6239
rect 20125 6187 20175 6213
rect 20333 6235 20383 6264
rect 20333 6211 20347 6235
rect 20371 6211 20383 6235
rect 20333 6187 20383 6211
rect 20541 6240 20591 6264
rect 20541 6216 20556 6240
rect 20580 6216 20591 6240
rect 20541 6187 20591 6216
rect 20754 6235 20804 6264
rect 20754 6215 20771 6235
rect 20791 6215 20804 6235
rect 20754 6187 20804 6215
rect 16296 6149 16346 6162
rect 16509 6149 16559 6162
rect 16717 6149 16767 6162
rect 16925 6149 16975 6162
rect 14844 6095 14894 6108
rect 15052 6095 15102 6108
rect 15260 6095 15310 6108
rect 15473 6095 15523 6108
rect 6264 5989 6282 6015
rect 6308 5989 6314 6015
rect 6264 5964 6314 5989
rect 8451 5997 8501 6022
rect 6647 5960 6697 5973
rect 6860 5960 6910 5973
rect 7068 5960 7118 5973
rect 7276 5960 7326 5973
rect 8451 5971 8457 5997
rect 8483 5971 8501 5997
rect 4182 5904 4232 5920
rect 4390 5904 4440 5920
rect 4598 5904 4648 5920
rect 4811 5904 4861 5920
rect 5635 5906 5685 5922
rect 5848 5906 5898 5922
rect 6056 5906 6106 5922
rect 6264 5906 6314 5922
rect 1995 5829 2013 5855
rect 2039 5829 2045 5855
rect 3170 5853 3220 5866
rect 3378 5853 3428 5866
rect 3586 5853 3636 5866
rect 3799 5853 3849 5866
rect 1995 5804 2045 5829
rect 4182 5837 4232 5862
rect 4182 5811 4188 5837
rect 4214 5811 4232 5837
rect 4182 5785 4232 5811
rect 4390 5833 4440 5862
rect 4390 5809 4404 5833
rect 4428 5809 4440 5833
rect 4390 5785 4440 5809
rect 4598 5838 4648 5862
rect 4598 5814 4613 5838
rect 4637 5814 4648 5838
rect 4598 5785 4648 5814
rect 4811 5833 4861 5862
rect 8451 5945 8501 5971
rect 8659 5993 8709 6022
rect 8659 5969 8673 5993
rect 8697 5969 8709 5993
rect 8659 5945 8709 5969
rect 8867 5998 8917 6022
rect 8867 5974 8882 5998
rect 8906 5974 8917 5998
rect 8867 5945 8917 5974
rect 9080 5993 9130 6022
rect 11015 6042 11065 6070
rect 11015 6022 11028 6042
rect 11048 6022 11065 6042
rect 9080 5973 9097 5993
rect 9117 5973 9130 5993
rect 9080 5945 9130 5973
rect 11015 5993 11065 6022
rect 11228 6041 11278 6070
rect 11228 6017 11239 6041
rect 11263 6017 11278 6041
rect 11228 5993 11278 6017
rect 11436 6046 11486 6070
rect 11436 6022 11448 6046
rect 11472 6022 11486 6046
rect 11436 5993 11486 6022
rect 11644 6044 11694 6070
rect 11644 6018 11662 6044
rect 11688 6018 11694 6044
rect 11644 5993 11694 6018
rect 13831 6026 13881 6051
rect 12027 5989 12077 6002
rect 12240 5989 12290 6002
rect 12448 5989 12498 6002
rect 12656 5989 12706 6002
rect 13831 6000 13837 6026
rect 13863 6000 13881 6026
rect 4811 5813 4828 5833
rect 4848 5813 4861 5833
rect 4811 5785 4861 5813
rect 353 5747 403 5760
rect 566 5747 616 5760
rect 774 5747 824 5760
rect 982 5747 1032 5760
rect 1366 5746 1416 5762
rect 1579 5746 1629 5762
rect 1787 5746 1837 5762
rect 1995 5746 2045 5762
rect 6647 5832 6697 5860
rect 6647 5812 6660 5832
rect 6680 5812 6697 5832
rect 6647 5783 6697 5812
rect 6860 5831 6910 5860
rect 6860 5807 6871 5831
rect 6895 5807 6910 5831
rect 6860 5783 6910 5807
rect 7068 5836 7118 5860
rect 7068 5812 7080 5836
rect 7104 5812 7118 5836
rect 7068 5783 7118 5812
rect 7276 5834 7326 5860
rect 11015 5935 11065 5951
rect 11228 5935 11278 5951
rect 11436 5935 11486 5951
rect 11644 5935 11694 5951
rect 9463 5883 9513 5899
rect 9671 5883 9721 5899
rect 9879 5883 9929 5899
rect 10092 5883 10142 5899
rect 13831 5974 13881 6000
rect 14039 6022 14089 6051
rect 14039 5998 14053 6022
rect 14077 5998 14089 6022
rect 14039 5974 14089 5998
rect 14247 6027 14297 6051
rect 14247 6003 14262 6027
rect 14286 6003 14297 6027
rect 14247 5974 14297 6003
rect 14460 6022 14510 6051
rect 14460 6002 14477 6022
rect 14497 6002 14510 6022
rect 14460 5974 14510 6002
rect 19112 6072 19162 6088
rect 19320 6072 19370 6088
rect 19528 6072 19578 6088
rect 19741 6072 19791 6088
rect 20125 6074 20175 6087
rect 20333 6074 20383 6087
rect 20541 6074 20591 6087
rect 20754 6074 20804 6087
rect 16296 6021 16346 6049
rect 16296 6001 16309 6021
rect 16329 6001 16346 6021
rect 7276 5808 7294 5834
rect 7320 5808 7326 5834
rect 8451 5832 8501 5845
rect 8659 5832 8709 5845
rect 8867 5832 8917 5845
rect 9080 5832 9130 5845
rect 7276 5783 7326 5808
rect 9463 5816 9513 5841
rect 9463 5790 9469 5816
rect 9495 5790 9513 5816
rect 9463 5764 9513 5790
rect 9671 5812 9721 5841
rect 9671 5788 9685 5812
rect 9709 5788 9721 5812
rect 9671 5764 9721 5788
rect 9879 5817 9929 5841
rect 9879 5793 9894 5817
rect 9918 5793 9929 5817
rect 9879 5764 9929 5793
rect 10092 5812 10142 5841
rect 12027 5861 12077 5889
rect 12027 5841 12040 5861
rect 12060 5841 12077 5861
rect 10092 5792 10109 5812
rect 10129 5792 10142 5812
rect 10092 5764 10142 5792
rect 12027 5812 12077 5841
rect 12240 5860 12290 5889
rect 12240 5836 12251 5860
rect 12275 5836 12290 5860
rect 12240 5812 12290 5836
rect 12448 5865 12498 5889
rect 12448 5841 12460 5865
rect 12484 5841 12498 5865
rect 12448 5812 12498 5841
rect 12656 5863 12706 5889
rect 16296 5972 16346 6001
rect 16509 6020 16559 6049
rect 16509 5996 16520 6020
rect 16544 5996 16559 6020
rect 16509 5972 16559 5996
rect 16717 6025 16767 6049
rect 16717 6001 16729 6025
rect 16753 6001 16767 6025
rect 16717 5972 16767 6001
rect 16925 6023 16975 6049
rect 16925 5997 16943 6023
rect 16969 5997 16975 6023
rect 16925 5972 16975 5997
rect 19112 6005 19162 6030
rect 17308 5968 17358 5981
rect 17521 5968 17571 5981
rect 17729 5968 17779 5981
rect 17937 5968 17987 5981
rect 19112 5979 19118 6005
rect 19144 5979 19162 6005
rect 14843 5912 14893 5928
rect 15051 5912 15101 5928
rect 15259 5912 15309 5928
rect 15472 5912 15522 5928
rect 16296 5914 16346 5930
rect 16509 5914 16559 5930
rect 16717 5914 16767 5930
rect 16925 5914 16975 5930
rect 12656 5837 12674 5863
rect 12700 5837 12706 5863
rect 13831 5861 13881 5874
rect 14039 5861 14089 5874
rect 14247 5861 14297 5874
rect 14460 5861 14510 5874
rect 12656 5812 12706 5837
rect 14843 5845 14893 5870
rect 14843 5819 14849 5845
rect 14875 5819 14893 5845
rect 5634 5726 5684 5739
rect 5847 5726 5897 5739
rect 6055 5726 6105 5739
rect 6263 5726 6313 5739
rect 3120 5665 3170 5681
rect 3328 5665 3378 5681
rect 3536 5665 3586 5681
rect 3749 5665 3799 5681
rect 4182 5672 4232 5685
rect 4390 5672 4440 5685
rect 4598 5672 4648 5685
rect 4811 5672 4861 5685
rect 353 5619 403 5647
rect 353 5599 366 5619
rect 386 5599 403 5619
rect 353 5570 403 5599
rect 566 5618 616 5647
rect 566 5594 577 5618
rect 601 5594 616 5618
rect 566 5570 616 5594
rect 774 5623 824 5647
rect 774 5599 786 5623
rect 810 5599 824 5623
rect 774 5570 824 5599
rect 982 5621 1032 5647
rect 982 5595 1000 5621
rect 1026 5595 1032 5621
rect 982 5570 1032 5595
rect 3120 5598 3170 5623
rect 3120 5572 3126 5598
rect 3152 5572 3170 5598
rect 3120 5546 3170 5572
rect 3328 5594 3378 5623
rect 3328 5570 3342 5594
rect 3366 5570 3378 5594
rect 3328 5546 3378 5570
rect 3536 5599 3586 5623
rect 3536 5575 3551 5599
rect 3575 5575 3586 5599
rect 3536 5546 3586 5575
rect 3749 5594 3799 5623
rect 3749 5574 3766 5594
rect 3786 5574 3799 5594
rect 3749 5546 3799 5574
rect 6647 5725 6697 5741
rect 6860 5725 6910 5741
rect 7068 5725 7118 5741
rect 7276 5725 7326 5741
rect 14843 5793 14893 5819
rect 15051 5841 15101 5870
rect 15051 5817 15065 5841
rect 15089 5817 15101 5841
rect 15051 5793 15101 5817
rect 15259 5846 15309 5870
rect 15259 5822 15274 5846
rect 15298 5822 15309 5846
rect 15259 5793 15309 5822
rect 15472 5841 15522 5870
rect 19112 5953 19162 5979
rect 19320 6001 19370 6030
rect 19320 5977 19334 6001
rect 19358 5977 19370 6001
rect 19320 5953 19370 5977
rect 19528 6006 19578 6030
rect 19528 5982 19543 6006
rect 19567 5982 19578 6006
rect 19528 5953 19578 5982
rect 19741 6001 19791 6030
rect 19741 5981 19758 6001
rect 19778 5981 19791 6001
rect 19741 5953 19791 5981
rect 15472 5821 15489 5841
rect 15509 5821 15522 5841
rect 15472 5793 15522 5821
rect 11014 5755 11064 5768
rect 11227 5755 11277 5768
rect 11435 5755 11485 5768
rect 11643 5755 11693 5768
rect 8401 5644 8451 5660
rect 8609 5644 8659 5660
rect 8817 5644 8867 5660
rect 9030 5644 9080 5660
rect 9463 5651 9513 5664
rect 9671 5651 9721 5664
rect 9879 5651 9929 5664
rect 10092 5651 10142 5664
rect 12027 5754 12077 5770
rect 12240 5754 12290 5770
rect 12448 5754 12498 5770
rect 12656 5754 12706 5770
rect 17308 5840 17358 5868
rect 17308 5820 17321 5840
rect 17341 5820 17358 5840
rect 17308 5791 17358 5820
rect 17521 5839 17571 5868
rect 17521 5815 17532 5839
rect 17556 5815 17571 5839
rect 17521 5791 17571 5815
rect 17729 5844 17779 5868
rect 17729 5820 17741 5844
rect 17765 5820 17779 5844
rect 17729 5791 17779 5820
rect 17937 5842 17987 5868
rect 20124 5891 20174 5907
rect 20332 5891 20382 5907
rect 20540 5891 20590 5907
rect 20753 5891 20803 5907
rect 17937 5816 17955 5842
rect 17981 5816 17987 5842
rect 19112 5840 19162 5853
rect 19320 5840 19370 5853
rect 19528 5840 19578 5853
rect 19741 5840 19791 5853
rect 17937 5791 17987 5816
rect 20124 5824 20174 5849
rect 20124 5798 20130 5824
rect 20156 5798 20174 5824
rect 20124 5772 20174 5798
rect 20332 5820 20382 5849
rect 20332 5796 20346 5820
rect 20370 5796 20382 5820
rect 20332 5772 20382 5796
rect 20540 5825 20590 5849
rect 20540 5801 20555 5825
rect 20579 5801 20590 5825
rect 20540 5772 20590 5801
rect 20753 5820 20803 5849
rect 20753 5800 20770 5820
rect 20790 5800 20803 5820
rect 20753 5772 20803 5800
rect 16295 5734 16345 5747
rect 16508 5734 16558 5747
rect 16716 5734 16766 5747
rect 16924 5734 16974 5747
rect 13781 5673 13831 5689
rect 13989 5673 14039 5689
rect 14197 5673 14247 5689
rect 14410 5673 14460 5689
rect 14843 5680 14893 5693
rect 15051 5680 15101 5693
rect 15259 5680 15309 5693
rect 15472 5680 15522 5693
rect 5634 5598 5684 5626
rect 353 5512 403 5528
rect 566 5512 616 5528
rect 774 5512 824 5528
rect 982 5512 1032 5528
rect 5634 5578 5647 5598
rect 5667 5578 5684 5598
rect 5634 5549 5684 5578
rect 5847 5597 5897 5626
rect 5847 5573 5858 5597
rect 5882 5573 5897 5597
rect 5847 5549 5897 5573
rect 6055 5602 6105 5626
rect 6055 5578 6067 5602
rect 6091 5578 6105 5602
rect 6055 5549 6105 5578
rect 6263 5600 6313 5626
rect 11014 5627 11064 5655
rect 6263 5574 6281 5600
rect 6307 5574 6313 5600
rect 6263 5549 6313 5574
rect 8401 5577 8451 5602
rect 8401 5551 8407 5577
rect 8433 5551 8451 5577
rect 8401 5525 8451 5551
rect 8609 5573 8659 5602
rect 8609 5549 8623 5573
rect 8647 5549 8659 5573
rect 8609 5525 8659 5549
rect 8817 5578 8867 5602
rect 8817 5554 8832 5578
rect 8856 5554 8867 5578
rect 8817 5525 8867 5554
rect 9030 5573 9080 5602
rect 9030 5553 9047 5573
rect 9067 5553 9080 5573
rect 9030 5525 9080 5553
rect 11014 5607 11027 5627
rect 11047 5607 11064 5627
rect 11014 5578 11064 5607
rect 11227 5626 11277 5655
rect 11227 5602 11238 5626
rect 11262 5602 11277 5626
rect 11227 5578 11277 5602
rect 11435 5631 11485 5655
rect 11435 5607 11447 5631
rect 11471 5607 11485 5631
rect 11435 5578 11485 5607
rect 11643 5629 11693 5655
rect 11643 5603 11661 5629
rect 11687 5603 11693 5629
rect 11643 5578 11693 5603
rect 13781 5606 13831 5631
rect 13781 5580 13787 5606
rect 13813 5580 13831 5606
rect 5634 5491 5684 5507
rect 5847 5491 5897 5507
rect 6055 5491 6105 5507
rect 6263 5491 6313 5507
rect 3120 5433 3170 5446
rect 3328 5433 3378 5446
rect 3536 5433 3586 5446
rect 3749 5433 3799 5446
rect 1421 5420 1471 5433
rect 1634 5420 1684 5433
rect 1842 5420 1892 5433
rect 2050 5420 2100 5433
rect 13781 5554 13831 5580
rect 13989 5602 14039 5631
rect 13989 5578 14003 5602
rect 14027 5578 14039 5602
rect 13989 5554 14039 5578
rect 14197 5607 14247 5631
rect 14197 5583 14212 5607
rect 14236 5583 14247 5607
rect 14197 5554 14247 5583
rect 14410 5602 14460 5631
rect 14410 5582 14427 5602
rect 14447 5582 14460 5602
rect 14410 5554 14460 5582
rect 17308 5733 17358 5749
rect 17521 5733 17571 5749
rect 17729 5733 17779 5749
rect 17937 5733 17987 5749
rect 19062 5652 19112 5668
rect 19270 5652 19320 5668
rect 19478 5652 19528 5668
rect 19691 5652 19741 5668
rect 20124 5659 20174 5672
rect 20332 5659 20382 5672
rect 20540 5659 20590 5672
rect 20753 5659 20803 5672
rect 16295 5606 16345 5634
rect 11014 5520 11064 5536
rect 11227 5520 11277 5536
rect 11435 5520 11485 5536
rect 11643 5520 11693 5536
rect 16295 5586 16308 5606
rect 16328 5586 16345 5606
rect 16295 5557 16345 5586
rect 16508 5605 16558 5634
rect 16508 5581 16519 5605
rect 16543 5581 16558 5605
rect 16508 5557 16558 5581
rect 16716 5610 16766 5634
rect 16716 5586 16728 5610
rect 16752 5586 16766 5610
rect 16716 5557 16766 5586
rect 16924 5608 16974 5634
rect 16924 5582 16942 5608
rect 16968 5582 16974 5608
rect 16924 5557 16974 5582
rect 19062 5585 19112 5610
rect 19062 5559 19068 5585
rect 19094 5559 19112 5585
rect 19062 5533 19112 5559
rect 19270 5581 19320 5610
rect 19270 5557 19284 5581
rect 19308 5557 19320 5581
rect 19270 5533 19320 5557
rect 19478 5586 19528 5610
rect 19478 5562 19493 5586
rect 19517 5562 19528 5586
rect 19478 5533 19528 5562
rect 19691 5581 19741 5610
rect 19691 5561 19708 5581
rect 19728 5561 19741 5581
rect 19691 5533 19741 5561
rect 16295 5499 16345 5515
rect 16508 5499 16558 5515
rect 16716 5499 16766 5515
rect 16924 5499 16974 5515
rect 13781 5441 13831 5454
rect 13989 5441 14039 5454
rect 14197 5441 14247 5454
rect 14410 5441 14460 5454
rect 12082 5428 12132 5441
rect 12295 5428 12345 5441
rect 12503 5428 12553 5441
rect 12711 5428 12761 5441
rect 8401 5412 8451 5425
rect 8609 5412 8659 5425
rect 8817 5412 8867 5425
rect 9030 5412 9080 5425
rect 6702 5399 6752 5412
rect 6915 5399 6965 5412
rect 7123 5399 7173 5412
rect 7331 5399 7381 5412
rect 4188 5338 4238 5354
rect 4396 5338 4446 5354
rect 4604 5338 4654 5354
rect 4817 5338 4867 5354
rect 1421 5292 1471 5320
rect 1421 5272 1434 5292
rect 1454 5272 1471 5292
rect 1421 5243 1471 5272
rect 1634 5291 1684 5320
rect 1634 5267 1645 5291
rect 1669 5267 1684 5291
rect 1634 5243 1684 5267
rect 1842 5296 1892 5320
rect 1842 5272 1854 5296
rect 1878 5272 1892 5296
rect 1842 5243 1892 5272
rect 2050 5294 2100 5320
rect 2050 5268 2068 5294
rect 2094 5268 2100 5294
rect 2050 5243 2100 5268
rect 4188 5271 4238 5296
rect 4188 5245 4194 5271
rect 4220 5245 4238 5271
rect 4188 5219 4238 5245
rect 4396 5267 4446 5296
rect 4396 5243 4410 5267
rect 4434 5243 4446 5267
rect 4396 5219 4446 5243
rect 4604 5272 4654 5296
rect 4604 5248 4619 5272
rect 4643 5248 4654 5272
rect 4604 5219 4654 5248
rect 4817 5267 4867 5296
rect 4817 5247 4834 5267
rect 4854 5247 4867 5267
rect 9469 5317 9519 5333
rect 9677 5317 9727 5333
rect 9885 5317 9935 5333
rect 10098 5317 10148 5333
rect 4817 5219 4867 5247
rect 359 5181 409 5194
rect 572 5181 622 5194
rect 780 5181 830 5194
rect 988 5181 1038 5194
rect 1421 5185 1471 5201
rect 1634 5185 1684 5201
rect 1842 5185 1892 5201
rect 2050 5185 2100 5201
rect 3175 5104 3225 5120
rect 3383 5104 3433 5120
rect 3591 5104 3641 5120
rect 3804 5104 3854 5120
rect 6702 5271 6752 5299
rect 6702 5251 6715 5271
rect 6735 5251 6752 5271
rect 6702 5222 6752 5251
rect 6915 5270 6965 5299
rect 6915 5246 6926 5270
rect 6950 5246 6965 5270
rect 6915 5222 6965 5246
rect 7123 5275 7173 5299
rect 7123 5251 7135 5275
rect 7159 5251 7173 5275
rect 7123 5222 7173 5251
rect 7331 5273 7381 5299
rect 19062 5420 19112 5433
rect 19270 5420 19320 5433
rect 19478 5420 19528 5433
rect 19691 5420 19741 5433
rect 17363 5407 17413 5420
rect 17576 5407 17626 5420
rect 17784 5407 17834 5420
rect 17992 5407 18042 5420
rect 14849 5346 14899 5362
rect 15057 5346 15107 5362
rect 15265 5346 15315 5362
rect 15478 5346 15528 5362
rect 7331 5247 7349 5273
rect 7375 5247 7381 5273
rect 7331 5222 7381 5247
rect 9469 5250 9519 5275
rect 9469 5224 9475 5250
rect 9501 5224 9519 5250
rect 9469 5198 9519 5224
rect 9677 5246 9727 5275
rect 9677 5222 9691 5246
rect 9715 5222 9727 5246
rect 9677 5198 9727 5222
rect 9885 5251 9935 5275
rect 9885 5227 9900 5251
rect 9924 5227 9935 5251
rect 9885 5198 9935 5227
rect 10098 5246 10148 5275
rect 10098 5226 10115 5246
rect 10135 5226 10148 5246
rect 12082 5300 12132 5328
rect 12082 5280 12095 5300
rect 12115 5280 12132 5300
rect 12082 5251 12132 5280
rect 12295 5299 12345 5328
rect 12295 5275 12306 5299
rect 12330 5275 12345 5299
rect 12295 5251 12345 5275
rect 12503 5304 12553 5328
rect 12503 5280 12515 5304
rect 12539 5280 12553 5304
rect 12503 5251 12553 5280
rect 12711 5302 12761 5328
rect 12711 5276 12729 5302
rect 12755 5276 12761 5302
rect 12711 5251 12761 5276
rect 14849 5279 14899 5304
rect 14849 5253 14855 5279
rect 14881 5253 14899 5279
rect 10098 5198 10148 5226
rect 14849 5227 14899 5253
rect 15057 5275 15107 5304
rect 15057 5251 15071 5275
rect 15095 5251 15107 5275
rect 15057 5227 15107 5251
rect 15265 5280 15315 5304
rect 15265 5256 15280 5280
rect 15304 5256 15315 5280
rect 15265 5227 15315 5256
rect 15478 5275 15528 5304
rect 15478 5255 15495 5275
rect 15515 5255 15528 5275
rect 20130 5325 20180 5341
rect 20338 5325 20388 5341
rect 20546 5325 20596 5341
rect 20759 5325 20809 5341
rect 15478 5227 15528 5255
rect 5640 5160 5690 5173
rect 5853 5160 5903 5173
rect 6061 5160 6111 5173
rect 6269 5160 6319 5173
rect 6702 5164 6752 5180
rect 6915 5164 6965 5180
rect 7123 5164 7173 5180
rect 7331 5164 7381 5180
rect 4188 5106 4238 5119
rect 4396 5106 4446 5119
rect 4604 5106 4654 5119
rect 4817 5106 4867 5119
rect 359 5053 409 5081
rect 359 5033 372 5053
rect 392 5033 409 5053
rect 359 5004 409 5033
rect 572 5052 622 5081
rect 572 5028 583 5052
rect 607 5028 622 5052
rect 572 5004 622 5028
rect 780 5057 830 5081
rect 780 5033 792 5057
rect 816 5033 830 5057
rect 780 5004 830 5033
rect 988 5055 1038 5081
rect 988 5029 1006 5055
rect 1032 5029 1038 5055
rect 988 5004 1038 5029
rect 3175 5037 3225 5062
rect 1371 5000 1421 5013
rect 1584 5000 1634 5013
rect 1792 5000 1842 5013
rect 2000 5000 2050 5013
rect 3175 5011 3181 5037
rect 3207 5011 3225 5037
rect 359 4946 409 4962
rect 572 4946 622 4962
rect 780 4946 830 4962
rect 988 4946 1038 4962
rect 3175 4985 3225 5011
rect 3383 5033 3433 5062
rect 3383 5009 3397 5033
rect 3421 5009 3433 5033
rect 3383 4985 3433 5009
rect 3591 5038 3641 5062
rect 3591 5014 3606 5038
rect 3630 5014 3641 5038
rect 3591 4985 3641 5014
rect 3804 5033 3854 5062
rect 3804 5013 3821 5033
rect 3841 5013 3854 5033
rect 3804 4985 3854 5013
rect 8456 5083 8506 5099
rect 8664 5083 8714 5099
rect 8872 5083 8922 5099
rect 9085 5083 9135 5099
rect 11020 5189 11070 5202
rect 11233 5189 11283 5202
rect 11441 5189 11491 5202
rect 11649 5189 11699 5202
rect 12082 5193 12132 5209
rect 12295 5193 12345 5209
rect 12503 5193 12553 5209
rect 12711 5193 12761 5209
rect 9469 5085 9519 5098
rect 9677 5085 9727 5098
rect 9885 5085 9935 5098
rect 10098 5085 10148 5098
rect 5640 5032 5690 5060
rect 5640 5012 5653 5032
rect 5673 5012 5690 5032
rect 1371 4872 1421 4900
rect 1371 4852 1384 4872
rect 1404 4852 1421 4872
rect 1371 4823 1421 4852
rect 1584 4871 1634 4900
rect 1584 4847 1595 4871
rect 1619 4847 1634 4871
rect 1584 4823 1634 4847
rect 1792 4876 1842 4900
rect 1792 4852 1804 4876
rect 1828 4852 1842 4876
rect 1792 4823 1842 4852
rect 2000 4874 2050 4900
rect 5640 4983 5690 5012
rect 5853 5031 5903 5060
rect 5853 5007 5864 5031
rect 5888 5007 5903 5031
rect 5853 4983 5903 5007
rect 6061 5036 6111 5060
rect 6061 5012 6073 5036
rect 6097 5012 6111 5036
rect 6061 4983 6111 5012
rect 6269 5034 6319 5060
rect 13836 5112 13886 5128
rect 14044 5112 14094 5128
rect 14252 5112 14302 5128
rect 14465 5112 14515 5128
rect 17363 5279 17413 5307
rect 17363 5259 17376 5279
rect 17396 5259 17413 5279
rect 17363 5230 17413 5259
rect 17576 5278 17626 5307
rect 17576 5254 17587 5278
rect 17611 5254 17626 5278
rect 17576 5230 17626 5254
rect 17784 5283 17834 5307
rect 17784 5259 17796 5283
rect 17820 5259 17834 5283
rect 17784 5230 17834 5259
rect 17992 5281 18042 5307
rect 17992 5255 18010 5281
rect 18036 5255 18042 5281
rect 17992 5230 18042 5255
rect 20130 5258 20180 5283
rect 20130 5232 20136 5258
rect 20162 5232 20180 5258
rect 20130 5206 20180 5232
rect 20338 5254 20388 5283
rect 20338 5230 20352 5254
rect 20376 5230 20388 5254
rect 20338 5206 20388 5230
rect 20546 5259 20596 5283
rect 20546 5235 20561 5259
rect 20585 5235 20596 5259
rect 20546 5206 20596 5235
rect 20759 5254 20809 5283
rect 20759 5234 20776 5254
rect 20796 5234 20809 5254
rect 20759 5206 20809 5234
rect 16301 5168 16351 5181
rect 16514 5168 16564 5181
rect 16722 5168 16772 5181
rect 16930 5168 16980 5181
rect 17363 5172 17413 5188
rect 17576 5172 17626 5188
rect 17784 5172 17834 5188
rect 17992 5172 18042 5188
rect 14849 5114 14899 5127
rect 15057 5114 15107 5127
rect 15265 5114 15315 5127
rect 15478 5114 15528 5127
rect 6269 5008 6287 5034
rect 6313 5008 6319 5034
rect 6269 4983 6319 5008
rect 8456 5016 8506 5041
rect 6652 4979 6702 4992
rect 6865 4979 6915 4992
rect 7073 4979 7123 4992
rect 7281 4979 7331 4992
rect 8456 4990 8462 5016
rect 8488 4990 8506 5016
rect 4187 4923 4237 4939
rect 4395 4923 4445 4939
rect 4603 4923 4653 4939
rect 4816 4923 4866 4939
rect 5640 4925 5690 4941
rect 5853 4925 5903 4941
rect 6061 4925 6111 4941
rect 6269 4925 6319 4941
rect 2000 4848 2018 4874
rect 2044 4848 2050 4874
rect 3175 4872 3225 4885
rect 3383 4872 3433 4885
rect 3591 4872 3641 4885
rect 3804 4872 3854 4885
rect 2000 4823 2050 4848
rect 4187 4856 4237 4881
rect 4187 4830 4193 4856
rect 4219 4830 4237 4856
rect 4187 4804 4237 4830
rect 4395 4852 4445 4881
rect 4395 4828 4409 4852
rect 4433 4828 4445 4852
rect 4395 4804 4445 4828
rect 4603 4857 4653 4881
rect 4603 4833 4618 4857
rect 4642 4833 4653 4857
rect 4603 4804 4653 4833
rect 4816 4852 4866 4881
rect 8456 4964 8506 4990
rect 8664 5012 8714 5041
rect 8664 4988 8678 5012
rect 8702 4988 8714 5012
rect 8664 4964 8714 4988
rect 8872 5017 8922 5041
rect 8872 4993 8887 5017
rect 8911 4993 8922 5017
rect 8872 4964 8922 4993
rect 9085 5012 9135 5041
rect 11020 5061 11070 5089
rect 11020 5041 11033 5061
rect 11053 5041 11070 5061
rect 9085 4992 9102 5012
rect 9122 4992 9135 5012
rect 9085 4964 9135 4992
rect 11020 5012 11070 5041
rect 11233 5060 11283 5089
rect 11233 5036 11244 5060
rect 11268 5036 11283 5060
rect 11233 5012 11283 5036
rect 11441 5065 11491 5089
rect 11441 5041 11453 5065
rect 11477 5041 11491 5065
rect 11441 5012 11491 5041
rect 11649 5063 11699 5089
rect 11649 5037 11667 5063
rect 11693 5037 11699 5063
rect 11649 5012 11699 5037
rect 13836 5045 13886 5070
rect 12032 5008 12082 5021
rect 12245 5008 12295 5021
rect 12453 5008 12503 5021
rect 12661 5008 12711 5021
rect 13836 5019 13842 5045
rect 13868 5019 13886 5045
rect 4816 4832 4833 4852
rect 4853 4832 4866 4852
rect 4816 4804 4866 4832
rect 358 4766 408 4779
rect 571 4766 621 4779
rect 779 4766 829 4779
rect 987 4766 1037 4779
rect 1371 4765 1421 4781
rect 1584 4765 1634 4781
rect 1792 4765 1842 4781
rect 2000 4765 2050 4781
rect 6652 4851 6702 4879
rect 6652 4831 6665 4851
rect 6685 4831 6702 4851
rect 6652 4802 6702 4831
rect 6865 4850 6915 4879
rect 6865 4826 6876 4850
rect 6900 4826 6915 4850
rect 6865 4802 6915 4826
rect 7073 4855 7123 4879
rect 7073 4831 7085 4855
rect 7109 4831 7123 4855
rect 7073 4802 7123 4831
rect 7281 4853 7331 4879
rect 11020 4954 11070 4970
rect 11233 4954 11283 4970
rect 11441 4954 11491 4970
rect 11649 4954 11699 4970
rect 9468 4902 9518 4918
rect 9676 4902 9726 4918
rect 9884 4902 9934 4918
rect 10097 4902 10147 4918
rect 13836 4993 13886 5019
rect 14044 5041 14094 5070
rect 14044 5017 14058 5041
rect 14082 5017 14094 5041
rect 14044 4993 14094 5017
rect 14252 5046 14302 5070
rect 14252 5022 14267 5046
rect 14291 5022 14302 5046
rect 14252 4993 14302 5022
rect 14465 5041 14515 5070
rect 14465 5021 14482 5041
rect 14502 5021 14515 5041
rect 14465 4993 14515 5021
rect 19117 5091 19167 5107
rect 19325 5091 19375 5107
rect 19533 5091 19583 5107
rect 19746 5091 19796 5107
rect 20130 5093 20180 5106
rect 20338 5093 20388 5106
rect 20546 5093 20596 5106
rect 20759 5093 20809 5106
rect 16301 5040 16351 5068
rect 16301 5020 16314 5040
rect 16334 5020 16351 5040
rect 7281 4827 7299 4853
rect 7325 4827 7331 4853
rect 8456 4851 8506 4864
rect 8664 4851 8714 4864
rect 8872 4851 8922 4864
rect 9085 4851 9135 4864
rect 7281 4802 7331 4827
rect 9468 4835 9518 4860
rect 9468 4809 9474 4835
rect 9500 4809 9518 4835
rect 9468 4783 9518 4809
rect 9676 4831 9726 4860
rect 9676 4807 9690 4831
rect 9714 4807 9726 4831
rect 9676 4783 9726 4807
rect 9884 4836 9934 4860
rect 9884 4812 9899 4836
rect 9923 4812 9934 4836
rect 9884 4783 9934 4812
rect 10097 4831 10147 4860
rect 12032 4880 12082 4908
rect 12032 4860 12045 4880
rect 12065 4860 12082 4880
rect 10097 4811 10114 4831
rect 10134 4811 10147 4831
rect 10097 4783 10147 4811
rect 12032 4831 12082 4860
rect 12245 4879 12295 4908
rect 12245 4855 12256 4879
rect 12280 4855 12295 4879
rect 12245 4831 12295 4855
rect 12453 4884 12503 4908
rect 12453 4860 12465 4884
rect 12489 4860 12503 4884
rect 12453 4831 12503 4860
rect 12661 4882 12711 4908
rect 16301 4991 16351 5020
rect 16514 5039 16564 5068
rect 16514 5015 16525 5039
rect 16549 5015 16564 5039
rect 16514 4991 16564 5015
rect 16722 5044 16772 5068
rect 16722 5020 16734 5044
rect 16758 5020 16772 5044
rect 16722 4991 16772 5020
rect 16930 5042 16980 5068
rect 16930 5016 16948 5042
rect 16974 5016 16980 5042
rect 16930 4991 16980 5016
rect 19117 5024 19167 5049
rect 17313 4987 17363 5000
rect 17526 4987 17576 5000
rect 17734 4987 17784 5000
rect 17942 4987 17992 5000
rect 19117 4998 19123 5024
rect 19149 4998 19167 5024
rect 14848 4931 14898 4947
rect 15056 4931 15106 4947
rect 15264 4931 15314 4947
rect 15477 4931 15527 4947
rect 16301 4933 16351 4949
rect 16514 4933 16564 4949
rect 16722 4933 16772 4949
rect 16930 4933 16980 4949
rect 12661 4856 12679 4882
rect 12705 4856 12711 4882
rect 13836 4880 13886 4893
rect 14044 4880 14094 4893
rect 14252 4880 14302 4893
rect 14465 4880 14515 4893
rect 12661 4831 12711 4856
rect 14848 4864 14898 4889
rect 14848 4838 14854 4864
rect 14880 4838 14898 4864
rect 5639 4745 5689 4758
rect 5852 4745 5902 4758
rect 6060 4745 6110 4758
rect 6268 4745 6318 4758
rect 4187 4691 4237 4704
rect 4395 4691 4445 4704
rect 4603 4691 4653 4704
rect 4816 4691 4866 4704
rect 2880 4672 2930 4688
rect 3088 4672 3138 4688
rect 3296 4672 3346 4688
rect 3509 4672 3559 4688
rect 358 4638 408 4666
rect 358 4618 371 4638
rect 391 4618 408 4638
rect 358 4589 408 4618
rect 571 4637 621 4666
rect 571 4613 582 4637
rect 606 4613 621 4637
rect 571 4589 621 4613
rect 779 4642 829 4666
rect 779 4618 791 4642
rect 815 4618 829 4642
rect 779 4589 829 4618
rect 987 4640 1037 4666
rect 987 4614 1005 4640
rect 1031 4614 1037 4640
rect 6652 4744 6702 4760
rect 6865 4744 6915 4760
rect 7073 4744 7123 4760
rect 7281 4744 7331 4760
rect 14848 4812 14898 4838
rect 15056 4860 15106 4889
rect 15056 4836 15070 4860
rect 15094 4836 15106 4860
rect 15056 4812 15106 4836
rect 15264 4865 15314 4889
rect 15264 4841 15279 4865
rect 15303 4841 15314 4865
rect 15264 4812 15314 4841
rect 15477 4860 15527 4889
rect 19117 4972 19167 4998
rect 19325 5020 19375 5049
rect 19325 4996 19339 5020
rect 19363 4996 19375 5020
rect 19325 4972 19375 4996
rect 19533 5025 19583 5049
rect 19533 5001 19548 5025
rect 19572 5001 19583 5025
rect 19533 4972 19583 5001
rect 19746 5020 19796 5049
rect 19746 5000 19763 5020
rect 19783 5000 19796 5020
rect 19746 4972 19796 5000
rect 15477 4840 15494 4860
rect 15514 4840 15527 4860
rect 15477 4812 15527 4840
rect 11019 4774 11069 4787
rect 11232 4774 11282 4787
rect 11440 4774 11490 4787
rect 11648 4774 11698 4787
rect 9468 4670 9518 4683
rect 9676 4670 9726 4683
rect 9884 4670 9934 4683
rect 10097 4670 10147 4683
rect 12032 4773 12082 4789
rect 12245 4773 12295 4789
rect 12453 4773 12503 4789
rect 12661 4773 12711 4789
rect 17313 4859 17363 4887
rect 17313 4839 17326 4859
rect 17346 4839 17363 4859
rect 17313 4810 17363 4839
rect 17526 4858 17576 4887
rect 17526 4834 17537 4858
rect 17561 4834 17576 4858
rect 17526 4810 17576 4834
rect 17734 4863 17784 4887
rect 17734 4839 17746 4863
rect 17770 4839 17784 4863
rect 17734 4810 17784 4839
rect 17942 4861 17992 4887
rect 20129 4910 20179 4926
rect 20337 4910 20387 4926
rect 20545 4910 20595 4926
rect 20758 4910 20808 4926
rect 17942 4835 17960 4861
rect 17986 4835 17992 4861
rect 19117 4859 19167 4872
rect 19325 4859 19375 4872
rect 19533 4859 19583 4872
rect 19746 4859 19796 4872
rect 17942 4810 17992 4835
rect 20129 4843 20179 4868
rect 20129 4817 20135 4843
rect 20161 4817 20179 4843
rect 20129 4791 20179 4817
rect 20337 4839 20387 4868
rect 20337 4815 20351 4839
rect 20375 4815 20387 4839
rect 20337 4791 20387 4815
rect 20545 4844 20595 4868
rect 20545 4820 20560 4844
rect 20584 4820 20595 4844
rect 20545 4791 20595 4820
rect 20758 4839 20808 4868
rect 20758 4819 20775 4839
rect 20795 4819 20808 4839
rect 20758 4791 20808 4819
rect 16300 4753 16350 4766
rect 16513 4753 16563 4766
rect 16721 4753 16771 4766
rect 16929 4753 16979 4766
rect 14848 4699 14898 4712
rect 15056 4699 15106 4712
rect 15264 4699 15314 4712
rect 15477 4699 15527 4712
rect 13541 4680 13591 4696
rect 13749 4680 13799 4696
rect 13957 4680 14007 4696
rect 14170 4680 14220 4696
rect 8161 4651 8211 4667
rect 8369 4651 8419 4667
rect 8577 4651 8627 4667
rect 8790 4651 8840 4667
rect 987 4589 1037 4614
rect 2880 4605 2930 4630
rect 2880 4579 2886 4605
rect 2912 4579 2930 4605
rect 2880 4553 2930 4579
rect 3088 4601 3138 4630
rect 3088 4577 3102 4601
rect 3126 4577 3138 4601
rect 3088 4553 3138 4577
rect 3296 4606 3346 4630
rect 3296 4582 3311 4606
rect 3335 4582 3346 4606
rect 3296 4553 3346 4582
rect 3509 4601 3559 4630
rect 3509 4581 3526 4601
rect 3546 4581 3559 4601
rect 5639 4617 5689 4645
rect 3509 4553 3559 4581
rect 358 4531 408 4547
rect 571 4531 621 4547
rect 779 4531 829 4547
rect 987 4531 1037 4547
rect 1669 4456 1719 4469
rect 1882 4456 1932 4469
rect 2090 4456 2140 4469
rect 2298 4456 2348 4469
rect 5639 4597 5652 4617
rect 5672 4597 5689 4617
rect 5639 4568 5689 4597
rect 5852 4616 5902 4645
rect 5852 4592 5863 4616
rect 5887 4592 5902 4616
rect 5852 4568 5902 4592
rect 6060 4621 6110 4645
rect 6060 4597 6072 4621
rect 6096 4597 6110 4621
rect 6060 4568 6110 4597
rect 6268 4619 6318 4645
rect 6268 4593 6286 4619
rect 6312 4593 6318 4619
rect 11019 4646 11069 4674
rect 11019 4626 11032 4646
rect 11052 4626 11069 4646
rect 6268 4568 6318 4593
rect 8161 4584 8211 4609
rect 8161 4558 8167 4584
rect 8193 4558 8211 4584
rect 8161 4532 8211 4558
rect 8369 4580 8419 4609
rect 8369 4556 8383 4580
rect 8407 4556 8419 4580
rect 8369 4532 8419 4556
rect 8577 4585 8627 4609
rect 8577 4561 8592 4585
rect 8616 4561 8627 4585
rect 8577 4532 8627 4561
rect 8790 4580 8840 4609
rect 8790 4560 8807 4580
rect 8827 4560 8840 4580
rect 11019 4597 11069 4626
rect 11232 4645 11282 4674
rect 11232 4621 11243 4645
rect 11267 4621 11282 4645
rect 11232 4597 11282 4621
rect 11440 4650 11490 4674
rect 11440 4626 11452 4650
rect 11476 4626 11490 4650
rect 11440 4597 11490 4626
rect 11648 4648 11698 4674
rect 11648 4622 11666 4648
rect 11692 4622 11698 4648
rect 17313 4752 17363 4768
rect 17526 4752 17576 4768
rect 17734 4752 17784 4768
rect 17942 4752 17992 4768
rect 20129 4678 20179 4691
rect 20337 4678 20387 4691
rect 20545 4678 20595 4691
rect 20758 4678 20808 4691
rect 18822 4659 18872 4675
rect 19030 4659 19080 4675
rect 19238 4659 19288 4675
rect 19451 4659 19501 4675
rect 11648 4597 11698 4622
rect 13541 4613 13591 4638
rect 8790 4532 8840 4560
rect 5639 4510 5689 4526
rect 5852 4510 5902 4526
rect 6060 4510 6110 4526
rect 6268 4510 6318 4526
rect 2880 4440 2930 4453
rect 3088 4440 3138 4453
rect 3296 4440 3346 4453
rect 3509 4440 3559 4453
rect 6950 4435 7000 4448
rect 7163 4435 7213 4448
rect 7371 4435 7421 4448
rect 7579 4435 7629 4448
rect 4191 4362 4241 4378
rect 4399 4362 4449 4378
rect 4607 4362 4657 4378
rect 4820 4362 4870 4378
rect 1669 4328 1719 4356
rect 1669 4308 1682 4328
rect 1702 4308 1719 4328
rect 1669 4279 1719 4308
rect 1882 4327 1932 4356
rect 1882 4303 1893 4327
rect 1917 4303 1932 4327
rect 1882 4279 1932 4303
rect 2090 4332 2140 4356
rect 2090 4308 2102 4332
rect 2126 4308 2140 4332
rect 2090 4279 2140 4308
rect 2298 4330 2348 4356
rect 2298 4304 2316 4330
rect 2342 4304 2348 4330
rect 2298 4279 2348 4304
rect 4191 4295 4241 4320
rect 4191 4269 4197 4295
rect 4223 4269 4241 4295
rect 4191 4243 4241 4269
rect 4399 4291 4449 4320
rect 4399 4267 4413 4291
rect 4437 4267 4449 4291
rect 4399 4243 4449 4267
rect 4607 4296 4657 4320
rect 4607 4272 4622 4296
rect 4646 4272 4657 4296
rect 4607 4243 4657 4272
rect 4820 4291 4870 4320
rect 4820 4271 4837 4291
rect 4857 4271 4870 4291
rect 13541 4587 13547 4613
rect 13573 4587 13591 4613
rect 13541 4561 13591 4587
rect 13749 4609 13799 4638
rect 13749 4585 13763 4609
rect 13787 4585 13799 4609
rect 13749 4561 13799 4585
rect 13957 4614 14007 4638
rect 13957 4590 13972 4614
rect 13996 4590 14007 4614
rect 13957 4561 14007 4590
rect 14170 4609 14220 4638
rect 14170 4589 14187 4609
rect 14207 4589 14220 4609
rect 16300 4625 16350 4653
rect 14170 4561 14220 4589
rect 11019 4539 11069 4555
rect 11232 4539 11282 4555
rect 11440 4539 11490 4555
rect 11648 4539 11698 4555
rect 12330 4464 12380 4477
rect 12543 4464 12593 4477
rect 12751 4464 12801 4477
rect 12959 4464 13009 4477
rect 8161 4419 8211 4432
rect 8369 4419 8419 4432
rect 8577 4419 8627 4432
rect 8790 4419 8840 4432
rect 9472 4341 9522 4357
rect 9680 4341 9730 4357
rect 9888 4341 9938 4357
rect 10101 4341 10151 4357
rect 6950 4307 7000 4335
rect 4820 4243 4870 4271
rect 6950 4287 6963 4307
rect 6983 4287 7000 4307
rect 6950 4258 7000 4287
rect 7163 4306 7213 4335
rect 7163 4282 7174 4306
rect 7198 4282 7213 4306
rect 7163 4258 7213 4282
rect 7371 4311 7421 4335
rect 7371 4287 7383 4311
rect 7407 4287 7421 4311
rect 7371 4258 7421 4287
rect 7579 4309 7629 4335
rect 7579 4283 7597 4309
rect 7623 4283 7629 4309
rect 16300 4605 16313 4625
rect 16333 4605 16350 4625
rect 16300 4576 16350 4605
rect 16513 4624 16563 4653
rect 16513 4600 16524 4624
rect 16548 4600 16563 4624
rect 16513 4576 16563 4600
rect 16721 4629 16771 4653
rect 16721 4605 16733 4629
rect 16757 4605 16771 4629
rect 16721 4576 16771 4605
rect 16929 4627 16979 4653
rect 16929 4601 16947 4627
rect 16973 4601 16979 4627
rect 16929 4576 16979 4601
rect 18822 4592 18872 4617
rect 18822 4566 18828 4592
rect 18854 4566 18872 4592
rect 18822 4540 18872 4566
rect 19030 4588 19080 4617
rect 19030 4564 19044 4588
rect 19068 4564 19080 4588
rect 19030 4540 19080 4564
rect 19238 4593 19288 4617
rect 19238 4569 19253 4593
rect 19277 4569 19288 4593
rect 19238 4540 19288 4569
rect 19451 4588 19501 4617
rect 19451 4568 19468 4588
rect 19488 4568 19501 4588
rect 19451 4540 19501 4568
rect 16300 4518 16350 4534
rect 16513 4518 16563 4534
rect 16721 4518 16771 4534
rect 16929 4518 16979 4534
rect 13541 4448 13591 4461
rect 13749 4448 13799 4461
rect 13957 4448 14007 4461
rect 14170 4448 14220 4461
rect 17611 4443 17661 4456
rect 17824 4443 17874 4456
rect 18032 4443 18082 4456
rect 18240 4443 18290 4456
rect 14852 4370 14902 4386
rect 15060 4370 15110 4386
rect 15268 4370 15318 4386
rect 15481 4370 15531 4386
rect 12330 4336 12380 4364
rect 7579 4258 7629 4283
rect 9472 4274 9522 4299
rect 1669 4221 1719 4237
rect 1882 4221 1932 4237
rect 2090 4221 2140 4237
rect 2298 4221 2348 4237
rect 362 4205 412 4218
rect 575 4205 625 4218
rect 783 4205 833 4218
rect 991 4205 1041 4218
rect 3178 4128 3228 4144
rect 3386 4128 3436 4144
rect 3594 4128 3644 4144
rect 3807 4128 3857 4144
rect 9472 4248 9478 4274
rect 9504 4248 9522 4274
rect 9472 4222 9522 4248
rect 9680 4270 9730 4299
rect 9680 4246 9694 4270
rect 9718 4246 9730 4270
rect 9680 4222 9730 4246
rect 9888 4275 9938 4299
rect 9888 4251 9903 4275
rect 9927 4251 9938 4275
rect 9888 4222 9938 4251
rect 10101 4270 10151 4299
rect 12330 4316 12343 4336
rect 12363 4316 12380 4336
rect 12330 4287 12380 4316
rect 12543 4335 12593 4364
rect 12543 4311 12554 4335
rect 12578 4311 12593 4335
rect 12543 4287 12593 4311
rect 12751 4340 12801 4364
rect 12751 4316 12763 4340
rect 12787 4316 12801 4340
rect 12751 4287 12801 4316
rect 12959 4338 13009 4364
rect 12959 4312 12977 4338
rect 13003 4312 13009 4338
rect 12959 4287 13009 4312
rect 14852 4303 14902 4328
rect 10101 4250 10118 4270
rect 10138 4250 10151 4270
rect 10101 4222 10151 4250
rect 14852 4277 14858 4303
rect 14884 4277 14902 4303
rect 14852 4251 14902 4277
rect 15060 4299 15110 4328
rect 15060 4275 15074 4299
rect 15098 4275 15110 4299
rect 15060 4251 15110 4275
rect 15268 4304 15318 4328
rect 15268 4280 15283 4304
rect 15307 4280 15318 4304
rect 15268 4251 15318 4280
rect 15481 4299 15531 4328
rect 15481 4279 15498 4299
rect 15518 4279 15531 4299
rect 18822 4427 18872 4440
rect 19030 4427 19080 4440
rect 19238 4427 19288 4440
rect 19451 4427 19501 4440
rect 20133 4349 20183 4365
rect 20341 4349 20391 4365
rect 20549 4349 20599 4365
rect 20762 4349 20812 4365
rect 17611 4315 17661 4343
rect 15481 4251 15531 4279
rect 17611 4295 17624 4315
rect 17644 4295 17661 4315
rect 17611 4266 17661 4295
rect 17824 4314 17874 4343
rect 17824 4290 17835 4314
rect 17859 4290 17874 4314
rect 17824 4266 17874 4290
rect 18032 4319 18082 4343
rect 18032 4295 18044 4319
rect 18068 4295 18082 4319
rect 18032 4266 18082 4295
rect 18240 4317 18290 4343
rect 18240 4291 18258 4317
rect 18284 4291 18290 4317
rect 18240 4266 18290 4291
rect 20133 4282 20183 4307
rect 12330 4229 12380 4245
rect 12543 4229 12593 4245
rect 12751 4229 12801 4245
rect 12959 4229 13009 4245
rect 6950 4200 7000 4216
rect 7163 4200 7213 4216
rect 7371 4200 7421 4216
rect 7579 4200 7629 4216
rect 5643 4184 5693 4197
rect 5856 4184 5906 4197
rect 6064 4184 6114 4197
rect 6272 4184 6322 4197
rect 4191 4130 4241 4143
rect 4399 4130 4449 4143
rect 4607 4130 4657 4143
rect 4820 4130 4870 4143
rect 362 4077 412 4105
rect 362 4057 375 4077
rect 395 4057 412 4077
rect 362 4028 412 4057
rect 575 4076 625 4105
rect 575 4052 586 4076
rect 610 4052 625 4076
rect 575 4028 625 4052
rect 783 4081 833 4105
rect 783 4057 795 4081
rect 819 4057 833 4081
rect 783 4028 833 4057
rect 991 4079 1041 4105
rect 991 4053 1009 4079
rect 1035 4053 1041 4079
rect 991 4028 1041 4053
rect 3178 4061 3228 4086
rect 1374 4024 1424 4037
rect 1587 4024 1637 4037
rect 1795 4024 1845 4037
rect 2003 4024 2053 4037
rect 3178 4035 3184 4061
rect 3210 4035 3228 4061
rect 362 3970 412 3986
rect 575 3970 625 3986
rect 783 3970 833 3986
rect 991 3970 1041 3986
rect 3178 4009 3228 4035
rect 3386 4057 3436 4086
rect 3386 4033 3400 4057
rect 3424 4033 3436 4057
rect 3386 4009 3436 4033
rect 3594 4062 3644 4086
rect 3594 4038 3609 4062
rect 3633 4038 3644 4062
rect 3594 4009 3644 4038
rect 3807 4057 3857 4086
rect 3807 4037 3824 4057
rect 3844 4037 3857 4057
rect 3807 4009 3857 4037
rect 8459 4107 8509 4123
rect 8667 4107 8717 4123
rect 8875 4107 8925 4123
rect 9088 4107 9138 4123
rect 11023 4213 11073 4226
rect 11236 4213 11286 4226
rect 11444 4213 11494 4226
rect 11652 4213 11702 4226
rect 9472 4109 9522 4122
rect 9680 4109 9730 4122
rect 9888 4109 9938 4122
rect 10101 4109 10151 4122
rect 5643 4056 5693 4084
rect 5643 4036 5656 4056
rect 5676 4036 5693 4056
rect 1374 3896 1424 3924
rect 1374 3876 1387 3896
rect 1407 3876 1424 3896
rect 1374 3847 1424 3876
rect 1587 3895 1637 3924
rect 1587 3871 1598 3895
rect 1622 3871 1637 3895
rect 1587 3847 1637 3871
rect 1795 3900 1845 3924
rect 1795 3876 1807 3900
rect 1831 3876 1845 3900
rect 1795 3847 1845 3876
rect 2003 3898 2053 3924
rect 5643 4007 5693 4036
rect 5856 4055 5906 4084
rect 5856 4031 5867 4055
rect 5891 4031 5906 4055
rect 5856 4007 5906 4031
rect 6064 4060 6114 4084
rect 6064 4036 6076 4060
rect 6100 4036 6114 4060
rect 6064 4007 6114 4036
rect 6272 4058 6322 4084
rect 13839 4136 13889 4152
rect 14047 4136 14097 4152
rect 14255 4136 14305 4152
rect 14468 4136 14518 4152
rect 20133 4256 20139 4282
rect 20165 4256 20183 4282
rect 20133 4230 20183 4256
rect 20341 4278 20391 4307
rect 20341 4254 20355 4278
rect 20379 4254 20391 4278
rect 20341 4230 20391 4254
rect 20549 4283 20599 4307
rect 20549 4259 20564 4283
rect 20588 4259 20599 4283
rect 20549 4230 20599 4259
rect 20762 4278 20812 4307
rect 20762 4258 20779 4278
rect 20799 4258 20812 4278
rect 20762 4230 20812 4258
rect 17611 4208 17661 4224
rect 17824 4208 17874 4224
rect 18032 4208 18082 4224
rect 18240 4208 18290 4224
rect 16304 4192 16354 4205
rect 16517 4192 16567 4205
rect 16725 4192 16775 4205
rect 16933 4192 16983 4205
rect 14852 4138 14902 4151
rect 15060 4138 15110 4151
rect 15268 4138 15318 4151
rect 15481 4138 15531 4151
rect 6272 4032 6290 4058
rect 6316 4032 6322 4058
rect 6272 4007 6322 4032
rect 8459 4040 8509 4065
rect 6655 4003 6705 4016
rect 6868 4003 6918 4016
rect 7076 4003 7126 4016
rect 7284 4003 7334 4016
rect 8459 4014 8465 4040
rect 8491 4014 8509 4040
rect 4190 3947 4240 3963
rect 4398 3947 4448 3963
rect 4606 3947 4656 3963
rect 4819 3947 4869 3963
rect 5643 3949 5693 3965
rect 5856 3949 5906 3965
rect 6064 3949 6114 3965
rect 6272 3949 6322 3965
rect 2003 3872 2021 3898
rect 2047 3872 2053 3898
rect 3178 3896 3228 3909
rect 3386 3896 3436 3909
rect 3594 3896 3644 3909
rect 3807 3896 3857 3909
rect 2003 3847 2053 3872
rect 4190 3880 4240 3905
rect 4190 3854 4196 3880
rect 4222 3854 4240 3880
rect 4190 3828 4240 3854
rect 4398 3876 4448 3905
rect 4398 3852 4412 3876
rect 4436 3852 4448 3876
rect 4398 3828 4448 3852
rect 4606 3881 4656 3905
rect 4606 3857 4621 3881
rect 4645 3857 4656 3881
rect 4606 3828 4656 3857
rect 4819 3876 4869 3905
rect 8459 3988 8509 4014
rect 8667 4036 8717 4065
rect 8667 4012 8681 4036
rect 8705 4012 8717 4036
rect 8667 3988 8717 4012
rect 8875 4041 8925 4065
rect 8875 4017 8890 4041
rect 8914 4017 8925 4041
rect 8875 3988 8925 4017
rect 9088 4036 9138 4065
rect 11023 4085 11073 4113
rect 11023 4065 11036 4085
rect 11056 4065 11073 4085
rect 9088 4016 9105 4036
rect 9125 4016 9138 4036
rect 9088 3988 9138 4016
rect 11023 4036 11073 4065
rect 11236 4084 11286 4113
rect 11236 4060 11247 4084
rect 11271 4060 11286 4084
rect 11236 4036 11286 4060
rect 11444 4089 11494 4113
rect 11444 4065 11456 4089
rect 11480 4065 11494 4089
rect 11444 4036 11494 4065
rect 11652 4087 11702 4113
rect 11652 4061 11670 4087
rect 11696 4061 11702 4087
rect 11652 4036 11702 4061
rect 13839 4069 13889 4094
rect 12035 4032 12085 4045
rect 12248 4032 12298 4045
rect 12456 4032 12506 4045
rect 12664 4032 12714 4045
rect 13839 4043 13845 4069
rect 13871 4043 13889 4069
rect 4819 3856 4836 3876
rect 4856 3856 4869 3876
rect 4819 3828 4869 3856
rect 361 3790 411 3803
rect 574 3790 624 3803
rect 782 3790 832 3803
rect 990 3790 1040 3803
rect 1374 3789 1424 3805
rect 1587 3789 1637 3805
rect 1795 3789 1845 3805
rect 2003 3789 2053 3805
rect 6655 3875 6705 3903
rect 6655 3855 6668 3875
rect 6688 3855 6705 3875
rect 6655 3826 6705 3855
rect 6868 3874 6918 3903
rect 6868 3850 6879 3874
rect 6903 3850 6918 3874
rect 6868 3826 6918 3850
rect 7076 3879 7126 3903
rect 7076 3855 7088 3879
rect 7112 3855 7126 3879
rect 7076 3826 7126 3855
rect 7284 3877 7334 3903
rect 11023 3978 11073 3994
rect 11236 3978 11286 3994
rect 11444 3978 11494 3994
rect 11652 3978 11702 3994
rect 9471 3926 9521 3942
rect 9679 3926 9729 3942
rect 9887 3926 9937 3942
rect 10100 3926 10150 3942
rect 13839 4017 13889 4043
rect 14047 4065 14097 4094
rect 14047 4041 14061 4065
rect 14085 4041 14097 4065
rect 14047 4017 14097 4041
rect 14255 4070 14305 4094
rect 14255 4046 14270 4070
rect 14294 4046 14305 4070
rect 14255 4017 14305 4046
rect 14468 4065 14518 4094
rect 14468 4045 14485 4065
rect 14505 4045 14518 4065
rect 14468 4017 14518 4045
rect 19120 4115 19170 4131
rect 19328 4115 19378 4131
rect 19536 4115 19586 4131
rect 19749 4115 19799 4131
rect 20133 4117 20183 4130
rect 20341 4117 20391 4130
rect 20549 4117 20599 4130
rect 20762 4117 20812 4130
rect 16304 4064 16354 4092
rect 16304 4044 16317 4064
rect 16337 4044 16354 4064
rect 7284 3851 7302 3877
rect 7328 3851 7334 3877
rect 8459 3875 8509 3888
rect 8667 3875 8717 3888
rect 8875 3875 8925 3888
rect 9088 3875 9138 3888
rect 7284 3826 7334 3851
rect 9471 3859 9521 3884
rect 9471 3833 9477 3859
rect 9503 3833 9521 3859
rect 9471 3807 9521 3833
rect 9679 3855 9729 3884
rect 9679 3831 9693 3855
rect 9717 3831 9729 3855
rect 9679 3807 9729 3831
rect 9887 3860 9937 3884
rect 9887 3836 9902 3860
rect 9926 3836 9937 3860
rect 9887 3807 9937 3836
rect 10100 3855 10150 3884
rect 12035 3904 12085 3932
rect 12035 3884 12048 3904
rect 12068 3884 12085 3904
rect 10100 3835 10117 3855
rect 10137 3835 10150 3855
rect 10100 3807 10150 3835
rect 12035 3855 12085 3884
rect 12248 3903 12298 3932
rect 12248 3879 12259 3903
rect 12283 3879 12298 3903
rect 12248 3855 12298 3879
rect 12456 3908 12506 3932
rect 12456 3884 12468 3908
rect 12492 3884 12506 3908
rect 12456 3855 12506 3884
rect 12664 3906 12714 3932
rect 16304 4015 16354 4044
rect 16517 4063 16567 4092
rect 16517 4039 16528 4063
rect 16552 4039 16567 4063
rect 16517 4015 16567 4039
rect 16725 4068 16775 4092
rect 16725 4044 16737 4068
rect 16761 4044 16775 4068
rect 16725 4015 16775 4044
rect 16933 4066 16983 4092
rect 16933 4040 16951 4066
rect 16977 4040 16983 4066
rect 16933 4015 16983 4040
rect 19120 4048 19170 4073
rect 17316 4011 17366 4024
rect 17529 4011 17579 4024
rect 17737 4011 17787 4024
rect 17945 4011 17995 4024
rect 19120 4022 19126 4048
rect 19152 4022 19170 4048
rect 14851 3955 14901 3971
rect 15059 3955 15109 3971
rect 15267 3955 15317 3971
rect 15480 3955 15530 3971
rect 16304 3957 16354 3973
rect 16517 3957 16567 3973
rect 16725 3957 16775 3973
rect 16933 3957 16983 3973
rect 12664 3880 12682 3906
rect 12708 3880 12714 3906
rect 13839 3904 13889 3917
rect 14047 3904 14097 3917
rect 14255 3904 14305 3917
rect 14468 3904 14518 3917
rect 12664 3855 12714 3880
rect 14851 3888 14901 3913
rect 14851 3862 14857 3888
rect 14883 3862 14901 3888
rect 5642 3769 5692 3782
rect 5855 3769 5905 3782
rect 6063 3769 6113 3782
rect 6271 3769 6321 3782
rect 3128 3708 3178 3724
rect 3336 3708 3386 3724
rect 3544 3708 3594 3724
rect 3757 3708 3807 3724
rect 4190 3715 4240 3728
rect 4398 3715 4448 3728
rect 4606 3715 4656 3728
rect 4819 3715 4869 3728
rect 361 3662 411 3690
rect 361 3642 374 3662
rect 394 3642 411 3662
rect 361 3613 411 3642
rect 574 3661 624 3690
rect 574 3637 585 3661
rect 609 3637 624 3661
rect 574 3613 624 3637
rect 782 3666 832 3690
rect 782 3642 794 3666
rect 818 3642 832 3666
rect 782 3613 832 3642
rect 990 3664 1040 3690
rect 990 3638 1008 3664
rect 1034 3638 1040 3664
rect 990 3613 1040 3638
rect 3128 3641 3178 3666
rect 3128 3615 3134 3641
rect 3160 3615 3178 3641
rect 3128 3589 3178 3615
rect 3336 3637 3386 3666
rect 3336 3613 3350 3637
rect 3374 3613 3386 3637
rect 3336 3589 3386 3613
rect 3544 3642 3594 3666
rect 3544 3618 3559 3642
rect 3583 3618 3594 3642
rect 3544 3589 3594 3618
rect 3757 3637 3807 3666
rect 3757 3617 3774 3637
rect 3794 3617 3807 3637
rect 3757 3589 3807 3617
rect 6655 3768 6705 3784
rect 6868 3768 6918 3784
rect 7076 3768 7126 3784
rect 7284 3768 7334 3784
rect 14851 3836 14901 3862
rect 15059 3884 15109 3913
rect 15059 3860 15073 3884
rect 15097 3860 15109 3884
rect 15059 3836 15109 3860
rect 15267 3889 15317 3913
rect 15267 3865 15282 3889
rect 15306 3865 15317 3889
rect 15267 3836 15317 3865
rect 15480 3884 15530 3913
rect 19120 3996 19170 4022
rect 19328 4044 19378 4073
rect 19328 4020 19342 4044
rect 19366 4020 19378 4044
rect 19328 3996 19378 4020
rect 19536 4049 19586 4073
rect 19536 4025 19551 4049
rect 19575 4025 19586 4049
rect 19536 3996 19586 4025
rect 19749 4044 19799 4073
rect 19749 4024 19766 4044
rect 19786 4024 19799 4044
rect 19749 3996 19799 4024
rect 15480 3864 15497 3884
rect 15517 3864 15530 3884
rect 15480 3836 15530 3864
rect 11022 3798 11072 3811
rect 11235 3798 11285 3811
rect 11443 3798 11493 3811
rect 11651 3798 11701 3811
rect 8409 3687 8459 3703
rect 8617 3687 8667 3703
rect 8825 3687 8875 3703
rect 9038 3687 9088 3703
rect 9471 3694 9521 3707
rect 9679 3694 9729 3707
rect 9887 3694 9937 3707
rect 10100 3694 10150 3707
rect 12035 3797 12085 3813
rect 12248 3797 12298 3813
rect 12456 3797 12506 3813
rect 12664 3797 12714 3813
rect 17316 3883 17366 3911
rect 17316 3863 17329 3883
rect 17349 3863 17366 3883
rect 17316 3834 17366 3863
rect 17529 3882 17579 3911
rect 17529 3858 17540 3882
rect 17564 3858 17579 3882
rect 17529 3834 17579 3858
rect 17737 3887 17787 3911
rect 17737 3863 17749 3887
rect 17773 3863 17787 3887
rect 17737 3834 17787 3863
rect 17945 3885 17995 3911
rect 20132 3934 20182 3950
rect 20340 3934 20390 3950
rect 20548 3934 20598 3950
rect 20761 3934 20811 3950
rect 17945 3859 17963 3885
rect 17989 3859 17995 3885
rect 19120 3883 19170 3896
rect 19328 3883 19378 3896
rect 19536 3883 19586 3896
rect 19749 3883 19799 3896
rect 17945 3834 17995 3859
rect 20132 3867 20182 3892
rect 20132 3841 20138 3867
rect 20164 3841 20182 3867
rect 20132 3815 20182 3841
rect 20340 3863 20390 3892
rect 20340 3839 20354 3863
rect 20378 3839 20390 3863
rect 20340 3815 20390 3839
rect 20548 3868 20598 3892
rect 20548 3844 20563 3868
rect 20587 3844 20598 3868
rect 20548 3815 20598 3844
rect 20761 3863 20811 3892
rect 20761 3843 20778 3863
rect 20798 3843 20811 3863
rect 20761 3815 20811 3843
rect 16303 3777 16353 3790
rect 16516 3777 16566 3790
rect 16724 3777 16774 3790
rect 16932 3777 16982 3790
rect 13789 3716 13839 3732
rect 13997 3716 14047 3732
rect 14205 3716 14255 3732
rect 14418 3716 14468 3732
rect 14851 3723 14901 3736
rect 15059 3723 15109 3736
rect 15267 3723 15317 3736
rect 15480 3723 15530 3736
rect 5642 3641 5692 3669
rect 361 3555 411 3571
rect 574 3555 624 3571
rect 782 3555 832 3571
rect 990 3555 1040 3571
rect 5642 3621 5655 3641
rect 5675 3621 5692 3641
rect 5642 3592 5692 3621
rect 5855 3640 5905 3669
rect 5855 3616 5866 3640
rect 5890 3616 5905 3640
rect 5855 3592 5905 3616
rect 6063 3645 6113 3669
rect 6063 3621 6075 3645
rect 6099 3621 6113 3645
rect 6063 3592 6113 3621
rect 6271 3643 6321 3669
rect 11022 3670 11072 3698
rect 6271 3617 6289 3643
rect 6315 3617 6321 3643
rect 6271 3592 6321 3617
rect 8409 3620 8459 3645
rect 8409 3594 8415 3620
rect 8441 3594 8459 3620
rect 8409 3568 8459 3594
rect 8617 3616 8667 3645
rect 8617 3592 8631 3616
rect 8655 3592 8667 3616
rect 8617 3568 8667 3592
rect 8825 3621 8875 3645
rect 8825 3597 8840 3621
rect 8864 3597 8875 3621
rect 8825 3568 8875 3597
rect 9038 3616 9088 3645
rect 9038 3596 9055 3616
rect 9075 3596 9088 3616
rect 9038 3568 9088 3596
rect 11022 3650 11035 3670
rect 11055 3650 11072 3670
rect 11022 3621 11072 3650
rect 11235 3669 11285 3698
rect 11235 3645 11246 3669
rect 11270 3645 11285 3669
rect 11235 3621 11285 3645
rect 11443 3674 11493 3698
rect 11443 3650 11455 3674
rect 11479 3650 11493 3674
rect 11443 3621 11493 3650
rect 11651 3672 11701 3698
rect 11651 3646 11669 3672
rect 11695 3646 11701 3672
rect 11651 3621 11701 3646
rect 13789 3649 13839 3674
rect 13789 3623 13795 3649
rect 13821 3623 13839 3649
rect 5642 3534 5692 3550
rect 5855 3534 5905 3550
rect 6063 3534 6113 3550
rect 6271 3534 6321 3550
rect 3128 3476 3178 3489
rect 3336 3476 3386 3489
rect 3544 3476 3594 3489
rect 3757 3476 3807 3489
rect 1429 3463 1479 3476
rect 1642 3463 1692 3476
rect 1850 3463 1900 3476
rect 2058 3463 2108 3476
rect 13789 3597 13839 3623
rect 13997 3645 14047 3674
rect 13997 3621 14011 3645
rect 14035 3621 14047 3645
rect 13997 3597 14047 3621
rect 14205 3650 14255 3674
rect 14205 3626 14220 3650
rect 14244 3626 14255 3650
rect 14205 3597 14255 3626
rect 14418 3645 14468 3674
rect 14418 3625 14435 3645
rect 14455 3625 14468 3645
rect 14418 3597 14468 3625
rect 17316 3776 17366 3792
rect 17529 3776 17579 3792
rect 17737 3776 17787 3792
rect 17945 3776 17995 3792
rect 19070 3695 19120 3711
rect 19278 3695 19328 3711
rect 19486 3695 19536 3711
rect 19699 3695 19749 3711
rect 20132 3702 20182 3715
rect 20340 3702 20390 3715
rect 20548 3702 20598 3715
rect 20761 3702 20811 3715
rect 16303 3649 16353 3677
rect 11022 3563 11072 3579
rect 11235 3563 11285 3579
rect 11443 3563 11493 3579
rect 11651 3563 11701 3579
rect 16303 3629 16316 3649
rect 16336 3629 16353 3649
rect 16303 3600 16353 3629
rect 16516 3648 16566 3677
rect 16516 3624 16527 3648
rect 16551 3624 16566 3648
rect 16516 3600 16566 3624
rect 16724 3653 16774 3677
rect 16724 3629 16736 3653
rect 16760 3629 16774 3653
rect 16724 3600 16774 3629
rect 16932 3651 16982 3677
rect 16932 3625 16950 3651
rect 16976 3625 16982 3651
rect 16932 3600 16982 3625
rect 19070 3628 19120 3653
rect 19070 3602 19076 3628
rect 19102 3602 19120 3628
rect 19070 3576 19120 3602
rect 19278 3624 19328 3653
rect 19278 3600 19292 3624
rect 19316 3600 19328 3624
rect 19278 3576 19328 3600
rect 19486 3629 19536 3653
rect 19486 3605 19501 3629
rect 19525 3605 19536 3629
rect 19486 3576 19536 3605
rect 19699 3624 19749 3653
rect 19699 3604 19716 3624
rect 19736 3604 19749 3624
rect 19699 3576 19749 3604
rect 16303 3542 16353 3558
rect 16516 3542 16566 3558
rect 16724 3542 16774 3558
rect 16932 3542 16982 3558
rect 13789 3484 13839 3497
rect 13997 3484 14047 3497
rect 14205 3484 14255 3497
rect 14418 3484 14468 3497
rect 12090 3471 12140 3484
rect 12303 3471 12353 3484
rect 12511 3471 12561 3484
rect 12719 3471 12769 3484
rect 8409 3455 8459 3468
rect 8617 3455 8667 3468
rect 8825 3455 8875 3468
rect 9038 3455 9088 3468
rect 6710 3442 6760 3455
rect 6923 3442 6973 3455
rect 7131 3442 7181 3455
rect 7339 3442 7389 3455
rect 4196 3381 4246 3397
rect 4404 3381 4454 3397
rect 4612 3381 4662 3397
rect 4825 3381 4875 3397
rect 1429 3335 1479 3363
rect 1429 3315 1442 3335
rect 1462 3315 1479 3335
rect 1429 3286 1479 3315
rect 1642 3334 1692 3363
rect 1642 3310 1653 3334
rect 1677 3310 1692 3334
rect 1642 3286 1692 3310
rect 1850 3339 1900 3363
rect 1850 3315 1862 3339
rect 1886 3315 1900 3339
rect 1850 3286 1900 3315
rect 2058 3337 2108 3363
rect 2058 3311 2076 3337
rect 2102 3311 2108 3337
rect 2058 3286 2108 3311
rect 4196 3314 4246 3339
rect 4196 3288 4202 3314
rect 4228 3288 4246 3314
rect 4196 3262 4246 3288
rect 4404 3310 4454 3339
rect 4404 3286 4418 3310
rect 4442 3286 4454 3310
rect 4404 3262 4454 3286
rect 4612 3315 4662 3339
rect 4612 3291 4627 3315
rect 4651 3291 4662 3315
rect 4612 3262 4662 3291
rect 4825 3310 4875 3339
rect 4825 3290 4842 3310
rect 4862 3290 4875 3310
rect 9477 3360 9527 3376
rect 9685 3360 9735 3376
rect 9893 3360 9943 3376
rect 10106 3360 10156 3376
rect 4825 3262 4875 3290
rect 367 3224 417 3237
rect 580 3224 630 3237
rect 788 3224 838 3237
rect 996 3224 1046 3237
rect 1429 3228 1479 3244
rect 1642 3228 1692 3244
rect 1850 3228 1900 3244
rect 2058 3228 2108 3244
rect 3183 3147 3233 3163
rect 3391 3147 3441 3163
rect 3599 3147 3649 3163
rect 3812 3147 3862 3163
rect 6710 3314 6760 3342
rect 6710 3294 6723 3314
rect 6743 3294 6760 3314
rect 6710 3265 6760 3294
rect 6923 3313 6973 3342
rect 6923 3289 6934 3313
rect 6958 3289 6973 3313
rect 6923 3265 6973 3289
rect 7131 3318 7181 3342
rect 7131 3294 7143 3318
rect 7167 3294 7181 3318
rect 7131 3265 7181 3294
rect 7339 3316 7389 3342
rect 19070 3463 19120 3476
rect 19278 3463 19328 3476
rect 19486 3463 19536 3476
rect 19699 3463 19749 3476
rect 17371 3450 17421 3463
rect 17584 3450 17634 3463
rect 17792 3450 17842 3463
rect 18000 3450 18050 3463
rect 14857 3389 14907 3405
rect 15065 3389 15115 3405
rect 15273 3389 15323 3405
rect 15486 3389 15536 3405
rect 7339 3290 7357 3316
rect 7383 3290 7389 3316
rect 7339 3265 7389 3290
rect 9477 3293 9527 3318
rect 9477 3267 9483 3293
rect 9509 3267 9527 3293
rect 9477 3241 9527 3267
rect 9685 3289 9735 3318
rect 9685 3265 9699 3289
rect 9723 3265 9735 3289
rect 9685 3241 9735 3265
rect 9893 3294 9943 3318
rect 9893 3270 9908 3294
rect 9932 3270 9943 3294
rect 9893 3241 9943 3270
rect 10106 3289 10156 3318
rect 10106 3269 10123 3289
rect 10143 3269 10156 3289
rect 12090 3343 12140 3371
rect 12090 3323 12103 3343
rect 12123 3323 12140 3343
rect 12090 3294 12140 3323
rect 12303 3342 12353 3371
rect 12303 3318 12314 3342
rect 12338 3318 12353 3342
rect 12303 3294 12353 3318
rect 12511 3347 12561 3371
rect 12511 3323 12523 3347
rect 12547 3323 12561 3347
rect 12511 3294 12561 3323
rect 12719 3345 12769 3371
rect 12719 3319 12737 3345
rect 12763 3319 12769 3345
rect 12719 3294 12769 3319
rect 14857 3322 14907 3347
rect 14857 3296 14863 3322
rect 14889 3296 14907 3322
rect 10106 3241 10156 3269
rect 14857 3270 14907 3296
rect 15065 3318 15115 3347
rect 15065 3294 15079 3318
rect 15103 3294 15115 3318
rect 15065 3270 15115 3294
rect 15273 3323 15323 3347
rect 15273 3299 15288 3323
rect 15312 3299 15323 3323
rect 15273 3270 15323 3299
rect 15486 3318 15536 3347
rect 15486 3298 15503 3318
rect 15523 3298 15536 3318
rect 20138 3368 20188 3384
rect 20346 3368 20396 3384
rect 20554 3368 20604 3384
rect 20767 3368 20817 3384
rect 15486 3270 15536 3298
rect 5648 3203 5698 3216
rect 5861 3203 5911 3216
rect 6069 3203 6119 3216
rect 6277 3203 6327 3216
rect 6710 3207 6760 3223
rect 6923 3207 6973 3223
rect 7131 3207 7181 3223
rect 7339 3207 7389 3223
rect 4196 3149 4246 3162
rect 4404 3149 4454 3162
rect 4612 3149 4662 3162
rect 4825 3149 4875 3162
rect 367 3096 417 3124
rect 367 3076 380 3096
rect 400 3076 417 3096
rect 367 3047 417 3076
rect 580 3095 630 3124
rect 580 3071 591 3095
rect 615 3071 630 3095
rect 580 3047 630 3071
rect 788 3100 838 3124
rect 788 3076 800 3100
rect 824 3076 838 3100
rect 788 3047 838 3076
rect 996 3098 1046 3124
rect 996 3072 1014 3098
rect 1040 3072 1046 3098
rect 996 3047 1046 3072
rect 3183 3080 3233 3105
rect 1379 3043 1429 3056
rect 1592 3043 1642 3056
rect 1800 3043 1850 3056
rect 2008 3043 2058 3056
rect 3183 3054 3189 3080
rect 3215 3054 3233 3080
rect 367 2989 417 3005
rect 580 2989 630 3005
rect 788 2989 838 3005
rect 996 2989 1046 3005
rect 3183 3028 3233 3054
rect 3391 3076 3441 3105
rect 3391 3052 3405 3076
rect 3429 3052 3441 3076
rect 3391 3028 3441 3052
rect 3599 3081 3649 3105
rect 3599 3057 3614 3081
rect 3638 3057 3649 3081
rect 3599 3028 3649 3057
rect 3812 3076 3862 3105
rect 3812 3056 3829 3076
rect 3849 3056 3862 3076
rect 3812 3028 3862 3056
rect 8464 3126 8514 3142
rect 8672 3126 8722 3142
rect 8880 3126 8930 3142
rect 9093 3126 9143 3142
rect 11028 3232 11078 3245
rect 11241 3232 11291 3245
rect 11449 3232 11499 3245
rect 11657 3232 11707 3245
rect 12090 3236 12140 3252
rect 12303 3236 12353 3252
rect 12511 3236 12561 3252
rect 12719 3236 12769 3252
rect 9477 3128 9527 3141
rect 9685 3128 9735 3141
rect 9893 3128 9943 3141
rect 10106 3128 10156 3141
rect 5648 3075 5698 3103
rect 5648 3055 5661 3075
rect 5681 3055 5698 3075
rect 1379 2915 1429 2943
rect 1379 2895 1392 2915
rect 1412 2895 1429 2915
rect 1379 2866 1429 2895
rect 1592 2914 1642 2943
rect 1592 2890 1603 2914
rect 1627 2890 1642 2914
rect 1592 2866 1642 2890
rect 1800 2919 1850 2943
rect 1800 2895 1812 2919
rect 1836 2895 1850 2919
rect 1800 2866 1850 2895
rect 2008 2917 2058 2943
rect 5648 3026 5698 3055
rect 5861 3074 5911 3103
rect 5861 3050 5872 3074
rect 5896 3050 5911 3074
rect 5861 3026 5911 3050
rect 6069 3079 6119 3103
rect 6069 3055 6081 3079
rect 6105 3055 6119 3079
rect 6069 3026 6119 3055
rect 6277 3077 6327 3103
rect 13844 3155 13894 3171
rect 14052 3155 14102 3171
rect 14260 3155 14310 3171
rect 14473 3155 14523 3171
rect 17371 3322 17421 3350
rect 17371 3302 17384 3322
rect 17404 3302 17421 3322
rect 17371 3273 17421 3302
rect 17584 3321 17634 3350
rect 17584 3297 17595 3321
rect 17619 3297 17634 3321
rect 17584 3273 17634 3297
rect 17792 3326 17842 3350
rect 17792 3302 17804 3326
rect 17828 3302 17842 3326
rect 17792 3273 17842 3302
rect 18000 3324 18050 3350
rect 18000 3298 18018 3324
rect 18044 3298 18050 3324
rect 18000 3273 18050 3298
rect 20138 3301 20188 3326
rect 20138 3275 20144 3301
rect 20170 3275 20188 3301
rect 20138 3249 20188 3275
rect 20346 3297 20396 3326
rect 20346 3273 20360 3297
rect 20384 3273 20396 3297
rect 20346 3249 20396 3273
rect 20554 3302 20604 3326
rect 20554 3278 20569 3302
rect 20593 3278 20604 3302
rect 20554 3249 20604 3278
rect 20767 3297 20817 3326
rect 20767 3277 20784 3297
rect 20804 3277 20817 3297
rect 20767 3249 20817 3277
rect 16309 3211 16359 3224
rect 16522 3211 16572 3224
rect 16730 3211 16780 3224
rect 16938 3211 16988 3224
rect 17371 3215 17421 3231
rect 17584 3215 17634 3231
rect 17792 3215 17842 3231
rect 18000 3215 18050 3231
rect 14857 3157 14907 3170
rect 15065 3157 15115 3170
rect 15273 3157 15323 3170
rect 15486 3157 15536 3170
rect 6277 3051 6295 3077
rect 6321 3051 6327 3077
rect 6277 3026 6327 3051
rect 8464 3059 8514 3084
rect 6660 3022 6710 3035
rect 6873 3022 6923 3035
rect 7081 3022 7131 3035
rect 7289 3022 7339 3035
rect 8464 3033 8470 3059
rect 8496 3033 8514 3059
rect 4195 2966 4245 2982
rect 4403 2966 4453 2982
rect 4611 2966 4661 2982
rect 4824 2966 4874 2982
rect 5648 2968 5698 2984
rect 5861 2968 5911 2984
rect 6069 2968 6119 2984
rect 6277 2968 6327 2984
rect 2008 2891 2026 2917
rect 2052 2891 2058 2917
rect 3183 2915 3233 2928
rect 3391 2915 3441 2928
rect 3599 2915 3649 2928
rect 3812 2915 3862 2928
rect 2008 2866 2058 2891
rect 4195 2899 4245 2924
rect 4195 2873 4201 2899
rect 4227 2873 4245 2899
rect 4195 2847 4245 2873
rect 4403 2895 4453 2924
rect 4403 2871 4417 2895
rect 4441 2871 4453 2895
rect 4403 2847 4453 2871
rect 4611 2900 4661 2924
rect 4611 2876 4626 2900
rect 4650 2876 4661 2900
rect 4611 2847 4661 2876
rect 4824 2895 4874 2924
rect 8464 3007 8514 3033
rect 8672 3055 8722 3084
rect 8672 3031 8686 3055
rect 8710 3031 8722 3055
rect 8672 3007 8722 3031
rect 8880 3060 8930 3084
rect 8880 3036 8895 3060
rect 8919 3036 8930 3060
rect 8880 3007 8930 3036
rect 9093 3055 9143 3084
rect 11028 3104 11078 3132
rect 11028 3084 11041 3104
rect 11061 3084 11078 3104
rect 9093 3035 9110 3055
rect 9130 3035 9143 3055
rect 9093 3007 9143 3035
rect 11028 3055 11078 3084
rect 11241 3103 11291 3132
rect 11241 3079 11252 3103
rect 11276 3079 11291 3103
rect 11241 3055 11291 3079
rect 11449 3108 11499 3132
rect 11449 3084 11461 3108
rect 11485 3084 11499 3108
rect 11449 3055 11499 3084
rect 11657 3106 11707 3132
rect 11657 3080 11675 3106
rect 11701 3080 11707 3106
rect 11657 3055 11707 3080
rect 13844 3088 13894 3113
rect 12040 3051 12090 3064
rect 12253 3051 12303 3064
rect 12461 3051 12511 3064
rect 12669 3051 12719 3064
rect 13844 3062 13850 3088
rect 13876 3062 13894 3088
rect 4824 2875 4841 2895
rect 4861 2875 4874 2895
rect 4824 2847 4874 2875
rect 366 2809 416 2822
rect 579 2809 629 2822
rect 787 2809 837 2822
rect 995 2809 1045 2822
rect 1379 2808 1429 2824
rect 1592 2808 1642 2824
rect 1800 2808 1850 2824
rect 2008 2808 2058 2824
rect 6660 2894 6710 2922
rect 6660 2874 6673 2894
rect 6693 2874 6710 2894
rect 6660 2845 6710 2874
rect 6873 2893 6923 2922
rect 6873 2869 6884 2893
rect 6908 2869 6923 2893
rect 6873 2845 6923 2869
rect 7081 2898 7131 2922
rect 7081 2874 7093 2898
rect 7117 2874 7131 2898
rect 7081 2845 7131 2874
rect 7289 2896 7339 2922
rect 11028 2997 11078 3013
rect 11241 2997 11291 3013
rect 11449 2997 11499 3013
rect 11657 2997 11707 3013
rect 9476 2945 9526 2961
rect 9684 2945 9734 2961
rect 9892 2945 9942 2961
rect 10105 2945 10155 2961
rect 13844 3036 13894 3062
rect 14052 3084 14102 3113
rect 14052 3060 14066 3084
rect 14090 3060 14102 3084
rect 14052 3036 14102 3060
rect 14260 3089 14310 3113
rect 14260 3065 14275 3089
rect 14299 3065 14310 3089
rect 14260 3036 14310 3065
rect 14473 3084 14523 3113
rect 14473 3064 14490 3084
rect 14510 3064 14523 3084
rect 14473 3036 14523 3064
rect 19125 3134 19175 3150
rect 19333 3134 19383 3150
rect 19541 3134 19591 3150
rect 19754 3134 19804 3150
rect 20138 3136 20188 3149
rect 20346 3136 20396 3149
rect 20554 3136 20604 3149
rect 20767 3136 20817 3149
rect 16309 3083 16359 3111
rect 16309 3063 16322 3083
rect 16342 3063 16359 3083
rect 7289 2870 7307 2896
rect 7333 2870 7339 2896
rect 8464 2894 8514 2907
rect 8672 2894 8722 2907
rect 8880 2894 8930 2907
rect 9093 2894 9143 2907
rect 7289 2845 7339 2870
rect 9476 2878 9526 2903
rect 9476 2852 9482 2878
rect 9508 2852 9526 2878
rect 9476 2826 9526 2852
rect 9684 2874 9734 2903
rect 9684 2850 9698 2874
rect 9722 2850 9734 2874
rect 9684 2826 9734 2850
rect 9892 2879 9942 2903
rect 9892 2855 9907 2879
rect 9931 2855 9942 2879
rect 9892 2826 9942 2855
rect 10105 2874 10155 2903
rect 12040 2923 12090 2951
rect 12040 2903 12053 2923
rect 12073 2903 12090 2923
rect 10105 2854 10122 2874
rect 10142 2854 10155 2874
rect 10105 2826 10155 2854
rect 12040 2874 12090 2903
rect 12253 2922 12303 2951
rect 12253 2898 12264 2922
rect 12288 2898 12303 2922
rect 12253 2874 12303 2898
rect 12461 2927 12511 2951
rect 12461 2903 12473 2927
rect 12497 2903 12511 2927
rect 12461 2874 12511 2903
rect 12669 2925 12719 2951
rect 16309 3034 16359 3063
rect 16522 3082 16572 3111
rect 16522 3058 16533 3082
rect 16557 3058 16572 3082
rect 16522 3034 16572 3058
rect 16730 3087 16780 3111
rect 16730 3063 16742 3087
rect 16766 3063 16780 3087
rect 16730 3034 16780 3063
rect 16938 3085 16988 3111
rect 16938 3059 16956 3085
rect 16982 3059 16988 3085
rect 16938 3034 16988 3059
rect 19125 3067 19175 3092
rect 17321 3030 17371 3043
rect 17534 3030 17584 3043
rect 17742 3030 17792 3043
rect 17950 3030 18000 3043
rect 19125 3041 19131 3067
rect 19157 3041 19175 3067
rect 14856 2974 14906 2990
rect 15064 2974 15114 2990
rect 15272 2974 15322 2990
rect 15485 2974 15535 2990
rect 16309 2976 16359 2992
rect 16522 2976 16572 2992
rect 16730 2976 16780 2992
rect 16938 2976 16988 2992
rect 12669 2899 12687 2925
rect 12713 2899 12719 2925
rect 13844 2923 13894 2936
rect 14052 2923 14102 2936
rect 14260 2923 14310 2936
rect 14473 2923 14523 2936
rect 12669 2874 12719 2899
rect 14856 2907 14906 2932
rect 14856 2881 14862 2907
rect 14888 2881 14906 2907
rect 5647 2788 5697 2801
rect 5860 2788 5910 2801
rect 6068 2788 6118 2801
rect 6276 2788 6326 2801
rect 4195 2734 4245 2747
rect 4403 2734 4453 2747
rect 4611 2734 4661 2747
rect 4824 2734 4874 2747
rect 366 2681 416 2709
rect 366 2661 379 2681
rect 399 2661 416 2681
rect 366 2632 416 2661
rect 579 2680 629 2709
rect 579 2656 590 2680
rect 614 2656 629 2680
rect 579 2632 629 2656
rect 787 2685 837 2709
rect 787 2661 799 2685
rect 823 2661 837 2685
rect 787 2632 837 2661
rect 995 2683 1045 2709
rect 995 2657 1013 2683
rect 1039 2657 1045 2683
rect 2975 2680 3025 2696
rect 3183 2680 3233 2696
rect 3391 2680 3441 2696
rect 3604 2680 3654 2696
rect 995 2632 1045 2657
rect 6660 2787 6710 2803
rect 6873 2787 6923 2803
rect 7081 2787 7131 2803
rect 7289 2787 7339 2803
rect 14856 2855 14906 2881
rect 15064 2903 15114 2932
rect 15064 2879 15078 2903
rect 15102 2879 15114 2903
rect 15064 2855 15114 2879
rect 15272 2908 15322 2932
rect 15272 2884 15287 2908
rect 15311 2884 15322 2908
rect 15272 2855 15322 2884
rect 15485 2903 15535 2932
rect 19125 3015 19175 3041
rect 19333 3063 19383 3092
rect 19333 3039 19347 3063
rect 19371 3039 19383 3063
rect 19333 3015 19383 3039
rect 19541 3068 19591 3092
rect 19541 3044 19556 3068
rect 19580 3044 19591 3068
rect 19541 3015 19591 3044
rect 19754 3063 19804 3092
rect 19754 3043 19771 3063
rect 19791 3043 19804 3063
rect 19754 3015 19804 3043
rect 15485 2883 15502 2903
rect 15522 2883 15535 2903
rect 15485 2855 15535 2883
rect 11027 2817 11077 2830
rect 11240 2817 11290 2830
rect 11448 2817 11498 2830
rect 11656 2817 11706 2830
rect 9476 2713 9526 2726
rect 9684 2713 9734 2726
rect 9892 2713 9942 2726
rect 10105 2713 10155 2726
rect 12040 2816 12090 2832
rect 12253 2816 12303 2832
rect 12461 2816 12511 2832
rect 12669 2816 12719 2832
rect 17321 2902 17371 2930
rect 17321 2882 17334 2902
rect 17354 2882 17371 2902
rect 17321 2853 17371 2882
rect 17534 2901 17584 2930
rect 17534 2877 17545 2901
rect 17569 2877 17584 2901
rect 17534 2853 17584 2877
rect 17742 2906 17792 2930
rect 17742 2882 17754 2906
rect 17778 2882 17792 2906
rect 17742 2853 17792 2882
rect 17950 2904 18000 2930
rect 20137 2953 20187 2969
rect 20345 2953 20395 2969
rect 20553 2953 20603 2969
rect 20766 2953 20816 2969
rect 17950 2878 17968 2904
rect 17994 2878 18000 2904
rect 19125 2902 19175 2915
rect 19333 2902 19383 2915
rect 19541 2902 19591 2915
rect 19754 2902 19804 2915
rect 17950 2853 18000 2878
rect 20137 2886 20187 2911
rect 20137 2860 20143 2886
rect 20169 2860 20187 2886
rect 20137 2834 20187 2860
rect 20345 2882 20395 2911
rect 20345 2858 20359 2882
rect 20383 2858 20395 2882
rect 20345 2834 20395 2858
rect 20553 2887 20603 2911
rect 20553 2863 20568 2887
rect 20592 2863 20603 2887
rect 20553 2834 20603 2863
rect 20766 2882 20816 2911
rect 20766 2862 20783 2882
rect 20803 2862 20816 2882
rect 20766 2834 20816 2862
rect 16308 2796 16358 2809
rect 16521 2796 16571 2809
rect 16729 2796 16779 2809
rect 16937 2796 16987 2809
rect 14856 2742 14906 2755
rect 15064 2742 15114 2755
rect 15272 2742 15322 2755
rect 15485 2742 15535 2755
rect 11027 2689 11077 2717
rect 2975 2613 3025 2638
rect 366 2574 416 2590
rect 579 2574 629 2590
rect 787 2574 837 2590
rect 995 2574 1045 2590
rect 2975 2587 2981 2613
rect 3007 2587 3025 2613
rect 2975 2561 3025 2587
rect 3183 2609 3233 2638
rect 3183 2585 3197 2609
rect 3221 2585 3233 2609
rect 3183 2561 3233 2585
rect 3391 2614 3441 2638
rect 3391 2590 3406 2614
rect 3430 2590 3441 2614
rect 3391 2561 3441 2590
rect 3604 2609 3654 2638
rect 5647 2660 5697 2688
rect 3604 2589 3621 2609
rect 3641 2589 3654 2609
rect 5647 2640 5660 2660
rect 5680 2640 5697 2660
rect 3604 2561 3654 2589
rect 5647 2611 5697 2640
rect 5860 2659 5910 2688
rect 5860 2635 5871 2659
rect 5895 2635 5910 2659
rect 5860 2611 5910 2635
rect 6068 2664 6118 2688
rect 6068 2640 6080 2664
rect 6104 2640 6118 2664
rect 6068 2611 6118 2640
rect 6276 2662 6326 2688
rect 6276 2636 6294 2662
rect 6320 2636 6326 2662
rect 8256 2659 8306 2675
rect 8464 2659 8514 2675
rect 8672 2659 8722 2675
rect 8885 2659 8935 2675
rect 6276 2611 6326 2636
rect 11027 2669 11040 2689
rect 11060 2669 11077 2689
rect 1594 2531 1644 2544
rect 1807 2531 1857 2544
rect 2015 2531 2065 2544
rect 2223 2531 2273 2544
rect 8256 2592 8306 2617
rect 5647 2553 5697 2569
rect 5860 2553 5910 2569
rect 6068 2553 6118 2569
rect 6276 2553 6326 2569
rect 8256 2566 8262 2592
rect 8288 2566 8306 2592
rect 8256 2540 8306 2566
rect 8464 2588 8514 2617
rect 8464 2564 8478 2588
rect 8502 2564 8514 2588
rect 8464 2540 8514 2564
rect 8672 2593 8722 2617
rect 8672 2569 8687 2593
rect 8711 2569 8722 2593
rect 8672 2540 8722 2569
rect 8885 2588 8935 2617
rect 11027 2640 11077 2669
rect 11240 2688 11290 2717
rect 11240 2664 11251 2688
rect 11275 2664 11290 2688
rect 11240 2640 11290 2664
rect 11448 2693 11498 2717
rect 11448 2669 11460 2693
rect 11484 2669 11498 2693
rect 11448 2640 11498 2669
rect 11656 2691 11706 2717
rect 11656 2665 11674 2691
rect 11700 2665 11706 2691
rect 13636 2688 13686 2704
rect 13844 2688 13894 2704
rect 14052 2688 14102 2704
rect 14265 2688 14315 2704
rect 11656 2640 11706 2665
rect 17321 2795 17371 2811
rect 17534 2795 17584 2811
rect 17742 2795 17792 2811
rect 17950 2795 18000 2811
rect 20137 2721 20187 2734
rect 20345 2721 20395 2734
rect 20553 2721 20603 2734
rect 20766 2721 20816 2734
rect 8885 2568 8902 2588
rect 8922 2568 8935 2588
rect 13636 2621 13686 2646
rect 11027 2582 11077 2598
rect 11240 2582 11290 2598
rect 11448 2582 11498 2598
rect 11656 2582 11706 2598
rect 13636 2595 13642 2621
rect 13668 2595 13686 2621
rect 8885 2540 8935 2568
rect 13636 2569 13686 2595
rect 13844 2617 13894 2646
rect 13844 2593 13858 2617
rect 13882 2593 13894 2617
rect 13844 2569 13894 2593
rect 14052 2622 14102 2646
rect 14052 2598 14067 2622
rect 14091 2598 14102 2622
rect 14052 2569 14102 2598
rect 14265 2617 14315 2646
rect 16308 2668 16358 2696
rect 14265 2597 14282 2617
rect 14302 2597 14315 2617
rect 16308 2648 16321 2668
rect 16341 2648 16358 2668
rect 14265 2569 14315 2597
rect 16308 2619 16358 2648
rect 16521 2667 16571 2696
rect 16521 2643 16532 2667
rect 16556 2643 16571 2667
rect 16521 2619 16571 2643
rect 16729 2672 16779 2696
rect 16729 2648 16741 2672
rect 16765 2648 16779 2672
rect 16729 2619 16779 2648
rect 16937 2670 16987 2696
rect 16937 2644 16955 2670
rect 16981 2644 16987 2670
rect 18917 2667 18967 2683
rect 19125 2667 19175 2683
rect 19333 2667 19383 2683
rect 19546 2667 19596 2683
rect 16937 2619 16987 2644
rect 6875 2510 6925 2523
rect 7088 2510 7138 2523
rect 7296 2510 7346 2523
rect 7504 2510 7554 2523
rect 2975 2448 3025 2461
rect 3183 2448 3233 2461
rect 3391 2448 3441 2461
rect 3604 2448 3654 2461
rect 1594 2403 1644 2431
rect 1594 2383 1607 2403
rect 1627 2383 1644 2403
rect 1594 2354 1644 2383
rect 1807 2402 1857 2431
rect 1807 2378 1818 2402
rect 1842 2378 1857 2402
rect 1807 2354 1857 2378
rect 2015 2407 2065 2431
rect 2015 2383 2027 2407
rect 2051 2383 2065 2407
rect 2015 2354 2065 2383
rect 2223 2405 2273 2431
rect 2223 2379 2241 2405
rect 2267 2379 2273 2405
rect 4203 2402 4253 2418
rect 4411 2402 4461 2418
rect 4619 2402 4669 2418
rect 4832 2402 4882 2418
rect 2223 2354 2273 2379
rect 12255 2539 12305 2552
rect 12468 2539 12518 2552
rect 12676 2539 12726 2552
rect 12884 2539 12934 2552
rect 8256 2427 8306 2440
rect 8464 2427 8514 2440
rect 8672 2427 8722 2440
rect 8885 2427 8935 2440
rect 18917 2600 18967 2625
rect 16308 2561 16358 2577
rect 16521 2561 16571 2577
rect 16729 2561 16779 2577
rect 16937 2561 16987 2577
rect 18917 2574 18923 2600
rect 18949 2574 18967 2600
rect 18917 2548 18967 2574
rect 19125 2596 19175 2625
rect 19125 2572 19139 2596
rect 19163 2572 19175 2596
rect 19125 2548 19175 2572
rect 19333 2601 19383 2625
rect 19333 2577 19348 2601
rect 19372 2577 19383 2601
rect 19333 2548 19383 2577
rect 19546 2596 19596 2625
rect 19546 2576 19563 2596
rect 19583 2576 19596 2596
rect 19546 2548 19596 2576
rect 17536 2518 17586 2531
rect 17749 2518 17799 2531
rect 17957 2518 18007 2531
rect 18165 2518 18215 2531
rect 13636 2456 13686 2469
rect 13844 2456 13894 2469
rect 14052 2456 14102 2469
rect 14265 2456 14315 2469
rect 4203 2335 4253 2360
rect 1594 2296 1644 2312
rect 1807 2296 1857 2312
rect 2015 2296 2065 2312
rect 2223 2296 2273 2312
rect 4203 2309 4209 2335
rect 4235 2309 4253 2335
rect 4203 2283 4253 2309
rect 4411 2331 4461 2360
rect 4411 2307 4425 2331
rect 4449 2307 4461 2331
rect 4411 2283 4461 2307
rect 4619 2336 4669 2360
rect 4619 2312 4634 2336
rect 4658 2312 4669 2336
rect 4619 2283 4669 2312
rect 4832 2331 4882 2360
rect 6875 2382 6925 2410
rect 4832 2311 4849 2331
rect 4869 2311 4882 2331
rect 6875 2362 6888 2382
rect 6908 2362 6925 2382
rect 4832 2283 4882 2311
rect 6875 2333 6925 2362
rect 7088 2381 7138 2410
rect 7088 2357 7099 2381
rect 7123 2357 7138 2381
rect 7088 2333 7138 2357
rect 7296 2386 7346 2410
rect 7296 2362 7308 2386
rect 7332 2362 7346 2386
rect 7296 2333 7346 2362
rect 7504 2384 7554 2410
rect 12255 2411 12305 2439
rect 7504 2358 7522 2384
rect 7548 2358 7554 2384
rect 9484 2381 9534 2397
rect 9692 2381 9742 2397
rect 9900 2381 9950 2397
rect 10113 2381 10163 2397
rect 7504 2333 7554 2358
rect 12255 2391 12268 2411
rect 12288 2391 12305 2411
rect 374 2245 424 2258
rect 587 2245 637 2258
rect 795 2245 845 2258
rect 1003 2245 1053 2258
rect 3190 2168 3240 2184
rect 3398 2168 3448 2184
rect 3606 2168 3656 2184
rect 3819 2168 3869 2184
rect 9484 2314 9534 2339
rect 6875 2275 6925 2291
rect 7088 2275 7138 2291
rect 7296 2275 7346 2291
rect 7504 2275 7554 2291
rect 9484 2288 9490 2314
rect 9516 2288 9534 2314
rect 9484 2262 9534 2288
rect 9692 2310 9742 2339
rect 9692 2286 9706 2310
rect 9730 2286 9742 2310
rect 9692 2262 9742 2286
rect 9900 2315 9950 2339
rect 9900 2291 9915 2315
rect 9939 2291 9950 2315
rect 9900 2262 9950 2291
rect 10113 2310 10163 2339
rect 12255 2362 12305 2391
rect 12468 2410 12518 2439
rect 12468 2386 12479 2410
rect 12503 2386 12518 2410
rect 12468 2362 12518 2386
rect 12676 2415 12726 2439
rect 12676 2391 12688 2415
rect 12712 2391 12726 2415
rect 12676 2362 12726 2391
rect 12884 2413 12934 2439
rect 12884 2387 12902 2413
rect 12928 2387 12934 2413
rect 14864 2410 14914 2426
rect 15072 2410 15122 2426
rect 15280 2410 15330 2426
rect 15493 2410 15543 2426
rect 12884 2362 12934 2387
rect 18917 2435 18967 2448
rect 19125 2435 19175 2448
rect 19333 2435 19383 2448
rect 19546 2435 19596 2448
rect 10113 2290 10130 2310
rect 10150 2290 10163 2310
rect 14864 2343 14914 2368
rect 12255 2304 12305 2320
rect 12468 2304 12518 2320
rect 12676 2304 12726 2320
rect 12884 2304 12934 2320
rect 14864 2317 14870 2343
rect 14896 2317 14914 2343
rect 14864 2291 14914 2317
rect 15072 2339 15122 2368
rect 15072 2315 15086 2339
rect 15110 2315 15122 2339
rect 15072 2291 15122 2315
rect 15280 2344 15330 2368
rect 15280 2320 15295 2344
rect 15319 2320 15330 2344
rect 15280 2291 15330 2320
rect 15493 2339 15543 2368
rect 17536 2390 17586 2418
rect 15493 2319 15510 2339
rect 15530 2319 15543 2339
rect 17536 2370 17549 2390
rect 17569 2370 17586 2390
rect 15493 2291 15543 2319
rect 17536 2341 17586 2370
rect 17749 2389 17799 2418
rect 17749 2365 17760 2389
rect 17784 2365 17799 2389
rect 17749 2341 17799 2365
rect 17957 2394 18007 2418
rect 17957 2370 17969 2394
rect 17993 2370 18007 2394
rect 17957 2341 18007 2370
rect 18165 2392 18215 2418
rect 18165 2366 18183 2392
rect 18209 2366 18215 2392
rect 20145 2389 20195 2405
rect 20353 2389 20403 2405
rect 20561 2389 20611 2405
rect 20774 2389 20824 2405
rect 18165 2341 18215 2366
rect 10113 2262 10163 2290
rect 5655 2224 5705 2237
rect 5868 2224 5918 2237
rect 6076 2224 6126 2237
rect 6284 2224 6334 2237
rect 4203 2170 4253 2183
rect 4411 2170 4461 2183
rect 4619 2170 4669 2183
rect 4832 2170 4882 2183
rect 374 2117 424 2145
rect 374 2097 387 2117
rect 407 2097 424 2117
rect 374 2068 424 2097
rect 587 2116 637 2145
rect 587 2092 598 2116
rect 622 2092 637 2116
rect 587 2068 637 2092
rect 795 2121 845 2145
rect 795 2097 807 2121
rect 831 2097 845 2121
rect 795 2068 845 2097
rect 1003 2119 1053 2145
rect 1003 2093 1021 2119
rect 1047 2093 1053 2119
rect 1003 2068 1053 2093
rect 3190 2101 3240 2126
rect 1386 2064 1436 2077
rect 1599 2064 1649 2077
rect 1807 2064 1857 2077
rect 2015 2064 2065 2077
rect 3190 2075 3196 2101
rect 3222 2075 3240 2101
rect 374 2010 424 2026
rect 587 2010 637 2026
rect 795 2010 845 2026
rect 1003 2010 1053 2026
rect 3190 2049 3240 2075
rect 3398 2097 3448 2126
rect 3398 2073 3412 2097
rect 3436 2073 3448 2097
rect 3398 2049 3448 2073
rect 3606 2102 3656 2126
rect 3606 2078 3621 2102
rect 3645 2078 3656 2102
rect 3606 2049 3656 2078
rect 3819 2097 3869 2126
rect 3819 2077 3836 2097
rect 3856 2077 3869 2097
rect 3819 2049 3869 2077
rect 8471 2147 8521 2163
rect 8679 2147 8729 2163
rect 8887 2147 8937 2163
rect 9100 2147 9150 2163
rect 11035 2253 11085 2266
rect 11248 2253 11298 2266
rect 11456 2253 11506 2266
rect 11664 2253 11714 2266
rect 9484 2149 9534 2162
rect 9692 2149 9742 2162
rect 9900 2149 9950 2162
rect 10113 2149 10163 2162
rect 5655 2096 5705 2124
rect 5655 2076 5668 2096
rect 5688 2076 5705 2096
rect 1386 1936 1436 1964
rect 1386 1916 1399 1936
rect 1419 1916 1436 1936
rect 1386 1887 1436 1916
rect 1599 1935 1649 1964
rect 1599 1911 1610 1935
rect 1634 1911 1649 1935
rect 1599 1887 1649 1911
rect 1807 1940 1857 1964
rect 1807 1916 1819 1940
rect 1843 1916 1857 1940
rect 1807 1887 1857 1916
rect 2015 1938 2065 1964
rect 5655 2047 5705 2076
rect 5868 2095 5918 2124
rect 5868 2071 5879 2095
rect 5903 2071 5918 2095
rect 5868 2047 5918 2071
rect 6076 2100 6126 2124
rect 6076 2076 6088 2100
rect 6112 2076 6126 2100
rect 6076 2047 6126 2076
rect 6284 2098 6334 2124
rect 13851 2176 13901 2192
rect 14059 2176 14109 2192
rect 14267 2176 14317 2192
rect 14480 2176 14530 2192
rect 20145 2322 20195 2347
rect 17536 2283 17586 2299
rect 17749 2283 17799 2299
rect 17957 2283 18007 2299
rect 18165 2283 18215 2299
rect 20145 2296 20151 2322
rect 20177 2296 20195 2322
rect 20145 2270 20195 2296
rect 20353 2318 20403 2347
rect 20353 2294 20367 2318
rect 20391 2294 20403 2318
rect 20353 2270 20403 2294
rect 20561 2323 20611 2347
rect 20561 2299 20576 2323
rect 20600 2299 20611 2323
rect 20561 2270 20611 2299
rect 20774 2318 20824 2347
rect 20774 2298 20791 2318
rect 20811 2298 20824 2318
rect 20774 2270 20824 2298
rect 16316 2232 16366 2245
rect 16529 2232 16579 2245
rect 16737 2232 16787 2245
rect 16945 2232 16995 2245
rect 14864 2178 14914 2191
rect 15072 2178 15122 2191
rect 15280 2178 15330 2191
rect 15493 2178 15543 2191
rect 6284 2072 6302 2098
rect 6328 2072 6334 2098
rect 6284 2047 6334 2072
rect 8471 2080 8521 2105
rect 6667 2043 6717 2056
rect 6880 2043 6930 2056
rect 7088 2043 7138 2056
rect 7296 2043 7346 2056
rect 8471 2054 8477 2080
rect 8503 2054 8521 2080
rect 4202 1987 4252 2003
rect 4410 1987 4460 2003
rect 4618 1987 4668 2003
rect 4831 1987 4881 2003
rect 5655 1989 5705 2005
rect 5868 1989 5918 2005
rect 6076 1989 6126 2005
rect 6284 1989 6334 2005
rect 2015 1912 2033 1938
rect 2059 1912 2065 1938
rect 3190 1936 3240 1949
rect 3398 1936 3448 1949
rect 3606 1936 3656 1949
rect 3819 1936 3869 1949
rect 2015 1887 2065 1912
rect 4202 1920 4252 1945
rect 4202 1894 4208 1920
rect 4234 1894 4252 1920
rect 4202 1868 4252 1894
rect 4410 1916 4460 1945
rect 4410 1892 4424 1916
rect 4448 1892 4460 1916
rect 4410 1868 4460 1892
rect 4618 1921 4668 1945
rect 4618 1897 4633 1921
rect 4657 1897 4668 1921
rect 4618 1868 4668 1897
rect 4831 1916 4881 1945
rect 8471 2028 8521 2054
rect 8679 2076 8729 2105
rect 8679 2052 8693 2076
rect 8717 2052 8729 2076
rect 8679 2028 8729 2052
rect 8887 2081 8937 2105
rect 8887 2057 8902 2081
rect 8926 2057 8937 2081
rect 8887 2028 8937 2057
rect 9100 2076 9150 2105
rect 11035 2125 11085 2153
rect 11035 2105 11048 2125
rect 11068 2105 11085 2125
rect 9100 2056 9117 2076
rect 9137 2056 9150 2076
rect 9100 2028 9150 2056
rect 11035 2076 11085 2105
rect 11248 2124 11298 2153
rect 11248 2100 11259 2124
rect 11283 2100 11298 2124
rect 11248 2076 11298 2100
rect 11456 2129 11506 2153
rect 11456 2105 11468 2129
rect 11492 2105 11506 2129
rect 11456 2076 11506 2105
rect 11664 2127 11714 2153
rect 11664 2101 11682 2127
rect 11708 2101 11714 2127
rect 11664 2076 11714 2101
rect 13851 2109 13901 2134
rect 12047 2072 12097 2085
rect 12260 2072 12310 2085
rect 12468 2072 12518 2085
rect 12676 2072 12726 2085
rect 13851 2083 13857 2109
rect 13883 2083 13901 2109
rect 4831 1896 4848 1916
rect 4868 1896 4881 1916
rect 4831 1868 4881 1896
rect 373 1830 423 1843
rect 586 1830 636 1843
rect 794 1830 844 1843
rect 1002 1830 1052 1843
rect 1386 1829 1436 1845
rect 1599 1829 1649 1845
rect 1807 1829 1857 1845
rect 2015 1829 2065 1845
rect 6667 1915 6717 1943
rect 6667 1895 6680 1915
rect 6700 1895 6717 1915
rect 6667 1866 6717 1895
rect 6880 1914 6930 1943
rect 6880 1890 6891 1914
rect 6915 1890 6930 1914
rect 6880 1866 6930 1890
rect 7088 1919 7138 1943
rect 7088 1895 7100 1919
rect 7124 1895 7138 1919
rect 7088 1866 7138 1895
rect 7296 1917 7346 1943
rect 11035 2018 11085 2034
rect 11248 2018 11298 2034
rect 11456 2018 11506 2034
rect 11664 2018 11714 2034
rect 9483 1966 9533 1982
rect 9691 1966 9741 1982
rect 9899 1966 9949 1982
rect 10112 1966 10162 1982
rect 13851 2057 13901 2083
rect 14059 2105 14109 2134
rect 14059 2081 14073 2105
rect 14097 2081 14109 2105
rect 14059 2057 14109 2081
rect 14267 2110 14317 2134
rect 14267 2086 14282 2110
rect 14306 2086 14317 2110
rect 14267 2057 14317 2086
rect 14480 2105 14530 2134
rect 14480 2085 14497 2105
rect 14517 2085 14530 2105
rect 14480 2057 14530 2085
rect 19132 2155 19182 2171
rect 19340 2155 19390 2171
rect 19548 2155 19598 2171
rect 19761 2155 19811 2171
rect 20145 2157 20195 2170
rect 20353 2157 20403 2170
rect 20561 2157 20611 2170
rect 20774 2157 20824 2170
rect 16316 2104 16366 2132
rect 16316 2084 16329 2104
rect 16349 2084 16366 2104
rect 7296 1891 7314 1917
rect 7340 1891 7346 1917
rect 8471 1915 8521 1928
rect 8679 1915 8729 1928
rect 8887 1915 8937 1928
rect 9100 1915 9150 1928
rect 7296 1866 7346 1891
rect 9483 1899 9533 1924
rect 9483 1873 9489 1899
rect 9515 1873 9533 1899
rect 9483 1847 9533 1873
rect 9691 1895 9741 1924
rect 9691 1871 9705 1895
rect 9729 1871 9741 1895
rect 9691 1847 9741 1871
rect 9899 1900 9949 1924
rect 9899 1876 9914 1900
rect 9938 1876 9949 1900
rect 9899 1847 9949 1876
rect 10112 1895 10162 1924
rect 12047 1944 12097 1972
rect 12047 1924 12060 1944
rect 12080 1924 12097 1944
rect 10112 1875 10129 1895
rect 10149 1875 10162 1895
rect 10112 1847 10162 1875
rect 12047 1895 12097 1924
rect 12260 1943 12310 1972
rect 12260 1919 12271 1943
rect 12295 1919 12310 1943
rect 12260 1895 12310 1919
rect 12468 1948 12518 1972
rect 12468 1924 12480 1948
rect 12504 1924 12518 1948
rect 12468 1895 12518 1924
rect 12676 1946 12726 1972
rect 16316 2055 16366 2084
rect 16529 2103 16579 2132
rect 16529 2079 16540 2103
rect 16564 2079 16579 2103
rect 16529 2055 16579 2079
rect 16737 2108 16787 2132
rect 16737 2084 16749 2108
rect 16773 2084 16787 2108
rect 16737 2055 16787 2084
rect 16945 2106 16995 2132
rect 16945 2080 16963 2106
rect 16989 2080 16995 2106
rect 16945 2055 16995 2080
rect 19132 2088 19182 2113
rect 17328 2051 17378 2064
rect 17541 2051 17591 2064
rect 17749 2051 17799 2064
rect 17957 2051 18007 2064
rect 19132 2062 19138 2088
rect 19164 2062 19182 2088
rect 14863 1995 14913 2011
rect 15071 1995 15121 2011
rect 15279 1995 15329 2011
rect 15492 1995 15542 2011
rect 16316 1997 16366 2013
rect 16529 1997 16579 2013
rect 16737 1997 16787 2013
rect 16945 1997 16995 2013
rect 12676 1920 12694 1946
rect 12720 1920 12726 1946
rect 13851 1944 13901 1957
rect 14059 1944 14109 1957
rect 14267 1944 14317 1957
rect 14480 1944 14530 1957
rect 12676 1895 12726 1920
rect 14863 1928 14913 1953
rect 14863 1902 14869 1928
rect 14895 1902 14913 1928
rect 5654 1809 5704 1822
rect 5867 1809 5917 1822
rect 6075 1809 6125 1822
rect 6283 1809 6333 1822
rect 3140 1748 3190 1764
rect 3348 1748 3398 1764
rect 3556 1748 3606 1764
rect 3769 1748 3819 1764
rect 4202 1755 4252 1768
rect 4410 1755 4460 1768
rect 4618 1755 4668 1768
rect 4831 1755 4881 1768
rect 373 1702 423 1730
rect 373 1682 386 1702
rect 406 1682 423 1702
rect 373 1653 423 1682
rect 586 1701 636 1730
rect 586 1677 597 1701
rect 621 1677 636 1701
rect 586 1653 636 1677
rect 794 1706 844 1730
rect 794 1682 806 1706
rect 830 1682 844 1706
rect 794 1653 844 1682
rect 1002 1704 1052 1730
rect 1002 1678 1020 1704
rect 1046 1678 1052 1704
rect 1002 1653 1052 1678
rect 3140 1681 3190 1706
rect 3140 1655 3146 1681
rect 3172 1655 3190 1681
rect 3140 1629 3190 1655
rect 3348 1677 3398 1706
rect 3348 1653 3362 1677
rect 3386 1653 3398 1677
rect 3348 1629 3398 1653
rect 3556 1682 3606 1706
rect 3556 1658 3571 1682
rect 3595 1658 3606 1682
rect 3556 1629 3606 1658
rect 3769 1677 3819 1706
rect 3769 1657 3786 1677
rect 3806 1657 3819 1677
rect 3769 1629 3819 1657
rect 6667 1808 6717 1824
rect 6880 1808 6930 1824
rect 7088 1808 7138 1824
rect 7296 1808 7346 1824
rect 14863 1876 14913 1902
rect 15071 1924 15121 1953
rect 15071 1900 15085 1924
rect 15109 1900 15121 1924
rect 15071 1876 15121 1900
rect 15279 1929 15329 1953
rect 15279 1905 15294 1929
rect 15318 1905 15329 1929
rect 15279 1876 15329 1905
rect 15492 1924 15542 1953
rect 19132 2036 19182 2062
rect 19340 2084 19390 2113
rect 19340 2060 19354 2084
rect 19378 2060 19390 2084
rect 19340 2036 19390 2060
rect 19548 2089 19598 2113
rect 19548 2065 19563 2089
rect 19587 2065 19598 2089
rect 19548 2036 19598 2065
rect 19761 2084 19811 2113
rect 19761 2064 19778 2084
rect 19798 2064 19811 2084
rect 19761 2036 19811 2064
rect 15492 1904 15509 1924
rect 15529 1904 15542 1924
rect 15492 1876 15542 1904
rect 11034 1838 11084 1851
rect 11247 1838 11297 1851
rect 11455 1838 11505 1851
rect 11663 1838 11713 1851
rect 8421 1727 8471 1743
rect 8629 1727 8679 1743
rect 8837 1727 8887 1743
rect 9050 1727 9100 1743
rect 9483 1734 9533 1747
rect 9691 1734 9741 1747
rect 9899 1734 9949 1747
rect 10112 1734 10162 1747
rect 12047 1837 12097 1853
rect 12260 1837 12310 1853
rect 12468 1837 12518 1853
rect 12676 1837 12726 1853
rect 17328 1923 17378 1951
rect 17328 1903 17341 1923
rect 17361 1903 17378 1923
rect 17328 1874 17378 1903
rect 17541 1922 17591 1951
rect 17541 1898 17552 1922
rect 17576 1898 17591 1922
rect 17541 1874 17591 1898
rect 17749 1927 17799 1951
rect 17749 1903 17761 1927
rect 17785 1903 17799 1927
rect 17749 1874 17799 1903
rect 17957 1925 18007 1951
rect 20144 1974 20194 1990
rect 20352 1974 20402 1990
rect 20560 1974 20610 1990
rect 20773 1974 20823 1990
rect 17957 1899 17975 1925
rect 18001 1899 18007 1925
rect 19132 1923 19182 1936
rect 19340 1923 19390 1936
rect 19548 1923 19598 1936
rect 19761 1923 19811 1936
rect 17957 1874 18007 1899
rect 20144 1907 20194 1932
rect 20144 1881 20150 1907
rect 20176 1881 20194 1907
rect 20144 1855 20194 1881
rect 20352 1903 20402 1932
rect 20352 1879 20366 1903
rect 20390 1879 20402 1903
rect 20352 1855 20402 1879
rect 20560 1908 20610 1932
rect 20560 1884 20575 1908
rect 20599 1884 20610 1908
rect 20560 1855 20610 1884
rect 20773 1903 20823 1932
rect 20773 1883 20790 1903
rect 20810 1883 20823 1903
rect 20773 1855 20823 1883
rect 16315 1817 16365 1830
rect 16528 1817 16578 1830
rect 16736 1817 16786 1830
rect 16944 1817 16994 1830
rect 13801 1756 13851 1772
rect 14009 1756 14059 1772
rect 14217 1756 14267 1772
rect 14430 1756 14480 1772
rect 14863 1763 14913 1776
rect 15071 1763 15121 1776
rect 15279 1763 15329 1776
rect 15492 1763 15542 1776
rect 5654 1681 5704 1709
rect 373 1595 423 1611
rect 586 1595 636 1611
rect 794 1595 844 1611
rect 1002 1595 1052 1611
rect 5654 1661 5667 1681
rect 5687 1661 5704 1681
rect 5654 1632 5704 1661
rect 5867 1680 5917 1709
rect 5867 1656 5878 1680
rect 5902 1656 5917 1680
rect 5867 1632 5917 1656
rect 6075 1685 6125 1709
rect 6075 1661 6087 1685
rect 6111 1661 6125 1685
rect 6075 1632 6125 1661
rect 6283 1683 6333 1709
rect 11034 1710 11084 1738
rect 6283 1657 6301 1683
rect 6327 1657 6333 1683
rect 6283 1632 6333 1657
rect 8421 1660 8471 1685
rect 8421 1634 8427 1660
rect 8453 1634 8471 1660
rect 8421 1608 8471 1634
rect 8629 1656 8679 1685
rect 8629 1632 8643 1656
rect 8667 1632 8679 1656
rect 8629 1608 8679 1632
rect 8837 1661 8887 1685
rect 8837 1637 8852 1661
rect 8876 1637 8887 1661
rect 8837 1608 8887 1637
rect 9050 1656 9100 1685
rect 9050 1636 9067 1656
rect 9087 1636 9100 1656
rect 9050 1608 9100 1636
rect 11034 1690 11047 1710
rect 11067 1690 11084 1710
rect 11034 1661 11084 1690
rect 11247 1709 11297 1738
rect 11247 1685 11258 1709
rect 11282 1685 11297 1709
rect 11247 1661 11297 1685
rect 11455 1714 11505 1738
rect 11455 1690 11467 1714
rect 11491 1690 11505 1714
rect 11455 1661 11505 1690
rect 11663 1712 11713 1738
rect 11663 1686 11681 1712
rect 11707 1686 11713 1712
rect 11663 1661 11713 1686
rect 13801 1689 13851 1714
rect 13801 1663 13807 1689
rect 13833 1663 13851 1689
rect 5654 1574 5704 1590
rect 5867 1574 5917 1590
rect 6075 1574 6125 1590
rect 6283 1574 6333 1590
rect 3140 1516 3190 1529
rect 3348 1516 3398 1529
rect 3556 1516 3606 1529
rect 3769 1516 3819 1529
rect 1441 1503 1491 1516
rect 1654 1503 1704 1516
rect 1862 1503 1912 1516
rect 2070 1503 2120 1516
rect 13801 1637 13851 1663
rect 14009 1685 14059 1714
rect 14009 1661 14023 1685
rect 14047 1661 14059 1685
rect 14009 1637 14059 1661
rect 14217 1690 14267 1714
rect 14217 1666 14232 1690
rect 14256 1666 14267 1690
rect 14217 1637 14267 1666
rect 14430 1685 14480 1714
rect 14430 1665 14447 1685
rect 14467 1665 14480 1685
rect 14430 1637 14480 1665
rect 17328 1816 17378 1832
rect 17541 1816 17591 1832
rect 17749 1816 17799 1832
rect 17957 1816 18007 1832
rect 19082 1735 19132 1751
rect 19290 1735 19340 1751
rect 19498 1735 19548 1751
rect 19711 1735 19761 1751
rect 20144 1742 20194 1755
rect 20352 1742 20402 1755
rect 20560 1742 20610 1755
rect 20773 1742 20823 1755
rect 16315 1689 16365 1717
rect 11034 1603 11084 1619
rect 11247 1603 11297 1619
rect 11455 1603 11505 1619
rect 11663 1603 11713 1619
rect 16315 1669 16328 1689
rect 16348 1669 16365 1689
rect 16315 1640 16365 1669
rect 16528 1688 16578 1717
rect 16528 1664 16539 1688
rect 16563 1664 16578 1688
rect 16528 1640 16578 1664
rect 16736 1693 16786 1717
rect 16736 1669 16748 1693
rect 16772 1669 16786 1693
rect 16736 1640 16786 1669
rect 16944 1691 16994 1717
rect 16944 1665 16962 1691
rect 16988 1665 16994 1691
rect 16944 1640 16994 1665
rect 19082 1668 19132 1693
rect 19082 1642 19088 1668
rect 19114 1642 19132 1668
rect 19082 1616 19132 1642
rect 19290 1664 19340 1693
rect 19290 1640 19304 1664
rect 19328 1640 19340 1664
rect 19290 1616 19340 1640
rect 19498 1669 19548 1693
rect 19498 1645 19513 1669
rect 19537 1645 19548 1669
rect 19498 1616 19548 1645
rect 19711 1664 19761 1693
rect 19711 1644 19728 1664
rect 19748 1644 19761 1664
rect 19711 1616 19761 1644
rect 16315 1582 16365 1598
rect 16528 1582 16578 1598
rect 16736 1582 16786 1598
rect 16944 1582 16994 1598
rect 13801 1524 13851 1537
rect 14009 1524 14059 1537
rect 14217 1524 14267 1537
rect 14430 1524 14480 1537
rect 12102 1511 12152 1524
rect 12315 1511 12365 1524
rect 12523 1511 12573 1524
rect 12731 1511 12781 1524
rect 8421 1495 8471 1508
rect 8629 1495 8679 1508
rect 8837 1495 8887 1508
rect 9050 1495 9100 1508
rect 6722 1482 6772 1495
rect 6935 1482 6985 1495
rect 7143 1482 7193 1495
rect 7351 1482 7401 1495
rect 4208 1421 4258 1437
rect 4416 1421 4466 1437
rect 4624 1421 4674 1437
rect 4837 1421 4887 1437
rect 1441 1375 1491 1403
rect 1441 1355 1454 1375
rect 1474 1355 1491 1375
rect 1441 1326 1491 1355
rect 1654 1374 1704 1403
rect 1654 1350 1665 1374
rect 1689 1350 1704 1374
rect 1654 1326 1704 1350
rect 1862 1379 1912 1403
rect 1862 1355 1874 1379
rect 1898 1355 1912 1379
rect 1862 1326 1912 1355
rect 2070 1377 2120 1403
rect 2070 1351 2088 1377
rect 2114 1351 2120 1377
rect 2070 1326 2120 1351
rect 4208 1354 4258 1379
rect 4208 1328 4214 1354
rect 4240 1328 4258 1354
rect 4208 1302 4258 1328
rect 4416 1350 4466 1379
rect 4416 1326 4430 1350
rect 4454 1326 4466 1350
rect 4416 1302 4466 1326
rect 4624 1355 4674 1379
rect 4624 1331 4639 1355
rect 4663 1331 4674 1355
rect 4624 1302 4674 1331
rect 4837 1350 4887 1379
rect 4837 1330 4854 1350
rect 4874 1330 4887 1350
rect 9489 1400 9539 1416
rect 9697 1400 9747 1416
rect 9905 1400 9955 1416
rect 10118 1400 10168 1416
rect 4837 1302 4887 1330
rect 379 1264 429 1277
rect 592 1264 642 1277
rect 800 1264 850 1277
rect 1008 1264 1058 1277
rect 1441 1268 1491 1284
rect 1654 1268 1704 1284
rect 1862 1268 1912 1284
rect 2070 1268 2120 1284
rect 3195 1187 3245 1203
rect 3403 1187 3453 1203
rect 3611 1187 3661 1203
rect 3824 1187 3874 1203
rect 6722 1354 6772 1382
rect 6722 1334 6735 1354
rect 6755 1334 6772 1354
rect 6722 1305 6772 1334
rect 6935 1353 6985 1382
rect 6935 1329 6946 1353
rect 6970 1329 6985 1353
rect 6935 1305 6985 1329
rect 7143 1358 7193 1382
rect 7143 1334 7155 1358
rect 7179 1334 7193 1358
rect 7143 1305 7193 1334
rect 7351 1356 7401 1382
rect 19082 1503 19132 1516
rect 19290 1503 19340 1516
rect 19498 1503 19548 1516
rect 19711 1503 19761 1516
rect 17383 1490 17433 1503
rect 17596 1490 17646 1503
rect 17804 1490 17854 1503
rect 18012 1490 18062 1503
rect 14869 1429 14919 1445
rect 15077 1429 15127 1445
rect 15285 1429 15335 1445
rect 15498 1429 15548 1445
rect 7351 1330 7369 1356
rect 7395 1330 7401 1356
rect 7351 1305 7401 1330
rect 9489 1333 9539 1358
rect 9489 1307 9495 1333
rect 9521 1307 9539 1333
rect 9489 1281 9539 1307
rect 9697 1329 9747 1358
rect 9697 1305 9711 1329
rect 9735 1305 9747 1329
rect 9697 1281 9747 1305
rect 9905 1334 9955 1358
rect 9905 1310 9920 1334
rect 9944 1310 9955 1334
rect 9905 1281 9955 1310
rect 10118 1329 10168 1358
rect 10118 1309 10135 1329
rect 10155 1309 10168 1329
rect 12102 1383 12152 1411
rect 12102 1363 12115 1383
rect 12135 1363 12152 1383
rect 12102 1334 12152 1363
rect 12315 1382 12365 1411
rect 12315 1358 12326 1382
rect 12350 1358 12365 1382
rect 12315 1334 12365 1358
rect 12523 1387 12573 1411
rect 12523 1363 12535 1387
rect 12559 1363 12573 1387
rect 12523 1334 12573 1363
rect 12731 1385 12781 1411
rect 12731 1359 12749 1385
rect 12775 1359 12781 1385
rect 12731 1334 12781 1359
rect 14869 1362 14919 1387
rect 14869 1336 14875 1362
rect 14901 1336 14919 1362
rect 10118 1281 10168 1309
rect 14869 1310 14919 1336
rect 15077 1358 15127 1387
rect 15077 1334 15091 1358
rect 15115 1334 15127 1358
rect 15077 1310 15127 1334
rect 15285 1363 15335 1387
rect 15285 1339 15300 1363
rect 15324 1339 15335 1363
rect 15285 1310 15335 1339
rect 15498 1358 15548 1387
rect 15498 1338 15515 1358
rect 15535 1338 15548 1358
rect 20150 1408 20200 1424
rect 20358 1408 20408 1424
rect 20566 1408 20616 1424
rect 20779 1408 20829 1424
rect 15498 1310 15548 1338
rect 5660 1243 5710 1256
rect 5873 1243 5923 1256
rect 6081 1243 6131 1256
rect 6289 1243 6339 1256
rect 6722 1247 6772 1263
rect 6935 1247 6985 1263
rect 7143 1247 7193 1263
rect 7351 1247 7401 1263
rect 4208 1189 4258 1202
rect 4416 1189 4466 1202
rect 4624 1189 4674 1202
rect 4837 1189 4887 1202
rect 379 1136 429 1164
rect 379 1116 392 1136
rect 412 1116 429 1136
rect 379 1087 429 1116
rect 592 1135 642 1164
rect 592 1111 603 1135
rect 627 1111 642 1135
rect 592 1087 642 1111
rect 800 1140 850 1164
rect 800 1116 812 1140
rect 836 1116 850 1140
rect 800 1087 850 1116
rect 1008 1138 1058 1164
rect 1008 1112 1026 1138
rect 1052 1112 1058 1138
rect 1008 1087 1058 1112
rect 3195 1120 3245 1145
rect 1391 1083 1441 1096
rect 1604 1083 1654 1096
rect 1812 1083 1862 1096
rect 2020 1083 2070 1096
rect 3195 1094 3201 1120
rect 3227 1094 3245 1120
rect 379 1029 429 1045
rect 592 1029 642 1045
rect 800 1029 850 1045
rect 1008 1029 1058 1045
rect 3195 1068 3245 1094
rect 3403 1116 3453 1145
rect 3403 1092 3417 1116
rect 3441 1092 3453 1116
rect 3403 1068 3453 1092
rect 3611 1121 3661 1145
rect 3611 1097 3626 1121
rect 3650 1097 3661 1121
rect 3611 1068 3661 1097
rect 3824 1116 3874 1145
rect 3824 1096 3841 1116
rect 3861 1096 3874 1116
rect 3824 1068 3874 1096
rect 8476 1166 8526 1182
rect 8684 1166 8734 1182
rect 8892 1166 8942 1182
rect 9105 1166 9155 1182
rect 11040 1272 11090 1285
rect 11253 1272 11303 1285
rect 11461 1272 11511 1285
rect 11669 1272 11719 1285
rect 12102 1276 12152 1292
rect 12315 1276 12365 1292
rect 12523 1276 12573 1292
rect 12731 1276 12781 1292
rect 9489 1168 9539 1181
rect 9697 1168 9747 1181
rect 9905 1168 9955 1181
rect 10118 1168 10168 1181
rect 5660 1115 5710 1143
rect 5660 1095 5673 1115
rect 5693 1095 5710 1115
rect 1391 955 1441 983
rect 1391 935 1404 955
rect 1424 935 1441 955
rect 1391 906 1441 935
rect 1604 954 1654 983
rect 1604 930 1615 954
rect 1639 930 1654 954
rect 1604 906 1654 930
rect 1812 959 1862 983
rect 1812 935 1824 959
rect 1848 935 1862 959
rect 1812 906 1862 935
rect 2020 957 2070 983
rect 5660 1066 5710 1095
rect 5873 1114 5923 1143
rect 5873 1090 5884 1114
rect 5908 1090 5923 1114
rect 5873 1066 5923 1090
rect 6081 1119 6131 1143
rect 6081 1095 6093 1119
rect 6117 1095 6131 1119
rect 6081 1066 6131 1095
rect 6289 1117 6339 1143
rect 13856 1195 13906 1211
rect 14064 1195 14114 1211
rect 14272 1195 14322 1211
rect 14485 1195 14535 1211
rect 17383 1362 17433 1390
rect 17383 1342 17396 1362
rect 17416 1342 17433 1362
rect 17383 1313 17433 1342
rect 17596 1361 17646 1390
rect 17596 1337 17607 1361
rect 17631 1337 17646 1361
rect 17596 1313 17646 1337
rect 17804 1366 17854 1390
rect 17804 1342 17816 1366
rect 17840 1342 17854 1366
rect 17804 1313 17854 1342
rect 18012 1364 18062 1390
rect 18012 1338 18030 1364
rect 18056 1338 18062 1364
rect 18012 1313 18062 1338
rect 20150 1341 20200 1366
rect 20150 1315 20156 1341
rect 20182 1315 20200 1341
rect 20150 1289 20200 1315
rect 20358 1337 20408 1366
rect 20358 1313 20372 1337
rect 20396 1313 20408 1337
rect 20358 1289 20408 1313
rect 20566 1342 20616 1366
rect 20566 1318 20581 1342
rect 20605 1318 20616 1342
rect 20566 1289 20616 1318
rect 20779 1337 20829 1366
rect 20779 1317 20796 1337
rect 20816 1317 20829 1337
rect 20779 1289 20829 1317
rect 16321 1251 16371 1264
rect 16534 1251 16584 1264
rect 16742 1251 16792 1264
rect 16950 1251 17000 1264
rect 17383 1255 17433 1271
rect 17596 1255 17646 1271
rect 17804 1255 17854 1271
rect 18012 1255 18062 1271
rect 14869 1197 14919 1210
rect 15077 1197 15127 1210
rect 15285 1197 15335 1210
rect 15498 1197 15548 1210
rect 6289 1091 6307 1117
rect 6333 1091 6339 1117
rect 6289 1066 6339 1091
rect 8476 1099 8526 1124
rect 6672 1062 6722 1075
rect 6885 1062 6935 1075
rect 7093 1062 7143 1075
rect 7301 1062 7351 1075
rect 8476 1073 8482 1099
rect 8508 1073 8526 1099
rect 4207 1006 4257 1022
rect 4415 1006 4465 1022
rect 4623 1006 4673 1022
rect 4836 1006 4886 1022
rect 5660 1008 5710 1024
rect 5873 1008 5923 1024
rect 6081 1008 6131 1024
rect 6289 1008 6339 1024
rect 2020 931 2038 957
rect 2064 931 2070 957
rect 3195 955 3245 968
rect 3403 955 3453 968
rect 3611 955 3661 968
rect 3824 955 3874 968
rect 2020 906 2070 931
rect 4207 939 4257 964
rect 4207 913 4213 939
rect 4239 913 4257 939
rect 4207 887 4257 913
rect 4415 935 4465 964
rect 4415 911 4429 935
rect 4453 911 4465 935
rect 4415 887 4465 911
rect 4623 940 4673 964
rect 4623 916 4638 940
rect 4662 916 4673 940
rect 4623 887 4673 916
rect 4836 935 4886 964
rect 8476 1047 8526 1073
rect 8684 1095 8734 1124
rect 8684 1071 8698 1095
rect 8722 1071 8734 1095
rect 8684 1047 8734 1071
rect 8892 1100 8942 1124
rect 8892 1076 8907 1100
rect 8931 1076 8942 1100
rect 8892 1047 8942 1076
rect 9105 1095 9155 1124
rect 11040 1144 11090 1172
rect 11040 1124 11053 1144
rect 11073 1124 11090 1144
rect 9105 1075 9122 1095
rect 9142 1075 9155 1095
rect 9105 1047 9155 1075
rect 11040 1095 11090 1124
rect 11253 1143 11303 1172
rect 11253 1119 11264 1143
rect 11288 1119 11303 1143
rect 11253 1095 11303 1119
rect 11461 1148 11511 1172
rect 11461 1124 11473 1148
rect 11497 1124 11511 1148
rect 11461 1095 11511 1124
rect 11669 1146 11719 1172
rect 11669 1120 11687 1146
rect 11713 1120 11719 1146
rect 11669 1095 11719 1120
rect 13856 1128 13906 1153
rect 12052 1091 12102 1104
rect 12265 1091 12315 1104
rect 12473 1091 12523 1104
rect 12681 1091 12731 1104
rect 13856 1102 13862 1128
rect 13888 1102 13906 1128
rect 4836 915 4853 935
rect 4873 915 4886 935
rect 4836 887 4886 915
rect 378 849 428 862
rect 591 849 641 862
rect 799 849 849 862
rect 1007 849 1057 862
rect 1391 848 1441 864
rect 1604 848 1654 864
rect 1812 848 1862 864
rect 2020 848 2070 864
rect 6672 934 6722 962
rect 6672 914 6685 934
rect 6705 914 6722 934
rect 6672 885 6722 914
rect 6885 933 6935 962
rect 6885 909 6896 933
rect 6920 909 6935 933
rect 6885 885 6935 909
rect 7093 938 7143 962
rect 7093 914 7105 938
rect 7129 914 7143 938
rect 7093 885 7143 914
rect 7301 936 7351 962
rect 11040 1037 11090 1053
rect 11253 1037 11303 1053
rect 11461 1037 11511 1053
rect 11669 1037 11719 1053
rect 9488 985 9538 1001
rect 9696 985 9746 1001
rect 9904 985 9954 1001
rect 10117 985 10167 1001
rect 13856 1076 13906 1102
rect 14064 1124 14114 1153
rect 14064 1100 14078 1124
rect 14102 1100 14114 1124
rect 14064 1076 14114 1100
rect 14272 1129 14322 1153
rect 14272 1105 14287 1129
rect 14311 1105 14322 1129
rect 14272 1076 14322 1105
rect 14485 1124 14535 1153
rect 14485 1104 14502 1124
rect 14522 1104 14535 1124
rect 14485 1076 14535 1104
rect 19137 1174 19187 1190
rect 19345 1174 19395 1190
rect 19553 1174 19603 1190
rect 19766 1174 19816 1190
rect 20150 1176 20200 1189
rect 20358 1176 20408 1189
rect 20566 1176 20616 1189
rect 20779 1176 20829 1189
rect 16321 1123 16371 1151
rect 16321 1103 16334 1123
rect 16354 1103 16371 1123
rect 7301 910 7319 936
rect 7345 910 7351 936
rect 8476 934 8526 947
rect 8684 934 8734 947
rect 8892 934 8942 947
rect 9105 934 9155 947
rect 7301 885 7351 910
rect 9488 918 9538 943
rect 9488 892 9494 918
rect 9520 892 9538 918
rect 9488 866 9538 892
rect 9696 914 9746 943
rect 9696 890 9710 914
rect 9734 890 9746 914
rect 9696 866 9746 890
rect 9904 919 9954 943
rect 9904 895 9919 919
rect 9943 895 9954 919
rect 9904 866 9954 895
rect 10117 914 10167 943
rect 12052 963 12102 991
rect 12052 943 12065 963
rect 12085 943 12102 963
rect 10117 894 10134 914
rect 10154 894 10167 914
rect 10117 866 10167 894
rect 12052 914 12102 943
rect 12265 962 12315 991
rect 12265 938 12276 962
rect 12300 938 12315 962
rect 12265 914 12315 938
rect 12473 967 12523 991
rect 12473 943 12485 967
rect 12509 943 12523 967
rect 12473 914 12523 943
rect 12681 965 12731 991
rect 16321 1074 16371 1103
rect 16534 1122 16584 1151
rect 16534 1098 16545 1122
rect 16569 1098 16584 1122
rect 16534 1074 16584 1098
rect 16742 1127 16792 1151
rect 16742 1103 16754 1127
rect 16778 1103 16792 1127
rect 16742 1074 16792 1103
rect 16950 1125 17000 1151
rect 16950 1099 16968 1125
rect 16994 1099 17000 1125
rect 16950 1074 17000 1099
rect 19137 1107 19187 1132
rect 17333 1070 17383 1083
rect 17546 1070 17596 1083
rect 17754 1070 17804 1083
rect 17962 1070 18012 1083
rect 19137 1081 19143 1107
rect 19169 1081 19187 1107
rect 14868 1014 14918 1030
rect 15076 1014 15126 1030
rect 15284 1014 15334 1030
rect 15497 1014 15547 1030
rect 16321 1016 16371 1032
rect 16534 1016 16584 1032
rect 16742 1016 16792 1032
rect 16950 1016 17000 1032
rect 12681 939 12699 965
rect 12725 939 12731 965
rect 13856 963 13906 976
rect 14064 963 14114 976
rect 14272 963 14322 976
rect 14485 963 14535 976
rect 12681 914 12731 939
rect 14868 947 14918 972
rect 14868 921 14874 947
rect 14900 921 14918 947
rect 5659 828 5709 841
rect 5872 828 5922 841
rect 6080 828 6130 841
rect 6288 828 6338 841
rect 4207 774 4257 787
rect 4415 774 4465 787
rect 4623 774 4673 787
rect 4836 774 4886 787
rect 378 721 428 749
rect 378 701 391 721
rect 411 701 428 721
rect 378 672 428 701
rect 591 720 641 749
rect 591 696 602 720
rect 626 696 641 720
rect 591 672 641 696
rect 799 725 849 749
rect 799 701 811 725
rect 835 701 849 725
rect 799 672 849 701
rect 1007 723 1057 749
rect 1007 697 1025 723
rect 1051 697 1057 723
rect 1007 672 1057 697
rect 6672 827 6722 843
rect 6885 827 6935 843
rect 7093 827 7143 843
rect 7301 827 7351 843
rect 14868 895 14918 921
rect 15076 943 15126 972
rect 15076 919 15090 943
rect 15114 919 15126 943
rect 15076 895 15126 919
rect 15284 948 15334 972
rect 15284 924 15299 948
rect 15323 924 15334 948
rect 15284 895 15334 924
rect 15497 943 15547 972
rect 19137 1055 19187 1081
rect 19345 1103 19395 1132
rect 19345 1079 19359 1103
rect 19383 1079 19395 1103
rect 19345 1055 19395 1079
rect 19553 1108 19603 1132
rect 19553 1084 19568 1108
rect 19592 1084 19603 1108
rect 19553 1055 19603 1084
rect 19766 1103 19816 1132
rect 19766 1083 19783 1103
rect 19803 1083 19816 1103
rect 19766 1055 19816 1083
rect 15497 923 15514 943
rect 15534 923 15547 943
rect 15497 895 15547 923
rect 11039 857 11089 870
rect 11252 857 11302 870
rect 11460 857 11510 870
rect 11668 857 11718 870
rect 9488 753 9538 766
rect 9696 753 9746 766
rect 9904 753 9954 766
rect 10117 753 10167 766
rect 12052 856 12102 872
rect 12265 856 12315 872
rect 12473 856 12523 872
rect 12681 856 12731 872
rect 17333 942 17383 970
rect 17333 922 17346 942
rect 17366 922 17383 942
rect 17333 893 17383 922
rect 17546 941 17596 970
rect 17546 917 17557 941
rect 17581 917 17596 941
rect 17546 893 17596 917
rect 17754 946 17804 970
rect 17754 922 17766 946
rect 17790 922 17804 946
rect 17754 893 17804 922
rect 17962 944 18012 970
rect 20149 993 20199 1009
rect 20357 993 20407 1009
rect 20565 993 20615 1009
rect 20778 993 20828 1009
rect 17962 918 17980 944
rect 18006 918 18012 944
rect 19137 942 19187 955
rect 19345 942 19395 955
rect 19553 942 19603 955
rect 19766 942 19816 955
rect 17962 893 18012 918
rect 20149 926 20199 951
rect 20149 900 20155 926
rect 20181 900 20199 926
rect 20149 874 20199 900
rect 20357 922 20407 951
rect 20357 898 20371 922
rect 20395 898 20407 922
rect 20357 874 20407 898
rect 20565 927 20615 951
rect 20565 903 20580 927
rect 20604 903 20615 927
rect 20565 874 20615 903
rect 20778 922 20828 951
rect 20778 902 20795 922
rect 20815 902 20828 922
rect 20778 874 20828 902
rect 16320 836 16370 849
rect 16533 836 16583 849
rect 16741 836 16791 849
rect 16949 836 16999 849
rect 14868 782 14918 795
rect 15076 782 15126 795
rect 15284 782 15334 795
rect 15497 782 15547 795
rect 11039 729 11089 757
rect 5659 700 5709 728
rect 5659 680 5672 700
rect 5692 680 5709 700
rect 378 614 428 630
rect 591 614 641 630
rect 799 614 849 630
rect 1007 614 1057 630
rect 5659 651 5709 680
rect 5872 699 5922 728
rect 5872 675 5883 699
rect 5907 675 5922 699
rect 5872 651 5922 675
rect 6080 704 6130 728
rect 6080 680 6092 704
rect 6116 680 6130 704
rect 6080 651 6130 680
rect 6288 702 6338 728
rect 6288 676 6306 702
rect 6332 676 6338 702
rect 6288 651 6338 676
rect 11039 709 11052 729
rect 11072 709 11089 729
rect 11039 680 11089 709
rect 11252 728 11302 757
rect 11252 704 11263 728
rect 11287 704 11302 728
rect 11252 680 11302 704
rect 11460 733 11510 757
rect 11460 709 11472 733
rect 11496 709 11510 733
rect 11460 680 11510 709
rect 11668 731 11718 757
rect 11668 705 11686 731
rect 11712 705 11718 731
rect 11668 680 11718 705
rect 17333 835 17383 851
rect 17546 835 17596 851
rect 17754 835 17804 851
rect 17962 835 18012 851
rect 20149 761 20199 774
rect 20357 761 20407 774
rect 20565 761 20615 774
rect 20778 761 20828 774
rect 16320 708 16370 736
rect 16320 688 16333 708
rect 16353 688 16370 708
rect 11039 622 11089 638
rect 11252 622 11302 638
rect 11460 622 11510 638
rect 11668 622 11718 638
rect 5659 593 5709 609
rect 5872 593 5922 609
rect 6080 593 6130 609
rect 6288 593 6338 609
rect 16320 659 16370 688
rect 16533 707 16583 736
rect 16533 683 16544 707
rect 16568 683 16583 707
rect 16533 659 16583 683
rect 16741 712 16791 736
rect 16741 688 16753 712
rect 16777 688 16791 712
rect 16741 659 16791 688
rect 16949 710 16999 736
rect 16949 684 16967 710
rect 16993 684 16999 710
rect 16949 659 16999 684
rect 16320 601 16370 617
rect 16533 601 16583 617
rect 16741 601 16791 617
rect 16949 601 16999 617
rect 1781 368 1831 381
rect 1994 368 2044 381
rect 2202 368 2252 381
rect 2410 368 2460 381
rect 12442 376 12492 389
rect 12655 376 12705 389
rect 12863 376 12913 389
rect 13071 376 13121 389
rect 7062 347 7112 360
rect 7275 347 7325 360
rect 7483 347 7533 360
rect 7691 347 7741 360
rect 4871 280 4921 293
rect 5084 280 5134 293
rect 5292 280 5342 293
rect 5500 280 5550 293
rect 1781 240 1831 268
rect 1781 220 1794 240
rect 1814 220 1831 240
rect 1781 191 1831 220
rect 1994 239 2044 268
rect 1994 215 2005 239
rect 2029 215 2044 239
rect 1994 191 2044 215
rect 2202 244 2252 268
rect 2202 220 2214 244
rect 2238 220 2252 244
rect 2202 191 2252 220
rect 2410 242 2460 268
rect 2410 216 2428 242
rect 2454 216 2460 242
rect 2410 191 2460 216
rect 10132 273 10182 286
rect 10345 273 10395 286
rect 10553 273 10603 286
rect 10761 273 10811 286
rect 17723 355 17773 368
rect 17936 355 17986 368
rect 18144 355 18194 368
rect 18352 355 18402 368
rect 15532 288 15582 301
rect 15745 288 15795 301
rect 15953 288 16003 301
rect 16161 288 16211 301
rect 7062 219 7112 247
rect 7062 199 7075 219
rect 7095 199 7112 219
rect 4871 152 4921 180
rect 1781 133 1831 149
rect 1994 133 2044 149
rect 2202 133 2252 149
rect 2410 133 2460 149
rect 4871 132 4884 152
rect 4904 132 4921 152
rect 4871 103 4921 132
rect 5084 151 5134 180
rect 5084 127 5095 151
rect 5119 127 5134 151
rect 5084 103 5134 127
rect 5292 156 5342 180
rect 5292 132 5304 156
rect 5328 132 5342 156
rect 5292 103 5342 132
rect 5500 154 5550 180
rect 7062 170 7112 199
rect 7275 218 7325 247
rect 7275 194 7286 218
rect 7310 194 7325 218
rect 7275 170 7325 194
rect 7483 223 7533 247
rect 7483 199 7495 223
rect 7519 199 7533 223
rect 7483 170 7533 199
rect 7691 221 7741 247
rect 7691 195 7709 221
rect 7735 195 7741 221
rect 7691 170 7741 195
rect 12442 248 12492 276
rect 12442 228 12455 248
rect 12475 228 12492 248
rect 12442 199 12492 228
rect 12655 247 12705 276
rect 12655 223 12666 247
rect 12690 223 12705 247
rect 12655 199 12705 223
rect 12863 252 12913 276
rect 12863 228 12875 252
rect 12899 228 12913 252
rect 12863 199 12913 228
rect 13071 250 13121 276
rect 13071 224 13089 250
rect 13115 224 13121 250
rect 13071 199 13121 224
rect 5500 128 5518 154
rect 5544 128 5550 154
rect 10132 145 10182 173
rect 5500 103 5550 128
rect 7062 112 7112 128
rect 7275 112 7325 128
rect 7483 112 7533 128
rect 7691 112 7741 128
rect 10132 125 10145 145
rect 10165 125 10182 145
rect 10132 96 10182 125
rect 10345 144 10395 173
rect 10345 120 10356 144
rect 10380 120 10395 144
rect 10345 96 10395 120
rect 10553 149 10603 173
rect 10553 125 10565 149
rect 10589 125 10603 149
rect 10553 96 10603 125
rect 10761 147 10811 173
rect 17723 227 17773 255
rect 17723 207 17736 227
rect 17756 207 17773 227
rect 15532 160 15582 188
rect 10761 121 10779 147
rect 10805 121 10811 147
rect 12442 141 12492 157
rect 12655 141 12705 157
rect 12863 141 12913 157
rect 13071 141 13121 157
rect 10761 96 10811 121
rect 15532 140 15545 160
rect 15565 140 15582 160
rect 15532 111 15582 140
rect 15745 159 15795 188
rect 15745 135 15756 159
rect 15780 135 15795 159
rect 15745 111 15795 135
rect 15953 164 16003 188
rect 15953 140 15965 164
rect 15989 140 16003 164
rect 15953 111 16003 140
rect 16161 162 16211 188
rect 17723 178 17773 207
rect 17936 226 17986 255
rect 17936 202 17947 226
rect 17971 202 17986 226
rect 17936 178 17986 202
rect 18144 231 18194 255
rect 18144 207 18156 231
rect 18180 207 18194 231
rect 18144 178 18194 207
rect 18352 229 18402 255
rect 18352 203 18370 229
rect 18396 203 18402 229
rect 18352 178 18402 203
rect 16161 136 16179 162
rect 16205 136 16211 162
rect 16161 111 16211 136
rect 17723 120 17773 136
rect 17936 120 17986 136
rect 18144 120 18194 136
rect 18352 120 18402 136
rect 4871 45 4921 61
rect 5084 45 5134 61
rect 5292 45 5342 61
rect 5500 45 5550 61
rect 10132 38 10182 54
rect 10345 38 10395 54
rect 10553 38 10603 54
rect 10761 38 10811 54
rect 15532 53 15582 69
rect 15745 53 15795 69
rect 15953 53 16003 69
rect 16161 53 16211 69
<< polycont >>
rect 4177 8186 4203 8212
rect 4393 8184 4417 8208
rect 4602 8189 4626 8213
rect 4817 8188 4837 8208
rect 9458 8165 9484 8191
rect 9674 8163 9698 8187
rect 9883 8168 9907 8192
rect 10098 8167 10118 8187
rect 14838 8194 14864 8220
rect 15054 8192 15078 8216
rect 15263 8197 15287 8221
rect 15478 8196 15498 8216
rect 355 7974 375 7994
rect 566 7969 590 7993
rect 775 7974 799 7998
rect 989 7970 1015 7996
rect 3164 7952 3190 7978
rect 3380 7950 3404 7974
rect 3589 7955 3613 7979
rect 3804 7954 3824 7974
rect 5636 7953 5656 7973
rect 1367 7793 1387 7813
rect 1578 7788 1602 7812
rect 1787 7793 1811 7817
rect 5847 7948 5871 7972
rect 6056 7953 6080 7977
rect 20119 8173 20145 8199
rect 20335 8171 20359 8195
rect 20544 8176 20568 8200
rect 20759 8175 20779 8195
rect 6270 7949 6296 7975
rect 8445 7931 8471 7957
rect 2001 7789 2027 7815
rect 4176 7771 4202 7797
rect 4392 7769 4416 7793
rect 4601 7774 4625 7798
rect 8661 7929 8685 7953
rect 8870 7934 8894 7958
rect 11016 7982 11036 8002
rect 9085 7933 9105 7953
rect 11227 7977 11251 8001
rect 11436 7982 11460 8006
rect 11650 7978 11676 8004
rect 13825 7960 13851 7986
rect 4816 7773 4836 7793
rect 6648 7772 6668 7792
rect 6859 7767 6883 7791
rect 7068 7772 7092 7796
rect 14041 7958 14065 7982
rect 14250 7963 14274 7987
rect 14465 7962 14485 7982
rect 16297 7961 16317 7981
rect 7282 7768 7308 7794
rect 9457 7750 9483 7776
rect 9673 7748 9697 7772
rect 9882 7753 9906 7777
rect 12028 7801 12048 7821
rect 10097 7752 10117 7772
rect 12239 7796 12263 7820
rect 12448 7801 12472 7825
rect 16508 7956 16532 7980
rect 16717 7961 16741 7985
rect 16931 7957 16957 7983
rect 19106 7939 19132 7965
rect 12662 7797 12688 7823
rect 14837 7779 14863 7805
rect 354 7559 374 7579
rect 565 7554 589 7578
rect 774 7559 798 7583
rect 988 7555 1014 7581
rect 3114 7532 3140 7558
rect 3330 7530 3354 7554
rect 3539 7535 3563 7559
rect 3754 7534 3774 7554
rect 15053 7777 15077 7801
rect 15262 7782 15286 7806
rect 19322 7937 19346 7961
rect 19531 7942 19555 7966
rect 19746 7941 19766 7961
rect 15477 7781 15497 7801
rect 17309 7780 17329 7800
rect 17520 7775 17544 7799
rect 17729 7780 17753 7804
rect 17943 7776 17969 7802
rect 20118 7758 20144 7784
rect 20334 7756 20358 7780
rect 20543 7761 20567 7785
rect 20758 7760 20778 7780
rect 5635 7538 5655 7558
rect 5846 7533 5870 7557
rect 6055 7538 6079 7562
rect 6269 7534 6295 7560
rect 8395 7511 8421 7537
rect 8611 7509 8635 7533
rect 8820 7514 8844 7538
rect 9035 7513 9055 7533
rect 11015 7567 11035 7587
rect 11226 7562 11250 7586
rect 11435 7567 11459 7591
rect 11649 7563 11675 7589
rect 13775 7540 13801 7566
rect 13991 7538 14015 7562
rect 14200 7543 14224 7567
rect 14415 7542 14435 7562
rect 16296 7546 16316 7566
rect 16507 7541 16531 7565
rect 16716 7546 16740 7570
rect 16930 7542 16956 7568
rect 19056 7519 19082 7545
rect 19272 7517 19296 7541
rect 19481 7522 19505 7546
rect 19696 7521 19716 7541
rect 1422 7232 1442 7252
rect 1633 7227 1657 7251
rect 1842 7232 1866 7256
rect 2056 7228 2082 7254
rect 4182 7205 4208 7231
rect 4398 7203 4422 7227
rect 4607 7208 4631 7232
rect 4822 7207 4842 7227
rect 6703 7211 6723 7231
rect 6914 7206 6938 7230
rect 7123 7211 7147 7235
rect 7337 7207 7363 7233
rect 9463 7184 9489 7210
rect 9679 7182 9703 7206
rect 9888 7187 9912 7211
rect 10103 7186 10123 7206
rect 12083 7240 12103 7260
rect 12294 7235 12318 7259
rect 12503 7240 12527 7264
rect 12717 7236 12743 7262
rect 14843 7213 14869 7239
rect 15059 7211 15083 7235
rect 15268 7216 15292 7240
rect 15483 7215 15503 7235
rect 360 6993 380 7013
rect 571 6988 595 7012
rect 780 6993 804 7017
rect 994 6989 1020 7015
rect 3169 6971 3195 6997
rect 3385 6969 3409 6993
rect 3594 6974 3618 6998
rect 3809 6973 3829 6993
rect 5641 6972 5661 6992
rect 1372 6812 1392 6832
rect 1583 6807 1607 6831
rect 1792 6812 1816 6836
rect 5852 6967 5876 6991
rect 6061 6972 6085 6996
rect 17364 7219 17384 7239
rect 17575 7214 17599 7238
rect 17784 7219 17808 7243
rect 17998 7215 18024 7241
rect 20124 7192 20150 7218
rect 20340 7190 20364 7214
rect 20549 7195 20573 7219
rect 20764 7194 20784 7214
rect 6275 6968 6301 6994
rect 8450 6950 8476 6976
rect 2006 6808 2032 6834
rect 4181 6790 4207 6816
rect 4397 6788 4421 6812
rect 4606 6793 4630 6817
rect 8666 6948 8690 6972
rect 8875 6953 8899 6977
rect 11021 7001 11041 7021
rect 9090 6952 9110 6972
rect 11232 6996 11256 7020
rect 11441 7001 11465 7025
rect 11655 6997 11681 7023
rect 13830 6979 13856 7005
rect 4821 6792 4841 6812
rect 6653 6791 6673 6811
rect 6864 6786 6888 6810
rect 7073 6791 7097 6815
rect 14046 6977 14070 7001
rect 14255 6982 14279 7006
rect 14470 6981 14490 7001
rect 16302 6980 16322 7000
rect 7287 6787 7313 6813
rect 9462 6769 9488 6795
rect 9678 6767 9702 6791
rect 9887 6772 9911 6796
rect 12033 6820 12053 6840
rect 10102 6771 10122 6791
rect 12244 6815 12268 6839
rect 12453 6820 12477 6844
rect 16513 6975 16537 6999
rect 16722 6980 16746 7004
rect 16936 6976 16962 7002
rect 19111 6958 19137 6984
rect 12667 6816 12693 6842
rect 14842 6798 14868 6824
rect 359 6578 379 6598
rect 570 6573 594 6597
rect 779 6578 803 6602
rect 993 6574 1019 6600
rect 15058 6796 15082 6820
rect 15267 6801 15291 6825
rect 19327 6956 19351 6980
rect 19536 6961 19560 6985
rect 19751 6960 19771 6980
rect 15482 6800 15502 6820
rect 17314 6799 17334 6819
rect 17525 6794 17549 6818
rect 17734 6799 17758 6823
rect 17948 6795 17974 6821
rect 20123 6777 20149 6803
rect 20339 6775 20363 6799
rect 20548 6780 20572 6804
rect 20763 6779 20783 6799
rect 2961 6504 2987 6530
rect 3177 6502 3201 6526
rect 3386 6507 3410 6531
rect 3601 6506 3621 6526
rect 5640 6557 5660 6577
rect 5851 6552 5875 6576
rect 6060 6557 6084 6581
rect 6274 6553 6300 6579
rect 11020 6586 11040 6606
rect 8242 6483 8268 6509
rect 8458 6481 8482 6505
rect 8667 6486 8691 6510
rect 11231 6581 11255 6605
rect 11440 6586 11464 6610
rect 11654 6582 11680 6608
rect 8882 6485 8902 6505
rect 13622 6512 13648 6538
rect 13838 6510 13862 6534
rect 14047 6515 14071 6539
rect 14262 6514 14282 6534
rect 16301 6565 16321 6585
rect 16512 6560 16536 6584
rect 16721 6565 16745 6589
rect 16935 6561 16961 6587
rect 1587 6300 1607 6320
rect 1798 6295 1822 6319
rect 2007 6300 2031 6324
rect 2221 6296 2247 6322
rect 18903 6491 18929 6517
rect 19119 6489 19143 6513
rect 19328 6494 19352 6518
rect 19543 6493 19563 6513
rect 4189 6226 4215 6252
rect 4405 6224 4429 6248
rect 4614 6229 4638 6253
rect 4829 6228 4849 6248
rect 6868 6279 6888 6299
rect 7079 6274 7103 6298
rect 7288 6279 7312 6303
rect 7502 6275 7528 6301
rect 12248 6308 12268 6328
rect 9470 6205 9496 6231
rect 9686 6203 9710 6227
rect 9895 6208 9919 6232
rect 12459 6303 12483 6327
rect 12668 6308 12692 6332
rect 12882 6304 12908 6330
rect 10110 6207 10130 6227
rect 14850 6234 14876 6260
rect 15066 6232 15090 6256
rect 15275 6237 15299 6261
rect 15490 6236 15510 6256
rect 17529 6287 17549 6307
rect 17740 6282 17764 6306
rect 17949 6287 17973 6311
rect 18163 6283 18189 6309
rect 367 6014 387 6034
rect 578 6009 602 6033
rect 787 6014 811 6038
rect 1001 6010 1027 6036
rect 3176 5992 3202 6018
rect 3392 5990 3416 6014
rect 3601 5995 3625 6019
rect 3816 5994 3836 6014
rect 5648 5993 5668 6013
rect 1379 5833 1399 5853
rect 1590 5828 1614 5852
rect 1799 5833 1823 5857
rect 5859 5988 5883 6012
rect 6068 5993 6092 6017
rect 20131 6213 20157 6239
rect 20347 6211 20371 6235
rect 20556 6216 20580 6240
rect 20771 6215 20791 6235
rect 6282 5989 6308 6015
rect 8457 5971 8483 5997
rect 2013 5829 2039 5855
rect 4188 5811 4214 5837
rect 4404 5809 4428 5833
rect 4613 5814 4637 5838
rect 8673 5969 8697 5993
rect 8882 5974 8906 5998
rect 11028 6022 11048 6042
rect 9097 5973 9117 5993
rect 11239 6017 11263 6041
rect 11448 6022 11472 6046
rect 11662 6018 11688 6044
rect 13837 6000 13863 6026
rect 4828 5813 4848 5833
rect 6660 5812 6680 5832
rect 6871 5807 6895 5831
rect 7080 5812 7104 5836
rect 14053 5998 14077 6022
rect 14262 6003 14286 6027
rect 14477 6002 14497 6022
rect 16309 6001 16329 6021
rect 7294 5808 7320 5834
rect 9469 5790 9495 5816
rect 9685 5788 9709 5812
rect 9894 5793 9918 5817
rect 12040 5841 12060 5861
rect 10109 5792 10129 5812
rect 12251 5836 12275 5860
rect 12460 5841 12484 5865
rect 16520 5996 16544 6020
rect 16729 6001 16753 6025
rect 16943 5997 16969 6023
rect 19118 5979 19144 6005
rect 12674 5837 12700 5863
rect 14849 5819 14875 5845
rect 366 5599 386 5619
rect 577 5594 601 5618
rect 786 5599 810 5623
rect 1000 5595 1026 5621
rect 3126 5572 3152 5598
rect 3342 5570 3366 5594
rect 3551 5575 3575 5599
rect 3766 5574 3786 5594
rect 15065 5817 15089 5841
rect 15274 5822 15298 5846
rect 19334 5977 19358 6001
rect 19543 5982 19567 6006
rect 19758 5981 19778 6001
rect 15489 5821 15509 5841
rect 17321 5820 17341 5840
rect 17532 5815 17556 5839
rect 17741 5820 17765 5844
rect 17955 5816 17981 5842
rect 20130 5798 20156 5824
rect 20346 5796 20370 5820
rect 20555 5801 20579 5825
rect 20770 5800 20790 5820
rect 5647 5578 5667 5598
rect 5858 5573 5882 5597
rect 6067 5578 6091 5602
rect 6281 5574 6307 5600
rect 8407 5551 8433 5577
rect 8623 5549 8647 5573
rect 8832 5554 8856 5578
rect 9047 5553 9067 5573
rect 11027 5607 11047 5627
rect 11238 5602 11262 5626
rect 11447 5607 11471 5631
rect 11661 5603 11687 5629
rect 13787 5580 13813 5606
rect 14003 5578 14027 5602
rect 14212 5583 14236 5607
rect 14427 5582 14447 5602
rect 16308 5586 16328 5606
rect 16519 5581 16543 5605
rect 16728 5586 16752 5610
rect 16942 5582 16968 5608
rect 19068 5559 19094 5585
rect 19284 5557 19308 5581
rect 19493 5562 19517 5586
rect 19708 5561 19728 5581
rect 1434 5272 1454 5292
rect 1645 5267 1669 5291
rect 1854 5272 1878 5296
rect 2068 5268 2094 5294
rect 4194 5245 4220 5271
rect 4410 5243 4434 5267
rect 4619 5248 4643 5272
rect 4834 5247 4854 5267
rect 6715 5251 6735 5271
rect 6926 5246 6950 5270
rect 7135 5251 7159 5275
rect 7349 5247 7375 5273
rect 9475 5224 9501 5250
rect 9691 5222 9715 5246
rect 9900 5227 9924 5251
rect 10115 5226 10135 5246
rect 12095 5280 12115 5300
rect 12306 5275 12330 5299
rect 12515 5280 12539 5304
rect 12729 5276 12755 5302
rect 14855 5253 14881 5279
rect 15071 5251 15095 5275
rect 15280 5256 15304 5280
rect 15495 5255 15515 5275
rect 372 5033 392 5053
rect 583 5028 607 5052
rect 792 5033 816 5057
rect 1006 5029 1032 5055
rect 3181 5011 3207 5037
rect 3397 5009 3421 5033
rect 3606 5014 3630 5038
rect 3821 5013 3841 5033
rect 5653 5012 5673 5032
rect 1384 4852 1404 4872
rect 1595 4847 1619 4871
rect 1804 4852 1828 4876
rect 5864 5007 5888 5031
rect 6073 5012 6097 5036
rect 17376 5259 17396 5279
rect 17587 5254 17611 5278
rect 17796 5259 17820 5283
rect 18010 5255 18036 5281
rect 20136 5232 20162 5258
rect 20352 5230 20376 5254
rect 20561 5235 20585 5259
rect 20776 5234 20796 5254
rect 6287 5008 6313 5034
rect 8462 4990 8488 5016
rect 2018 4848 2044 4874
rect 4193 4830 4219 4856
rect 4409 4828 4433 4852
rect 4618 4833 4642 4857
rect 8678 4988 8702 5012
rect 8887 4993 8911 5017
rect 11033 5041 11053 5061
rect 9102 4992 9122 5012
rect 11244 5036 11268 5060
rect 11453 5041 11477 5065
rect 11667 5037 11693 5063
rect 13842 5019 13868 5045
rect 4833 4832 4853 4852
rect 6665 4831 6685 4851
rect 6876 4826 6900 4850
rect 7085 4831 7109 4855
rect 14058 5017 14082 5041
rect 14267 5022 14291 5046
rect 14482 5021 14502 5041
rect 16314 5020 16334 5040
rect 7299 4827 7325 4853
rect 9474 4809 9500 4835
rect 9690 4807 9714 4831
rect 9899 4812 9923 4836
rect 12045 4860 12065 4880
rect 10114 4811 10134 4831
rect 12256 4855 12280 4879
rect 12465 4860 12489 4884
rect 16525 5015 16549 5039
rect 16734 5020 16758 5044
rect 16948 5016 16974 5042
rect 19123 4998 19149 5024
rect 12679 4856 12705 4882
rect 14854 4838 14880 4864
rect 371 4618 391 4638
rect 582 4613 606 4637
rect 791 4618 815 4642
rect 1005 4614 1031 4640
rect 15070 4836 15094 4860
rect 15279 4841 15303 4865
rect 19339 4996 19363 5020
rect 19548 5001 19572 5025
rect 19763 5000 19783 5020
rect 15494 4840 15514 4860
rect 17326 4839 17346 4859
rect 17537 4834 17561 4858
rect 17746 4839 17770 4863
rect 17960 4835 17986 4861
rect 20135 4817 20161 4843
rect 20351 4815 20375 4839
rect 20560 4820 20584 4844
rect 20775 4819 20795 4839
rect 2886 4579 2912 4605
rect 3102 4577 3126 4601
rect 3311 4582 3335 4606
rect 3526 4581 3546 4601
rect 5652 4597 5672 4617
rect 5863 4592 5887 4616
rect 6072 4597 6096 4621
rect 6286 4593 6312 4619
rect 11032 4626 11052 4646
rect 8167 4558 8193 4584
rect 8383 4556 8407 4580
rect 8592 4561 8616 4585
rect 8807 4560 8827 4580
rect 11243 4621 11267 4645
rect 11452 4626 11476 4650
rect 11666 4622 11692 4648
rect 1682 4308 1702 4328
rect 1893 4303 1917 4327
rect 2102 4308 2126 4332
rect 2316 4304 2342 4330
rect 4197 4269 4223 4295
rect 4413 4267 4437 4291
rect 4622 4272 4646 4296
rect 4837 4271 4857 4291
rect 13547 4587 13573 4613
rect 13763 4585 13787 4609
rect 13972 4590 13996 4614
rect 14187 4589 14207 4609
rect 6963 4287 6983 4307
rect 7174 4282 7198 4306
rect 7383 4287 7407 4311
rect 7597 4283 7623 4309
rect 16313 4605 16333 4625
rect 16524 4600 16548 4624
rect 16733 4605 16757 4629
rect 16947 4601 16973 4627
rect 18828 4566 18854 4592
rect 19044 4564 19068 4588
rect 19253 4569 19277 4593
rect 19468 4568 19488 4588
rect 9478 4248 9504 4274
rect 9694 4246 9718 4270
rect 9903 4251 9927 4275
rect 12343 4316 12363 4336
rect 12554 4311 12578 4335
rect 12763 4316 12787 4340
rect 12977 4312 13003 4338
rect 10118 4250 10138 4270
rect 14858 4277 14884 4303
rect 15074 4275 15098 4299
rect 15283 4280 15307 4304
rect 15498 4279 15518 4299
rect 17624 4295 17644 4315
rect 17835 4290 17859 4314
rect 18044 4295 18068 4319
rect 18258 4291 18284 4317
rect 375 4057 395 4077
rect 586 4052 610 4076
rect 795 4057 819 4081
rect 1009 4053 1035 4079
rect 3184 4035 3210 4061
rect 3400 4033 3424 4057
rect 3609 4038 3633 4062
rect 3824 4037 3844 4057
rect 5656 4036 5676 4056
rect 1387 3876 1407 3896
rect 1598 3871 1622 3895
rect 1807 3876 1831 3900
rect 5867 4031 5891 4055
rect 6076 4036 6100 4060
rect 20139 4256 20165 4282
rect 20355 4254 20379 4278
rect 20564 4259 20588 4283
rect 20779 4258 20799 4278
rect 6290 4032 6316 4058
rect 8465 4014 8491 4040
rect 2021 3872 2047 3898
rect 4196 3854 4222 3880
rect 4412 3852 4436 3876
rect 4621 3857 4645 3881
rect 8681 4012 8705 4036
rect 8890 4017 8914 4041
rect 11036 4065 11056 4085
rect 9105 4016 9125 4036
rect 11247 4060 11271 4084
rect 11456 4065 11480 4089
rect 11670 4061 11696 4087
rect 13845 4043 13871 4069
rect 4836 3856 4856 3876
rect 6668 3855 6688 3875
rect 6879 3850 6903 3874
rect 7088 3855 7112 3879
rect 14061 4041 14085 4065
rect 14270 4046 14294 4070
rect 14485 4045 14505 4065
rect 16317 4044 16337 4064
rect 7302 3851 7328 3877
rect 9477 3833 9503 3859
rect 9693 3831 9717 3855
rect 9902 3836 9926 3860
rect 12048 3884 12068 3904
rect 10117 3835 10137 3855
rect 12259 3879 12283 3903
rect 12468 3884 12492 3908
rect 16528 4039 16552 4063
rect 16737 4044 16761 4068
rect 16951 4040 16977 4066
rect 19126 4022 19152 4048
rect 12682 3880 12708 3906
rect 14857 3862 14883 3888
rect 374 3642 394 3662
rect 585 3637 609 3661
rect 794 3642 818 3666
rect 1008 3638 1034 3664
rect 3134 3615 3160 3641
rect 3350 3613 3374 3637
rect 3559 3618 3583 3642
rect 3774 3617 3794 3637
rect 15073 3860 15097 3884
rect 15282 3865 15306 3889
rect 19342 4020 19366 4044
rect 19551 4025 19575 4049
rect 19766 4024 19786 4044
rect 15497 3864 15517 3884
rect 17329 3863 17349 3883
rect 17540 3858 17564 3882
rect 17749 3863 17773 3887
rect 17963 3859 17989 3885
rect 20138 3841 20164 3867
rect 20354 3839 20378 3863
rect 20563 3844 20587 3868
rect 20778 3843 20798 3863
rect 5655 3621 5675 3641
rect 5866 3616 5890 3640
rect 6075 3621 6099 3645
rect 6289 3617 6315 3643
rect 8415 3594 8441 3620
rect 8631 3592 8655 3616
rect 8840 3597 8864 3621
rect 9055 3596 9075 3616
rect 11035 3650 11055 3670
rect 11246 3645 11270 3669
rect 11455 3650 11479 3674
rect 11669 3646 11695 3672
rect 13795 3623 13821 3649
rect 14011 3621 14035 3645
rect 14220 3626 14244 3650
rect 14435 3625 14455 3645
rect 16316 3629 16336 3649
rect 16527 3624 16551 3648
rect 16736 3629 16760 3653
rect 16950 3625 16976 3651
rect 19076 3602 19102 3628
rect 19292 3600 19316 3624
rect 19501 3605 19525 3629
rect 19716 3604 19736 3624
rect 1442 3315 1462 3335
rect 1653 3310 1677 3334
rect 1862 3315 1886 3339
rect 2076 3311 2102 3337
rect 4202 3288 4228 3314
rect 4418 3286 4442 3310
rect 4627 3291 4651 3315
rect 4842 3290 4862 3310
rect 6723 3294 6743 3314
rect 6934 3289 6958 3313
rect 7143 3294 7167 3318
rect 7357 3290 7383 3316
rect 9483 3267 9509 3293
rect 9699 3265 9723 3289
rect 9908 3270 9932 3294
rect 10123 3269 10143 3289
rect 12103 3323 12123 3343
rect 12314 3318 12338 3342
rect 12523 3323 12547 3347
rect 12737 3319 12763 3345
rect 14863 3296 14889 3322
rect 15079 3294 15103 3318
rect 15288 3299 15312 3323
rect 15503 3298 15523 3318
rect 380 3076 400 3096
rect 591 3071 615 3095
rect 800 3076 824 3100
rect 1014 3072 1040 3098
rect 3189 3054 3215 3080
rect 3405 3052 3429 3076
rect 3614 3057 3638 3081
rect 3829 3056 3849 3076
rect 5661 3055 5681 3075
rect 1392 2895 1412 2915
rect 1603 2890 1627 2914
rect 1812 2895 1836 2919
rect 5872 3050 5896 3074
rect 6081 3055 6105 3079
rect 17384 3302 17404 3322
rect 17595 3297 17619 3321
rect 17804 3302 17828 3326
rect 18018 3298 18044 3324
rect 20144 3275 20170 3301
rect 20360 3273 20384 3297
rect 20569 3278 20593 3302
rect 20784 3277 20804 3297
rect 6295 3051 6321 3077
rect 8470 3033 8496 3059
rect 2026 2891 2052 2917
rect 4201 2873 4227 2899
rect 4417 2871 4441 2895
rect 4626 2876 4650 2900
rect 8686 3031 8710 3055
rect 8895 3036 8919 3060
rect 11041 3084 11061 3104
rect 9110 3035 9130 3055
rect 11252 3079 11276 3103
rect 11461 3084 11485 3108
rect 11675 3080 11701 3106
rect 13850 3062 13876 3088
rect 4841 2875 4861 2895
rect 6673 2874 6693 2894
rect 6884 2869 6908 2893
rect 7093 2874 7117 2898
rect 14066 3060 14090 3084
rect 14275 3065 14299 3089
rect 14490 3064 14510 3084
rect 16322 3063 16342 3083
rect 7307 2870 7333 2896
rect 9482 2852 9508 2878
rect 9698 2850 9722 2874
rect 9907 2855 9931 2879
rect 12053 2903 12073 2923
rect 10122 2854 10142 2874
rect 12264 2898 12288 2922
rect 12473 2903 12497 2927
rect 16533 3058 16557 3082
rect 16742 3063 16766 3087
rect 16956 3059 16982 3085
rect 19131 3041 19157 3067
rect 12687 2899 12713 2925
rect 14862 2881 14888 2907
rect 379 2661 399 2681
rect 590 2656 614 2680
rect 799 2661 823 2685
rect 1013 2657 1039 2683
rect 15078 2879 15102 2903
rect 15287 2884 15311 2908
rect 19347 3039 19371 3063
rect 19556 3044 19580 3068
rect 19771 3043 19791 3063
rect 15502 2883 15522 2903
rect 17334 2882 17354 2902
rect 17545 2877 17569 2901
rect 17754 2882 17778 2906
rect 17968 2878 17994 2904
rect 20143 2860 20169 2886
rect 20359 2858 20383 2882
rect 20568 2863 20592 2887
rect 20783 2862 20803 2882
rect 2981 2587 3007 2613
rect 3197 2585 3221 2609
rect 3406 2590 3430 2614
rect 3621 2589 3641 2609
rect 5660 2640 5680 2660
rect 5871 2635 5895 2659
rect 6080 2640 6104 2664
rect 6294 2636 6320 2662
rect 11040 2669 11060 2689
rect 8262 2566 8288 2592
rect 8478 2564 8502 2588
rect 8687 2569 8711 2593
rect 11251 2664 11275 2688
rect 11460 2669 11484 2693
rect 11674 2665 11700 2691
rect 8902 2568 8922 2588
rect 13642 2595 13668 2621
rect 13858 2593 13882 2617
rect 14067 2598 14091 2622
rect 14282 2597 14302 2617
rect 16321 2648 16341 2668
rect 16532 2643 16556 2667
rect 16741 2648 16765 2672
rect 16955 2644 16981 2670
rect 1607 2383 1627 2403
rect 1818 2378 1842 2402
rect 2027 2383 2051 2407
rect 2241 2379 2267 2405
rect 18923 2574 18949 2600
rect 19139 2572 19163 2596
rect 19348 2577 19372 2601
rect 19563 2576 19583 2596
rect 4209 2309 4235 2335
rect 4425 2307 4449 2331
rect 4634 2312 4658 2336
rect 4849 2311 4869 2331
rect 6888 2362 6908 2382
rect 7099 2357 7123 2381
rect 7308 2362 7332 2386
rect 7522 2358 7548 2384
rect 12268 2391 12288 2411
rect 9490 2288 9516 2314
rect 9706 2286 9730 2310
rect 9915 2291 9939 2315
rect 12479 2386 12503 2410
rect 12688 2391 12712 2415
rect 12902 2387 12928 2413
rect 10130 2290 10150 2310
rect 14870 2317 14896 2343
rect 15086 2315 15110 2339
rect 15295 2320 15319 2344
rect 15510 2319 15530 2339
rect 17549 2370 17569 2390
rect 17760 2365 17784 2389
rect 17969 2370 17993 2394
rect 18183 2366 18209 2392
rect 387 2097 407 2117
rect 598 2092 622 2116
rect 807 2097 831 2121
rect 1021 2093 1047 2119
rect 3196 2075 3222 2101
rect 3412 2073 3436 2097
rect 3621 2078 3645 2102
rect 3836 2077 3856 2097
rect 5668 2076 5688 2096
rect 1399 1916 1419 1936
rect 1610 1911 1634 1935
rect 1819 1916 1843 1940
rect 5879 2071 5903 2095
rect 6088 2076 6112 2100
rect 20151 2296 20177 2322
rect 20367 2294 20391 2318
rect 20576 2299 20600 2323
rect 20791 2298 20811 2318
rect 6302 2072 6328 2098
rect 8477 2054 8503 2080
rect 2033 1912 2059 1938
rect 4208 1894 4234 1920
rect 4424 1892 4448 1916
rect 4633 1897 4657 1921
rect 8693 2052 8717 2076
rect 8902 2057 8926 2081
rect 11048 2105 11068 2125
rect 9117 2056 9137 2076
rect 11259 2100 11283 2124
rect 11468 2105 11492 2129
rect 11682 2101 11708 2127
rect 13857 2083 13883 2109
rect 4848 1896 4868 1916
rect 6680 1895 6700 1915
rect 6891 1890 6915 1914
rect 7100 1895 7124 1919
rect 14073 2081 14097 2105
rect 14282 2086 14306 2110
rect 14497 2085 14517 2105
rect 16329 2084 16349 2104
rect 7314 1891 7340 1917
rect 9489 1873 9515 1899
rect 9705 1871 9729 1895
rect 9914 1876 9938 1900
rect 12060 1924 12080 1944
rect 10129 1875 10149 1895
rect 12271 1919 12295 1943
rect 12480 1924 12504 1948
rect 16540 2079 16564 2103
rect 16749 2084 16773 2108
rect 16963 2080 16989 2106
rect 19138 2062 19164 2088
rect 12694 1920 12720 1946
rect 14869 1902 14895 1928
rect 386 1682 406 1702
rect 597 1677 621 1701
rect 806 1682 830 1706
rect 1020 1678 1046 1704
rect 3146 1655 3172 1681
rect 3362 1653 3386 1677
rect 3571 1658 3595 1682
rect 3786 1657 3806 1677
rect 15085 1900 15109 1924
rect 15294 1905 15318 1929
rect 19354 2060 19378 2084
rect 19563 2065 19587 2089
rect 19778 2064 19798 2084
rect 15509 1904 15529 1924
rect 17341 1903 17361 1923
rect 17552 1898 17576 1922
rect 17761 1903 17785 1927
rect 17975 1899 18001 1925
rect 20150 1881 20176 1907
rect 20366 1879 20390 1903
rect 20575 1884 20599 1908
rect 20790 1883 20810 1903
rect 5667 1661 5687 1681
rect 5878 1656 5902 1680
rect 6087 1661 6111 1685
rect 6301 1657 6327 1683
rect 8427 1634 8453 1660
rect 8643 1632 8667 1656
rect 8852 1637 8876 1661
rect 9067 1636 9087 1656
rect 11047 1690 11067 1710
rect 11258 1685 11282 1709
rect 11467 1690 11491 1714
rect 11681 1686 11707 1712
rect 13807 1663 13833 1689
rect 14023 1661 14047 1685
rect 14232 1666 14256 1690
rect 14447 1665 14467 1685
rect 16328 1669 16348 1689
rect 16539 1664 16563 1688
rect 16748 1669 16772 1693
rect 16962 1665 16988 1691
rect 19088 1642 19114 1668
rect 19304 1640 19328 1664
rect 19513 1645 19537 1669
rect 19728 1644 19748 1664
rect 1454 1355 1474 1375
rect 1665 1350 1689 1374
rect 1874 1355 1898 1379
rect 2088 1351 2114 1377
rect 4214 1328 4240 1354
rect 4430 1326 4454 1350
rect 4639 1331 4663 1355
rect 4854 1330 4874 1350
rect 6735 1334 6755 1354
rect 6946 1329 6970 1353
rect 7155 1334 7179 1358
rect 7369 1330 7395 1356
rect 9495 1307 9521 1333
rect 9711 1305 9735 1329
rect 9920 1310 9944 1334
rect 10135 1309 10155 1329
rect 12115 1363 12135 1383
rect 12326 1358 12350 1382
rect 12535 1363 12559 1387
rect 12749 1359 12775 1385
rect 14875 1336 14901 1362
rect 15091 1334 15115 1358
rect 15300 1339 15324 1363
rect 15515 1338 15535 1358
rect 392 1116 412 1136
rect 603 1111 627 1135
rect 812 1116 836 1140
rect 1026 1112 1052 1138
rect 3201 1094 3227 1120
rect 3417 1092 3441 1116
rect 3626 1097 3650 1121
rect 3841 1096 3861 1116
rect 5673 1095 5693 1115
rect 1404 935 1424 955
rect 1615 930 1639 954
rect 1824 935 1848 959
rect 5884 1090 5908 1114
rect 6093 1095 6117 1119
rect 17396 1342 17416 1362
rect 17607 1337 17631 1361
rect 17816 1342 17840 1366
rect 18030 1338 18056 1364
rect 20156 1315 20182 1341
rect 20372 1313 20396 1337
rect 20581 1318 20605 1342
rect 20796 1317 20816 1337
rect 6307 1091 6333 1117
rect 8482 1073 8508 1099
rect 2038 931 2064 957
rect 4213 913 4239 939
rect 4429 911 4453 935
rect 4638 916 4662 940
rect 8698 1071 8722 1095
rect 8907 1076 8931 1100
rect 11053 1124 11073 1144
rect 9122 1075 9142 1095
rect 11264 1119 11288 1143
rect 11473 1124 11497 1148
rect 11687 1120 11713 1146
rect 13862 1102 13888 1128
rect 4853 915 4873 935
rect 6685 914 6705 934
rect 6896 909 6920 933
rect 7105 914 7129 938
rect 14078 1100 14102 1124
rect 14287 1105 14311 1129
rect 14502 1104 14522 1124
rect 16334 1103 16354 1123
rect 7319 910 7345 936
rect 9494 892 9520 918
rect 9710 890 9734 914
rect 9919 895 9943 919
rect 12065 943 12085 963
rect 10134 894 10154 914
rect 12276 938 12300 962
rect 12485 943 12509 967
rect 16545 1098 16569 1122
rect 16754 1103 16778 1127
rect 16968 1099 16994 1125
rect 19143 1081 19169 1107
rect 12699 939 12725 965
rect 14874 921 14900 947
rect 391 701 411 721
rect 602 696 626 720
rect 811 701 835 725
rect 1025 697 1051 723
rect 15090 919 15114 943
rect 15299 924 15323 948
rect 19359 1079 19383 1103
rect 19568 1084 19592 1108
rect 19783 1083 19803 1103
rect 15514 923 15534 943
rect 17346 922 17366 942
rect 17557 917 17581 941
rect 17766 922 17790 946
rect 17980 918 18006 944
rect 20155 900 20181 926
rect 20371 898 20395 922
rect 20580 903 20604 927
rect 20795 902 20815 922
rect 5672 680 5692 700
rect 5883 675 5907 699
rect 6092 680 6116 704
rect 6306 676 6332 702
rect 11052 709 11072 729
rect 11263 704 11287 728
rect 11472 709 11496 733
rect 11686 705 11712 731
rect 16333 688 16353 708
rect 16544 683 16568 707
rect 16753 688 16777 712
rect 16967 684 16993 710
rect 1794 220 1814 240
rect 2005 215 2029 239
rect 2214 220 2238 244
rect 2428 216 2454 242
rect 7075 199 7095 219
rect 4884 132 4904 152
rect 5095 127 5119 151
rect 5304 132 5328 156
rect 7286 194 7310 218
rect 7495 199 7519 223
rect 7709 195 7735 221
rect 12455 228 12475 248
rect 12666 223 12690 247
rect 12875 228 12899 252
rect 13089 224 13115 250
rect 5518 128 5544 154
rect 10145 125 10165 145
rect 10356 120 10380 144
rect 10565 125 10589 149
rect 17736 207 17756 227
rect 10779 121 10805 147
rect 15545 140 15565 160
rect 15756 135 15780 159
rect 15965 140 15989 164
rect 17947 202 17971 226
rect 18156 207 18180 231
rect 18370 203 18396 229
rect 16179 136 16205 162
<< ndiffres >>
rect 97 8317 154 8336
rect 10758 8325 10815 8344
rect 10758 8322 10779 8325
rect 97 8314 118 8317
rect 3 8299 118 8314
rect 136 8299 154 8317
rect 3 8276 154 8299
rect 5378 8296 5435 8315
rect 5378 8293 5399 8296
rect 3 8240 45 8276
rect 2 8239 102 8240
rect 2 8218 158 8239
rect 5028 8268 5089 8284
rect 5284 8278 5399 8293
rect 5417 8278 5435 8296
rect 5028 8264 5184 8268
rect 5028 8246 5048 8264
rect 5066 8246 5184 8264
rect 2 8200 120 8218
rect 138 8200 158 8218
rect 2 8196 158 8200
rect 97 8180 158 8196
rect 5028 8225 5184 8246
rect 5084 8224 5184 8225
rect 5284 8255 5435 8278
rect 10664 8307 10779 8322
rect 10797 8307 10815 8325
rect 10664 8284 10815 8307
rect 16039 8304 16096 8323
rect 16039 8301 16060 8304
rect 5141 8188 5183 8224
rect 5284 8219 5326 8255
rect 5032 8165 5183 8188
rect 5283 8218 5383 8219
rect 5283 8197 5439 8218
rect 10309 8247 10370 8263
rect 10664 8248 10706 8284
rect 10663 8247 10763 8248
rect 10309 8243 10465 8247
rect 10309 8225 10329 8243
rect 10347 8225 10465 8243
rect 5283 8179 5401 8197
rect 5419 8179 5439 8197
rect 5283 8175 5439 8179
rect 95 8103 152 8122
rect 95 8100 116 8103
rect 1 8085 116 8100
rect 134 8085 152 8103
rect 1 8062 152 8085
rect 1 8026 43 8062
rect 0 8025 100 8026
rect 0 8004 156 8025
rect 5032 8147 5050 8165
rect 5068 8150 5183 8165
rect 5378 8159 5439 8175
rect 5068 8147 5089 8150
rect 5032 8128 5089 8147
rect 10309 8204 10465 8225
rect 10663 8226 10819 8247
rect 15689 8276 15750 8292
rect 15945 8286 16060 8301
rect 16078 8286 16096 8304
rect 15689 8272 15845 8276
rect 15689 8254 15709 8272
rect 15727 8254 15845 8272
rect 10663 8208 10781 8226
rect 10799 8208 10819 8226
rect 10663 8204 10819 8208
rect 10365 8203 10465 8204
rect 10422 8167 10464 8203
rect 10758 8188 10819 8204
rect 15689 8233 15845 8254
rect 15745 8232 15845 8233
rect 15945 8263 16096 8286
rect 15802 8196 15844 8232
rect 15945 8227 15987 8263
rect 15693 8173 15844 8196
rect 15944 8226 16044 8227
rect 15944 8205 16100 8226
rect 20970 8255 21031 8271
rect 20970 8251 21126 8255
rect 20970 8233 20990 8251
rect 21008 8233 21126 8251
rect 15944 8187 16062 8205
rect 16080 8187 16100 8205
rect 15944 8183 16100 8187
rect 10313 8144 10464 8167
rect 5035 8067 5096 8083
rect 5376 8082 5433 8101
rect 5376 8079 5397 8082
rect 5035 8063 5191 8067
rect 5035 8045 5055 8063
rect 5073 8045 5191 8063
rect 0 7986 118 8004
rect 136 7986 156 8004
rect 0 7982 156 7986
rect 95 7966 156 7982
rect 5035 8024 5191 8045
rect 5091 8023 5191 8024
rect 5282 8064 5397 8079
rect 5415 8064 5433 8082
rect 5282 8041 5433 8064
rect 5148 7987 5190 8023
rect 5282 8005 5324 8041
rect 5039 7964 5190 7987
rect 5039 7946 5057 7964
rect 5075 7949 5190 7964
rect 5281 8004 5381 8005
rect 5281 7983 5437 8004
rect 10313 8126 10331 8144
rect 10349 8129 10464 8144
rect 10349 8126 10370 8129
rect 10313 8107 10370 8126
rect 10756 8111 10813 8130
rect 10756 8108 10777 8111
rect 10662 8093 10777 8108
rect 10795 8093 10813 8111
rect 10662 8070 10813 8093
rect 10316 8046 10377 8062
rect 10316 8042 10472 8046
rect 10316 8024 10336 8042
rect 10354 8024 10472 8042
rect 10662 8034 10704 8070
rect 5281 7965 5399 7983
rect 5417 7965 5437 7983
rect 5281 7961 5437 7965
rect 5075 7946 5096 7949
rect 5039 7927 5096 7946
rect 5376 7945 5437 7961
rect 95 7821 152 7840
rect 95 7818 116 7821
rect 1 7803 116 7818
rect 134 7803 152 7821
rect 1 7780 152 7803
rect 1 7744 43 7780
rect 10316 8003 10472 8024
rect 10372 8002 10472 8003
rect 10661 8033 10761 8034
rect 10661 8012 10817 8033
rect 15693 8155 15711 8173
rect 15729 8158 15844 8173
rect 16039 8167 16100 8183
rect 15729 8155 15750 8158
rect 15693 8136 15750 8155
rect 20970 8212 21126 8233
rect 21026 8211 21126 8212
rect 21083 8175 21125 8211
rect 20974 8152 21125 8175
rect 15696 8075 15757 8091
rect 16037 8090 16094 8109
rect 16037 8087 16058 8090
rect 15696 8071 15852 8075
rect 15696 8053 15716 8071
rect 15734 8053 15852 8071
rect 0 7743 100 7744
rect 0 7722 156 7743
rect 10429 7966 10471 8002
rect 10661 7994 10779 8012
rect 10797 7994 10817 8012
rect 10661 7990 10817 7994
rect 10756 7974 10817 7990
rect 10320 7943 10471 7966
rect 15696 8032 15852 8053
rect 15752 8031 15852 8032
rect 15943 8072 16058 8087
rect 16076 8072 16094 8090
rect 15943 8049 16094 8072
rect 10320 7925 10338 7943
rect 10356 7928 10471 7943
rect 10356 7925 10377 7928
rect 10320 7906 10377 7925
rect 5035 7785 5096 7801
rect 5376 7800 5433 7819
rect 5376 7797 5397 7800
rect 5035 7781 5191 7785
rect 5035 7763 5055 7781
rect 5073 7763 5191 7781
rect 0 7704 118 7722
rect 136 7704 156 7722
rect 0 7700 156 7704
rect 95 7684 156 7700
rect 102 7620 159 7639
rect 102 7617 123 7620
rect 8 7602 123 7617
rect 141 7602 159 7620
rect 5035 7742 5191 7763
rect 5091 7741 5191 7742
rect 5282 7782 5397 7797
rect 5415 7782 5433 7800
rect 5282 7759 5433 7782
rect 5148 7705 5190 7741
rect 5282 7723 5324 7759
rect 15809 7995 15851 8031
rect 15943 8013 15985 8049
rect 15700 7972 15851 7995
rect 15700 7954 15718 7972
rect 15736 7957 15851 7972
rect 15942 8012 16042 8013
rect 15942 7991 16098 8012
rect 20974 8134 20992 8152
rect 21010 8137 21125 8152
rect 21010 8134 21031 8137
rect 20974 8115 21031 8134
rect 20977 8054 21038 8070
rect 20977 8050 21133 8054
rect 20977 8032 20997 8050
rect 21015 8032 21133 8050
rect 15942 7973 16060 7991
rect 16078 7973 16098 7991
rect 15942 7969 16098 7973
rect 15736 7954 15757 7957
rect 15700 7935 15757 7954
rect 16037 7953 16098 7969
rect 10756 7829 10813 7848
rect 10756 7826 10777 7829
rect 10662 7811 10777 7826
rect 10795 7811 10813 7829
rect 5039 7682 5190 7705
rect 5039 7664 5057 7682
rect 5075 7667 5190 7682
rect 5281 7722 5381 7723
rect 5281 7701 5437 7722
rect 10662 7788 10813 7811
rect 10316 7764 10377 7780
rect 10316 7760 10472 7764
rect 10316 7742 10336 7760
rect 10354 7742 10472 7760
rect 10662 7752 10704 7788
rect 20977 8011 21133 8032
rect 21033 8010 21133 8011
rect 5281 7683 5399 7701
rect 5417 7683 5437 7701
rect 5281 7679 5437 7683
rect 5075 7664 5096 7667
rect 5039 7645 5096 7664
rect 5376 7663 5437 7679
rect 8 7579 159 7602
rect 8 7543 50 7579
rect 7 7542 107 7543
rect 7 7521 163 7542
rect 5383 7599 5440 7618
rect 5383 7596 5404 7599
rect 7 7503 125 7521
rect 143 7503 163 7521
rect 7 7499 163 7503
rect 102 7483 163 7499
rect 5033 7571 5094 7587
rect 5289 7581 5404 7596
rect 5422 7581 5440 7599
rect 10316 7721 10472 7742
rect 10372 7720 10472 7721
rect 10661 7751 10761 7752
rect 10661 7730 10817 7751
rect 21090 7974 21132 8010
rect 20981 7951 21132 7974
rect 20981 7933 20999 7951
rect 21017 7936 21132 7951
rect 21017 7933 21038 7936
rect 20981 7914 21038 7933
rect 15696 7793 15757 7809
rect 16037 7808 16094 7827
rect 16037 7805 16058 7808
rect 15696 7789 15852 7793
rect 15696 7771 15716 7789
rect 15734 7771 15852 7789
rect 10429 7684 10471 7720
rect 10661 7712 10779 7730
rect 10797 7712 10817 7730
rect 10661 7708 10817 7712
rect 10756 7692 10817 7708
rect 10320 7661 10471 7684
rect 10320 7643 10338 7661
rect 10356 7646 10471 7661
rect 10356 7643 10377 7646
rect 10320 7624 10377 7643
rect 10763 7628 10820 7647
rect 10763 7625 10784 7628
rect 10669 7610 10784 7625
rect 10802 7610 10820 7628
rect 15696 7750 15852 7771
rect 15752 7749 15852 7750
rect 15943 7790 16058 7805
rect 16076 7790 16094 7808
rect 15943 7767 16094 7790
rect 15809 7713 15851 7749
rect 15943 7731 15985 7767
rect 15700 7690 15851 7713
rect 15700 7672 15718 7690
rect 15736 7675 15851 7690
rect 15942 7730 16042 7731
rect 15942 7709 16098 7730
rect 20977 7772 21038 7788
rect 20977 7768 21133 7772
rect 20977 7750 20997 7768
rect 21015 7750 21133 7768
rect 15942 7691 16060 7709
rect 16078 7691 16098 7709
rect 15942 7687 16098 7691
rect 15736 7672 15757 7675
rect 15700 7653 15757 7672
rect 16037 7671 16098 7687
rect 5033 7567 5189 7571
rect 5033 7549 5053 7567
rect 5071 7549 5189 7567
rect 5033 7528 5189 7549
rect 5089 7527 5189 7528
rect 5289 7558 5440 7581
rect 5146 7491 5188 7527
rect 5289 7522 5331 7558
rect 5037 7468 5188 7491
rect 5288 7521 5388 7522
rect 5288 7500 5444 7521
rect 10669 7587 10820 7610
rect 5288 7482 5406 7500
rect 5424 7482 5444 7500
rect 5288 7478 5444 7482
rect 5037 7450 5055 7468
rect 5073 7453 5188 7468
rect 5383 7462 5444 7478
rect 10314 7550 10375 7566
rect 10669 7551 10711 7587
rect 10668 7550 10768 7551
rect 10314 7546 10470 7550
rect 10314 7528 10334 7546
rect 10352 7528 10470 7546
rect 10314 7507 10470 7528
rect 10668 7529 10824 7550
rect 16044 7607 16101 7626
rect 16044 7604 16065 7607
rect 10668 7511 10786 7529
rect 10804 7511 10824 7529
rect 10668 7507 10824 7511
rect 10370 7506 10470 7507
rect 5073 7450 5094 7453
rect 5037 7431 5094 7450
rect 10427 7470 10469 7506
rect 10763 7491 10824 7507
rect 15694 7579 15755 7595
rect 15950 7589 16065 7604
rect 16083 7589 16101 7607
rect 20977 7729 21133 7750
rect 21033 7728 21133 7729
rect 21090 7692 21132 7728
rect 20981 7669 21132 7692
rect 20981 7651 20999 7669
rect 21017 7654 21132 7669
rect 21017 7651 21038 7654
rect 20981 7632 21038 7651
rect 15694 7575 15850 7579
rect 15694 7557 15714 7575
rect 15732 7557 15850 7575
rect 15694 7536 15850 7557
rect 15750 7535 15850 7536
rect 15950 7566 16101 7589
rect 10318 7447 10469 7470
rect 10318 7429 10336 7447
rect 10354 7432 10469 7447
rect 10354 7429 10375 7432
rect 10318 7410 10375 7429
rect 15807 7499 15849 7535
rect 15950 7530 15992 7566
rect 15698 7476 15849 7499
rect 15949 7529 16049 7530
rect 15949 7508 16105 7529
rect 15949 7490 16067 7508
rect 16085 7490 16105 7508
rect 15949 7486 16105 7490
rect 15698 7458 15716 7476
rect 15734 7461 15849 7476
rect 16044 7470 16105 7486
rect 20975 7558 21036 7574
rect 20975 7554 21131 7558
rect 20975 7536 20995 7554
rect 21013 7536 21131 7554
rect 20975 7515 21131 7536
rect 21031 7514 21131 7515
rect 15734 7458 15755 7461
rect 15698 7439 15755 7458
rect 21088 7478 21130 7514
rect 20979 7455 21130 7478
rect 20979 7437 20997 7455
rect 21015 7440 21130 7455
rect 21015 7437 21036 7440
rect 20979 7418 21036 7437
rect 102 7336 159 7355
rect 102 7333 123 7336
rect 8 7318 123 7333
rect 141 7318 159 7336
rect 8 7295 159 7318
rect 8 7259 50 7295
rect 5383 7315 5440 7334
rect 5383 7312 5404 7315
rect 7 7258 107 7259
rect 7 7237 163 7258
rect 7 7219 125 7237
rect 143 7219 163 7237
rect 7 7215 163 7219
rect 102 7199 163 7215
rect 5033 7287 5094 7303
rect 5289 7297 5404 7312
rect 5422 7297 5440 7315
rect 5033 7283 5189 7287
rect 5033 7265 5053 7283
rect 5071 7265 5189 7283
rect 5033 7244 5189 7265
rect 5089 7243 5189 7244
rect 5289 7274 5440 7297
rect 5146 7207 5188 7243
rect 5289 7238 5331 7274
rect 10763 7344 10820 7363
rect 10763 7341 10784 7344
rect 10669 7326 10784 7341
rect 10802 7326 10820 7344
rect 10669 7303 10820 7326
rect 5037 7184 5188 7207
rect 5288 7237 5388 7238
rect 5288 7216 5444 7237
rect 5288 7198 5406 7216
rect 5424 7198 5444 7216
rect 5288 7194 5444 7198
rect 100 7122 157 7141
rect 100 7119 121 7122
rect 6 7104 121 7119
rect 139 7104 157 7122
rect 6 7081 157 7104
rect 6 7045 48 7081
rect 5 7044 105 7045
rect 5 7023 161 7044
rect 5037 7166 5055 7184
rect 5073 7169 5188 7184
rect 5383 7178 5444 7194
rect 10314 7266 10375 7282
rect 10669 7267 10711 7303
rect 16044 7323 16101 7342
rect 16044 7320 16065 7323
rect 10668 7266 10768 7267
rect 10314 7262 10470 7266
rect 10314 7244 10334 7262
rect 10352 7244 10470 7262
rect 5073 7166 5094 7169
rect 5037 7147 5094 7166
rect 10314 7223 10470 7244
rect 10668 7245 10824 7266
rect 10668 7227 10786 7245
rect 10804 7227 10824 7245
rect 10668 7223 10824 7227
rect 10370 7222 10470 7223
rect 10427 7186 10469 7222
rect 10763 7207 10824 7223
rect 15694 7295 15755 7311
rect 15950 7305 16065 7320
rect 16083 7305 16101 7323
rect 15694 7291 15850 7295
rect 15694 7273 15714 7291
rect 15732 7273 15850 7291
rect 10318 7163 10469 7186
rect 15694 7252 15850 7273
rect 15750 7251 15850 7252
rect 15950 7282 16101 7305
rect 15807 7215 15849 7251
rect 15950 7246 15992 7282
rect 15698 7192 15849 7215
rect 15949 7245 16049 7246
rect 15949 7224 16105 7245
rect 15949 7206 16067 7224
rect 16085 7206 16105 7224
rect 15949 7202 16105 7206
rect 5040 7086 5101 7102
rect 5381 7101 5438 7120
rect 5381 7098 5402 7101
rect 5040 7082 5196 7086
rect 5040 7064 5060 7082
rect 5078 7064 5196 7082
rect 5 7005 123 7023
rect 141 7005 161 7023
rect 5 7001 161 7005
rect 100 6985 161 7001
rect 5040 7043 5196 7064
rect 5096 7042 5196 7043
rect 5287 7083 5402 7098
rect 5420 7083 5438 7101
rect 5287 7060 5438 7083
rect 5153 7006 5195 7042
rect 5287 7024 5329 7060
rect 5044 6983 5195 7006
rect 5044 6965 5062 6983
rect 5080 6968 5195 6983
rect 5286 7023 5386 7024
rect 5286 7002 5442 7023
rect 10318 7145 10336 7163
rect 10354 7148 10469 7163
rect 10354 7145 10375 7148
rect 10318 7126 10375 7145
rect 10761 7130 10818 7149
rect 10761 7127 10782 7130
rect 10667 7112 10782 7127
rect 10800 7112 10818 7130
rect 10667 7089 10818 7112
rect 10321 7065 10382 7081
rect 10321 7061 10477 7065
rect 10321 7043 10341 7061
rect 10359 7043 10477 7061
rect 10667 7053 10709 7089
rect 5286 6984 5404 7002
rect 5422 6984 5442 7002
rect 5286 6980 5442 6984
rect 5080 6965 5101 6968
rect 5044 6946 5101 6965
rect 5381 6964 5442 6980
rect 100 6840 157 6859
rect 100 6837 121 6840
rect 6 6822 121 6837
rect 139 6822 157 6840
rect 6 6799 157 6822
rect 6 6763 48 6799
rect 10321 7022 10477 7043
rect 10377 7021 10477 7022
rect 10666 7052 10766 7053
rect 10666 7031 10822 7052
rect 15698 7174 15716 7192
rect 15734 7177 15849 7192
rect 16044 7186 16105 7202
rect 20975 7274 21036 7290
rect 20975 7270 21131 7274
rect 20975 7252 20995 7270
rect 21013 7252 21131 7270
rect 15734 7174 15755 7177
rect 15698 7155 15755 7174
rect 20975 7231 21131 7252
rect 21031 7230 21131 7231
rect 21088 7194 21130 7230
rect 20979 7171 21130 7194
rect 15701 7094 15762 7110
rect 16042 7109 16099 7128
rect 16042 7106 16063 7109
rect 15701 7090 15857 7094
rect 15701 7072 15721 7090
rect 15739 7072 15857 7090
rect 5 6762 105 6763
rect 5 6741 161 6762
rect 10434 6985 10476 7021
rect 10666 7013 10784 7031
rect 10802 7013 10822 7031
rect 10666 7009 10822 7013
rect 10761 6993 10822 7009
rect 10325 6962 10476 6985
rect 15701 7051 15857 7072
rect 15757 7050 15857 7051
rect 15948 7091 16063 7106
rect 16081 7091 16099 7109
rect 15948 7068 16099 7091
rect 10325 6944 10343 6962
rect 10361 6947 10476 6962
rect 10361 6944 10382 6947
rect 10325 6925 10382 6944
rect 5040 6804 5101 6820
rect 5381 6819 5438 6838
rect 5381 6816 5402 6819
rect 5040 6800 5196 6804
rect 5040 6782 5060 6800
rect 5078 6782 5196 6800
rect 5 6723 123 6741
rect 141 6723 161 6741
rect 5 6719 161 6723
rect 100 6703 161 6719
rect 107 6639 164 6658
rect 107 6636 128 6639
rect 13 6621 128 6636
rect 146 6621 164 6639
rect 5040 6761 5196 6782
rect 5096 6760 5196 6761
rect 5287 6801 5402 6816
rect 5420 6801 5438 6819
rect 5287 6778 5438 6801
rect 5153 6724 5195 6760
rect 5287 6742 5329 6778
rect 15814 7014 15856 7050
rect 15948 7032 15990 7068
rect 15705 6991 15856 7014
rect 15705 6973 15723 6991
rect 15741 6976 15856 6991
rect 15947 7031 16047 7032
rect 15947 7010 16103 7031
rect 20979 7153 20997 7171
rect 21015 7156 21130 7171
rect 21015 7153 21036 7156
rect 20979 7134 21036 7153
rect 20982 7073 21043 7089
rect 20982 7069 21138 7073
rect 20982 7051 21002 7069
rect 21020 7051 21138 7069
rect 15947 6992 16065 7010
rect 16083 6992 16103 7010
rect 15947 6988 16103 6992
rect 15741 6973 15762 6976
rect 15705 6954 15762 6973
rect 16042 6972 16103 6988
rect 10761 6848 10818 6867
rect 10761 6845 10782 6848
rect 10667 6830 10782 6845
rect 10800 6830 10818 6848
rect 5044 6701 5195 6724
rect 5044 6683 5062 6701
rect 5080 6686 5195 6701
rect 5286 6741 5386 6742
rect 5286 6720 5442 6741
rect 10667 6807 10818 6830
rect 10321 6783 10382 6799
rect 10321 6779 10477 6783
rect 10321 6761 10341 6779
rect 10359 6761 10477 6779
rect 10667 6771 10709 6807
rect 20982 7030 21138 7051
rect 21038 7029 21138 7030
rect 5286 6702 5404 6720
rect 5422 6702 5442 6720
rect 5286 6698 5442 6702
rect 5080 6683 5101 6686
rect 5044 6664 5101 6683
rect 5381 6682 5442 6698
rect 13 6598 164 6621
rect 13 6562 55 6598
rect 12 6561 112 6562
rect 12 6540 168 6561
rect 5388 6618 5445 6637
rect 5388 6615 5409 6618
rect 5038 6590 5099 6606
rect 5294 6600 5409 6615
rect 5427 6600 5445 6618
rect 10321 6740 10477 6761
rect 10377 6739 10477 6740
rect 10666 6770 10766 6771
rect 10666 6749 10822 6770
rect 21095 6993 21137 7029
rect 20986 6970 21137 6993
rect 20986 6952 21004 6970
rect 21022 6955 21137 6970
rect 21022 6952 21043 6955
rect 20986 6933 21043 6952
rect 15701 6812 15762 6828
rect 16042 6827 16099 6846
rect 16042 6824 16063 6827
rect 15701 6808 15857 6812
rect 15701 6790 15721 6808
rect 15739 6790 15857 6808
rect 10434 6703 10476 6739
rect 10666 6731 10784 6749
rect 10802 6731 10822 6749
rect 10666 6727 10822 6731
rect 10761 6711 10822 6727
rect 10325 6680 10476 6703
rect 10325 6662 10343 6680
rect 10361 6665 10476 6680
rect 10361 6662 10382 6665
rect 10325 6643 10382 6662
rect 10768 6647 10825 6666
rect 10768 6644 10789 6647
rect 10674 6629 10789 6644
rect 10807 6629 10825 6647
rect 15701 6769 15857 6790
rect 15757 6768 15857 6769
rect 15948 6809 16063 6824
rect 16081 6809 16099 6827
rect 15948 6786 16099 6809
rect 15814 6732 15856 6768
rect 15948 6750 15990 6786
rect 15705 6709 15856 6732
rect 15705 6691 15723 6709
rect 15741 6694 15856 6709
rect 15947 6749 16047 6750
rect 15947 6728 16103 6749
rect 20982 6791 21043 6807
rect 20982 6787 21138 6791
rect 20982 6769 21002 6787
rect 21020 6769 21138 6787
rect 15947 6710 16065 6728
rect 16083 6710 16103 6728
rect 15947 6706 16103 6710
rect 15741 6691 15762 6694
rect 15705 6672 15762 6691
rect 16042 6690 16103 6706
rect 10674 6606 10825 6629
rect 5038 6586 5194 6590
rect 5038 6568 5058 6586
rect 5076 6568 5194 6586
rect 12 6522 130 6540
rect 148 6522 168 6540
rect 12 6518 168 6522
rect 107 6502 168 6518
rect 5038 6547 5194 6568
rect 5094 6546 5194 6547
rect 5294 6577 5445 6600
rect 5151 6510 5193 6546
rect 5294 6541 5336 6577
rect 5042 6487 5193 6510
rect 5293 6540 5393 6541
rect 5293 6519 5449 6540
rect 10319 6569 10380 6585
rect 10674 6570 10716 6606
rect 10673 6569 10773 6570
rect 10319 6565 10475 6569
rect 10319 6547 10339 6565
rect 10357 6547 10475 6565
rect 5293 6501 5411 6519
rect 5429 6501 5449 6519
rect 5293 6497 5449 6501
rect 109 6357 166 6376
rect 109 6354 130 6357
rect 15 6339 130 6354
rect 148 6339 166 6357
rect 5042 6469 5060 6487
rect 5078 6472 5193 6487
rect 5388 6481 5449 6497
rect 5078 6469 5099 6472
rect 5042 6450 5099 6469
rect 10319 6526 10475 6547
rect 10673 6548 10829 6569
rect 16049 6626 16106 6645
rect 16049 6623 16070 6626
rect 15699 6598 15760 6614
rect 15955 6608 16070 6623
rect 16088 6608 16106 6626
rect 20982 6748 21138 6769
rect 21038 6747 21138 6748
rect 21095 6711 21137 6747
rect 20986 6688 21137 6711
rect 20986 6670 21004 6688
rect 21022 6673 21137 6688
rect 21022 6670 21043 6673
rect 20986 6651 21043 6670
rect 15699 6594 15855 6598
rect 15699 6576 15719 6594
rect 15737 6576 15855 6594
rect 10673 6530 10791 6548
rect 10809 6530 10829 6548
rect 10673 6526 10829 6530
rect 10375 6525 10475 6526
rect 10432 6489 10474 6525
rect 10768 6510 10829 6526
rect 10323 6466 10474 6489
rect 15699 6555 15855 6576
rect 15755 6554 15855 6555
rect 15955 6585 16106 6608
rect 15812 6518 15854 6554
rect 15955 6549 15997 6585
rect 15703 6495 15854 6518
rect 15954 6548 16054 6549
rect 15954 6527 16110 6548
rect 20980 6577 21041 6593
rect 20980 6573 21136 6577
rect 20980 6555 21000 6573
rect 21018 6555 21136 6573
rect 15954 6509 16072 6527
rect 16090 6509 16110 6527
rect 15954 6505 16110 6509
rect 15 6316 166 6339
rect 15 6280 57 6316
rect 14 6279 114 6280
rect 14 6258 170 6279
rect 5390 6336 5447 6355
rect 5390 6333 5411 6336
rect 5040 6308 5101 6324
rect 5296 6318 5411 6333
rect 5429 6318 5447 6336
rect 10323 6448 10341 6466
rect 10359 6451 10474 6466
rect 10359 6448 10380 6451
rect 10323 6429 10380 6448
rect 10770 6365 10827 6384
rect 10770 6362 10791 6365
rect 10676 6347 10791 6362
rect 10809 6347 10827 6365
rect 15703 6477 15721 6495
rect 15739 6480 15854 6495
rect 16049 6489 16110 6505
rect 15739 6477 15760 6480
rect 15703 6458 15760 6477
rect 20980 6534 21136 6555
rect 21036 6533 21136 6534
rect 21093 6497 21135 6533
rect 20984 6474 21135 6497
rect 5040 6304 5196 6308
rect 5040 6286 5060 6304
rect 5078 6286 5196 6304
rect 14 6240 132 6258
rect 150 6240 170 6258
rect 14 6236 170 6240
rect 109 6220 170 6236
rect 5040 6265 5196 6286
rect 5096 6264 5196 6265
rect 5296 6295 5447 6318
rect 5153 6228 5195 6264
rect 5296 6259 5338 6295
rect 5044 6205 5195 6228
rect 5295 6258 5395 6259
rect 5295 6237 5451 6258
rect 10676 6324 10827 6347
rect 10321 6287 10382 6303
rect 10676 6288 10718 6324
rect 10675 6287 10775 6288
rect 10321 6283 10477 6287
rect 10321 6265 10341 6283
rect 10359 6265 10477 6283
rect 5295 6219 5413 6237
rect 5431 6219 5451 6237
rect 5295 6215 5451 6219
rect 107 6143 164 6162
rect 107 6140 128 6143
rect 13 6125 128 6140
rect 146 6125 164 6143
rect 13 6102 164 6125
rect 13 6066 55 6102
rect 12 6065 112 6066
rect 12 6044 168 6065
rect 5044 6187 5062 6205
rect 5080 6190 5195 6205
rect 5390 6199 5451 6215
rect 5080 6187 5101 6190
rect 5044 6168 5101 6187
rect 10321 6244 10477 6265
rect 10675 6266 10831 6287
rect 16051 6344 16108 6363
rect 16051 6341 16072 6344
rect 15701 6316 15762 6332
rect 15957 6326 16072 6341
rect 16090 6326 16108 6344
rect 20984 6456 21002 6474
rect 21020 6459 21135 6474
rect 21020 6456 21041 6459
rect 20984 6437 21041 6456
rect 15701 6312 15857 6316
rect 15701 6294 15721 6312
rect 15739 6294 15857 6312
rect 10675 6248 10793 6266
rect 10811 6248 10831 6266
rect 10675 6244 10831 6248
rect 10377 6243 10477 6244
rect 10434 6207 10476 6243
rect 10770 6228 10831 6244
rect 15701 6273 15857 6294
rect 15757 6272 15857 6273
rect 15957 6303 16108 6326
rect 15814 6236 15856 6272
rect 15957 6267 15999 6303
rect 15705 6213 15856 6236
rect 15956 6266 16056 6267
rect 15956 6245 16112 6266
rect 20982 6295 21043 6311
rect 20982 6291 21138 6295
rect 20982 6273 21002 6291
rect 21020 6273 21138 6291
rect 15956 6227 16074 6245
rect 16092 6227 16112 6245
rect 15956 6223 16112 6227
rect 10325 6184 10476 6207
rect 5047 6107 5108 6123
rect 5388 6122 5445 6141
rect 5388 6119 5409 6122
rect 5047 6103 5203 6107
rect 5047 6085 5067 6103
rect 5085 6085 5203 6103
rect 12 6026 130 6044
rect 148 6026 168 6044
rect 12 6022 168 6026
rect 107 6006 168 6022
rect 5047 6064 5203 6085
rect 5103 6063 5203 6064
rect 5294 6104 5409 6119
rect 5427 6104 5445 6122
rect 5294 6081 5445 6104
rect 5160 6027 5202 6063
rect 5294 6045 5336 6081
rect 5051 6004 5202 6027
rect 5051 5986 5069 6004
rect 5087 5989 5202 6004
rect 5293 6044 5393 6045
rect 5293 6023 5449 6044
rect 10325 6166 10343 6184
rect 10361 6169 10476 6184
rect 10361 6166 10382 6169
rect 10325 6147 10382 6166
rect 10768 6151 10825 6170
rect 10768 6148 10789 6151
rect 10674 6133 10789 6148
rect 10807 6133 10825 6151
rect 10674 6110 10825 6133
rect 10328 6086 10389 6102
rect 10328 6082 10484 6086
rect 10328 6064 10348 6082
rect 10366 6064 10484 6082
rect 10674 6074 10716 6110
rect 5293 6005 5411 6023
rect 5429 6005 5449 6023
rect 5293 6001 5449 6005
rect 5087 5986 5108 5989
rect 5051 5967 5108 5986
rect 5388 5985 5449 6001
rect 107 5861 164 5880
rect 107 5858 128 5861
rect 13 5843 128 5858
rect 146 5843 164 5861
rect 13 5820 164 5843
rect 13 5784 55 5820
rect 10328 6043 10484 6064
rect 10384 6042 10484 6043
rect 10673 6073 10773 6074
rect 10673 6052 10829 6073
rect 15705 6195 15723 6213
rect 15741 6198 15856 6213
rect 16051 6207 16112 6223
rect 15741 6195 15762 6198
rect 15705 6176 15762 6195
rect 20982 6252 21138 6273
rect 21038 6251 21138 6252
rect 21095 6215 21137 6251
rect 20986 6192 21137 6215
rect 15708 6115 15769 6131
rect 16049 6130 16106 6149
rect 16049 6127 16070 6130
rect 15708 6111 15864 6115
rect 15708 6093 15728 6111
rect 15746 6093 15864 6111
rect 12 5783 112 5784
rect 12 5762 168 5783
rect 10441 6006 10483 6042
rect 10673 6034 10791 6052
rect 10809 6034 10829 6052
rect 10673 6030 10829 6034
rect 10768 6014 10829 6030
rect 10332 5983 10483 6006
rect 15708 6072 15864 6093
rect 15764 6071 15864 6072
rect 15955 6112 16070 6127
rect 16088 6112 16106 6130
rect 15955 6089 16106 6112
rect 10332 5965 10350 5983
rect 10368 5968 10483 5983
rect 10368 5965 10389 5968
rect 10332 5946 10389 5965
rect 5047 5825 5108 5841
rect 5388 5840 5445 5859
rect 5388 5837 5409 5840
rect 5047 5821 5203 5825
rect 5047 5803 5067 5821
rect 5085 5803 5203 5821
rect 12 5744 130 5762
rect 148 5744 168 5762
rect 12 5740 168 5744
rect 107 5724 168 5740
rect 114 5660 171 5679
rect 114 5657 135 5660
rect 20 5642 135 5657
rect 153 5642 171 5660
rect 5047 5782 5203 5803
rect 5103 5781 5203 5782
rect 5294 5822 5409 5837
rect 5427 5822 5445 5840
rect 5294 5799 5445 5822
rect 5160 5745 5202 5781
rect 5294 5763 5336 5799
rect 15821 6035 15863 6071
rect 15955 6053 15997 6089
rect 15712 6012 15863 6035
rect 15712 5994 15730 6012
rect 15748 5997 15863 6012
rect 15954 6052 16054 6053
rect 15954 6031 16110 6052
rect 20986 6174 21004 6192
rect 21022 6177 21137 6192
rect 21022 6174 21043 6177
rect 20986 6155 21043 6174
rect 20989 6094 21050 6110
rect 20989 6090 21145 6094
rect 20989 6072 21009 6090
rect 21027 6072 21145 6090
rect 15954 6013 16072 6031
rect 16090 6013 16110 6031
rect 15954 6009 16110 6013
rect 15748 5994 15769 5997
rect 15712 5975 15769 5994
rect 16049 5993 16110 6009
rect 10768 5869 10825 5888
rect 10768 5866 10789 5869
rect 10674 5851 10789 5866
rect 10807 5851 10825 5869
rect 5051 5722 5202 5745
rect 5051 5704 5069 5722
rect 5087 5707 5202 5722
rect 5293 5762 5393 5763
rect 5293 5741 5449 5762
rect 10674 5828 10825 5851
rect 10328 5804 10389 5820
rect 10328 5800 10484 5804
rect 10328 5782 10348 5800
rect 10366 5782 10484 5800
rect 10674 5792 10716 5828
rect 20989 6051 21145 6072
rect 21045 6050 21145 6051
rect 5293 5723 5411 5741
rect 5429 5723 5449 5741
rect 5293 5719 5449 5723
rect 5087 5704 5108 5707
rect 5051 5685 5108 5704
rect 5388 5703 5449 5719
rect 20 5619 171 5642
rect 20 5583 62 5619
rect 19 5582 119 5583
rect 19 5561 175 5582
rect 5395 5639 5452 5658
rect 5395 5636 5416 5639
rect 19 5543 137 5561
rect 155 5543 175 5561
rect 19 5539 175 5543
rect 114 5523 175 5539
rect 5045 5611 5106 5627
rect 5301 5621 5416 5636
rect 5434 5621 5452 5639
rect 10328 5761 10484 5782
rect 10384 5760 10484 5761
rect 10673 5791 10773 5792
rect 10673 5770 10829 5791
rect 21102 6014 21144 6050
rect 20993 5991 21144 6014
rect 20993 5973 21011 5991
rect 21029 5976 21144 5991
rect 21029 5973 21050 5976
rect 20993 5954 21050 5973
rect 15708 5833 15769 5849
rect 16049 5848 16106 5867
rect 16049 5845 16070 5848
rect 15708 5829 15864 5833
rect 15708 5811 15728 5829
rect 15746 5811 15864 5829
rect 10441 5724 10483 5760
rect 10673 5752 10791 5770
rect 10809 5752 10829 5770
rect 10673 5748 10829 5752
rect 10768 5732 10829 5748
rect 10332 5701 10483 5724
rect 10332 5683 10350 5701
rect 10368 5686 10483 5701
rect 10368 5683 10389 5686
rect 10332 5664 10389 5683
rect 10775 5668 10832 5687
rect 10775 5665 10796 5668
rect 10681 5650 10796 5665
rect 10814 5650 10832 5668
rect 15708 5790 15864 5811
rect 15764 5789 15864 5790
rect 15955 5830 16070 5845
rect 16088 5830 16106 5848
rect 15955 5807 16106 5830
rect 15821 5753 15863 5789
rect 15955 5771 15997 5807
rect 15712 5730 15863 5753
rect 15712 5712 15730 5730
rect 15748 5715 15863 5730
rect 15954 5770 16054 5771
rect 15954 5749 16110 5770
rect 20989 5812 21050 5828
rect 20989 5808 21145 5812
rect 20989 5790 21009 5808
rect 21027 5790 21145 5808
rect 15954 5731 16072 5749
rect 16090 5731 16110 5749
rect 15954 5727 16110 5731
rect 15748 5712 15769 5715
rect 15712 5693 15769 5712
rect 16049 5711 16110 5727
rect 5045 5607 5201 5611
rect 5045 5589 5065 5607
rect 5083 5589 5201 5607
rect 5045 5568 5201 5589
rect 5101 5567 5201 5568
rect 5301 5598 5452 5621
rect 5158 5531 5200 5567
rect 5301 5562 5343 5598
rect 5049 5508 5200 5531
rect 5300 5561 5400 5562
rect 5300 5540 5456 5561
rect 10681 5627 10832 5650
rect 5300 5522 5418 5540
rect 5436 5522 5456 5540
rect 5300 5518 5456 5522
rect 5049 5490 5067 5508
rect 5085 5493 5200 5508
rect 5395 5502 5456 5518
rect 10326 5590 10387 5606
rect 10681 5591 10723 5627
rect 10680 5590 10780 5591
rect 10326 5586 10482 5590
rect 10326 5568 10346 5586
rect 10364 5568 10482 5586
rect 10326 5547 10482 5568
rect 10680 5569 10836 5590
rect 16056 5647 16113 5666
rect 16056 5644 16077 5647
rect 10680 5551 10798 5569
rect 10816 5551 10836 5569
rect 10680 5547 10836 5551
rect 10382 5546 10482 5547
rect 5085 5490 5106 5493
rect 5049 5471 5106 5490
rect 10439 5510 10481 5546
rect 10775 5531 10836 5547
rect 15706 5619 15767 5635
rect 15962 5629 16077 5644
rect 16095 5629 16113 5647
rect 20989 5769 21145 5790
rect 21045 5768 21145 5769
rect 21102 5732 21144 5768
rect 20993 5709 21144 5732
rect 20993 5691 21011 5709
rect 21029 5694 21144 5709
rect 21029 5691 21050 5694
rect 20993 5672 21050 5691
rect 15706 5615 15862 5619
rect 15706 5597 15726 5615
rect 15744 5597 15862 5615
rect 15706 5576 15862 5597
rect 15762 5575 15862 5576
rect 15962 5606 16113 5629
rect 10330 5487 10481 5510
rect 10330 5469 10348 5487
rect 10366 5472 10481 5487
rect 10366 5469 10387 5472
rect 10330 5450 10387 5469
rect 15819 5539 15861 5575
rect 15962 5570 16004 5606
rect 15710 5516 15861 5539
rect 15961 5569 16061 5570
rect 15961 5548 16117 5569
rect 15961 5530 16079 5548
rect 16097 5530 16117 5548
rect 15961 5526 16117 5530
rect 15710 5498 15728 5516
rect 15746 5501 15861 5516
rect 16056 5510 16117 5526
rect 20987 5598 21048 5614
rect 20987 5594 21143 5598
rect 20987 5576 21007 5594
rect 21025 5576 21143 5594
rect 20987 5555 21143 5576
rect 21043 5554 21143 5555
rect 15746 5498 15767 5501
rect 15710 5479 15767 5498
rect 21100 5518 21142 5554
rect 20991 5495 21142 5518
rect 20991 5477 21009 5495
rect 21027 5480 21142 5495
rect 21027 5477 21048 5480
rect 20991 5458 21048 5477
rect 114 5376 171 5395
rect 114 5373 135 5376
rect 20 5358 135 5373
rect 153 5358 171 5376
rect 20 5335 171 5358
rect 20 5299 62 5335
rect 5395 5355 5452 5374
rect 5395 5352 5416 5355
rect 19 5298 119 5299
rect 19 5277 175 5298
rect 19 5259 137 5277
rect 155 5259 175 5277
rect 19 5255 175 5259
rect 114 5239 175 5255
rect 5045 5327 5106 5343
rect 5301 5337 5416 5352
rect 5434 5337 5452 5355
rect 5045 5323 5201 5327
rect 5045 5305 5065 5323
rect 5083 5305 5201 5323
rect 5045 5284 5201 5305
rect 5101 5283 5201 5284
rect 5301 5314 5452 5337
rect 5158 5247 5200 5283
rect 5301 5278 5343 5314
rect 10775 5384 10832 5403
rect 10775 5381 10796 5384
rect 10681 5366 10796 5381
rect 10814 5366 10832 5384
rect 10681 5343 10832 5366
rect 5049 5224 5200 5247
rect 5300 5277 5400 5278
rect 5300 5256 5456 5277
rect 5300 5238 5418 5256
rect 5436 5238 5456 5256
rect 5300 5234 5456 5238
rect 112 5162 169 5181
rect 112 5159 133 5162
rect 18 5144 133 5159
rect 151 5144 169 5162
rect 18 5121 169 5144
rect 18 5085 60 5121
rect 17 5084 117 5085
rect 17 5063 173 5084
rect 5049 5206 5067 5224
rect 5085 5209 5200 5224
rect 5395 5218 5456 5234
rect 10326 5306 10387 5322
rect 10681 5307 10723 5343
rect 16056 5363 16113 5382
rect 16056 5360 16077 5363
rect 10680 5306 10780 5307
rect 10326 5302 10482 5306
rect 10326 5284 10346 5302
rect 10364 5284 10482 5302
rect 5085 5206 5106 5209
rect 5049 5187 5106 5206
rect 10326 5263 10482 5284
rect 10680 5285 10836 5306
rect 10680 5267 10798 5285
rect 10816 5267 10836 5285
rect 10680 5263 10836 5267
rect 10382 5262 10482 5263
rect 10439 5226 10481 5262
rect 10775 5247 10836 5263
rect 15706 5335 15767 5351
rect 15962 5345 16077 5360
rect 16095 5345 16113 5363
rect 15706 5331 15862 5335
rect 15706 5313 15726 5331
rect 15744 5313 15862 5331
rect 10330 5203 10481 5226
rect 15706 5292 15862 5313
rect 15762 5291 15862 5292
rect 15962 5322 16113 5345
rect 15819 5255 15861 5291
rect 15962 5286 16004 5322
rect 15710 5232 15861 5255
rect 15961 5285 16061 5286
rect 15961 5264 16117 5285
rect 15961 5246 16079 5264
rect 16097 5246 16117 5264
rect 15961 5242 16117 5246
rect 5052 5126 5113 5142
rect 5393 5141 5450 5160
rect 5393 5138 5414 5141
rect 5052 5122 5208 5126
rect 5052 5104 5072 5122
rect 5090 5104 5208 5122
rect 17 5045 135 5063
rect 153 5045 173 5063
rect 17 5041 173 5045
rect 112 5025 173 5041
rect 5052 5083 5208 5104
rect 5108 5082 5208 5083
rect 5299 5123 5414 5138
rect 5432 5123 5450 5141
rect 5299 5100 5450 5123
rect 5165 5046 5207 5082
rect 5299 5064 5341 5100
rect 5056 5023 5207 5046
rect 5056 5005 5074 5023
rect 5092 5008 5207 5023
rect 5298 5063 5398 5064
rect 5298 5042 5454 5063
rect 10330 5185 10348 5203
rect 10366 5188 10481 5203
rect 10366 5185 10387 5188
rect 10330 5166 10387 5185
rect 10773 5170 10830 5189
rect 10773 5167 10794 5170
rect 10679 5152 10794 5167
rect 10812 5152 10830 5170
rect 10679 5129 10830 5152
rect 10333 5105 10394 5121
rect 10333 5101 10489 5105
rect 10333 5083 10353 5101
rect 10371 5083 10489 5101
rect 10679 5093 10721 5129
rect 5298 5024 5416 5042
rect 5434 5024 5454 5042
rect 5298 5020 5454 5024
rect 5092 5005 5113 5008
rect 5056 4986 5113 5005
rect 5393 5004 5454 5020
rect 112 4880 169 4899
rect 112 4877 133 4880
rect 18 4862 133 4877
rect 151 4862 169 4880
rect 18 4839 169 4862
rect 18 4803 60 4839
rect 10333 5062 10489 5083
rect 10389 5061 10489 5062
rect 10678 5092 10778 5093
rect 10678 5071 10834 5092
rect 15710 5214 15728 5232
rect 15746 5217 15861 5232
rect 16056 5226 16117 5242
rect 20987 5314 21048 5330
rect 20987 5310 21143 5314
rect 20987 5292 21007 5310
rect 21025 5292 21143 5310
rect 15746 5214 15767 5217
rect 15710 5195 15767 5214
rect 20987 5271 21143 5292
rect 21043 5270 21143 5271
rect 21100 5234 21142 5270
rect 20991 5211 21142 5234
rect 15713 5134 15774 5150
rect 16054 5149 16111 5168
rect 16054 5146 16075 5149
rect 15713 5130 15869 5134
rect 15713 5112 15733 5130
rect 15751 5112 15869 5130
rect 17 4802 117 4803
rect 17 4781 173 4802
rect 10446 5025 10488 5061
rect 10678 5053 10796 5071
rect 10814 5053 10834 5071
rect 10678 5049 10834 5053
rect 10773 5033 10834 5049
rect 10337 5002 10488 5025
rect 15713 5091 15869 5112
rect 15769 5090 15869 5091
rect 15960 5131 16075 5146
rect 16093 5131 16111 5149
rect 15960 5108 16111 5131
rect 10337 4984 10355 5002
rect 10373 4987 10488 5002
rect 10373 4984 10394 4987
rect 10337 4965 10394 4984
rect 5052 4844 5113 4860
rect 5393 4859 5450 4878
rect 5393 4856 5414 4859
rect 5052 4840 5208 4844
rect 5052 4822 5072 4840
rect 5090 4822 5208 4840
rect 17 4763 135 4781
rect 153 4763 173 4781
rect 17 4759 173 4763
rect 112 4743 173 4759
rect 119 4679 176 4698
rect 119 4676 140 4679
rect 25 4661 140 4676
rect 158 4661 176 4679
rect 5052 4801 5208 4822
rect 5108 4800 5208 4801
rect 5299 4841 5414 4856
rect 5432 4841 5450 4859
rect 5299 4818 5450 4841
rect 5165 4764 5207 4800
rect 5299 4782 5341 4818
rect 15826 5054 15868 5090
rect 15960 5072 16002 5108
rect 15717 5031 15868 5054
rect 15717 5013 15735 5031
rect 15753 5016 15868 5031
rect 15959 5071 16059 5072
rect 15959 5050 16115 5071
rect 20991 5193 21009 5211
rect 21027 5196 21142 5211
rect 21027 5193 21048 5196
rect 20991 5174 21048 5193
rect 20994 5113 21055 5129
rect 20994 5109 21150 5113
rect 20994 5091 21014 5109
rect 21032 5091 21150 5109
rect 15959 5032 16077 5050
rect 16095 5032 16115 5050
rect 15959 5028 16115 5032
rect 15753 5013 15774 5016
rect 15717 4994 15774 5013
rect 16054 5012 16115 5028
rect 10773 4888 10830 4907
rect 10773 4885 10794 4888
rect 10679 4870 10794 4885
rect 10812 4870 10830 4888
rect 5056 4741 5207 4764
rect 5056 4723 5074 4741
rect 5092 4726 5207 4741
rect 5298 4781 5398 4782
rect 5298 4760 5454 4781
rect 10679 4847 10830 4870
rect 10333 4823 10394 4839
rect 10333 4819 10489 4823
rect 10333 4801 10353 4819
rect 10371 4801 10489 4819
rect 10679 4811 10721 4847
rect 20994 5070 21150 5091
rect 21050 5069 21150 5070
rect 5298 4742 5416 4760
rect 5434 4742 5454 4760
rect 5298 4738 5454 4742
rect 5092 4723 5113 4726
rect 5056 4704 5113 4723
rect 5393 4722 5454 4738
rect 25 4638 176 4661
rect 25 4602 67 4638
rect 24 4601 124 4602
rect 24 4580 180 4601
rect 5400 4658 5457 4677
rect 5400 4655 5421 4658
rect 5050 4630 5111 4646
rect 5306 4640 5421 4655
rect 5439 4640 5457 4658
rect 10333 4780 10489 4801
rect 10389 4779 10489 4780
rect 10678 4810 10778 4811
rect 10678 4789 10834 4810
rect 21107 5033 21149 5069
rect 20998 5010 21149 5033
rect 20998 4992 21016 5010
rect 21034 4995 21149 5010
rect 21034 4992 21055 4995
rect 20998 4973 21055 4992
rect 15713 4852 15774 4868
rect 16054 4867 16111 4886
rect 16054 4864 16075 4867
rect 15713 4848 15869 4852
rect 15713 4830 15733 4848
rect 15751 4830 15869 4848
rect 10446 4743 10488 4779
rect 10678 4771 10796 4789
rect 10814 4771 10834 4789
rect 10678 4767 10834 4771
rect 10773 4751 10834 4767
rect 10337 4720 10488 4743
rect 10337 4702 10355 4720
rect 10373 4705 10488 4720
rect 10373 4702 10394 4705
rect 10337 4683 10394 4702
rect 10780 4687 10837 4706
rect 10780 4684 10801 4687
rect 10686 4669 10801 4684
rect 10819 4669 10837 4687
rect 15713 4809 15869 4830
rect 15769 4808 15869 4809
rect 15960 4849 16075 4864
rect 16093 4849 16111 4867
rect 15960 4826 16111 4849
rect 15826 4772 15868 4808
rect 15960 4790 16002 4826
rect 15717 4749 15868 4772
rect 15717 4731 15735 4749
rect 15753 4734 15868 4749
rect 15959 4789 16059 4790
rect 15959 4768 16115 4789
rect 20994 4831 21055 4847
rect 20994 4827 21150 4831
rect 20994 4809 21014 4827
rect 21032 4809 21150 4827
rect 15959 4750 16077 4768
rect 16095 4750 16115 4768
rect 15959 4746 16115 4750
rect 15753 4731 15774 4734
rect 15717 4712 15774 4731
rect 16054 4730 16115 4746
rect 24 4562 142 4580
rect 160 4562 180 4580
rect 24 4558 180 4562
rect 119 4542 180 4558
rect 5050 4626 5206 4630
rect 5050 4608 5070 4626
rect 5088 4608 5206 4626
rect 5050 4587 5206 4608
rect 5106 4586 5206 4587
rect 5306 4617 5457 4640
rect 117 4400 174 4419
rect 117 4397 138 4400
rect 23 4382 138 4397
rect 156 4382 174 4400
rect 23 4359 174 4382
rect 23 4323 65 4359
rect 5163 4550 5205 4586
rect 5306 4581 5348 4617
rect 5054 4527 5205 4550
rect 5305 4580 5405 4581
rect 5305 4559 5461 4580
rect 10686 4646 10837 4669
rect 10331 4609 10392 4625
rect 10686 4610 10728 4646
rect 10685 4609 10785 4610
rect 5305 4541 5423 4559
rect 5441 4541 5461 4559
rect 5305 4537 5461 4541
rect 5054 4509 5072 4527
rect 5090 4512 5205 4527
rect 5400 4521 5461 4537
rect 10331 4605 10487 4609
rect 10331 4587 10351 4605
rect 10369 4587 10487 4605
rect 10331 4566 10487 4587
rect 10685 4588 10841 4609
rect 16061 4666 16118 4685
rect 16061 4663 16082 4666
rect 15711 4638 15772 4654
rect 15967 4648 16082 4663
rect 16100 4648 16118 4666
rect 20994 4788 21150 4809
rect 21050 4787 21150 4788
rect 21107 4751 21149 4787
rect 20998 4728 21149 4751
rect 20998 4710 21016 4728
rect 21034 4713 21149 4728
rect 21034 4710 21055 4713
rect 20998 4691 21055 4710
rect 10685 4570 10803 4588
rect 10821 4570 10841 4588
rect 10685 4566 10841 4570
rect 10387 4565 10487 4566
rect 5090 4509 5111 4512
rect 5054 4490 5111 4509
rect 5398 4379 5455 4398
rect 5398 4376 5419 4379
rect 22 4322 122 4323
rect 22 4301 178 4322
rect 22 4283 140 4301
rect 158 4283 178 4301
rect 22 4279 178 4283
rect 5048 4351 5109 4367
rect 5304 4361 5419 4376
rect 5437 4361 5455 4379
rect 5048 4347 5204 4351
rect 5048 4329 5068 4347
rect 5086 4329 5204 4347
rect 117 4263 178 4279
rect 5048 4308 5204 4329
rect 5104 4307 5204 4308
rect 5304 4338 5455 4361
rect 5161 4271 5203 4307
rect 5304 4302 5346 4338
rect 10444 4529 10486 4565
rect 10780 4550 10841 4566
rect 15711 4634 15867 4638
rect 15711 4616 15731 4634
rect 15749 4616 15867 4634
rect 15711 4595 15867 4616
rect 15767 4594 15867 4595
rect 15967 4625 16118 4648
rect 10335 4506 10486 4529
rect 10335 4488 10353 4506
rect 10371 4491 10486 4506
rect 10371 4488 10392 4491
rect 10335 4469 10392 4488
rect 10778 4408 10835 4427
rect 10778 4405 10799 4408
rect 10684 4390 10799 4405
rect 10817 4390 10835 4408
rect 10684 4367 10835 4390
rect 5052 4248 5203 4271
rect 5303 4301 5403 4302
rect 5303 4280 5459 4301
rect 5303 4262 5421 4280
rect 5439 4262 5459 4280
rect 5303 4258 5459 4262
rect 10329 4330 10390 4346
rect 10684 4331 10726 4367
rect 15824 4558 15866 4594
rect 15967 4589 16009 4625
rect 15715 4535 15866 4558
rect 15966 4588 16066 4589
rect 15966 4567 16122 4588
rect 20992 4617 21053 4633
rect 15966 4549 16084 4567
rect 16102 4549 16122 4567
rect 15966 4545 16122 4549
rect 15715 4517 15733 4535
rect 15751 4520 15866 4535
rect 16061 4529 16122 4545
rect 20992 4613 21148 4617
rect 20992 4595 21012 4613
rect 21030 4595 21148 4613
rect 20992 4574 21148 4595
rect 21048 4573 21148 4574
rect 15751 4517 15772 4520
rect 15715 4498 15772 4517
rect 16059 4387 16116 4406
rect 16059 4384 16080 4387
rect 10683 4330 10783 4331
rect 10329 4326 10485 4330
rect 10329 4308 10349 4326
rect 10367 4308 10485 4326
rect 115 4186 172 4205
rect 115 4183 136 4186
rect 21 4168 136 4183
rect 154 4168 172 4186
rect 21 4145 172 4168
rect 21 4109 63 4145
rect 20 4108 120 4109
rect 20 4087 176 4108
rect 5052 4230 5070 4248
rect 5088 4233 5203 4248
rect 5398 4242 5459 4258
rect 5088 4230 5109 4233
rect 5052 4211 5109 4230
rect 10329 4287 10485 4308
rect 10683 4309 10839 4330
rect 10683 4291 10801 4309
rect 10819 4291 10839 4309
rect 10683 4287 10839 4291
rect 15709 4359 15770 4375
rect 15965 4369 16080 4384
rect 16098 4369 16116 4387
rect 15709 4355 15865 4359
rect 15709 4337 15729 4355
rect 15747 4337 15865 4355
rect 10385 4286 10485 4287
rect 10442 4250 10484 4286
rect 10778 4271 10839 4287
rect 10333 4227 10484 4250
rect 15709 4316 15865 4337
rect 15765 4315 15865 4316
rect 15965 4346 16116 4369
rect 15822 4279 15864 4315
rect 15965 4310 16007 4346
rect 21105 4537 21147 4573
rect 20996 4514 21147 4537
rect 20996 4496 21014 4514
rect 21032 4499 21147 4514
rect 21032 4496 21053 4499
rect 20996 4477 21053 4496
rect 15713 4256 15864 4279
rect 15964 4309 16064 4310
rect 15964 4288 16120 4309
rect 15964 4270 16082 4288
rect 16100 4270 16120 4288
rect 15964 4266 16120 4270
rect 20990 4338 21051 4354
rect 20990 4334 21146 4338
rect 20990 4316 21010 4334
rect 21028 4316 21146 4334
rect 5055 4150 5116 4166
rect 5396 4165 5453 4184
rect 5396 4162 5417 4165
rect 5055 4146 5211 4150
rect 5055 4128 5075 4146
rect 5093 4128 5211 4146
rect 20 4069 138 4087
rect 156 4069 176 4087
rect 20 4065 176 4069
rect 115 4049 176 4065
rect 5055 4107 5211 4128
rect 5111 4106 5211 4107
rect 5302 4147 5417 4162
rect 5435 4147 5453 4165
rect 5302 4124 5453 4147
rect 5168 4070 5210 4106
rect 5302 4088 5344 4124
rect 5059 4047 5210 4070
rect 5059 4029 5077 4047
rect 5095 4032 5210 4047
rect 5301 4087 5401 4088
rect 5301 4066 5457 4087
rect 10333 4209 10351 4227
rect 10369 4212 10484 4227
rect 10369 4209 10390 4212
rect 10333 4190 10390 4209
rect 10776 4194 10833 4213
rect 10776 4191 10797 4194
rect 10682 4176 10797 4191
rect 10815 4176 10833 4194
rect 10682 4153 10833 4176
rect 10336 4129 10397 4145
rect 10336 4125 10492 4129
rect 10336 4107 10356 4125
rect 10374 4107 10492 4125
rect 10682 4117 10724 4153
rect 5301 4048 5419 4066
rect 5437 4048 5457 4066
rect 5301 4044 5457 4048
rect 5095 4029 5116 4032
rect 5059 4010 5116 4029
rect 5396 4028 5457 4044
rect 115 3904 172 3923
rect 115 3901 136 3904
rect 21 3886 136 3901
rect 154 3886 172 3904
rect 21 3863 172 3886
rect 21 3827 63 3863
rect 10336 4086 10492 4107
rect 10392 4085 10492 4086
rect 10681 4116 10781 4117
rect 10681 4095 10837 4116
rect 15713 4238 15731 4256
rect 15749 4241 15864 4256
rect 16059 4250 16120 4266
rect 15749 4238 15770 4241
rect 15713 4219 15770 4238
rect 20990 4295 21146 4316
rect 21046 4294 21146 4295
rect 21103 4258 21145 4294
rect 20994 4235 21145 4258
rect 15716 4158 15777 4174
rect 16057 4173 16114 4192
rect 16057 4170 16078 4173
rect 15716 4154 15872 4158
rect 15716 4136 15736 4154
rect 15754 4136 15872 4154
rect 20 3826 120 3827
rect 20 3805 176 3826
rect 10449 4049 10491 4085
rect 10681 4077 10799 4095
rect 10817 4077 10837 4095
rect 10681 4073 10837 4077
rect 10776 4057 10837 4073
rect 10340 4026 10491 4049
rect 15716 4115 15872 4136
rect 15772 4114 15872 4115
rect 15963 4155 16078 4170
rect 16096 4155 16114 4173
rect 15963 4132 16114 4155
rect 10340 4008 10358 4026
rect 10376 4011 10491 4026
rect 10376 4008 10397 4011
rect 10340 3989 10397 4008
rect 5055 3868 5116 3884
rect 5396 3883 5453 3902
rect 5396 3880 5417 3883
rect 5055 3864 5211 3868
rect 5055 3846 5075 3864
rect 5093 3846 5211 3864
rect 20 3787 138 3805
rect 156 3787 176 3805
rect 20 3783 176 3787
rect 115 3767 176 3783
rect 122 3703 179 3722
rect 122 3700 143 3703
rect 28 3685 143 3700
rect 161 3685 179 3703
rect 5055 3825 5211 3846
rect 5111 3824 5211 3825
rect 5302 3865 5417 3880
rect 5435 3865 5453 3883
rect 5302 3842 5453 3865
rect 5168 3788 5210 3824
rect 5302 3806 5344 3842
rect 15829 4078 15871 4114
rect 15963 4096 16005 4132
rect 15720 4055 15871 4078
rect 15720 4037 15738 4055
rect 15756 4040 15871 4055
rect 15962 4095 16062 4096
rect 15962 4074 16118 4095
rect 20994 4217 21012 4235
rect 21030 4220 21145 4235
rect 21030 4217 21051 4220
rect 20994 4198 21051 4217
rect 20997 4137 21058 4153
rect 20997 4133 21153 4137
rect 20997 4115 21017 4133
rect 21035 4115 21153 4133
rect 15962 4056 16080 4074
rect 16098 4056 16118 4074
rect 15962 4052 16118 4056
rect 15756 4037 15777 4040
rect 15720 4018 15777 4037
rect 16057 4036 16118 4052
rect 10776 3912 10833 3931
rect 10776 3909 10797 3912
rect 10682 3894 10797 3909
rect 10815 3894 10833 3912
rect 5059 3765 5210 3788
rect 5059 3747 5077 3765
rect 5095 3750 5210 3765
rect 5301 3805 5401 3806
rect 5301 3784 5457 3805
rect 10682 3871 10833 3894
rect 10336 3847 10397 3863
rect 10336 3843 10492 3847
rect 10336 3825 10356 3843
rect 10374 3825 10492 3843
rect 10682 3835 10724 3871
rect 20997 4094 21153 4115
rect 21053 4093 21153 4094
rect 5301 3766 5419 3784
rect 5437 3766 5457 3784
rect 5301 3762 5457 3766
rect 5095 3747 5116 3750
rect 5059 3728 5116 3747
rect 5396 3746 5457 3762
rect 28 3662 179 3685
rect 28 3626 70 3662
rect 27 3625 127 3626
rect 27 3604 183 3625
rect 5403 3682 5460 3701
rect 5403 3679 5424 3682
rect 27 3586 145 3604
rect 163 3586 183 3604
rect 27 3582 183 3586
rect 122 3566 183 3582
rect 5053 3654 5114 3670
rect 5309 3664 5424 3679
rect 5442 3664 5460 3682
rect 10336 3804 10492 3825
rect 10392 3803 10492 3804
rect 10681 3834 10781 3835
rect 10681 3813 10837 3834
rect 21110 4057 21152 4093
rect 21001 4034 21152 4057
rect 21001 4016 21019 4034
rect 21037 4019 21152 4034
rect 21037 4016 21058 4019
rect 21001 3997 21058 4016
rect 15716 3876 15777 3892
rect 16057 3891 16114 3910
rect 16057 3888 16078 3891
rect 15716 3872 15872 3876
rect 15716 3854 15736 3872
rect 15754 3854 15872 3872
rect 10449 3767 10491 3803
rect 10681 3795 10799 3813
rect 10817 3795 10837 3813
rect 10681 3791 10837 3795
rect 10776 3775 10837 3791
rect 10340 3744 10491 3767
rect 10340 3726 10358 3744
rect 10376 3729 10491 3744
rect 10376 3726 10397 3729
rect 10340 3707 10397 3726
rect 10783 3711 10840 3730
rect 10783 3708 10804 3711
rect 10689 3693 10804 3708
rect 10822 3693 10840 3711
rect 15716 3833 15872 3854
rect 15772 3832 15872 3833
rect 15963 3873 16078 3888
rect 16096 3873 16114 3891
rect 15963 3850 16114 3873
rect 15829 3796 15871 3832
rect 15963 3814 16005 3850
rect 15720 3773 15871 3796
rect 15720 3755 15738 3773
rect 15756 3758 15871 3773
rect 15962 3813 16062 3814
rect 15962 3792 16118 3813
rect 20997 3855 21058 3871
rect 20997 3851 21153 3855
rect 20997 3833 21017 3851
rect 21035 3833 21153 3851
rect 15962 3774 16080 3792
rect 16098 3774 16118 3792
rect 15962 3770 16118 3774
rect 15756 3755 15777 3758
rect 15720 3736 15777 3755
rect 16057 3754 16118 3770
rect 5053 3650 5209 3654
rect 5053 3632 5073 3650
rect 5091 3632 5209 3650
rect 5053 3611 5209 3632
rect 5109 3610 5209 3611
rect 5309 3641 5460 3664
rect 5166 3574 5208 3610
rect 5309 3605 5351 3641
rect 5057 3551 5208 3574
rect 5308 3604 5408 3605
rect 5308 3583 5464 3604
rect 10689 3670 10840 3693
rect 5308 3565 5426 3583
rect 5444 3565 5464 3583
rect 5308 3561 5464 3565
rect 5057 3533 5075 3551
rect 5093 3536 5208 3551
rect 5403 3545 5464 3561
rect 10334 3633 10395 3649
rect 10689 3634 10731 3670
rect 10688 3633 10788 3634
rect 10334 3629 10490 3633
rect 10334 3611 10354 3629
rect 10372 3611 10490 3629
rect 10334 3590 10490 3611
rect 10688 3612 10844 3633
rect 16064 3690 16121 3709
rect 16064 3687 16085 3690
rect 10688 3594 10806 3612
rect 10824 3594 10844 3612
rect 10688 3590 10844 3594
rect 10390 3589 10490 3590
rect 5093 3533 5114 3536
rect 5057 3514 5114 3533
rect 10447 3553 10489 3589
rect 10783 3574 10844 3590
rect 15714 3662 15775 3678
rect 15970 3672 16085 3687
rect 16103 3672 16121 3690
rect 20997 3812 21153 3833
rect 21053 3811 21153 3812
rect 21110 3775 21152 3811
rect 21001 3752 21152 3775
rect 21001 3734 21019 3752
rect 21037 3737 21152 3752
rect 21037 3734 21058 3737
rect 21001 3715 21058 3734
rect 15714 3658 15870 3662
rect 15714 3640 15734 3658
rect 15752 3640 15870 3658
rect 15714 3619 15870 3640
rect 15770 3618 15870 3619
rect 15970 3649 16121 3672
rect 10338 3530 10489 3553
rect 10338 3512 10356 3530
rect 10374 3515 10489 3530
rect 10374 3512 10395 3515
rect 10338 3493 10395 3512
rect 15827 3582 15869 3618
rect 15970 3613 16012 3649
rect 15718 3559 15869 3582
rect 15969 3612 16069 3613
rect 15969 3591 16125 3612
rect 15969 3573 16087 3591
rect 16105 3573 16125 3591
rect 15969 3569 16125 3573
rect 15718 3541 15736 3559
rect 15754 3544 15869 3559
rect 16064 3553 16125 3569
rect 20995 3641 21056 3657
rect 20995 3637 21151 3641
rect 20995 3619 21015 3637
rect 21033 3619 21151 3637
rect 20995 3598 21151 3619
rect 21051 3597 21151 3598
rect 15754 3541 15775 3544
rect 15718 3522 15775 3541
rect 21108 3561 21150 3597
rect 20999 3538 21150 3561
rect 20999 3520 21017 3538
rect 21035 3523 21150 3538
rect 21035 3520 21056 3523
rect 20999 3501 21056 3520
rect 122 3419 179 3438
rect 122 3416 143 3419
rect 28 3401 143 3416
rect 161 3401 179 3419
rect 28 3378 179 3401
rect 28 3342 70 3378
rect 5403 3398 5460 3417
rect 5403 3395 5424 3398
rect 27 3341 127 3342
rect 27 3320 183 3341
rect 27 3302 145 3320
rect 163 3302 183 3320
rect 27 3298 183 3302
rect 122 3282 183 3298
rect 5053 3370 5114 3386
rect 5309 3380 5424 3395
rect 5442 3380 5460 3398
rect 5053 3366 5209 3370
rect 5053 3348 5073 3366
rect 5091 3348 5209 3366
rect 5053 3327 5209 3348
rect 5109 3326 5209 3327
rect 5309 3357 5460 3380
rect 5166 3290 5208 3326
rect 5309 3321 5351 3357
rect 10783 3427 10840 3446
rect 10783 3424 10804 3427
rect 10689 3409 10804 3424
rect 10822 3409 10840 3427
rect 10689 3386 10840 3409
rect 5057 3267 5208 3290
rect 5308 3320 5408 3321
rect 5308 3299 5464 3320
rect 5308 3281 5426 3299
rect 5444 3281 5464 3299
rect 5308 3277 5464 3281
rect 120 3205 177 3224
rect 120 3202 141 3205
rect 26 3187 141 3202
rect 159 3187 177 3205
rect 26 3164 177 3187
rect 26 3128 68 3164
rect 25 3127 125 3128
rect 25 3106 181 3127
rect 5057 3249 5075 3267
rect 5093 3252 5208 3267
rect 5403 3261 5464 3277
rect 10334 3349 10395 3365
rect 10689 3350 10731 3386
rect 16064 3406 16121 3425
rect 16064 3403 16085 3406
rect 10688 3349 10788 3350
rect 10334 3345 10490 3349
rect 10334 3327 10354 3345
rect 10372 3327 10490 3345
rect 5093 3249 5114 3252
rect 5057 3230 5114 3249
rect 10334 3306 10490 3327
rect 10688 3328 10844 3349
rect 10688 3310 10806 3328
rect 10824 3310 10844 3328
rect 10688 3306 10844 3310
rect 10390 3305 10490 3306
rect 10447 3269 10489 3305
rect 10783 3290 10844 3306
rect 15714 3378 15775 3394
rect 15970 3388 16085 3403
rect 16103 3388 16121 3406
rect 15714 3374 15870 3378
rect 15714 3356 15734 3374
rect 15752 3356 15870 3374
rect 10338 3246 10489 3269
rect 15714 3335 15870 3356
rect 15770 3334 15870 3335
rect 15970 3365 16121 3388
rect 15827 3298 15869 3334
rect 15970 3329 16012 3365
rect 15718 3275 15869 3298
rect 15969 3328 16069 3329
rect 15969 3307 16125 3328
rect 15969 3289 16087 3307
rect 16105 3289 16125 3307
rect 15969 3285 16125 3289
rect 5060 3169 5121 3185
rect 5401 3184 5458 3203
rect 5401 3181 5422 3184
rect 5060 3165 5216 3169
rect 5060 3147 5080 3165
rect 5098 3147 5216 3165
rect 25 3088 143 3106
rect 161 3088 181 3106
rect 25 3084 181 3088
rect 120 3068 181 3084
rect 5060 3126 5216 3147
rect 5116 3125 5216 3126
rect 5307 3166 5422 3181
rect 5440 3166 5458 3184
rect 5307 3143 5458 3166
rect 5173 3089 5215 3125
rect 5307 3107 5349 3143
rect 5064 3066 5215 3089
rect 5064 3048 5082 3066
rect 5100 3051 5215 3066
rect 5306 3106 5406 3107
rect 5306 3085 5462 3106
rect 10338 3228 10356 3246
rect 10374 3231 10489 3246
rect 10374 3228 10395 3231
rect 10338 3209 10395 3228
rect 10781 3213 10838 3232
rect 10781 3210 10802 3213
rect 10687 3195 10802 3210
rect 10820 3195 10838 3213
rect 10687 3172 10838 3195
rect 10341 3148 10402 3164
rect 10341 3144 10497 3148
rect 10341 3126 10361 3144
rect 10379 3126 10497 3144
rect 10687 3136 10729 3172
rect 5306 3067 5424 3085
rect 5442 3067 5462 3085
rect 5306 3063 5462 3067
rect 5100 3048 5121 3051
rect 5064 3029 5121 3048
rect 5401 3047 5462 3063
rect 120 2923 177 2942
rect 120 2920 141 2923
rect 26 2905 141 2920
rect 159 2905 177 2923
rect 26 2882 177 2905
rect 26 2846 68 2882
rect 10341 3105 10497 3126
rect 10397 3104 10497 3105
rect 10686 3135 10786 3136
rect 10686 3114 10842 3135
rect 15718 3257 15736 3275
rect 15754 3260 15869 3275
rect 16064 3269 16125 3285
rect 20995 3357 21056 3373
rect 20995 3353 21151 3357
rect 20995 3335 21015 3353
rect 21033 3335 21151 3353
rect 15754 3257 15775 3260
rect 15718 3238 15775 3257
rect 20995 3314 21151 3335
rect 21051 3313 21151 3314
rect 21108 3277 21150 3313
rect 20999 3254 21150 3277
rect 15721 3177 15782 3193
rect 16062 3192 16119 3211
rect 16062 3189 16083 3192
rect 15721 3173 15877 3177
rect 15721 3155 15741 3173
rect 15759 3155 15877 3173
rect 25 2845 125 2846
rect 25 2824 181 2845
rect 10454 3068 10496 3104
rect 10686 3096 10804 3114
rect 10822 3096 10842 3114
rect 10686 3092 10842 3096
rect 10781 3076 10842 3092
rect 10345 3045 10496 3068
rect 15721 3134 15877 3155
rect 15777 3133 15877 3134
rect 15968 3174 16083 3189
rect 16101 3174 16119 3192
rect 15968 3151 16119 3174
rect 10345 3027 10363 3045
rect 10381 3030 10496 3045
rect 10381 3027 10402 3030
rect 10345 3008 10402 3027
rect 5060 2887 5121 2903
rect 5401 2902 5458 2921
rect 5401 2899 5422 2902
rect 5060 2883 5216 2887
rect 5060 2865 5080 2883
rect 5098 2865 5216 2883
rect 25 2806 143 2824
rect 161 2806 181 2824
rect 25 2802 181 2806
rect 120 2786 181 2802
rect 127 2722 184 2741
rect 127 2719 148 2722
rect 33 2704 148 2719
rect 166 2704 184 2722
rect 5060 2844 5216 2865
rect 5116 2843 5216 2844
rect 5307 2884 5422 2899
rect 5440 2884 5458 2902
rect 5307 2861 5458 2884
rect 5173 2807 5215 2843
rect 5307 2825 5349 2861
rect 15834 3097 15876 3133
rect 15968 3115 16010 3151
rect 15725 3074 15876 3097
rect 15725 3056 15743 3074
rect 15761 3059 15876 3074
rect 15967 3114 16067 3115
rect 15967 3093 16123 3114
rect 20999 3236 21017 3254
rect 21035 3239 21150 3254
rect 21035 3236 21056 3239
rect 20999 3217 21056 3236
rect 21002 3156 21063 3172
rect 21002 3152 21158 3156
rect 21002 3134 21022 3152
rect 21040 3134 21158 3152
rect 15967 3075 16085 3093
rect 16103 3075 16123 3093
rect 15967 3071 16123 3075
rect 15761 3056 15782 3059
rect 15725 3037 15782 3056
rect 16062 3055 16123 3071
rect 10781 2931 10838 2950
rect 10781 2928 10802 2931
rect 10687 2913 10802 2928
rect 10820 2913 10838 2931
rect 5064 2784 5215 2807
rect 5064 2766 5082 2784
rect 5100 2769 5215 2784
rect 5306 2824 5406 2825
rect 5306 2803 5462 2824
rect 10687 2890 10838 2913
rect 10341 2866 10402 2882
rect 10341 2862 10497 2866
rect 10341 2844 10361 2862
rect 10379 2844 10497 2862
rect 10687 2854 10729 2890
rect 21002 3113 21158 3134
rect 21058 3112 21158 3113
rect 5306 2785 5424 2803
rect 5442 2785 5462 2803
rect 5306 2781 5462 2785
rect 5100 2766 5121 2769
rect 5064 2747 5121 2766
rect 5401 2765 5462 2781
rect 33 2681 184 2704
rect 33 2645 75 2681
rect 32 2644 132 2645
rect 32 2623 188 2644
rect 5408 2701 5465 2720
rect 5408 2698 5429 2701
rect 5058 2673 5119 2689
rect 5314 2683 5429 2698
rect 5447 2683 5465 2701
rect 10341 2823 10497 2844
rect 10397 2822 10497 2823
rect 10686 2853 10786 2854
rect 10686 2832 10842 2853
rect 21115 3076 21157 3112
rect 21006 3053 21157 3076
rect 21006 3035 21024 3053
rect 21042 3038 21157 3053
rect 21042 3035 21063 3038
rect 21006 3016 21063 3035
rect 15721 2895 15782 2911
rect 16062 2910 16119 2929
rect 16062 2907 16083 2910
rect 15721 2891 15877 2895
rect 15721 2873 15741 2891
rect 15759 2873 15877 2891
rect 10454 2786 10496 2822
rect 10686 2814 10804 2832
rect 10822 2814 10842 2832
rect 10686 2810 10842 2814
rect 10781 2794 10842 2810
rect 10345 2763 10496 2786
rect 10345 2745 10363 2763
rect 10381 2748 10496 2763
rect 10381 2745 10402 2748
rect 10345 2726 10402 2745
rect 10788 2730 10845 2749
rect 10788 2727 10809 2730
rect 10694 2712 10809 2727
rect 10827 2712 10845 2730
rect 15721 2852 15877 2873
rect 15777 2851 15877 2852
rect 15968 2892 16083 2907
rect 16101 2892 16119 2910
rect 15968 2869 16119 2892
rect 15834 2815 15876 2851
rect 15968 2833 16010 2869
rect 15725 2792 15876 2815
rect 15725 2774 15743 2792
rect 15761 2777 15876 2792
rect 15967 2832 16067 2833
rect 15967 2811 16123 2832
rect 21002 2874 21063 2890
rect 21002 2870 21158 2874
rect 21002 2852 21022 2870
rect 21040 2852 21158 2870
rect 15967 2793 16085 2811
rect 16103 2793 16123 2811
rect 15967 2789 16123 2793
rect 15761 2774 15782 2777
rect 15725 2755 15782 2774
rect 16062 2773 16123 2789
rect 10694 2689 10845 2712
rect 5058 2669 5214 2673
rect 5058 2651 5078 2669
rect 5096 2651 5214 2669
rect 32 2605 150 2623
rect 168 2605 188 2623
rect 32 2601 188 2605
rect 127 2585 188 2601
rect 5058 2630 5214 2651
rect 5114 2629 5214 2630
rect 5314 2660 5465 2683
rect 5171 2593 5213 2629
rect 5314 2624 5356 2660
rect 5062 2570 5213 2593
rect 5313 2623 5413 2624
rect 5313 2602 5469 2623
rect 10339 2652 10400 2668
rect 10694 2653 10736 2689
rect 10693 2652 10793 2653
rect 10339 2648 10495 2652
rect 10339 2630 10359 2648
rect 10377 2630 10495 2648
rect 5313 2584 5431 2602
rect 5449 2584 5469 2602
rect 5313 2580 5469 2584
rect 129 2440 186 2459
rect 129 2437 150 2440
rect 35 2422 150 2437
rect 168 2422 186 2440
rect 5062 2552 5080 2570
rect 5098 2555 5213 2570
rect 5408 2564 5469 2580
rect 5098 2552 5119 2555
rect 5062 2533 5119 2552
rect 10339 2609 10495 2630
rect 10693 2631 10849 2652
rect 16069 2709 16126 2728
rect 16069 2706 16090 2709
rect 15719 2681 15780 2697
rect 15975 2691 16090 2706
rect 16108 2691 16126 2709
rect 21002 2831 21158 2852
rect 21058 2830 21158 2831
rect 21115 2794 21157 2830
rect 21006 2771 21157 2794
rect 21006 2753 21024 2771
rect 21042 2756 21157 2771
rect 21042 2753 21063 2756
rect 21006 2734 21063 2753
rect 15719 2677 15875 2681
rect 15719 2659 15739 2677
rect 15757 2659 15875 2677
rect 10693 2613 10811 2631
rect 10829 2613 10849 2631
rect 10693 2609 10849 2613
rect 10395 2608 10495 2609
rect 10452 2572 10494 2608
rect 10788 2593 10849 2609
rect 10343 2549 10494 2572
rect 15719 2638 15875 2659
rect 15775 2637 15875 2638
rect 15975 2668 16126 2691
rect 15832 2601 15874 2637
rect 15975 2632 16017 2668
rect 15723 2578 15874 2601
rect 15974 2631 16074 2632
rect 15974 2610 16130 2631
rect 21000 2660 21061 2676
rect 21000 2656 21156 2660
rect 21000 2638 21020 2656
rect 21038 2638 21156 2656
rect 15974 2592 16092 2610
rect 16110 2592 16130 2610
rect 15974 2588 16130 2592
rect 35 2399 186 2422
rect 35 2363 77 2399
rect 34 2362 134 2363
rect 34 2341 190 2362
rect 5410 2419 5467 2438
rect 5410 2416 5431 2419
rect 5060 2391 5121 2407
rect 5316 2401 5431 2416
rect 5449 2401 5467 2419
rect 10343 2531 10361 2549
rect 10379 2534 10494 2549
rect 10379 2531 10400 2534
rect 10343 2512 10400 2531
rect 10790 2448 10847 2467
rect 10790 2445 10811 2448
rect 10696 2430 10811 2445
rect 10829 2430 10847 2448
rect 15723 2560 15741 2578
rect 15759 2563 15874 2578
rect 16069 2572 16130 2588
rect 15759 2560 15780 2563
rect 15723 2541 15780 2560
rect 21000 2617 21156 2638
rect 21056 2616 21156 2617
rect 21113 2580 21155 2616
rect 21004 2557 21155 2580
rect 5060 2387 5216 2391
rect 5060 2369 5080 2387
rect 5098 2369 5216 2387
rect 34 2323 152 2341
rect 170 2323 190 2341
rect 34 2319 190 2323
rect 129 2303 190 2319
rect 5060 2348 5216 2369
rect 5116 2347 5216 2348
rect 5316 2378 5467 2401
rect 5173 2311 5215 2347
rect 5316 2342 5358 2378
rect 5064 2288 5215 2311
rect 5315 2341 5415 2342
rect 5315 2320 5471 2341
rect 10696 2407 10847 2430
rect 10341 2370 10402 2386
rect 10696 2371 10738 2407
rect 10695 2370 10795 2371
rect 10341 2366 10497 2370
rect 10341 2348 10361 2366
rect 10379 2348 10497 2366
rect 5315 2302 5433 2320
rect 5451 2302 5471 2320
rect 5315 2298 5471 2302
rect 127 2226 184 2245
rect 127 2223 148 2226
rect 33 2208 148 2223
rect 166 2208 184 2226
rect 33 2185 184 2208
rect 33 2149 75 2185
rect 32 2148 132 2149
rect 32 2127 188 2148
rect 5064 2270 5082 2288
rect 5100 2273 5215 2288
rect 5410 2282 5471 2298
rect 5100 2270 5121 2273
rect 5064 2251 5121 2270
rect 10341 2327 10497 2348
rect 10695 2349 10851 2370
rect 16071 2427 16128 2446
rect 16071 2424 16092 2427
rect 15721 2399 15782 2415
rect 15977 2409 16092 2424
rect 16110 2409 16128 2427
rect 21004 2539 21022 2557
rect 21040 2542 21155 2557
rect 21040 2539 21061 2542
rect 21004 2520 21061 2539
rect 15721 2395 15877 2399
rect 15721 2377 15741 2395
rect 15759 2377 15877 2395
rect 10695 2331 10813 2349
rect 10831 2331 10851 2349
rect 10695 2327 10851 2331
rect 10397 2326 10497 2327
rect 10454 2290 10496 2326
rect 10790 2311 10851 2327
rect 15721 2356 15877 2377
rect 15777 2355 15877 2356
rect 15977 2386 16128 2409
rect 15834 2319 15876 2355
rect 15977 2350 16019 2386
rect 15725 2296 15876 2319
rect 15976 2349 16076 2350
rect 15976 2328 16132 2349
rect 21002 2378 21063 2394
rect 21002 2374 21158 2378
rect 21002 2356 21022 2374
rect 21040 2356 21158 2374
rect 15976 2310 16094 2328
rect 16112 2310 16132 2328
rect 15976 2306 16132 2310
rect 10345 2267 10496 2290
rect 5067 2190 5128 2206
rect 5408 2205 5465 2224
rect 5408 2202 5429 2205
rect 5067 2186 5223 2190
rect 5067 2168 5087 2186
rect 5105 2168 5223 2186
rect 32 2109 150 2127
rect 168 2109 188 2127
rect 32 2105 188 2109
rect 127 2089 188 2105
rect 5067 2147 5223 2168
rect 5123 2146 5223 2147
rect 5314 2187 5429 2202
rect 5447 2187 5465 2205
rect 5314 2164 5465 2187
rect 5180 2110 5222 2146
rect 5314 2128 5356 2164
rect 5071 2087 5222 2110
rect 5071 2069 5089 2087
rect 5107 2072 5222 2087
rect 5313 2127 5413 2128
rect 5313 2106 5469 2127
rect 10345 2249 10363 2267
rect 10381 2252 10496 2267
rect 10381 2249 10402 2252
rect 10345 2230 10402 2249
rect 10788 2234 10845 2253
rect 10788 2231 10809 2234
rect 10694 2216 10809 2231
rect 10827 2216 10845 2234
rect 10694 2193 10845 2216
rect 10348 2169 10409 2185
rect 10348 2165 10504 2169
rect 10348 2147 10368 2165
rect 10386 2147 10504 2165
rect 10694 2157 10736 2193
rect 5313 2088 5431 2106
rect 5449 2088 5469 2106
rect 5313 2084 5469 2088
rect 5107 2069 5128 2072
rect 5071 2050 5128 2069
rect 5408 2068 5469 2084
rect 127 1944 184 1963
rect 127 1941 148 1944
rect 33 1926 148 1941
rect 166 1926 184 1944
rect 33 1903 184 1926
rect 33 1867 75 1903
rect 10348 2126 10504 2147
rect 10404 2125 10504 2126
rect 10693 2156 10793 2157
rect 10693 2135 10849 2156
rect 15725 2278 15743 2296
rect 15761 2281 15876 2296
rect 16071 2290 16132 2306
rect 15761 2278 15782 2281
rect 15725 2259 15782 2278
rect 21002 2335 21158 2356
rect 21058 2334 21158 2335
rect 21115 2298 21157 2334
rect 21006 2275 21157 2298
rect 15728 2198 15789 2214
rect 16069 2213 16126 2232
rect 16069 2210 16090 2213
rect 15728 2194 15884 2198
rect 15728 2176 15748 2194
rect 15766 2176 15884 2194
rect 32 1866 132 1867
rect 32 1845 188 1866
rect 10461 2089 10503 2125
rect 10693 2117 10811 2135
rect 10829 2117 10849 2135
rect 10693 2113 10849 2117
rect 10788 2097 10849 2113
rect 10352 2066 10503 2089
rect 15728 2155 15884 2176
rect 15784 2154 15884 2155
rect 15975 2195 16090 2210
rect 16108 2195 16126 2213
rect 15975 2172 16126 2195
rect 10352 2048 10370 2066
rect 10388 2051 10503 2066
rect 10388 2048 10409 2051
rect 10352 2029 10409 2048
rect 5067 1908 5128 1924
rect 5408 1923 5465 1942
rect 5408 1920 5429 1923
rect 5067 1904 5223 1908
rect 5067 1886 5087 1904
rect 5105 1886 5223 1904
rect 32 1827 150 1845
rect 168 1827 188 1845
rect 32 1823 188 1827
rect 127 1807 188 1823
rect 134 1743 191 1762
rect 134 1740 155 1743
rect 40 1725 155 1740
rect 173 1725 191 1743
rect 5067 1865 5223 1886
rect 5123 1864 5223 1865
rect 5314 1905 5429 1920
rect 5447 1905 5465 1923
rect 5314 1882 5465 1905
rect 5180 1828 5222 1864
rect 5314 1846 5356 1882
rect 15841 2118 15883 2154
rect 15975 2136 16017 2172
rect 15732 2095 15883 2118
rect 15732 2077 15750 2095
rect 15768 2080 15883 2095
rect 15974 2135 16074 2136
rect 15974 2114 16130 2135
rect 21006 2257 21024 2275
rect 21042 2260 21157 2275
rect 21042 2257 21063 2260
rect 21006 2238 21063 2257
rect 21009 2177 21070 2193
rect 21009 2173 21165 2177
rect 21009 2155 21029 2173
rect 21047 2155 21165 2173
rect 15974 2096 16092 2114
rect 16110 2096 16130 2114
rect 15974 2092 16130 2096
rect 15768 2077 15789 2080
rect 15732 2058 15789 2077
rect 16069 2076 16130 2092
rect 10788 1952 10845 1971
rect 10788 1949 10809 1952
rect 10694 1934 10809 1949
rect 10827 1934 10845 1952
rect 5071 1805 5222 1828
rect 5071 1787 5089 1805
rect 5107 1790 5222 1805
rect 5313 1845 5413 1846
rect 5313 1824 5469 1845
rect 10694 1911 10845 1934
rect 10348 1887 10409 1903
rect 10348 1883 10504 1887
rect 10348 1865 10368 1883
rect 10386 1865 10504 1883
rect 10694 1875 10736 1911
rect 21009 2134 21165 2155
rect 21065 2133 21165 2134
rect 5313 1806 5431 1824
rect 5449 1806 5469 1824
rect 5313 1802 5469 1806
rect 5107 1787 5128 1790
rect 5071 1768 5128 1787
rect 5408 1786 5469 1802
rect 40 1702 191 1725
rect 40 1666 82 1702
rect 39 1665 139 1666
rect 39 1644 195 1665
rect 5415 1722 5472 1741
rect 5415 1719 5436 1722
rect 39 1626 157 1644
rect 175 1626 195 1644
rect 39 1622 195 1626
rect 134 1606 195 1622
rect 5065 1694 5126 1710
rect 5321 1704 5436 1719
rect 5454 1704 5472 1722
rect 10348 1844 10504 1865
rect 10404 1843 10504 1844
rect 10693 1874 10793 1875
rect 10693 1853 10849 1874
rect 21122 2097 21164 2133
rect 21013 2074 21164 2097
rect 21013 2056 21031 2074
rect 21049 2059 21164 2074
rect 21049 2056 21070 2059
rect 21013 2037 21070 2056
rect 15728 1916 15789 1932
rect 16069 1931 16126 1950
rect 16069 1928 16090 1931
rect 15728 1912 15884 1916
rect 15728 1894 15748 1912
rect 15766 1894 15884 1912
rect 10461 1807 10503 1843
rect 10693 1835 10811 1853
rect 10829 1835 10849 1853
rect 10693 1831 10849 1835
rect 10788 1815 10849 1831
rect 10352 1784 10503 1807
rect 10352 1766 10370 1784
rect 10388 1769 10503 1784
rect 10388 1766 10409 1769
rect 10352 1747 10409 1766
rect 10795 1751 10852 1770
rect 10795 1748 10816 1751
rect 10701 1733 10816 1748
rect 10834 1733 10852 1751
rect 15728 1873 15884 1894
rect 15784 1872 15884 1873
rect 15975 1913 16090 1928
rect 16108 1913 16126 1931
rect 15975 1890 16126 1913
rect 15841 1836 15883 1872
rect 15975 1854 16017 1890
rect 15732 1813 15883 1836
rect 15732 1795 15750 1813
rect 15768 1798 15883 1813
rect 15974 1853 16074 1854
rect 15974 1832 16130 1853
rect 21009 1895 21070 1911
rect 21009 1891 21165 1895
rect 21009 1873 21029 1891
rect 21047 1873 21165 1891
rect 15974 1814 16092 1832
rect 16110 1814 16130 1832
rect 15974 1810 16130 1814
rect 15768 1795 15789 1798
rect 15732 1776 15789 1795
rect 16069 1794 16130 1810
rect 5065 1690 5221 1694
rect 5065 1672 5085 1690
rect 5103 1672 5221 1690
rect 5065 1651 5221 1672
rect 5121 1650 5221 1651
rect 5321 1681 5472 1704
rect 5178 1614 5220 1650
rect 5321 1645 5363 1681
rect 5069 1591 5220 1614
rect 5320 1644 5420 1645
rect 5320 1623 5476 1644
rect 10701 1710 10852 1733
rect 5320 1605 5438 1623
rect 5456 1605 5476 1623
rect 5320 1601 5476 1605
rect 5069 1573 5087 1591
rect 5105 1576 5220 1591
rect 5415 1585 5476 1601
rect 10346 1673 10407 1689
rect 10701 1674 10743 1710
rect 10700 1673 10800 1674
rect 10346 1669 10502 1673
rect 10346 1651 10366 1669
rect 10384 1651 10502 1669
rect 10346 1630 10502 1651
rect 10700 1652 10856 1673
rect 16076 1730 16133 1749
rect 16076 1727 16097 1730
rect 10700 1634 10818 1652
rect 10836 1634 10856 1652
rect 10700 1630 10856 1634
rect 10402 1629 10502 1630
rect 5105 1573 5126 1576
rect 5069 1554 5126 1573
rect 10459 1593 10501 1629
rect 10795 1614 10856 1630
rect 15726 1702 15787 1718
rect 15982 1712 16097 1727
rect 16115 1712 16133 1730
rect 21009 1852 21165 1873
rect 21065 1851 21165 1852
rect 21122 1815 21164 1851
rect 21013 1792 21164 1815
rect 21013 1774 21031 1792
rect 21049 1777 21164 1792
rect 21049 1774 21070 1777
rect 21013 1755 21070 1774
rect 15726 1698 15882 1702
rect 15726 1680 15746 1698
rect 15764 1680 15882 1698
rect 15726 1659 15882 1680
rect 15782 1658 15882 1659
rect 15982 1689 16133 1712
rect 10350 1570 10501 1593
rect 10350 1552 10368 1570
rect 10386 1555 10501 1570
rect 10386 1552 10407 1555
rect 10350 1533 10407 1552
rect 15839 1622 15881 1658
rect 15982 1653 16024 1689
rect 15730 1599 15881 1622
rect 15981 1652 16081 1653
rect 15981 1631 16137 1652
rect 15981 1613 16099 1631
rect 16117 1613 16137 1631
rect 15981 1609 16137 1613
rect 15730 1581 15748 1599
rect 15766 1584 15881 1599
rect 16076 1593 16137 1609
rect 21007 1681 21068 1697
rect 21007 1677 21163 1681
rect 21007 1659 21027 1677
rect 21045 1659 21163 1677
rect 21007 1638 21163 1659
rect 21063 1637 21163 1638
rect 15766 1581 15787 1584
rect 15730 1562 15787 1581
rect 21120 1601 21162 1637
rect 21011 1578 21162 1601
rect 21011 1560 21029 1578
rect 21047 1563 21162 1578
rect 21047 1560 21068 1563
rect 21011 1541 21068 1560
rect 134 1459 191 1478
rect 134 1456 155 1459
rect 40 1441 155 1456
rect 173 1441 191 1459
rect 40 1418 191 1441
rect 40 1382 82 1418
rect 5415 1438 5472 1457
rect 5415 1435 5436 1438
rect 39 1381 139 1382
rect 39 1360 195 1381
rect 39 1342 157 1360
rect 175 1342 195 1360
rect 39 1338 195 1342
rect 134 1322 195 1338
rect 5065 1410 5126 1426
rect 5321 1420 5436 1435
rect 5454 1420 5472 1438
rect 5065 1406 5221 1410
rect 5065 1388 5085 1406
rect 5103 1388 5221 1406
rect 5065 1367 5221 1388
rect 5121 1366 5221 1367
rect 5321 1397 5472 1420
rect 5178 1330 5220 1366
rect 5321 1361 5363 1397
rect 10795 1467 10852 1486
rect 10795 1464 10816 1467
rect 10701 1449 10816 1464
rect 10834 1449 10852 1467
rect 10701 1426 10852 1449
rect 5069 1307 5220 1330
rect 5320 1360 5420 1361
rect 5320 1339 5476 1360
rect 5320 1321 5438 1339
rect 5456 1321 5476 1339
rect 5320 1317 5476 1321
rect 132 1245 189 1264
rect 132 1242 153 1245
rect 38 1227 153 1242
rect 171 1227 189 1245
rect 38 1204 189 1227
rect 38 1168 80 1204
rect 37 1167 137 1168
rect 37 1146 193 1167
rect 5069 1289 5087 1307
rect 5105 1292 5220 1307
rect 5415 1301 5476 1317
rect 10346 1389 10407 1405
rect 10701 1390 10743 1426
rect 16076 1446 16133 1465
rect 16076 1443 16097 1446
rect 10700 1389 10800 1390
rect 10346 1385 10502 1389
rect 10346 1367 10366 1385
rect 10384 1367 10502 1385
rect 5105 1289 5126 1292
rect 5069 1270 5126 1289
rect 10346 1346 10502 1367
rect 10700 1368 10856 1389
rect 10700 1350 10818 1368
rect 10836 1350 10856 1368
rect 10700 1346 10856 1350
rect 10402 1345 10502 1346
rect 10459 1309 10501 1345
rect 10795 1330 10856 1346
rect 15726 1418 15787 1434
rect 15982 1428 16097 1443
rect 16115 1428 16133 1446
rect 15726 1414 15882 1418
rect 15726 1396 15746 1414
rect 15764 1396 15882 1414
rect 10350 1286 10501 1309
rect 15726 1375 15882 1396
rect 15782 1374 15882 1375
rect 15982 1405 16133 1428
rect 15839 1338 15881 1374
rect 15982 1369 16024 1405
rect 15730 1315 15881 1338
rect 15981 1368 16081 1369
rect 15981 1347 16137 1368
rect 15981 1329 16099 1347
rect 16117 1329 16137 1347
rect 15981 1325 16137 1329
rect 5072 1209 5133 1225
rect 5413 1224 5470 1243
rect 5413 1221 5434 1224
rect 5072 1205 5228 1209
rect 5072 1187 5092 1205
rect 5110 1187 5228 1205
rect 37 1128 155 1146
rect 173 1128 193 1146
rect 37 1124 193 1128
rect 132 1108 193 1124
rect 5072 1166 5228 1187
rect 5128 1165 5228 1166
rect 5319 1206 5434 1221
rect 5452 1206 5470 1224
rect 5319 1183 5470 1206
rect 5185 1129 5227 1165
rect 5319 1147 5361 1183
rect 5076 1106 5227 1129
rect 5076 1088 5094 1106
rect 5112 1091 5227 1106
rect 5318 1146 5418 1147
rect 5318 1125 5474 1146
rect 10350 1268 10368 1286
rect 10386 1271 10501 1286
rect 10386 1268 10407 1271
rect 10350 1249 10407 1268
rect 10793 1253 10850 1272
rect 10793 1250 10814 1253
rect 10699 1235 10814 1250
rect 10832 1235 10850 1253
rect 10699 1212 10850 1235
rect 10353 1188 10414 1204
rect 10353 1184 10509 1188
rect 10353 1166 10373 1184
rect 10391 1166 10509 1184
rect 10699 1176 10741 1212
rect 5318 1107 5436 1125
rect 5454 1107 5474 1125
rect 5318 1103 5474 1107
rect 5112 1088 5133 1091
rect 5076 1069 5133 1088
rect 5413 1087 5474 1103
rect 132 963 189 982
rect 132 960 153 963
rect 38 945 153 960
rect 171 945 189 963
rect 38 922 189 945
rect 38 886 80 922
rect 10353 1145 10509 1166
rect 10409 1144 10509 1145
rect 10698 1175 10798 1176
rect 10698 1154 10854 1175
rect 15730 1297 15748 1315
rect 15766 1300 15881 1315
rect 16076 1309 16137 1325
rect 21007 1397 21068 1413
rect 21007 1393 21163 1397
rect 21007 1375 21027 1393
rect 21045 1375 21163 1393
rect 15766 1297 15787 1300
rect 15730 1278 15787 1297
rect 21007 1354 21163 1375
rect 21063 1353 21163 1354
rect 21120 1317 21162 1353
rect 21011 1294 21162 1317
rect 15733 1217 15794 1233
rect 16074 1232 16131 1251
rect 16074 1229 16095 1232
rect 15733 1213 15889 1217
rect 15733 1195 15753 1213
rect 15771 1195 15889 1213
rect 37 885 137 886
rect 37 864 193 885
rect 10466 1108 10508 1144
rect 10698 1136 10816 1154
rect 10834 1136 10854 1154
rect 10698 1132 10854 1136
rect 10793 1116 10854 1132
rect 10357 1085 10508 1108
rect 15733 1174 15889 1195
rect 15789 1173 15889 1174
rect 15980 1214 16095 1229
rect 16113 1214 16131 1232
rect 15980 1191 16131 1214
rect 10357 1067 10375 1085
rect 10393 1070 10508 1085
rect 10393 1067 10414 1070
rect 10357 1048 10414 1067
rect 5072 927 5133 943
rect 5413 942 5470 961
rect 5413 939 5434 942
rect 5072 923 5228 927
rect 5072 905 5092 923
rect 5110 905 5228 923
rect 37 846 155 864
rect 173 846 193 864
rect 37 842 193 846
rect 132 826 193 842
rect 139 762 196 781
rect 139 759 160 762
rect 45 744 160 759
rect 178 744 196 762
rect 5072 884 5228 905
rect 5128 883 5228 884
rect 5319 924 5434 939
rect 5452 924 5470 942
rect 5319 901 5470 924
rect 5185 847 5227 883
rect 5319 865 5361 901
rect 15846 1137 15888 1173
rect 15980 1155 16022 1191
rect 15737 1114 15888 1137
rect 15737 1096 15755 1114
rect 15773 1099 15888 1114
rect 15979 1154 16079 1155
rect 15979 1133 16135 1154
rect 21011 1276 21029 1294
rect 21047 1279 21162 1294
rect 21047 1276 21068 1279
rect 21011 1257 21068 1276
rect 21014 1196 21075 1212
rect 21014 1192 21170 1196
rect 21014 1174 21034 1192
rect 21052 1174 21170 1192
rect 15979 1115 16097 1133
rect 16115 1115 16135 1133
rect 15979 1111 16135 1115
rect 15773 1096 15794 1099
rect 15737 1077 15794 1096
rect 16074 1095 16135 1111
rect 10793 971 10850 990
rect 10793 968 10814 971
rect 10699 953 10814 968
rect 10832 953 10850 971
rect 5076 824 5227 847
rect 5076 806 5094 824
rect 5112 809 5227 824
rect 5318 864 5418 865
rect 5318 843 5474 864
rect 10699 930 10850 953
rect 10353 906 10414 922
rect 10353 902 10509 906
rect 10353 884 10373 902
rect 10391 884 10509 902
rect 10699 894 10741 930
rect 21014 1153 21170 1174
rect 21070 1152 21170 1153
rect 5318 825 5436 843
rect 5454 825 5474 843
rect 5318 821 5474 825
rect 5112 806 5133 809
rect 5076 787 5133 806
rect 5413 805 5474 821
rect 45 721 196 744
rect 45 685 87 721
rect 44 684 144 685
rect 44 663 200 684
rect 5420 741 5477 760
rect 5420 738 5441 741
rect 5070 713 5131 729
rect 5326 723 5441 738
rect 5459 723 5477 741
rect 10353 863 10509 884
rect 10409 862 10509 863
rect 10698 893 10798 894
rect 10698 872 10854 893
rect 21127 1116 21169 1152
rect 21018 1093 21169 1116
rect 21018 1075 21036 1093
rect 21054 1078 21169 1093
rect 21054 1075 21075 1078
rect 21018 1056 21075 1075
rect 15733 935 15794 951
rect 16074 950 16131 969
rect 16074 947 16095 950
rect 15733 931 15889 935
rect 15733 913 15753 931
rect 15771 913 15889 931
rect 10466 826 10508 862
rect 10698 854 10816 872
rect 10834 854 10854 872
rect 10698 850 10854 854
rect 10793 834 10854 850
rect 10357 803 10508 826
rect 10357 785 10375 803
rect 10393 788 10508 803
rect 10393 785 10414 788
rect 10357 766 10414 785
rect 10800 770 10857 789
rect 10800 767 10821 770
rect 10706 752 10821 767
rect 10839 752 10857 770
rect 15733 892 15889 913
rect 15789 891 15889 892
rect 15980 932 16095 947
rect 16113 932 16131 950
rect 15980 909 16131 932
rect 15846 855 15888 891
rect 15980 873 16022 909
rect 15737 832 15888 855
rect 15737 814 15755 832
rect 15773 817 15888 832
rect 15979 872 16079 873
rect 15979 851 16135 872
rect 21014 914 21075 930
rect 21014 910 21170 914
rect 21014 892 21034 910
rect 21052 892 21170 910
rect 15979 833 16097 851
rect 16115 833 16135 851
rect 15979 829 16135 833
rect 15773 814 15794 817
rect 15737 795 15794 814
rect 16074 813 16135 829
rect 10706 729 10857 752
rect 5070 709 5226 713
rect 5070 691 5090 709
rect 5108 691 5226 709
rect 44 645 162 663
rect 180 645 200 663
rect 44 641 200 645
rect 139 625 200 641
rect 5070 670 5226 691
rect 5126 669 5226 670
rect 5326 700 5477 723
rect 5183 633 5225 669
rect 5326 664 5368 700
rect 5074 610 5225 633
rect 5325 663 5425 664
rect 5325 642 5481 663
rect 10351 692 10412 708
rect 10706 693 10748 729
rect 10705 692 10805 693
rect 10351 688 10507 692
rect 10351 670 10371 688
rect 10389 670 10507 688
rect 5325 624 5443 642
rect 5461 624 5481 642
rect 5325 620 5481 624
rect 5074 592 5092 610
rect 5110 595 5225 610
rect 5420 604 5481 620
rect 10351 649 10507 670
rect 10705 671 10861 692
rect 16081 749 16138 768
rect 16081 746 16102 749
rect 15731 721 15792 737
rect 15987 731 16102 746
rect 16120 731 16138 749
rect 21014 871 21170 892
rect 21070 870 21170 871
rect 21127 834 21169 870
rect 21018 811 21169 834
rect 21018 793 21036 811
rect 21054 796 21169 811
rect 21054 793 21075 796
rect 21018 774 21075 793
rect 15731 717 15887 721
rect 15731 699 15751 717
rect 15769 699 15887 717
rect 10705 653 10823 671
rect 10841 653 10861 671
rect 10705 649 10861 653
rect 10407 648 10507 649
rect 10464 612 10506 648
rect 10800 633 10861 649
rect 15731 678 15887 699
rect 15787 677 15887 678
rect 15987 708 16138 731
rect 15844 641 15886 677
rect 15987 672 16029 708
rect 5110 592 5131 595
rect 5074 573 5131 592
rect 10355 589 10506 612
rect 10355 571 10373 589
rect 10391 574 10506 589
rect 15735 618 15886 641
rect 15986 671 16086 672
rect 15986 650 16142 671
rect 21012 700 21073 716
rect 21012 696 21168 700
rect 21012 678 21032 696
rect 21050 678 21168 696
rect 15986 632 16104 650
rect 16122 632 16142 650
rect 15986 628 16142 632
rect 15735 600 15753 618
rect 15771 603 15886 618
rect 16081 612 16142 628
rect 21012 657 21168 678
rect 21068 656 21168 657
rect 21125 620 21167 656
rect 15771 600 15792 603
rect 15735 581 15792 600
rect 21016 597 21167 620
rect 21016 579 21034 597
rect 21052 582 21167 597
rect 21052 579 21073 582
rect 10391 571 10412 574
rect 10355 552 10412 571
rect 21016 560 21073 579
<< locali >>
rect 110 8326 145 8374
rect 5038 8368 5434 8374
rect 4449 8350 5434 8368
rect 108 8317 145 8326
rect 108 8299 118 8317
rect 136 8299 145 8317
rect 108 8289 145 8299
rect 4031 8333 4199 8334
rect 4450 8333 4474 8350
rect 5038 8342 5434 8350
rect 10319 8358 10806 8388
rect 15699 8376 16095 8382
rect 15110 8358 16095 8376
rect 10319 8347 10355 8358
rect 4031 8307 4475 8333
rect 4031 8305 4199 8307
rect 111 8225 148 8227
rect 111 8224 759 8225
rect 110 8218 759 8224
rect 110 8200 120 8218
rect 138 8204 759 8218
rect 138 8200 148 8204
rect 589 8203 759 8204
rect 110 8190 148 8200
rect 110 8112 145 8190
rect 722 8180 759 8203
rect 106 8103 145 8112
rect 106 8085 116 8103
rect 134 8085 145 8103
rect 106 8079 145 8085
rect 301 8155 551 8179
rect 301 8084 338 8155
rect 453 8094 484 8095
rect 106 8075 143 8079
rect 301 8064 310 8084
rect 330 8064 338 8084
rect 301 8054 338 8064
rect 397 8084 484 8094
rect 397 8064 406 8084
rect 426 8064 484 8084
rect 397 8055 484 8064
rect 397 8054 434 8055
rect 109 8004 146 8013
rect 107 7986 118 8004
rect 136 7986 146 8004
rect 453 8002 484 8055
rect 514 8084 551 8155
rect 722 8160 1115 8180
rect 1135 8160 1138 8180
rect 722 8155 1138 8160
rect 722 8154 1063 8155
rect 666 8094 697 8095
rect 514 8064 523 8084
rect 543 8064 551 8084
rect 514 8054 551 8064
rect 610 8087 697 8094
rect 610 8084 671 8087
rect 610 8064 619 8084
rect 639 8067 671 8084
rect 692 8067 697 8087
rect 639 8064 697 8067
rect 610 8057 697 8064
rect 722 8084 759 8154
rect 1025 8153 1062 8154
rect 4031 8127 4058 8305
rect 4098 8267 4162 8279
rect 4438 8275 4475 8307
rect 4646 8306 4895 8328
rect 4646 8275 4683 8306
rect 4859 8304 4895 8306
rect 5038 8309 5076 8342
rect 4859 8275 4896 8304
rect 4098 8266 4133 8267
rect 4075 8261 4133 8266
rect 4075 8241 4078 8261
rect 4098 8247 4133 8261
rect 4153 8247 4162 8267
rect 4098 8239 4162 8247
rect 4124 8238 4162 8239
rect 4125 8237 4162 8238
rect 4228 8271 4264 8272
rect 4336 8271 4372 8272
rect 4228 8265 4372 8271
rect 4228 8263 4294 8265
rect 4228 8243 4236 8263
rect 4256 8244 4294 8263
rect 4316 8263 4372 8265
rect 4316 8244 4344 8263
rect 4256 8243 4344 8244
rect 4364 8243 4372 8263
rect 4228 8237 4372 8243
rect 4438 8267 4476 8275
rect 4544 8271 4580 8272
rect 4438 8247 4447 8267
rect 4467 8247 4476 8267
rect 4438 8238 4476 8247
rect 4495 8264 4580 8271
rect 4495 8244 4502 8264
rect 4523 8263 4580 8264
rect 4523 8244 4552 8263
rect 4495 8243 4552 8244
rect 4572 8243 4580 8263
rect 4438 8237 4475 8238
rect 4495 8237 4580 8243
rect 4646 8267 4684 8275
rect 4757 8271 4793 8272
rect 4646 8247 4655 8267
rect 4675 8247 4684 8267
rect 4646 8238 4684 8247
rect 4708 8263 4793 8271
rect 4708 8243 4765 8263
rect 4785 8243 4793 8263
rect 4646 8237 4683 8238
rect 4708 8237 4793 8243
rect 4859 8267 4897 8275
rect 4859 8247 4868 8267
rect 4888 8247 4897 8267
rect 4859 8238 4897 8247
rect 5038 8274 5074 8309
rect 5391 8305 5426 8342
rect 9730 8329 10355 8347
rect 10771 8334 10806 8358
rect 5389 8296 5426 8305
rect 5389 8278 5399 8296
rect 5417 8278 5426 8296
rect 5038 8264 5075 8274
rect 5389 8268 5426 8278
rect 9312 8312 9480 8313
rect 9731 8312 9755 8329
rect 9312 8286 9756 8312
rect 9312 8284 9480 8286
rect 5038 8246 5048 8264
rect 5066 8246 5075 8264
rect 4859 8237 4896 8238
rect 5038 8237 5075 8246
rect 4282 8216 4318 8237
rect 4708 8216 4739 8237
rect 4115 8212 4215 8216
rect 4115 8208 4177 8212
rect 4115 8182 4122 8208
rect 4148 8186 4177 8208
rect 4203 8186 4215 8212
rect 4148 8182 4215 8186
rect 4115 8179 4215 8182
rect 4283 8179 4318 8216
rect 4380 8213 4739 8216
rect 4380 8208 4602 8213
rect 4380 8184 4393 8208
rect 4417 8189 4602 8208
rect 4626 8189 4739 8213
rect 4417 8184 4739 8189
rect 4380 8180 4739 8184
rect 4806 8208 4955 8216
rect 4806 8188 4817 8208
rect 4837 8188 4955 8208
rect 5392 8204 5429 8206
rect 5392 8203 6040 8204
rect 4806 8181 4955 8188
rect 5391 8197 6040 8203
rect 4806 8180 4847 8181
rect 4130 8127 4167 8128
rect 4226 8127 4263 8128
rect 4282 8127 4318 8179
rect 4337 8127 4374 8128
rect 4030 8118 4168 8127
rect 2966 8100 2997 8103
rect 874 8094 910 8095
rect 722 8064 731 8084
rect 751 8064 759 8084
rect 610 8055 666 8057
rect 610 8054 647 8055
rect 722 8054 759 8064
rect 818 8084 966 8094
rect 1066 8091 1162 8093
rect 818 8064 827 8084
rect 847 8064 937 8084
rect 957 8064 966 8084
rect 818 8055 966 8064
rect 1024 8084 1162 8091
rect 1024 8064 1033 8084
rect 1053 8064 1162 8084
rect 1024 8055 1162 8064
rect 2966 8074 2973 8100
rect 2992 8074 2997 8100
rect 818 8054 855 8055
rect 874 8003 910 8055
rect 929 8054 966 8055
rect 1025 8054 1062 8055
rect 345 8001 386 8002
rect 107 7837 146 7986
rect 237 7994 386 8001
rect 237 7974 355 7994
rect 375 7974 386 7994
rect 237 7966 386 7974
rect 453 7998 812 8002
rect 453 7993 775 7998
rect 453 7969 566 7993
rect 590 7974 775 7993
rect 799 7974 812 7998
rect 590 7969 812 7974
rect 453 7966 812 7969
rect 874 7966 909 8003
rect 977 8000 1077 8003
rect 977 7996 1044 8000
rect 977 7970 989 7996
rect 1015 7974 1044 7996
rect 1070 7974 1077 8000
rect 1015 7970 1077 7974
rect 977 7966 1077 7970
rect 453 7945 484 7966
rect 874 7945 910 7966
rect 296 7944 333 7945
rect 295 7935 333 7944
rect 295 7915 304 7935
rect 324 7915 333 7935
rect 295 7907 333 7915
rect 399 7939 484 7945
rect 509 7944 546 7945
rect 399 7919 407 7939
rect 427 7919 484 7939
rect 399 7911 484 7919
rect 508 7935 546 7944
rect 508 7915 517 7935
rect 537 7915 546 7935
rect 399 7910 435 7911
rect 508 7907 546 7915
rect 612 7939 697 7945
rect 717 7944 754 7945
rect 612 7919 620 7939
rect 640 7938 697 7939
rect 640 7919 669 7938
rect 612 7918 669 7919
rect 690 7918 697 7938
rect 612 7911 697 7918
rect 716 7935 754 7944
rect 716 7915 725 7935
rect 745 7915 754 7935
rect 612 7910 648 7911
rect 716 7907 754 7915
rect 820 7940 964 7945
rect 820 7939 885 7940
rect 820 7919 828 7939
rect 848 7919 885 7939
rect 907 7939 964 7940
rect 907 7919 936 7939
rect 956 7919 964 7939
rect 820 7911 964 7919
rect 820 7910 856 7911
rect 928 7910 964 7911
rect 1030 7944 1067 7945
rect 1030 7943 1068 7944
rect 1030 7935 1094 7943
rect 1030 7915 1039 7935
rect 1059 7921 1094 7935
rect 1114 7921 1117 7941
rect 1059 7916 1117 7921
rect 1059 7915 1094 7916
rect 296 7878 333 7907
rect 297 7876 333 7878
rect 509 7876 546 7907
rect 297 7854 546 7876
rect 717 7875 754 7907
rect 1030 7903 1094 7915
rect 1134 7877 1161 8055
rect 993 7875 1161 7877
rect 717 7849 1161 7875
rect 1313 7974 1563 7998
rect 1313 7903 1350 7974
rect 1465 7913 1496 7914
rect 1313 7883 1322 7903
rect 1342 7883 1350 7903
rect 1313 7873 1350 7883
rect 1409 7903 1496 7913
rect 1409 7883 1418 7903
rect 1438 7883 1496 7903
rect 1409 7874 1496 7883
rect 1409 7873 1446 7874
rect 717 7839 739 7849
rect 993 7848 1161 7849
rect 677 7837 739 7839
rect 107 7830 739 7837
rect 106 7821 739 7830
rect 1465 7821 1496 7874
rect 1526 7903 1563 7974
rect 1734 7979 2127 7999
rect 2147 7979 2150 7999
rect 1734 7974 2150 7979
rect 1734 7973 2075 7974
rect 1678 7913 1709 7914
rect 1526 7883 1535 7903
rect 1555 7883 1563 7903
rect 1526 7873 1563 7883
rect 1622 7906 1709 7913
rect 1622 7903 1683 7906
rect 1622 7883 1631 7903
rect 1651 7886 1683 7903
rect 1704 7886 1709 7906
rect 1651 7883 1709 7886
rect 1622 7876 1709 7883
rect 1734 7903 1771 7973
rect 2037 7972 2074 7973
rect 1886 7913 1922 7914
rect 1734 7883 1743 7903
rect 1763 7883 1771 7903
rect 1622 7874 1678 7876
rect 1622 7873 1659 7874
rect 1734 7873 1771 7883
rect 1830 7903 1978 7913
rect 2078 7910 2174 7912
rect 1830 7883 1839 7903
rect 1859 7883 1949 7903
rect 1969 7883 1978 7903
rect 1830 7874 1978 7883
rect 2036 7903 2174 7910
rect 2036 7883 2045 7903
rect 2065 7883 2174 7903
rect 2036 7874 2174 7883
rect 1830 7873 1867 7874
rect 1886 7822 1922 7874
rect 1941 7873 1978 7874
rect 2037 7873 2074 7874
rect 106 7803 116 7821
rect 134 7820 739 7821
rect 1357 7820 1398 7821
rect 134 7815 155 7820
rect 134 7803 146 7815
rect 1249 7813 1398 7820
rect 106 7795 146 7803
rect 189 7802 215 7803
rect 106 7793 143 7795
rect 189 7784 743 7802
rect 1249 7793 1367 7813
rect 1387 7793 1398 7813
rect 1249 7785 1398 7793
rect 1465 7817 1824 7821
rect 1465 7812 1787 7817
rect 1465 7788 1578 7812
rect 1602 7793 1787 7812
rect 1811 7793 1824 7817
rect 1602 7788 1824 7793
rect 1465 7785 1824 7788
rect 1886 7785 1921 7822
rect 1989 7819 2089 7822
rect 1989 7815 2056 7819
rect 1989 7789 2001 7815
rect 2027 7793 2056 7815
rect 2082 7793 2089 7819
rect 2027 7789 2089 7793
rect 1989 7785 2089 7789
rect 109 7725 146 7731
rect 189 7725 215 7784
rect 722 7765 743 7784
rect 109 7722 215 7725
rect 109 7704 118 7722
rect 136 7708 215 7722
rect 300 7740 550 7764
rect 136 7706 212 7708
rect 136 7704 146 7706
rect 109 7694 146 7704
rect 114 7629 145 7694
rect 300 7669 337 7740
rect 452 7679 483 7680
rect 300 7649 309 7669
rect 329 7649 337 7669
rect 300 7639 337 7649
rect 396 7669 483 7679
rect 396 7649 405 7669
rect 425 7649 483 7669
rect 396 7640 483 7649
rect 396 7639 433 7640
rect 113 7620 150 7629
rect 113 7602 123 7620
rect 141 7602 150 7620
rect 113 7592 150 7602
rect 452 7587 483 7640
rect 513 7669 550 7740
rect 721 7745 1114 7765
rect 1134 7745 1137 7765
rect 1465 7764 1496 7785
rect 1886 7764 1922 7785
rect 1308 7763 1345 7764
rect 721 7740 1137 7745
rect 1307 7754 1345 7763
rect 721 7739 1062 7740
rect 665 7679 696 7680
rect 513 7649 522 7669
rect 542 7649 550 7669
rect 513 7639 550 7649
rect 609 7672 696 7679
rect 609 7669 670 7672
rect 609 7649 618 7669
rect 638 7652 670 7669
rect 691 7652 696 7672
rect 638 7649 696 7652
rect 609 7642 696 7649
rect 721 7669 758 7739
rect 1024 7738 1061 7739
rect 1307 7734 1316 7754
rect 1336 7734 1345 7754
rect 1307 7726 1345 7734
rect 1411 7758 1496 7764
rect 1521 7763 1558 7764
rect 1411 7738 1419 7758
rect 1439 7738 1496 7758
rect 1411 7730 1496 7738
rect 1520 7754 1558 7763
rect 1520 7734 1529 7754
rect 1549 7734 1558 7754
rect 1411 7729 1447 7730
rect 1520 7726 1558 7734
rect 1624 7758 1709 7764
rect 1729 7763 1766 7764
rect 1624 7738 1632 7758
rect 1652 7757 1709 7758
rect 1652 7738 1681 7757
rect 1624 7737 1681 7738
rect 1702 7737 1709 7757
rect 1624 7730 1709 7737
rect 1728 7754 1766 7763
rect 1728 7734 1737 7754
rect 1757 7734 1766 7754
rect 1624 7729 1660 7730
rect 1728 7726 1766 7734
rect 1832 7758 1976 7764
rect 1832 7738 1840 7758
rect 1860 7738 1892 7758
rect 1916 7738 1948 7758
rect 1968 7738 1976 7758
rect 1832 7730 1976 7738
rect 1832 7729 1868 7730
rect 1940 7729 1976 7730
rect 2042 7763 2079 7764
rect 2042 7762 2080 7763
rect 2042 7754 2106 7762
rect 2042 7734 2051 7754
rect 2071 7740 2106 7754
rect 2126 7740 2129 7760
rect 2071 7735 2129 7740
rect 2071 7734 2106 7735
rect 1308 7697 1345 7726
rect 1309 7695 1345 7697
rect 1521 7695 1558 7726
rect 873 7679 909 7680
rect 721 7649 730 7669
rect 750 7649 758 7669
rect 609 7640 665 7642
rect 609 7639 646 7640
rect 721 7639 758 7649
rect 817 7669 965 7679
rect 1065 7676 1161 7678
rect 817 7649 826 7669
rect 846 7649 936 7669
rect 956 7649 965 7669
rect 817 7640 965 7649
rect 1023 7669 1161 7676
rect 1309 7673 1558 7695
rect 1729 7694 1766 7726
rect 2042 7722 2106 7734
rect 2146 7696 2173 7874
rect 2005 7694 2173 7696
rect 1729 7690 2173 7694
rect 1023 7649 1032 7669
rect 1052 7649 1161 7669
rect 1729 7671 1778 7690
rect 1798 7671 2173 7690
rect 1729 7668 2173 7671
rect 2005 7667 2173 7668
rect 2873 7681 2902 7683
rect 2873 7676 2905 7681
rect 2873 7658 2880 7676
rect 2900 7658 2905 7676
rect 2966 7680 2997 8074
rect 3018 8099 3186 8100
rect 3018 8096 3462 8099
rect 3018 8077 3393 8096
rect 3413 8077 3462 8096
rect 4030 8098 4139 8118
rect 4159 8098 4168 8118
rect 3018 8073 3462 8077
rect 3018 8071 3186 8073
rect 3018 7893 3045 8071
rect 3085 8033 3149 8045
rect 3425 8041 3462 8073
rect 3633 8072 3882 8094
rect 4030 8091 4168 8098
rect 4226 8118 4374 8127
rect 4226 8098 4235 8118
rect 4255 8098 4345 8118
rect 4365 8098 4374 8118
rect 4030 8089 4126 8091
rect 4226 8088 4374 8098
rect 4433 8118 4470 8128
rect 4545 8127 4582 8128
rect 4526 8125 4582 8127
rect 4433 8098 4441 8118
rect 4461 8098 4470 8118
rect 4282 8087 4318 8088
rect 3633 8041 3670 8072
rect 3846 8070 3882 8072
rect 3846 8041 3883 8070
rect 3085 8032 3120 8033
rect 3062 8027 3120 8032
rect 3062 8007 3065 8027
rect 3085 8013 3120 8027
rect 3140 8013 3149 8033
rect 3085 8005 3149 8013
rect 3111 8004 3149 8005
rect 3112 8003 3149 8004
rect 3215 8037 3251 8038
rect 3323 8037 3359 8038
rect 3215 8029 3359 8037
rect 3215 8009 3223 8029
rect 3243 8028 3331 8029
rect 3243 8009 3276 8028
rect 3215 8008 3276 8009
rect 3300 8009 3331 8028
rect 3351 8009 3359 8029
rect 3300 8008 3359 8009
rect 3215 8003 3359 8008
rect 3425 8033 3463 8041
rect 3531 8037 3567 8038
rect 3425 8013 3434 8033
rect 3454 8013 3463 8033
rect 3425 8004 3463 8013
rect 3482 8030 3567 8037
rect 3482 8010 3489 8030
rect 3510 8029 3567 8030
rect 3510 8010 3539 8029
rect 3482 8009 3539 8010
rect 3559 8009 3567 8029
rect 3425 8003 3462 8004
rect 3482 8003 3567 8009
rect 3633 8033 3671 8041
rect 3744 8037 3780 8038
rect 3633 8013 3642 8033
rect 3662 8013 3671 8033
rect 3633 8004 3671 8013
rect 3695 8029 3780 8037
rect 3695 8009 3752 8029
rect 3772 8009 3780 8029
rect 3633 8003 3670 8004
rect 3695 8003 3780 8009
rect 3846 8033 3884 8041
rect 3846 8013 3855 8033
rect 3875 8013 3884 8033
rect 4130 8028 4167 8029
rect 4433 8028 4470 8098
rect 4495 8118 4582 8125
rect 4495 8115 4553 8118
rect 4495 8095 4500 8115
rect 4521 8098 4553 8115
rect 4573 8098 4582 8118
rect 4521 8095 4582 8098
rect 4495 8088 4582 8095
rect 4641 8118 4678 8128
rect 4641 8098 4649 8118
rect 4669 8098 4678 8118
rect 4495 8087 4526 8088
rect 4129 8027 4470 8028
rect 3846 8004 3884 8013
rect 4054 8022 4470 8027
rect 3846 8003 3883 8004
rect 3269 7982 3305 8003
rect 3695 7982 3726 8003
rect 4054 8002 4057 8022
rect 4077 8002 4470 8022
rect 4641 8027 4678 8098
rect 4708 8127 4739 8180
rect 5391 8179 5401 8197
rect 5419 8183 6040 8197
rect 5419 8179 5429 8183
rect 5870 8182 6040 8183
rect 5041 8165 5078 8175
rect 5041 8147 5050 8165
rect 5068 8147 5078 8165
rect 5041 8138 5078 8147
rect 5391 8169 5429 8179
rect 4758 8127 4795 8128
rect 4708 8118 4795 8127
rect 4708 8098 4766 8118
rect 4786 8098 4795 8118
rect 4708 8088 4795 8098
rect 4854 8118 4891 8128
rect 4854 8098 4862 8118
rect 4882 8098 4891 8118
rect 4708 8087 4739 8088
rect 4854 8027 4891 8098
rect 5046 8073 5077 8138
rect 5391 8091 5426 8169
rect 6003 8159 6040 8182
rect 5387 8082 5426 8091
rect 5045 8063 5082 8073
rect 5045 8061 5055 8063
rect 4979 8059 5055 8061
rect 4641 8003 4891 8027
rect 4976 8045 5055 8059
rect 5073 8045 5082 8063
rect 5387 8064 5397 8082
rect 5415 8064 5426 8082
rect 5387 8058 5426 8064
rect 5582 8134 5832 8158
rect 5582 8063 5619 8134
rect 5734 8073 5765 8074
rect 5387 8054 5424 8058
rect 4976 8042 5082 8045
rect 4448 7983 4469 8002
rect 4976 7983 5002 8042
rect 5045 8036 5082 8042
rect 5582 8043 5591 8063
rect 5611 8043 5619 8063
rect 5582 8033 5619 8043
rect 5678 8063 5765 8073
rect 5678 8043 5687 8063
rect 5707 8043 5765 8063
rect 5678 8034 5765 8043
rect 5678 8033 5715 8034
rect 5390 7983 5427 7992
rect 3102 7978 3202 7982
rect 3102 7974 3164 7978
rect 3102 7948 3109 7974
rect 3135 7952 3164 7974
rect 3190 7952 3202 7978
rect 3135 7948 3202 7952
rect 3102 7945 3202 7948
rect 3270 7945 3305 7982
rect 3367 7979 3726 7982
rect 3367 7974 3589 7979
rect 3367 7950 3380 7974
rect 3404 7955 3589 7974
rect 3613 7955 3726 7979
rect 3404 7950 3726 7955
rect 3367 7946 3726 7950
rect 3793 7974 3942 7982
rect 3793 7954 3804 7974
rect 3824 7954 3942 7974
rect 4448 7965 5002 7983
rect 5048 7972 5085 7974
rect 4976 7964 5002 7965
rect 5045 7964 5085 7972
rect 3793 7947 3942 7954
rect 5045 7952 5057 7964
rect 5036 7947 5057 7952
rect 3793 7946 3834 7947
rect 4452 7946 5057 7947
rect 5075 7946 5085 7964
rect 3117 7893 3154 7894
rect 3213 7893 3250 7894
rect 3269 7893 3305 7945
rect 3324 7893 3361 7894
rect 3017 7884 3155 7893
rect 3017 7864 3126 7884
rect 3146 7864 3155 7884
rect 3017 7857 3155 7864
rect 3213 7884 3361 7893
rect 3213 7864 3222 7884
rect 3242 7864 3332 7884
rect 3352 7864 3361 7884
rect 3017 7855 3113 7857
rect 3213 7854 3361 7864
rect 3420 7884 3457 7894
rect 3532 7893 3569 7894
rect 3513 7891 3569 7893
rect 3420 7864 3428 7884
rect 3448 7864 3457 7884
rect 3269 7853 3305 7854
rect 3117 7794 3154 7795
rect 3420 7794 3457 7864
rect 3482 7884 3569 7891
rect 3482 7881 3540 7884
rect 3482 7861 3487 7881
rect 3508 7864 3540 7881
rect 3560 7864 3569 7884
rect 3508 7861 3569 7864
rect 3482 7854 3569 7861
rect 3628 7884 3665 7894
rect 3628 7864 3636 7884
rect 3656 7864 3665 7884
rect 3482 7853 3513 7854
rect 3116 7793 3457 7794
rect 3041 7788 3457 7793
rect 3041 7768 3044 7788
rect 3064 7768 3457 7788
rect 3628 7793 3665 7864
rect 3695 7893 3726 7946
rect 4452 7937 5085 7946
rect 5388 7965 5399 7983
rect 5417 7965 5427 7983
rect 5734 7981 5765 8034
rect 5795 8063 5832 8134
rect 6003 8139 6396 8159
rect 6416 8139 6419 8159
rect 6003 8134 6419 8139
rect 6003 8133 6344 8134
rect 5947 8073 5978 8074
rect 5795 8043 5804 8063
rect 5824 8043 5832 8063
rect 5795 8033 5832 8043
rect 5891 8066 5978 8073
rect 5891 8063 5952 8066
rect 5891 8043 5900 8063
rect 5920 8046 5952 8063
rect 5973 8046 5978 8066
rect 5920 8043 5978 8046
rect 5891 8036 5978 8043
rect 6003 8063 6040 8133
rect 6306 8132 6343 8133
rect 9312 8106 9339 8284
rect 9379 8246 9443 8258
rect 9719 8254 9756 8286
rect 9927 8285 10176 8307
rect 9927 8254 9964 8285
rect 10140 8283 10176 8285
rect 10140 8254 10177 8283
rect 9379 8245 9414 8246
rect 9356 8240 9414 8245
rect 9356 8220 9359 8240
rect 9379 8226 9414 8240
rect 9434 8226 9443 8246
rect 9379 8218 9443 8226
rect 9405 8217 9443 8218
rect 9406 8216 9443 8217
rect 9509 8250 9545 8251
rect 9617 8250 9653 8251
rect 9509 8244 9653 8250
rect 9509 8242 9575 8244
rect 9509 8222 9517 8242
rect 9537 8223 9575 8242
rect 9597 8242 9653 8244
rect 9597 8223 9625 8242
rect 9537 8222 9625 8223
rect 9645 8222 9653 8242
rect 9509 8216 9653 8222
rect 9719 8246 9757 8254
rect 9825 8250 9861 8251
rect 9719 8226 9728 8246
rect 9748 8226 9757 8246
rect 9719 8217 9757 8226
rect 9776 8243 9861 8250
rect 9776 8223 9783 8243
rect 9804 8242 9861 8243
rect 9804 8223 9833 8242
rect 9776 8222 9833 8223
rect 9853 8222 9861 8242
rect 9719 8216 9756 8217
rect 9776 8216 9861 8222
rect 9927 8246 9965 8254
rect 10038 8250 10074 8251
rect 9927 8226 9936 8246
rect 9956 8226 9965 8246
rect 9927 8217 9965 8226
rect 9989 8242 10074 8250
rect 9989 8222 10046 8242
rect 10066 8222 10074 8242
rect 9927 8216 9964 8217
rect 9989 8216 10074 8222
rect 10140 8246 10178 8254
rect 10140 8226 10149 8246
rect 10169 8226 10178 8246
rect 10140 8217 10178 8226
rect 10319 8253 10355 8329
rect 10769 8325 10806 8334
rect 10769 8307 10779 8325
rect 10797 8307 10806 8325
rect 10769 8297 10806 8307
rect 14692 8341 14860 8342
rect 15111 8341 15135 8358
rect 15699 8350 16095 8358
rect 20980 8355 21018 8361
rect 14692 8315 15136 8341
rect 14692 8313 14860 8315
rect 10319 8243 10356 8253
rect 10319 8225 10329 8243
rect 10347 8225 10356 8243
rect 10772 8233 10809 8235
rect 10772 8232 11420 8233
rect 10140 8216 10177 8217
rect 10319 8216 10356 8225
rect 10771 8226 11420 8232
rect 9563 8195 9599 8216
rect 9989 8195 10020 8216
rect 10771 8208 10781 8226
rect 10799 8212 11420 8226
rect 10799 8208 10809 8212
rect 11250 8211 11420 8212
rect 10771 8198 10809 8208
rect 9396 8191 9496 8195
rect 9396 8187 9458 8191
rect 9396 8161 9403 8187
rect 9429 8165 9458 8187
rect 9484 8165 9496 8191
rect 9429 8161 9496 8165
rect 9396 8158 9496 8161
rect 9564 8158 9599 8195
rect 9661 8192 10020 8195
rect 9661 8187 9883 8192
rect 9661 8163 9674 8187
rect 9698 8168 9883 8187
rect 9907 8168 10020 8192
rect 9698 8163 10020 8168
rect 9661 8159 10020 8163
rect 10087 8187 10236 8195
rect 10087 8167 10098 8187
rect 10118 8167 10236 8187
rect 10087 8160 10236 8167
rect 10087 8159 10128 8160
rect 9411 8106 9448 8107
rect 9507 8106 9544 8107
rect 9563 8106 9599 8158
rect 9618 8106 9655 8107
rect 9311 8097 9449 8106
rect 8247 8079 8278 8082
rect 6155 8073 6191 8074
rect 6003 8043 6012 8063
rect 6032 8043 6040 8063
rect 5891 8034 5947 8036
rect 5891 8033 5928 8034
rect 6003 8033 6040 8043
rect 6099 8063 6247 8073
rect 6347 8070 6443 8072
rect 6099 8043 6108 8063
rect 6128 8043 6218 8063
rect 6238 8043 6247 8063
rect 6099 8034 6247 8043
rect 6305 8063 6443 8070
rect 6305 8043 6314 8063
rect 6334 8043 6443 8063
rect 6305 8034 6443 8043
rect 8247 8053 8254 8079
rect 8273 8053 8278 8079
rect 6099 8033 6136 8034
rect 6155 7982 6191 8034
rect 6210 8033 6247 8034
rect 6306 8033 6343 8034
rect 5626 7980 5667 7981
rect 4452 7930 5084 7937
rect 4452 7928 4514 7930
rect 4030 7918 4198 7919
rect 4452 7918 4474 7928
rect 3745 7893 3782 7894
rect 3695 7884 3782 7893
rect 3695 7864 3753 7884
rect 3773 7864 3782 7884
rect 3695 7854 3782 7864
rect 3841 7884 3878 7894
rect 3841 7864 3849 7884
rect 3869 7864 3878 7884
rect 3695 7853 3726 7854
rect 3841 7793 3878 7864
rect 3628 7769 3878 7793
rect 4030 7892 4474 7918
rect 4030 7890 4198 7892
rect 4030 7712 4057 7890
rect 4097 7852 4161 7864
rect 4437 7860 4474 7892
rect 4645 7891 4894 7913
rect 4645 7860 4682 7891
rect 4858 7889 4894 7891
rect 4858 7860 4895 7889
rect 4097 7851 4132 7852
rect 4074 7846 4132 7851
rect 4074 7826 4077 7846
rect 4097 7832 4132 7846
rect 4152 7832 4161 7852
rect 4097 7824 4161 7832
rect 4123 7823 4161 7824
rect 4124 7822 4161 7823
rect 4227 7856 4263 7857
rect 4335 7856 4371 7857
rect 4227 7848 4371 7856
rect 4227 7828 4235 7848
rect 4255 7828 4284 7848
rect 4227 7827 4284 7828
rect 4306 7828 4343 7848
rect 4363 7828 4371 7848
rect 4306 7827 4371 7828
rect 4227 7822 4371 7827
rect 4437 7852 4475 7860
rect 4543 7856 4579 7857
rect 4437 7832 4446 7852
rect 4466 7832 4475 7852
rect 4437 7823 4475 7832
rect 4494 7849 4579 7856
rect 4494 7829 4501 7849
rect 4522 7848 4579 7849
rect 4522 7829 4551 7848
rect 4494 7828 4551 7829
rect 4571 7828 4579 7848
rect 4437 7822 4474 7823
rect 4494 7822 4579 7828
rect 4645 7852 4683 7860
rect 4756 7856 4792 7857
rect 4645 7832 4654 7852
rect 4674 7832 4683 7852
rect 4645 7823 4683 7832
rect 4707 7848 4792 7856
rect 4707 7828 4764 7848
rect 4784 7828 4792 7848
rect 4645 7822 4682 7823
rect 4707 7822 4792 7828
rect 4858 7852 4896 7860
rect 4858 7832 4867 7852
rect 4887 7832 4896 7852
rect 4858 7823 4896 7832
rect 4858 7822 4895 7823
rect 4281 7801 4317 7822
rect 4707 7801 4738 7822
rect 4114 7797 4214 7801
rect 4114 7793 4176 7797
rect 4114 7767 4121 7793
rect 4147 7771 4176 7793
rect 4202 7771 4214 7797
rect 4147 7767 4214 7771
rect 4114 7764 4214 7767
rect 4282 7764 4317 7801
rect 4379 7798 4738 7801
rect 4379 7793 4601 7798
rect 4379 7769 4392 7793
rect 4416 7774 4601 7793
rect 4625 7774 4738 7798
rect 4416 7769 4738 7774
rect 4379 7765 4738 7769
rect 4805 7793 4954 7801
rect 4805 7773 4816 7793
rect 4836 7773 4954 7793
rect 4805 7766 4954 7773
rect 5045 7781 5084 7930
rect 5388 7816 5427 7965
rect 5518 7973 5667 7980
rect 5518 7953 5636 7973
rect 5656 7953 5667 7973
rect 5518 7945 5667 7953
rect 5734 7977 6093 7981
rect 5734 7972 6056 7977
rect 5734 7948 5847 7972
rect 5871 7953 6056 7972
rect 6080 7953 6093 7977
rect 5871 7948 6093 7953
rect 5734 7945 6093 7948
rect 6155 7945 6190 7982
rect 6258 7979 6358 7982
rect 6258 7975 6325 7979
rect 6258 7949 6270 7975
rect 6296 7953 6325 7975
rect 6351 7953 6358 7979
rect 6296 7949 6358 7953
rect 6258 7945 6358 7949
rect 5734 7924 5765 7945
rect 6155 7924 6191 7945
rect 5577 7923 5614 7924
rect 5576 7914 5614 7923
rect 5576 7894 5585 7914
rect 5605 7894 5614 7914
rect 5576 7886 5614 7894
rect 5680 7918 5765 7924
rect 5790 7923 5827 7924
rect 5680 7898 5688 7918
rect 5708 7898 5765 7918
rect 5680 7890 5765 7898
rect 5789 7914 5827 7923
rect 5789 7894 5798 7914
rect 5818 7894 5827 7914
rect 5680 7889 5716 7890
rect 5789 7886 5827 7894
rect 5893 7918 5978 7924
rect 5998 7923 6035 7924
rect 5893 7898 5901 7918
rect 5921 7917 5978 7918
rect 5921 7898 5950 7917
rect 5893 7897 5950 7898
rect 5971 7897 5978 7917
rect 5893 7890 5978 7897
rect 5997 7914 6035 7923
rect 5997 7894 6006 7914
rect 6026 7894 6035 7914
rect 5893 7889 5929 7890
rect 5997 7886 6035 7894
rect 6101 7919 6245 7924
rect 6101 7918 6166 7919
rect 6101 7898 6109 7918
rect 6129 7898 6166 7918
rect 6188 7918 6245 7919
rect 6188 7898 6217 7918
rect 6237 7898 6245 7918
rect 6101 7890 6245 7898
rect 6101 7889 6137 7890
rect 6209 7889 6245 7890
rect 6311 7923 6348 7924
rect 6311 7922 6349 7923
rect 6311 7914 6375 7922
rect 6311 7894 6320 7914
rect 6340 7900 6375 7914
rect 6395 7900 6398 7920
rect 6340 7895 6398 7900
rect 6340 7894 6375 7895
rect 5577 7857 5614 7886
rect 5578 7855 5614 7857
rect 5790 7855 5827 7886
rect 5578 7833 5827 7855
rect 5998 7854 6035 7886
rect 6311 7882 6375 7894
rect 6415 7856 6442 8034
rect 6274 7854 6442 7856
rect 5998 7828 6442 7854
rect 6594 7953 6844 7977
rect 6594 7882 6631 7953
rect 6746 7892 6777 7893
rect 6594 7862 6603 7882
rect 6623 7862 6631 7882
rect 6594 7852 6631 7862
rect 6690 7882 6777 7892
rect 6690 7862 6699 7882
rect 6719 7862 6777 7882
rect 6690 7853 6777 7862
rect 6690 7852 6727 7853
rect 5998 7818 6020 7828
rect 6274 7827 6442 7828
rect 5958 7816 6020 7818
rect 5388 7809 6020 7816
rect 4805 7765 4846 7766
rect 4129 7712 4166 7713
rect 4225 7712 4262 7713
rect 4281 7712 4317 7764
rect 4336 7712 4373 7713
rect 4029 7703 4167 7712
rect 4029 7683 4138 7703
rect 4158 7683 4167 7703
rect 2966 7679 3136 7680
rect 2966 7664 3412 7679
rect 4029 7676 4167 7683
rect 4225 7703 4373 7712
rect 4225 7683 4234 7703
rect 4254 7683 4344 7703
rect 4364 7683 4373 7703
rect 4029 7674 4125 7676
rect 2873 7653 2905 7658
rect 1023 7640 1161 7649
rect 817 7639 854 7640
rect 873 7588 909 7640
rect 928 7639 965 7640
rect 1024 7639 1061 7640
rect 344 7586 385 7587
rect 236 7579 385 7586
rect 236 7559 354 7579
rect 374 7559 385 7579
rect 236 7551 385 7559
rect 452 7583 811 7587
rect 452 7578 774 7583
rect 452 7554 565 7578
rect 589 7559 774 7578
rect 798 7559 811 7583
rect 589 7554 811 7559
rect 452 7551 811 7554
rect 873 7551 908 7588
rect 976 7585 1076 7588
rect 976 7581 1043 7585
rect 976 7555 988 7581
rect 1014 7559 1043 7581
rect 1069 7559 1076 7585
rect 1014 7555 1076 7559
rect 976 7551 1076 7555
rect 452 7530 483 7551
rect 873 7530 909 7551
rect 116 7521 153 7530
rect 295 7529 332 7530
rect 116 7503 125 7521
rect 143 7503 153 7521
rect 116 7493 153 7503
rect 117 7458 153 7493
rect 294 7520 332 7529
rect 294 7500 303 7520
rect 323 7500 332 7520
rect 294 7492 332 7500
rect 398 7524 483 7530
rect 508 7529 545 7530
rect 398 7504 406 7524
rect 426 7504 483 7524
rect 398 7496 483 7504
rect 507 7520 545 7529
rect 507 7500 516 7520
rect 536 7500 545 7520
rect 398 7495 434 7496
rect 507 7492 545 7500
rect 611 7524 696 7530
rect 716 7529 753 7530
rect 611 7504 619 7524
rect 639 7523 696 7524
rect 639 7504 668 7523
rect 611 7503 668 7504
rect 689 7503 696 7523
rect 611 7496 696 7503
rect 715 7520 753 7529
rect 715 7500 724 7520
rect 744 7500 753 7520
rect 611 7495 647 7496
rect 715 7492 753 7500
rect 819 7524 963 7530
rect 819 7504 827 7524
rect 847 7523 935 7524
rect 847 7504 875 7523
rect 819 7502 875 7504
rect 897 7504 935 7523
rect 955 7504 963 7524
rect 897 7502 963 7504
rect 819 7496 963 7502
rect 819 7495 855 7496
rect 927 7495 963 7496
rect 1029 7529 1066 7530
rect 1029 7528 1067 7529
rect 1029 7520 1093 7528
rect 1029 7500 1038 7520
rect 1058 7506 1093 7520
rect 1113 7506 1116 7526
rect 1058 7501 1116 7506
rect 1058 7500 1093 7501
rect 295 7463 332 7492
rect 115 7417 153 7458
rect 296 7461 332 7463
rect 508 7461 545 7492
rect 296 7439 545 7461
rect 716 7460 753 7492
rect 1029 7488 1093 7500
rect 1133 7462 1160 7640
rect 992 7460 1160 7462
rect 716 7434 1160 7460
rect 717 7417 741 7434
rect 992 7433 1160 7434
rect 115 7399 742 7417
rect 1368 7413 1618 7437
rect 115 7393 153 7399
rect 115 7369 152 7393
rect 115 7345 150 7369
rect 113 7336 150 7345
rect 113 7318 123 7336
rect 141 7318 150 7336
rect 113 7308 150 7318
rect 1368 7342 1405 7413
rect 1520 7352 1551 7353
rect 1368 7322 1377 7342
rect 1397 7322 1405 7342
rect 1368 7312 1405 7322
rect 1464 7342 1551 7352
rect 1464 7322 1473 7342
rect 1493 7322 1551 7342
rect 1464 7313 1551 7322
rect 1464 7312 1501 7313
rect 1520 7260 1551 7313
rect 1581 7342 1618 7413
rect 1789 7418 2182 7438
rect 2202 7418 2205 7438
rect 1789 7413 2205 7418
rect 1789 7412 2130 7413
rect 1733 7352 1764 7353
rect 1581 7322 1590 7342
rect 1610 7322 1618 7342
rect 1581 7312 1618 7322
rect 1677 7345 1764 7352
rect 1677 7342 1738 7345
rect 1677 7322 1686 7342
rect 1706 7325 1738 7342
rect 1759 7325 1764 7345
rect 1706 7322 1764 7325
rect 1677 7315 1764 7322
rect 1789 7342 1826 7412
rect 2092 7411 2129 7412
rect 1941 7352 1977 7353
rect 1789 7322 1798 7342
rect 1818 7322 1826 7342
rect 1677 7313 1733 7315
rect 1677 7312 1714 7313
rect 1789 7312 1826 7322
rect 1885 7342 2033 7352
rect 2133 7349 2229 7351
rect 1885 7322 1894 7342
rect 1914 7322 2004 7342
rect 2024 7322 2033 7342
rect 1885 7313 2033 7322
rect 2091 7342 2229 7349
rect 2091 7322 2100 7342
rect 2120 7322 2229 7342
rect 2091 7313 2229 7322
rect 1885 7312 1922 7313
rect 1941 7261 1977 7313
rect 1996 7312 2033 7313
rect 2092 7312 2129 7313
rect 1412 7259 1453 7260
rect 1304 7252 1453 7259
rect 116 7244 153 7246
rect 116 7243 764 7244
rect 115 7237 764 7243
rect 115 7219 125 7237
rect 143 7223 764 7237
rect 1304 7232 1422 7252
rect 1442 7232 1453 7252
rect 1304 7224 1453 7232
rect 1520 7256 1879 7260
rect 1520 7251 1842 7256
rect 1520 7227 1633 7251
rect 1657 7232 1842 7251
rect 1866 7232 1879 7256
rect 1657 7227 1879 7232
rect 1520 7224 1879 7227
rect 1941 7224 1976 7261
rect 2044 7258 2144 7261
rect 2044 7254 2111 7258
rect 2044 7228 2056 7254
rect 2082 7232 2111 7254
rect 2137 7232 2144 7258
rect 2082 7228 2144 7232
rect 2044 7224 2144 7228
rect 143 7219 153 7223
rect 594 7222 764 7223
rect 115 7209 153 7219
rect 115 7131 150 7209
rect 727 7199 764 7222
rect 1520 7203 1551 7224
rect 1941 7203 1977 7224
rect 1363 7202 1400 7203
rect 111 7122 150 7131
rect 111 7104 121 7122
rect 139 7104 150 7122
rect 111 7098 150 7104
rect 306 7174 556 7198
rect 306 7103 343 7174
rect 458 7113 489 7114
rect 111 7094 148 7098
rect 306 7083 315 7103
rect 335 7083 343 7103
rect 306 7073 343 7083
rect 402 7103 489 7113
rect 402 7083 411 7103
rect 431 7083 489 7103
rect 402 7074 489 7083
rect 402 7073 439 7074
rect 114 7023 151 7032
rect 112 7005 123 7023
rect 141 7005 151 7023
rect 458 7021 489 7074
rect 519 7103 556 7174
rect 727 7179 1120 7199
rect 1140 7179 1143 7199
rect 727 7174 1143 7179
rect 1362 7193 1400 7202
rect 727 7173 1068 7174
rect 1362 7173 1371 7193
rect 1391 7173 1400 7193
rect 671 7113 702 7114
rect 519 7083 528 7103
rect 548 7083 556 7103
rect 519 7073 556 7083
rect 615 7106 702 7113
rect 615 7103 676 7106
rect 615 7083 624 7103
rect 644 7086 676 7103
rect 697 7086 702 7106
rect 644 7083 702 7086
rect 615 7076 702 7083
rect 727 7103 764 7173
rect 1030 7172 1067 7173
rect 1362 7165 1400 7173
rect 1466 7197 1551 7203
rect 1576 7202 1613 7203
rect 1466 7177 1474 7197
rect 1494 7177 1551 7197
rect 1466 7169 1551 7177
rect 1575 7193 1613 7202
rect 1575 7173 1584 7193
rect 1604 7173 1613 7193
rect 1466 7168 1502 7169
rect 1575 7165 1613 7173
rect 1679 7197 1764 7203
rect 1784 7202 1821 7203
rect 1679 7177 1687 7197
rect 1707 7196 1764 7197
rect 1707 7177 1736 7196
rect 1679 7176 1736 7177
rect 1757 7176 1764 7196
rect 1679 7169 1764 7176
rect 1783 7193 1821 7202
rect 1783 7173 1792 7193
rect 1812 7173 1821 7193
rect 1679 7168 1715 7169
rect 1783 7165 1821 7173
rect 1887 7197 2031 7203
rect 1887 7177 1895 7197
rect 1915 7195 2003 7197
rect 1915 7178 1951 7195
rect 1975 7178 2003 7195
rect 1915 7177 2003 7178
rect 2023 7177 2031 7197
rect 1887 7169 2031 7177
rect 1887 7168 1923 7169
rect 1995 7168 2031 7169
rect 2097 7202 2134 7203
rect 2097 7201 2135 7202
rect 2097 7193 2161 7201
rect 2097 7173 2106 7193
rect 2126 7179 2161 7193
rect 2181 7179 2184 7199
rect 2126 7174 2184 7179
rect 2126 7173 2161 7174
rect 1363 7136 1400 7165
rect 1364 7134 1400 7136
rect 1576 7134 1613 7165
rect 879 7113 915 7114
rect 727 7083 736 7103
rect 756 7083 764 7103
rect 615 7074 671 7076
rect 615 7073 652 7074
rect 727 7073 764 7083
rect 823 7103 971 7113
rect 1364 7112 1613 7134
rect 1784 7133 1821 7165
rect 2097 7161 2161 7173
rect 2201 7135 2228 7313
rect 2060 7133 2228 7135
rect 1784 7122 2228 7133
rect 1071 7110 1167 7112
rect 823 7083 832 7103
rect 852 7083 942 7103
rect 962 7083 971 7103
rect 823 7074 971 7083
rect 1029 7103 1167 7110
rect 1784 7107 2230 7122
rect 2060 7106 2230 7107
rect 1029 7083 1038 7103
rect 1058 7083 1167 7103
rect 1029 7074 1167 7083
rect 823 7073 860 7074
rect 879 7022 915 7074
rect 934 7073 971 7074
rect 1030 7073 1067 7074
rect 350 7020 391 7021
rect 112 6856 151 7005
rect 242 7013 391 7020
rect 242 6993 360 7013
rect 380 6993 391 7013
rect 242 6985 391 6993
rect 458 7017 817 7021
rect 458 7012 780 7017
rect 458 6988 571 7012
rect 595 6993 780 7012
rect 804 6993 817 7017
rect 595 6988 817 6993
rect 458 6985 817 6988
rect 879 6985 914 7022
rect 982 7019 1082 7022
rect 982 7015 1049 7019
rect 982 6989 994 7015
rect 1020 6993 1049 7015
rect 1075 6993 1082 7019
rect 1020 6989 1082 6993
rect 982 6985 1082 6989
rect 458 6964 489 6985
rect 879 6964 915 6985
rect 301 6963 338 6964
rect 300 6954 338 6963
rect 300 6934 309 6954
rect 329 6934 338 6954
rect 300 6926 338 6934
rect 404 6958 489 6964
rect 514 6963 551 6964
rect 404 6938 412 6958
rect 432 6938 489 6958
rect 404 6930 489 6938
rect 513 6954 551 6963
rect 513 6934 522 6954
rect 542 6934 551 6954
rect 404 6929 440 6930
rect 513 6926 551 6934
rect 617 6958 702 6964
rect 722 6963 759 6964
rect 617 6938 625 6958
rect 645 6957 702 6958
rect 645 6938 674 6957
rect 617 6937 674 6938
rect 695 6937 702 6957
rect 617 6930 702 6937
rect 721 6954 759 6963
rect 721 6934 730 6954
rect 750 6934 759 6954
rect 617 6929 653 6930
rect 721 6926 759 6934
rect 825 6959 969 6964
rect 825 6958 890 6959
rect 825 6938 833 6958
rect 853 6938 890 6958
rect 912 6958 969 6959
rect 912 6938 941 6958
rect 961 6938 969 6958
rect 825 6930 969 6938
rect 825 6929 861 6930
rect 933 6929 969 6930
rect 1035 6963 1072 6964
rect 1035 6962 1073 6963
rect 1035 6954 1099 6962
rect 1035 6934 1044 6954
rect 1064 6940 1099 6954
rect 1119 6940 1122 6960
rect 1064 6935 1122 6940
rect 1064 6934 1099 6935
rect 301 6897 338 6926
rect 302 6895 338 6897
rect 514 6895 551 6926
rect 302 6873 551 6895
rect 722 6894 759 6926
rect 1035 6922 1099 6934
rect 1139 6896 1166 7074
rect 998 6894 1166 6896
rect 722 6868 1166 6894
rect 1318 6993 1568 7017
rect 1318 6922 1355 6993
rect 1470 6932 1501 6933
rect 1318 6902 1327 6922
rect 1347 6902 1355 6922
rect 1318 6892 1355 6902
rect 1414 6922 1501 6932
rect 1414 6902 1423 6922
rect 1443 6902 1501 6922
rect 1414 6893 1501 6902
rect 1414 6892 1451 6893
rect 722 6858 744 6868
rect 998 6867 1166 6868
rect 682 6856 744 6858
rect 112 6849 744 6856
rect 111 6840 744 6849
rect 1470 6840 1501 6893
rect 1531 6922 1568 6993
rect 1739 6998 2132 7018
rect 2152 6998 2155 7018
rect 1739 6993 2155 6998
rect 1739 6992 2080 6993
rect 1683 6932 1714 6933
rect 1531 6902 1540 6922
rect 1560 6902 1568 6922
rect 1531 6892 1568 6902
rect 1627 6925 1714 6932
rect 1627 6922 1688 6925
rect 1627 6902 1636 6922
rect 1656 6905 1688 6922
rect 1709 6905 1714 6925
rect 1656 6902 1714 6905
rect 1627 6895 1714 6902
rect 1739 6922 1776 6992
rect 2042 6991 2079 6992
rect 1891 6932 1927 6933
rect 1739 6902 1748 6922
rect 1768 6902 1776 6922
rect 1627 6893 1683 6895
rect 1627 6892 1664 6893
rect 1739 6892 1776 6902
rect 1835 6922 1983 6932
rect 2083 6929 2179 6931
rect 1835 6902 1844 6922
rect 1864 6902 1954 6922
rect 1974 6902 1983 6922
rect 1835 6893 1983 6902
rect 2041 6922 2179 6929
rect 2041 6902 2050 6922
rect 2070 6902 2179 6922
rect 2041 6893 2179 6902
rect 1835 6892 1872 6893
rect 1891 6841 1927 6893
rect 1946 6892 1983 6893
rect 2042 6892 2079 6893
rect 111 6822 121 6840
rect 139 6839 744 6840
rect 1362 6839 1403 6840
rect 139 6834 160 6839
rect 139 6822 151 6834
rect 1254 6832 1403 6839
rect 111 6814 151 6822
rect 194 6821 220 6822
rect 111 6812 148 6814
rect 194 6803 748 6821
rect 1254 6812 1372 6832
rect 1392 6812 1403 6832
rect 1254 6804 1403 6812
rect 1470 6836 1829 6840
rect 1470 6831 1792 6836
rect 1470 6807 1583 6831
rect 1607 6812 1792 6831
rect 1816 6812 1829 6836
rect 1607 6807 1829 6812
rect 1470 6804 1829 6807
rect 1891 6804 1926 6841
rect 1994 6838 2094 6841
rect 1994 6834 2061 6838
rect 1994 6808 2006 6834
rect 2032 6812 2061 6834
rect 2087 6812 2094 6838
rect 2032 6808 2094 6812
rect 1994 6804 2094 6808
rect 114 6744 151 6750
rect 194 6744 220 6803
rect 727 6784 748 6803
rect 114 6741 220 6744
rect 114 6723 123 6741
rect 141 6727 220 6741
rect 305 6759 555 6783
rect 141 6725 217 6727
rect 141 6723 151 6725
rect 114 6713 151 6723
rect 119 6648 150 6713
rect 305 6688 342 6759
rect 457 6698 488 6699
rect 305 6668 314 6688
rect 334 6668 342 6688
rect 305 6658 342 6668
rect 401 6688 488 6698
rect 401 6668 410 6688
rect 430 6668 488 6688
rect 401 6659 488 6668
rect 401 6658 438 6659
rect 118 6639 155 6648
rect 118 6621 128 6639
rect 146 6621 155 6639
rect 118 6611 155 6621
rect 457 6606 488 6659
rect 518 6688 555 6759
rect 726 6764 1119 6784
rect 1139 6764 1142 6784
rect 1470 6783 1501 6804
rect 1891 6783 1927 6804
rect 1313 6782 1350 6783
rect 726 6759 1142 6764
rect 1312 6773 1350 6782
rect 726 6758 1067 6759
rect 670 6698 701 6699
rect 518 6668 527 6688
rect 547 6668 555 6688
rect 518 6658 555 6668
rect 614 6691 701 6698
rect 614 6688 675 6691
rect 614 6668 623 6688
rect 643 6671 675 6688
rect 696 6671 701 6691
rect 643 6668 701 6671
rect 614 6661 701 6668
rect 726 6688 763 6758
rect 1029 6757 1066 6758
rect 1312 6753 1321 6773
rect 1341 6753 1350 6773
rect 1312 6745 1350 6753
rect 1416 6777 1501 6783
rect 1526 6782 1563 6783
rect 1416 6757 1424 6777
rect 1444 6757 1501 6777
rect 1416 6749 1501 6757
rect 1525 6773 1563 6782
rect 1525 6753 1534 6773
rect 1554 6753 1563 6773
rect 1416 6748 1452 6749
rect 1525 6745 1563 6753
rect 1629 6777 1714 6783
rect 1734 6782 1771 6783
rect 1629 6757 1637 6777
rect 1657 6776 1714 6777
rect 1657 6757 1686 6776
rect 1629 6756 1686 6757
rect 1707 6756 1714 6776
rect 1629 6749 1714 6756
rect 1733 6773 1771 6782
rect 1733 6753 1742 6773
rect 1762 6753 1771 6773
rect 1629 6748 1665 6749
rect 1733 6745 1771 6753
rect 1837 6778 1981 6783
rect 1837 6777 1896 6778
rect 1837 6757 1845 6777
rect 1865 6758 1896 6777
rect 1920 6777 1981 6778
rect 1920 6758 1953 6777
rect 1865 6757 1953 6758
rect 1973 6757 1981 6777
rect 1837 6749 1981 6757
rect 1837 6748 1873 6749
rect 1945 6748 1981 6749
rect 2047 6782 2084 6783
rect 2047 6781 2085 6782
rect 2047 6773 2111 6781
rect 2047 6753 2056 6773
rect 2076 6759 2111 6773
rect 2131 6759 2134 6779
rect 2076 6754 2134 6759
rect 2076 6753 2111 6754
rect 1313 6716 1350 6745
rect 1314 6714 1350 6716
rect 1526 6714 1563 6745
rect 878 6698 914 6699
rect 726 6668 735 6688
rect 755 6668 763 6688
rect 614 6659 670 6661
rect 614 6658 651 6659
rect 726 6658 763 6668
rect 822 6688 970 6698
rect 1070 6695 1166 6697
rect 822 6668 831 6688
rect 851 6668 941 6688
rect 961 6668 970 6688
rect 822 6659 970 6668
rect 1028 6688 1166 6695
rect 1314 6692 1563 6714
rect 1734 6713 1771 6745
rect 2047 6741 2111 6753
rect 2151 6715 2178 6893
rect 2010 6713 2178 6715
rect 1734 6709 2178 6713
rect 1028 6668 1037 6688
rect 1057 6668 1166 6688
rect 1734 6690 1783 6709
rect 1803 6690 2178 6709
rect 1734 6687 2178 6690
rect 2010 6686 2178 6687
rect 2199 6712 2230 7106
rect 2199 6686 2204 6712
rect 2223 6686 2230 6712
rect 2199 6683 2230 6686
rect 1028 6659 1166 6668
rect 822 6658 859 6659
rect 878 6607 914 6659
rect 933 6658 970 6659
rect 1029 6658 1066 6659
rect 349 6605 390 6606
rect 241 6598 390 6605
rect 241 6578 359 6598
rect 379 6578 390 6598
rect 241 6570 390 6578
rect 457 6602 816 6606
rect 457 6597 779 6602
rect 457 6573 570 6597
rect 594 6578 779 6597
rect 803 6578 816 6602
rect 594 6573 816 6578
rect 457 6570 816 6573
rect 878 6570 913 6607
rect 981 6604 1081 6607
rect 981 6600 1048 6604
rect 981 6574 993 6600
rect 1019 6578 1048 6600
rect 1074 6578 1081 6604
rect 1019 6574 1081 6578
rect 981 6570 1081 6574
rect 457 6549 488 6570
rect 878 6549 914 6570
rect 121 6540 158 6549
rect 300 6548 337 6549
rect 121 6522 130 6540
rect 148 6522 158 6540
rect 121 6512 158 6522
rect 122 6477 158 6512
rect 299 6539 337 6548
rect 299 6519 308 6539
rect 328 6519 337 6539
rect 299 6511 337 6519
rect 403 6543 488 6549
rect 513 6548 550 6549
rect 403 6523 411 6543
rect 431 6523 488 6543
rect 403 6515 488 6523
rect 512 6539 550 6548
rect 512 6519 521 6539
rect 541 6519 550 6539
rect 403 6514 439 6515
rect 512 6511 550 6519
rect 616 6543 701 6549
rect 721 6548 758 6549
rect 616 6523 624 6543
rect 644 6542 701 6543
rect 644 6523 673 6542
rect 616 6522 673 6523
rect 694 6522 701 6542
rect 616 6515 701 6522
rect 720 6539 758 6548
rect 720 6519 729 6539
rect 749 6519 758 6539
rect 616 6514 652 6515
rect 720 6511 758 6519
rect 824 6543 968 6549
rect 824 6523 832 6543
rect 852 6542 940 6543
rect 852 6523 880 6542
rect 824 6521 880 6523
rect 902 6523 940 6542
rect 960 6523 968 6543
rect 902 6521 968 6523
rect 824 6515 968 6521
rect 824 6514 860 6515
rect 932 6514 968 6515
rect 1034 6548 1071 6549
rect 1034 6547 1072 6548
rect 1034 6539 1098 6547
rect 1034 6519 1043 6539
rect 1063 6525 1098 6539
rect 1118 6525 1121 6545
rect 1063 6520 1121 6525
rect 1063 6519 1098 6520
rect 300 6482 337 6511
rect 120 6436 158 6477
rect 301 6480 337 6482
rect 513 6480 550 6511
rect 301 6458 550 6480
rect 721 6479 758 6511
rect 1034 6507 1098 6519
rect 1138 6481 1165 6659
rect 2749 6648 2786 6659
rect 2875 6652 2905 7653
rect 2968 7653 3412 7664
rect 2968 7651 3136 7653
rect 2968 7473 2995 7651
rect 3035 7613 3099 7625
rect 3375 7621 3412 7653
rect 3583 7652 3832 7674
rect 4225 7673 4373 7683
rect 4432 7703 4469 7713
rect 4544 7712 4581 7713
rect 4525 7710 4581 7712
rect 4432 7683 4440 7703
rect 4460 7683 4469 7703
rect 4281 7672 4317 7673
rect 3583 7621 3620 7652
rect 3796 7650 3832 7652
rect 3796 7621 3833 7650
rect 3035 7612 3070 7613
rect 3012 7607 3070 7612
rect 3012 7587 3015 7607
rect 3035 7593 3070 7607
rect 3090 7593 3099 7613
rect 3035 7585 3099 7593
rect 3061 7584 3099 7585
rect 3062 7583 3099 7584
rect 3165 7617 3201 7618
rect 3273 7617 3309 7618
rect 3165 7609 3309 7617
rect 3165 7589 3173 7609
rect 3193 7590 3225 7609
rect 3248 7590 3281 7609
rect 3193 7589 3281 7590
rect 3301 7589 3309 7609
rect 3165 7583 3309 7589
rect 3375 7613 3413 7621
rect 3481 7617 3517 7618
rect 3375 7593 3384 7613
rect 3404 7593 3413 7613
rect 3375 7584 3413 7593
rect 3432 7610 3517 7617
rect 3432 7590 3439 7610
rect 3460 7609 3517 7610
rect 3460 7590 3489 7609
rect 3432 7589 3489 7590
rect 3509 7589 3517 7609
rect 3375 7583 3412 7584
rect 3432 7583 3517 7589
rect 3583 7613 3621 7621
rect 3694 7617 3730 7618
rect 3583 7593 3592 7613
rect 3612 7593 3621 7613
rect 3583 7584 3621 7593
rect 3645 7609 3730 7617
rect 3645 7589 3702 7609
rect 3722 7589 3730 7609
rect 3583 7583 3620 7584
rect 3645 7583 3730 7589
rect 3796 7613 3834 7621
rect 4129 7613 4166 7614
rect 4432 7613 4469 7683
rect 4494 7703 4581 7710
rect 4494 7700 4552 7703
rect 4494 7680 4499 7700
rect 4520 7683 4552 7700
rect 4572 7683 4581 7703
rect 4520 7680 4581 7683
rect 4494 7673 4581 7680
rect 4640 7703 4677 7713
rect 4640 7683 4648 7703
rect 4668 7683 4677 7703
rect 4494 7672 4525 7673
rect 3796 7593 3805 7613
rect 3825 7593 3834 7613
rect 4128 7612 4469 7613
rect 3796 7584 3834 7593
rect 4053 7607 4469 7612
rect 4053 7587 4056 7607
rect 4076 7587 4469 7607
rect 4640 7612 4677 7683
rect 4707 7712 4738 7765
rect 5045 7763 5055 7781
rect 5073 7763 5084 7781
rect 5387 7800 6020 7809
rect 6746 7800 6777 7853
rect 6807 7882 6844 7953
rect 7015 7958 7408 7978
rect 7428 7958 7431 7978
rect 7015 7953 7431 7958
rect 7015 7952 7356 7953
rect 6959 7892 6990 7893
rect 6807 7862 6816 7882
rect 6836 7862 6844 7882
rect 6807 7852 6844 7862
rect 6903 7885 6990 7892
rect 6903 7882 6964 7885
rect 6903 7862 6912 7882
rect 6932 7865 6964 7882
rect 6985 7865 6990 7885
rect 6932 7862 6990 7865
rect 6903 7855 6990 7862
rect 7015 7882 7052 7952
rect 7318 7951 7355 7952
rect 7167 7892 7203 7893
rect 7015 7862 7024 7882
rect 7044 7862 7052 7882
rect 6903 7853 6959 7855
rect 6903 7852 6940 7853
rect 7015 7852 7052 7862
rect 7111 7882 7259 7892
rect 7359 7889 7455 7891
rect 7111 7862 7120 7882
rect 7140 7862 7230 7882
rect 7250 7862 7259 7882
rect 7111 7853 7259 7862
rect 7317 7882 7455 7889
rect 7317 7862 7326 7882
rect 7346 7862 7455 7882
rect 7317 7853 7455 7862
rect 7111 7852 7148 7853
rect 7167 7801 7203 7853
rect 7222 7852 7259 7853
rect 7318 7852 7355 7853
rect 5387 7782 5397 7800
rect 5415 7799 6020 7800
rect 6638 7799 6679 7800
rect 5415 7794 5436 7799
rect 5415 7782 5427 7794
rect 6530 7792 6679 7799
rect 5387 7774 5427 7782
rect 5470 7781 5496 7782
rect 5387 7772 5424 7774
rect 5470 7763 6024 7781
rect 6530 7772 6648 7792
rect 6668 7772 6679 7792
rect 6530 7764 6679 7772
rect 6746 7796 7105 7800
rect 6746 7791 7068 7796
rect 6746 7767 6859 7791
rect 6883 7772 7068 7791
rect 7092 7772 7105 7796
rect 6883 7767 7105 7772
rect 6746 7764 7105 7767
rect 7167 7764 7202 7801
rect 7270 7798 7370 7801
rect 7270 7794 7337 7798
rect 7270 7768 7282 7794
rect 7308 7772 7337 7794
rect 7363 7772 7370 7798
rect 7308 7768 7370 7772
rect 7270 7764 7370 7768
rect 5045 7754 5082 7763
rect 4757 7712 4794 7713
rect 4707 7703 4794 7712
rect 4707 7683 4765 7703
rect 4785 7683 4794 7703
rect 4707 7673 4794 7683
rect 4853 7703 4890 7713
rect 4853 7683 4861 7703
rect 4881 7683 4890 7703
rect 5390 7704 5427 7710
rect 5470 7704 5496 7763
rect 6003 7744 6024 7763
rect 5390 7701 5496 7704
rect 5048 7688 5085 7692
rect 4707 7672 4738 7673
rect 4853 7612 4890 7683
rect 4640 7588 4890 7612
rect 5046 7682 5085 7688
rect 5046 7664 5057 7682
rect 5075 7664 5085 7682
rect 5390 7683 5399 7701
rect 5417 7687 5496 7701
rect 5581 7719 5831 7743
rect 5417 7685 5493 7687
rect 5417 7683 5427 7685
rect 5390 7673 5427 7683
rect 5046 7655 5085 7664
rect 3796 7583 3833 7584
rect 3219 7562 3255 7583
rect 3645 7562 3676 7583
rect 4432 7564 4469 7587
rect 5046 7577 5081 7655
rect 5395 7608 5426 7673
rect 5581 7648 5618 7719
rect 5733 7658 5764 7659
rect 5581 7628 5590 7648
rect 5610 7628 5618 7648
rect 5581 7618 5618 7628
rect 5677 7648 5764 7658
rect 5677 7628 5686 7648
rect 5706 7628 5764 7648
rect 5677 7619 5764 7628
rect 5677 7618 5714 7619
rect 5043 7567 5081 7577
rect 5394 7599 5431 7608
rect 5394 7581 5404 7599
rect 5422 7581 5431 7599
rect 5394 7571 5431 7581
rect 4432 7563 4602 7564
rect 5043 7563 5053 7567
rect 3052 7558 3152 7562
rect 3052 7554 3114 7558
rect 3052 7528 3059 7554
rect 3085 7532 3114 7554
rect 3140 7532 3152 7558
rect 3085 7528 3152 7532
rect 3052 7525 3152 7528
rect 3220 7525 3255 7562
rect 3317 7559 3676 7562
rect 3317 7554 3539 7559
rect 3317 7530 3330 7554
rect 3354 7535 3539 7554
rect 3563 7535 3676 7559
rect 3354 7530 3676 7535
rect 3317 7526 3676 7530
rect 3743 7554 3892 7562
rect 3743 7534 3754 7554
rect 3774 7534 3892 7554
rect 4432 7549 5053 7563
rect 5071 7549 5081 7567
rect 5733 7566 5764 7619
rect 5794 7648 5831 7719
rect 6002 7724 6395 7744
rect 6415 7724 6418 7744
rect 6746 7743 6777 7764
rect 7167 7743 7203 7764
rect 6589 7742 6626 7743
rect 6002 7719 6418 7724
rect 6588 7733 6626 7742
rect 6002 7718 6343 7719
rect 5946 7658 5977 7659
rect 5794 7628 5803 7648
rect 5823 7628 5831 7648
rect 5794 7618 5831 7628
rect 5890 7651 5977 7658
rect 5890 7648 5951 7651
rect 5890 7628 5899 7648
rect 5919 7631 5951 7648
rect 5972 7631 5977 7651
rect 5919 7628 5977 7631
rect 5890 7621 5977 7628
rect 6002 7648 6039 7718
rect 6305 7717 6342 7718
rect 6588 7713 6597 7733
rect 6617 7713 6626 7733
rect 6588 7705 6626 7713
rect 6692 7737 6777 7743
rect 6802 7742 6839 7743
rect 6692 7717 6700 7737
rect 6720 7717 6777 7737
rect 6692 7709 6777 7717
rect 6801 7733 6839 7742
rect 6801 7713 6810 7733
rect 6830 7713 6839 7733
rect 6692 7708 6728 7709
rect 6801 7705 6839 7713
rect 6905 7737 6990 7743
rect 7010 7742 7047 7743
rect 6905 7717 6913 7737
rect 6933 7736 6990 7737
rect 6933 7717 6962 7736
rect 6905 7716 6962 7717
rect 6983 7716 6990 7736
rect 6905 7709 6990 7716
rect 7009 7733 7047 7742
rect 7009 7713 7018 7733
rect 7038 7713 7047 7733
rect 6905 7708 6941 7709
rect 7009 7705 7047 7713
rect 7113 7737 7257 7743
rect 7113 7717 7121 7737
rect 7141 7717 7173 7737
rect 7197 7717 7229 7737
rect 7249 7717 7257 7737
rect 7113 7709 7257 7717
rect 7113 7708 7149 7709
rect 7221 7708 7257 7709
rect 7323 7742 7360 7743
rect 7323 7741 7361 7742
rect 7323 7733 7387 7741
rect 7323 7713 7332 7733
rect 7352 7719 7387 7733
rect 7407 7719 7410 7739
rect 7352 7714 7410 7719
rect 7352 7713 7387 7714
rect 6589 7676 6626 7705
rect 6590 7674 6626 7676
rect 6802 7674 6839 7705
rect 6154 7658 6190 7659
rect 6002 7628 6011 7648
rect 6031 7628 6039 7648
rect 5890 7619 5946 7621
rect 5890 7618 5927 7619
rect 6002 7618 6039 7628
rect 6098 7648 6246 7658
rect 6346 7655 6442 7657
rect 6098 7628 6107 7648
rect 6127 7628 6217 7648
rect 6237 7628 6246 7648
rect 6098 7619 6246 7628
rect 6304 7648 6442 7655
rect 6590 7652 6839 7674
rect 7010 7673 7047 7705
rect 7323 7701 7387 7713
rect 7427 7675 7454 7853
rect 7286 7673 7454 7675
rect 7010 7669 7454 7673
rect 6304 7628 6313 7648
rect 6333 7628 6442 7648
rect 7010 7650 7059 7669
rect 7079 7650 7454 7669
rect 7010 7647 7454 7650
rect 7286 7646 7454 7647
rect 8154 7660 8183 7662
rect 8154 7655 8186 7660
rect 8154 7637 8161 7655
rect 8181 7637 8186 7655
rect 8247 7659 8278 8053
rect 8299 8078 8467 8079
rect 8299 8075 8743 8078
rect 8299 8056 8674 8075
rect 8694 8056 8743 8075
rect 9311 8077 9420 8097
rect 9440 8077 9449 8097
rect 8299 8052 8743 8056
rect 8299 8050 8467 8052
rect 8299 7872 8326 8050
rect 8366 8012 8430 8024
rect 8706 8020 8743 8052
rect 8914 8051 9163 8073
rect 9311 8070 9449 8077
rect 9507 8097 9655 8106
rect 9507 8077 9516 8097
rect 9536 8077 9626 8097
rect 9646 8077 9655 8097
rect 9311 8068 9407 8070
rect 9507 8067 9655 8077
rect 9714 8097 9751 8107
rect 9826 8106 9863 8107
rect 9807 8104 9863 8106
rect 9714 8077 9722 8097
rect 9742 8077 9751 8097
rect 9563 8066 9599 8067
rect 8914 8020 8951 8051
rect 9127 8049 9163 8051
rect 9127 8020 9164 8049
rect 8366 8011 8401 8012
rect 8343 8006 8401 8011
rect 8343 7986 8346 8006
rect 8366 7992 8401 8006
rect 8421 7992 8430 8012
rect 8366 7984 8430 7992
rect 8392 7983 8430 7984
rect 8393 7982 8430 7983
rect 8496 8016 8532 8017
rect 8604 8016 8640 8017
rect 8496 8008 8640 8016
rect 8496 7988 8504 8008
rect 8524 8007 8612 8008
rect 8524 7988 8557 8007
rect 8496 7987 8557 7988
rect 8581 7988 8612 8007
rect 8632 7988 8640 8008
rect 8581 7987 8640 7988
rect 8496 7982 8640 7987
rect 8706 8012 8744 8020
rect 8812 8016 8848 8017
rect 8706 7992 8715 8012
rect 8735 7992 8744 8012
rect 8706 7983 8744 7992
rect 8763 8009 8848 8016
rect 8763 7989 8770 8009
rect 8791 8008 8848 8009
rect 8791 7989 8820 8008
rect 8763 7988 8820 7989
rect 8840 7988 8848 8008
rect 8706 7982 8743 7983
rect 8763 7982 8848 7988
rect 8914 8012 8952 8020
rect 9025 8016 9061 8017
rect 8914 7992 8923 8012
rect 8943 7992 8952 8012
rect 8914 7983 8952 7992
rect 8976 8008 9061 8016
rect 8976 7988 9033 8008
rect 9053 7988 9061 8008
rect 8914 7982 8951 7983
rect 8976 7982 9061 7988
rect 9127 8012 9165 8020
rect 9127 7992 9136 8012
rect 9156 7992 9165 8012
rect 9411 8007 9448 8008
rect 9714 8007 9751 8077
rect 9776 8097 9863 8104
rect 9776 8094 9834 8097
rect 9776 8074 9781 8094
rect 9802 8077 9834 8094
rect 9854 8077 9863 8097
rect 9802 8074 9863 8077
rect 9776 8067 9863 8074
rect 9922 8097 9959 8107
rect 9922 8077 9930 8097
rect 9950 8077 9959 8097
rect 9776 8066 9807 8067
rect 9410 8006 9751 8007
rect 9127 7983 9165 7992
rect 9335 8001 9751 8006
rect 9127 7982 9164 7983
rect 8550 7961 8586 7982
rect 8976 7961 9007 7982
rect 9335 7981 9338 8001
rect 9358 7981 9751 8001
rect 9922 8006 9959 8077
rect 9989 8106 10020 8159
rect 10322 8144 10359 8154
rect 10322 8126 10331 8144
rect 10349 8126 10359 8144
rect 10322 8117 10359 8126
rect 10771 8120 10806 8198
rect 11383 8188 11420 8211
rect 10039 8106 10076 8107
rect 9989 8097 10076 8106
rect 9989 8077 10047 8097
rect 10067 8077 10076 8097
rect 9989 8067 10076 8077
rect 10135 8097 10172 8107
rect 10135 8077 10143 8097
rect 10163 8077 10172 8097
rect 9989 8066 10020 8067
rect 10135 8006 10172 8077
rect 10327 8052 10358 8117
rect 10767 8111 10806 8120
rect 10767 8093 10777 8111
rect 10795 8093 10806 8111
rect 10767 8087 10806 8093
rect 10962 8163 11212 8187
rect 10962 8092 10999 8163
rect 11114 8102 11145 8103
rect 10767 8083 10804 8087
rect 10962 8072 10971 8092
rect 10991 8072 10999 8092
rect 10962 8062 10999 8072
rect 11058 8092 11145 8102
rect 11058 8072 11067 8092
rect 11087 8072 11145 8092
rect 11058 8063 11145 8072
rect 11058 8062 11095 8063
rect 10326 8042 10363 8052
rect 10326 8040 10336 8042
rect 10260 8038 10336 8040
rect 9922 7982 10172 8006
rect 10257 8024 10336 8038
rect 10354 8024 10363 8042
rect 10257 8021 10363 8024
rect 9729 7962 9750 7981
rect 10257 7962 10283 8021
rect 10326 8015 10363 8021
rect 10770 8012 10807 8021
rect 8383 7957 8483 7961
rect 8383 7953 8445 7957
rect 8383 7927 8390 7953
rect 8416 7931 8445 7953
rect 8471 7931 8483 7957
rect 8416 7927 8483 7931
rect 8383 7924 8483 7927
rect 8551 7924 8586 7961
rect 8648 7958 9007 7961
rect 8648 7953 8870 7958
rect 8648 7929 8661 7953
rect 8685 7934 8870 7953
rect 8894 7934 9007 7958
rect 8685 7929 9007 7934
rect 8648 7925 9007 7929
rect 9074 7953 9223 7961
rect 9074 7933 9085 7953
rect 9105 7933 9223 7953
rect 9729 7944 10283 7962
rect 10768 7994 10779 8012
rect 10797 7994 10807 8012
rect 11114 8010 11145 8063
rect 11175 8092 11212 8163
rect 11383 8168 11776 8188
rect 11796 8168 11799 8188
rect 11383 8163 11799 8168
rect 11383 8162 11724 8163
rect 11327 8102 11358 8103
rect 11175 8072 11184 8092
rect 11204 8072 11212 8092
rect 11175 8062 11212 8072
rect 11271 8095 11358 8102
rect 11271 8092 11332 8095
rect 11271 8072 11280 8092
rect 11300 8075 11332 8092
rect 11353 8075 11358 8095
rect 11300 8072 11358 8075
rect 11271 8065 11358 8072
rect 11383 8092 11420 8162
rect 11686 8161 11723 8162
rect 14692 8135 14719 8313
rect 14759 8275 14823 8287
rect 15099 8283 15136 8315
rect 15307 8314 15556 8336
rect 15307 8283 15344 8314
rect 15520 8312 15556 8314
rect 15699 8317 15737 8350
rect 15520 8283 15557 8312
rect 14759 8274 14794 8275
rect 14736 8269 14794 8274
rect 14736 8249 14739 8269
rect 14759 8255 14794 8269
rect 14814 8255 14823 8275
rect 14759 8247 14823 8255
rect 14785 8246 14823 8247
rect 14786 8245 14823 8246
rect 14889 8279 14925 8280
rect 14997 8279 15033 8280
rect 14889 8273 15033 8279
rect 14889 8271 14955 8273
rect 14889 8251 14897 8271
rect 14917 8252 14955 8271
rect 14977 8271 15033 8273
rect 14977 8252 15005 8271
rect 14917 8251 15005 8252
rect 15025 8251 15033 8271
rect 14889 8245 15033 8251
rect 15099 8275 15137 8283
rect 15205 8279 15241 8280
rect 15099 8255 15108 8275
rect 15128 8255 15137 8275
rect 15099 8246 15137 8255
rect 15156 8272 15241 8279
rect 15156 8252 15163 8272
rect 15184 8271 15241 8272
rect 15184 8252 15213 8271
rect 15156 8251 15213 8252
rect 15233 8251 15241 8271
rect 15099 8245 15136 8246
rect 15156 8245 15241 8251
rect 15307 8275 15345 8283
rect 15418 8279 15454 8280
rect 15307 8255 15316 8275
rect 15336 8255 15345 8275
rect 15307 8246 15345 8255
rect 15369 8271 15454 8279
rect 15369 8251 15426 8271
rect 15446 8251 15454 8271
rect 15307 8245 15344 8246
rect 15369 8245 15454 8251
rect 15520 8275 15558 8283
rect 15520 8255 15529 8275
rect 15549 8255 15558 8275
rect 15520 8246 15558 8255
rect 15699 8282 15735 8317
rect 16052 8313 16087 8350
rect 20391 8337 21018 8355
rect 16050 8304 16087 8313
rect 16050 8286 16060 8304
rect 16078 8286 16087 8304
rect 15699 8272 15736 8282
rect 16050 8276 16087 8286
rect 19973 8320 20141 8321
rect 20392 8320 20416 8337
rect 19973 8294 20417 8320
rect 19973 8292 20141 8294
rect 15699 8254 15709 8272
rect 15727 8254 15736 8272
rect 15520 8245 15557 8246
rect 15699 8245 15736 8254
rect 14943 8224 14979 8245
rect 15369 8224 15400 8245
rect 14776 8220 14876 8224
rect 14776 8216 14838 8220
rect 14776 8190 14783 8216
rect 14809 8194 14838 8216
rect 14864 8194 14876 8220
rect 14809 8190 14876 8194
rect 14776 8187 14876 8190
rect 14944 8187 14979 8224
rect 15041 8221 15400 8224
rect 15041 8216 15263 8221
rect 15041 8192 15054 8216
rect 15078 8197 15263 8216
rect 15287 8197 15400 8221
rect 15078 8192 15400 8197
rect 15041 8188 15400 8192
rect 15467 8216 15616 8224
rect 15467 8196 15478 8216
rect 15498 8196 15616 8216
rect 16053 8212 16090 8214
rect 16053 8211 16701 8212
rect 15467 8189 15616 8196
rect 16052 8205 16701 8211
rect 15467 8188 15508 8189
rect 14791 8135 14828 8136
rect 14887 8135 14924 8136
rect 14943 8135 14979 8187
rect 14998 8135 15035 8136
rect 14691 8126 14829 8135
rect 13627 8108 13658 8111
rect 11535 8102 11571 8103
rect 11383 8072 11392 8092
rect 11412 8072 11420 8092
rect 11271 8063 11327 8065
rect 11271 8062 11308 8063
rect 11383 8062 11420 8072
rect 11479 8092 11627 8102
rect 11727 8099 11823 8101
rect 11479 8072 11488 8092
rect 11508 8072 11598 8092
rect 11618 8072 11627 8092
rect 11479 8063 11627 8072
rect 11685 8092 11823 8099
rect 11685 8072 11694 8092
rect 11714 8072 11823 8092
rect 11685 8063 11823 8072
rect 13627 8082 13634 8108
rect 13653 8082 13658 8108
rect 11479 8062 11516 8063
rect 11535 8011 11571 8063
rect 11590 8062 11627 8063
rect 11686 8062 11723 8063
rect 11006 8009 11047 8010
rect 10329 7951 10366 7953
rect 10257 7943 10283 7944
rect 10326 7943 10366 7951
rect 9074 7926 9223 7933
rect 10326 7931 10338 7943
rect 10317 7926 10338 7931
rect 9074 7925 9115 7926
rect 9733 7925 10338 7926
rect 10356 7925 10366 7943
rect 8398 7872 8435 7873
rect 8494 7872 8531 7873
rect 8550 7872 8586 7924
rect 8605 7872 8642 7873
rect 8298 7863 8436 7872
rect 8298 7843 8407 7863
rect 8427 7843 8436 7863
rect 8298 7836 8436 7843
rect 8494 7863 8642 7872
rect 8494 7843 8503 7863
rect 8523 7843 8613 7863
rect 8633 7843 8642 7863
rect 8298 7834 8394 7836
rect 8494 7833 8642 7843
rect 8701 7863 8738 7873
rect 8813 7872 8850 7873
rect 8794 7870 8850 7872
rect 8701 7843 8709 7863
rect 8729 7843 8738 7863
rect 8550 7832 8586 7833
rect 8398 7773 8435 7774
rect 8701 7773 8738 7843
rect 8763 7863 8850 7870
rect 8763 7860 8821 7863
rect 8763 7840 8768 7860
rect 8789 7843 8821 7860
rect 8841 7843 8850 7863
rect 8789 7840 8850 7843
rect 8763 7833 8850 7840
rect 8909 7863 8946 7873
rect 8909 7843 8917 7863
rect 8937 7843 8946 7863
rect 8763 7832 8794 7833
rect 8397 7772 8738 7773
rect 8322 7767 8738 7772
rect 8322 7747 8325 7767
rect 8345 7747 8738 7767
rect 8909 7772 8946 7843
rect 8976 7872 9007 7925
rect 9733 7916 10366 7925
rect 9733 7909 10365 7916
rect 9733 7907 9795 7909
rect 9311 7897 9479 7898
rect 9733 7897 9755 7907
rect 9026 7872 9063 7873
rect 8976 7863 9063 7872
rect 8976 7843 9034 7863
rect 9054 7843 9063 7863
rect 8976 7833 9063 7843
rect 9122 7863 9159 7873
rect 9122 7843 9130 7863
rect 9150 7843 9159 7863
rect 8976 7832 9007 7833
rect 9122 7772 9159 7843
rect 8909 7748 9159 7772
rect 9311 7871 9755 7897
rect 9311 7869 9479 7871
rect 9311 7691 9338 7869
rect 9378 7831 9442 7843
rect 9718 7839 9755 7871
rect 9926 7870 10175 7892
rect 9926 7839 9963 7870
rect 10139 7868 10175 7870
rect 10139 7839 10176 7868
rect 9378 7830 9413 7831
rect 9355 7825 9413 7830
rect 9355 7805 9358 7825
rect 9378 7811 9413 7825
rect 9433 7811 9442 7831
rect 9378 7803 9442 7811
rect 9404 7802 9442 7803
rect 9405 7801 9442 7802
rect 9508 7835 9544 7836
rect 9616 7835 9652 7836
rect 9508 7827 9652 7835
rect 9508 7807 9516 7827
rect 9536 7807 9565 7827
rect 9508 7806 9565 7807
rect 9587 7807 9624 7827
rect 9644 7807 9652 7827
rect 9587 7806 9652 7807
rect 9508 7801 9652 7806
rect 9718 7831 9756 7839
rect 9824 7835 9860 7836
rect 9718 7811 9727 7831
rect 9747 7811 9756 7831
rect 9718 7802 9756 7811
rect 9775 7828 9860 7835
rect 9775 7808 9782 7828
rect 9803 7827 9860 7828
rect 9803 7808 9832 7827
rect 9775 7807 9832 7808
rect 9852 7807 9860 7827
rect 9718 7801 9755 7802
rect 9775 7801 9860 7807
rect 9926 7831 9964 7839
rect 10037 7835 10073 7836
rect 9926 7811 9935 7831
rect 9955 7811 9964 7831
rect 9926 7802 9964 7811
rect 9988 7827 10073 7835
rect 9988 7807 10045 7827
rect 10065 7807 10073 7827
rect 9926 7801 9963 7802
rect 9988 7801 10073 7807
rect 10139 7831 10177 7839
rect 10139 7811 10148 7831
rect 10168 7811 10177 7831
rect 10139 7802 10177 7811
rect 10139 7801 10176 7802
rect 9562 7780 9598 7801
rect 9988 7780 10019 7801
rect 9395 7776 9495 7780
rect 9395 7772 9457 7776
rect 9395 7746 9402 7772
rect 9428 7750 9457 7772
rect 9483 7750 9495 7776
rect 9428 7746 9495 7750
rect 9395 7743 9495 7746
rect 9563 7743 9598 7780
rect 9660 7777 10019 7780
rect 9660 7772 9882 7777
rect 9660 7748 9673 7772
rect 9697 7753 9882 7772
rect 9906 7753 10019 7777
rect 9697 7748 10019 7753
rect 9660 7744 10019 7748
rect 10086 7772 10235 7780
rect 10086 7752 10097 7772
rect 10117 7752 10235 7772
rect 10086 7745 10235 7752
rect 10326 7760 10365 7909
rect 10768 7845 10807 7994
rect 10898 8002 11047 8009
rect 10898 7982 11016 8002
rect 11036 7982 11047 8002
rect 10898 7974 11047 7982
rect 11114 8006 11473 8010
rect 11114 8001 11436 8006
rect 11114 7977 11227 8001
rect 11251 7982 11436 8001
rect 11460 7982 11473 8006
rect 11251 7977 11473 7982
rect 11114 7974 11473 7977
rect 11535 7974 11570 8011
rect 11638 8008 11738 8011
rect 11638 8004 11705 8008
rect 11638 7978 11650 8004
rect 11676 7982 11705 8004
rect 11731 7982 11738 8008
rect 11676 7978 11738 7982
rect 11638 7974 11738 7978
rect 11114 7953 11145 7974
rect 11535 7953 11571 7974
rect 10957 7952 10994 7953
rect 10956 7943 10994 7952
rect 10956 7923 10965 7943
rect 10985 7923 10994 7943
rect 10956 7915 10994 7923
rect 11060 7947 11145 7953
rect 11170 7952 11207 7953
rect 11060 7927 11068 7947
rect 11088 7927 11145 7947
rect 11060 7919 11145 7927
rect 11169 7943 11207 7952
rect 11169 7923 11178 7943
rect 11198 7923 11207 7943
rect 11060 7918 11096 7919
rect 11169 7915 11207 7923
rect 11273 7947 11358 7953
rect 11378 7952 11415 7953
rect 11273 7927 11281 7947
rect 11301 7946 11358 7947
rect 11301 7927 11330 7946
rect 11273 7926 11330 7927
rect 11351 7926 11358 7946
rect 11273 7919 11358 7926
rect 11377 7943 11415 7952
rect 11377 7923 11386 7943
rect 11406 7923 11415 7943
rect 11273 7918 11309 7919
rect 11377 7915 11415 7923
rect 11481 7948 11625 7953
rect 11481 7947 11546 7948
rect 11481 7927 11489 7947
rect 11509 7927 11546 7947
rect 11568 7947 11625 7948
rect 11568 7927 11597 7947
rect 11617 7927 11625 7947
rect 11481 7919 11625 7927
rect 11481 7918 11517 7919
rect 11589 7918 11625 7919
rect 11691 7952 11728 7953
rect 11691 7951 11729 7952
rect 11691 7943 11755 7951
rect 11691 7923 11700 7943
rect 11720 7929 11755 7943
rect 11775 7929 11778 7949
rect 11720 7924 11778 7929
rect 11720 7923 11755 7924
rect 10957 7886 10994 7915
rect 10958 7884 10994 7886
rect 11170 7884 11207 7915
rect 10958 7862 11207 7884
rect 11378 7883 11415 7915
rect 11691 7911 11755 7923
rect 11795 7885 11822 8063
rect 11654 7883 11822 7885
rect 11378 7857 11822 7883
rect 11974 7982 12224 8006
rect 11974 7911 12011 7982
rect 12126 7921 12157 7922
rect 11974 7891 11983 7911
rect 12003 7891 12011 7911
rect 11974 7881 12011 7891
rect 12070 7911 12157 7921
rect 12070 7891 12079 7911
rect 12099 7891 12157 7911
rect 12070 7882 12157 7891
rect 12070 7881 12107 7882
rect 11378 7847 11400 7857
rect 11654 7856 11822 7857
rect 11338 7845 11400 7847
rect 10768 7838 11400 7845
rect 10767 7829 11400 7838
rect 12126 7829 12157 7882
rect 12187 7911 12224 7982
rect 12395 7987 12788 8007
rect 12808 7987 12811 8007
rect 12395 7982 12811 7987
rect 12395 7981 12736 7982
rect 12339 7921 12370 7922
rect 12187 7891 12196 7911
rect 12216 7891 12224 7911
rect 12187 7881 12224 7891
rect 12283 7914 12370 7921
rect 12283 7911 12344 7914
rect 12283 7891 12292 7911
rect 12312 7894 12344 7911
rect 12365 7894 12370 7914
rect 12312 7891 12370 7894
rect 12283 7884 12370 7891
rect 12395 7911 12432 7981
rect 12698 7980 12735 7981
rect 12547 7921 12583 7922
rect 12395 7891 12404 7911
rect 12424 7891 12432 7911
rect 12283 7882 12339 7884
rect 12283 7881 12320 7882
rect 12395 7881 12432 7891
rect 12491 7911 12639 7921
rect 12739 7918 12835 7920
rect 12491 7891 12500 7911
rect 12520 7891 12610 7911
rect 12630 7891 12639 7911
rect 12491 7882 12639 7891
rect 12697 7911 12835 7918
rect 12697 7891 12706 7911
rect 12726 7891 12835 7911
rect 12697 7882 12835 7891
rect 12491 7881 12528 7882
rect 12547 7830 12583 7882
rect 12602 7881 12639 7882
rect 12698 7881 12735 7882
rect 10767 7811 10777 7829
rect 10795 7828 11400 7829
rect 12018 7828 12059 7829
rect 10795 7823 10816 7828
rect 10795 7811 10807 7823
rect 11910 7821 12059 7828
rect 10767 7803 10807 7811
rect 10850 7810 10876 7811
rect 10767 7801 10804 7803
rect 10086 7744 10127 7745
rect 9410 7691 9447 7692
rect 9506 7691 9543 7692
rect 9562 7691 9598 7743
rect 9617 7691 9654 7692
rect 9310 7682 9448 7691
rect 9310 7662 9419 7682
rect 9439 7662 9448 7682
rect 8247 7658 8417 7659
rect 8247 7643 8693 7658
rect 9310 7655 9448 7662
rect 9506 7682 9654 7691
rect 9506 7662 9515 7682
rect 9535 7662 9625 7682
rect 9645 7662 9654 7682
rect 9310 7653 9406 7655
rect 8154 7632 8186 7637
rect 6304 7619 6442 7628
rect 6098 7618 6135 7619
rect 6154 7567 6190 7619
rect 6209 7618 6246 7619
rect 6305 7618 6342 7619
rect 5625 7565 5666 7566
rect 4432 7543 5081 7549
rect 5517 7558 5666 7565
rect 4432 7542 5080 7543
rect 5043 7540 5080 7542
rect 3743 7527 3892 7534
rect 5517 7538 5635 7558
rect 5655 7538 5666 7558
rect 5517 7530 5666 7538
rect 5733 7562 6092 7566
rect 5733 7557 6055 7562
rect 5733 7533 5846 7557
rect 5870 7538 6055 7557
rect 6079 7538 6092 7562
rect 5870 7533 6092 7538
rect 5733 7530 6092 7533
rect 6154 7530 6189 7567
rect 6257 7564 6357 7567
rect 6257 7560 6324 7564
rect 6257 7534 6269 7560
rect 6295 7538 6324 7560
rect 6350 7538 6357 7564
rect 6295 7534 6357 7538
rect 6257 7530 6357 7534
rect 3743 7526 3784 7527
rect 3067 7473 3104 7474
rect 3163 7473 3200 7474
rect 3219 7473 3255 7525
rect 3274 7473 3311 7474
rect 2967 7464 3105 7473
rect 2967 7444 3076 7464
rect 3096 7444 3105 7464
rect 2967 7437 3105 7444
rect 3163 7464 3311 7473
rect 3163 7444 3172 7464
rect 3192 7444 3282 7464
rect 3302 7444 3311 7464
rect 2967 7435 3063 7437
rect 3163 7434 3311 7444
rect 3370 7464 3407 7474
rect 3482 7473 3519 7474
rect 3463 7471 3519 7473
rect 3370 7444 3378 7464
rect 3398 7444 3407 7464
rect 3219 7433 3255 7434
rect 3067 7374 3104 7375
rect 3370 7374 3407 7444
rect 3432 7464 3519 7471
rect 3432 7461 3490 7464
rect 3432 7441 3437 7461
rect 3458 7444 3490 7461
rect 3510 7444 3519 7464
rect 3458 7441 3519 7444
rect 3432 7434 3519 7441
rect 3578 7464 3615 7474
rect 3578 7444 3586 7464
rect 3606 7444 3615 7464
rect 3432 7433 3463 7434
rect 3066 7373 3407 7374
rect 2991 7368 3407 7373
rect 2991 7348 2994 7368
rect 3014 7348 3407 7368
rect 3578 7373 3615 7444
rect 3645 7473 3676 7526
rect 5733 7509 5764 7530
rect 6154 7509 6190 7530
rect 5397 7500 5434 7509
rect 5576 7508 5613 7509
rect 5397 7482 5406 7500
rect 5424 7482 5434 7500
rect 3695 7473 3732 7474
rect 3645 7464 3732 7473
rect 3645 7444 3703 7464
rect 3723 7444 3732 7464
rect 3645 7434 3732 7444
rect 3791 7464 3828 7474
rect 3791 7444 3799 7464
rect 3819 7444 3828 7464
rect 3645 7433 3676 7434
rect 3791 7373 3828 7444
rect 5046 7468 5083 7478
rect 5397 7472 5434 7482
rect 5046 7450 5055 7468
rect 5073 7450 5083 7468
rect 5046 7441 5083 7450
rect 5046 7417 5081 7441
rect 5398 7437 5434 7472
rect 5575 7499 5613 7508
rect 5575 7479 5584 7499
rect 5604 7479 5613 7499
rect 5575 7471 5613 7479
rect 5679 7503 5764 7509
rect 5789 7508 5826 7509
rect 5679 7483 5687 7503
rect 5707 7483 5764 7503
rect 5679 7475 5764 7483
rect 5788 7499 5826 7508
rect 5788 7479 5797 7499
rect 5817 7479 5826 7499
rect 5679 7474 5715 7475
rect 5788 7471 5826 7479
rect 5892 7503 5977 7509
rect 5997 7508 6034 7509
rect 5892 7483 5900 7503
rect 5920 7502 5977 7503
rect 5920 7483 5949 7502
rect 5892 7482 5949 7483
rect 5970 7482 5977 7502
rect 5892 7475 5977 7482
rect 5996 7499 6034 7508
rect 5996 7479 6005 7499
rect 6025 7479 6034 7499
rect 5892 7474 5928 7475
rect 5996 7471 6034 7479
rect 6100 7503 6244 7509
rect 6100 7483 6108 7503
rect 6128 7502 6216 7503
rect 6128 7483 6156 7502
rect 6100 7481 6156 7483
rect 6178 7483 6216 7502
rect 6236 7483 6244 7503
rect 6178 7481 6244 7483
rect 6100 7475 6244 7481
rect 6100 7474 6136 7475
rect 6208 7474 6244 7475
rect 6310 7508 6347 7509
rect 6310 7507 6348 7508
rect 6310 7499 6374 7507
rect 6310 7479 6319 7499
rect 6339 7485 6374 7499
rect 6394 7485 6397 7505
rect 6339 7480 6397 7485
rect 6339 7479 6374 7480
rect 5576 7442 5613 7471
rect 5044 7393 5081 7417
rect 5043 7387 5081 7393
rect 3578 7349 3828 7373
rect 4454 7369 5081 7387
rect 4036 7352 4204 7353
rect 4455 7352 4479 7369
rect 4036 7326 4480 7352
rect 4036 7324 4204 7326
rect 4036 7146 4063 7324
rect 4103 7286 4167 7298
rect 4443 7294 4480 7326
rect 4651 7325 4900 7347
rect 4651 7294 4688 7325
rect 4864 7323 4900 7325
rect 5043 7328 5081 7369
rect 5396 7396 5434 7437
rect 5577 7440 5613 7442
rect 5789 7440 5826 7471
rect 5577 7418 5826 7440
rect 5997 7439 6034 7471
rect 6310 7467 6374 7479
rect 6414 7441 6441 7619
rect 6273 7439 6441 7441
rect 5997 7413 6441 7439
rect 5998 7396 6022 7413
rect 6273 7412 6441 7413
rect 5396 7378 6023 7396
rect 6649 7392 6899 7416
rect 5396 7372 5434 7378
rect 5396 7348 5433 7372
rect 4864 7294 4901 7323
rect 4103 7285 4138 7286
rect 4080 7280 4138 7285
rect 4080 7260 4083 7280
rect 4103 7266 4138 7280
rect 4158 7266 4167 7286
rect 4103 7258 4167 7266
rect 4129 7257 4167 7258
rect 4130 7256 4167 7257
rect 4233 7290 4269 7291
rect 4341 7290 4377 7291
rect 4233 7284 4377 7290
rect 4233 7282 4299 7284
rect 4233 7262 4241 7282
rect 4261 7263 4299 7282
rect 4321 7282 4377 7284
rect 4321 7263 4349 7282
rect 4261 7262 4349 7263
rect 4369 7262 4377 7282
rect 4233 7256 4377 7262
rect 4443 7286 4481 7294
rect 4549 7290 4585 7291
rect 4443 7266 4452 7286
rect 4472 7266 4481 7286
rect 4443 7257 4481 7266
rect 4500 7283 4585 7290
rect 4500 7263 4507 7283
rect 4528 7282 4585 7283
rect 4528 7263 4557 7282
rect 4500 7262 4557 7263
rect 4577 7262 4585 7282
rect 4443 7256 4480 7257
rect 4500 7256 4585 7262
rect 4651 7286 4689 7294
rect 4762 7290 4798 7291
rect 4651 7266 4660 7286
rect 4680 7266 4689 7286
rect 4651 7257 4689 7266
rect 4713 7282 4798 7290
rect 4713 7262 4770 7282
rect 4790 7262 4798 7282
rect 4651 7256 4688 7257
rect 4713 7256 4798 7262
rect 4864 7286 4902 7294
rect 4864 7266 4873 7286
rect 4893 7266 4902 7286
rect 4864 7257 4902 7266
rect 5043 7293 5079 7328
rect 5396 7324 5431 7348
rect 5394 7315 5431 7324
rect 5394 7297 5404 7315
rect 5422 7297 5431 7315
rect 5043 7283 5080 7293
rect 5394 7287 5431 7297
rect 6649 7321 6686 7392
rect 6801 7331 6832 7332
rect 6649 7301 6658 7321
rect 6678 7301 6686 7321
rect 6649 7291 6686 7301
rect 6745 7321 6832 7331
rect 6745 7301 6754 7321
rect 6774 7301 6832 7321
rect 6745 7292 6832 7301
rect 6745 7291 6782 7292
rect 5043 7265 5053 7283
rect 5071 7265 5080 7283
rect 4864 7256 4901 7257
rect 5043 7256 5080 7265
rect 4287 7235 4323 7256
rect 4713 7235 4744 7256
rect 6801 7239 6832 7292
rect 6862 7321 6899 7392
rect 7070 7397 7463 7417
rect 7483 7397 7486 7417
rect 7070 7392 7486 7397
rect 7070 7391 7411 7392
rect 7014 7331 7045 7332
rect 6862 7301 6871 7321
rect 6891 7301 6899 7321
rect 6862 7291 6899 7301
rect 6958 7324 7045 7331
rect 6958 7321 7019 7324
rect 6958 7301 6967 7321
rect 6987 7304 7019 7321
rect 7040 7304 7045 7324
rect 6987 7301 7045 7304
rect 6958 7294 7045 7301
rect 7070 7321 7107 7391
rect 7373 7390 7410 7391
rect 7222 7331 7258 7332
rect 7070 7301 7079 7321
rect 7099 7301 7107 7321
rect 6958 7292 7014 7294
rect 6958 7291 6995 7292
rect 7070 7291 7107 7301
rect 7166 7321 7314 7331
rect 7414 7328 7510 7330
rect 7166 7301 7175 7321
rect 7195 7301 7285 7321
rect 7305 7301 7314 7321
rect 7166 7292 7314 7301
rect 7372 7321 7510 7328
rect 7372 7301 7381 7321
rect 7401 7301 7510 7321
rect 7372 7292 7510 7301
rect 7166 7291 7203 7292
rect 7222 7240 7258 7292
rect 7277 7291 7314 7292
rect 7373 7291 7410 7292
rect 6693 7238 6734 7239
rect 4120 7231 4220 7235
rect 4120 7227 4182 7231
rect 4120 7201 4127 7227
rect 4153 7205 4182 7227
rect 4208 7205 4220 7231
rect 4153 7201 4220 7205
rect 4120 7198 4220 7201
rect 4288 7198 4323 7235
rect 4385 7232 4744 7235
rect 4385 7227 4607 7232
rect 4385 7203 4398 7227
rect 4422 7208 4607 7227
rect 4631 7208 4744 7232
rect 4422 7203 4744 7208
rect 4385 7199 4744 7203
rect 4811 7227 4960 7235
rect 4811 7207 4822 7227
rect 4842 7207 4960 7227
rect 6585 7231 6734 7238
rect 5397 7223 5434 7225
rect 5397 7222 6045 7223
rect 4811 7200 4960 7207
rect 5396 7216 6045 7222
rect 4811 7199 4852 7200
rect 4135 7146 4172 7147
rect 4231 7146 4268 7147
rect 4287 7146 4323 7198
rect 4342 7146 4379 7147
rect 4035 7137 4173 7146
rect 3023 7118 3191 7119
rect 3023 7115 3467 7118
rect 3023 7096 3398 7115
rect 3418 7096 3467 7115
rect 4035 7117 4144 7137
rect 4164 7117 4173 7137
rect 3023 7092 3467 7096
rect 3023 7090 3191 7092
rect 3023 6912 3050 7090
rect 3090 7052 3154 7064
rect 3430 7060 3467 7092
rect 3638 7091 3887 7113
rect 4035 7110 4173 7117
rect 4231 7137 4379 7146
rect 4231 7117 4240 7137
rect 4260 7117 4350 7137
rect 4370 7117 4379 7137
rect 4035 7108 4131 7110
rect 4231 7107 4379 7117
rect 4438 7137 4475 7147
rect 4550 7146 4587 7147
rect 4531 7144 4587 7146
rect 4438 7117 4446 7137
rect 4466 7117 4475 7137
rect 4287 7106 4323 7107
rect 3638 7060 3675 7091
rect 3851 7089 3887 7091
rect 3851 7060 3888 7089
rect 3090 7051 3125 7052
rect 3067 7046 3125 7051
rect 3067 7026 3070 7046
rect 3090 7032 3125 7046
rect 3145 7032 3154 7052
rect 3090 7024 3154 7032
rect 3116 7023 3154 7024
rect 3117 7022 3154 7023
rect 3220 7056 3256 7057
rect 3328 7056 3364 7057
rect 3220 7048 3364 7056
rect 3220 7028 3228 7048
rect 3248 7028 3280 7048
rect 3304 7028 3336 7048
rect 3356 7028 3364 7048
rect 3220 7022 3364 7028
rect 3430 7052 3468 7060
rect 3536 7056 3572 7057
rect 3430 7032 3439 7052
rect 3459 7032 3468 7052
rect 3430 7023 3468 7032
rect 3487 7049 3572 7056
rect 3487 7029 3494 7049
rect 3515 7048 3572 7049
rect 3515 7029 3544 7048
rect 3487 7028 3544 7029
rect 3564 7028 3572 7048
rect 3430 7022 3467 7023
rect 3487 7022 3572 7028
rect 3638 7052 3676 7060
rect 3749 7056 3785 7057
rect 3638 7032 3647 7052
rect 3667 7032 3676 7052
rect 3638 7023 3676 7032
rect 3700 7048 3785 7056
rect 3700 7028 3757 7048
rect 3777 7028 3785 7048
rect 3638 7022 3675 7023
rect 3700 7022 3785 7028
rect 3851 7052 3889 7060
rect 3851 7032 3860 7052
rect 3880 7032 3889 7052
rect 4135 7047 4172 7048
rect 4438 7047 4475 7117
rect 4500 7137 4587 7144
rect 4500 7134 4558 7137
rect 4500 7114 4505 7134
rect 4526 7117 4558 7134
rect 4578 7117 4587 7137
rect 4526 7114 4587 7117
rect 4500 7107 4587 7114
rect 4646 7137 4683 7147
rect 4646 7117 4654 7137
rect 4674 7117 4683 7137
rect 4500 7106 4531 7107
rect 4134 7046 4475 7047
rect 3851 7023 3889 7032
rect 4059 7041 4475 7046
rect 3851 7022 3888 7023
rect 3274 7001 3310 7022
rect 3700 7001 3731 7022
rect 4059 7021 4062 7041
rect 4082 7021 4475 7041
rect 4646 7046 4683 7117
rect 4713 7146 4744 7199
rect 5396 7198 5406 7216
rect 5424 7202 6045 7216
rect 6585 7211 6703 7231
rect 6723 7211 6734 7231
rect 6585 7203 6734 7211
rect 6801 7235 7160 7239
rect 6801 7230 7123 7235
rect 6801 7206 6914 7230
rect 6938 7211 7123 7230
rect 7147 7211 7160 7235
rect 6938 7206 7160 7211
rect 6801 7203 7160 7206
rect 7222 7203 7257 7240
rect 7325 7237 7425 7240
rect 7325 7233 7392 7237
rect 7325 7207 7337 7233
rect 7363 7211 7392 7233
rect 7418 7211 7425 7237
rect 7363 7207 7425 7211
rect 7325 7203 7425 7207
rect 5424 7198 5434 7202
rect 5875 7201 6045 7202
rect 5046 7184 5083 7194
rect 5046 7166 5055 7184
rect 5073 7166 5083 7184
rect 5046 7157 5083 7166
rect 5396 7188 5434 7198
rect 4763 7146 4800 7147
rect 4713 7137 4800 7146
rect 4713 7117 4771 7137
rect 4791 7117 4800 7137
rect 4713 7107 4800 7117
rect 4859 7137 4896 7147
rect 4859 7117 4867 7137
rect 4887 7117 4896 7137
rect 4713 7106 4744 7107
rect 4859 7046 4896 7117
rect 5051 7092 5082 7157
rect 5396 7110 5431 7188
rect 6008 7178 6045 7201
rect 6801 7182 6832 7203
rect 7222 7182 7258 7203
rect 6644 7181 6681 7182
rect 5392 7101 5431 7110
rect 5050 7082 5087 7092
rect 5050 7080 5060 7082
rect 4984 7078 5060 7080
rect 4646 7022 4896 7046
rect 4981 7064 5060 7078
rect 5078 7064 5087 7082
rect 5392 7083 5402 7101
rect 5420 7083 5431 7101
rect 5392 7077 5431 7083
rect 5587 7153 5837 7177
rect 5587 7082 5624 7153
rect 5739 7092 5770 7093
rect 5392 7073 5429 7077
rect 4981 7061 5087 7064
rect 4453 7002 4474 7021
rect 4981 7002 5007 7061
rect 5050 7055 5087 7061
rect 5587 7062 5596 7082
rect 5616 7062 5624 7082
rect 5587 7052 5624 7062
rect 5683 7082 5770 7092
rect 5683 7062 5692 7082
rect 5712 7062 5770 7082
rect 5683 7053 5770 7062
rect 5683 7052 5720 7053
rect 5395 7002 5432 7011
rect 3107 6997 3207 7001
rect 3107 6993 3169 6997
rect 3107 6967 3114 6993
rect 3140 6971 3169 6993
rect 3195 6971 3207 6997
rect 3140 6967 3207 6971
rect 3107 6964 3207 6967
rect 3275 6964 3310 7001
rect 3372 6998 3731 7001
rect 3372 6993 3594 6998
rect 3372 6969 3385 6993
rect 3409 6974 3594 6993
rect 3618 6974 3731 6998
rect 3409 6969 3731 6974
rect 3372 6965 3731 6969
rect 3798 6993 3947 7001
rect 3798 6973 3809 6993
rect 3829 6973 3947 6993
rect 4453 6984 5007 7002
rect 5053 6991 5090 6993
rect 4981 6983 5007 6984
rect 5050 6983 5090 6991
rect 3798 6966 3947 6973
rect 5050 6971 5062 6983
rect 5041 6966 5062 6971
rect 3798 6965 3839 6966
rect 4457 6965 5062 6966
rect 5080 6965 5090 6983
rect 3122 6912 3159 6913
rect 3218 6912 3255 6913
rect 3274 6912 3310 6964
rect 3329 6912 3366 6913
rect 3022 6903 3160 6912
rect 3022 6883 3131 6903
rect 3151 6883 3160 6903
rect 3022 6876 3160 6883
rect 3218 6903 3366 6912
rect 3218 6883 3227 6903
rect 3247 6883 3337 6903
rect 3357 6883 3366 6903
rect 3022 6874 3118 6876
rect 3218 6873 3366 6883
rect 3425 6903 3462 6913
rect 3537 6912 3574 6913
rect 3518 6910 3574 6912
rect 3425 6883 3433 6903
rect 3453 6883 3462 6903
rect 3274 6872 3310 6873
rect 3122 6813 3159 6814
rect 3425 6813 3462 6883
rect 3487 6903 3574 6910
rect 3487 6900 3545 6903
rect 3487 6880 3492 6900
rect 3513 6883 3545 6900
rect 3565 6883 3574 6903
rect 3513 6880 3574 6883
rect 3487 6873 3574 6880
rect 3633 6903 3670 6913
rect 3633 6883 3641 6903
rect 3661 6883 3670 6903
rect 3487 6872 3518 6873
rect 3121 6812 3462 6813
rect 3046 6807 3462 6812
rect 3046 6787 3049 6807
rect 3069 6787 3462 6807
rect 3633 6812 3670 6883
rect 3700 6912 3731 6965
rect 4457 6956 5090 6965
rect 5393 6984 5404 7002
rect 5422 6984 5432 7002
rect 5739 7000 5770 7053
rect 5800 7082 5837 7153
rect 6008 7158 6401 7178
rect 6421 7158 6424 7178
rect 6008 7153 6424 7158
rect 6643 7172 6681 7181
rect 6008 7152 6349 7153
rect 6643 7152 6652 7172
rect 6672 7152 6681 7172
rect 5952 7092 5983 7093
rect 5800 7062 5809 7082
rect 5829 7062 5837 7082
rect 5800 7052 5837 7062
rect 5896 7085 5983 7092
rect 5896 7082 5957 7085
rect 5896 7062 5905 7082
rect 5925 7065 5957 7082
rect 5978 7065 5983 7085
rect 5925 7062 5983 7065
rect 5896 7055 5983 7062
rect 6008 7082 6045 7152
rect 6311 7151 6348 7152
rect 6643 7144 6681 7152
rect 6747 7176 6832 7182
rect 6857 7181 6894 7182
rect 6747 7156 6755 7176
rect 6775 7156 6832 7176
rect 6747 7148 6832 7156
rect 6856 7172 6894 7181
rect 6856 7152 6865 7172
rect 6885 7152 6894 7172
rect 6747 7147 6783 7148
rect 6856 7144 6894 7152
rect 6960 7176 7045 7182
rect 7065 7181 7102 7182
rect 6960 7156 6968 7176
rect 6988 7175 7045 7176
rect 6988 7156 7017 7175
rect 6960 7155 7017 7156
rect 7038 7155 7045 7175
rect 6960 7148 7045 7155
rect 7064 7172 7102 7181
rect 7064 7152 7073 7172
rect 7093 7152 7102 7172
rect 6960 7147 6996 7148
rect 7064 7144 7102 7152
rect 7168 7176 7312 7182
rect 7168 7156 7176 7176
rect 7196 7174 7284 7176
rect 7196 7157 7232 7174
rect 7256 7157 7284 7174
rect 7196 7156 7284 7157
rect 7304 7156 7312 7176
rect 7168 7148 7312 7156
rect 7168 7147 7204 7148
rect 7276 7147 7312 7148
rect 7378 7181 7415 7182
rect 7378 7180 7416 7181
rect 7378 7172 7442 7180
rect 7378 7152 7387 7172
rect 7407 7158 7442 7172
rect 7462 7158 7465 7178
rect 7407 7153 7465 7158
rect 7407 7152 7442 7153
rect 6644 7115 6681 7144
rect 6645 7113 6681 7115
rect 6857 7113 6894 7144
rect 6160 7092 6196 7093
rect 6008 7062 6017 7082
rect 6037 7062 6045 7082
rect 5896 7053 5952 7055
rect 5896 7052 5933 7053
rect 6008 7052 6045 7062
rect 6104 7082 6252 7092
rect 6645 7091 6894 7113
rect 7065 7112 7102 7144
rect 7378 7140 7442 7152
rect 7482 7114 7509 7292
rect 7341 7112 7509 7114
rect 7065 7101 7509 7112
rect 6352 7089 6448 7091
rect 6104 7062 6113 7082
rect 6133 7062 6223 7082
rect 6243 7062 6252 7082
rect 6104 7053 6252 7062
rect 6310 7082 6448 7089
rect 7065 7086 7511 7101
rect 7341 7085 7511 7086
rect 6310 7062 6319 7082
rect 6339 7062 6448 7082
rect 6310 7053 6448 7062
rect 6104 7052 6141 7053
rect 6160 7001 6196 7053
rect 6215 7052 6252 7053
rect 6311 7052 6348 7053
rect 5631 6999 5672 7000
rect 4457 6949 5089 6956
rect 4457 6947 4519 6949
rect 4035 6937 4203 6938
rect 4457 6937 4479 6947
rect 3750 6912 3787 6913
rect 3700 6903 3787 6912
rect 3700 6883 3758 6903
rect 3778 6883 3787 6903
rect 3700 6873 3787 6883
rect 3846 6903 3883 6913
rect 3846 6883 3854 6903
rect 3874 6883 3883 6903
rect 3700 6872 3731 6873
rect 3846 6812 3883 6883
rect 3633 6788 3883 6812
rect 4035 6911 4479 6937
rect 4035 6909 4203 6911
rect 4035 6731 4062 6909
rect 4102 6871 4166 6883
rect 4442 6879 4479 6911
rect 4650 6910 4899 6932
rect 4650 6879 4687 6910
rect 4863 6908 4899 6910
rect 4863 6879 4900 6908
rect 4102 6870 4137 6871
rect 4079 6865 4137 6870
rect 4079 6845 4082 6865
rect 4102 6851 4137 6865
rect 4157 6851 4166 6871
rect 4102 6843 4166 6851
rect 4128 6842 4166 6843
rect 4129 6841 4166 6842
rect 4232 6875 4268 6876
rect 4340 6875 4376 6876
rect 4232 6867 4376 6875
rect 4232 6847 4240 6867
rect 4260 6847 4289 6867
rect 4232 6846 4289 6847
rect 4311 6847 4348 6867
rect 4368 6847 4376 6867
rect 4311 6846 4376 6847
rect 4232 6841 4376 6846
rect 4442 6871 4480 6879
rect 4548 6875 4584 6876
rect 4442 6851 4451 6871
rect 4471 6851 4480 6871
rect 4442 6842 4480 6851
rect 4499 6868 4584 6875
rect 4499 6848 4506 6868
rect 4527 6867 4584 6868
rect 4527 6848 4556 6867
rect 4499 6847 4556 6848
rect 4576 6847 4584 6867
rect 4442 6841 4479 6842
rect 4499 6841 4584 6847
rect 4650 6871 4688 6879
rect 4761 6875 4797 6876
rect 4650 6851 4659 6871
rect 4679 6851 4688 6871
rect 4650 6842 4688 6851
rect 4712 6867 4797 6875
rect 4712 6847 4769 6867
rect 4789 6847 4797 6867
rect 4650 6841 4687 6842
rect 4712 6841 4797 6847
rect 4863 6871 4901 6879
rect 4863 6851 4872 6871
rect 4892 6851 4901 6871
rect 4863 6842 4901 6851
rect 4863 6841 4900 6842
rect 4286 6820 4322 6841
rect 4712 6820 4743 6841
rect 4119 6816 4219 6820
rect 4119 6812 4181 6816
rect 4119 6786 4126 6812
rect 4152 6790 4181 6812
rect 4207 6790 4219 6816
rect 4152 6786 4219 6790
rect 4119 6783 4219 6786
rect 4287 6783 4322 6820
rect 4384 6817 4743 6820
rect 4384 6812 4606 6817
rect 4384 6788 4397 6812
rect 4421 6793 4606 6812
rect 4630 6793 4743 6817
rect 4421 6788 4743 6793
rect 4384 6784 4743 6788
rect 4810 6812 4959 6820
rect 4810 6792 4821 6812
rect 4841 6792 4959 6812
rect 4810 6785 4959 6792
rect 5050 6800 5089 6949
rect 5393 6835 5432 6984
rect 5523 6992 5672 6999
rect 5523 6972 5641 6992
rect 5661 6972 5672 6992
rect 5523 6964 5672 6972
rect 5739 6996 6098 7000
rect 5739 6991 6061 6996
rect 5739 6967 5852 6991
rect 5876 6972 6061 6991
rect 6085 6972 6098 6996
rect 5876 6967 6098 6972
rect 5739 6964 6098 6967
rect 6160 6964 6195 7001
rect 6263 6998 6363 7001
rect 6263 6994 6330 6998
rect 6263 6968 6275 6994
rect 6301 6972 6330 6994
rect 6356 6972 6363 6998
rect 6301 6968 6363 6972
rect 6263 6964 6363 6968
rect 5739 6943 5770 6964
rect 6160 6943 6196 6964
rect 5582 6942 5619 6943
rect 5581 6933 5619 6942
rect 5581 6913 5590 6933
rect 5610 6913 5619 6933
rect 5581 6905 5619 6913
rect 5685 6937 5770 6943
rect 5795 6942 5832 6943
rect 5685 6917 5693 6937
rect 5713 6917 5770 6937
rect 5685 6909 5770 6917
rect 5794 6933 5832 6942
rect 5794 6913 5803 6933
rect 5823 6913 5832 6933
rect 5685 6908 5721 6909
rect 5794 6905 5832 6913
rect 5898 6937 5983 6943
rect 6003 6942 6040 6943
rect 5898 6917 5906 6937
rect 5926 6936 5983 6937
rect 5926 6917 5955 6936
rect 5898 6916 5955 6917
rect 5976 6916 5983 6936
rect 5898 6909 5983 6916
rect 6002 6933 6040 6942
rect 6002 6913 6011 6933
rect 6031 6913 6040 6933
rect 5898 6908 5934 6909
rect 6002 6905 6040 6913
rect 6106 6938 6250 6943
rect 6106 6937 6171 6938
rect 6106 6917 6114 6937
rect 6134 6917 6171 6937
rect 6193 6937 6250 6938
rect 6193 6917 6222 6937
rect 6242 6917 6250 6937
rect 6106 6909 6250 6917
rect 6106 6908 6142 6909
rect 6214 6908 6250 6909
rect 6316 6942 6353 6943
rect 6316 6941 6354 6942
rect 6316 6933 6380 6941
rect 6316 6913 6325 6933
rect 6345 6919 6380 6933
rect 6400 6919 6403 6939
rect 6345 6914 6403 6919
rect 6345 6913 6380 6914
rect 5582 6876 5619 6905
rect 5583 6874 5619 6876
rect 5795 6874 5832 6905
rect 5583 6852 5832 6874
rect 6003 6873 6040 6905
rect 6316 6901 6380 6913
rect 6420 6875 6447 7053
rect 6279 6873 6447 6875
rect 6003 6847 6447 6873
rect 6599 6972 6849 6996
rect 6599 6901 6636 6972
rect 6751 6911 6782 6912
rect 6599 6881 6608 6901
rect 6628 6881 6636 6901
rect 6599 6871 6636 6881
rect 6695 6901 6782 6911
rect 6695 6881 6704 6901
rect 6724 6881 6782 6901
rect 6695 6872 6782 6881
rect 6695 6871 6732 6872
rect 6003 6837 6025 6847
rect 6279 6846 6447 6847
rect 5963 6835 6025 6837
rect 5393 6828 6025 6835
rect 4810 6784 4851 6785
rect 4134 6731 4171 6732
rect 4230 6731 4267 6732
rect 4286 6731 4322 6783
rect 4341 6731 4378 6732
rect 4034 6722 4172 6731
rect 4034 6702 4143 6722
rect 4163 6702 4172 6722
rect 4034 6695 4172 6702
rect 4230 6722 4378 6731
rect 4230 6702 4239 6722
rect 4259 6702 4349 6722
rect 4369 6702 4378 6722
rect 4034 6693 4130 6695
rect 4230 6692 4378 6702
rect 4437 6722 4474 6732
rect 4549 6731 4586 6732
rect 4530 6729 4586 6731
rect 4437 6702 4445 6722
rect 4465 6702 4474 6722
rect 4286 6691 4322 6692
rect 2749 6629 2757 6648
rect 2780 6629 2786 6648
rect 2749 6618 2786 6629
rect 2815 6651 2983 6652
rect 2815 6625 3259 6651
rect 2815 6623 2983 6625
rect 2752 6558 2785 6618
rect 997 6479 1165 6481
rect 721 6453 1165 6479
rect 722 6436 746 6453
rect 997 6452 1165 6453
rect 1533 6481 1783 6505
rect 120 6418 747 6436
rect 120 6412 158 6418
rect 122 6366 157 6412
rect 1533 6410 1570 6481
rect 1685 6420 1716 6421
rect 1533 6390 1542 6410
rect 1562 6390 1570 6410
rect 1533 6380 1570 6390
rect 1629 6410 1716 6420
rect 1629 6390 1638 6410
rect 1658 6390 1716 6410
rect 1629 6381 1716 6390
rect 1629 6380 1666 6381
rect 120 6357 157 6366
rect 120 6339 130 6357
rect 148 6339 157 6357
rect 120 6329 157 6339
rect 1685 6328 1716 6381
rect 1746 6410 1783 6481
rect 1954 6486 2347 6506
rect 2367 6486 2370 6506
rect 1954 6481 2370 6486
rect 1954 6480 2295 6481
rect 1898 6420 1929 6421
rect 1746 6390 1755 6410
rect 1775 6390 1783 6410
rect 1746 6380 1783 6390
rect 1842 6413 1929 6420
rect 1842 6410 1903 6413
rect 1842 6390 1851 6410
rect 1871 6393 1903 6410
rect 1924 6393 1929 6413
rect 1871 6390 1929 6393
rect 1842 6383 1929 6390
rect 1954 6410 1991 6480
rect 2257 6479 2294 6480
rect 2106 6420 2142 6421
rect 1954 6390 1963 6410
rect 1983 6390 1991 6410
rect 1842 6381 1898 6383
rect 1842 6380 1879 6381
rect 1954 6380 1991 6390
rect 2050 6410 2198 6420
rect 2298 6417 2394 6419
rect 2050 6390 2059 6410
rect 2079 6390 2169 6410
rect 2189 6390 2198 6410
rect 2050 6381 2198 6390
rect 2256 6410 2394 6417
rect 2256 6390 2265 6410
rect 2285 6390 2394 6410
rect 2256 6381 2394 6390
rect 2050 6380 2087 6381
rect 2106 6329 2142 6381
rect 2161 6380 2198 6381
rect 2257 6380 2294 6381
rect 1577 6327 1618 6328
rect 1469 6320 1618 6327
rect 1469 6300 1587 6320
rect 1607 6300 1618 6320
rect 1469 6292 1618 6300
rect 1685 6324 2044 6328
rect 1685 6319 2007 6324
rect 1685 6295 1798 6319
rect 1822 6300 2007 6319
rect 2031 6300 2044 6324
rect 1822 6295 2044 6300
rect 1685 6292 2044 6295
rect 2106 6292 2141 6329
rect 2209 6326 2309 6329
rect 2209 6322 2276 6326
rect 2209 6296 2221 6322
rect 2247 6300 2276 6322
rect 2302 6300 2309 6326
rect 2247 6296 2309 6300
rect 2209 6292 2309 6296
rect 1685 6271 1716 6292
rect 2106 6271 2142 6292
rect 1528 6270 1565 6271
rect 123 6265 160 6267
rect 123 6264 771 6265
rect 122 6258 771 6264
rect 122 6240 132 6258
rect 150 6244 771 6258
rect 150 6240 160 6244
rect 601 6243 771 6244
rect 122 6230 160 6240
rect 122 6152 157 6230
rect 734 6220 771 6243
rect 1527 6261 1565 6270
rect 1527 6241 1536 6261
rect 1556 6241 1565 6261
rect 1527 6233 1565 6241
rect 1631 6265 1716 6271
rect 1741 6270 1778 6271
rect 1631 6245 1639 6265
rect 1659 6245 1716 6265
rect 1631 6237 1716 6245
rect 1740 6261 1778 6270
rect 1740 6241 1749 6261
rect 1769 6241 1778 6261
rect 1631 6236 1667 6237
rect 1740 6233 1778 6241
rect 1844 6265 1929 6271
rect 1949 6270 1986 6271
rect 1844 6245 1852 6265
rect 1872 6264 1929 6265
rect 1872 6245 1901 6264
rect 1844 6244 1901 6245
rect 1922 6244 1929 6264
rect 1844 6237 1929 6244
rect 1948 6261 1986 6270
rect 1948 6241 1957 6261
rect 1977 6241 1986 6261
rect 1844 6236 1880 6237
rect 1948 6233 1986 6241
rect 2052 6269 2196 6271
rect 2052 6265 2110 6269
rect 2052 6245 2060 6265
rect 2080 6245 2110 6265
rect 2052 6243 2110 6245
rect 2135 6265 2196 6269
rect 2135 6245 2168 6265
rect 2188 6245 2196 6265
rect 2135 6243 2196 6245
rect 2052 6237 2196 6243
rect 2052 6236 2088 6237
rect 2160 6236 2196 6237
rect 2262 6270 2299 6271
rect 2262 6269 2300 6270
rect 2262 6261 2326 6269
rect 2262 6241 2271 6261
rect 2291 6247 2326 6261
rect 2346 6247 2349 6267
rect 2291 6242 2349 6247
rect 2291 6241 2326 6242
rect 118 6143 157 6152
rect 118 6125 128 6143
rect 146 6125 157 6143
rect 118 6119 157 6125
rect 313 6195 563 6219
rect 313 6124 350 6195
rect 465 6134 496 6135
rect 118 6115 155 6119
rect 313 6104 322 6124
rect 342 6104 350 6124
rect 313 6094 350 6104
rect 409 6124 496 6134
rect 409 6104 418 6124
rect 438 6104 496 6124
rect 409 6095 496 6104
rect 409 6094 446 6095
rect 121 6044 158 6053
rect 119 6026 130 6044
rect 148 6026 158 6044
rect 465 6042 496 6095
rect 526 6124 563 6195
rect 734 6200 1127 6220
rect 1147 6200 1150 6220
rect 1528 6204 1565 6233
rect 734 6195 1150 6200
rect 1529 6202 1565 6204
rect 1741 6202 1778 6233
rect 734 6194 1075 6195
rect 678 6134 709 6135
rect 526 6104 535 6124
rect 555 6104 563 6124
rect 526 6094 563 6104
rect 622 6127 709 6134
rect 622 6124 683 6127
rect 622 6104 631 6124
rect 651 6107 683 6124
rect 704 6107 709 6127
rect 651 6104 709 6107
rect 622 6097 709 6104
rect 734 6124 771 6194
rect 1037 6193 1074 6194
rect 1529 6180 1778 6202
rect 1949 6201 1986 6233
rect 2262 6229 2326 6241
rect 2366 6203 2393 6381
rect 2225 6201 2393 6203
rect 1949 6175 2393 6201
rect 2225 6174 2393 6175
rect 886 6134 922 6135
rect 734 6104 743 6124
rect 763 6104 771 6124
rect 622 6095 678 6097
rect 622 6094 659 6095
rect 734 6094 771 6104
rect 830 6124 978 6134
rect 1078 6131 1174 6133
rect 830 6104 839 6124
rect 859 6104 949 6124
rect 969 6104 978 6124
rect 830 6095 978 6104
rect 1036 6124 1174 6131
rect 1036 6104 1045 6124
rect 1065 6104 1174 6124
rect 1036 6095 1174 6104
rect 830 6094 867 6095
rect 886 6043 922 6095
rect 941 6094 978 6095
rect 1037 6094 1074 6095
rect 357 6041 398 6042
rect 119 5877 158 6026
rect 249 6034 398 6041
rect 249 6014 367 6034
rect 387 6014 398 6034
rect 249 6006 398 6014
rect 465 6038 824 6042
rect 465 6033 787 6038
rect 465 6009 578 6033
rect 602 6014 787 6033
rect 811 6014 824 6038
rect 602 6009 824 6014
rect 465 6006 824 6009
rect 886 6006 921 6043
rect 989 6040 1089 6043
rect 989 6036 1056 6040
rect 989 6010 1001 6036
rect 1027 6014 1056 6036
rect 1082 6014 1089 6040
rect 1027 6010 1089 6014
rect 989 6006 1089 6010
rect 465 5985 496 6006
rect 886 5985 922 6006
rect 308 5984 345 5985
rect 307 5975 345 5984
rect 307 5955 316 5975
rect 336 5955 345 5975
rect 307 5947 345 5955
rect 411 5979 496 5985
rect 521 5984 558 5985
rect 411 5959 419 5979
rect 439 5959 496 5979
rect 411 5951 496 5959
rect 520 5975 558 5984
rect 520 5955 529 5975
rect 549 5955 558 5975
rect 411 5950 447 5951
rect 520 5947 558 5955
rect 624 5979 709 5985
rect 729 5984 766 5985
rect 624 5959 632 5979
rect 652 5978 709 5979
rect 652 5959 681 5978
rect 624 5958 681 5959
rect 702 5958 709 5978
rect 624 5951 709 5958
rect 728 5975 766 5984
rect 728 5955 737 5975
rect 757 5955 766 5975
rect 624 5950 660 5951
rect 728 5947 766 5955
rect 832 5980 976 5985
rect 832 5979 897 5980
rect 832 5959 840 5979
rect 860 5959 897 5979
rect 919 5979 976 5980
rect 919 5959 948 5979
rect 968 5959 976 5979
rect 832 5951 976 5959
rect 832 5950 868 5951
rect 940 5950 976 5951
rect 1042 5984 1079 5985
rect 1042 5983 1080 5984
rect 1042 5975 1106 5983
rect 1042 5955 1051 5975
rect 1071 5961 1106 5975
rect 1126 5961 1129 5981
rect 1071 5956 1129 5961
rect 1071 5955 1106 5956
rect 308 5918 345 5947
rect 309 5916 345 5918
rect 521 5916 558 5947
rect 309 5894 558 5916
rect 729 5915 766 5947
rect 1042 5943 1106 5955
rect 1146 5917 1173 6095
rect 1005 5915 1173 5917
rect 729 5889 1173 5915
rect 1325 6014 1575 6038
rect 1325 5943 1362 6014
rect 1477 5953 1508 5954
rect 1325 5923 1334 5943
rect 1354 5923 1362 5943
rect 1325 5913 1362 5923
rect 1421 5943 1508 5953
rect 1421 5923 1430 5943
rect 1450 5923 1508 5943
rect 1421 5914 1508 5923
rect 1421 5913 1458 5914
rect 729 5879 751 5889
rect 1005 5888 1173 5889
rect 689 5877 751 5879
rect 119 5870 751 5877
rect 118 5861 751 5870
rect 1477 5861 1508 5914
rect 1538 5943 1575 6014
rect 1746 6019 2139 6039
rect 2159 6019 2162 6039
rect 1746 6014 2162 6019
rect 1746 6013 2087 6014
rect 1690 5953 1721 5954
rect 1538 5923 1547 5943
rect 1567 5923 1575 5943
rect 1538 5913 1575 5923
rect 1634 5946 1721 5953
rect 1634 5943 1695 5946
rect 1634 5923 1643 5943
rect 1663 5926 1695 5943
rect 1716 5926 1721 5946
rect 1663 5923 1721 5926
rect 1634 5916 1721 5923
rect 1746 5943 1783 6013
rect 2049 6012 2086 6013
rect 1898 5953 1934 5954
rect 1746 5923 1755 5943
rect 1775 5923 1783 5943
rect 1634 5914 1690 5916
rect 1634 5913 1671 5914
rect 1746 5913 1783 5923
rect 1842 5943 1990 5953
rect 2090 5950 2186 5952
rect 1842 5923 1851 5943
rect 1871 5923 1961 5943
rect 1981 5923 1990 5943
rect 1842 5914 1990 5923
rect 2048 5943 2186 5950
rect 2048 5923 2057 5943
rect 2077 5923 2186 5943
rect 2048 5914 2186 5923
rect 1842 5913 1879 5914
rect 1898 5862 1934 5914
rect 1953 5913 1990 5914
rect 2049 5913 2086 5914
rect 118 5843 128 5861
rect 146 5860 751 5861
rect 1369 5860 1410 5861
rect 146 5855 167 5860
rect 146 5843 158 5855
rect 1261 5853 1410 5860
rect 118 5835 158 5843
rect 201 5842 227 5843
rect 118 5833 155 5835
rect 201 5824 755 5842
rect 1261 5833 1379 5853
rect 1399 5833 1410 5853
rect 1261 5825 1410 5833
rect 1477 5857 1836 5861
rect 1477 5852 1799 5857
rect 1477 5828 1590 5852
rect 1614 5833 1799 5852
rect 1823 5833 1836 5857
rect 1614 5828 1836 5833
rect 1477 5825 1836 5828
rect 1898 5825 1933 5862
rect 2001 5859 2101 5862
rect 2001 5855 2068 5859
rect 2001 5829 2013 5855
rect 2039 5833 2068 5855
rect 2094 5833 2101 5859
rect 2039 5829 2101 5833
rect 2001 5825 2101 5829
rect 121 5765 158 5771
rect 201 5765 227 5824
rect 734 5805 755 5824
rect 121 5762 227 5765
rect 121 5744 130 5762
rect 148 5748 227 5762
rect 312 5780 562 5804
rect 148 5746 224 5748
rect 148 5744 158 5746
rect 121 5734 158 5744
rect 126 5669 157 5734
rect 312 5709 349 5780
rect 464 5719 495 5720
rect 312 5689 321 5709
rect 341 5689 349 5709
rect 312 5679 349 5689
rect 408 5709 495 5719
rect 408 5689 417 5709
rect 437 5689 495 5709
rect 408 5680 495 5689
rect 408 5679 445 5680
rect 125 5660 162 5669
rect 125 5642 135 5660
rect 153 5642 162 5660
rect 125 5632 162 5642
rect 464 5627 495 5680
rect 525 5709 562 5780
rect 733 5785 1126 5805
rect 1146 5785 1149 5805
rect 1477 5804 1508 5825
rect 1898 5804 1934 5825
rect 1320 5803 1357 5804
rect 733 5780 1149 5785
rect 1319 5794 1357 5803
rect 733 5779 1074 5780
rect 677 5719 708 5720
rect 525 5689 534 5709
rect 554 5689 562 5709
rect 525 5679 562 5689
rect 621 5712 708 5719
rect 621 5709 682 5712
rect 621 5689 630 5709
rect 650 5692 682 5709
rect 703 5692 708 5712
rect 650 5689 708 5692
rect 621 5682 708 5689
rect 733 5709 770 5779
rect 1036 5778 1073 5779
rect 1319 5774 1328 5794
rect 1348 5774 1357 5794
rect 1319 5766 1357 5774
rect 1423 5798 1508 5804
rect 1533 5803 1570 5804
rect 1423 5778 1431 5798
rect 1451 5778 1508 5798
rect 1423 5770 1508 5778
rect 1532 5794 1570 5803
rect 1532 5774 1541 5794
rect 1561 5774 1570 5794
rect 1423 5769 1459 5770
rect 1532 5766 1570 5774
rect 1636 5798 1721 5804
rect 1741 5803 1778 5804
rect 1636 5778 1644 5798
rect 1664 5797 1721 5798
rect 1664 5778 1693 5797
rect 1636 5777 1693 5778
rect 1714 5777 1721 5797
rect 1636 5770 1721 5777
rect 1740 5794 1778 5803
rect 1740 5774 1749 5794
rect 1769 5774 1778 5794
rect 1636 5769 1672 5770
rect 1740 5766 1778 5774
rect 1844 5798 1988 5804
rect 1844 5778 1852 5798
rect 1872 5778 1904 5798
rect 1928 5778 1960 5798
rect 1980 5778 1988 5798
rect 1844 5770 1988 5778
rect 1844 5769 1880 5770
rect 1952 5769 1988 5770
rect 2054 5803 2091 5804
rect 2054 5802 2092 5803
rect 2054 5794 2118 5802
rect 2054 5774 2063 5794
rect 2083 5780 2118 5794
rect 2138 5780 2141 5800
rect 2083 5775 2141 5780
rect 2083 5774 2118 5775
rect 1320 5737 1357 5766
rect 1321 5735 1357 5737
rect 1533 5735 1570 5766
rect 885 5719 921 5720
rect 733 5689 742 5709
rect 762 5689 770 5709
rect 621 5680 677 5682
rect 621 5679 658 5680
rect 733 5679 770 5689
rect 829 5709 977 5719
rect 1077 5716 1173 5718
rect 829 5689 838 5709
rect 858 5689 948 5709
rect 968 5689 977 5709
rect 829 5680 977 5689
rect 1035 5709 1173 5716
rect 1321 5713 1570 5735
rect 1741 5734 1778 5766
rect 2054 5762 2118 5774
rect 2158 5736 2185 5914
rect 2017 5734 2185 5736
rect 1741 5730 2185 5734
rect 1035 5689 1044 5709
rect 1064 5689 1173 5709
rect 1741 5711 1790 5730
rect 1810 5711 2185 5730
rect 1741 5708 2185 5711
rect 2017 5707 2185 5708
rect 1035 5680 1173 5689
rect 829 5679 866 5680
rect 885 5628 921 5680
rect 940 5679 977 5680
rect 1036 5679 1073 5680
rect 356 5626 397 5627
rect 248 5619 397 5626
rect 248 5599 366 5619
rect 386 5599 397 5619
rect 248 5591 397 5599
rect 464 5623 823 5627
rect 464 5618 786 5623
rect 464 5594 577 5618
rect 601 5599 786 5618
rect 810 5599 823 5623
rect 601 5594 823 5599
rect 464 5591 823 5594
rect 885 5591 920 5628
rect 988 5625 1088 5628
rect 988 5621 1055 5625
rect 988 5595 1000 5621
rect 1026 5599 1055 5621
rect 1081 5599 1088 5625
rect 1026 5595 1088 5599
rect 988 5591 1088 5595
rect 464 5570 495 5591
rect 885 5570 921 5591
rect 128 5561 165 5570
rect 307 5569 344 5570
rect 128 5543 137 5561
rect 155 5543 165 5561
rect 128 5533 165 5543
rect 129 5498 165 5533
rect 306 5560 344 5569
rect 306 5540 315 5560
rect 335 5540 344 5560
rect 306 5532 344 5540
rect 410 5564 495 5570
rect 520 5569 557 5570
rect 410 5544 418 5564
rect 438 5544 495 5564
rect 410 5536 495 5544
rect 519 5560 557 5569
rect 519 5540 528 5560
rect 548 5540 557 5560
rect 410 5535 446 5536
rect 519 5532 557 5540
rect 623 5564 708 5570
rect 728 5569 765 5570
rect 623 5544 631 5564
rect 651 5563 708 5564
rect 651 5544 680 5563
rect 623 5543 680 5544
rect 701 5543 708 5563
rect 623 5536 708 5543
rect 727 5560 765 5569
rect 727 5540 736 5560
rect 756 5540 765 5560
rect 623 5535 659 5536
rect 727 5532 765 5540
rect 831 5564 975 5570
rect 831 5544 839 5564
rect 859 5563 947 5564
rect 859 5544 887 5563
rect 831 5542 887 5544
rect 909 5544 947 5563
rect 967 5544 975 5564
rect 909 5542 975 5544
rect 831 5536 975 5542
rect 831 5535 867 5536
rect 939 5535 975 5536
rect 1041 5569 1078 5570
rect 1041 5568 1079 5569
rect 1041 5560 1105 5568
rect 1041 5540 1050 5560
rect 1070 5546 1105 5560
rect 1125 5546 1128 5566
rect 1070 5541 1128 5546
rect 1070 5540 1105 5541
rect 307 5503 344 5532
rect 127 5457 165 5498
rect 308 5501 344 5503
rect 520 5501 557 5532
rect 308 5479 557 5501
rect 728 5500 765 5532
rect 1041 5528 1105 5540
rect 1145 5502 1172 5680
rect 1004 5500 1172 5502
rect 728 5474 1172 5500
rect 729 5457 753 5474
rect 1004 5473 1172 5474
rect 127 5439 754 5457
rect 1380 5453 1630 5477
rect 127 5433 165 5439
rect 127 5409 164 5433
rect 127 5385 162 5409
rect 125 5376 162 5385
rect 125 5358 135 5376
rect 153 5358 162 5376
rect 125 5348 162 5358
rect 1380 5382 1417 5453
rect 1532 5392 1563 5393
rect 1380 5362 1389 5382
rect 1409 5362 1417 5382
rect 1380 5352 1417 5362
rect 1476 5382 1563 5392
rect 1476 5362 1485 5382
rect 1505 5362 1563 5382
rect 1476 5353 1563 5362
rect 1476 5352 1513 5353
rect 1532 5300 1563 5353
rect 1593 5382 1630 5453
rect 1801 5458 2194 5478
rect 2214 5458 2217 5478
rect 1801 5453 2217 5458
rect 1801 5452 2142 5453
rect 1745 5392 1776 5393
rect 1593 5362 1602 5382
rect 1622 5362 1630 5382
rect 1593 5352 1630 5362
rect 1689 5385 1776 5392
rect 1689 5382 1750 5385
rect 1689 5362 1698 5382
rect 1718 5365 1750 5382
rect 1771 5365 1776 5385
rect 1718 5362 1776 5365
rect 1689 5355 1776 5362
rect 1801 5382 1838 5452
rect 2104 5451 2141 5452
rect 1953 5392 1989 5393
rect 1801 5362 1810 5382
rect 1830 5362 1838 5382
rect 1689 5353 1745 5355
rect 1689 5352 1726 5353
rect 1801 5352 1838 5362
rect 1897 5382 2045 5392
rect 2145 5389 2241 5391
rect 1897 5362 1906 5382
rect 1926 5362 2016 5382
rect 2036 5362 2045 5382
rect 1897 5353 2045 5362
rect 2103 5382 2241 5389
rect 2103 5362 2112 5382
rect 2132 5362 2241 5382
rect 2103 5353 2241 5362
rect 1897 5352 1934 5353
rect 1953 5301 1989 5353
rect 2008 5352 2045 5353
rect 2104 5352 2141 5353
rect 1424 5299 1465 5300
rect 1316 5292 1465 5299
rect 128 5284 165 5286
rect 128 5283 776 5284
rect 127 5277 776 5283
rect 127 5259 137 5277
rect 155 5263 776 5277
rect 1316 5272 1434 5292
rect 1454 5272 1465 5292
rect 1316 5264 1465 5272
rect 1532 5296 1891 5300
rect 1532 5291 1854 5296
rect 1532 5267 1645 5291
rect 1669 5272 1854 5291
rect 1878 5272 1891 5296
rect 1669 5267 1891 5272
rect 1532 5264 1891 5267
rect 1953 5264 1988 5301
rect 2056 5298 2156 5301
rect 2056 5294 2123 5298
rect 2056 5268 2068 5294
rect 2094 5272 2123 5294
rect 2149 5272 2156 5298
rect 2094 5268 2156 5272
rect 2056 5264 2156 5268
rect 155 5259 165 5263
rect 606 5262 776 5263
rect 127 5249 165 5259
rect 127 5171 162 5249
rect 739 5239 776 5262
rect 1532 5243 1563 5264
rect 1953 5243 1989 5264
rect 1375 5242 1412 5243
rect 123 5162 162 5171
rect 123 5144 133 5162
rect 151 5144 162 5162
rect 123 5138 162 5144
rect 318 5214 568 5238
rect 318 5143 355 5214
rect 470 5153 501 5154
rect 123 5134 160 5138
rect 318 5123 327 5143
rect 347 5123 355 5143
rect 318 5113 355 5123
rect 414 5143 501 5153
rect 414 5123 423 5143
rect 443 5123 501 5143
rect 414 5114 501 5123
rect 414 5113 451 5114
rect 126 5063 163 5072
rect 124 5045 135 5063
rect 153 5045 163 5063
rect 470 5061 501 5114
rect 531 5143 568 5214
rect 739 5219 1132 5239
rect 1152 5219 1155 5239
rect 739 5214 1155 5219
rect 1374 5233 1412 5242
rect 739 5213 1080 5214
rect 1374 5213 1383 5233
rect 1403 5213 1412 5233
rect 683 5153 714 5154
rect 531 5123 540 5143
rect 560 5123 568 5143
rect 531 5113 568 5123
rect 627 5146 714 5153
rect 627 5143 688 5146
rect 627 5123 636 5143
rect 656 5126 688 5143
rect 709 5126 714 5146
rect 656 5123 714 5126
rect 627 5116 714 5123
rect 739 5143 776 5213
rect 1042 5212 1079 5213
rect 1374 5205 1412 5213
rect 1478 5237 1563 5243
rect 1588 5242 1625 5243
rect 1478 5217 1486 5237
rect 1506 5217 1563 5237
rect 1478 5209 1563 5217
rect 1587 5233 1625 5242
rect 1587 5213 1596 5233
rect 1616 5213 1625 5233
rect 1478 5208 1514 5209
rect 1587 5205 1625 5213
rect 1691 5237 1776 5243
rect 1796 5242 1833 5243
rect 1691 5217 1699 5237
rect 1719 5236 1776 5237
rect 1719 5217 1748 5236
rect 1691 5216 1748 5217
rect 1769 5216 1776 5236
rect 1691 5209 1776 5216
rect 1795 5233 1833 5242
rect 1795 5213 1804 5233
rect 1824 5213 1833 5233
rect 1691 5208 1727 5209
rect 1795 5205 1833 5213
rect 1899 5237 2043 5243
rect 1899 5217 1907 5237
rect 1927 5236 2015 5237
rect 1927 5217 1960 5236
rect 1983 5217 2015 5236
rect 2035 5217 2043 5237
rect 1899 5209 2043 5217
rect 1899 5208 1935 5209
rect 2007 5208 2043 5209
rect 2109 5242 2146 5243
rect 2109 5241 2147 5242
rect 2109 5233 2173 5241
rect 2109 5213 2118 5233
rect 2138 5219 2173 5233
rect 2193 5219 2196 5239
rect 2138 5214 2196 5219
rect 2138 5213 2173 5214
rect 1375 5176 1412 5205
rect 1376 5174 1412 5176
rect 1588 5174 1625 5205
rect 891 5153 927 5154
rect 739 5123 748 5143
rect 768 5123 776 5143
rect 627 5114 683 5116
rect 627 5113 664 5114
rect 739 5113 776 5123
rect 835 5143 983 5153
rect 1376 5152 1625 5174
rect 1796 5173 1833 5205
rect 2109 5201 2173 5213
rect 2213 5175 2240 5353
rect 2072 5173 2240 5175
rect 1796 5162 2240 5173
rect 2303 5173 2333 6174
rect 2303 5168 2335 5173
rect 1083 5150 1179 5152
rect 835 5123 844 5143
rect 864 5123 954 5143
rect 974 5123 983 5143
rect 835 5114 983 5123
rect 1041 5143 1179 5150
rect 1796 5147 2242 5162
rect 2072 5146 2242 5147
rect 1041 5123 1050 5143
rect 1070 5123 1179 5143
rect 1041 5114 1179 5123
rect 835 5113 872 5114
rect 891 5062 927 5114
rect 946 5113 983 5114
rect 1042 5113 1079 5114
rect 362 5060 403 5061
rect 124 4896 163 5045
rect 254 5053 403 5060
rect 254 5033 372 5053
rect 392 5033 403 5053
rect 254 5025 403 5033
rect 470 5057 829 5061
rect 470 5052 792 5057
rect 470 5028 583 5052
rect 607 5033 792 5052
rect 816 5033 829 5057
rect 607 5028 829 5033
rect 470 5025 829 5028
rect 891 5025 926 5062
rect 994 5059 1094 5062
rect 994 5055 1061 5059
rect 994 5029 1006 5055
rect 1032 5033 1061 5055
rect 1087 5033 1094 5059
rect 1032 5029 1094 5033
rect 994 5025 1094 5029
rect 470 5004 501 5025
rect 891 5004 927 5025
rect 313 5003 350 5004
rect 312 4994 350 5003
rect 312 4974 321 4994
rect 341 4974 350 4994
rect 312 4966 350 4974
rect 416 4998 501 5004
rect 526 5003 563 5004
rect 416 4978 424 4998
rect 444 4978 501 4998
rect 416 4970 501 4978
rect 525 4994 563 5003
rect 525 4974 534 4994
rect 554 4974 563 4994
rect 416 4969 452 4970
rect 525 4966 563 4974
rect 629 4998 714 5004
rect 734 5003 771 5004
rect 629 4978 637 4998
rect 657 4997 714 4998
rect 657 4978 686 4997
rect 629 4977 686 4978
rect 707 4977 714 4997
rect 629 4970 714 4977
rect 733 4994 771 5003
rect 733 4974 742 4994
rect 762 4974 771 4994
rect 629 4969 665 4970
rect 733 4966 771 4974
rect 837 4999 981 5004
rect 837 4998 902 4999
rect 837 4978 845 4998
rect 865 4978 902 4998
rect 924 4998 981 4999
rect 924 4978 953 4998
rect 973 4978 981 4998
rect 837 4970 981 4978
rect 837 4969 873 4970
rect 945 4969 981 4970
rect 1047 5003 1084 5004
rect 1047 5002 1085 5003
rect 1047 4994 1111 5002
rect 1047 4974 1056 4994
rect 1076 4980 1111 4994
rect 1131 4980 1134 5000
rect 1076 4975 1134 4980
rect 1076 4974 1111 4975
rect 313 4937 350 4966
rect 314 4935 350 4937
rect 526 4935 563 4966
rect 314 4913 563 4935
rect 734 4934 771 4966
rect 1047 4962 1111 4974
rect 1151 4936 1178 5114
rect 1010 4934 1178 4936
rect 734 4908 1178 4934
rect 1330 5033 1580 5057
rect 1330 4962 1367 5033
rect 1482 4972 1513 4973
rect 1330 4942 1339 4962
rect 1359 4942 1367 4962
rect 1330 4932 1367 4942
rect 1426 4962 1513 4972
rect 1426 4942 1435 4962
rect 1455 4942 1513 4962
rect 1426 4933 1513 4942
rect 1426 4932 1463 4933
rect 734 4898 756 4908
rect 1010 4907 1178 4908
rect 694 4896 756 4898
rect 124 4889 756 4896
rect 123 4880 756 4889
rect 1482 4880 1513 4933
rect 1543 4962 1580 5033
rect 1751 5038 2144 5058
rect 2164 5038 2167 5058
rect 1751 5033 2167 5038
rect 1751 5032 2092 5033
rect 1695 4972 1726 4973
rect 1543 4942 1552 4962
rect 1572 4942 1580 4962
rect 1543 4932 1580 4942
rect 1639 4965 1726 4972
rect 1639 4962 1700 4965
rect 1639 4942 1648 4962
rect 1668 4945 1700 4962
rect 1721 4945 1726 4965
rect 1668 4942 1726 4945
rect 1639 4935 1726 4942
rect 1751 4962 1788 5032
rect 2054 5031 2091 5032
rect 1903 4972 1939 4973
rect 1751 4942 1760 4962
rect 1780 4942 1788 4962
rect 1639 4933 1695 4935
rect 1639 4932 1676 4933
rect 1751 4932 1788 4942
rect 1847 4962 1995 4972
rect 2095 4969 2191 4971
rect 1847 4942 1856 4962
rect 1876 4942 1966 4962
rect 1986 4942 1995 4962
rect 1847 4933 1995 4942
rect 2053 4962 2191 4969
rect 2053 4942 2062 4962
rect 2082 4942 2191 4962
rect 2053 4933 2191 4942
rect 1847 4932 1884 4933
rect 1903 4881 1939 4933
rect 1958 4932 1995 4933
rect 2054 4932 2091 4933
rect 123 4862 133 4880
rect 151 4879 756 4880
rect 1374 4879 1415 4880
rect 151 4874 172 4879
rect 151 4862 163 4874
rect 1266 4872 1415 4879
rect 123 4854 163 4862
rect 206 4861 232 4862
rect 123 4852 160 4854
rect 206 4843 760 4861
rect 1266 4852 1384 4872
rect 1404 4852 1415 4872
rect 1266 4844 1415 4852
rect 1482 4876 1841 4880
rect 1482 4871 1804 4876
rect 1482 4847 1595 4871
rect 1619 4852 1804 4871
rect 1828 4852 1841 4876
rect 1619 4847 1841 4852
rect 1482 4844 1841 4847
rect 1903 4844 1938 4881
rect 2006 4878 2106 4881
rect 2006 4874 2073 4878
rect 2006 4848 2018 4874
rect 2044 4852 2073 4874
rect 2099 4852 2106 4878
rect 2044 4848 2106 4852
rect 2006 4844 2106 4848
rect 126 4784 163 4790
rect 206 4784 232 4843
rect 739 4824 760 4843
rect 126 4781 232 4784
rect 126 4763 135 4781
rect 153 4767 232 4781
rect 317 4799 567 4823
rect 153 4765 229 4767
rect 153 4763 163 4765
rect 126 4753 163 4763
rect 131 4688 162 4753
rect 317 4728 354 4799
rect 469 4738 500 4739
rect 317 4708 326 4728
rect 346 4708 354 4728
rect 317 4698 354 4708
rect 413 4728 500 4738
rect 413 4708 422 4728
rect 442 4708 500 4728
rect 413 4699 500 4708
rect 413 4698 450 4699
rect 130 4679 167 4688
rect 130 4661 140 4679
rect 158 4661 167 4679
rect 130 4651 167 4661
rect 469 4646 500 4699
rect 530 4728 567 4799
rect 738 4804 1131 4824
rect 1151 4804 1154 4824
rect 1482 4823 1513 4844
rect 1903 4823 1939 4844
rect 1325 4822 1362 4823
rect 738 4799 1154 4804
rect 1324 4813 1362 4822
rect 738 4798 1079 4799
rect 682 4738 713 4739
rect 530 4708 539 4728
rect 559 4708 567 4728
rect 530 4698 567 4708
rect 626 4731 713 4738
rect 626 4728 687 4731
rect 626 4708 635 4728
rect 655 4711 687 4728
rect 708 4711 713 4731
rect 655 4708 713 4711
rect 626 4701 713 4708
rect 738 4728 775 4798
rect 1041 4797 1078 4798
rect 1324 4793 1333 4813
rect 1353 4793 1362 4813
rect 1324 4785 1362 4793
rect 1428 4817 1513 4823
rect 1538 4822 1575 4823
rect 1428 4797 1436 4817
rect 1456 4797 1513 4817
rect 1428 4789 1513 4797
rect 1537 4813 1575 4822
rect 1537 4793 1546 4813
rect 1566 4793 1575 4813
rect 1428 4788 1464 4789
rect 1537 4785 1575 4793
rect 1641 4817 1726 4823
rect 1746 4822 1783 4823
rect 1641 4797 1649 4817
rect 1669 4816 1726 4817
rect 1669 4797 1698 4816
rect 1641 4796 1698 4797
rect 1719 4796 1726 4816
rect 1641 4789 1726 4796
rect 1745 4813 1783 4822
rect 1745 4793 1754 4813
rect 1774 4793 1783 4813
rect 1641 4788 1677 4789
rect 1745 4785 1783 4793
rect 1849 4818 1993 4823
rect 1849 4817 1908 4818
rect 1849 4797 1857 4817
rect 1877 4798 1908 4817
rect 1932 4817 1993 4818
rect 1932 4798 1965 4817
rect 1877 4797 1965 4798
rect 1985 4797 1993 4817
rect 1849 4789 1993 4797
rect 1849 4788 1885 4789
rect 1957 4788 1993 4789
rect 2059 4822 2096 4823
rect 2059 4821 2097 4822
rect 2059 4813 2123 4821
rect 2059 4793 2068 4813
rect 2088 4799 2123 4813
rect 2143 4799 2146 4819
rect 2088 4794 2146 4799
rect 2088 4793 2123 4794
rect 1325 4756 1362 4785
rect 1326 4754 1362 4756
rect 1538 4754 1575 4785
rect 890 4738 926 4739
rect 738 4708 747 4728
rect 767 4708 775 4728
rect 626 4699 682 4701
rect 626 4698 663 4699
rect 738 4698 775 4708
rect 834 4728 982 4738
rect 1082 4735 1178 4737
rect 834 4708 843 4728
rect 863 4708 953 4728
rect 973 4708 982 4728
rect 834 4699 982 4708
rect 1040 4728 1178 4735
rect 1326 4732 1575 4754
rect 1746 4753 1783 4785
rect 2059 4781 2123 4793
rect 2163 4755 2190 4933
rect 2022 4753 2190 4755
rect 1746 4749 2190 4753
rect 1040 4708 1049 4728
rect 1069 4708 1178 4728
rect 1746 4730 1795 4749
rect 1815 4730 2190 4749
rect 1746 4727 2190 4730
rect 2022 4726 2190 4727
rect 2211 4752 2242 5146
rect 2303 5150 2308 5168
rect 2328 5150 2335 5168
rect 2303 5145 2335 5150
rect 2306 5143 2335 5145
rect 2211 4726 2216 4752
rect 2235 4726 2242 4752
rect 2749 4727 2787 6558
rect 2815 6445 2842 6623
rect 2882 6585 2946 6597
rect 3222 6593 3259 6625
rect 3430 6624 3679 6646
rect 4134 6632 4171 6633
rect 4437 6632 4474 6702
rect 4499 6722 4586 6729
rect 4499 6719 4557 6722
rect 4499 6699 4504 6719
rect 4525 6702 4557 6719
rect 4577 6702 4586 6722
rect 4525 6699 4586 6702
rect 4499 6692 4586 6699
rect 4645 6722 4682 6732
rect 4645 6702 4653 6722
rect 4673 6702 4682 6722
rect 4499 6691 4530 6692
rect 4133 6631 4474 6632
rect 3430 6593 3467 6624
rect 3643 6622 3679 6624
rect 4058 6626 4474 6631
rect 3643 6593 3680 6622
rect 4058 6606 4061 6626
rect 4081 6606 4474 6626
rect 4645 6631 4682 6702
rect 4712 6731 4743 6784
rect 5050 6782 5060 6800
rect 5078 6782 5089 6800
rect 5392 6819 6025 6828
rect 6751 6819 6782 6872
rect 6812 6901 6849 6972
rect 7020 6977 7413 6997
rect 7433 6977 7436 6997
rect 7020 6972 7436 6977
rect 7020 6971 7361 6972
rect 6964 6911 6995 6912
rect 6812 6881 6821 6901
rect 6841 6881 6849 6901
rect 6812 6871 6849 6881
rect 6908 6904 6995 6911
rect 6908 6901 6969 6904
rect 6908 6881 6917 6901
rect 6937 6884 6969 6901
rect 6990 6884 6995 6904
rect 6937 6881 6995 6884
rect 6908 6874 6995 6881
rect 7020 6901 7057 6971
rect 7323 6970 7360 6971
rect 7172 6911 7208 6912
rect 7020 6881 7029 6901
rect 7049 6881 7057 6901
rect 6908 6872 6964 6874
rect 6908 6871 6945 6872
rect 7020 6871 7057 6881
rect 7116 6901 7264 6911
rect 7364 6908 7460 6910
rect 7116 6881 7125 6901
rect 7145 6881 7235 6901
rect 7255 6881 7264 6901
rect 7116 6872 7264 6881
rect 7322 6901 7460 6908
rect 7322 6881 7331 6901
rect 7351 6881 7460 6901
rect 7322 6872 7460 6881
rect 7116 6871 7153 6872
rect 7172 6820 7208 6872
rect 7227 6871 7264 6872
rect 7323 6871 7360 6872
rect 5392 6801 5402 6819
rect 5420 6818 6025 6819
rect 6643 6818 6684 6819
rect 5420 6813 5441 6818
rect 5420 6801 5432 6813
rect 6535 6811 6684 6818
rect 5392 6793 5432 6801
rect 5475 6800 5501 6801
rect 5392 6791 5429 6793
rect 5475 6782 6029 6800
rect 6535 6791 6653 6811
rect 6673 6791 6684 6811
rect 6535 6783 6684 6791
rect 6751 6815 7110 6819
rect 6751 6810 7073 6815
rect 6751 6786 6864 6810
rect 6888 6791 7073 6810
rect 7097 6791 7110 6815
rect 6888 6786 7110 6791
rect 6751 6783 7110 6786
rect 7172 6783 7207 6820
rect 7275 6817 7375 6820
rect 7275 6813 7342 6817
rect 7275 6787 7287 6813
rect 7313 6791 7342 6813
rect 7368 6791 7375 6817
rect 7313 6787 7375 6791
rect 7275 6783 7375 6787
rect 5050 6773 5087 6782
rect 4762 6731 4799 6732
rect 4712 6722 4799 6731
rect 4712 6702 4770 6722
rect 4790 6702 4799 6722
rect 4712 6692 4799 6702
rect 4858 6722 4895 6732
rect 4858 6702 4866 6722
rect 4886 6702 4895 6722
rect 5395 6723 5432 6729
rect 5475 6723 5501 6782
rect 6008 6763 6029 6782
rect 5395 6720 5501 6723
rect 5053 6707 5090 6711
rect 4712 6691 4743 6692
rect 4858 6631 4895 6702
rect 4645 6607 4895 6631
rect 5051 6701 5090 6707
rect 5051 6683 5062 6701
rect 5080 6683 5090 6701
rect 5395 6702 5404 6720
rect 5422 6706 5501 6720
rect 5586 6738 5836 6762
rect 5422 6704 5498 6706
rect 5422 6702 5432 6704
rect 5395 6692 5432 6702
rect 5051 6674 5090 6683
rect 2882 6584 2917 6585
rect 2859 6579 2917 6584
rect 2859 6559 2862 6579
rect 2882 6565 2917 6579
rect 2937 6565 2946 6585
rect 2882 6557 2946 6565
rect 2908 6556 2946 6557
rect 2909 6555 2946 6556
rect 3012 6589 3048 6590
rect 3120 6589 3156 6590
rect 3012 6581 3156 6589
rect 3012 6561 3020 6581
rect 3040 6580 3128 6581
rect 3040 6561 3069 6580
rect 3092 6561 3128 6580
rect 3148 6561 3156 6581
rect 3012 6555 3156 6561
rect 3222 6585 3260 6593
rect 3328 6589 3364 6590
rect 3222 6565 3231 6585
rect 3251 6565 3260 6585
rect 3222 6556 3260 6565
rect 3279 6582 3364 6589
rect 3279 6562 3286 6582
rect 3307 6581 3364 6582
rect 3307 6562 3336 6581
rect 3279 6561 3336 6562
rect 3356 6561 3364 6581
rect 3222 6555 3259 6556
rect 3279 6555 3364 6561
rect 3430 6585 3468 6593
rect 3541 6589 3577 6590
rect 3430 6565 3439 6585
rect 3459 6565 3468 6585
rect 3430 6556 3468 6565
rect 3492 6581 3577 6589
rect 3492 6561 3549 6581
rect 3569 6561 3577 6581
rect 3430 6555 3467 6556
rect 3492 6555 3577 6561
rect 3643 6585 3681 6593
rect 3643 6565 3652 6585
rect 3672 6565 3681 6585
rect 3643 6556 3681 6565
rect 4437 6583 4474 6606
rect 5051 6596 5086 6674
rect 5400 6627 5431 6692
rect 5586 6667 5623 6738
rect 5738 6677 5769 6678
rect 5586 6647 5595 6667
rect 5615 6647 5623 6667
rect 5586 6637 5623 6647
rect 5682 6667 5769 6677
rect 5682 6647 5691 6667
rect 5711 6647 5769 6667
rect 5682 6638 5769 6647
rect 5682 6637 5719 6638
rect 5048 6586 5086 6596
rect 5399 6618 5436 6627
rect 5399 6600 5409 6618
rect 5427 6600 5436 6618
rect 5399 6590 5436 6600
rect 4437 6582 4607 6583
rect 5048 6582 5058 6586
rect 4437 6568 5058 6582
rect 5076 6568 5086 6586
rect 5738 6585 5769 6638
rect 5799 6667 5836 6738
rect 6007 6743 6400 6763
rect 6420 6743 6423 6763
rect 6751 6762 6782 6783
rect 7172 6762 7208 6783
rect 6594 6761 6631 6762
rect 6007 6738 6423 6743
rect 6593 6752 6631 6761
rect 6007 6737 6348 6738
rect 5951 6677 5982 6678
rect 5799 6647 5808 6667
rect 5828 6647 5836 6667
rect 5799 6637 5836 6647
rect 5895 6670 5982 6677
rect 5895 6667 5956 6670
rect 5895 6647 5904 6667
rect 5924 6650 5956 6667
rect 5977 6650 5982 6670
rect 5924 6647 5982 6650
rect 5895 6640 5982 6647
rect 6007 6667 6044 6737
rect 6310 6736 6347 6737
rect 6593 6732 6602 6752
rect 6622 6732 6631 6752
rect 6593 6724 6631 6732
rect 6697 6756 6782 6762
rect 6807 6761 6844 6762
rect 6697 6736 6705 6756
rect 6725 6736 6782 6756
rect 6697 6728 6782 6736
rect 6806 6752 6844 6761
rect 6806 6732 6815 6752
rect 6835 6732 6844 6752
rect 6697 6727 6733 6728
rect 6806 6724 6844 6732
rect 6910 6756 6995 6762
rect 7015 6761 7052 6762
rect 6910 6736 6918 6756
rect 6938 6755 6995 6756
rect 6938 6736 6967 6755
rect 6910 6735 6967 6736
rect 6988 6735 6995 6755
rect 6910 6728 6995 6735
rect 7014 6752 7052 6761
rect 7014 6732 7023 6752
rect 7043 6732 7052 6752
rect 6910 6727 6946 6728
rect 7014 6724 7052 6732
rect 7118 6757 7262 6762
rect 7118 6756 7177 6757
rect 7118 6736 7126 6756
rect 7146 6737 7177 6756
rect 7201 6756 7262 6757
rect 7201 6737 7234 6756
rect 7146 6736 7234 6737
rect 7254 6736 7262 6756
rect 7118 6728 7262 6736
rect 7118 6727 7154 6728
rect 7226 6727 7262 6728
rect 7328 6761 7365 6762
rect 7328 6760 7366 6761
rect 7328 6752 7392 6760
rect 7328 6732 7337 6752
rect 7357 6738 7392 6752
rect 7412 6738 7415 6758
rect 7357 6733 7415 6738
rect 7357 6732 7392 6733
rect 6594 6695 6631 6724
rect 6595 6693 6631 6695
rect 6807 6693 6844 6724
rect 6159 6677 6195 6678
rect 6007 6647 6016 6667
rect 6036 6647 6044 6667
rect 5895 6638 5951 6640
rect 5895 6637 5932 6638
rect 6007 6637 6044 6647
rect 6103 6667 6251 6677
rect 6351 6674 6447 6676
rect 6103 6647 6112 6667
rect 6132 6647 6222 6667
rect 6242 6647 6251 6667
rect 6103 6638 6251 6647
rect 6309 6667 6447 6674
rect 6595 6671 6844 6693
rect 7015 6692 7052 6724
rect 7328 6720 7392 6732
rect 7432 6694 7459 6872
rect 7291 6692 7459 6694
rect 7015 6688 7459 6692
rect 6309 6647 6318 6667
rect 6338 6647 6447 6667
rect 7015 6669 7064 6688
rect 7084 6669 7459 6688
rect 7015 6666 7459 6669
rect 7291 6665 7459 6666
rect 7480 6691 7511 7085
rect 7480 6665 7485 6691
rect 7504 6665 7511 6691
rect 7480 6662 7511 6665
rect 6309 6638 6447 6647
rect 6103 6637 6140 6638
rect 6159 6586 6195 6638
rect 6214 6637 6251 6638
rect 6310 6637 6347 6638
rect 5630 6584 5671 6585
rect 4437 6562 5086 6568
rect 5522 6577 5671 6584
rect 4437 6561 5085 6562
rect 5048 6559 5085 6561
rect 5522 6557 5640 6577
rect 5660 6557 5671 6577
rect 3643 6555 3680 6556
rect 3066 6534 3102 6555
rect 3492 6534 3523 6555
rect 5522 6549 5671 6557
rect 5738 6581 6097 6585
rect 5738 6576 6060 6581
rect 5738 6552 5851 6576
rect 5875 6557 6060 6576
rect 6084 6557 6097 6581
rect 5875 6552 6097 6557
rect 5738 6549 6097 6552
rect 6159 6549 6194 6586
rect 6262 6583 6362 6586
rect 6262 6579 6329 6583
rect 6262 6553 6274 6579
rect 6300 6557 6329 6579
rect 6355 6557 6362 6583
rect 6300 6553 6362 6557
rect 6262 6549 6362 6553
rect 2899 6530 2999 6534
rect 2899 6526 2961 6530
rect 2899 6500 2906 6526
rect 2932 6504 2961 6526
rect 2987 6504 2999 6530
rect 2932 6500 2999 6504
rect 2899 6497 2999 6500
rect 3067 6497 3102 6534
rect 3164 6531 3523 6534
rect 3164 6526 3386 6531
rect 3164 6502 3177 6526
rect 3201 6507 3386 6526
rect 3410 6507 3523 6531
rect 3201 6502 3523 6507
rect 3164 6498 3523 6502
rect 3590 6526 3739 6534
rect 5738 6528 5769 6549
rect 6159 6528 6195 6549
rect 3590 6506 3601 6526
rect 3621 6506 3739 6526
rect 3590 6499 3739 6506
rect 5402 6519 5439 6528
rect 5581 6527 5618 6528
rect 5402 6501 5411 6519
rect 5429 6501 5439 6519
rect 3590 6498 3631 6499
rect 2914 6445 2951 6446
rect 3010 6445 3047 6446
rect 3066 6445 3102 6497
rect 3121 6445 3158 6446
rect 2814 6436 2952 6445
rect 2814 6416 2923 6436
rect 2943 6416 2952 6436
rect 2814 6409 2952 6416
rect 3010 6436 3158 6445
rect 3010 6416 3019 6436
rect 3039 6416 3129 6436
rect 3149 6416 3158 6436
rect 2814 6407 2910 6409
rect 3010 6406 3158 6416
rect 3217 6436 3254 6446
rect 3329 6445 3366 6446
rect 3310 6443 3366 6445
rect 3217 6416 3225 6436
rect 3245 6416 3254 6436
rect 3066 6405 3102 6406
rect 2914 6346 2951 6347
rect 3217 6346 3254 6416
rect 3279 6436 3366 6443
rect 3279 6433 3337 6436
rect 3279 6413 3284 6433
rect 3305 6416 3337 6433
rect 3357 6416 3366 6436
rect 3305 6413 3366 6416
rect 3279 6406 3366 6413
rect 3425 6436 3462 6446
rect 3425 6416 3433 6436
rect 3453 6416 3462 6436
rect 3279 6405 3310 6406
rect 2913 6345 3254 6346
rect 2838 6340 3254 6345
rect 2838 6320 2841 6340
rect 2861 6320 3254 6340
rect 3425 6345 3462 6416
rect 3492 6445 3523 6498
rect 5051 6487 5088 6497
rect 5402 6491 5439 6501
rect 5051 6469 5060 6487
rect 5078 6469 5088 6487
rect 5051 6460 5088 6469
rect 3542 6445 3579 6446
rect 3492 6436 3579 6445
rect 3492 6416 3550 6436
rect 3570 6416 3579 6436
rect 3492 6406 3579 6416
rect 3638 6436 3675 6446
rect 3638 6416 3646 6436
rect 3666 6416 3675 6436
rect 3492 6405 3523 6406
rect 3638 6345 3675 6416
rect 5051 6414 5086 6460
rect 5403 6456 5439 6491
rect 5580 6518 5618 6527
rect 5580 6498 5589 6518
rect 5609 6498 5618 6518
rect 5580 6490 5618 6498
rect 5684 6522 5769 6528
rect 5794 6527 5831 6528
rect 5684 6502 5692 6522
rect 5712 6502 5769 6522
rect 5684 6494 5769 6502
rect 5793 6518 5831 6527
rect 5793 6498 5802 6518
rect 5822 6498 5831 6518
rect 5684 6493 5720 6494
rect 5793 6490 5831 6498
rect 5897 6522 5982 6528
rect 6002 6527 6039 6528
rect 5897 6502 5905 6522
rect 5925 6521 5982 6522
rect 5925 6502 5954 6521
rect 5897 6501 5954 6502
rect 5975 6501 5982 6521
rect 5897 6494 5982 6501
rect 6001 6518 6039 6527
rect 6001 6498 6010 6518
rect 6030 6498 6039 6518
rect 5897 6493 5933 6494
rect 6001 6490 6039 6498
rect 6105 6522 6249 6528
rect 6105 6502 6113 6522
rect 6133 6521 6221 6522
rect 6133 6502 6161 6521
rect 6105 6500 6161 6502
rect 6183 6502 6221 6521
rect 6241 6502 6249 6522
rect 6183 6500 6249 6502
rect 6105 6494 6249 6500
rect 6105 6493 6141 6494
rect 6213 6493 6249 6494
rect 6315 6527 6352 6528
rect 6315 6526 6353 6527
rect 6315 6518 6379 6526
rect 6315 6498 6324 6518
rect 6344 6504 6379 6518
rect 6399 6504 6402 6524
rect 6344 6499 6402 6504
rect 6344 6498 6379 6499
rect 5581 6461 5618 6490
rect 5401 6415 5439 6456
rect 5582 6459 5618 6461
rect 5794 6459 5831 6490
rect 5582 6437 5831 6459
rect 6002 6458 6039 6490
rect 6315 6486 6379 6498
rect 6419 6460 6446 6638
rect 8030 6627 8067 6638
rect 8156 6631 8186 7632
rect 8249 7632 8693 7643
rect 8249 7630 8417 7632
rect 8249 7452 8276 7630
rect 8316 7592 8380 7604
rect 8656 7600 8693 7632
rect 8864 7631 9113 7653
rect 9506 7652 9654 7662
rect 9713 7682 9750 7692
rect 9825 7691 9862 7692
rect 9806 7689 9862 7691
rect 9713 7662 9721 7682
rect 9741 7662 9750 7682
rect 9562 7651 9598 7652
rect 8864 7600 8901 7631
rect 9077 7629 9113 7631
rect 9077 7600 9114 7629
rect 8316 7591 8351 7592
rect 8293 7586 8351 7591
rect 8293 7566 8296 7586
rect 8316 7572 8351 7586
rect 8371 7572 8380 7592
rect 8316 7564 8380 7572
rect 8342 7563 8380 7564
rect 8343 7562 8380 7563
rect 8446 7596 8482 7597
rect 8554 7596 8590 7597
rect 8446 7588 8590 7596
rect 8446 7568 8454 7588
rect 8474 7569 8506 7588
rect 8529 7569 8562 7588
rect 8474 7568 8562 7569
rect 8582 7568 8590 7588
rect 8446 7562 8590 7568
rect 8656 7592 8694 7600
rect 8762 7596 8798 7597
rect 8656 7572 8665 7592
rect 8685 7572 8694 7592
rect 8656 7563 8694 7572
rect 8713 7589 8798 7596
rect 8713 7569 8720 7589
rect 8741 7588 8798 7589
rect 8741 7569 8770 7588
rect 8713 7568 8770 7569
rect 8790 7568 8798 7588
rect 8656 7562 8693 7563
rect 8713 7562 8798 7568
rect 8864 7592 8902 7600
rect 8975 7596 9011 7597
rect 8864 7572 8873 7592
rect 8893 7572 8902 7592
rect 8864 7563 8902 7572
rect 8926 7588 9011 7596
rect 8926 7568 8983 7588
rect 9003 7568 9011 7588
rect 8864 7562 8901 7563
rect 8926 7562 9011 7568
rect 9077 7592 9115 7600
rect 9410 7592 9447 7593
rect 9713 7592 9750 7662
rect 9775 7682 9862 7689
rect 9775 7679 9833 7682
rect 9775 7659 9780 7679
rect 9801 7662 9833 7679
rect 9853 7662 9862 7682
rect 9801 7659 9862 7662
rect 9775 7652 9862 7659
rect 9921 7682 9958 7692
rect 9921 7662 9929 7682
rect 9949 7662 9958 7682
rect 9775 7651 9806 7652
rect 9077 7572 9086 7592
rect 9106 7572 9115 7592
rect 9409 7591 9750 7592
rect 9077 7563 9115 7572
rect 9334 7586 9750 7591
rect 9334 7566 9337 7586
rect 9357 7566 9750 7586
rect 9921 7591 9958 7662
rect 9988 7691 10019 7744
rect 10326 7742 10336 7760
rect 10354 7742 10365 7760
rect 10850 7792 11404 7810
rect 11910 7801 12028 7821
rect 12048 7801 12059 7821
rect 11910 7793 12059 7801
rect 12126 7825 12485 7829
rect 12126 7820 12448 7825
rect 12126 7796 12239 7820
rect 12263 7801 12448 7820
rect 12472 7801 12485 7825
rect 12263 7796 12485 7801
rect 12126 7793 12485 7796
rect 12547 7793 12582 7830
rect 12650 7827 12750 7830
rect 12650 7823 12717 7827
rect 12650 7797 12662 7823
rect 12688 7801 12717 7823
rect 12743 7801 12750 7827
rect 12688 7797 12750 7801
rect 12650 7793 12750 7797
rect 10326 7733 10363 7742
rect 10770 7733 10807 7739
rect 10850 7733 10876 7792
rect 11383 7773 11404 7792
rect 10770 7730 10876 7733
rect 10770 7712 10779 7730
rect 10797 7716 10876 7730
rect 10961 7748 11211 7772
rect 10797 7714 10873 7716
rect 10797 7712 10807 7714
rect 10770 7702 10807 7712
rect 10038 7691 10075 7692
rect 9988 7682 10075 7691
rect 9988 7662 10046 7682
rect 10066 7662 10075 7682
rect 9988 7652 10075 7662
rect 10134 7682 10171 7692
rect 10134 7662 10142 7682
rect 10162 7662 10171 7682
rect 10329 7667 10366 7671
rect 9988 7651 10019 7652
rect 10134 7591 10171 7662
rect 9921 7567 10171 7591
rect 10327 7661 10366 7667
rect 10327 7643 10338 7661
rect 10356 7643 10366 7661
rect 10327 7634 10366 7643
rect 10775 7637 10806 7702
rect 10961 7677 10998 7748
rect 11113 7687 11144 7688
rect 10961 7657 10970 7677
rect 10990 7657 10998 7677
rect 10961 7647 10998 7657
rect 11057 7677 11144 7687
rect 11057 7657 11066 7677
rect 11086 7657 11144 7677
rect 11057 7648 11144 7657
rect 11057 7647 11094 7648
rect 9077 7562 9114 7563
rect 8500 7541 8536 7562
rect 8926 7541 8957 7562
rect 9713 7543 9750 7566
rect 10327 7556 10362 7634
rect 10774 7628 10811 7637
rect 10774 7610 10784 7628
rect 10802 7610 10811 7628
rect 10774 7600 10811 7610
rect 11113 7595 11144 7648
rect 11174 7677 11211 7748
rect 11382 7753 11775 7773
rect 11795 7753 11798 7773
rect 12126 7772 12157 7793
rect 12547 7772 12583 7793
rect 11969 7771 12006 7772
rect 11382 7748 11798 7753
rect 11968 7762 12006 7771
rect 11382 7747 11723 7748
rect 11326 7687 11357 7688
rect 11174 7657 11183 7677
rect 11203 7657 11211 7677
rect 11174 7647 11211 7657
rect 11270 7680 11357 7687
rect 11270 7677 11331 7680
rect 11270 7657 11279 7677
rect 11299 7660 11331 7677
rect 11352 7660 11357 7680
rect 11299 7657 11357 7660
rect 11270 7650 11357 7657
rect 11382 7677 11419 7747
rect 11685 7746 11722 7747
rect 11968 7742 11977 7762
rect 11997 7742 12006 7762
rect 11968 7734 12006 7742
rect 12072 7766 12157 7772
rect 12182 7771 12219 7772
rect 12072 7746 12080 7766
rect 12100 7746 12157 7766
rect 12072 7738 12157 7746
rect 12181 7762 12219 7771
rect 12181 7742 12190 7762
rect 12210 7742 12219 7762
rect 12072 7737 12108 7738
rect 12181 7734 12219 7742
rect 12285 7766 12370 7772
rect 12390 7771 12427 7772
rect 12285 7746 12293 7766
rect 12313 7765 12370 7766
rect 12313 7746 12342 7765
rect 12285 7745 12342 7746
rect 12363 7745 12370 7765
rect 12285 7738 12370 7745
rect 12389 7762 12427 7771
rect 12389 7742 12398 7762
rect 12418 7742 12427 7762
rect 12285 7737 12321 7738
rect 12389 7734 12427 7742
rect 12493 7766 12637 7772
rect 12493 7746 12501 7766
rect 12521 7746 12553 7766
rect 12577 7746 12609 7766
rect 12629 7746 12637 7766
rect 12493 7738 12637 7746
rect 12493 7737 12529 7738
rect 12601 7737 12637 7738
rect 12703 7771 12740 7772
rect 12703 7770 12741 7771
rect 12703 7762 12767 7770
rect 12703 7742 12712 7762
rect 12732 7748 12767 7762
rect 12787 7748 12790 7768
rect 12732 7743 12790 7748
rect 12732 7742 12767 7743
rect 11969 7705 12006 7734
rect 11970 7703 12006 7705
rect 12182 7703 12219 7734
rect 11534 7687 11570 7688
rect 11382 7657 11391 7677
rect 11411 7657 11419 7677
rect 11270 7648 11326 7650
rect 11270 7647 11307 7648
rect 11382 7647 11419 7657
rect 11478 7677 11626 7687
rect 11726 7684 11822 7686
rect 11478 7657 11487 7677
rect 11507 7657 11597 7677
rect 11617 7657 11626 7677
rect 11478 7648 11626 7657
rect 11684 7677 11822 7684
rect 11970 7681 12219 7703
rect 12390 7702 12427 7734
rect 12703 7730 12767 7742
rect 12807 7704 12834 7882
rect 12666 7702 12834 7704
rect 12390 7698 12834 7702
rect 11684 7657 11693 7677
rect 11713 7657 11822 7677
rect 12390 7679 12439 7698
rect 12459 7679 12834 7698
rect 12390 7676 12834 7679
rect 12666 7675 12834 7676
rect 13534 7689 13563 7691
rect 13534 7684 13566 7689
rect 13534 7666 13541 7684
rect 13561 7666 13566 7684
rect 13627 7688 13658 8082
rect 13679 8107 13847 8108
rect 13679 8104 14123 8107
rect 13679 8085 14054 8104
rect 14074 8085 14123 8104
rect 14691 8106 14800 8126
rect 14820 8106 14829 8126
rect 13679 8081 14123 8085
rect 13679 8079 13847 8081
rect 13679 7901 13706 8079
rect 13746 8041 13810 8053
rect 14086 8049 14123 8081
rect 14294 8080 14543 8102
rect 14691 8099 14829 8106
rect 14887 8126 15035 8135
rect 14887 8106 14896 8126
rect 14916 8106 15006 8126
rect 15026 8106 15035 8126
rect 14691 8097 14787 8099
rect 14887 8096 15035 8106
rect 15094 8126 15131 8136
rect 15206 8135 15243 8136
rect 15187 8133 15243 8135
rect 15094 8106 15102 8126
rect 15122 8106 15131 8126
rect 14943 8095 14979 8096
rect 14294 8049 14331 8080
rect 14507 8078 14543 8080
rect 14507 8049 14544 8078
rect 13746 8040 13781 8041
rect 13723 8035 13781 8040
rect 13723 8015 13726 8035
rect 13746 8021 13781 8035
rect 13801 8021 13810 8041
rect 13746 8013 13810 8021
rect 13772 8012 13810 8013
rect 13773 8011 13810 8012
rect 13876 8045 13912 8046
rect 13984 8045 14020 8046
rect 13876 8037 14020 8045
rect 13876 8017 13884 8037
rect 13904 8036 13992 8037
rect 13904 8017 13937 8036
rect 13876 8016 13937 8017
rect 13961 8017 13992 8036
rect 14012 8017 14020 8037
rect 13961 8016 14020 8017
rect 13876 8011 14020 8016
rect 14086 8041 14124 8049
rect 14192 8045 14228 8046
rect 14086 8021 14095 8041
rect 14115 8021 14124 8041
rect 14086 8012 14124 8021
rect 14143 8038 14228 8045
rect 14143 8018 14150 8038
rect 14171 8037 14228 8038
rect 14171 8018 14200 8037
rect 14143 8017 14200 8018
rect 14220 8017 14228 8037
rect 14086 8011 14123 8012
rect 14143 8011 14228 8017
rect 14294 8041 14332 8049
rect 14405 8045 14441 8046
rect 14294 8021 14303 8041
rect 14323 8021 14332 8041
rect 14294 8012 14332 8021
rect 14356 8037 14441 8045
rect 14356 8017 14413 8037
rect 14433 8017 14441 8037
rect 14294 8011 14331 8012
rect 14356 8011 14441 8017
rect 14507 8041 14545 8049
rect 14507 8021 14516 8041
rect 14536 8021 14545 8041
rect 14791 8036 14828 8037
rect 15094 8036 15131 8106
rect 15156 8126 15243 8133
rect 15156 8123 15214 8126
rect 15156 8103 15161 8123
rect 15182 8106 15214 8123
rect 15234 8106 15243 8126
rect 15182 8103 15243 8106
rect 15156 8096 15243 8103
rect 15302 8126 15339 8136
rect 15302 8106 15310 8126
rect 15330 8106 15339 8126
rect 15156 8095 15187 8096
rect 14790 8035 15131 8036
rect 14507 8012 14545 8021
rect 14715 8030 15131 8035
rect 14507 8011 14544 8012
rect 13930 7990 13966 8011
rect 14356 7990 14387 8011
rect 14715 8010 14718 8030
rect 14738 8010 15131 8030
rect 15302 8035 15339 8106
rect 15369 8135 15400 8188
rect 16052 8187 16062 8205
rect 16080 8191 16701 8205
rect 16080 8187 16090 8191
rect 16531 8190 16701 8191
rect 15702 8173 15739 8183
rect 15702 8155 15711 8173
rect 15729 8155 15739 8173
rect 15702 8146 15739 8155
rect 16052 8177 16090 8187
rect 15419 8135 15456 8136
rect 15369 8126 15456 8135
rect 15369 8106 15427 8126
rect 15447 8106 15456 8126
rect 15369 8096 15456 8106
rect 15515 8126 15552 8136
rect 15515 8106 15523 8126
rect 15543 8106 15552 8126
rect 15369 8095 15400 8096
rect 15515 8035 15552 8106
rect 15707 8081 15738 8146
rect 16052 8099 16087 8177
rect 16664 8167 16701 8190
rect 16048 8090 16087 8099
rect 15706 8071 15743 8081
rect 15706 8069 15716 8071
rect 15640 8067 15716 8069
rect 15302 8011 15552 8035
rect 15637 8053 15716 8067
rect 15734 8053 15743 8071
rect 16048 8072 16058 8090
rect 16076 8072 16087 8090
rect 16048 8066 16087 8072
rect 16243 8142 16493 8166
rect 16243 8071 16280 8142
rect 16395 8081 16426 8082
rect 16048 8062 16085 8066
rect 15637 8050 15743 8053
rect 15109 7991 15130 8010
rect 15637 7991 15663 8050
rect 15706 8044 15743 8050
rect 16243 8051 16252 8071
rect 16272 8051 16280 8071
rect 16243 8041 16280 8051
rect 16339 8071 16426 8081
rect 16339 8051 16348 8071
rect 16368 8051 16426 8071
rect 16339 8042 16426 8051
rect 16339 8041 16376 8042
rect 16051 7991 16088 8000
rect 13763 7986 13863 7990
rect 13763 7982 13825 7986
rect 13763 7956 13770 7982
rect 13796 7960 13825 7982
rect 13851 7960 13863 7986
rect 13796 7956 13863 7960
rect 13763 7953 13863 7956
rect 13931 7953 13966 7990
rect 14028 7987 14387 7990
rect 14028 7982 14250 7987
rect 14028 7958 14041 7982
rect 14065 7963 14250 7982
rect 14274 7963 14387 7987
rect 14065 7958 14387 7963
rect 14028 7954 14387 7958
rect 14454 7982 14603 7990
rect 14454 7962 14465 7982
rect 14485 7962 14603 7982
rect 15109 7973 15663 7991
rect 15709 7980 15746 7982
rect 15637 7972 15663 7973
rect 15706 7972 15746 7980
rect 14454 7955 14603 7962
rect 15706 7960 15718 7972
rect 15697 7955 15718 7960
rect 14454 7954 14495 7955
rect 15113 7954 15718 7955
rect 15736 7954 15746 7972
rect 13778 7901 13815 7902
rect 13874 7901 13911 7902
rect 13930 7901 13966 7953
rect 13985 7901 14022 7902
rect 13678 7892 13816 7901
rect 13678 7872 13787 7892
rect 13807 7872 13816 7892
rect 13678 7865 13816 7872
rect 13874 7892 14022 7901
rect 13874 7872 13883 7892
rect 13903 7872 13993 7892
rect 14013 7872 14022 7892
rect 13678 7863 13774 7865
rect 13874 7862 14022 7872
rect 14081 7892 14118 7902
rect 14193 7901 14230 7902
rect 14174 7899 14230 7901
rect 14081 7872 14089 7892
rect 14109 7872 14118 7892
rect 13930 7861 13966 7862
rect 13778 7802 13815 7803
rect 14081 7802 14118 7872
rect 14143 7892 14230 7899
rect 14143 7889 14201 7892
rect 14143 7869 14148 7889
rect 14169 7872 14201 7889
rect 14221 7872 14230 7892
rect 14169 7869 14230 7872
rect 14143 7862 14230 7869
rect 14289 7892 14326 7902
rect 14289 7872 14297 7892
rect 14317 7872 14326 7892
rect 14143 7861 14174 7862
rect 13777 7801 14118 7802
rect 13702 7796 14118 7801
rect 13702 7776 13705 7796
rect 13725 7776 14118 7796
rect 14289 7801 14326 7872
rect 14356 7901 14387 7954
rect 15113 7945 15746 7954
rect 16049 7973 16060 7991
rect 16078 7973 16088 7991
rect 16395 7989 16426 8042
rect 16456 8071 16493 8142
rect 16664 8147 17057 8167
rect 17077 8147 17080 8167
rect 16664 8142 17080 8147
rect 16664 8141 17005 8142
rect 16608 8081 16639 8082
rect 16456 8051 16465 8071
rect 16485 8051 16493 8071
rect 16456 8041 16493 8051
rect 16552 8074 16639 8081
rect 16552 8071 16613 8074
rect 16552 8051 16561 8071
rect 16581 8054 16613 8071
rect 16634 8054 16639 8074
rect 16581 8051 16639 8054
rect 16552 8044 16639 8051
rect 16664 8071 16701 8141
rect 16967 8140 17004 8141
rect 19973 8114 20000 8292
rect 20040 8254 20104 8266
rect 20380 8262 20417 8294
rect 20588 8293 20837 8315
rect 20588 8262 20625 8293
rect 20801 8291 20837 8293
rect 20980 8296 21018 8337
rect 20801 8262 20838 8291
rect 20040 8253 20075 8254
rect 20017 8248 20075 8253
rect 20017 8228 20020 8248
rect 20040 8234 20075 8248
rect 20095 8234 20104 8254
rect 20040 8226 20104 8234
rect 20066 8225 20104 8226
rect 20067 8224 20104 8225
rect 20170 8258 20206 8259
rect 20278 8258 20314 8259
rect 20170 8252 20314 8258
rect 20170 8250 20236 8252
rect 20170 8230 20178 8250
rect 20198 8231 20236 8250
rect 20258 8250 20314 8252
rect 20258 8231 20286 8250
rect 20198 8230 20286 8231
rect 20306 8230 20314 8250
rect 20170 8224 20314 8230
rect 20380 8254 20418 8262
rect 20486 8258 20522 8259
rect 20380 8234 20389 8254
rect 20409 8234 20418 8254
rect 20380 8225 20418 8234
rect 20437 8251 20522 8258
rect 20437 8231 20444 8251
rect 20465 8250 20522 8251
rect 20465 8231 20494 8250
rect 20437 8230 20494 8231
rect 20514 8230 20522 8250
rect 20380 8224 20417 8225
rect 20437 8224 20522 8230
rect 20588 8254 20626 8262
rect 20699 8258 20735 8259
rect 20588 8234 20597 8254
rect 20617 8234 20626 8254
rect 20588 8225 20626 8234
rect 20650 8250 20735 8258
rect 20650 8230 20707 8250
rect 20727 8230 20735 8250
rect 20588 8224 20625 8225
rect 20650 8224 20735 8230
rect 20801 8254 20839 8262
rect 20801 8234 20810 8254
rect 20830 8234 20839 8254
rect 20801 8225 20839 8234
rect 20980 8261 21016 8296
rect 20980 8251 21017 8261
rect 20980 8233 20990 8251
rect 21008 8233 21017 8251
rect 20801 8224 20838 8225
rect 20980 8224 21017 8233
rect 20224 8203 20260 8224
rect 20650 8203 20681 8224
rect 20057 8199 20157 8203
rect 20057 8195 20119 8199
rect 20057 8169 20064 8195
rect 20090 8173 20119 8195
rect 20145 8173 20157 8199
rect 20090 8169 20157 8173
rect 20057 8166 20157 8169
rect 20225 8166 20260 8203
rect 20322 8200 20681 8203
rect 20322 8195 20544 8200
rect 20322 8171 20335 8195
rect 20359 8176 20544 8195
rect 20568 8176 20681 8200
rect 20359 8171 20681 8176
rect 20322 8167 20681 8171
rect 20748 8195 20897 8203
rect 20748 8175 20759 8195
rect 20779 8175 20897 8195
rect 20748 8168 20897 8175
rect 20748 8167 20789 8168
rect 20072 8114 20109 8115
rect 20168 8114 20205 8115
rect 20224 8114 20260 8166
rect 20279 8114 20316 8115
rect 19972 8105 20110 8114
rect 18908 8087 18939 8090
rect 16816 8081 16852 8082
rect 16664 8051 16673 8071
rect 16693 8051 16701 8071
rect 16552 8042 16608 8044
rect 16552 8041 16589 8042
rect 16664 8041 16701 8051
rect 16760 8071 16908 8081
rect 17008 8078 17104 8080
rect 16760 8051 16769 8071
rect 16789 8051 16879 8071
rect 16899 8051 16908 8071
rect 16760 8042 16908 8051
rect 16966 8071 17104 8078
rect 16966 8051 16975 8071
rect 16995 8051 17104 8071
rect 16966 8042 17104 8051
rect 18908 8061 18915 8087
rect 18934 8061 18939 8087
rect 16760 8041 16797 8042
rect 16816 7990 16852 8042
rect 16871 8041 16908 8042
rect 16967 8041 17004 8042
rect 16287 7988 16328 7989
rect 15113 7938 15745 7945
rect 15113 7936 15175 7938
rect 14691 7926 14859 7927
rect 15113 7926 15135 7936
rect 14406 7901 14443 7902
rect 14356 7892 14443 7901
rect 14356 7872 14414 7892
rect 14434 7872 14443 7892
rect 14356 7862 14443 7872
rect 14502 7892 14539 7902
rect 14502 7872 14510 7892
rect 14530 7872 14539 7892
rect 14356 7861 14387 7862
rect 14502 7801 14539 7872
rect 14289 7777 14539 7801
rect 14691 7900 15135 7926
rect 14691 7898 14859 7900
rect 14691 7720 14718 7898
rect 14758 7860 14822 7872
rect 15098 7868 15135 7900
rect 15306 7899 15555 7921
rect 15306 7868 15343 7899
rect 15519 7897 15555 7899
rect 15519 7868 15556 7897
rect 14758 7859 14793 7860
rect 14735 7854 14793 7859
rect 14735 7834 14738 7854
rect 14758 7840 14793 7854
rect 14813 7840 14822 7860
rect 14758 7832 14822 7840
rect 14784 7831 14822 7832
rect 14785 7830 14822 7831
rect 14888 7864 14924 7865
rect 14996 7864 15032 7865
rect 14888 7856 15032 7864
rect 14888 7836 14896 7856
rect 14916 7836 14945 7856
rect 14888 7835 14945 7836
rect 14967 7836 15004 7856
rect 15024 7836 15032 7856
rect 14967 7835 15032 7836
rect 14888 7830 15032 7835
rect 15098 7860 15136 7868
rect 15204 7864 15240 7865
rect 15098 7840 15107 7860
rect 15127 7840 15136 7860
rect 15098 7831 15136 7840
rect 15155 7857 15240 7864
rect 15155 7837 15162 7857
rect 15183 7856 15240 7857
rect 15183 7837 15212 7856
rect 15155 7836 15212 7837
rect 15232 7836 15240 7856
rect 15098 7830 15135 7831
rect 15155 7830 15240 7836
rect 15306 7860 15344 7868
rect 15417 7864 15453 7865
rect 15306 7840 15315 7860
rect 15335 7840 15344 7860
rect 15306 7831 15344 7840
rect 15368 7856 15453 7864
rect 15368 7836 15425 7856
rect 15445 7836 15453 7856
rect 15306 7830 15343 7831
rect 15368 7830 15453 7836
rect 15519 7860 15557 7868
rect 15519 7840 15528 7860
rect 15548 7840 15557 7860
rect 15519 7831 15557 7840
rect 15519 7830 15556 7831
rect 14942 7809 14978 7830
rect 15368 7809 15399 7830
rect 14775 7805 14875 7809
rect 14775 7801 14837 7805
rect 14775 7775 14782 7801
rect 14808 7779 14837 7801
rect 14863 7779 14875 7805
rect 14808 7775 14875 7779
rect 14775 7772 14875 7775
rect 14943 7772 14978 7809
rect 15040 7806 15399 7809
rect 15040 7801 15262 7806
rect 15040 7777 15053 7801
rect 15077 7782 15262 7801
rect 15286 7782 15399 7806
rect 15077 7777 15399 7782
rect 15040 7773 15399 7777
rect 15466 7801 15615 7809
rect 15466 7781 15477 7801
rect 15497 7781 15615 7801
rect 15466 7774 15615 7781
rect 15706 7789 15745 7938
rect 16049 7824 16088 7973
rect 16179 7981 16328 7988
rect 16179 7961 16297 7981
rect 16317 7961 16328 7981
rect 16179 7953 16328 7961
rect 16395 7985 16754 7989
rect 16395 7980 16717 7985
rect 16395 7956 16508 7980
rect 16532 7961 16717 7980
rect 16741 7961 16754 7985
rect 16532 7956 16754 7961
rect 16395 7953 16754 7956
rect 16816 7953 16851 7990
rect 16919 7987 17019 7990
rect 16919 7983 16986 7987
rect 16919 7957 16931 7983
rect 16957 7961 16986 7983
rect 17012 7961 17019 7987
rect 16957 7957 17019 7961
rect 16919 7953 17019 7957
rect 16395 7932 16426 7953
rect 16816 7932 16852 7953
rect 16238 7931 16275 7932
rect 16237 7922 16275 7931
rect 16237 7902 16246 7922
rect 16266 7902 16275 7922
rect 16237 7894 16275 7902
rect 16341 7926 16426 7932
rect 16451 7931 16488 7932
rect 16341 7906 16349 7926
rect 16369 7906 16426 7926
rect 16341 7898 16426 7906
rect 16450 7922 16488 7931
rect 16450 7902 16459 7922
rect 16479 7902 16488 7922
rect 16341 7897 16377 7898
rect 16450 7894 16488 7902
rect 16554 7926 16639 7932
rect 16659 7931 16696 7932
rect 16554 7906 16562 7926
rect 16582 7925 16639 7926
rect 16582 7906 16611 7925
rect 16554 7905 16611 7906
rect 16632 7905 16639 7925
rect 16554 7898 16639 7905
rect 16658 7922 16696 7931
rect 16658 7902 16667 7922
rect 16687 7902 16696 7922
rect 16554 7897 16590 7898
rect 16658 7894 16696 7902
rect 16762 7927 16906 7932
rect 16762 7926 16827 7927
rect 16762 7906 16770 7926
rect 16790 7906 16827 7926
rect 16849 7926 16906 7927
rect 16849 7906 16878 7926
rect 16898 7906 16906 7926
rect 16762 7898 16906 7906
rect 16762 7897 16798 7898
rect 16870 7897 16906 7898
rect 16972 7931 17009 7932
rect 16972 7930 17010 7931
rect 16972 7922 17036 7930
rect 16972 7902 16981 7922
rect 17001 7908 17036 7922
rect 17056 7908 17059 7928
rect 17001 7903 17059 7908
rect 17001 7902 17036 7903
rect 16238 7865 16275 7894
rect 16239 7863 16275 7865
rect 16451 7863 16488 7894
rect 16239 7841 16488 7863
rect 16659 7862 16696 7894
rect 16972 7890 17036 7902
rect 17076 7864 17103 8042
rect 16935 7862 17103 7864
rect 16659 7836 17103 7862
rect 17255 7961 17505 7985
rect 17255 7890 17292 7961
rect 17407 7900 17438 7901
rect 17255 7870 17264 7890
rect 17284 7870 17292 7890
rect 17255 7860 17292 7870
rect 17351 7890 17438 7900
rect 17351 7870 17360 7890
rect 17380 7870 17438 7890
rect 17351 7861 17438 7870
rect 17351 7860 17388 7861
rect 16659 7826 16681 7836
rect 16935 7835 17103 7836
rect 16619 7824 16681 7826
rect 16049 7817 16681 7824
rect 15466 7773 15507 7774
rect 14790 7720 14827 7721
rect 14886 7720 14923 7721
rect 14942 7720 14978 7772
rect 14997 7720 15034 7721
rect 14690 7711 14828 7720
rect 14690 7691 14799 7711
rect 14819 7691 14828 7711
rect 13627 7687 13797 7688
rect 13627 7672 14073 7687
rect 14690 7684 14828 7691
rect 14886 7711 15034 7720
rect 14886 7691 14895 7711
rect 14915 7691 15005 7711
rect 15025 7691 15034 7711
rect 14690 7682 14786 7684
rect 13534 7661 13566 7666
rect 11684 7648 11822 7657
rect 11478 7647 11515 7648
rect 11534 7596 11570 7648
rect 11589 7647 11626 7648
rect 11685 7647 11722 7648
rect 11005 7594 11046 7595
rect 10897 7587 11046 7594
rect 10897 7567 11015 7587
rect 11035 7567 11046 7587
rect 10897 7559 11046 7567
rect 11113 7591 11472 7595
rect 11113 7586 11435 7591
rect 11113 7562 11226 7586
rect 11250 7567 11435 7586
rect 11459 7567 11472 7591
rect 11250 7562 11472 7567
rect 11113 7559 11472 7562
rect 11534 7559 11569 7596
rect 11637 7593 11737 7596
rect 11637 7589 11704 7593
rect 11637 7563 11649 7589
rect 11675 7567 11704 7589
rect 11730 7567 11737 7593
rect 11675 7563 11737 7567
rect 11637 7559 11737 7563
rect 10324 7546 10362 7556
rect 9713 7542 9883 7543
rect 10324 7542 10334 7546
rect 8333 7537 8433 7541
rect 8333 7533 8395 7537
rect 8333 7507 8340 7533
rect 8366 7511 8395 7533
rect 8421 7511 8433 7537
rect 8366 7507 8433 7511
rect 8333 7504 8433 7507
rect 8501 7504 8536 7541
rect 8598 7538 8957 7541
rect 8598 7533 8820 7538
rect 8598 7509 8611 7533
rect 8635 7514 8820 7533
rect 8844 7514 8957 7538
rect 8635 7509 8957 7514
rect 8598 7505 8957 7509
rect 9024 7533 9173 7541
rect 9024 7513 9035 7533
rect 9055 7513 9173 7533
rect 9713 7528 10334 7542
rect 10352 7528 10362 7546
rect 11113 7538 11144 7559
rect 11534 7538 11570 7559
rect 9713 7522 10362 7528
rect 10777 7529 10814 7538
rect 10956 7537 10993 7538
rect 9713 7521 10361 7522
rect 10324 7519 10361 7521
rect 9024 7506 9173 7513
rect 10777 7511 10786 7529
rect 10804 7511 10814 7529
rect 9024 7505 9065 7506
rect 8348 7452 8385 7453
rect 8444 7452 8481 7453
rect 8500 7452 8536 7504
rect 8555 7452 8592 7453
rect 8248 7443 8386 7452
rect 8248 7423 8357 7443
rect 8377 7423 8386 7443
rect 8248 7416 8386 7423
rect 8444 7443 8592 7452
rect 8444 7423 8453 7443
rect 8473 7423 8563 7443
rect 8583 7423 8592 7443
rect 8248 7414 8344 7416
rect 8444 7413 8592 7423
rect 8651 7443 8688 7453
rect 8763 7452 8800 7453
rect 8744 7450 8800 7452
rect 8651 7423 8659 7443
rect 8679 7423 8688 7443
rect 8500 7412 8536 7413
rect 8348 7353 8385 7354
rect 8651 7353 8688 7423
rect 8713 7443 8800 7450
rect 8713 7440 8771 7443
rect 8713 7420 8718 7440
rect 8739 7423 8771 7440
rect 8791 7423 8800 7443
rect 8739 7420 8800 7423
rect 8713 7413 8800 7420
rect 8859 7443 8896 7453
rect 8859 7423 8867 7443
rect 8887 7423 8896 7443
rect 8713 7412 8744 7413
rect 8347 7352 8688 7353
rect 8272 7347 8688 7352
rect 8272 7327 8275 7347
rect 8295 7327 8688 7347
rect 8859 7352 8896 7423
rect 8926 7452 8957 7505
rect 10777 7501 10814 7511
rect 10778 7466 10814 7501
rect 10955 7528 10993 7537
rect 10955 7508 10964 7528
rect 10984 7508 10993 7528
rect 10955 7500 10993 7508
rect 11059 7532 11144 7538
rect 11169 7537 11206 7538
rect 11059 7512 11067 7532
rect 11087 7512 11144 7532
rect 11059 7504 11144 7512
rect 11168 7528 11206 7537
rect 11168 7508 11177 7528
rect 11197 7508 11206 7528
rect 11059 7503 11095 7504
rect 11168 7500 11206 7508
rect 11272 7532 11357 7538
rect 11377 7537 11414 7538
rect 11272 7512 11280 7532
rect 11300 7531 11357 7532
rect 11300 7512 11329 7531
rect 11272 7511 11329 7512
rect 11350 7511 11357 7531
rect 11272 7504 11357 7511
rect 11376 7528 11414 7537
rect 11376 7508 11385 7528
rect 11405 7508 11414 7528
rect 11272 7503 11308 7504
rect 11376 7500 11414 7508
rect 11480 7532 11624 7538
rect 11480 7512 11488 7532
rect 11508 7531 11596 7532
rect 11508 7512 11536 7531
rect 11480 7510 11536 7512
rect 11558 7512 11596 7531
rect 11616 7512 11624 7532
rect 11558 7510 11624 7512
rect 11480 7504 11624 7510
rect 11480 7503 11516 7504
rect 11588 7503 11624 7504
rect 11690 7537 11727 7538
rect 11690 7536 11728 7537
rect 11690 7528 11754 7536
rect 11690 7508 11699 7528
rect 11719 7514 11754 7528
rect 11774 7514 11777 7534
rect 11719 7509 11777 7514
rect 11719 7508 11754 7509
rect 10956 7471 10993 7500
rect 8976 7452 9013 7453
rect 8926 7443 9013 7452
rect 8926 7423 8984 7443
rect 9004 7423 9013 7443
rect 8926 7413 9013 7423
rect 9072 7443 9109 7453
rect 9072 7423 9080 7443
rect 9100 7423 9109 7443
rect 8926 7412 8957 7413
rect 9072 7352 9109 7423
rect 10327 7447 10364 7457
rect 10327 7429 10336 7447
rect 10354 7429 10364 7447
rect 10327 7420 10364 7429
rect 10776 7425 10814 7466
rect 10957 7469 10993 7471
rect 11169 7469 11206 7500
rect 10957 7447 11206 7469
rect 11377 7468 11414 7500
rect 11690 7496 11754 7508
rect 11794 7470 11821 7648
rect 11653 7468 11821 7470
rect 11377 7442 11821 7468
rect 11378 7425 11402 7442
rect 11653 7441 11821 7442
rect 10327 7396 10362 7420
rect 10325 7372 10362 7396
rect 10324 7366 10362 7372
rect 8859 7328 9109 7352
rect 9735 7348 10362 7366
rect 10776 7407 11403 7425
rect 12029 7421 12279 7445
rect 10776 7401 10814 7407
rect 10776 7377 10813 7401
rect 10776 7353 10811 7377
rect 9317 7331 9485 7332
rect 9736 7331 9760 7348
rect 9317 7305 9761 7331
rect 9317 7303 9485 7305
rect 9317 7125 9344 7303
rect 9384 7265 9448 7277
rect 9724 7273 9761 7305
rect 9932 7304 10181 7326
rect 9932 7273 9969 7304
rect 10145 7302 10181 7304
rect 10324 7307 10362 7348
rect 10774 7344 10811 7353
rect 10774 7326 10784 7344
rect 10802 7326 10811 7344
rect 10774 7316 10811 7326
rect 12029 7350 12066 7421
rect 12181 7360 12212 7361
rect 12029 7330 12038 7350
rect 12058 7330 12066 7350
rect 12029 7320 12066 7330
rect 12125 7350 12212 7360
rect 12125 7330 12134 7350
rect 12154 7330 12212 7350
rect 12125 7321 12212 7330
rect 12125 7320 12162 7321
rect 10145 7273 10182 7302
rect 9384 7264 9419 7265
rect 9361 7259 9419 7264
rect 9361 7239 9364 7259
rect 9384 7245 9419 7259
rect 9439 7245 9448 7265
rect 9384 7237 9448 7245
rect 9410 7236 9448 7237
rect 9411 7235 9448 7236
rect 9514 7269 9550 7270
rect 9622 7269 9658 7270
rect 9514 7263 9658 7269
rect 9514 7261 9580 7263
rect 9514 7241 9522 7261
rect 9542 7242 9580 7261
rect 9602 7261 9658 7263
rect 9602 7242 9630 7261
rect 9542 7241 9630 7242
rect 9650 7241 9658 7261
rect 9514 7235 9658 7241
rect 9724 7265 9762 7273
rect 9830 7269 9866 7270
rect 9724 7245 9733 7265
rect 9753 7245 9762 7265
rect 9724 7236 9762 7245
rect 9781 7262 9866 7269
rect 9781 7242 9788 7262
rect 9809 7261 9866 7262
rect 9809 7242 9838 7261
rect 9781 7241 9838 7242
rect 9858 7241 9866 7261
rect 9724 7235 9761 7236
rect 9781 7235 9866 7241
rect 9932 7265 9970 7273
rect 10043 7269 10079 7270
rect 9932 7245 9941 7265
rect 9961 7245 9970 7265
rect 9932 7236 9970 7245
rect 9994 7261 10079 7269
rect 9994 7241 10051 7261
rect 10071 7241 10079 7261
rect 9932 7235 9969 7236
rect 9994 7235 10079 7241
rect 10145 7265 10183 7273
rect 10145 7245 10154 7265
rect 10174 7245 10183 7265
rect 10145 7236 10183 7245
rect 10324 7272 10360 7307
rect 10324 7262 10361 7272
rect 12181 7268 12212 7321
rect 12242 7350 12279 7421
rect 12450 7426 12843 7446
rect 12863 7426 12866 7446
rect 12450 7421 12866 7426
rect 12450 7420 12791 7421
rect 12394 7360 12425 7361
rect 12242 7330 12251 7350
rect 12271 7330 12279 7350
rect 12242 7320 12279 7330
rect 12338 7353 12425 7360
rect 12338 7350 12399 7353
rect 12338 7330 12347 7350
rect 12367 7333 12399 7350
rect 12420 7333 12425 7353
rect 12367 7330 12425 7333
rect 12338 7323 12425 7330
rect 12450 7350 12487 7420
rect 12753 7419 12790 7420
rect 12602 7360 12638 7361
rect 12450 7330 12459 7350
rect 12479 7330 12487 7350
rect 12338 7321 12394 7323
rect 12338 7320 12375 7321
rect 12450 7320 12487 7330
rect 12546 7350 12694 7360
rect 12794 7357 12890 7359
rect 12546 7330 12555 7350
rect 12575 7330 12665 7350
rect 12685 7330 12694 7350
rect 12546 7321 12694 7330
rect 12752 7350 12890 7357
rect 12752 7330 12761 7350
rect 12781 7330 12890 7350
rect 12752 7321 12890 7330
rect 12546 7320 12583 7321
rect 12602 7269 12638 7321
rect 12657 7320 12694 7321
rect 12753 7320 12790 7321
rect 12073 7267 12114 7268
rect 10324 7244 10334 7262
rect 10352 7244 10361 7262
rect 11965 7260 12114 7267
rect 10777 7252 10814 7254
rect 10777 7251 11425 7252
rect 10145 7235 10182 7236
rect 10324 7235 10361 7244
rect 10776 7245 11425 7251
rect 9568 7214 9604 7235
rect 9994 7214 10025 7235
rect 10776 7227 10786 7245
rect 10804 7231 11425 7245
rect 11965 7240 12083 7260
rect 12103 7240 12114 7260
rect 11965 7232 12114 7240
rect 12181 7264 12540 7268
rect 12181 7259 12503 7264
rect 12181 7235 12294 7259
rect 12318 7240 12503 7259
rect 12527 7240 12540 7264
rect 12318 7235 12540 7240
rect 12181 7232 12540 7235
rect 12602 7232 12637 7269
rect 12705 7266 12805 7269
rect 12705 7262 12772 7266
rect 12705 7236 12717 7262
rect 12743 7240 12772 7262
rect 12798 7240 12805 7266
rect 12743 7236 12805 7240
rect 12705 7232 12805 7236
rect 10804 7227 10814 7231
rect 11255 7230 11425 7231
rect 10776 7217 10814 7227
rect 9401 7210 9501 7214
rect 9401 7206 9463 7210
rect 9401 7180 9408 7206
rect 9434 7184 9463 7206
rect 9489 7184 9501 7210
rect 9434 7180 9501 7184
rect 9401 7177 9501 7180
rect 9569 7177 9604 7214
rect 9666 7211 10025 7214
rect 9666 7206 9888 7211
rect 9666 7182 9679 7206
rect 9703 7187 9888 7206
rect 9912 7187 10025 7211
rect 9703 7182 10025 7187
rect 9666 7178 10025 7182
rect 10092 7206 10241 7214
rect 10092 7186 10103 7206
rect 10123 7186 10241 7206
rect 10092 7179 10241 7186
rect 10092 7178 10133 7179
rect 9416 7125 9453 7126
rect 9512 7125 9549 7126
rect 9568 7125 9604 7177
rect 9623 7125 9660 7126
rect 9316 7116 9454 7125
rect 8304 7097 8472 7098
rect 8304 7094 8748 7097
rect 8304 7075 8679 7094
rect 8699 7075 8748 7094
rect 9316 7096 9425 7116
rect 9445 7096 9454 7116
rect 8304 7071 8748 7075
rect 8304 7069 8472 7071
rect 8304 6891 8331 7069
rect 8371 7031 8435 7043
rect 8711 7039 8748 7071
rect 8919 7070 9168 7092
rect 9316 7089 9454 7096
rect 9512 7116 9660 7125
rect 9512 7096 9521 7116
rect 9541 7096 9631 7116
rect 9651 7096 9660 7116
rect 9316 7087 9412 7089
rect 9512 7086 9660 7096
rect 9719 7116 9756 7126
rect 9831 7125 9868 7126
rect 9812 7123 9868 7125
rect 9719 7096 9727 7116
rect 9747 7096 9756 7116
rect 9568 7085 9604 7086
rect 8919 7039 8956 7070
rect 9132 7068 9168 7070
rect 9132 7039 9169 7068
rect 8371 7030 8406 7031
rect 8348 7025 8406 7030
rect 8348 7005 8351 7025
rect 8371 7011 8406 7025
rect 8426 7011 8435 7031
rect 8371 7003 8435 7011
rect 8397 7002 8435 7003
rect 8398 7001 8435 7002
rect 8501 7035 8537 7036
rect 8609 7035 8645 7036
rect 8501 7027 8645 7035
rect 8501 7007 8509 7027
rect 8529 7007 8561 7027
rect 8585 7007 8617 7027
rect 8637 7007 8645 7027
rect 8501 7001 8645 7007
rect 8711 7031 8749 7039
rect 8817 7035 8853 7036
rect 8711 7011 8720 7031
rect 8740 7011 8749 7031
rect 8711 7002 8749 7011
rect 8768 7028 8853 7035
rect 8768 7008 8775 7028
rect 8796 7027 8853 7028
rect 8796 7008 8825 7027
rect 8768 7007 8825 7008
rect 8845 7007 8853 7027
rect 8711 7001 8748 7002
rect 8768 7001 8853 7007
rect 8919 7031 8957 7039
rect 9030 7035 9066 7036
rect 8919 7011 8928 7031
rect 8948 7011 8957 7031
rect 8919 7002 8957 7011
rect 8981 7027 9066 7035
rect 8981 7007 9038 7027
rect 9058 7007 9066 7027
rect 8919 7001 8956 7002
rect 8981 7001 9066 7007
rect 9132 7031 9170 7039
rect 9132 7011 9141 7031
rect 9161 7011 9170 7031
rect 9416 7026 9453 7027
rect 9719 7026 9756 7096
rect 9781 7116 9868 7123
rect 9781 7113 9839 7116
rect 9781 7093 9786 7113
rect 9807 7096 9839 7113
rect 9859 7096 9868 7116
rect 9807 7093 9868 7096
rect 9781 7086 9868 7093
rect 9927 7116 9964 7126
rect 9927 7096 9935 7116
rect 9955 7096 9964 7116
rect 9781 7085 9812 7086
rect 9415 7025 9756 7026
rect 9132 7002 9170 7011
rect 9340 7020 9756 7025
rect 9132 7001 9169 7002
rect 8555 6980 8591 7001
rect 8981 6980 9012 7001
rect 9340 7000 9343 7020
rect 9363 7000 9756 7020
rect 9927 7025 9964 7096
rect 9994 7125 10025 7178
rect 10327 7163 10364 7173
rect 10327 7145 10336 7163
rect 10354 7145 10364 7163
rect 10327 7136 10364 7145
rect 10776 7139 10811 7217
rect 11388 7207 11425 7230
rect 12181 7211 12212 7232
rect 12602 7211 12638 7232
rect 12024 7210 12061 7211
rect 10044 7125 10081 7126
rect 9994 7116 10081 7125
rect 9994 7096 10052 7116
rect 10072 7096 10081 7116
rect 9994 7086 10081 7096
rect 10140 7116 10177 7126
rect 10140 7096 10148 7116
rect 10168 7096 10177 7116
rect 9994 7085 10025 7086
rect 10140 7025 10177 7096
rect 10332 7071 10363 7136
rect 10772 7130 10811 7139
rect 10772 7112 10782 7130
rect 10800 7112 10811 7130
rect 10772 7106 10811 7112
rect 10967 7182 11217 7206
rect 10967 7111 11004 7182
rect 11119 7121 11150 7122
rect 10772 7102 10809 7106
rect 10967 7091 10976 7111
rect 10996 7091 11004 7111
rect 10967 7081 11004 7091
rect 11063 7111 11150 7121
rect 11063 7091 11072 7111
rect 11092 7091 11150 7111
rect 11063 7082 11150 7091
rect 11063 7081 11100 7082
rect 10331 7061 10368 7071
rect 10331 7059 10341 7061
rect 10265 7057 10341 7059
rect 9927 7001 10177 7025
rect 10262 7043 10341 7057
rect 10359 7043 10368 7061
rect 10262 7040 10368 7043
rect 9734 6981 9755 7000
rect 10262 6981 10288 7040
rect 10331 7034 10368 7040
rect 10775 7031 10812 7040
rect 8388 6976 8488 6980
rect 8388 6972 8450 6976
rect 8388 6946 8395 6972
rect 8421 6950 8450 6972
rect 8476 6950 8488 6976
rect 8421 6946 8488 6950
rect 8388 6943 8488 6946
rect 8556 6943 8591 6980
rect 8653 6977 9012 6980
rect 8653 6972 8875 6977
rect 8653 6948 8666 6972
rect 8690 6953 8875 6972
rect 8899 6953 9012 6977
rect 8690 6948 9012 6953
rect 8653 6944 9012 6948
rect 9079 6972 9228 6980
rect 9079 6952 9090 6972
rect 9110 6952 9228 6972
rect 9734 6963 10288 6981
rect 10773 7013 10784 7031
rect 10802 7013 10812 7031
rect 11119 7029 11150 7082
rect 11180 7111 11217 7182
rect 11388 7187 11781 7207
rect 11801 7187 11804 7207
rect 11388 7182 11804 7187
rect 12023 7201 12061 7210
rect 11388 7181 11729 7182
rect 12023 7181 12032 7201
rect 12052 7181 12061 7201
rect 11332 7121 11363 7122
rect 11180 7091 11189 7111
rect 11209 7091 11217 7111
rect 11180 7081 11217 7091
rect 11276 7114 11363 7121
rect 11276 7111 11337 7114
rect 11276 7091 11285 7111
rect 11305 7094 11337 7111
rect 11358 7094 11363 7114
rect 11305 7091 11363 7094
rect 11276 7084 11363 7091
rect 11388 7111 11425 7181
rect 11691 7180 11728 7181
rect 12023 7173 12061 7181
rect 12127 7205 12212 7211
rect 12237 7210 12274 7211
rect 12127 7185 12135 7205
rect 12155 7185 12212 7205
rect 12127 7177 12212 7185
rect 12236 7201 12274 7210
rect 12236 7181 12245 7201
rect 12265 7181 12274 7201
rect 12127 7176 12163 7177
rect 12236 7173 12274 7181
rect 12340 7205 12425 7211
rect 12445 7210 12482 7211
rect 12340 7185 12348 7205
rect 12368 7204 12425 7205
rect 12368 7185 12397 7204
rect 12340 7184 12397 7185
rect 12418 7184 12425 7204
rect 12340 7177 12425 7184
rect 12444 7201 12482 7210
rect 12444 7181 12453 7201
rect 12473 7181 12482 7201
rect 12340 7176 12376 7177
rect 12444 7173 12482 7181
rect 12548 7205 12692 7211
rect 12548 7185 12556 7205
rect 12576 7203 12664 7205
rect 12576 7186 12612 7203
rect 12636 7186 12664 7203
rect 12576 7185 12664 7186
rect 12684 7185 12692 7205
rect 12548 7177 12692 7185
rect 12548 7176 12584 7177
rect 12656 7176 12692 7177
rect 12758 7210 12795 7211
rect 12758 7209 12796 7210
rect 12758 7201 12822 7209
rect 12758 7181 12767 7201
rect 12787 7187 12822 7201
rect 12842 7187 12845 7207
rect 12787 7182 12845 7187
rect 12787 7181 12822 7182
rect 12024 7144 12061 7173
rect 12025 7142 12061 7144
rect 12237 7142 12274 7173
rect 11540 7121 11576 7122
rect 11388 7091 11397 7111
rect 11417 7091 11425 7111
rect 11276 7082 11332 7084
rect 11276 7081 11313 7082
rect 11388 7081 11425 7091
rect 11484 7111 11632 7121
rect 12025 7120 12274 7142
rect 12445 7141 12482 7173
rect 12758 7169 12822 7181
rect 12862 7143 12889 7321
rect 12721 7141 12889 7143
rect 12445 7130 12889 7141
rect 11732 7118 11828 7120
rect 11484 7091 11493 7111
rect 11513 7091 11603 7111
rect 11623 7091 11632 7111
rect 11484 7082 11632 7091
rect 11690 7111 11828 7118
rect 12445 7115 12891 7130
rect 12721 7114 12891 7115
rect 11690 7091 11699 7111
rect 11719 7091 11828 7111
rect 11690 7082 11828 7091
rect 11484 7081 11521 7082
rect 11540 7030 11576 7082
rect 11595 7081 11632 7082
rect 11691 7081 11728 7082
rect 11011 7028 11052 7029
rect 10334 6970 10371 6972
rect 10262 6962 10288 6963
rect 10331 6962 10371 6970
rect 9079 6945 9228 6952
rect 10331 6950 10343 6962
rect 10322 6945 10343 6950
rect 9079 6944 9120 6945
rect 9738 6944 10343 6945
rect 10361 6944 10371 6962
rect 8403 6891 8440 6892
rect 8499 6891 8536 6892
rect 8555 6891 8591 6943
rect 8610 6891 8647 6892
rect 8303 6882 8441 6891
rect 8303 6862 8412 6882
rect 8432 6862 8441 6882
rect 8303 6855 8441 6862
rect 8499 6882 8647 6891
rect 8499 6862 8508 6882
rect 8528 6862 8618 6882
rect 8638 6862 8647 6882
rect 8303 6853 8399 6855
rect 8499 6852 8647 6862
rect 8706 6882 8743 6892
rect 8818 6891 8855 6892
rect 8799 6889 8855 6891
rect 8706 6862 8714 6882
rect 8734 6862 8743 6882
rect 8555 6851 8591 6852
rect 8403 6792 8440 6793
rect 8706 6792 8743 6862
rect 8768 6882 8855 6889
rect 8768 6879 8826 6882
rect 8768 6859 8773 6879
rect 8794 6862 8826 6879
rect 8846 6862 8855 6882
rect 8794 6859 8855 6862
rect 8768 6852 8855 6859
rect 8914 6882 8951 6892
rect 8914 6862 8922 6882
rect 8942 6862 8951 6882
rect 8768 6851 8799 6852
rect 8402 6791 8743 6792
rect 8327 6786 8743 6791
rect 8327 6766 8330 6786
rect 8350 6766 8743 6786
rect 8914 6791 8951 6862
rect 8981 6891 9012 6944
rect 9738 6935 10371 6944
rect 9738 6928 10370 6935
rect 9738 6926 9800 6928
rect 9316 6916 9484 6917
rect 9738 6916 9760 6926
rect 9031 6891 9068 6892
rect 8981 6882 9068 6891
rect 8981 6862 9039 6882
rect 9059 6862 9068 6882
rect 8981 6852 9068 6862
rect 9127 6882 9164 6892
rect 9127 6862 9135 6882
rect 9155 6862 9164 6882
rect 8981 6851 9012 6852
rect 9127 6791 9164 6862
rect 8914 6767 9164 6791
rect 9316 6890 9760 6916
rect 9316 6888 9484 6890
rect 9316 6710 9343 6888
rect 9383 6850 9447 6862
rect 9723 6858 9760 6890
rect 9931 6889 10180 6911
rect 9931 6858 9968 6889
rect 10144 6887 10180 6889
rect 10144 6858 10181 6887
rect 9383 6849 9418 6850
rect 9360 6844 9418 6849
rect 9360 6824 9363 6844
rect 9383 6830 9418 6844
rect 9438 6830 9447 6850
rect 9383 6822 9447 6830
rect 9409 6821 9447 6822
rect 9410 6820 9447 6821
rect 9513 6854 9549 6855
rect 9621 6854 9657 6855
rect 9513 6846 9657 6854
rect 9513 6826 9521 6846
rect 9541 6826 9570 6846
rect 9513 6825 9570 6826
rect 9592 6826 9629 6846
rect 9649 6826 9657 6846
rect 9592 6825 9657 6826
rect 9513 6820 9657 6825
rect 9723 6850 9761 6858
rect 9829 6854 9865 6855
rect 9723 6830 9732 6850
rect 9752 6830 9761 6850
rect 9723 6821 9761 6830
rect 9780 6847 9865 6854
rect 9780 6827 9787 6847
rect 9808 6846 9865 6847
rect 9808 6827 9837 6846
rect 9780 6826 9837 6827
rect 9857 6826 9865 6846
rect 9723 6820 9760 6821
rect 9780 6820 9865 6826
rect 9931 6850 9969 6858
rect 10042 6854 10078 6855
rect 9931 6830 9940 6850
rect 9960 6830 9969 6850
rect 9931 6821 9969 6830
rect 9993 6846 10078 6854
rect 9993 6826 10050 6846
rect 10070 6826 10078 6846
rect 9931 6820 9968 6821
rect 9993 6820 10078 6826
rect 10144 6850 10182 6858
rect 10144 6830 10153 6850
rect 10173 6830 10182 6850
rect 10144 6821 10182 6830
rect 10144 6820 10181 6821
rect 9567 6799 9603 6820
rect 9993 6799 10024 6820
rect 9400 6795 9500 6799
rect 9400 6791 9462 6795
rect 9400 6765 9407 6791
rect 9433 6769 9462 6791
rect 9488 6769 9500 6795
rect 9433 6765 9500 6769
rect 9400 6762 9500 6765
rect 9568 6762 9603 6799
rect 9665 6796 10024 6799
rect 9665 6791 9887 6796
rect 9665 6767 9678 6791
rect 9702 6772 9887 6791
rect 9911 6772 10024 6796
rect 9702 6767 10024 6772
rect 9665 6763 10024 6767
rect 10091 6791 10240 6799
rect 10091 6771 10102 6791
rect 10122 6771 10240 6791
rect 10091 6764 10240 6771
rect 10331 6779 10370 6928
rect 10773 6864 10812 7013
rect 10903 7021 11052 7028
rect 10903 7001 11021 7021
rect 11041 7001 11052 7021
rect 10903 6993 11052 7001
rect 11119 7025 11478 7029
rect 11119 7020 11441 7025
rect 11119 6996 11232 7020
rect 11256 7001 11441 7020
rect 11465 7001 11478 7025
rect 11256 6996 11478 7001
rect 11119 6993 11478 6996
rect 11540 6993 11575 7030
rect 11643 7027 11743 7030
rect 11643 7023 11710 7027
rect 11643 6997 11655 7023
rect 11681 7001 11710 7023
rect 11736 7001 11743 7027
rect 11681 6997 11743 7001
rect 11643 6993 11743 6997
rect 11119 6972 11150 6993
rect 11540 6972 11576 6993
rect 10962 6971 10999 6972
rect 10961 6962 10999 6971
rect 10961 6942 10970 6962
rect 10990 6942 10999 6962
rect 10961 6934 10999 6942
rect 11065 6966 11150 6972
rect 11175 6971 11212 6972
rect 11065 6946 11073 6966
rect 11093 6946 11150 6966
rect 11065 6938 11150 6946
rect 11174 6962 11212 6971
rect 11174 6942 11183 6962
rect 11203 6942 11212 6962
rect 11065 6937 11101 6938
rect 11174 6934 11212 6942
rect 11278 6966 11363 6972
rect 11383 6971 11420 6972
rect 11278 6946 11286 6966
rect 11306 6965 11363 6966
rect 11306 6946 11335 6965
rect 11278 6945 11335 6946
rect 11356 6945 11363 6965
rect 11278 6938 11363 6945
rect 11382 6962 11420 6971
rect 11382 6942 11391 6962
rect 11411 6942 11420 6962
rect 11278 6937 11314 6938
rect 11382 6934 11420 6942
rect 11486 6967 11630 6972
rect 11486 6966 11551 6967
rect 11486 6946 11494 6966
rect 11514 6946 11551 6966
rect 11573 6966 11630 6967
rect 11573 6946 11602 6966
rect 11622 6946 11630 6966
rect 11486 6938 11630 6946
rect 11486 6937 11522 6938
rect 11594 6937 11630 6938
rect 11696 6971 11733 6972
rect 11696 6970 11734 6971
rect 11696 6962 11760 6970
rect 11696 6942 11705 6962
rect 11725 6948 11760 6962
rect 11780 6948 11783 6968
rect 11725 6943 11783 6948
rect 11725 6942 11760 6943
rect 10962 6905 10999 6934
rect 10963 6903 10999 6905
rect 11175 6903 11212 6934
rect 10963 6881 11212 6903
rect 11383 6902 11420 6934
rect 11696 6930 11760 6942
rect 11800 6904 11827 7082
rect 11659 6902 11827 6904
rect 11383 6876 11827 6902
rect 11979 7001 12229 7025
rect 11979 6930 12016 7001
rect 12131 6940 12162 6941
rect 11979 6910 11988 6930
rect 12008 6910 12016 6930
rect 11979 6900 12016 6910
rect 12075 6930 12162 6940
rect 12075 6910 12084 6930
rect 12104 6910 12162 6930
rect 12075 6901 12162 6910
rect 12075 6900 12112 6901
rect 11383 6866 11405 6876
rect 11659 6875 11827 6876
rect 11343 6864 11405 6866
rect 10773 6857 11405 6864
rect 10772 6848 11405 6857
rect 12131 6848 12162 6901
rect 12192 6930 12229 7001
rect 12400 7006 12793 7026
rect 12813 7006 12816 7026
rect 12400 7001 12816 7006
rect 12400 7000 12741 7001
rect 12344 6940 12375 6941
rect 12192 6910 12201 6930
rect 12221 6910 12229 6930
rect 12192 6900 12229 6910
rect 12288 6933 12375 6940
rect 12288 6930 12349 6933
rect 12288 6910 12297 6930
rect 12317 6913 12349 6930
rect 12370 6913 12375 6933
rect 12317 6910 12375 6913
rect 12288 6903 12375 6910
rect 12400 6930 12437 7000
rect 12703 6999 12740 7000
rect 12552 6940 12588 6941
rect 12400 6910 12409 6930
rect 12429 6910 12437 6930
rect 12288 6901 12344 6903
rect 12288 6900 12325 6901
rect 12400 6900 12437 6910
rect 12496 6930 12644 6940
rect 12744 6937 12840 6939
rect 12496 6910 12505 6930
rect 12525 6910 12615 6930
rect 12635 6910 12644 6930
rect 12496 6901 12644 6910
rect 12702 6930 12840 6937
rect 12702 6910 12711 6930
rect 12731 6910 12840 6930
rect 12702 6901 12840 6910
rect 12496 6900 12533 6901
rect 12552 6849 12588 6901
rect 12607 6900 12644 6901
rect 12703 6900 12740 6901
rect 10772 6830 10782 6848
rect 10800 6847 11405 6848
rect 12023 6847 12064 6848
rect 10800 6842 10821 6847
rect 10800 6830 10812 6842
rect 11915 6840 12064 6847
rect 10772 6822 10812 6830
rect 10855 6829 10881 6830
rect 10772 6820 10809 6822
rect 10091 6763 10132 6764
rect 9415 6710 9452 6711
rect 9511 6710 9548 6711
rect 9567 6710 9603 6762
rect 9622 6710 9659 6711
rect 9315 6701 9453 6710
rect 9315 6681 9424 6701
rect 9444 6681 9453 6701
rect 9315 6674 9453 6681
rect 9511 6701 9659 6710
rect 9511 6681 9520 6701
rect 9540 6681 9630 6701
rect 9650 6681 9659 6701
rect 9315 6672 9411 6674
rect 9511 6671 9659 6681
rect 9718 6701 9755 6711
rect 9830 6710 9867 6711
rect 9811 6708 9867 6710
rect 9718 6681 9726 6701
rect 9746 6681 9755 6701
rect 9567 6670 9603 6671
rect 8030 6608 8038 6627
rect 8061 6608 8067 6627
rect 8030 6597 8067 6608
rect 8096 6630 8264 6631
rect 8096 6604 8540 6630
rect 8096 6602 8264 6604
rect 8033 6537 8066 6597
rect 6278 6458 6446 6460
rect 6002 6432 6446 6458
rect 6003 6415 6027 6432
rect 6278 6431 6446 6432
rect 6814 6460 7064 6484
rect 5050 6408 5088 6414
rect 4461 6390 5088 6408
rect 5401 6397 6028 6415
rect 5401 6391 5439 6397
rect 3425 6321 3675 6345
rect 4043 6373 4211 6374
rect 4462 6373 4486 6390
rect 4043 6347 4487 6373
rect 4043 6345 4211 6347
rect 4043 6167 4070 6345
rect 4110 6307 4174 6319
rect 4450 6315 4487 6347
rect 4658 6346 4907 6368
rect 4658 6315 4695 6346
rect 4871 6344 4907 6346
rect 5050 6349 5088 6390
rect 4871 6315 4908 6344
rect 4110 6306 4145 6307
rect 4087 6301 4145 6306
rect 4087 6281 4090 6301
rect 4110 6287 4145 6301
rect 4165 6287 4174 6307
rect 4110 6279 4174 6287
rect 4136 6278 4174 6279
rect 4137 6277 4174 6278
rect 4240 6311 4276 6312
rect 4348 6311 4384 6312
rect 4240 6305 4384 6311
rect 4240 6303 4306 6305
rect 4240 6283 4248 6303
rect 4268 6284 4306 6303
rect 4328 6303 4384 6305
rect 4328 6284 4356 6303
rect 4268 6283 4356 6284
rect 4376 6283 4384 6303
rect 4240 6277 4384 6283
rect 4450 6307 4488 6315
rect 4556 6311 4592 6312
rect 4450 6287 4459 6307
rect 4479 6287 4488 6307
rect 4450 6278 4488 6287
rect 4507 6304 4592 6311
rect 4507 6284 4514 6304
rect 4535 6303 4592 6304
rect 4535 6284 4564 6303
rect 4507 6283 4564 6284
rect 4584 6283 4592 6303
rect 4450 6277 4487 6278
rect 4507 6277 4592 6283
rect 4658 6307 4696 6315
rect 4769 6311 4805 6312
rect 4658 6287 4667 6307
rect 4687 6287 4696 6307
rect 4658 6278 4696 6287
rect 4720 6303 4805 6311
rect 4720 6283 4777 6303
rect 4797 6283 4805 6303
rect 4658 6277 4695 6278
rect 4720 6277 4805 6283
rect 4871 6307 4909 6315
rect 4871 6287 4880 6307
rect 4900 6287 4909 6307
rect 4871 6278 4909 6287
rect 5050 6314 5086 6349
rect 5403 6345 5438 6391
rect 6814 6389 6851 6460
rect 6966 6399 6997 6400
rect 6814 6369 6823 6389
rect 6843 6369 6851 6389
rect 6814 6359 6851 6369
rect 6910 6389 6997 6399
rect 6910 6369 6919 6389
rect 6939 6369 6997 6389
rect 6910 6360 6997 6369
rect 6910 6359 6947 6360
rect 5401 6336 5438 6345
rect 5401 6318 5411 6336
rect 5429 6318 5438 6336
rect 5050 6304 5087 6314
rect 5401 6308 5438 6318
rect 6966 6307 6997 6360
rect 7027 6389 7064 6460
rect 7235 6465 7628 6485
rect 7648 6465 7651 6485
rect 7235 6460 7651 6465
rect 7235 6459 7576 6460
rect 7179 6399 7210 6400
rect 7027 6369 7036 6389
rect 7056 6369 7064 6389
rect 7027 6359 7064 6369
rect 7123 6392 7210 6399
rect 7123 6389 7184 6392
rect 7123 6369 7132 6389
rect 7152 6372 7184 6389
rect 7205 6372 7210 6392
rect 7152 6369 7210 6372
rect 7123 6362 7210 6369
rect 7235 6389 7272 6459
rect 7538 6458 7575 6459
rect 7387 6399 7423 6400
rect 7235 6369 7244 6389
rect 7264 6369 7272 6389
rect 7123 6360 7179 6362
rect 7123 6359 7160 6360
rect 7235 6359 7272 6369
rect 7331 6389 7479 6399
rect 7579 6396 7675 6398
rect 7331 6369 7340 6389
rect 7360 6369 7450 6389
rect 7470 6369 7479 6389
rect 7331 6360 7479 6369
rect 7537 6389 7675 6396
rect 7537 6369 7546 6389
rect 7566 6369 7675 6389
rect 7537 6360 7675 6369
rect 7331 6359 7368 6360
rect 7387 6308 7423 6360
rect 7442 6359 7479 6360
rect 7538 6359 7575 6360
rect 6858 6306 6899 6307
rect 5050 6286 5060 6304
rect 5078 6286 5087 6304
rect 4871 6277 4908 6278
rect 5050 6277 5087 6286
rect 6750 6299 6899 6306
rect 6750 6279 6868 6299
rect 6888 6279 6899 6299
rect 4294 6256 4330 6277
rect 4720 6256 4751 6277
rect 6750 6271 6899 6279
rect 6966 6303 7325 6307
rect 6966 6298 7288 6303
rect 6966 6274 7079 6298
rect 7103 6279 7288 6298
rect 7312 6279 7325 6303
rect 7103 6274 7325 6279
rect 6966 6271 7325 6274
rect 7387 6271 7422 6308
rect 7490 6305 7590 6308
rect 7490 6301 7557 6305
rect 7490 6275 7502 6301
rect 7528 6279 7557 6301
rect 7583 6279 7590 6305
rect 7528 6275 7590 6279
rect 7490 6271 7590 6275
rect 4127 6252 4227 6256
rect 4127 6248 4189 6252
rect 4127 6222 4134 6248
rect 4160 6226 4189 6248
rect 4215 6226 4227 6252
rect 4160 6222 4227 6226
rect 4127 6219 4227 6222
rect 4295 6219 4330 6256
rect 4392 6253 4751 6256
rect 4392 6248 4614 6253
rect 4392 6224 4405 6248
rect 4429 6229 4614 6248
rect 4638 6229 4751 6253
rect 4429 6224 4751 6229
rect 4392 6220 4751 6224
rect 4818 6248 4967 6256
rect 6966 6250 6997 6271
rect 7387 6250 7423 6271
rect 6809 6249 6846 6250
rect 4818 6228 4829 6248
rect 4849 6228 4967 6248
rect 5404 6244 5441 6246
rect 5404 6243 6052 6244
rect 4818 6221 4967 6228
rect 5403 6237 6052 6243
rect 4818 6220 4859 6221
rect 4142 6167 4179 6168
rect 4238 6167 4275 6168
rect 4294 6167 4330 6219
rect 4349 6167 4386 6168
rect 4042 6158 4180 6167
rect 2978 6140 3009 6143
rect 2978 6114 2985 6140
rect 3004 6114 3009 6140
rect 2978 5720 3009 6114
rect 3030 6139 3198 6140
rect 3030 6136 3474 6139
rect 3030 6117 3405 6136
rect 3425 6117 3474 6136
rect 4042 6138 4151 6158
rect 4171 6138 4180 6158
rect 3030 6113 3474 6117
rect 3030 6111 3198 6113
rect 3030 5933 3057 6111
rect 3097 6073 3161 6085
rect 3437 6081 3474 6113
rect 3645 6112 3894 6134
rect 4042 6131 4180 6138
rect 4238 6158 4386 6167
rect 4238 6138 4247 6158
rect 4267 6138 4357 6158
rect 4377 6138 4386 6158
rect 4042 6129 4138 6131
rect 4238 6128 4386 6138
rect 4445 6158 4482 6168
rect 4557 6167 4594 6168
rect 4538 6165 4594 6167
rect 4445 6138 4453 6158
rect 4473 6138 4482 6158
rect 4294 6127 4330 6128
rect 3645 6081 3682 6112
rect 3858 6110 3894 6112
rect 3858 6081 3895 6110
rect 3097 6072 3132 6073
rect 3074 6067 3132 6072
rect 3074 6047 3077 6067
rect 3097 6053 3132 6067
rect 3152 6053 3161 6073
rect 3097 6045 3161 6053
rect 3123 6044 3161 6045
rect 3124 6043 3161 6044
rect 3227 6077 3263 6078
rect 3335 6077 3371 6078
rect 3227 6069 3371 6077
rect 3227 6049 3235 6069
rect 3255 6068 3343 6069
rect 3255 6049 3288 6068
rect 3227 6048 3288 6049
rect 3312 6049 3343 6068
rect 3363 6049 3371 6069
rect 3312 6048 3371 6049
rect 3227 6043 3371 6048
rect 3437 6073 3475 6081
rect 3543 6077 3579 6078
rect 3437 6053 3446 6073
rect 3466 6053 3475 6073
rect 3437 6044 3475 6053
rect 3494 6070 3579 6077
rect 3494 6050 3501 6070
rect 3522 6069 3579 6070
rect 3522 6050 3551 6069
rect 3494 6049 3551 6050
rect 3571 6049 3579 6069
rect 3437 6043 3474 6044
rect 3494 6043 3579 6049
rect 3645 6073 3683 6081
rect 3756 6077 3792 6078
rect 3645 6053 3654 6073
rect 3674 6053 3683 6073
rect 3645 6044 3683 6053
rect 3707 6069 3792 6077
rect 3707 6049 3764 6069
rect 3784 6049 3792 6069
rect 3645 6043 3682 6044
rect 3707 6043 3792 6049
rect 3858 6073 3896 6081
rect 3858 6053 3867 6073
rect 3887 6053 3896 6073
rect 4142 6068 4179 6069
rect 4445 6068 4482 6138
rect 4507 6158 4594 6165
rect 4507 6155 4565 6158
rect 4507 6135 4512 6155
rect 4533 6138 4565 6155
rect 4585 6138 4594 6158
rect 4533 6135 4594 6138
rect 4507 6128 4594 6135
rect 4653 6158 4690 6168
rect 4653 6138 4661 6158
rect 4681 6138 4690 6158
rect 4507 6127 4538 6128
rect 4141 6067 4482 6068
rect 3858 6044 3896 6053
rect 4066 6062 4482 6067
rect 3858 6043 3895 6044
rect 3281 6022 3317 6043
rect 3707 6022 3738 6043
rect 4066 6042 4069 6062
rect 4089 6042 4482 6062
rect 4653 6067 4690 6138
rect 4720 6167 4751 6220
rect 5403 6219 5413 6237
rect 5431 6223 6052 6237
rect 5431 6219 5441 6223
rect 5882 6222 6052 6223
rect 5053 6205 5090 6215
rect 5053 6187 5062 6205
rect 5080 6187 5090 6205
rect 5053 6178 5090 6187
rect 5403 6209 5441 6219
rect 4770 6167 4807 6168
rect 4720 6158 4807 6167
rect 4720 6138 4778 6158
rect 4798 6138 4807 6158
rect 4720 6128 4807 6138
rect 4866 6158 4903 6168
rect 4866 6138 4874 6158
rect 4894 6138 4903 6158
rect 4720 6127 4751 6128
rect 4866 6067 4903 6138
rect 5058 6113 5089 6178
rect 5403 6131 5438 6209
rect 6015 6199 6052 6222
rect 6808 6240 6846 6249
rect 6808 6220 6817 6240
rect 6837 6220 6846 6240
rect 6808 6212 6846 6220
rect 6912 6244 6997 6250
rect 7022 6249 7059 6250
rect 6912 6224 6920 6244
rect 6940 6224 6997 6244
rect 6912 6216 6997 6224
rect 7021 6240 7059 6249
rect 7021 6220 7030 6240
rect 7050 6220 7059 6240
rect 6912 6215 6948 6216
rect 7021 6212 7059 6220
rect 7125 6244 7210 6250
rect 7230 6249 7267 6250
rect 7125 6224 7133 6244
rect 7153 6243 7210 6244
rect 7153 6224 7182 6243
rect 7125 6223 7182 6224
rect 7203 6223 7210 6243
rect 7125 6216 7210 6223
rect 7229 6240 7267 6249
rect 7229 6220 7238 6240
rect 7258 6220 7267 6240
rect 7125 6215 7161 6216
rect 7229 6212 7267 6220
rect 7333 6248 7477 6250
rect 7333 6244 7391 6248
rect 7333 6224 7341 6244
rect 7361 6224 7391 6244
rect 7333 6222 7391 6224
rect 7416 6244 7477 6248
rect 7416 6224 7449 6244
rect 7469 6224 7477 6244
rect 7416 6222 7477 6224
rect 7333 6216 7477 6222
rect 7333 6215 7369 6216
rect 7441 6215 7477 6216
rect 7543 6249 7580 6250
rect 7543 6248 7581 6249
rect 7543 6240 7607 6248
rect 7543 6220 7552 6240
rect 7572 6226 7607 6240
rect 7627 6226 7630 6246
rect 7572 6221 7630 6226
rect 7572 6220 7607 6221
rect 5399 6122 5438 6131
rect 5057 6103 5094 6113
rect 5057 6101 5067 6103
rect 4991 6099 5067 6101
rect 4653 6043 4903 6067
rect 4988 6085 5067 6099
rect 5085 6085 5094 6103
rect 5399 6104 5409 6122
rect 5427 6104 5438 6122
rect 5399 6098 5438 6104
rect 5594 6174 5844 6198
rect 5594 6103 5631 6174
rect 5746 6113 5777 6114
rect 5399 6094 5436 6098
rect 4988 6082 5094 6085
rect 4460 6023 4481 6042
rect 4988 6023 5014 6082
rect 5057 6076 5094 6082
rect 5594 6083 5603 6103
rect 5623 6083 5631 6103
rect 5594 6073 5631 6083
rect 5690 6103 5777 6113
rect 5690 6083 5699 6103
rect 5719 6083 5777 6103
rect 5690 6074 5777 6083
rect 5690 6073 5727 6074
rect 5402 6023 5439 6032
rect 3114 6018 3214 6022
rect 3114 6014 3176 6018
rect 3114 5988 3121 6014
rect 3147 5992 3176 6014
rect 3202 5992 3214 6018
rect 3147 5988 3214 5992
rect 3114 5985 3214 5988
rect 3282 5985 3317 6022
rect 3379 6019 3738 6022
rect 3379 6014 3601 6019
rect 3379 5990 3392 6014
rect 3416 5995 3601 6014
rect 3625 5995 3738 6019
rect 3416 5990 3738 5995
rect 3379 5986 3738 5990
rect 3805 6014 3954 6022
rect 3805 5994 3816 6014
rect 3836 5994 3954 6014
rect 4460 6005 5014 6023
rect 5060 6012 5097 6014
rect 4988 6004 5014 6005
rect 5057 6004 5097 6012
rect 3805 5987 3954 5994
rect 5057 5992 5069 6004
rect 5048 5987 5069 5992
rect 3805 5986 3846 5987
rect 4464 5986 5069 5987
rect 5087 5986 5097 6004
rect 3129 5933 3166 5934
rect 3225 5933 3262 5934
rect 3281 5933 3317 5985
rect 3336 5933 3373 5934
rect 3029 5924 3167 5933
rect 3029 5904 3138 5924
rect 3158 5904 3167 5924
rect 3029 5897 3167 5904
rect 3225 5924 3373 5933
rect 3225 5904 3234 5924
rect 3254 5904 3344 5924
rect 3364 5904 3373 5924
rect 3029 5895 3125 5897
rect 3225 5894 3373 5904
rect 3432 5924 3469 5934
rect 3544 5933 3581 5934
rect 3525 5931 3581 5933
rect 3432 5904 3440 5924
rect 3460 5904 3469 5924
rect 3281 5893 3317 5894
rect 3129 5834 3166 5835
rect 3432 5834 3469 5904
rect 3494 5924 3581 5931
rect 3494 5921 3552 5924
rect 3494 5901 3499 5921
rect 3520 5904 3552 5921
rect 3572 5904 3581 5924
rect 3520 5901 3581 5904
rect 3494 5894 3581 5901
rect 3640 5924 3677 5934
rect 3640 5904 3648 5924
rect 3668 5904 3677 5924
rect 3494 5893 3525 5894
rect 3128 5833 3469 5834
rect 3053 5828 3469 5833
rect 3053 5808 3056 5828
rect 3076 5808 3469 5828
rect 3640 5833 3677 5904
rect 3707 5933 3738 5986
rect 4464 5977 5097 5986
rect 5400 6005 5411 6023
rect 5429 6005 5439 6023
rect 5746 6021 5777 6074
rect 5807 6103 5844 6174
rect 6015 6179 6408 6199
rect 6428 6179 6431 6199
rect 6809 6183 6846 6212
rect 6015 6174 6431 6179
rect 6810 6181 6846 6183
rect 7022 6181 7059 6212
rect 6015 6173 6356 6174
rect 5959 6113 5990 6114
rect 5807 6083 5816 6103
rect 5836 6083 5844 6103
rect 5807 6073 5844 6083
rect 5903 6106 5990 6113
rect 5903 6103 5964 6106
rect 5903 6083 5912 6103
rect 5932 6086 5964 6103
rect 5985 6086 5990 6106
rect 5932 6083 5990 6086
rect 5903 6076 5990 6083
rect 6015 6103 6052 6173
rect 6318 6172 6355 6173
rect 6810 6159 7059 6181
rect 7230 6180 7267 6212
rect 7543 6208 7607 6220
rect 7647 6182 7674 6360
rect 7506 6180 7674 6182
rect 7230 6154 7674 6180
rect 7506 6153 7674 6154
rect 6167 6113 6203 6114
rect 6015 6083 6024 6103
rect 6044 6083 6052 6103
rect 5903 6074 5959 6076
rect 5903 6073 5940 6074
rect 6015 6073 6052 6083
rect 6111 6103 6259 6113
rect 6359 6110 6455 6112
rect 6111 6083 6120 6103
rect 6140 6083 6230 6103
rect 6250 6083 6259 6103
rect 6111 6074 6259 6083
rect 6317 6103 6455 6110
rect 6317 6083 6326 6103
rect 6346 6083 6455 6103
rect 6317 6074 6455 6083
rect 6111 6073 6148 6074
rect 6167 6022 6203 6074
rect 6222 6073 6259 6074
rect 6318 6073 6355 6074
rect 5638 6020 5679 6021
rect 4464 5970 5096 5977
rect 4464 5968 4526 5970
rect 4042 5958 4210 5959
rect 4464 5958 4486 5968
rect 3757 5933 3794 5934
rect 3707 5924 3794 5933
rect 3707 5904 3765 5924
rect 3785 5904 3794 5924
rect 3707 5894 3794 5904
rect 3853 5924 3890 5934
rect 3853 5904 3861 5924
rect 3881 5904 3890 5924
rect 3707 5893 3738 5894
rect 3853 5833 3890 5904
rect 3640 5809 3890 5833
rect 4042 5932 4486 5958
rect 4042 5930 4210 5932
rect 4042 5752 4069 5930
rect 4109 5892 4173 5904
rect 4449 5900 4486 5932
rect 4657 5931 4906 5953
rect 4657 5900 4694 5931
rect 4870 5929 4906 5931
rect 4870 5900 4907 5929
rect 4109 5891 4144 5892
rect 4086 5886 4144 5891
rect 4086 5866 4089 5886
rect 4109 5872 4144 5886
rect 4164 5872 4173 5892
rect 4109 5864 4173 5872
rect 4135 5863 4173 5864
rect 4136 5862 4173 5863
rect 4239 5896 4275 5897
rect 4347 5896 4383 5897
rect 4239 5888 4383 5896
rect 4239 5868 4247 5888
rect 4267 5868 4296 5888
rect 4239 5867 4296 5868
rect 4318 5868 4355 5888
rect 4375 5868 4383 5888
rect 4318 5867 4383 5868
rect 4239 5862 4383 5867
rect 4449 5892 4487 5900
rect 4555 5896 4591 5897
rect 4449 5872 4458 5892
rect 4478 5872 4487 5892
rect 4449 5863 4487 5872
rect 4506 5889 4591 5896
rect 4506 5869 4513 5889
rect 4534 5888 4591 5889
rect 4534 5869 4563 5888
rect 4506 5868 4563 5869
rect 4583 5868 4591 5888
rect 4449 5862 4486 5863
rect 4506 5862 4591 5868
rect 4657 5892 4695 5900
rect 4768 5896 4804 5897
rect 4657 5872 4666 5892
rect 4686 5872 4695 5892
rect 4657 5863 4695 5872
rect 4719 5888 4804 5896
rect 4719 5868 4776 5888
rect 4796 5868 4804 5888
rect 4657 5862 4694 5863
rect 4719 5862 4804 5868
rect 4870 5892 4908 5900
rect 4870 5872 4879 5892
rect 4899 5872 4908 5892
rect 4870 5863 4908 5872
rect 4870 5862 4907 5863
rect 4293 5841 4329 5862
rect 4719 5841 4750 5862
rect 4126 5837 4226 5841
rect 4126 5833 4188 5837
rect 4126 5807 4133 5833
rect 4159 5811 4188 5833
rect 4214 5811 4226 5837
rect 4159 5807 4226 5811
rect 4126 5804 4226 5807
rect 4294 5804 4329 5841
rect 4391 5838 4750 5841
rect 4391 5833 4613 5838
rect 4391 5809 4404 5833
rect 4428 5814 4613 5833
rect 4637 5814 4750 5838
rect 4428 5809 4750 5814
rect 4391 5805 4750 5809
rect 4817 5833 4966 5841
rect 4817 5813 4828 5833
rect 4848 5813 4966 5833
rect 4817 5806 4966 5813
rect 5057 5821 5096 5970
rect 5400 5856 5439 6005
rect 5530 6013 5679 6020
rect 5530 5993 5648 6013
rect 5668 5993 5679 6013
rect 5530 5985 5679 5993
rect 5746 6017 6105 6021
rect 5746 6012 6068 6017
rect 5746 5988 5859 6012
rect 5883 5993 6068 6012
rect 6092 5993 6105 6017
rect 5883 5988 6105 5993
rect 5746 5985 6105 5988
rect 6167 5985 6202 6022
rect 6270 6019 6370 6022
rect 6270 6015 6337 6019
rect 6270 5989 6282 6015
rect 6308 5993 6337 6015
rect 6363 5993 6370 6019
rect 6308 5989 6370 5993
rect 6270 5985 6370 5989
rect 5746 5964 5777 5985
rect 6167 5964 6203 5985
rect 5589 5963 5626 5964
rect 5588 5954 5626 5963
rect 5588 5934 5597 5954
rect 5617 5934 5626 5954
rect 5588 5926 5626 5934
rect 5692 5958 5777 5964
rect 5802 5963 5839 5964
rect 5692 5938 5700 5958
rect 5720 5938 5777 5958
rect 5692 5930 5777 5938
rect 5801 5954 5839 5963
rect 5801 5934 5810 5954
rect 5830 5934 5839 5954
rect 5692 5929 5728 5930
rect 5801 5926 5839 5934
rect 5905 5958 5990 5964
rect 6010 5963 6047 5964
rect 5905 5938 5913 5958
rect 5933 5957 5990 5958
rect 5933 5938 5962 5957
rect 5905 5937 5962 5938
rect 5983 5937 5990 5957
rect 5905 5930 5990 5937
rect 6009 5954 6047 5963
rect 6009 5934 6018 5954
rect 6038 5934 6047 5954
rect 5905 5929 5941 5930
rect 6009 5926 6047 5934
rect 6113 5959 6257 5964
rect 6113 5958 6178 5959
rect 6113 5938 6121 5958
rect 6141 5938 6178 5958
rect 6200 5958 6257 5959
rect 6200 5938 6229 5958
rect 6249 5938 6257 5958
rect 6113 5930 6257 5938
rect 6113 5929 6149 5930
rect 6221 5929 6257 5930
rect 6323 5963 6360 5964
rect 6323 5962 6361 5963
rect 6323 5954 6387 5962
rect 6323 5934 6332 5954
rect 6352 5940 6387 5954
rect 6407 5940 6410 5960
rect 6352 5935 6410 5940
rect 6352 5934 6387 5935
rect 5589 5897 5626 5926
rect 5590 5895 5626 5897
rect 5802 5895 5839 5926
rect 5590 5873 5839 5895
rect 6010 5894 6047 5926
rect 6323 5922 6387 5934
rect 6427 5896 6454 6074
rect 6286 5894 6454 5896
rect 6010 5868 6454 5894
rect 6606 5993 6856 6017
rect 6606 5922 6643 5993
rect 6758 5932 6789 5933
rect 6606 5902 6615 5922
rect 6635 5902 6643 5922
rect 6606 5892 6643 5902
rect 6702 5922 6789 5932
rect 6702 5902 6711 5922
rect 6731 5902 6789 5922
rect 6702 5893 6789 5902
rect 6702 5892 6739 5893
rect 6010 5858 6032 5868
rect 6286 5867 6454 5868
rect 5970 5856 6032 5858
rect 5400 5849 6032 5856
rect 4817 5805 4858 5806
rect 4141 5752 4178 5753
rect 4237 5752 4274 5753
rect 4293 5752 4329 5804
rect 4348 5752 4385 5753
rect 4041 5743 4179 5752
rect 4041 5723 4150 5743
rect 4170 5723 4179 5743
rect 2978 5719 3148 5720
rect 2978 5704 3424 5719
rect 4041 5716 4179 5723
rect 4237 5743 4385 5752
rect 4237 5723 4246 5743
rect 4266 5723 4356 5743
rect 4376 5723 4385 5743
rect 4041 5714 4137 5716
rect 2980 5693 3424 5704
rect 2980 5691 3148 5693
rect 2980 5513 3007 5691
rect 3047 5653 3111 5665
rect 3387 5661 3424 5693
rect 3595 5692 3844 5714
rect 4237 5713 4385 5723
rect 4444 5743 4481 5753
rect 4556 5752 4593 5753
rect 4537 5750 4593 5752
rect 4444 5723 4452 5743
rect 4472 5723 4481 5743
rect 4293 5712 4329 5713
rect 3595 5661 3632 5692
rect 3808 5690 3844 5692
rect 3808 5661 3845 5690
rect 3047 5652 3082 5653
rect 3024 5647 3082 5652
rect 3024 5627 3027 5647
rect 3047 5633 3082 5647
rect 3102 5633 3111 5653
rect 3047 5625 3111 5633
rect 3073 5624 3111 5625
rect 3074 5623 3111 5624
rect 3177 5657 3213 5658
rect 3285 5657 3321 5658
rect 3177 5649 3321 5657
rect 3177 5629 3185 5649
rect 3205 5648 3293 5649
rect 3205 5631 3233 5648
rect 3257 5631 3293 5648
rect 3205 5629 3293 5631
rect 3313 5629 3321 5649
rect 3177 5623 3321 5629
rect 3387 5653 3425 5661
rect 3493 5657 3529 5658
rect 3387 5633 3396 5653
rect 3416 5633 3425 5653
rect 3387 5624 3425 5633
rect 3444 5650 3529 5657
rect 3444 5630 3451 5650
rect 3472 5649 3529 5650
rect 3472 5630 3501 5649
rect 3444 5629 3501 5630
rect 3521 5629 3529 5649
rect 3387 5623 3424 5624
rect 3444 5623 3529 5629
rect 3595 5653 3633 5661
rect 3706 5657 3742 5658
rect 3595 5633 3604 5653
rect 3624 5633 3633 5653
rect 3595 5624 3633 5633
rect 3657 5649 3742 5657
rect 3657 5629 3714 5649
rect 3734 5629 3742 5649
rect 3595 5623 3632 5624
rect 3657 5623 3742 5629
rect 3808 5653 3846 5661
rect 4141 5653 4178 5654
rect 4444 5653 4481 5723
rect 4506 5743 4593 5750
rect 4506 5740 4564 5743
rect 4506 5720 4511 5740
rect 4532 5723 4564 5740
rect 4584 5723 4593 5743
rect 4532 5720 4593 5723
rect 4506 5713 4593 5720
rect 4652 5743 4689 5753
rect 4652 5723 4660 5743
rect 4680 5723 4689 5743
rect 4506 5712 4537 5713
rect 3808 5633 3817 5653
rect 3837 5633 3846 5653
rect 4140 5652 4481 5653
rect 3808 5624 3846 5633
rect 4065 5647 4481 5652
rect 4065 5627 4068 5647
rect 4088 5627 4481 5647
rect 4652 5652 4689 5723
rect 4719 5752 4750 5805
rect 5057 5803 5067 5821
rect 5085 5803 5096 5821
rect 5399 5840 6032 5849
rect 6758 5840 6789 5893
rect 6819 5922 6856 5993
rect 7027 5998 7420 6018
rect 7440 5998 7443 6018
rect 7027 5993 7443 5998
rect 7027 5992 7368 5993
rect 6971 5932 7002 5933
rect 6819 5902 6828 5922
rect 6848 5902 6856 5922
rect 6819 5892 6856 5902
rect 6915 5925 7002 5932
rect 6915 5922 6976 5925
rect 6915 5902 6924 5922
rect 6944 5905 6976 5922
rect 6997 5905 7002 5925
rect 6944 5902 7002 5905
rect 6915 5895 7002 5902
rect 7027 5922 7064 5992
rect 7330 5991 7367 5992
rect 7179 5932 7215 5933
rect 7027 5902 7036 5922
rect 7056 5902 7064 5922
rect 6915 5893 6971 5895
rect 6915 5892 6952 5893
rect 7027 5892 7064 5902
rect 7123 5922 7271 5932
rect 7371 5929 7467 5931
rect 7123 5902 7132 5922
rect 7152 5902 7242 5922
rect 7262 5902 7271 5922
rect 7123 5893 7271 5902
rect 7329 5922 7467 5929
rect 7329 5902 7338 5922
rect 7358 5902 7467 5922
rect 7329 5893 7467 5902
rect 7123 5892 7160 5893
rect 7179 5841 7215 5893
rect 7234 5892 7271 5893
rect 7330 5892 7367 5893
rect 5399 5822 5409 5840
rect 5427 5839 6032 5840
rect 6650 5839 6691 5840
rect 5427 5834 5448 5839
rect 5427 5822 5439 5834
rect 6542 5832 6691 5839
rect 5399 5814 5439 5822
rect 5482 5821 5508 5822
rect 5399 5812 5436 5814
rect 5482 5803 6036 5821
rect 6542 5812 6660 5832
rect 6680 5812 6691 5832
rect 6542 5804 6691 5812
rect 6758 5836 7117 5840
rect 6758 5831 7080 5836
rect 6758 5807 6871 5831
rect 6895 5812 7080 5831
rect 7104 5812 7117 5836
rect 6895 5807 7117 5812
rect 6758 5804 7117 5807
rect 7179 5804 7214 5841
rect 7282 5838 7382 5841
rect 7282 5834 7349 5838
rect 7282 5808 7294 5834
rect 7320 5812 7349 5834
rect 7375 5812 7382 5838
rect 7320 5808 7382 5812
rect 7282 5804 7382 5808
rect 5057 5794 5094 5803
rect 4769 5752 4806 5753
rect 4719 5743 4806 5752
rect 4719 5723 4777 5743
rect 4797 5723 4806 5743
rect 4719 5713 4806 5723
rect 4865 5743 4902 5753
rect 4865 5723 4873 5743
rect 4893 5723 4902 5743
rect 5402 5744 5439 5750
rect 5482 5744 5508 5803
rect 6015 5784 6036 5803
rect 5402 5741 5508 5744
rect 5060 5728 5097 5732
rect 4719 5712 4750 5713
rect 4865 5652 4902 5723
rect 4652 5628 4902 5652
rect 5058 5722 5097 5728
rect 5058 5704 5069 5722
rect 5087 5704 5097 5722
rect 5402 5723 5411 5741
rect 5429 5727 5508 5741
rect 5593 5759 5843 5783
rect 5429 5725 5505 5727
rect 5429 5723 5439 5725
rect 5402 5713 5439 5723
rect 5058 5695 5097 5704
rect 3808 5623 3845 5624
rect 3231 5602 3267 5623
rect 3657 5602 3688 5623
rect 4444 5604 4481 5627
rect 5058 5617 5093 5695
rect 5407 5648 5438 5713
rect 5593 5688 5630 5759
rect 5745 5698 5776 5699
rect 5593 5668 5602 5688
rect 5622 5668 5630 5688
rect 5593 5658 5630 5668
rect 5689 5688 5776 5698
rect 5689 5668 5698 5688
rect 5718 5668 5776 5688
rect 5689 5659 5776 5668
rect 5689 5658 5726 5659
rect 5055 5607 5093 5617
rect 5406 5639 5443 5648
rect 5406 5621 5416 5639
rect 5434 5621 5443 5639
rect 5406 5611 5443 5621
rect 4444 5603 4614 5604
rect 5055 5603 5065 5607
rect 3064 5598 3164 5602
rect 3064 5594 3126 5598
rect 3064 5568 3071 5594
rect 3097 5572 3126 5594
rect 3152 5572 3164 5598
rect 3097 5568 3164 5572
rect 3064 5565 3164 5568
rect 3232 5565 3267 5602
rect 3329 5599 3688 5602
rect 3329 5594 3551 5599
rect 3329 5570 3342 5594
rect 3366 5575 3551 5594
rect 3575 5575 3688 5599
rect 3366 5570 3688 5575
rect 3329 5566 3688 5570
rect 3755 5594 3904 5602
rect 3755 5574 3766 5594
rect 3786 5574 3904 5594
rect 4444 5589 5065 5603
rect 5083 5589 5093 5607
rect 5745 5606 5776 5659
rect 5806 5688 5843 5759
rect 6014 5764 6407 5784
rect 6427 5764 6430 5784
rect 6758 5783 6789 5804
rect 7179 5783 7215 5804
rect 6601 5782 6638 5783
rect 6014 5759 6430 5764
rect 6600 5773 6638 5782
rect 6014 5758 6355 5759
rect 5958 5698 5989 5699
rect 5806 5668 5815 5688
rect 5835 5668 5843 5688
rect 5806 5658 5843 5668
rect 5902 5691 5989 5698
rect 5902 5688 5963 5691
rect 5902 5668 5911 5688
rect 5931 5671 5963 5688
rect 5984 5671 5989 5691
rect 5931 5668 5989 5671
rect 5902 5661 5989 5668
rect 6014 5688 6051 5758
rect 6317 5757 6354 5758
rect 6600 5753 6609 5773
rect 6629 5753 6638 5773
rect 6600 5745 6638 5753
rect 6704 5777 6789 5783
rect 6814 5782 6851 5783
rect 6704 5757 6712 5777
rect 6732 5757 6789 5777
rect 6704 5749 6789 5757
rect 6813 5773 6851 5782
rect 6813 5753 6822 5773
rect 6842 5753 6851 5773
rect 6704 5748 6740 5749
rect 6813 5745 6851 5753
rect 6917 5777 7002 5783
rect 7022 5782 7059 5783
rect 6917 5757 6925 5777
rect 6945 5776 7002 5777
rect 6945 5757 6974 5776
rect 6917 5756 6974 5757
rect 6995 5756 7002 5776
rect 6917 5749 7002 5756
rect 7021 5773 7059 5782
rect 7021 5753 7030 5773
rect 7050 5753 7059 5773
rect 6917 5748 6953 5749
rect 7021 5745 7059 5753
rect 7125 5777 7269 5783
rect 7125 5757 7133 5777
rect 7153 5757 7185 5777
rect 7209 5757 7241 5777
rect 7261 5757 7269 5777
rect 7125 5749 7269 5757
rect 7125 5748 7161 5749
rect 7233 5748 7269 5749
rect 7335 5782 7372 5783
rect 7335 5781 7373 5782
rect 7335 5773 7399 5781
rect 7335 5753 7344 5773
rect 7364 5759 7399 5773
rect 7419 5759 7422 5779
rect 7364 5754 7422 5759
rect 7364 5753 7399 5754
rect 6601 5716 6638 5745
rect 6602 5714 6638 5716
rect 6814 5714 6851 5745
rect 6166 5698 6202 5699
rect 6014 5668 6023 5688
rect 6043 5668 6051 5688
rect 5902 5659 5958 5661
rect 5902 5658 5939 5659
rect 6014 5658 6051 5668
rect 6110 5688 6258 5698
rect 6358 5695 6454 5697
rect 6110 5668 6119 5688
rect 6139 5668 6229 5688
rect 6249 5668 6258 5688
rect 6110 5659 6258 5668
rect 6316 5688 6454 5695
rect 6602 5692 6851 5714
rect 7022 5713 7059 5745
rect 7335 5741 7399 5753
rect 7439 5715 7466 5893
rect 7298 5713 7466 5715
rect 7022 5709 7466 5713
rect 6316 5668 6325 5688
rect 6345 5668 6454 5688
rect 7022 5690 7071 5709
rect 7091 5690 7466 5709
rect 7022 5687 7466 5690
rect 7298 5686 7466 5687
rect 6316 5659 6454 5668
rect 6110 5658 6147 5659
rect 6166 5607 6202 5659
rect 6221 5658 6258 5659
rect 6317 5658 6354 5659
rect 5637 5605 5678 5606
rect 4444 5583 5093 5589
rect 5529 5598 5678 5605
rect 4444 5582 5092 5583
rect 5055 5580 5092 5582
rect 3755 5567 3904 5574
rect 5529 5578 5647 5598
rect 5667 5578 5678 5598
rect 5529 5570 5678 5578
rect 5745 5602 6104 5606
rect 5745 5597 6067 5602
rect 5745 5573 5858 5597
rect 5882 5578 6067 5597
rect 6091 5578 6104 5602
rect 5882 5573 6104 5578
rect 5745 5570 6104 5573
rect 6166 5570 6201 5607
rect 6269 5604 6369 5607
rect 6269 5600 6336 5604
rect 6269 5574 6281 5600
rect 6307 5578 6336 5600
rect 6362 5578 6369 5604
rect 6307 5574 6369 5578
rect 6269 5570 6369 5574
rect 3755 5566 3796 5567
rect 3079 5513 3116 5514
rect 3175 5513 3212 5514
rect 3231 5513 3267 5565
rect 3286 5513 3323 5514
rect 2979 5504 3117 5513
rect 2979 5484 3088 5504
rect 3108 5484 3117 5504
rect 2979 5477 3117 5484
rect 3175 5504 3323 5513
rect 3175 5484 3184 5504
rect 3204 5484 3294 5504
rect 3314 5484 3323 5504
rect 2979 5475 3075 5477
rect 3175 5474 3323 5484
rect 3382 5504 3419 5514
rect 3494 5513 3531 5514
rect 3475 5511 3531 5513
rect 3382 5484 3390 5504
rect 3410 5484 3419 5504
rect 3231 5473 3267 5474
rect 3079 5414 3116 5415
rect 3382 5414 3419 5484
rect 3444 5504 3531 5511
rect 3444 5501 3502 5504
rect 3444 5481 3449 5501
rect 3470 5484 3502 5501
rect 3522 5484 3531 5504
rect 3470 5481 3531 5484
rect 3444 5474 3531 5481
rect 3590 5504 3627 5514
rect 3590 5484 3598 5504
rect 3618 5484 3627 5504
rect 3444 5473 3475 5474
rect 3078 5413 3419 5414
rect 3003 5408 3419 5413
rect 3003 5388 3006 5408
rect 3026 5388 3419 5408
rect 3590 5413 3627 5484
rect 3657 5513 3688 5566
rect 5745 5549 5776 5570
rect 6166 5549 6202 5570
rect 5409 5540 5446 5549
rect 5588 5548 5625 5549
rect 5409 5522 5418 5540
rect 5436 5522 5446 5540
rect 3707 5513 3744 5514
rect 3657 5504 3744 5513
rect 3657 5484 3715 5504
rect 3735 5484 3744 5504
rect 3657 5474 3744 5484
rect 3803 5504 3840 5514
rect 3803 5484 3811 5504
rect 3831 5484 3840 5504
rect 3657 5473 3688 5474
rect 3803 5413 3840 5484
rect 5058 5508 5095 5518
rect 5409 5512 5446 5522
rect 5058 5490 5067 5508
rect 5085 5490 5095 5508
rect 5058 5481 5095 5490
rect 5058 5457 5093 5481
rect 5410 5477 5446 5512
rect 5587 5539 5625 5548
rect 5587 5519 5596 5539
rect 5616 5519 5625 5539
rect 5587 5511 5625 5519
rect 5691 5543 5776 5549
rect 5801 5548 5838 5549
rect 5691 5523 5699 5543
rect 5719 5523 5776 5543
rect 5691 5515 5776 5523
rect 5800 5539 5838 5548
rect 5800 5519 5809 5539
rect 5829 5519 5838 5539
rect 5691 5514 5727 5515
rect 5800 5511 5838 5519
rect 5904 5543 5989 5549
rect 6009 5548 6046 5549
rect 5904 5523 5912 5543
rect 5932 5542 5989 5543
rect 5932 5523 5961 5542
rect 5904 5522 5961 5523
rect 5982 5522 5989 5542
rect 5904 5515 5989 5522
rect 6008 5539 6046 5548
rect 6008 5519 6017 5539
rect 6037 5519 6046 5539
rect 5904 5514 5940 5515
rect 6008 5511 6046 5519
rect 6112 5543 6256 5549
rect 6112 5523 6120 5543
rect 6140 5542 6228 5543
rect 6140 5523 6168 5542
rect 6112 5521 6168 5523
rect 6190 5523 6228 5542
rect 6248 5523 6256 5543
rect 6190 5521 6256 5523
rect 6112 5515 6256 5521
rect 6112 5514 6148 5515
rect 6220 5514 6256 5515
rect 6322 5548 6359 5549
rect 6322 5547 6360 5548
rect 6322 5539 6386 5547
rect 6322 5519 6331 5539
rect 6351 5525 6386 5539
rect 6406 5525 6409 5545
rect 6351 5520 6409 5525
rect 6351 5519 6386 5520
rect 5588 5482 5625 5511
rect 5056 5433 5093 5457
rect 5055 5427 5093 5433
rect 3590 5389 3840 5413
rect 4466 5409 5093 5427
rect 4048 5392 4216 5393
rect 4467 5392 4491 5409
rect 4048 5366 4492 5392
rect 4048 5364 4216 5366
rect 4048 5186 4075 5364
rect 4115 5326 4179 5338
rect 4455 5334 4492 5366
rect 4663 5365 4912 5387
rect 4663 5334 4700 5365
rect 4876 5363 4912 5365
rect 5055 5368 5093 5409
rect 5408 5436 5446 5477
rect 5589 5480 5625 5482
rect 5801 5480 5838 5511
rect 5589 5458 5838 5480
rect 6009 5479 6046 5511
rect 6322 5507 6386 5519
rect 6426 5481 6453 5659
rect 6285 5479 6453 5481
rect 6009 5453 6453 5479
rect 6010 5436 6034 5453
rect 6285 5452 6453 5453
rect 5408 5418 6035 5436
rect 6661 5432 6911 5456
rect 5408 5412 5446 5418
rect 5408 5388 5445 5412
rect 4876 5334 4913 5363
rect 4115 5325 4150 5326
rect 4092 5320 4150 5325
rect 4092 5300 4095 5320
rect 4115 5306 4150 5320
rect 4170 5306 4179 5326
rect 4115 5298 4179 5306
rect 4141 5297 4179 5298
rect 4142 5296 4179 5297
rect 4245 5330 4281 5331
rect 4353 5330 4389 5331
rect 4245 5324 4389 5330
rect 4245 5322 4311 5324
rect 4245 5302 4253 5322
rect 4273 5303 4311 5322
rect 4333 5322 4389 5324
rect 4333 5303 4361 5322
rect 4273 5302 4361 5303
rect 4381 5302 4389 5322
rect 4245 5296 4389 5302
rect 4455 5326 4493 5334
rect 4561 5330 4597 5331
rect 4455 5306 4464 5326
rect 4484 5306 4493 5326
rect 4455 5297 4493 5306
rect 4512 5323 4597 5330
rect 4512 5303 4519 5323
rect 4540 5322 4597 5323
rect 4540 5303 4569 5322
rect 4512 5302 4569 5303
rect 4589 5302 4597 5322
rect 4455 5296 4492 5297
rect 4512 5296 4597 5302
rect 4663 5326 4701 5334
rect 4774 5330 4810 5331
rect 4663 5306 4672 5326
rect 4692 5306 4701 5326
rect 4663 5297 4701 5306
rect 4725 5322 4810 5330
rect 4725 5302 4782 5322
rect 4802 5302 4810 5322
rect 4663 5296 4700 5297
rect 4725 5296 4810 5302
rect 4876 5326 4914 5334
rect 4876 5306 4885 5326
rect 4905 5306 4914 5326
rect 4876 5297 4914 5306
rect 5055 5333 5091 5368
rect 5408 5364 5443 5388
rect 5406 5355 5443 5364
rect 5406 5337 5416 5355
rect 5434 5337 5443 5355
rect 5055 5323 5092 5333
rect 5406 5327 5443 5337
rect 6661 5361 6698 5432
rect 6813 5371 6844 5372
rect 6661 5341 6670 5361
rect 6690 5341 6698 5361
rect 6661 5331 6698 5341
rect 6757 5361 6844 5371
rect 6757 5341 6766 5361
rect 6786 5341 6844 5361
rect 6757 5332 6844 5341
rect 6757 5331 6794 5332
rect 5055 5305 5065 5323
rect 5083 5305 5092 5323
rect 4876 5296 4913 5297
rect 5055 5296 5092 5305
rect 4299 5275 4335 5296
rect 4725 5275 4756 5296
rect 6813 5279 6844 5332
rect 6874 5361 6911 5432
rect 7082 5437 7475 5457
rect 7495 5437 7498 5457
rect 7082 5432 7498 5437
rect 7082 5431 7423 5432
rect 7026 5371 7057 5372
rect 6874 5341 6883 5361
rect 6903 5341 6911 5361
rect 6874 5331 6911 5341
rect 6970 5364 7057 5371
rect 6970 5361 7031 5364
rect 6970 5341 6979 5361
rect 6999 5344 7031 5361
rect 7052 5344 7057 5364
rect 6999 5341 7057 5344
rect 6970 5334 7057 5341
rect 7082 5361 7119 5431
rect 7385 5430 7422 5431
rect 7234 5371 7270 5372
rect 7082 5341 7091 5361
rect 7111 5341 7119 5361
rect 6970 5332 7026 5334
rect 6970 5331 7007 5332
rect 7082 5331 7119 5341
rect 7178 5361 7326 5371
rect 7426 5368 7522 5370
rect 7178 5341 7187 5361
rect 7207 5341 7297 5361
rect 7317 5341 7326 5361
rect 7178 5332 7326 5341
rect 7384 5361 7522 5368
rect 7384 5341 7393 5361
rect 7413 5341 7522 5361
rect 7384 5332 7522 5341
rect 7178 5331 7215 5332
rect 7234 5280 7270 5332
rect 7289 5331 7326 5332
rect 7385 5331 7422 5332
rect 6705 5278 6746 5279
rect 4132 5271 4232 5275
rect 4132 5267 4194 5271
rect 4132 5241 4139 5267
rect 4165 5245 4194 5267
rect 4220 5245 4232 5271
rect 4165 5241 4232 5245
rect 4132 5238 4232 5241
rect 4300 5238 4335 5275
rect 4397 5272 4756 5275
rect 4397 5267 4619 5272
rect 4397 5243 4410 5267
rect 4434 5248 4619 5267
rect 4643 5248 4756 5272
rect 4434 5243 4756 5248
rect 4397 5239 4756 5243
rect 4823 5267 4972 5275
rect 4823 5247 4834 5267
rect 4854 5247 4972 5267
rect 6597 5271 6746 5278
rect 5409 5263 5446 5265
rect 5409 5262 6057 5263
rect 4823 5240 4972 5247
rect 5408 5256 6057 5262
rect 4823 5239 4864 5240
rect 4147 5186 4184 5187
rect 4243 5186 4280 5187
rect 4299 5186 4335 5238
rect 4354 5186 4391 5187
rect 4047 5177 4185 5186
rect 3035 5158 3203 5159
rect 3035 5155 3479 5158
rect 3035 5136 3410 5155
rect 3430 5136 3479 5155
rect 4047 5157 4156 5177
rect 4176 5157 4185 5177
rect 3035 5132 3479 5136
rect 3035 5130 3203 5132
rect 3035 4952 3062 5130
rect 3102 5092 3166 5104
rect 3442 5100 3479 5132
rect 3650 5131 3899 5153
rect 4047 5150 4185 5157
rect 4243 5177 4391 5186
rect 4243 5157 4252 5177
rect 4272 5157 4362 5177
rect 4382 5157 4391 5177
rect 4047 5148 4143 5150
rect 4243 5147 4391 5157
rect 4450 5177 4487 5187
rect 4562 5186 4599 5187
rect 4543 5184 4599 5186
rect 4450 5157 4458 5177
rect 4478 5157 4487 5177
rect 4299 5146 4335 5147
rect 3650 5100 3687 5131
rect 3863 5129 3899 5131
rect 3863 5100 3900 5129
rect 3102 5091 3137 5092
rect 3079 5086 3137 5091
rect 3079 5066 3082 5086
rect 3102 5072 3137 5086
rect 3157 5072 3166 5092
rect 3102 5064 3166 5072
rect 3128 5063 3166 5064
rect 3129 5062 3166 5063
rect 3232 5096 3268 5097
rect 3340 5096 3376 5097
rect 3232 5088 3376 5096
rect 3232 5068 3240 5088
rect 3260 5068 3292 5088
rect 3316 5068 3348 5088
rect 3368 5068 3376 5088
rect 3232 5062 3376 5068
rect 3442 5092 3480 5100
rect 3548 5096 3584 5097
rect 3442 5072 3451 5092
rect 3471 5072 3480 5092
rect 3442 5063 3480 5072
rect 3499 5089 3584 5096
rect 3499 5069 3506 5089
rect 3527 5088 3584 5089
rect 3527 5069 3556 5088
rect 3499 5068 3556 5069
rect 3576 5068 3584 5088
rect 3442 5062 3479 5063
rect 3499 5062 3584 5068
rect 3650 5092 3688 5100
rect 3761 5096 3797 5097
rect 3650 5072 3659 5092
rect 3679 5072 3688 5092
rect 3650 5063 3688 5072
rect 3712 5088 3797 5096
rect 3712 5068 3769 5088
rect 3789 5068 3797 5088
rect 3650 5062 3687 5063
rect 3712 5062 3797 5068
rect 3863 5092 3901 5100
rect 3863 5072 3872 5092
rect 3892 5072 3901 5092
rect 4147 5087 4184 5088
rect 4450 5087 4487 5157
rect 4512 5177 4599 5184
rect 4512 5174 4570 5177
rect 4512 5154 4517 5174
rect 4538 5157 4570 5174
rect 4590 5157 4599 5177
rect 4538 5154 4599 5157
rect 4512 5147 4599 5154
rect 4658 5177 4695 5187
rect 4658 5157 4666 5177
rect 4686 5157 4695 5177
rect 4512 5146 4543 5147
rect 4146 5086 4487 5087
rect 3863 5063 3901 5072
rect 4071 5081 4487 5086
rect 3863 5062 3900 5063
rect 3286 5041 3322 5062
rect 3712 5041 3743 5062
rect 4071 5061 4074 5081
rect 4094 5061 4487 5081
rect 4658 5086 4695 5157
rect 4725 5186 4756 5239
rect 5408 5238 5418 5256
rect 5436 5242 6057 5256
rect 6597 5251 6715 5271
rect 6735 5251 6746 5271
rect 6597 5243 6746 5251
rect 6813 5275 7172 5279
rect 6813 5270 7135 5275
rect 6813 5246 6926 5270
rect 6950 5251 7135 5270
rect 7159 5251 7172 5275
rect 6950 5246 7172 5251
rect 6813 5243 7172 5246
rect 7234 5243 7269 5280
rect 7337 5277 7437 5280
rect 7337 5273 7404 5277
rect 7337 5247 7349 5273
rect 7375 5251 7404 5273
rect 7430 5251 7437 5277
rect 7375 5247 7437 5251
rect 7337 5243 7437 5247
rect 5436 5238 5446 5242
rect 5887 5241 6057 5242
rect 5058 5224 5095 5234
rect 5058 5206 5067 5224
rect 5085 5206 5095 5224
rect 5058 5197 5095 5206
rect 5408 5228 5446 5238
rect 4775 5186 4812 5187
rect 4725 5177 4812 5186
rect 4725 5157 4783 5177
rect 4803 5157 4812 5177
rect 4725 5147 4812 5157
rect 4871 5177 4908 5187
rect 4871 5157 4879 5177
rect 4899 5157 4908 5177
rect 4725 5146 4756 5147
rect 4871 5086 4908 5157
rect 5063 5132 5094 5197
rect 5408 5150 5443 5228
rect 6020 5218 6057 5241
rect 6813 5222 6844 5243
rect 7234 5222 7270 5243
rect 6656 5221 6693 5222
rect 5404 5141 5443 5150
rect 5062 5122 5099 5132
rect 5062 5120 5072 5122
rect 4996 5118 5072 5120
rect 4658 5062 4908 5086
rect 4993 5104 5072 5118
rect 5090 5104 5099 5122
rect 5404 5123 5414 5141
rect 5432 5123 5443 5141
rect 5404 5117 5443 5123
rect 5599 5193 5849 5217
rect 5599 5122 5636 5193
rect 5751 5132 5782 5133
rect 5404 5113 5441 5117
rect 4993 5101 5099 5104
rect 4465 5042 4486 5061
rect 4993 5042 5019 5101
rect 5062 5095 5099 5101
rect 5599 5102 5608 5122
rect 5628 5102 5636 5122
rect 5599 5092 5636 5102
rect 5695 5122 5782 5132
rect 5695 5102 5704 5122
rect 5724 5102 5782 5122
rect 5695 5093 5782 5102
rect 5695 5092 5732 5093
rect 5407 5042 5444 5051
rect 3119 5037 3219 5041
rect 3119 5033 3181 5037
rect 3119 5007 3126 5033
rect 3152 5011 3181 5033
rect 3207 5011 3219 5037
rect 3152 5007 3219 5011
rect 3119 5004 3219 5007
rect 3287 5004 3322 5041
rect 3384 5038 3743 5041
rect 3384 5033 3606 5038
rect 3384 5009 3397 5033
rect 3421 5014 3606 5033
rect 3630 5014 3743 5038
rect 3421 5009 3743 5014
rect 3384 5005 3743 5009
rect 3810 5033 3959 5041
rect 3810 5013 3821 5033
rect 3841 5013 3959 5033
rect 4465 5024 5019 5042
rect 5065 5031 5102 5033
rect 4993 5023 5019 5024
rect 5062 5023 5102 5031
rect 3810 5006 3959 5013
rect 5062 5011 5074 5023
rect 5053 5006 5074 5011
rect 3810 5005 3851 5006
rect 4469 5005 5074 5006
rect 5092 5005 5102 5023
rect 3134 4952 3171 4953
rect 3230 4952 3267 4953
rect 3286 4952 3322 5004
rect 3341 4952 3378 4953
rect 3034 4943 3172 4952
rect 3034 4923 3143 4943
rect 3163 4923 3172 4943
rect 3034 4916 3172 4923
rect 3230 4943 3378 4952
rect 3230 4923 3239 4943
rect 3259 4923 3349 4943
rect 3369 4923 3378 4943
rect 3034 4914 3130 4916
rect 3230 4913 3378 4923
rect 3437 4943 3474 4953
rect 3549 4952 3586 4953
rect 3530 4950 3586 4952
rect 3437 4923 3445 4943
rect 3465 4923 3474 4943
rect 3286 4912 3322 4913
rect 3134 4853 3171 4854
rect 3437 4853 3474 4923
rect 3499 4943 3586 4950
rect 3499 4940 3557 4943
rect 3499 4920 3504 4940
rect 3525 4923 3557 4940
rect 3577 4923 3586 4943
rect 3525 4920 3586 4923
rect 3499 4913 3586 4920
rect 3645 4943 3682 4953
rect 3645 4923 3653 4943
rect 3673 4923 3682 4943
rect 3499 4912 3530 4913
rect 3133 4852 3474 4853
rect 3058 4847 3474 4852
rect 3058 4827 3061 4847
rect 3081 4827 3474 4847
rect 3645 4852 3682 4923
rect 3712 4952 3743 5005
rect 4469 4996 5102 5005
rect 5405 5024 5416 5042
rect 5434 5024 5444 5042
rect 5751 5040 5782 5093
rect 5812 5122 5849 5193
rect 6020 5198 6413 5218
rect 6433 5198 6436 5218
rect 6020 5193 6436 5198
rect 6655 5212 6693 5221
rect 6020 5192 6361 5193
rect 6655 5192 6664 5212
rect 6684 5192 6693 5212
rect 5964 5132 5995 5133
rect 5812 5102 5821 5122
rect 5841 5102 5849 5122
rect 5812 5092 5849 5102
rect 5908 5125 5995 5132
rect 5908 5122 5969 5125
rect 5908 5102 5917 5122
rect 5937 5105 5969 5122
rect 5990 5105 5995 5125
rect 5937 5102 5995 5105
rect 5908 5095 5995 5102
rect 6020 5122 6057 5192
rect 6323 5191 6360 5192
rect 6655 5184 6693 5192
rect 6759 5216 6844 5222
rect 6869 5221 6906 5222
rect 6759 5196 6767 5216
rect 6787 5196 6844 5216
rect 6759 5188 6844 5196
rect 6868 5212 6906 5221
rect 6868 5192 6877 5212
rect 6897 5192 6906 5212
rect 6759 5187 6795 5188
rect 6868 5184 6906 5192
rect 6972 5216 7057 5222
rect 7077 5221 7114 5222
rect 6972 5196 6980 5216
rect 7000 5215 7057 5216
rect 7000 5196 7029 5215
rect 6972 5195 7029 5196
rect 7050 5195 7057 5215
rect 6972 5188 7057 5195
rect 7076 5212 7114 5221
rect 7076 5192 7085 5212
rect 7105 5192 7114 5212
rect 6972 5187 7008 5188
rect 7076 5184 7114 5192
rect 7180 5216 7324 5222
rect 7180 5196 7188 5216
rect 7208 5215 7296 5216
rect 7208 5196 7241 5215
rect 7264 5196 7296 5215
rect 7316 5196 7324 5216
rect 7180 5188 7324 5196
rect 7180 5187 7216 5188
rect 7288 5187 7324 5188
rect 7390 5221 7427 5222
rect 7390 5220 7428 5221
rect 7390 5212 7454 5220
rect 7390 5192 7399 5212
rect 7419 5198 7454 5212
rect 7474 5198 7477 5218
rect 7419 5193 7477 5198
rect 7419 5192 7454 5193
rect 6656 5155 6693 5184
rect 6657 5153 6693 5155
rect 6869 5153 6906 5184
rect 6172 5132 6208 5133
rect 6020 5102 6029 5122
rect 6049 5102 6057 5122
rect 5908 5093 5964 5095
rect 5908 5092 5945 5093
rect 6020 5092 6057 5102
rect 6116 5122 6264 5132
rect 6657 5131 6906 5153
rect 7077 5152 7114 5184
rect 7390 5180 7454 5192
rect 7494 5154 7521 5332
rect 7353 5152 7521 5154
rect 7077 5141 7521 5152
rect 7584 5152 7614 6153
rect 7584 5147 7616 5152
rect 6364 5129 6460 5131
rect 6116 5102 6125 5122
rect 6145 5102 6235 5122
rect 6255 5102 6264 5122
rect 6116 5093 6264 5102
rect 6322 5122 6460 5129
rect 7077 5126 7523 5141
rect 7353 5125 7523 5126
rect 6322 5102 6331 5122
rect 6351 5102 6460 5122
rect 6322 5093 6460 5102
rect 6116 5092 6153 5093
rect 6172 5041 6208 5093
rect 6227 5092 6264 5093
rect 6323 5092 6360 5093
rect 5643 5039 5684 5040
rect 4469 4989 5101 4996
rect 4469 4987 4531 4989
rect 4047 4977 4215 4978
rect 4469 4977 4491 4987
rect 3762 4952 3799 4953
rect 3712 4943 3799 4952
rect 3712 4923 3770 4943
rect 3790 4923 3799 4943
rect 3712 4913 3799 4923
rect 3858 4943 3895 4953
rect 3858 4923 3866 4943
rect 3886 4923 3895 4943
rect 3712 4912 3743 4913
rect 3858 4852 3895 4923
rect 3645 4828 3895 4852
rect 4047 4951 4491 4977
rect 4047 4949 4215 4951
rect 4047 4771 4074 4949
rect 4114 4911 4178 4923
rect 4454 4919 4491 4951
rect 4662 4950 4911 4972
rect 4662 4919 4699 4950
rect 4875 4948 4911 4950
rect 4875 4919 4912 4948
rect 4114 4910 4149 4911
rect 4091 4905 4149 4910
rect 4091 4885 4094 4905
rect 4114 4891 4149 4905
rect 4169 4891 4178 4911
rect 4114 4883 4178 4891
rect 4140 4882 4178 4883
rect 4141 4881 4178 4882
rect 4244 4915 4280 4916
rect 4352 4915 4388 4916
rect 4244 4907 4388 4915
rect 4244 4887 4252 4907
rect 4272 4887 4301 4907
rect 4244 4886 4301 4887
rect 4323 4887 4360 4907
rect 4380 4887 4388 4907
rect 4323 4886 4388 4887
rect 4244 4881 4388 4886
rect 4454 4911 4492 4919
rect 4560 4915 4596 4916
rect 4454 4891 4463 4911
rect 4483 4891 4492 4911
rect 4454 4882 4492 4891
rect 4511 4908 4596 4915
rect 4511 4888 4518 4908
rect 4539 4907 4596 4908
rect 4539 4888 4568 4907
rect 4511 4887 4568 4888
rect 4588 4887 4596 4907
rect 4454 4881 4491 4882
rect 4511 4881 4596 4887
rect 4662 4911 4700 4919
rect 4773 4915 4809 4916
rect 4662 4891 4671 4911
rect 4691 4891 4700 4911
rect 4662 4882 4700 4891
rect 4724 4907 4809 4915
rect 4724 4887 4781 4907
rect 4801 4887 4809 4907
rect 4662 4881 4699 4882
rect 4724 4881 4809 4887
rect 4875 4911 4913 4919
rect 4875 4891 4884 4911
rect 4904 4891 4913 4911
rect 4875 4882 4913 4891
rect 4875 4881 4912 4882
rect 4298 4860 4334 4881
rect 4724 4860 4755 4881
rect 4131 4856 4231 4860
rect 4131 4852 4193 4856
rect 4131 4826 4138 4852
rect 4164 4830 4193 4852
rect 4219 4830 4231 4856
rect 4164 4826 4231 4830
rect 4131 4823 4231 4826
rect 4299 4823 4334 4860
rect 4396 4857 4755 4860
rect 4396 4852 4618 4857
rect 4396 4828 4409 4852
rect 4433 4833 4618 4852
rect 4642 4833 4755 4857
rect 4433 4828 4755 4833
rect 4396 4824 4755 4828
rect 4822 4852 4971 4860
rect 4822 4832 4833 4852
rect 4853 4832 4971 4852
rect 4822 4825 4971 4832
rect 5062 4840 5101 4989
rect 5405 4875 5444 5024
rect 5535 5032 5684 5039
rect 5535 5012 5653 5032
rect 5673 5012 5684 5032
rect 5535 5004 5684 5012
rect 5751 5036 6110 5040
rect 5751 5031 6073 5036
rect 5751 5007 5864 5031
rect 5888 5012 6073 5031
rect 6097 5012 6110 5036
rect 5888 5007 6110 5012
rect 5751 5004 6110 5007
rect 6172 5004 6207 5041
rect 6275 5038 6375 5041
rect 6275 5034 6342 5038
rect 6275 5008 6287 5034
rect 6313 5012 6342 5034
rect 6368 5012 6375 5038
rect 6313 5008 6375 5012
rect 6275 5004 6375 5008
rect 5751 4983 5782 5004
rect 6172 4983 6208 5004
rect 5594 4982 5631 4983
rect 5593 4973 5631 4982
rect 5593 4953 5602 4973
rect 5622 4953 5631 4973
rect 5593 4945 5631 4953
rect 5697 4977 5782 4983
rect 5807 4982 5844 4983
rect 5697 4957 5705 4977
rect 5725 4957 5782 4977
rect 5697 4949 5782 4957
rect 5806 4973 5844 4982
rect 5806 4953 5815 4973
rect 5835 4953 5844 4973
rect 5697 4948 5733 4949
rect 5806 4945 5844 4953
rect 5910 4977 5995 4983
rect 6015 4982 6052 4983
rect 5910 4957 5918 4977
rect 5938 4976 5995 4977
rect 5938 4957 5967 4976
rect 5910 4956 5967 4957
rect 5988 4956 5995 4976
rect 5910 4949 5995 4956
rect 6014 4973 6052 4982
rect 6014 4953 6023 4973
rect 6043 4953 6052 4973
rect 5910 4948 5946 4949
rect 6014 4945 6052 4953
rect 6118 4978 6262 4983
rect 6118 4977 6183 4978
rect 6118 4957 6126 4977
rect 6146 4957 6183 4977
rect 6205 4977 6262 4978
rect 6205 4957 6234 4977
rect 6254 4957 6262 4977
rect 6118 4949 6262 4957
rect 6118 4948 6154 4949
rect 6226 4948 6262 4949
rect 6328 4982 6365 4983
rect 6328 4981 6366 4982
rect 6328 4973 6392 4981
rect 6328 4953 6337 4973
rect 6357 4959 6392 4973
rect 6412 4959 6415 4979
rect 6357 4954 6415 4959
rect 6357 4953 6392 4954
rect 5594 4916 5631 4945
rect 5595 4914 5631 4916
rect 5807 4914 5844 4945
rect 5595 4892 5844 4914
rect 6015 4913 6052 4945
rect 6328 4941 6392 4953
rect 6432 4915 6459 5093
rect 6291 4913 6459 4915
rect 6015 4887 6459 4913
rect 6611 5012 6861 5036
rect 6611 4941 6648 5012
rect 6763 4951 6794 4952
rect 6611 4921 6620 4941
rect 6640 4921 6648 4941
rect 6611 4911 6648 4921
rect 6707 4941 6794 4951
rect 6707 4921 6716 4941
rect 6736 4921 6794 4941
rect 6707 4912 6794 4921
rect 6707 4911 6744 4912
rect 6015 4877 6037 4887
rect 6291 4886 6459 4887
rect 5975 4875 6037 4877
rect 5405 4868 6037 4875
rect 4822 4824 4863 4825
rect 4146 4771 4183 4772
rect 4242 4771 4279 4772
rect 4298 4771 4334 4823
rect 4353 4771 4390 4772
rect 4046 4762 4184 4771
rect 4046 4742 4155 4762
rect 4175 4742 4184 4762
rect 4046 4735 4184 4742
rect 4242 4762 4390 4771
rect 4242 4742 4251 4762
rect 4271 4742 4361 4762
rect 4381 4742 4390 4762
rect 4046 4733 4142 4735
rect 4242 4732 4390 4742
rect 4449 4762 4486 4772
rect 4561 4771 4598 4772
rect 4542 4769 4598 4771
rect 4449 4742 4457 4762
rect 4477 4742 4486 4762
rect 4298 4731 4334 4732
rect 2211 4723 2242 4726
rect 2740 4726 2908 4727
rect 1040 4699 1178 4708
rect 2740 4700 3184 4726
rect 834 4698 871 4699
rect 890 4647 926 4699
rect 945 4698 982 4699
rect 1041 4698 1078 4699
rect 361 4645 402 4646
rect 253 4638 402 4645
rect 253 4618 371 4638
rect 391 4618 402 4638
rect 253 4610 402 4618
rect 469 4642 828 4646
rect 469 4637 791 4642
rect 469 4613 582 4637
rect 606 4618 791 4637
rect 815 4618 828 4642
rect 606 4613 828 4618
rect 469 4610 828 4613
rect 890 4610 925 4647
rect 993 4644 1093 4647
rect 993 4640 1060 4644
rect 993 4614 1005 4640
rect 1031 4618 1060 4640
rect 1086 4618 1093 4644
rect 1031 4614 1093 4618
rect 993 4610 1093 4614
rect 469 4589 500 4610
rect 890 4589 926 4610
rect 133 4580 170 4589
rect 312 4588 349 4589
rect 133 4562 142 4580
rect 160 4562 170 4580
rect 133 4552 170 4562
rect 134 4517 170 4552
rect 311 4579 349 4588
rect 311 4559 320 4579
rect 340 4559 349 4579
rect 311 4551 349 4559
rect 415 4583 500 4589
rect 525 4588 562 4589
rect 415 4563 423 4583
rect 443 4563 500 4583
rect 415 4555 500 4563
rect 524 4579 562 4588
rect 524 4559 533 4579
rect 553 4559 562 4579
rect 415 4554 451 4555
rect 524 4551 562 4559
rect 628 4583 713 4589
rect 733 4588 770 4589
rect 628 4563 636 4583
rect 656 4582 713 4583
rect 656 4563 685 4582
rect 628 4562 685 4563
rect 706 4562 713 4582
rect 628 4555 713 4562
rect 732 4579 770 4588
rect 732 4559 741 4579
rect 761 4559 770 4579
rect 628 4554 664 4555
rect 732 4551 770 4559
rect 836 4583 980 4589
rect 836 4563 844 4583
rect 864 4582 952 4583
rect 864 4563 892 4582
rect 836 4561 892 4563
rect 914 4563 952 4582
rect 972 4563 980 4583
rect 914 4561 980 4563
rect 836 4555 980 4561
rect 836 4554 872 4555
rect 944 4554 980 4555
rect 1046 4588 1083 4589
rect 1046 4587 1084 4588
rect 1046 4579 1110 4587
rect 1046 4559 1055 4579
rect 1075 4565 1110 4579
rect 1130 4565 1133 4585
rect 1075 4560 1133 4565
rect 1075 4559 1110 4560
rect 312 4522 349 4551
rect 132 4476 170 4517
rect 313 4520 349 4522
rect 525 4520 562 4551
rect 313 4498 562 4520
rect 733 4519 770 4551
rect 1046 4547 1110 4559
rect 1150 4521 1177 4699
rect 1009 4519 1177 4521
rect 2740 4698 2908 4700
rect 2740 4695 2787 4698
rect 2740 4520 2767 4695
rect 2807 4660 2871 4672
rect 3147 4668 3184 4700
rect 3355 4699 3604 4721
rect 3355 4668 3392 4699
rect 3568 4697 3604 4699
rect 3568 4668 3605 4697
rect 4146 4672 4183 4673
rect 4449 4672 4486 4742
rect 4511 4762 4598 4769
rect 4511 4759 4569 4762
rect 4511 4739 4516 4759
rect 4537 4742 4569 4759
rect 4589 4742 4598 4762
rect 4537 4739 4598 4742
rect 4511 4732 4598 4739
rect 4657 4762 4694 4772
rect 4657 4742 4665 4762
rect 4685 4742 4694 4762
rect 4511 4731 4542 4732
rect 4145 4671 4486 4672
rect 2807 4659 2842 4660
rect 2784 4654 2842 4659
rect 2784 4634 2787 4654
rect 2807 4640 2842 4654
rect 2862 4640 2871 4660
rect 2807 4632 2871 4640
rect 2833 4631 2871 4632
rect 2834 4630 2871 4631
rect 2937 4664 2973 4665
rect 3045 4664 3081 4665
rect 2937 4656 3081 4664
rect 2937 4636 2945 4656
rect 2965 4654 3053 4656
rect 2965 4636 2991 4654
rect 2937 4635 2991 4636
rect 3017 4636 3053 4654
rect 3073 4636 3081 4656
rect 3017 4635 3081 4636
rect 2937 4630 3081 4635
rect 3147 4660 3185 4668
rect 3253 4664 3289 4665
rect 3147 4640 3156 4660
rect 3176 4640 3185 4660
rect 3147 4631 3185 4640
rect 3204 4657 3289 4664
rect 3204 4637 3211 4657
rect 3232 4656 3289 4657
rect 3232 4637 3261 4656
rect 3204 4636 3261 4637
rect 3281 4636 3289 4656
rect 3147 4630 3184 4631
rect 3204 4630 3289 4636
rect 3355 4660 3393 4668
rect 3466 4664 3502 4665
rect 3355 4640 3364 4660
rect 3384 4640 3393 4660
rect 3355 4631 3393 4640
rect 3417 4656 3502 4664
rect 3417 4636 3474 4656
rect 3494 4636 3502 4656
rect 3355 4630 3392 4631
rect 3417 4630 3502 4636
rect 3568 4660 3606 4668
rect 3568 4640 3577 4660
rect 3597 4640 3606 4660
rect 4070 4666 4486 4671
rect 4070 4646 4073 4666
rect 4093 4646 4486 4666
rect 4657 4671 4694 4742
rect 4724 4771 4755 4824
rect 5062 4822 5072 4840
rect 5090 4822 5101 4840
rect 5404 4859 6037 4868
rect 6763 4859 6794 4912
rect 6824 4941 6861 5012
rect 7032 5017 7425 5037
rect 7445 5017 7448 5037
rect 7032 5012 7448 5017
rect 7032 5011 7373 5012
rect 6976 4951 7007 4952
rect 6824 4921 6833 4941
rect 6853 4921 6861 4941
rect 6824 4911 6861 4921
rect 6920 4944 7007 4951
rect 6920 4941 6981 4944
rect 6920 4921 6929 4941
rect 6949 4924 6981 4941
rect 7002 4924 7007 4944
rect 6949 4921 7007 4924
rect 6920 4914 7007 4921
rect 7032 4941 7069 5011
rect 7335 5010 7372 5011
rect 7184 4951 7220 4952
rect 7032 4921 7041 4941
rect 7061 4921 7069 4941
rect 6920 4912 6976 4914
rect 6920 4911 6957 4912
rect 7032 4911 7069 4921
rect 7128 4941 7276 4951
rect 7376 4948 7472 4950
rect 7128 4921 7137 4941
rect 7157 4921 7247 4941
rect 7267 4921 7276 4941
rect 7128 4912 7276 4921
rect 7334 4941 7472 4948
rect 7334 4921 7343 4941
rect 7363 4921 7472 4941
rect 7334 4912 7472 4921
rect 7128 4911 7165 4912
rect 7184 4860 7220 4912
rect 7239 4911 7276 4912
rect 7335 4911 7372 4912
rect 5404 4841 5414 4859
rect 5432 4858 6037 4859
rect 6655 4858 6696 4859
rect 5432 4853 5453 4858
rect 5432 4841 5444 4853
rect 6547 4851 6696 4858
rect 5404 4833 5444 4841
rect 5487 4840 5513 4841
rect 5404 4831 5441 4833
rect 5487 4822 6041 4840
rect 6547 4831 6665 4851
rect 6685 4831 6696 4851
rect 6547 4823 6696 4831
rect 6763 4855 7122 4859
rect 6763 4850 7085 4855
rect 6763 4826 6876 4850
rect 6900 4831 7085 4850
rect 7109 4831 7122 4855
rect 6900 4826 7122 4831
rect 6763 4823 7122 4826
rect 7184 4823 7219 4860
rect 7287 4857 7387 4860
rect 7287 4853 7354 4857
rect 7287 4827 7299 4853
rect 7325 4831 7354 4853
rect 7380 4831 7387 4857
rect 7325 4827 7387 4831
rect 7287 4823 7387 4827
rect 5062 4813 5099 4822
rect 4774 4771 4811 4772
rect 4724 4762 4811 4771
rect 4724 4742 4782 4762
rect 4802 4742 4811 4762
rect 4724 4732 4811 4742
rect 4870 4762 4907 4772
rect 4870 4742 4878 4762
rect 4898 4742 4907 4762
rect 5407 4763 5444 4769
rect 5487 4763 5513 4822
rect 6020 4803 6041 4822
rect 5407 4760 5513 4763
rect 5065 4747 5102 4751
rect 4724 4731 4755 4732
rect 4870 4671 4907 4742
rect 4657 4647 4907 4671
rect 5063 4741 5102 4747
rect 5063 4723 5074 4741
rect 5092 4723 5102 4741
rect 5407 4742 5416 4760
rect 5434 4746 5513 4760
rect 5598 4778 5848 4802
rect 5434 4744 5510 4746
rect 5434 4742 5444 4744
rect 5407 4732 5444 4742
rect 5063 4714 5102 4723
rect 3568 4631 3606 4640
rect 3568 4630 3605 4631
rect 2991 4609 3027 4630
rect 3417 4609 3448 4630
rect 4449 4623 4486 4646
rect 5063 4636 5098 4714
rect 5412 4667 5443 4732
rect 5598 4707 5635 4778
rect 5750 4717 5781 4718
rect 5598 4687 5607 4707
rect 5627 4687 5635 4707
rect 5598 4677 5635 4687
rect 5694 4707 5781 4717
rect 5694 4687 5703 4707
rect 5723 4687 5781 4707
rect 5694 4678 5781 4687
rect 5694 4677 5731 4678
rect 5060 4626 5098 4636
rect 5411 4658 5448 4667
rect 5411 4640 5421 4658
rect 5439 4640 5448 4658
rect 5411 4630 5448 4640
rect 4449 4622 4619 4623
rect 5060 4622 5070 4626
rect 2824 4605 2924 4609
rect 2824 4601 2886 4605
rect 2824 4575 2831 4601
rect 2857 4579 2886 4601
rect 2912 4579 2924 4605
rect 2857 4575 2924 4579
rect 2824 4572 2924 4575
rect 2992 4572 3027 4609
rect 3089 4606 3448 4609
rect 3089 4601 3311 4606
rect 3089 4577 3102 4601
rect 3126 4582 3311 4601
rect 3335 4582 3448 4606
rect 3126 4577 3448 4582
rect 3089 4573 3448 4577
rect 3515 4601 3664 4609
rect 4449 4608 5070 4622
rect 5088 4608 5098 4626
rect 5750 4625 5781 4678
rect 5811 4707 5848 4778
rect 6019 4783 6412 4803
rect 6432 4783 6435 4803
rect 6763 4802 6794 4823
rect 7184 4802 7220 4823
rect 6606 4801 6643 4802
rect 6019 4778 6435 4783
rect 6605 4792 6643 4801
rect 6019 4777 6360 4778
rect 5963 4717 5994 4718
rect 5811 4687 5820 4707
rect 5840 4687 5848 4707
rect 5811 4677 5848 4687
rect 5907 4710 5994 4717
rect 5907 4707 5968 4710
rect 5907 4687 5916 4707
rect 5936 4690 5968 4707
rect 5989 4690 5994 4710
rect 5936 4687 5994 4690
rect 5907 4680 5994 4687
rect 6019 4707 6056 4777
rect 6322 4776 6359 4777
rect 6605 4772 6614 4792
rect 6634 4772 6643 4792
rect 6605 4764 6643 4772
rect 6709 4796 6794 4802
rect 6819 4801 6856 4802
rect 6709 4776 6717 4796
rect 6737 4776 6794 4796
rect 6709 4768 6794 4776
rect 6818 4792 6856 4801
rect 6818 4772 6827 4792
rect 6847 4772 6856 4792
rect 6709 4767 6745 4768
rect 6818 4764 6856 4772
rect 6922 4796 7007 4802
rect 7027 4801 7064 4802
rect 6922 4776 6930 4796
rect 6950 4795 7007 4796
rect 6950 4776 6979 4795
rect 6922 4775 6979 4776
rect 7000 4775 7007 4795
rect 6922 4768 7007 4775
rect 7026 4792 7064 4801
rect 7026 4772 7035 4792
rect 7055 4772 7064 4792
rect 6922 4767 6958 4768
rect 7026 4764 7064 4772
rect 7130 4797 7274 4802
rect 7130 4796 7189 4797
rect 7130 4776 7138 4796
rect 7158 4777 7189 4796
rect 7213 4796 7274 4797
rect 7213 4777 7246 4796
rect 7158 4776 7246 4777
rect 7266 4776 7274 4796
rect 7130 4768 7274 4776
rect 7130 4767 7166 4768
rect 7238 4767 7274 4768
rect 7340 4801 7377 4802
rect 7340 4800 7378 4801
rect 7340 4792 7404 4800
rect 7340 4772 7349 4792
rect 7369 4778 7404 4792
rect 7424 4778 7427 4798
rect 7369 4773 7427 4778
rect 7369 4772 7404 4773
rect 6606 4735 6643 4764
rect 6607 4733 6643 4735
rect 6819 4733 6856 4764
rect 6171 4717 6207 4718
rect 6019 4687 6028 4707
rect 6048 4687 6056 4707
rect 5907 4678 5963 4680
rect 5907 4677 5944 4678
rect 6019 4677 6056 4687
rect 6115 4707 6263 4717
rect 6363 4714 6459 4716
rect 6115 4687 6124 4707
rect 6144 4687 6234 4707
rect 6254 4687 6263 4707
rect 6115 4678 6263 4687
rect 6321 4707 6459 4714
rect 6607 4711 6856 4733
rect 7027 4732 7064 4764
rect 7340 4760 7404 4772
rect 7444 4734 7471 4912
rect 7303 4732 7471 4734
rect 7027 4728 7471 4732
rect 6321 4687 6330 4707
rect 6350 4687 6459 4707
rect 7027 4709 7076 4728
rect 7096 4709 7471 4728
rect 7027 4706 7471 4709
rect 7303 4705 7471 4706
rect 7492 4731 7523 5125
rect 7584 5129 7589 5147
rect 7609 5129 7616 5147
rect 7584 5124 7616 5129
rect 7587 5122 7616 5124
rect 7492 4705 7497 4731
rect 7516 4705 7523 4731
rect 8030 4706 8068 6537
rect 8096 6424 8123 6602
rect 8163 6564 8227 6576
rect 8503 6572 8540 6604
rect 8711 6603 8960 6625
rect 9415 6611 9452 6612
rect 9718 6611 9755 6681
rect 9780 6701 9867 6708
rect 9780 6698 9838 6701
rect 9780 6678 9785 6698
rect 9806 6681 9838 6698
rect 9858 6681 9867 6701
rect 9806 6678 9867 6681
rect 9780 6671 9867 6678
rect 9926 6701 9963 6711
rect 9926 6681 9934 6701
rect 9954 6681 9963 6701
rect 9780 6670 9811 6671
rect 9414 6610 9755 6611
rect 8711 6572 8748 6603
rect 8924 6601 8960 6603
rect 9339 6605 9755 6610
rect 8924 6572 8961 6601
rect 9339 6585 9342 6605
rect 9362 6585 9755 6605
rect 9926 6610 9963 6681
rect 9993 6710 10024 6763
rect 10331 6761 10341 6779
rect 10359 6761 10370 6779
rect 10855 6811 11409 6829
rect 11915 6820 12033 6840
rect 12053 6820 12064 6840
rect 11915 6812 12064 6820
rect 12131 6844 12490 6848
rect 12131 6839 12453 6844
rect 12131 6815 12244 6839
rect 12268 6820 12453 6839
rect 12477 6820 12490 6844
rect 12268 6815 12490 6820
rect 12131 6812 12490 6815
rect 12552 6812 12587 6849
rect 12655 6846 12755 6849
rect 12655 6842 12722 6846
rect 12655 6816 12667 6842
rect 12693 6820 12722 6842
rect 12748 6820 12755 6846
rect 12693 6816 12755 6820
rect 12655 6812 12755 6816
rect 10331 6752 10368 6761
rect 10775 6752 10812 6758
rect 10855 6752 10881 6811
rect 11388 6792 11409 6811
rect 10775 6749 10881 6752
rect 10775 6731 10784 6749
rect 10802 6735 10881 6749
rect 10966 6767 11216 6791
rect 10802 6733 10878 6735
rect 10802 6731 10812 6733
rect 10775 6721 10812 6731
rect 10043 6710 10080 6711
rect 9993 6701 10080 6710
rect 9993 6681 10051 6701
rect 10071 6681 10080 6701
rect 9993 6671 10080 6681
rect 10139 6701 10176 6711
rect 10139 6681 10147 6701
rect 10167 6681 10176 6701
rect 10334 6686 10371 6690
rect 9993 6670 10024 6671
rect 10139 6610 10176 6681
rect 9926 6586 10176 6610
rect 10332 6680 10371 6686
rect 10332 6662 10343 6680
rect 10361 6662 10371 6680
rect 10332 6653 10371 6662
rect 10780 6656 10811 6721
rect 10966 6696 11003 6767
rect 11118 6706 11149 6707
rect 10966 6676 10975 6696
rect 10995 6676 11003 6696
rect 10966 6666 11003 6676
rect 11062 6696 11149 6706
rect 11062 6676 11071 6696
rect 11091 6676 11149 6696
rect 11062 6667 11149 6676
rect 11062 6666 11099 6667
rect 8163 6563 8198 6564
rect 8140 6558 8198 6563
rect 8140 6538 8143 6558
rect 8163 6544 8198 6558
rect 8218 6544 8227 6564
rect 8163 6536 8227 6544
rect 8189 6535 8227 6536
rect 8190 6534 8227 6535
rect 8293 6568 8329 6569
rect 8401 6568 8437 6569
rect 8293 6560 8437 6568
rect 8293 6540 8301 6560
rect 8321 6559 8409 6560
rect 8321 6540 8350 6559
rect 8373 6540 8409 6559
rect 8429 6540 8437 6560
rect 8293 6534 8437 6540
rect 8503 6564 8541 6572
rect 8609 6568 8645 6569
rect 8503 6544 8512 6564
rect 8532 6544 8541 6564
rect 8503 6535 8541 6544
rect 8560 6561 8645 6568
rect 8560 6541 8567 6561
rect 8588 6560 8645 6561
rect 8588 6541 8617 6560
rect 8560 6540 8617 6541
rect 8637 6540 8645 6560
rect 8503 6534 8540 6535
rect 8560 6534 8645 6540
rect 8711 6564 8749 6572
rect 8822 6568 8858 6569
rect 8711 6544 8720 6564
rect 8740 6544 8749 6564
rect 8711 6535 8749 6544
rect 8773 6560 8858 6568
rect 8773 6540 8830 6560
rect 8850 6540 8858 6560
rect 8711 6534 8748 6535
rect 8773 6534 8858 6540
rect 8924 6564 8962 6572
rect 8924 6544 8933 6564
rect 8953 6544 8962 6564
rect 8924 6535 8962 6544
rect 9718 6562 9755 6585
rect 10332 6575 10367 6653
rect 10779 6647 10816 6656
rect 10779 6629 10789 6647
rect 10807 6629 10816 6647
rect 10779 6619 10816 6629
rect 11118 6614 11149 6667
rect 11179 6696 11216 6767
rect 11387 6772 11780 6792
rect 11800 6772 11803 6792
rect 12131 6791 12162 6812
rect 12552 6791 12588 6812
rect 11974 6790 12011 6791
rect 11387 6767 11803 6772
rect 11973 6781 12011 6790
rect 11387 6766 11728 6767
rect 11331 6706 11362 6707
rect 11179 6676 11188 6696
rect 11208 6676 11216 6696
rect 11179 6666 11216 6676
rect 11275 6699 11362 6706
rect 11275 6696 11336 6699
rect 11275 6676 11284 6696
rect 11304 6679 11336 6696
rect 11357 6679 11362 6699
rect 11304 6676 11362 6679
rect 11275 6669 11362 6676
rect 11387 6696 11424 6766
rect 11690 6765 11727 6766
rect 11973 6761 11982 6781
rect 12002 6761 12011 6781
rect 11973 6753 12011 6761
rect 12077 6785 12162 6791
rect 12187 6790 12224 6791
rect 12077 6765 12085 6785
rect 12105 6765 12162 6785
rect 12077 6757 12162 6765
rect 12186 6781 12224 6790
rect 12186 6761 12195 6781
rect 12215 6761 12224 6781
rect 12077 6756 12113 6757
rect 12186 6753 12224 6761
rect 12290 6785 12375 6791
rect 12395 6790 12432 6791
rect 12290 6765 12298 6785
rect 12318 6784 12375 6785
rect 12318 6765 12347 6784
rect 12290 6764 12347 6765
rect 12368 6764 12375 6784
rect 12290 6757 12375 6764
rect 12394 6781 12432 6790
rect 12394 6761 12403 6781
rect 12423 6761 12432 6781
rect 12290 6756 12326 6757
rect 12394 6753 12432 6761
rect 12498 6786 12642 6791
rect 12498 6785 12557 6786
rect 12498 6765 12506 6785
rect 12526 6766 12557 6785
rect 12581 6785 12642 6786
rect 12581 6766 12614 6785
rect 12526 6765 12614 6766
rect 12634 6765 12642 6785
rect 12498 6757 12642 6765
rect 12498 6756 12534 6757
rect 12606 6756 12642 6757
rect 12708 6790 12745 6791
rect 12708 6789 12746 6790
rect 12708 6781 12772 6789
rect 12708 6761 12717 6781
rect 12737 6767 12772 6781
rect 12792 6767 12795 6787
rect 12737 6762 12795 6767
rect 12737 6761 12772 6762
rect 11974 6724 12011 6753
rect 11975 6722 12011 6724
rect 12187 6722 12224 6753
rect 11539 6706 11575 6707
rect 11387 6676 11396 6696
rect 11416 6676 11424 6696
rect 11275 6667 11331 6669
rect 11275 6666 11312 6667
rect 11387 6666 11424 6676
rect 11483 6696 11631 6706
rect 11731 6703 11827 6705
rect 11483 6676 11492 6696
rect 11512 6676 11602 6696
rect 11622 6676 11631 6696
rect 11483 6667 11631 6676
rect 11689 6696 11827 6703
rect 11975 6700 12224 6722
rect 12395 6721 12432 6753
rect 12708 6749 12772 6761
rect 12812 6723 12839 6901
rect 12671 6721 12839 6723
rect 12395 6717 12839 6721
rect 11689 6676 11698 6696
rect 11718 6676 11827 6696
rect 12395 6698 12444 6717
rect 12464 6698 12839 6717
rect 12395 6695 12839 6698
rect 12671 6694 12839 6695
rect 12860 6720 12891 7114
rect 12860 6694 12865 6720
rect 12884 6694 12891 6720
rect 12860 6691 12891 6694
rect 11689 6667 11827 6676
rect 11483 6666 11520 6667
rect 11539 6615 11575 6667
rect 11594 6666 11631 6667
rect 11690 6666 11727 6667
rect 11010 6613 11051 6614
rect 10902 6606 11051 6613
rect 10902 6586 11020 6606
rect 11040 6586 11051 6606
rect 10902 6578 11051 6586
rect 11118 6610 11477 6614
rect 11118 6605 11440 6610
rect 11118 6581 11231 6605
rect 11255 6586 11440 6605
rect 11464 6586 11477 6610
rect 11255 6581 11477 6586
rect 11118 6578 11477 6581
rect 11539 6578 11574 6615
rect 11642 6612 11742 6615
rect 11642 6608 11709 6612
rect 11642 6582 11654 6608
rect 11680 6586 11709 6608
rect 11735 6586 11742 6612
rect 11680 6582 11742 6586
rect 11642 6578 11742 6582
rect 10329 6565 10367 6575
rect 9718 6561 9888 6562
rect 10329 6561 10339 6565
rect 9718 6547 10339 6561
rect 10357 6547 10367 6565
rect 11118 6557 11149 6578
rect 11539 6557 11575 6578
rect 9718 6541 10367 6547
rect 10782 6548 10819 6557
rect 10961 6556 10998 6557
rect 9718 6540 10366 6541
rect 10329 6538 10366 6540
rect 8924 6534 8961 6535
rect 8347 6513 8383 6534
rect 8773 6513 8804 6534
rect 10782 6530 10791 6548
rect 10809 6530 10819 6548
rect 10782 6520 10819 6530
rect 8180 6509 8280 6513
rect 8180 6505 8242 6509
rect 8180 6479 8187 6505
rect 8213 6483 8242 6505
rect 8268 6483 8280 6509
rect 8213 6479 8280 6483
rect 8180 6476 8280 6479
rect 8348 6476 8383 6513
rect 8445 6510 8804 6513
rect 8445 6505 8667 6510
rect 8445 6481 8458 6505
rect 8482 6486 8667 6505
rect 8691 6486 8804 6510
rect 8482 6481 8804 6486
rect 8445 6477 8804 6481
rect 8871 6505 9020 6513
rect 8871 6485 8882 6505
rect 8902 6485 9020 6505
rect 10783 6485 10819 6520
rect 10960 6547 10998 6556
rect 10960 6527 10969 6547
rect 10989 6527 10998 6547
rect 10960 6519 10998 6527
rect 11064 6551 11149 6557
rect 11174 6556 11211 6557
rect 11064 6531 11072 6551
rect 11092 6531 11149 6551
rect 11064 6523 11149 6531
rect 11173 6547 11211 6556
rect 11173 6527 11182 6547
rect 11202 6527 11211 6547
rect 11064 6522 11100 6523
rect 11173 6519 11211 6527
rect 11277 6551 11362 6557
rect 11382 6556 11419 6557
rect 11277 6531 11285 6551
rect 11305 6550 11362 6551
rect 11305 6531 11334 6550
rect 11277 6530 11334 6531
rect 11355 6530 11362 6550
rect 11277 6523 11362 6530
rect 11381 6547 11419 6556
rect 11381 6527 11390 6547
rect 11410 6527 11419 6547
rect 11277 6522 11313 6523
rect 11381 6519 11419 6527
rect 11485 6551 11629 6557
rect 11485 6531 11493 6551
rect 11513 6550 11601 6551
rect 11513 6531 11541 6550
rect 11485 6529 11541 6531
rect 11563 6531 11601 6550
rect 11621 6531 11629 6551
rect 11563 6529 11629 6531
rect 11485 6523 11629 6529
rect 11485 6522 11521 6523
rect 11593 6522 11629 6523
rect 11695 6556 11732 6557
rect 11695 6555 11733 6556
rect 11695 6547 11759 6555
rect 11695 6527 11704 6547
rect 11724 6533 11759 6547
rect 11779 6533 11782 6553
rect 11724 6528 11782 6533
rect 11724 6527 11759 6528
rect 10961 6490 10998 6519
rect 8871 6478 9020 6485
rect 8871 6477 8912 6478
rect 8195 6424 8232 6425
rect 8291 6424 8328 6425
rect 8347 6424 8383 6476
rect 8402 6424 8439 6425
rect 8095 6415 8233 6424
rect 8095 6395 8204 6415
rect 8224 6395 8233 6415
rect 8095 6388 8233 6395
rect 8291 6415 8439 6424
rect 8291 6395 8300 6415
rect 8320 6395 8410 6415
rect 8430 6395 8439 6415
rect 8095 6386 8191 6388
rect 8291 6385 8439 6395
rect 8498 6415 8535 6425
rect 8610 6424 8647 6425
rect 8591 6422 8647 6424
rect 8498 6395 8506 6415
rect 8526 6395 8535 6415
rect 8347 6384 8383 6385
rect 8195 6325 8232 6326
rect 8498 6325 8535 6395
rect 8560 6415 8647 6422
rect 8560 6412 8618 6415
rect 8560 6392 8565 6412
rect 8586 6395 8618 6412
rect 8638 6395 8647 6415
rect 8586 6392 8647 6395
rect 8560 6385 8647 6392
rect 8706 6415 8743 6425
rect 8706 6395 8714 6415
rect 8734 6395 8743 6415
rect 8560 6384 8591 6385
rect 8194 6324 8535 6325
rect 8119 6319 8535 6324
rect 8119 6299 8122 6319
rect 8142 6299 8535 6319
rect 8706 6324 8743 6395
rect 8773 6424 8804 6477
rect 10332 6466 10369 6476
rect 10332 6448 10341 6466
rect 10359 6448 10369 6466
rect 10332 6439 10369 6448
rect 10781 6444 10819 6485
rect 10962 6488 10998 6490
rect 11174 6488 11211 6519
rect 10962 6466 11211 6488
rect 11382 6487 11419 6519
rect 11695 6515 11759 6527
rect 11799 6489 11826 6667
rect 13410 6656 13447 6667
rect 13536 6660 13566 7661
rect 13629 7661 14073 7672
rect 13629 7659 13797 7661
rect 13629 7481 13656 7659
rect 13696 7621 13760 7633
rect 14036 7629 14073 7661
rect 14244 7660 14493 7682
rect 14886 7681 15034 7691
rect 15093 7711 15130 7721
rect 15205 7720 15242 7721
rect 15186 7718 15242 7720
rect 15093 7691 15101 7711
rect 15121 7691 15130 7711
rect 14942 7680 14978 7681
rect 14244 7629 14281 7660
rect 14457 7658 14493 7660
rect 14457 7629 14494 7658
rect 13696 7620 13731 7621
rect 13673 7615 13731 7620
rect 13673 7595 13676 7615
rect 13696 7601 13731 7615
rect 13751 7601 13760 7621
rect 13696 7593 13760 7601
rect 13722 7592 13760 7593
rect 13723 7591 13760 7592
rect 13826 7625 13862 7626
rect 13934 7625 13970 7626
rect 13826 7617 13970 7625
rect 13826 7597 13834 7617
rect 13854 7598 13886 7617
rect 13909 7598 13942 7617
rect 13854 7597 13942 7598
rect 13962 7597 13970 7617
rect 13826 7591 13970 7597
rect 14036 7621 14074 7629
rect 14142 7625 14178 7626
rect 14036 7601 14045 7621
rect 14065 7601 14074 7621
rect 14036 7592 14074 7601
rect 14093 7618 14178 7625
rect 14093 7598 14100 7618
rect 14121 7617 14178 7618
rect 14121 7598 14150 7617
rect 14093 7597 14150 7598
rect 14170 7597 14178 7617
rect 14036 7591 14073 7592
rect 14093 7591 14178 7597
rect 14244 7621 14282 7629
rect 14355 7625 14391 7626
rect 14244 7601 14253 7621
rect 14273 7601 14282 7621
rect 14244 7592 14282 7601
rect 14306 7617 14391 7625
rect 14306 7597 14363 7617
rect 14383 7597 14391 7617
rect 14244 7591 14281 7592
rect 14306 7591 14391 7597
rect 14457 7621 14495 7629
rect 14790 7621 14827 7622
rect 15093 7621 15130 7691
rect 15155 7711 15242 7718
rect 15155 7708 15213 7711
rect 15155 7688 15160 7708
rect 15181 7691 15213 7708
rect 15233 7691 15242 7711
rect 15181 7688 15242 7691
rect 15155 7681 15242 7688
rect 15301 7711 15338 7721
rect 15301 7691 15309 7711
rect 15329 7691 15338 7711
rect 15155 7680 15186 7681
rect 14457 7601 14466 7621
rect 14486 7601 14495 7621
rect 14789 7620 15130 7621
rect 14457 7592 14495 7601
rect 14714 7615 15130 7620
rect 14714 7595 14717 7615
rect 14737 7595 15130 7615
rect 15301 7620 15338 7691
rect 15368 7720 15399 7773
rect 15706 7771 15716 7789
rect 15734 7771 15745 7789
rect 16048 7808 16681 7817
rect 17407 7808 17438 7861
rect 17468 7890 17505 7961
rect 17676 7966 18069 7986
rect 18089 7966 18092 7986
rect 17676 7961 18092 7966
rect 17676 7960 18017 7961
rect 17620 7900 17651 7901
rect 17468 7870 17477 7890
rect 17497 7870 17505 7890
rect 17468 7860 17505 7870
rect 17564 7893 17651 7900
rect 17564 7890 17625 7893
rect 17564 7870 17573 7890
rect 17593 7873 17625 7890
rect 17646 7873 17651 7893
rect 17593 7870 17651 7873
rect 17564 7863 17651 7870
rect 17676 7890 17713 7960
rect 17979 7959 18016 7960
rect 17828 7900 17864 7901
rect 17676 7870 17685 7890
rect 17705 7870 17713 7890
rect 17564 7861 17620 7863
rect 17564 7860 17601 7861
rect 17676 7860 17713 7870
rect 17772 7890 17920 7900
rect 18020 7897 18116 7899
rect 17772 7870 17781 7890
rect 17801 7870 17891 7890
rect 17911 7870 17920 7890
rect 17772 7861 17920 7870
rect 17978 7890 18116 7897
rect 17978 7870 17987 7890
rect 18007 7870 18116 7890
rect 17978 7861 18116 7870
rect 17772 7860 17809 7861
rect 17828 7809 17864 7861
rect 17883 7860 17920 7861
rect 17979 7860 18016 7861
rect 16048 7790 16058 7808
rect 16076 7807 16681 7808
rect 17299 7807 17340 7808
rect 16076 7802 16097 7807
rect 16076 7790 16088 7802
rect 17191 7800 17340 7807
rect 16048 7782 16088 7790
rect 16131 7789 16157 7790
rect 16048 7780 16085 7782
rect 16131 7771 16685 7789
rect 17191 7780 17309 7800
rect 17329 7780 17340 7800
rect 17191 7772 17340 7780
rect 17407 7804 17766 7808
rect 17407 7799 17729 7804
rect 17407 7775 17520 7799
rect 17544 7780 17729 7799
rect 17753 7780 17766 7804
rect 17544 7775 17766 7780
rect 17407 7772 17766 7775
rect 17828 7772 17863 7809
rect 17931 7806 18031 7809
rect 17931 7802 17998 7806
rect 17931 7776 17943 7802
rect 17969 7780 17998 7802
rect 18024 7780 18031 7806
rect 17969 7776 18031 7780
rect 17931 7772 18031 7776
rect 15706 7762 15743 7771
rect 15418 7720 15455 7721
rect 15368 7711 15455 7720
rect 15368 7691 15426 7711
rect 15446 7691 15455 7711
rect 15368 7681 15455 7691
rect 15514 7711 15551 7721
rect 15514 7691 15522 7711
rect 15542 7691 15551 7711
rect 16051 7712 16088 7718
rect 16131 7712 16157 7771
rect 16664 7752 16685 7771
rect 16051 7709 16157 7712
rect 15709 7696 15746 7700
rect 15368 7680 15399 7681
rect 15514 7620 15551 7691
rect 15301 7596 15551 7620
rect 15707 7690 15746 7696
rect 15707 7672 15718 7690
rect 15736 7672 15746 7690
rect 16051 7691 16060 7709
rect 16078 7695 16157 7709
rect 16242 7727 16492 7751
rect 16078 7693 16154 7695
rect 16078 7691 16088 7693
rect 16051 7681 16088 7691
rect 15707 7663 15746 7672
rect 14457 7591 14494 7592
rect 13880 7570 13916 7591
rect 14306 7570 14337 7591
rect 15093 7572 15130 7595
rect 15707 7585 15742 7663
rect 16056 7616 16087 7681
rect 16242 7656 16279 7727
rect 16394 7666 16425 7667
rect 16242 7636 16251 7656
rect 16271 7636 16279 7656
rect 16242 7626 16279 7636
rect 16338 7656 16425 7666
rect 16338 7636 16347 7656
rect 16367 7636 16425 7656
rect 16338 7627 16425 7636
rect 16338 7626 16375 7627
rect 15704 7575 15742 7585
rect 16055 7607 16092 7616
rect 16055 7589 16065 7607
rect 16083 7589 16092 7607
rect 16055 7579 16092 7589
rect 15093 7571 15263 7572
rect 15704 7571 15714 7575
rect 13713 7566 13813 7570
rect 13713 7562 13775 7566
rect 13713 7536 13720 7562
rect 13746 7540 13775 7562
rect 13801 7540 13813 7566
rect 13746 7536 13813 7540
rect 13713 7533 13813 7536
rect 13881 7533 13916 7570
rect 13978 7567 14337 7570
rect 13978 7562 14200 7567
rect 13978 7538 13991 7562
rect 14015 7543 14200 7562
rect 14224 7543 14337 7567
rect 14015 7538 14337 7543
rect 13978 7534 14337 7538
rect 14404 7562 14553 7570
rect 14404 7542 14415 7562
rect 14435 7542 14553 7562
rect 15093 7557 15714 7571
rect 15732 7557 15742 7575
rect 16394 7574 16425 7627
rect 16455 7656 16492 7727
rect 16663 7732 17056 7752
rect 17076 7732 17079 7752
rect 17407 7751 17438 7772
rect 17828 7751 17864 7772
rect 17250 7750 17287 7751
rect 16663 7727 17079 7732
rect 17249 7741 17287 7750
rect 16663 7726 17004 7727
rect 16607 7666 16638 7667
rect 16455 7636 16464 7656
rect 16484 7636 16492 7656
rect 16455 7626 16492 7636
rect 16551 7659 16638 7666
rect 16551 7656 16612 7659
rect 16551 7636 16560 7656
rect 16580 7639 16612 7656
rect 16633 7639 16638 7659
rect 16580 7636 16638 7639
rect 16551 7629 16638 7636
rect 16663 7656 16700 7726
rect 16966 7725 17003 7726
rect 17249 7721 17258 7741
rect 17278 7721 17287 7741
rect 17249 7713 17287 7721
rect 17353 7745 17438 7751
rect 17463 7750 17500 7751
rect 17353 7725 17361 7745
rect 17381 7725 17438 7745
rect 17353 7717 17438 7725
rect 17462 7741 17500 7750
rect 17462 7721 17471 7741
rect 17491 7721 17500 7741
rect 17353 7716 17389 7717
rect 17462 7713 17500 7721
rect 17566 7745 17651 7751
rect 17671 7750 17708 7751
rect 17566 7725 17574 7745
rect 17594 7744 17651 7745
rect 17594 7725 17623 7744
rect 17566 7724 17623 7725
rect 17644 7724 17651 7744
rect 17566 7717 17651 7724
rect 17670 7741 17708 7750
rect 17670 7721 17679 7741
rect 17699 7721 17708 7741
rect 17566 7716 17602 7717
rect 17670 7713 17708 7721
rect 17774 7745 17918 7751
rect 17774 7725 17782 7745
rect 17802 7725 17834 7745
rect 17858 7725 17890 7745
rect 17910 7725 17918 7745
rect 17774 7717 17918 7725
rect 17774 7716 17810 7717
rect 17882 7716 17918 7717
rect 17984 7750 18021 7751
rect 17984 7749 18022 7750
rect 17984 7741 18048 7749
rect 17984 7721 17993 7741
rect 18013 7727 18048 7741
rect 18068 7727 18071 7747
rect 18013 7722 18071 7727
rect 18013 7721 18048 7722
rect 17250 7684 17287 7713
rect 17251 7682 17287 7684
rect 17463 7682 17500 7713
rect 16815 7666 16851 7667
rect 16663 7636 16672 7656
rect 16692 7636 16700 7656
rect 16551 7627 16607 7629
rect 16551 7626 16588 7627
rect 16663 7626 16700 7636
rect 16759 7656 16907 7666
rect 17007 7663 17103 7665
rect 16759 7636 16768 7656
rect 16788 7636 16878 7656
rect 16898 7636 16907 7656
rect 16759 7627 16907 7636
rect 16965 7656 17103 7663
rect 17251 7660 17500 7682
rect 17671 7681 17708 7713
rect 17984 7709 18048 7721
rect 18088 7683 18115 7861
rect 17947 7681 18115 7683
rect 17671 7677 18115 7681
rect 16965 7636 16974 7656
rect 16994 7636 17103 7656
rect 17671 7658 17720 7677
rect 17740 7658 18115 7677
rect 17671 7655 18115 7658
rect 17947 7654 18115 7655
rect 18815 7668 18844 7670
rect 18815 7663 18847 7668
rect 18815 7645 18822 7663
rect 18842 7645 18847 7663
rect 18908 7667 18939 8061
rect 18960 8086 19128 8087
rect 18960 8083 19404 8086
rect 18960 8064 19335 8083
rect 19355 8064 19404 8083
rect 19972 8085 20081 8105
rect 20101 8085 20110 8105
rect 18960 8060 19404 8064
rect 18960 8058 19128 8060
rect 18960 7880 18987 8058
rect 19027 8020 19091 8032
rect 19367 8028 19404 8060
rect 19575 8059 19824 8081
rect 19972 8078 20110 8085
rect 20168 8105 20316 8114
rect 20168 8085 20177 8105
rect 20197 8085 20287 8105
rect 20307 8085 20316 8105
rect 19972 8076 20068 8078
rect 20168 8075 20316 8085
rect 20375 8105 20412 8115
rect 20487 8114 20524 8115
rect 20468 8112 20524 8114
rect 20375 8085 20383 8105
rect 20403 8085 20412 8105
rect 20224 8074 20260 8075
rect 19575 8028 19612 8059
rect 19788 8057 19824 8059
rect 19788 8028 19825 8057
rect 19027 8019 19062 8020
rect 19004 8014 19062 8019
rect 19004 7994 19007 8014
rect 19027 8000 19062 8014
rect 19082 8000 19091 8020
rect 19027 7992 19091 8000
rect 19053 7991 19091 7992
rect 19054 7990 19091 7991
rect 19157 8024 19193 8025
rect 19265 8024 19301 8025
rect 19157 8016 19301 8024
rect 19157 7996 19165 8016
rect 19185 8015 19273 8016
rect 19185 7996 19218 8015
rect 19157 7995 19218 7996
rect 19242 7996 19273 8015
rect 19293 7996 19301 8016
rect 19242 7995 19301 7996
rect 19157 7990 19301 7995
rect 19367 8020 19405 8028
rect 19473 8024 19509 8025
rect 19367 8000 19376 8020
rect 19396 8000 19405 8020
rect 19367 7991 19405 8000
rect 19424 8017 19509 8024
rect 19424 7997 19431 8017
rect 19452 8016 19509 8017
rect 19452 7997 19481 8016
rect 19424 7996 19481 7997
rect 19501 7996 19509 8016
rect 19367 7990 19404 7991
rect 19424 7990 19509 7996
rect 19575 8020 19613 8028
rect 19686 8024 19722 8025
rect 19575 8000 19584 8020
rect 19604 8000 19613 8020
rect 19575 7991 19613 8000
rect 19637 8016 19722 8024
rect 19637 7996 19694 8016
rect 19714 7996 19722 8016
rect 19575 7990 19612 7991
rect 19637 7990 19722 7996
rect 19788 8020 19826 8028
rect 19788 8000 19797 8020
rect 19817 8000 19826 8020
rect 20072 8015 20109 8016
rect 20375 8015 20412 8085
rect 20437 8105 20524 8112
rect 20437 8102 20495 8105
rect 20437 8082 20442 8102
rect 20463 8085 20495 8102
rect 20515 8085 20524 8105
rect 20463 8082 20524 8085
rect 20437 8075 20524 8082
rect 20583 8105 20620 8115
rect 20583 8085 20591 8105
rect 20611 8085 20620 8105
rect 20437 8074 20468 8075
rect 20071 8014 20412 8015
rect 19788 7991 19826 8000
rect 19996 8009 20412 8014
rect 19788 7990 19825 7991
rect 19211 7969 19247 7990
rect 19637 7969 19668 7990
rect 19996 7989 19999 8009
rect 20019 7989 20412 8009
rect 20583 8014 20620 8085
rect 20650 8114 20681 8167
rect 20983 8152 21020 8162
rect 20983 8134 20992 8152
rect 21010 8134 21020 8152
rect 20983 8125 21020 8134
rect 20700 8114 20737 8115
rect 20650 8105 20737 8114
rect 20650 8085 20708 8105
rect 20728 8085 20737 8105
rect 20650 8075 20737 8085
rect 20796 8105 20833 8115
rect 20796 8085 20804 8105
rect 20824 8085 20833 8105
rect 20650 8074 20681 8075
rect 20796 8014 20833 8085
rect 20988 8060 21019 8125
rect 20987 8050 21024 8060
rect 20987 8048 20997 8050
rect 20921 8046 20997 8048
rect 20583 7990 20833 8014
rect 20918 8032 20997 8046
rect 21015 8032 21024 8050
rect 20918 8029 21024 8032
rect 20390 7970 20411 7989
rect 20918 7970 20944 8029
rect 20987 8023 21024 8029
rect 19044 7965 19144 7969
rect 19044 7961 19106 7965
rect 19044 7935 19051 7961
rect 19077 7939 19106 7961
rect 19132 7939 19144 7965
rect 19077 7935 19144 7939
rect 19044 7932 19144 7935
rect 19212 7932 19247 7969
rect 19309 7966 19668 7969
rect 19309 7961 19531 7966
rect 19309 7937 19322 7961
rect 19346 7942 19531 7961
rect 19555 7942 19668 7966
rect 19346 7937 19668 7942
rect 19309 7933 19668 7937
rect 19735 7961 19884 7969
rect 19735 7941 19746 7961
rect 19766 7941 19884 7961
rect 20390 7952 20944 7970
rect 20990 7959 21027 7961
rect 20918 7951 20944 7952
rect 20987 7951 21027 7959
rect 19735 7934 19884 7941
rect 20987 7939 20999 7951
rect 20978 7934 20999 7939
rect 19735 7933 19776 7934
rect 20394 7933 20999 7934
rect 21017 7933 21027 7951
rect 19059 7880 19096 7881
rect 19155 7880 19192 7881
rect 19211 7880 19247 7932
rect 19266 7880 19303 7881
rect 18959 7871 19097 7880
rect 18959 7851 19068 7871
rect 19088 7851 19097 7871
rect 18959 7844 19097 7851
rect 19155 7871 19303 7880
rect 19155 7851 19164 7871
rect 19184 7851 19274 7871
rect 19294 7851 19303 7871
rect 18959 7842 19055 7844
rect 19155 7841 19303 7851
rect 19362 7871 19399 7881
rect 19474 7880 19511 7881
rect 19455 7878 19511 7880
rect 19362 7851 19370 7871
rect 19390 7851 19399 7871
rect 19211 7840 19247 7841
rect 19059 7781 19096 7782
rect 19362 7781 19399 7851
rect 19424 7871 19511 7878
rect 19424 7868 19482 7871
rect 19424 7848 19429 7868
rect 19450 7851 19482 7868
rect 19502 7851 19511 7871
rect 19450 7848 19511 7851
rect 19424 7841 19511 7848
rect 19570 7871 19607 7881
rect 19570 7851 19578 7871
rect 19598 7851 19607 7871
rect 19424 7840 19455 7841
rect 19058 7780 19399 7781
rect 18983 7775 19399 7780
rect 18983 7755 18986 7775
rect 19006 7755 19399 7775
rect 19570 7780 19607 7851
rect 19637 7880 19668 7933
rect 20394 7924 21027 7933
rect 20394 7917 21026 7924
rect 20394 7915 20456 7917
rect 19972 7905 20140 7906
rect 20394 7905 20416 7915
rect 19687 7880 19724 7881
rect 19637 7871 19724 7880
rect 19637 7851 19695 7871
rect 19715 7851 19724 7871
rect 19637 7841 19724 7851
rect 19783 7871 19820 7881
rect 19783 7851 19791 7871
rect 19811 7851 19820 7871
rect 19637 7840 19668 7841
rect 19783 7780 19820 7851
rect 19570 7756 19820 7780
rect 19972 7879 20416 7905
rect 19972 7877 20140 7879
rect 19972 7699 19999 7877
rect 20039 7839 20103 7851
rect 20379 7847 20416 7879
rect 20587 7878 20836 7900
rect 20587 7847 20624 7878
rect 20800 7876 20836 7878
rect 20800 7847 20837 7876
rect 20039 7838 20074 7839
rect 20016 7833 20074 7838
rect 20016 7813 20019 7833
rect 20039 7819 20074 7833
rect 20094 7819 20103 7839
rect 20039 7811 20103 7819
rect 20065 7810 20103 7811
rect 20066 7809 20103 7810
rect 20169 7843 20205 7844
rect 20277 7843 20313 7844
rect 20169 7835 20313 7843
rect 20169 7815 20177 7835
rect 20197 7815 20226 7835
rect 20169 7814 20226 7815
rect 20248 7815 20285 7835
rect 20305 7815 20313 7835
rect 20248 7814 20313 7815
rect 20169 7809 20313 7814
rect 20379 7839 20417 7847
rect 20485 7843 20521 7844
rect 20379 7819 20388 7839
rect 20408 7819 20417 7839
rect 20379 7810 20417 7819
rect 20436 7836 20521 7843
rect 20436 7816 20443 7836
rect 20464 7835 20521 7836
rect 20464 7816 20493 7835
rect 20436 7815 20493 7816
rect 20513 7815 20521 7835
rect 20379 7809 20416 7810
rect 20436 7809 20521 7815
rect 20587 7839 20625 7847
rect 20698 7843 20734 7844
rect 20587 7819 20596 7839
rect 20616 7819 20625 7839
rect 20587 7810 20625 7819
rect 20649 7835 20734 7843
rect 20649 7815 20706 7835
rect 20726 7815 20734 7835
rect 20587 7809 20624 7810
rect 20649 7809 20734 7815
rect 20800 7839 20838 7847
rect 20800 7819 20809 7839
rect 20829 7819 20838 7839
rect 20800 7810 20838 7819
rect 20800 7809 20837 7810
rect 20223 7788 20259 7809
rect 20649 7788 20680 7809
rect 20056 7784 20156 7788
rect 20056 7780 20118 7784
rect 20056 7754 20063 7780
rect 20089 7758 20118 7780
rect 20144 7758 20156 7784
rect 20089 7754 20156 7758
rect 20056 7751 20156 7754
rect 20224 7751 20259 7788
rect 20321 7785 20680 7788
rect 20321 7780 20543 7785
rect 20321 7756 20334 7780
rect 20358 7761 20543 7780
rect 20567 7761 20680 7785
rect 20358 7756 20680 7761
rect 20321 7752 20680 7756
rect 20747 7780 20896 7788
rect 20747 7760 20758 7780
rect 20778 7760 20896 7780
rect 20747 7753 20896 7760
rect 20987 7768 21026 7917
rect 20747 7752 20788 7753
rect 20071 7699 20108 7700
rect 20167 7699 20204 7700
rect 20223 7699 20259 7751
rect 20278 7699 20315 7700
rect 19971 7690 20109 7699
rect 19971 7670 20080 7690
rect 20100 7670 20109 7690
rect 18908 7666 19078 7667
rect 18908 7651 19354 7666
rect 19971 7663 20109 7670
rect 20167 7690 20315 7699
rect 20167 7670 20176 7690
rect 20196 7670 20286 7690
rect 20306 7670 20315 7690
rect 19971 7661 20067 7663
rect 18815 7640 18847 7645
rect 16965 7627 17103 7636
rect 16759 7626 16796 7627
rect 16815 7575 16851 7627
rect 16870 7626 16907 7627
rect 16966 7626 17003 7627
rect 16286 7573 16327 7574
rect 15093 7551 15742 7557
rect 16178 7566 16327 7573
rect 15093 7550 15741 7551
rect 15704 7548 15741 7550
rect 14404 7535 14553 7542
rect 16178 7546 16296 7566
rect 16316 7546 16327 7566
rect 16178 7538 16327 7546
rect 16394 7570 16753 7574
rect 16394 7565 16716 7570
rect 16394 7541 16507 7565
rect 16531 7546 16716 7565
rect 16740 7546 16753 7570
rect 16531 7541 16753 7546
rect 16394 7538 16753 7541
rect 16815 7538 16850 7575
rect 16918 7572 17018 7575
rect 16918 7568 16985 7572
rect 16918 7542 16930 7568
rect 16956 7546 16985 7568
rect 17011 7546 17018 7572
rect 16956 7542 17018 7546
rect 16918 7538 17018 7542
rect 14404 7534 14445 7535
rect 13728 7481 13765 7482
rect 13824 7481 13861 7482
rect 13880 7481 13916 7533
rect 13935 7481 13972 7482
rect 13628 7472 13766 7481
rect 13628 7452 13737 7472
rect 13757 7452 13766 7472
rect 13628 7445 13766 7452
rect 13824 7472 13972 7481
rect 13824 7452 13833 7472
rect 13853 7452 13943 7472
rect 13963 7452 13972 7472
rect 13628 7443 13724 7445
rect 13824 7442 13972 7452
rect 14031 7472 14068 7482
rect 14143 7481 14180 7482
rect 14124 7479 14180 7481
rect 14031 7452 14039 7472
rect 14059 7452 14068 7472
rect 13880 7441 13916 7442
rect 13728 7382 13765 7383
rect 14031 7382 14068 7452
rect 14093 7472 14180 7479
rect 14093 7469 14151 7472
rect 14093 7449 14098 7469
rect 14119 7452 14151 7469
rect 14171 7452 14180 7472
rect 14119 7449 14180 7452
rect 14093 7442 14180 7449
rect 14239 7472 14276 7482
rect 14239 7452 14247 7472
rect 14267 7452 14276 7472
rect 14093 7441 14124 7442
rect 13727 7381 14068 7382
rect 13652 7376 14068 7381
rect 13652 7356 13655 7376
rect 13675 7356 14068 7376
rect 14239 7381 14276 7452
rect 14306 7481 14337 7534
rect 16394 7517 16425 7538
rect 16815 7517 16851 7538
rect 16058 7508 16095 7517
rect 16237 7516 16274 7517
rect 16058 7490 16067 7508
rect 16085 7490 16095 7508
rect 14356 7481 14393 7482
rect 14306 7472 14393 7481
rect 14306 7452 14364 7472
rect 14384 7452 14393 7472
rect 14306 7442 14393 7452
rect 14452 7472 14489 7482
rect 14452 7452 14460 7472
rect 14480 7452 14489 7472
rect 14306 7441 14337 7442
rect 14452 7381 14489 7452
rect 15707 7476 15744 7486
rect 16058 7480 16095 7490
rect 15707 7458 15716 7476
rect 15734 7458 15744 7476
rect 15707 7449 15744 7458
rect 15707 7425 15742 7449
rect 16059 7445 16095 7480
rect 16236 7507 16274 7516
rect 16236 7487 16245 7507
rect 16265 7487 16274 7507
rect 16236 7479 16274 7487
rect 16340 7511 16425 7517
rect 16450 7516 16487 7517
rect 16340 7491 16348 7511
rect 16368 7491 16425 7511
rect 16340 7483 16425 7491
rect 16449 7507 16487 7516
rect 16449 7487 16458 7507
rect 16478 7487 16487 7507
rect 16340 7482 16376 7483
rect 16449 7479 16487 7487
rect 16553 7511 16638 7517
rect 16658 7516 16695 7517
rect 16553 7491 16561 7511
rect 16581 7510 16638 7511
rect 16581 7491 16610 7510
rect 16553 7490 16610 7491
rect 16631 7490 16638 7510
rect 16553 7483 16638 7490
rect 16657 7507 16695 7516
rect 16657 7487 16666 7507
rect 16686 7487 16695 7507
rect 16553 7482 16589 7483
rect 16657 7479 16695 7487
rect 16761 7511 16905 7517
rect 16761 7491 16769 7511
rect 16789 7510 16877 7511
rect 16789 7491 16817 7510
rect 16761 7489 16817 7491
rect 16839 7491 16877 7510
rect 16897 7491 16905 7511
rect 16839 7489 16905 7491
rect 16761 7483 16905 7489
rect 16761 7482 16797 7483
rect 16869 7482 16905 7483
rect 16971 7516 17008 7517
rect 16971 7515 17009 7516
rect 16971 7507 17035 7515
rect 16971 7487 16980 7507
rect 17000 7493 17035 7507
rect 17055 7493 17058 7513
rect 17000 7488 17058 7493
rect 17000 7487 17035 7488
rect 16237 7450 16274 7479
rect 15705 7401 15742 7425
rect 15704 7395 15742 7401
rect 14239 7357 14489 7381
rect 15115 7377 15742 7395
rect 14697 7360 14865 7361
rect 15116 7360 15140 7377
rect 14697 7334 15141 7360
rect 14697 7332 14865 7334
rect 14697 7154 14724 7332
rect 14764 7294 14828 7306
rect 15104 7302 15141 7334
rect 15312 7333 15561 7355
rect 15312 7302 15349 7333
rect 15525 7331 15561 7333
rect 15704 7336 15742 7377
rect 16057 7404 16095 7445
rect 16238 7448 16274 7450
rect 16450 7448 16487 7479
rect 16238 7426 16487 7448
rect 16658 7447 16695 7479
rect 16971 7475 17035 7487
rect 17075 7449 17102 7627
rect 16934 7447 17102 7449
rect 16658 7421 17102 7447
rect 16659 7404 16683 7421
rect 16934 7420 17102 7421
rect 16057 7386 16684 7404
rect 17310 7400 17560 7424
rect 16057 7380 16095 7386
rect 16057 7356 16094 7380
rect 15525 7302 15562 7331
rect 14764 7293 14799 7294
rect 14741 7288 14799 7293
rect 14741 7268 14744 7288
rect 14764 7274 14799 7288
rect 14819 7274 14828 7294
rect 14764 7266 14828 7274
rect 14790 7265 14828 7266
rect 14791 7264 14828 7265
rect 14894 7298 14930 7299
rect 15002 7298 15038 7299
rect 14894 7292 15038 7298
rect 14894 7290 14960 7292
rect 14894 7270 14902 7290
rect 14922 7271 14960 7290
rect 14982 7290 15038 7292
rect 14982 7271 15010 7290
rect 14922 7270 15010 7271
rect 15030 7270 15038 7290
rect 14894 7264 15038 7270
rect 15104 7294 15142 7302
rect 15210 7298 15246 7299
rect 15104 7274 15113 7294
rect 15133 7274 15142 7294
rect 15104 7265 15142 7274
rect 15161 7291 15246 7298
rect 15161 7271 15168 7291
rect 15189 7290 15246 7291
rect 15189 7271 15218 7290
rect 15161 7270 15218 7271
rect 15238 7270 15246 7290
rect 15104 7264 15141 7265
rect 15161 7264 15246 7270
rect 15312 7294 15350 7302
rect 15423 7298 15459 7299
rect 15312 7274 15321 7294
rect 15341 7274 15350 7294
rect 15312 7265 15350 7274
rect 15374 7290 15459 7298
rect 15374 7270 15431 7290
rect 15451 7270 15459 7290
rect 15312 7264 15349 7265
rect 15374 7264 15459 7270
rect 15525 7294 15563 7302
rect 15525 7274 15534 7294
rect 15554 7274 15563 7294
rect 15525 7265 15563 7274
rect 15704 7301 15740 7336
rect 16057 7332 16092 7356
rect 16055 7323 16092 7332
rect 16055 7305 16065 7323
rect 16083 7305 16092 7323
rect 15704 7291 15741 7301
rect 16055 7295 16092 7305
rect 17310 7329 17347 7400
rect 17462 7339 17493 7340
rect 17310 7309 17319 7329
rect 17339 7309 17347 7329
rect 17310 7299 17347 7309
rect 17406 7329 17493 7339
rect 17406 7309 17415 7329
rect 17435 7309 17493 7329
rect 17406 7300 17493 7309
rect 17406 7299 17443 7300
rect 15704 7273 15714 7291
rect 15732 7273 15741 7291
rect 15525 7264 15562 7265
rect 15704 7264 15741 7273
rect 14948 7243 14984 7264
rect 15374 7243 15405 7264
rect 17462 7247 17493 7300
rect 17523 7329 17560 7400
rect 17731 7405 18124 7425
rect 18144 7405 18147 7425
rect 17731 7400 18147 7405
rect 17731 7399 18072 7400
rect 17675 7339 17706 7340
rect 17523 7309 17532 7329
rect 17552 7309 17560 7329
rect 17523 7299 17560 7309
rect 17619 7332 17706 7339
rect 17619 7329 17680 7332
rect 17619 7309 17628 7329
rect 17648 7312 17680 7329
rect 17701 7312 17706 7332
rect 17648 7309 17706 7312
rect 17619 7302 17706 7309
rect 17731 7329 17768 7399
rect 18034 7398 18071 7399
rect 17883 7339 17919 7340
rect 17731 7309 17740 7329
rect 17760 7309 17768 7329
rect 17619 7300 17675 7302
rect 17619 7299 17656 7300
rect 17731 7299 17768 7309
rect 17827 7329 17975 7339
rect 18075 7336 18171 7338
rect 17827 7309 17836 7329
rect 17856 7309 17946 7329
rect 17966 7309 17975 7329
rect 17827 7300 17975 7309
rect 18033 7329 18171 7336
rect 18033 7309 18042 7329
rect 18062 7309 18171 7329
rect 18033 7300 18171 7309
rect 17827 7299 17864 7300
rect 17883 7248 17919 7300
rect 17938 7299 17975 7300
rect 18034 7299 18071 7300
rect 17354 7246 17395 7247
rect 14781 7239 14881 7243
rect 14781 7235 14843 7239
rect 14781 7209 14788 7235
rect 14814 7213 14843 7235
rect 14869 7213 14881 7239
rect 14814 7209 14881 7213
rect 14781 7206 14881 7209
rect 14949 7206 14984 7243
rect 15046 7240 15405 7243
rect 15046 7235 15268 7240
rect 15046 7211 15059 7235
rect 15083 7216 15268 7235
rect 15292 7216 15405 7240
rect 15083 7211 15405 7216
rect 15046 7207 15405 7211
rect 15472 7235 15621 7243
rect 15472 7215 15483 7235
rect 15503 7215 15621 7235
rect 17246 7239 17395 7246
rect 16058 7231 16095 7233
rect 16058 7230 16706 7231
rect 15472 7208 15621 7215
rect 16057 7224 16706 7230
rect 15472 7207 15513 7208
rect 14796 7154 14833 7155
rect 14892 7154 14929 7155
rect 14948 7154 14984 7206
rect 15003 7154 15040 7155
rect 14696 7145 14834 7154
rect 13684 7126 13852 7127
rect 13684 7123 14128 7126
rect 13684 7104 14059 7123
rect 14079 7104 14128 7123
rect 14696 7125 14805 7145
rect 14825 7125 14834 7145
rect 13684 7100 14128 7104
rect 13684 7098 13852 7100
rect 13684 6920 13711 7098
rect 13751 7060 13815 7072
rect 14091 7068 14128 7100
rect 14299 7099 14548 7121
rect 14696 7118 14834 7125
rect 14892 7145 15040 7154
rect 14892 7125 14901 7145
rect 14921 7125 15011 7145
rect 15031 7125 15040 7145
rect 14696 7116 14792 7118
rect 14892 7115 15040 7125
rect 15099 7145 15136 7155
rect 15211 7154 15248 7155
rect 15192 7152 15248 7154
rect 15099 7125 15107 7145
rect 15127 7125 15136 7145
rect 14948 7114 14984 7115
rect 14299 7068 14336 7099
rect 14512 7097 14548 7099
rect 14512 7068 14549 7097
rect 13751 7059 13786 7060
rect 13728 7054 13786 7059
rect 13728 7034 13731 7054
rect 13751 7040 13786 7054
rect 13806 7040 13815 7060
rect 13751 7032 13815 7040
rect 13777 7031 13815 7032
rect 13778 7030 13815 7031
rect 13881 7064 13917 7065
rect 13989 7064 14025 7065
rect 13881 7056 14025 7064
rect 13881 7036 13889 7056
rect 13909 7036 13941 7056
rect 13965 7036 13997 7056
rect 14017 7036 14025 7056
rect 13881 7030 14025 7036
rect 14091 7060 14129 7068
rect 14197 7064 14233 7065
rect 14091 7040 14100 7060
rect 14120 7040 14129 7060
rect 14091 7031 14129 7040
rect 14148 7057 14233 7064
rect 14148 7037 14155 7057
rect 14176 7056 14233 7057
rect 14176 7037 14205 7056
rect 14148 7036 14205 7037
rect 14225 7036 14233 7056
rect 14091 7030 14128 7031
rect 14148 7030 14233 7036
rect 14299 7060 14337 7068
rect 14410 7064 14446 7065
rect 14299 7040 14308 7060
rect 14328 7040 14337 7060
rect 14299 7031 14337 7040
rect 14361 7056 14446 7064
rect 14361 7036 14418 7056
rect 14438 7036 14446 7056
rect 14299 7030 14336 7031
rect 14361 7030 14446 7036
rect 14512 7060 14550 7068
rect 14512 7040 14521 7060
rect 14541 7040 14550 7060
rect 14796 7055 14833 7056
rect 15099 7055 15136 7125
rect 15161 7145 15248 7152
rect 15161 7142 15219 7145
rect 15161 7122 15166 7142
rect 15187 7125 15219 7142
rect 15239 7125 15248 7145
rect 15187 7122 15248 7125
rect 15161 7115 15248 7122
rect 15307 7145 15344 7155
rect 15307 7125 15315 7145
rect 15335 7125 15344 7145
rect 15161 7114 15192 7115
rect 14795 7054 15136 7055
rect 14512 7031 14550 7040
rect 14720 7049 15136 7054
rect 14512 7030 14549 7031
rect 13935 7009 13971 7030
rect 14361 7009 14392 7030
rect 14720 7029 14723 7049
rect 14743 7029 15136 7049
rect 15307 7054 15344 7125
rect 15374 7154 15405 7207
rect 16057 7206 16067 7224
rect 16085 7210 16706 7224
rect 17246 7219 17364 7239
rect 17384 7219 17395 7239
rect 17246 7211 17395 7219
rect 17462 7243 17821 7247
rect 17462 7238 17784 7243
rect 17462 7214 17575 7238
rect 17599 7219 17784 7238
rect 17808 7219 17821 7243
rect 17599 7214 17821 7219
rect 17462 7211 17821 7214
rect 17883 7211 17918 7248
rect 17986 7245 18086 7248
rect 17986 7241 18053 7245
rect 17986 7215 17998 7241
rect 18024 7219 18053 7241
rect 18079 7219 18086 7245
rect 18024 7215 18086 7219
rect 17986 7211 18086 7215
rect 16085 7206 16095 7210
rect 16536 7209 16706 7210
rect 15707 7192 15744 7202
rect 15707 7174 15716 7192
rect 15734 7174 15744 7192
rect 15707 7165 15744 7174
rect 16057 7196 16095 7206
rect 15424 7154 15461 7155
rect 15374 7145 15461 7154
rect 15374 7125 15432 7145
rect 15452 7125 15461 7145
rect 15374 7115 15461 7125
rect 15520 7145 15557 7155
rect 15520 7125 15528 7145
rect 15548 7125 15557 7145
rect 15374 7114 15405 7115
rect 15520 7054 15557 7125
rect 15712 7100 15743 7165
rect 16057 7118 16092 7196
rect 16669 7186 16706 7209
rect 17462 7190 17493 7211
rect 17883 7190 17919 7211
rect 17305 7189 17342 7190
rect 16053 7109 16092 7118
rect 15711 7090 15748 7100
rect 15711 7088 15721 7090
rect 15645 7086 15721 7088
rect 15307 7030 15557 7054
rect 15642 7072 15721 7086
rect 15739 7072 15748 7090
rect 16053 7091 16063 7109
rect 16081 7091 16092 7109
rect 16053 7085 16092 7091
rect 16248 7161 16498 7185
rect 16248 7090 16285 7161
rect 16400 7100 16431 7101
rect 16053 7081 16090 7085
rect 15642 7069 15748 7072
rect 15114 7010 15135 7029
rect 15642 7010 15668 7069
rect 15711 7063 15748 7069
rect 16248 7070 16257 7090
rect 16277 7070 16285 7090
rect 16248 7060 16285 7070
rect 16344 7090 16431 7100
rect 16344 7070 16353 7090
rect 16373 7070 16431 7090
rect 16344 7061 16431 7070
rect 16344 7060 16381 7061
rect 16056 7010 16093 7019
rect 13768 7005 13868 7009
rect 13768 7001 13830 7005
rect 13768 6975 13775 7001
rect 13801 6979 13830 7001
rect 13856 6979 13868 7005
rect 13801 6975 13868 6979
rect 13768 6972 13868 6975
rect 13936 6972 13971 7009
rect 14033 7006 14392 7009
rect 14033 7001 14255 7006
rect 14033 6977 14046 7001
rect 14070 6982 14255 7001
rect 14279 6982 14392 7006
rect 14070 6977 14392 6982
rect 14033 6973 14392 6977
rect 14459 7001 14608 7009
rect 14459 6981 14470 7001
rect 14490 6981 14608 7001
rect 15114 6992 15668 7010
rect 15714 6999 15751 7001
rect 15642 6991 15668 6992
rect 15711 6991 15751 6999
rect 14459 6974 14608 6981
rect 15711 6979 15723 6991
rect 15702 6974 15723 6979
rect 14459 6973 14500 6974
rect 15118 6973 15723 6974
rect 15741 6973 15751 6991
rect 13783 6920 13820 6921
rect 13879 6920 13916 6921
rect 13935 6920 13971 6972
rect 13990 6920 14027 6921
rect 13683 6911 13821 6920
rect 13683 6891 13792 6911
rect 13812 6891 13821 6911
rect 13683 6884 13821 6891
rect 13879 6911 14027 6920
rect 13879 6891 13888 6911
rect 13908 6891 13998 6911
rect 14018 6891 14027 6911
rect 13683 6882 13779 6884
rect 13879 6881 14027 6891
rect 14086 6911 14123 6921
rect 14198 6920 14235 6921
rect 14179 6918 14235 6920
rect 14086 6891 14094 6911
rect 14114 6891 14123 6911
rect 13935 6880 13971 6881
rect 13783 6821 13820 6822
rect 14086 6821 14123 6891
rect 14148 6911 14235 6918
rect 14148 6908 14206 6911
rect 14148 6888 14153 6908
rect 14174 6891 14206 6908
rect 14226 6891 14235 6911
rect 14174 6888 14235 6891
rect 14148 6881 14235 6888
rect 14294 6911 14331 6921
rect 14294 6891 14302 6911
rect 14322 6891 14331 6911
rect 14148 6880 14179 6881
rect 13782 6820 14123 6821
rect 13707 6815 14123 6820
rect 13707 6795 13710 6815
rect 13730 6795 14123 6815
rect 14294 6820 14331 6891
rect 14361 6920 14392 6973
rect 15118 6964 15751 6973
rect 16054 6992 16065 7010
rect 16083 6992 16093 7010
rect 16400 7008 16431 7061
rect 16461 7090 16498 7161
rect 16669 7166 17062 7186
rect 17082 7166 17085 7186
rect 16669 7161 17085 7166
rect 17304 7180 17342 7189
rect 16669 7160 17010 7161
rect 17304 7160 17313 7180
rect 17333 7160 17342 7180
rect 16613 7100 16644 7101
rect 16461 7070 16470 7090
rect 16490 7070 16498 7090
rect 16461 7060 16498 7070
rect 16557 7093 16644 7100
rect 16557 7090 16618 7093
rect 16557 7070 16566 7090
rect 16586 7073 16618 7090
rect 16639 7073 16644 7093
rect 16586 7070 16644 7073
rect 16557 7063 16644 7070
rect 16669 7090 16706 7160
rect 16972 7159 17009 7160
rect 17304 7152 17342 7160
rect 17408 7184 17493 7190
rect 17518 7189 17555 7190
rect 17408 7164 17416 7184
rect 17436 7164 17493 7184
rect 17408 7156 17493 7164
rect 17517 7180 17555 7189
rect 17517 7160 17526 7180
rect 17546 7160 17555 7180
rect 17408 7155 17444 7156
rect 17517 7152 17555 7160
rect 17621 7184 17706 7190
rect 17726 7189 17763 7190
rect 17621 7164 17629 7184
rect 17649 7183 17706 7184
rect 17649 7164 17678 7183
rect 17621 7163 17678 7164
rect 17699 7163 17706 7183
rect 17621 7156 17706 7163
rect 17725 7180 17763 7189
rect 17725 7160 17734 7180
rect 17754 7160 17763 7180
rect 17621 7155 17657 7156
rect 17725 7152 17763 7160
rect 17829 7184 17973 7190
rect 17829 7164 17837 7184
rect 17857 7182 17945 7184
rect 17857 7165 17893 7182
rect 17917 7165 17945 7182
rect 17857 7164 17945 7165
rect 17965 7164 17973 7184
rect 17829 7156 17973 7164
rect 17829 7155 17865 7156
rect 17937 7155 17973 7156
rect 18039 7189 18076 7190
rect 18039 7188 18077 7189
rect 18039 7180 18103 7188
rect 18039 7160 18048 7180
rect 18068 7166 18103 7180
rect 18123 7166 18126 7186
rect 18068 7161 18126 7166
rect 18068 7160 18103 7161
rect 17305 7123 17342 7152
rect 17306 7121 17342 7123
rect 17518 7121 17555 7152
rect 16821 7100 16857 7101
rect 16669 7070 16678 7090
rect 16698 7070 16706 7090
rect 16557 7061 16613 7063
rect 16557 7060 16594 7061
rect 16669 7060 16706 7070
rect 16765 7090 16913 7100
rect 17306 7099 17555 7121
rect 17726 7120 17763 7152
rect 18039 7148 18103 7160
rect 18143 7122 18170 7300
rect 18002 7120 18170 7122
rect 17726 7109 18170 7120
rect 17013 7097 17109 7099
rect 16765 7070 16774 7090
rect 16794 7070 16884 7090
rect 16904 7070 16913 7090
rect 16765 7061 16913 7070
rect 16971 7090 17109 7097
rect 17726 7094 18172 7109
rect 18002 7093 18172 7094
rect 16971 7070 16980 7090
rect 17000 7070 17109 7090
rect 16971 7061 17109 7070
rect 16765 7060 16802 7061
rect 16821 7009 16857 7061
rect 16876 7060 16913 7061
rect 16972 7060 17009 7061
rect 16292 7007 16333 7008
rect 15118 6957 15750 6964
rect 15118 6955 15180 6957
rect 14696 6945 14864 6946
rect 15118 6945 15140 6955
rect 14411 6920 14448 6921
rect 14361 6911 14448 6920
rect 14361 6891 14419 6911
rect 14439 6891 14448 6911
rect 14361 6881 14448 6891
rect 14507 6911 14544 6921
rect 14507 6891 14515 6911
rect 14535 6891 14544 6911
rect 14361 6880 14392 6881
rect 14507 6820 14544 6891
rect 14294 6796 14544 6820
rect 14696 6919 15140 6945
rect 14696 6917 14864 6919
rect 14696 6739 14723 6917
rect 14763 6879 14827 6891
rect 15103 6887 15140 6919
rect 15311 6918 15560 6940
rect 15311 6887 15348 6918
rect 15524 6916 15560 6918
rect 15524 6887 15561 6916
rect 14763 6878 14798 6879
rect 14740 6873 14798 6878
rect 14740 6853 14743 6873
rect 14763 6859 14798 6873
rect 14818 6859 14827 6879
rect 14763 6851 14827 6859
rect 14789 6850 14827 6851
rect 14790 6849 14827 6850
rect 14893 6883 14929 6884
rect 15001 6883 15037 6884
rect 14893 6875 15037 6883
rect 14893 6855 14901 6875
rect 14921 6855 14950 6875
rect 14893 6854 14950 6855
rect 14972 6855 15009 6875
rect 15029 6855 15037 6875
rect 14972 6854 15037 6855
rect 14893 6849 15037 6854
rect 15103 6879 15141 6887
rect 15209 6883 15245 6884
rect 15103 6859 15112 6879
rect 15132 6859 15141 6879
rect 15103 6850 15141 6859
rect 15160 6876 15245 6883
rect 15160 6856 15167 6876
rect 15188 6875 15245 6876
rect 15188 6856 15217 6875
rect 15160 6855 15217 6856
rect 15237 6855 15245 6875
rect 15103 6849 15140 6850
rect 15160 6849 15245 6855
rect 15311 6879 15349 6887
rect 15422 6883 15458 6884
rect 15311 6859 15320 6879
rect 15340 6859 15349 6879
rect 15311 6850 15349 6859
rect 15373 6875 15458 6883
rect 15373 6855 15430 6875
rect 15450 6855 15458 6875
rect 15311 6849 15348 6850
rect 15373 6849 15458 6855
rect 15524 6879 15562 6887
rect 15524 6859 15533 6879
rect 15553 6859 15562 6879
rect 15524 6850 15562 6859
rect 15524 6849 15561 6850
rect 14947 6828 14983 6849
rect 15373 6828 15404 6849
rect 14780 6824 14880 6828
rect 14780 6820 14842 6824
rect 14780 6794 14787 6820
rect 14813 6798 14842 6820
rect 14868 6798 14880 6824
rect 14813 6794 14880 6798
rect 14780 6791 14880 6794
rect 14948 6791 14983 6828
rect 15045 6825 15404 6828
rect 15045 6820 15267 6825
rect 15045 6796 15058 6820
rect 15082 6801 15267 6820
rect 15291 6801 15404 6825
rect 15082 6796 15404 6801
rect 15045 6792 15404 6796
rect 15471 6820 15620 6828
rect 15471 6800 15482 6820
rect 15502 6800 15620 6820
rect 15471 6793 15620 6800
rect 15711 6808 15750 6957
rect 16054 6843 16093 6992
rect 16184 7000 16333 7007
rect 16184 6980 16302 7000
rect 16322 6980 16333 7000
rect 16184 6972 16333 6980
rect 16400 7004 16759 7008
rect 16400 6999 16722 7004
rect 16400 6975 16513 6999
rect 16537 6980 16722 6999
rect 16746 6980 16759 7004
rect 16537 6975 16759 6980
rect 16400 6972 16759 6975
rect 16821 6972 16856 7009
rect 16924 7006 17024 7009
rect 16924 7002 16991 7006
rect 16924 6976 16936 7002
rect 16962 6980 16991 7002
rect 17017 6980 17024 7006
rect 16962 6976 17024 6980
rect 16924 6972 17024 6976
rect 16400 6951 16431 6972
rect 16821 6951 16857 6972
rect 16243 6950 16280 6951
rect 16242 6941 16280 6950
rect 16242 6921 16251 6941
rect 16271 6921 16280 6941
rect 16242 6913 16280 6921
rect 16346 6945 16431 6951
rect 16456 6950 16493 6951
rect 16346 6925 16354 6945
rect 16374 6925 16431 6945
rect 16346 6917 16431 6925
rect 16455 6941 16493 6950
rect 16455 6921 16464 6941
rect 16484 6921 16493 6941
rect 16346 6916 16382 6917
rect 16455 6913 16493 6921
rect 16559 6945 16644 6951
rect 16664 6950 16701 6951
rect 16559 6925 16567 6945
rect 16587 6944 16644 6945
rect 16587 6925 16616 6944
rect 16559 6924 16616 6925
rect 16637 6924 16644 6944
rect 16559 6917 16644 6924
rect 16663 6941 16701 6950
rect 16663 6921 16672 6941
rect 16692 6921 16701 6941
rect 16559 6916 16595 6917
rect 16663 6913 16701 6921
rect 16767 6946 16911 6951
rect 16767 6945 16832 6946
rect 16767 6925 16775 6945
rect 16795 6925 16832 6945
rect 16854 6945 16911 6946
rect 16854 6925 16883 6945
rect 16903 6925 16911 6945
rect 16767 6917 16911 6925
rect 16767 6916 16803 6917
rect 16875 6916 16911 6917
rect 16977 6950 17014 6951
rect 16977 6949 17015 6950
rect 16977 6941 17041 6949
rect 16977 6921 16986 6941
rect 17006 6927 17041 6941
rect 17061 6927 17064 6947
rect 17006 6922 17064 6927
rect 17006 6921 17041 6922
rect 16243 6884 16280 6913
rect 16244 6882 16280 6884
rect 16456 6882 16493 6913
rect 16244 6860 16493 6882
rect 16664 6881 16701 6913
rect 16977 6909 17041 6921
rect 17081 6883 17108 7061
rect 16940 6881 17108 6883
rect 16664 6855 17108 6881
rect 17260 6980 17510 7004
rect 17260 6909 17297 6980
rect 17412 6919 17443 6920
rect 17260 6889 17269 6909
rect 17289 6889 17297 6909
rect 17260 6879 17297 6889
rect 17356 6909 17443 6919
rect 17356 6889 17365 6909
rect 17385 6889 17443 6909
rect 17356 6880 17443 6889
rect 17356 6879 17393 6880
rect 16664 6845 16686 6855
rect 16940 6854 17108 6855
rect 16624 6843 16686 6845
rect 16054 6836 16686 6843
rect 15471 6792 15512 6793
rect 14795 6739 14832 6740
rect 14891 6739 14928 6740
rect 14947 6739 14983 6791
rect 15002 6739 15039 6740
rect 14695 6730 14833 6739
rect 14695 6710 14804 6730
rect 14824 6710 14833 6730
rect 14695 6703 14833 6710
rect 14891 6730 15039 6739
rect 14891 6710 14900 6730
rect 14920 6710 15010 6730
rect 15030 6710 15039 6730
rect 14695 6701 14791 6703
rect 14891 6700 15039 6710
rect 15098 6730 15135 6740
rect 15210 6739 15247 6740
rect 15191 6737 15247 6739
rect 15098 6710 15106 6730
rect 15126 6710 15135 6730
rect 14947 6699 14983 6700
rect 13410 6637 13418 6656
rect 13441 6637 13447 6656
rect 13410 6626 13447 6637
rect 13476 6659 13644 6660
rect 13476 6633 13920 6659
rect 13476 6631 13644 6633
rect 13413 6566 13446 6626
rect 11658 6487 11826 6489
rect 11382 6461 11826 6487
rect 11383 6444 11407 6461
rect 11658 6460 11826 6461
rect 12194 6489 12444 6513
rect 8823 6424 8860 6425
rect 8773 6415 8860 6424
rect 8773 6395 8831 6415
rect 8851 6395 8860 6415
rect 8773 6385 8860 6395
rect 8919 6415 8956 6425
rect 8919 6395 8927 6415
rect 8947 6395 8956 6415
rect 8773 6384 8804 6385
rect 8919 6324 8956 6395
rect 10332 6393 10367 6439
rect 10781 6426 11408 6444
rect 10781 6420 10819 6426
rect 10331 6387 10369 6393
rect 9742 6369 10369 6387
rect 10783 6374 10818 6420
rect 12194 6418 12231 6489
rect 12346 6428 12377 6429
rect 12194 6398 12203 6418
rect 12223 6398 12231 6418
rect 12194 6388 12231 6398
rect 12290 6418 12377 6428
rect 12290 6398 12299 6418
rect 12319 6398 12377 6418
rect 12290 6389 12377 6398
rect 12290 6388 12327 6389
rect 8706 6300 8956 6324
rect 9324 6352 9492 6353
rect 9743 6352 9767 6369
rect 9324 6326 9768 6352
rect 9324 6324 9492 6326
rect 9324 6146 9351 6324
rect 9391 6286 9455 6298
rect 9731 6294 9768 6326
rect 9939 6325 10188 6347
rect 9939 6294 9976 6325
rect 10152 6323 10188 6325
rect 10331 6328 10369 6369
rect 10781 6365 10818 6374
rect 10781 6347 10791 6365
rect 10809 6347 10818 6365
rect 10781 6337 10818 6347
rect 12346 6336 12377 6389
rect 12407 6418 12444 6489
rect 12615 6494 13008 6514
rect 13028 6494 13031 6514
rect 12615 6489 13031 6494
rect 12615 6488 12956 6489
rect 12559 6428 12590 6429
rect 12407 6398 12416 6418
rect 12436 6398 12444 6418
rect 12407 6388 12444 6398
rect 12503 6421 12590 6428
rect 12503 6418 12564 6421
rect 12503 6398 12512 6418
rect 12532 6401 12564 6418
rect 12585 6401 12590 6421
rect 12532 6398 12590 6401
rect 12503 6391 12590 6398
rect 12615 6418 12652 6488
rect 12918 6487 12955 6488
rect 12767 6428 12803 6429
rect 12615 6398 12624 6418
rect 12644 6398 12652 6418
rect 12503 6389 12559 6391
rect 12503 6388 12540 6389
rect 12615 6388 12652 6398
rect 12711 6418 12859 6428
rect 12959 6425 13055 6427
rect 12711 6398 12720 6418
rect 12740 6398 12830 6418
rect 12850 6398 12859 6418
rect 12711 6389 12859 6398
rect 12917 6418 13055 6425
rect 12917 6398 12926 6418
rect 12946 6398 13055 6418
rect 12917 6389 13055 6398
rect 12711 6388 12748 6389
rect 12767 6337 12803 6389
rect 12822 6388 12859 6389
rect 12918 6388 12955 6389
rect 12238 6335 12279 6336
rect 12130 6328 12279 6335
rect 10152 6294 10189 6323
rect 9391 6285 9426 6286
rect 9368 6280 9426 6285
rect 9368 6260 9371 6280
rect 9391 6266 9426 6280
rect 9446 6266 9455 6286
rect 9391 6258 9455 6266
rect 9417 6257 9455 6258
rect 9418 6256 9455 6257
rect 9521 6290 9557 6291
rect 9629 6290 9665 6291
rect 9521 6284 9665 6290
rect 9521 6282 9587 6284
rect 9521 6262 9529 6282
rect 9549 6263 9587 6282
rect 9609 6282 9665 6284
rect 9609 6263 9637 6282
rect 9549 6262 9637 6263
rect 9657 6262 9665 6282
rect 9521 6256 9665 6262
rect 9731 6286 9769 6294
rect 9837 6290 9873 6291
rect 9731 6266 9740 6286
rect 9760 6266 9769 6286
rect 9731 6257 9769 6266
rect 9788 6283 9873 6290
rect 9788 6263 9795 6283
rect 9816 6282 9873 6283
rect 9816 6263 9845 6282
rect 9788 6262 9845 6263
rect 9865 6262 9873 6282
rect 9731 6256 9768 6257
rect 9788 6256 9873 6262
rect 9939 6286 9977 6294
rect 10050 6290 10086 6291
rect 9939 6266 9948 6286
rect 9968 6266 9977 6286
rect 9939 6257 9977 6266
rect 10001 6282 10086 6290
rect 10001 6262 10058 6282
rect 10078 6262 10086 6282
rect 9939 6256 9976 6257
rect 10001 6256 10086 6262
rect 10152 6286 10190 6294
rect 10152 6266 10161 6286
rect 10181 6266 10190 6286
rect 10152 6257 10190 6266
rect 10331 6293 10367 6328
rect 12130 6308 12248 6328
rect 12268 6308 12279 6328
rect 12130 6300 12279 6308
rect 12346 6332 12705 6336
rect 12346 6327 12668 6332
rect 12346 6303 12459 6327
rect 12483 6308 12668 6327
rect 12692 6308 12705 6332
rect 12483 6303 12705 6308
rect 12346 6300 12705 6303
rect 12767 6300 12802 6337
rect 12870 6334 12970 6337
rect 12870 6330 12937 6334
rect 12870 6304 12882 6330
rect 12908 6308 12937 6330
rect 12963 6308 12970 6334
rect 12908 6304 12970 6308
rect 12870 6300 12970 6304
rect 10331 6283 10368 6293
rect 10331 6265 10341 6283
rect 10359 6265 10368 6283
rect 12346 6279 12377 6300
rect 12767 6279 12803 6300
rect 12189 6278 12226 6279
rect 10784 6273 10821 6275
rect 10784 6272 11432 6273
rect 10152 6256 10189 6257
rect 10331 6256 10368 6265
rect 10783 6266 11432 6272
rect 9575 6235 9611 6256
rect 10001 6235 10032 6256
rect 10783 6248 10793 6266
rect 10811 6252 11432 6266
rect 10811 6248 10821 6252
rect 11262 6251 11432 6252
rect 10783 6238 10821 6248
rect 9408 6231 9508 6235
rect 9408 6227 9470 6231
rect 9408 6201 9415 6227
rect 9441 6205 9470 6227
rect 9496 6205 9508 6231
rect 9441 6201 9508 6205
rect 9408 6198 9508 6201
rect 9576 6198 9611 6235
rect 9673 6232 10032 6235
rect 9673 6227 9895 6232
rect 9673 6203 9686 6227
rect 9710 6208 9895 6227
rect 9919 6208 10032 6232
rect 9710 6203 10032 6208
rect 9673 6199 10032 6203
rect 10099 6227 10248 6235
rect 10099 6207 10110 6227
rect 10130 6207 10248 6227
rect 10099 6200 10248 6207
rect 10099 6199 10140 6200
rect 9423 6146 9460 6147
rect 9519 6146 9556 6147
rect 9575 6146 9611 6198
rect 9630 6146 9667 6147
rect 9323 6137 9461 6146
rect 8259 6119 8290 6122
rect 8259 6093 8266 6119
rect 8285 6093 8290 6119
rect 8259 5699 8290 6093
rect 8311 6118 8479 6119
rect 8311 6115 8755 6118
rect 8311 6096 8686 6115
rect 8706 6096 8755 6115
rect 9323 6117 9432 6137
rect 9452 6117 9461 6137
rect 8311 6092 8755 6096
rect 8311 6090 8479 6092
rect 8311 5912 8338 6090
rect 8378 6052 8442 6064
rect 8718 6060 8755 6092
rect 8926 6091 9175 6113
rect 9323 6110 9461 6117
rect 9519 6137 9667 6146
rect 9519 6117 9528 6137
rect 9548 6117 9638 6137
rect 9658 6117 9667 6137
rect 9323 6108 9419 6110
rect 9519 6107 9667 6117
rect 9726 6137 9763 6147
rect 9838 6146 9875 6147
rect 9819 6144 9875 6146
rect 9726 6117 9734 6137
rect 9754 6117 9763 6137
rect 9575 6106 9611 6107
rect 8926 6060 8963 6091
rect 9139 6089 9175 6091
rect 9139 6060 9176 6089
rect 8378 6051 8413 6052
rect 8355 6046 8413 6051
rect 8355 6026 8358 6046
rect 8378 6032 8413 6046
rect 8433 6032 8442 6052
rect 8378 6024 8442 6032
rect 8404 6023 8442 6024
rect 8405 6022 8442 6023
rect 8508 6056 8544 6057
rect 8616 6056 8652 6057
rect 8508 6048 8652 6056
rect 8508 6028 8516 6048
rect 8536 6047 8624 6048
rect 8536 6028 8569 6047
rect 8508 6027 8569 6028
rect 8593 6028 8624 6047
rect 8644 6028 8652 6048
rect 8593 6027 8652 6028
rect 8508 6022 8652 6027
rect 8718 6052 8756 6060
rect 8824 6056 8860 6057
rect 8718 6032 8727 6052
rect 8747 6032 8756 6052
rect 8718 6023 8756 6032
rect 8775 6049 8860 6056
rect 8775 6029 8782 6049
rect 8803 6048 8860 6049
rect 8803 6029 8832 6048
rect 8775 6028 8832 6029
rect 8852 6028 8860 6048
rect 8718 6022 8755 6023
rect 8775 6022 8860 6028
rect 8926 6052 8964 6060
rect 9037 6056 9073 6057
rect 8926 6032 8935 6052
rect 8955 6032 8964 6052
rect 8926 6023 8964 6032
rect 8988 6048 9073 6056
rect 8988 6028 9045 6048
rect 9065 6028 9073 6048
rect 8926 6022 8963 6023
rect 8988 6022 9073 6028
rect 9139 6052 9177 6060
rect 9139 6032 9148 6052
rect 9168 6032 9177 6052
rect 9423 6047 9460 6048
rect 9726 6047 9763 6117
rect 9788 6137 9875 6144
rect 9788 6134 9846 6137
rect 9788 6114 9793 6134
rect 9814 6117 9846 6134
rect 9866 6117 9875 6137
rect 9814 6114 9875 6117
rect 9788 6107 9875 6114
rect 9934 6137 9971 6147
rect 9934 6117 9942 6137
rect 9962 6117 9971 6137
rect 9788 6106 9819 6107
rect 9422 6046 9763 6047
rect 9139 6023 9177 6032
rect 9347 6041 9763 6046
rect 9139 6022 9176 6023
rect 8562 6001 8598 6022
rect 8988 6001 9019 6022
rect 9347 6021 9350 6041
rect 9370 6021 9763 6041
rect 9934 6046 9971 6117
rect 10001 6146 10032 6199
rect 10334 6184 10371 6194
rect 10334 6166 10343 6184
rect 10361 6166 10371 6184
rect 10334 6157 10371 6166
rect 10783 6160 10818 6238
rect 11395 6228 11432 6251
rect 12188 6269 12226 6278
rect 12188 6249 12197 6269
rect 12217 6249 12226 6269
rect 12188 6241 12226 6249
rect 12292 6273 12377 6279
rect 12402 6278 12439 6279
rect 12292 6253 12300 6273
rect 12320 6253 12377 6273
rect 12292 6245 12377 6253
rect 12401 6269 12439 6278
rect 12401 6249 12410 6269
rect 12430 6249 12439 6269
rect 12292 6244 12328 6245
rect 12401 6241 12439 6249
rect 12505 6273 12590 6279
rect 12610 6278 12647 6279
rect 12505 6253 12513 6273
rect 12533 6272 12590 6273
rect 12533 6253 12562 6272
rect 12505 6252 12562 6253
rect 12583 6252 12590 6272
rect 12505 6245 12590 6252
rect 12609 6269 12647 6278
rect 12609 6249 12618 6269
rect 12638 6249 12647 6269
rect 12505 6244 12541 6245
rect 12609 6241 12647 6249
rect 12713 6277 12857 6279
rect 12713 6273 12771 6277
rect 12713 6253 12721 6273
rect 12741 6253 12771 6273
rect 12713 6251 12771 6253
rect 12796 6273 12857 6277
rect 12796 6253 12829 6273
rect 12849 6253 12857 6273
rect 12796 6251 12857 6253
rect 12713 6245 12857 6251
rect 12713 6244 12749 6245
rect 12821 6244 12857 6245
rect 12923 6278 12960 6279
rect 12923 6277 12961 6278
rect 12923 6269 12987 6277
rect 12923 6249 12932 6269
rect 12952 6255 12987 6269
rect 13007 6255 13010 6275
rect 12952 6250 13010 6255
rect 12952 6249 12987 6250
rect 10051 6146 10088 6147
rect 10001 6137 10088 6146
rect 10001 6117 10059 6137
rect 10079 6117 10088 6137
rect 10001 6107 10088 6117
rect 10147 6137 10184 6147
rect 10147 6117 10155 6137
rect 10175 6117 10184 6137
rect 10001 6106 10032 6107
rect 10147 6046 10184 6117
rect 10339 6092 10370 6157
rect 10779 6151 10818 6160
rect 10779 6133 10789 6151
rect 10807 6133 10818 6151
rect 10779 6127 10818 6133
rect 10974 6203 11224 6227
rect 10974 6132 11011 6203
rect 11126 6142 11157 6143
rect 10779 6123 10816 6127
rect 10974 6112 10983 6132
rect 11003 6112 11011 6132
rect 10974 6102 11011 6112
rect 11070 6132 11157 6142
rect 11070 6112 11079 6132
rect 11099 6112 11157 6132
rect 11070 6103 11157 6112
rect 11070 6102 11107 6103
rect 10338 6082 10375 6092
rect 10338 6080 10348 6082
rect 10272 6078 10348 6080
rect 9934 6022 10184 6046
rect 10269 6064 10348 6078
rect 10366 6064 10375 6082
rect 10269 6061 10375 6064
rect 9741 6002 9762 6021
rect 10269 6002 10295 6061
rect 10338 6055 10375 6061
rect 10782 6052 10819 6061
rect 8395 5997 8495 6001
rect 8395 5993 8457 5997
rect 8395 5967 8402 5993
rect 8428 5971 8457 5993
rect 8483 5971 8495 5997
rect 8428 5967 8495 5971
rect 8395 5964 8495 5967
rect 8563 5964 8598 6001
rect 8660 5998 9019 6001
rect 8660 5993 8882 5998
rect 8660 5969 8673 5993
rect 8697 5974 8882 5993
rect 8906 5974 9019 5998
rect 8697 5969 9019 5974
rect 8660 5965 9019 5969
rect 9086 5993 9235 6001
rect 9086 5973 9097 5993
rect 9117 5973 9235 5993
rect 9741 5984 10295 6002
rect 10780 6034 10791 6052
rect 10809 6034 10819 6052
rect 11126 6050 11157 6103
rect 11187 6132 11224 6203
rect 11395 6208 11788 6228
rect 11808 6208 11811 6228
rect 12189 6212 12226 6241
rect 11395 6203 11811 6208
rect 12190 6210 12226 6212
rect 12402 6210 12439 6241
rect 11395 6202 11736 6203
rect 11339 6142 11370 6143
rect 11187 6112 11196 6132
rect 11216 6112 11224 6132
rect 11187 6102 11224 6112
rect 11283 6135 11370 6142
rect 11283 6132 11344 6135
rect 11283 6112 11292 6132
rect 11312 6115 11344 6132
rect 11365 6115 11370 6135
rect 11312 6112 11370 6115
rect 11283 6105 11370 6112
rect 11395 6132 11432 6202
rect 11698 6201 11735 6202
rect 12190 6188 12439 6210
rect 12610 6209 12647 6241
rect 12923 6237 12987 6249
rect 13027 6211 13054 6389
rect 12886 6209 13054 6211
rect 12610 6183 13054 6209
rect 12886 6182 13054 6183
rect 11547 6142 11583 6143
rect 11395 6112 11404 6132
rect 11424 6112 11432 6132
rect 11283 6103 11339 6105
rect 11283 6102 11320 6103
rect 11395 6102 11432 6112
rect 11491 6132 11639 6142
rect 11739 6139 11835 6141
rect 11491 6112 11500 6132
rect 11520 6112 11610 6132
rect 11630 6112 11639 6132
rect 11491 6103 11639 6112
rect 11697 6132 11835 6139
rect 11697 6112 11706 6132
rect 11726 6112 11835 6132
rect 11697 6103 11835 6112
rect 11491 6102 11528 6103
rect 11547 6051 11583 6103
rect 11602 6102 11639 6103
rect 11698 6102 11735 6103
rect 11018 6049 11059 6050
rect 10341 5991 10378 5993
rect 10269 5983 10295 5984
rect 10338 5983 10378 5991
rect 9086 5966 9235 5973
rect 10338 5971 10350 5983
rect 10329 5966 10350 5971
rect 9086 5965 9127 5966
rect 9745 5965 10350 5966
rect 10368 5965 10378 5983
rect 8410 5912 8447 5913
rect 8506 5912 8543 5913
rect 8562 5912 8598 5964
rect 8617 5912 8654 5913
rect 8310 5903 8448 5912
rect 8310 5883 8419 5903
rect 8439 5883 8448 5903
rect 8310 5876 8448 5883
rect 8506 5903 8654 5912
rect 8506 5883 8515 5903
rect 8535 5883 8625 5903
rect 8645 5883 8654 5903
rect 8310 5874 8406 5876
rect 8506 5873 8654 5883
rect 8713 5903 8750 5913
rect 8825 5912 8862 5913
rect 8806 5910 8862 5912
rect 8713 5883 8721 5903
rect 8741 5883 8750 5903
rect 8562 5872 8598 5873
rect 8410 5813 8447 5814
rect 8713 5813 8750 5883
rect 8775 5903 8862 5910
rect 8775 5900 8833 5903
rect 8775 5880 8780 5900
rect 8801 5883 8833 5900
rect 8853 5883 8862 5903
rect 8801 5880 8862 5883
rect 8775 5873 8862 5880
rect 8921 5903 8958 5913
rect 8921 5883 8929 5903
rect 8949 5883 8958 5903
rect 8775 5872 8806 5873
rect 8409 5812 8750 5813
rect 8334 5807 8750 5812
rect 8334 5787 8337 5807
rect 8357 5787 8750 5807
rect 8921 5812 8958 5883
rect 8988 5912 9019 5965
rect 9745 5956 10378 5965
rect 9745 5949 10377 5956
rect 9745 5947 9807 5949
rect 9323 5937 9491 5938
rect 9745 5937 9767 5947
rect 9038 5912 9075 5913
rect 8988 5903 9075 5912
rect 8988 5883 9046 5903
rect 9066 5883 9075 5903
rect 8988 5873 9075 5883
rect 9134 5903 9171 5913
rect 9134 5883 9142 5903
rect 9162 5883 9171 5903
rect 8988 5872 9019 5873
rect 9134 5812 9171 5883
rect 8921 5788 9171 5812
rect 9323 5911 9767 5937
rect 9323 5909 9491 5911
rect 9323 5731 9350 5909
rect 9390 5871 9454 5883
rect 9730 5879 9767 5911
rect 9938 5910 10187 5932
rect 9938 5879 9975 5910
rect 10151 5908 10187 5910
rect 10151 5879 10188 5908
rect 9390 5870 9425 5871
rect 9367 5865 9425 5870
rect 9367 5845 9370 5865
rect 9390 5851 9425 5865
rect 9445 5851 9454 5871
rect 9390 5843 9454 5851
rect 9416 5842 9454 5843
rect 9417 5841 9454 5842
rect 9520 5875 9556 5876
rect 9628 5875 9664 5876
rect 9520 5867 9664 5875
rect 9520 5847 9528 5867
rect 9548 5847 9577 5867
rect 9520 5846 9577 5847
rect 9599 5847 9636 5867
rect 9656 5847 9664 5867
rect 9599 5846 9664 5847
rect 9520 5841 9664 5846
rect 9730 5871 9768 5879
rect 9836 5875 9872 5876
rect 9730 5851 9739 5871
rect 9759 5851 9768 5871
rect 9730 5842 9768 5851
rect 9787 5868 9872 5875
rect 9787 5848 9794 5868
rect 9815 5867 9872 5868
rect 9815 5848 9844 5867
rect 9787 5847 9844 5848
rect 9864 5847 9872 5867
rect 9730 5841 9767 5842
rect 9787 5841 9872 5847
rect 9938 5871 9976 5879
rect 10049 5875 10085 5876
rect 9938 5851 9947 5871
rect 9967 5851 9976 5871
rect 9938 5842 9976 5851
rect 10000 5867 10085 5875
rect 10000 5847 10057 5867
rect 10077 5847 10085 5867
rect 9938 5841 9975 5842
rect 10000 5841 10085 5847
rect 10151 5871 10189 5879
rect 10151 5851 10160 5871
rect 10180 5851 10189 5871
rect 10151 5842 10189 5851
rect 10151 5841 10188 5842
rect 9574 5820 9610 5841
rect 10000 5820 10031 5841
rect 9407 5816 9507 5820
rect 9407 5812 9469 5816
rect 9407 5786 9414 5812
rect 9440 5790 9469 5812
rect 9495 5790 9507 5816
rect 9440 5786 9507 5790
rect 9407 5783 9507 5786
rect 9575 5783 9610 5820
rect 9672 5817 10031 5820
rect 9672 5812 9894 5817
rect 9672 5788 9685 5812
rect 9709 5793 9894 5812
rect 9918 5793 10031 5817
rect 9709 5788 10031 5793
rect 9672 5784 10031 5788
rect 10098 5812 10247 5820
rect 10098 5792 10109 5812
rect 10129 5792 10247 5812
rect 10098 5785 10247 5792
rect 10338 5800 10377 5949
rect 10780 5885 10819 6034
rect 10910 6042 11059 6049
rect 10910 6022 11028 6042
rect 11048 6022 11059 6042
rect 10910 6014 11059 6022
rect 11126 6046 11485 6050
rect 11126 6041 11448 6046
rect 11126 6017 11239 6041
rect 11263 6022 11448 6041
rect 11472 6022 11485 6046
rect 11263 6017 11485 6022
rect 11126 6014 11485 6017
rect 11547 6014 11582 6051
rect 11650 6048 11750 6051
rect 11650 6044 11717 6048
rect 11650 6018 11662 6044
rect 11688 6022 11717 6044
rect 11743 6022 11750 6048
rect 11688 6018 11750 6022
rect 11650 6014 11750 6018
rect 11126 5993 11157 6014
rect 11547 5993 11583 6014
rect 10969 5992 11006 5993
rect 10968 5983 11006 5992
rect 10968 5963 10977 5983
rect 10997 5963 11006 5983
rect 10968 5955 11006 5963
rect 11072 5987 11157 5993
rect 11182 5992 11219 5993
rect 11072 5967 11080 5987
rect 11100 5967 11157 5987
rect 11072 5959 11157 5967
rect 11181 5983 11219 5992
rect 11181 5963 11190 5983
rect 11210 5963 11219 5983
rect 11072 5958 11108 5959
rect 11181 5955 11219 5963
rect 11285 5987 11370 5993
rect 11390 5992 11427 5993
rect 11285 5967 11293 5987
rect 11313 5986 11370 5987
rect 11313 5967 11342 5986
rect 11285 5966 11342 5967
rect 11363 5966 11370 5986
rect 11285 5959 11370 5966
rect 11389 5983 11427 5992
rect 11389 5963 11398 5983
rect 11418 5963 11427 5983
rect 11285 5958 11321 5959
rect 11389 5955 11427 5963
rect 11493 5988 11637 5993
rect 11493 5987 11558 5988
rect 11493 5967 11501 5987
rect 11521 5967 11558 5987
rect 11580 5987 11637 5988
rect 11580 5967 11609 5987
rect 11629 5967 11637 5987
rect 11493 5959 11637 5967
rect 11493 5958 11529 5959
rect 11601 5958 11637 5959
rect 11703 5992 11740 5993
rect 11703 5991 11741 5992
rect 11703 5983 11767 5991
rect 11703 5963 11712 5983
rect 11732 5969 11767 5983
rect 11787 5969 11790 5989
rect 11732 5964 11790 5969
rect 11732 5963 11767 5964
rect 10969 5926 11006 5955
rect 10970 5924 11006 5926
rect 11182 5924 11219 5955
rect 10970 5902 11219 5924
rect 11390 5923 11427 5955
rect 11703 5951 11767 5963
rect 11807 5925 11834 6103
rect 11666 5923 11834 5925
rect 11390 5897 11834 5923
rect 11986 6022 12236 6046
rect 11986 5951 12023 6022
rect 12138 5961 12169 5962
rect 11986 5931 11995 5951
rect 12015 5931 12023 5951
rect 11986 5921 12023 5931
rect 12082 5951 12169 5961
rect 12082 5931 12091 5951
rect 12111 5931 12169 5951
rect 12082 5922 12169 5931
rect 12082 5921 12119 5922
rect 11390 5887 11412 5897
rect 11666 5896 11834 5897
rect 11350 5885 11412 5887
rect 10780 5878 11412 5885
rect 10779 5869 11412 5878
rect 12138 5869 12169 5922
rect 12199 5951 12236 6022
rect 12407 6027 12800 6047
rect 12820 6027 12823 6047
rect 12407 6022 12823 6027
rect 12407 6021 12748 6022
rect 12351 5961 12382 5962
rect 12199 5931 12208 5951
rect 12228 5931 12236 5951
rect 12199 5921 12236 5931
rect 12295 5954 12382 5961
rect 12295 5951 12356 5954
rect 12295 5931 12304 5951
rect 12324 5934 12356 5951
rect 12377 5934 12382 5954
rect 12324 5931 12382 5934
rect 12295 5924 12382 5931
rect 12407 5951 12444 6021
rect 12710 6020 12747 6021
rect 12559 5961 12595 5962
rect 12407 5931 12416 5951
rect 12436 5931 12444 5951
rect 12295 5922 12351 5924
rect 12295 5921 12332 5922
rect 12407 5921 12444 5931
rect 12503 5951 12651 5961
rect 12751 5958 12847 5960
rect 12503 5931 12512 5951
rect 12532 5931 12622 5951
rect 12642 5931 12651 5951
rect 12503 5922 12651 5931
rect 12709 5951 12847 5958
rect 12709 5931 12718 5951
rect 12738 5931 12847 5951
rect 12709 5922 12847 5931
rect 12503 5921 12540 5922
rect 12559 5870 12595 5922
rect 12614 5921 12651 5922
rect 12710 5921 12747 5922
rect 10779 5851 10789 5869
rect 10807 5868 11412 5869
rect 12030 5868 12071 5869
rect 10807 5863 10828 5868
rect 10807 5851 10819 5863
rect 11922 5861 12071 5868
rect 10779 5843 10819 5851
rect 10862 5850 10888 5851
rect 10779 5841 10816 5843
rect 10098 5784 10139 5785
rect 9422 5731 9459 5732
rect 9518 5731 9555 5732
rect 9574 5731 9610 5783
rect 9629 5731 9666 5732
rect 9322 5722 9460 5731
rect 9322 5702 9431 5722
rect 9451 5702 9460 5722
rect 8259 5698 8429 5699
rect 8259 5683 8705 5698
rect 9322 5695 9460 5702
rect 9518 5722 9666 5731
rect 9518 5702 9527 5722
rect 9547 5702 9637 5722
rect 9657 5702 9666 5722
rect 9322 5693 9418 5695
rect 8261 5672 8705 5683
rect 8261 5670 8429 5672
rect 8261 5492 8288 5670
rect 8328 5632 8392 5644
rect 8668 5640 8705 5672
rect 8876 5671 9125 5693
rect 9518 5692 9666 5702
rect 9725 5722 9762 5732
rect 9837 5731 9874 5732
rect 9818 5729 9874 5731
rect 9725 5702 9733 5722
rect 9753 5702 9762 5722
rect 9574 5691 9610 5692
rect 8876 5640 8913 5671
rect 9089 5669 9125 5671
rect 9089 5640 9126 5669
rect 8328 5631 8363 5632
rect 8305 5626 8363 5631
rect 8305 5606 8308 5626
rect 8328 5612 8363 5626
rect 8383 5612 8392 5632
rect 8328 5604 8392 5612
rect 8354 5603 8392 5604
rect 8355 5602 8392 5603
rect 8458 5636 8494 5637
rect 8566 5636 8602 5637
rect 8458 5628 8602 5636
rect 8458 5608 8466 5628
rect 8486 5627 8574 5628
rect 8486 5610 8514 5627
rect 8538 5610 8574 5627
rect 8486 5608 8574 5610
rect 8594 5608 8602 5628
rect 8458 5602 8602 5608
rect 8668 5632 8706 5640
rect 8774 5636 8810 5637
rect 8668 5612 8677 5632
rect 8697 5612 8706 5632
rect 8668 5603 8706 5612
rect 8725 5629 8810 5636
rect 8725 5609 8732 5629
rect 8753 5628 8810 5629
rect 8753 5609 8782 5628
rect 8725 5608 8782 5609
rect 8802 5608 8810 5628
rect 8668 5602 8705 5603
rect 8725 5602 8810 5608
rect 8876 5632 8914 5640
rect 8987 5636 9023 5637
rect 8876 5612 8885 5632
rect 8905 5612 8914 5632
rect 8876 5603 8914 5612
rect 8938 5628 9023 5636
rect 8938 5608 8995 5628
rect 9015 5608 9023 5628
rect 8876 5602 8913 5603
rect 8938 5602 9023 5608
rect 9089 5632 9127 5640
rect 9422 5632 9459 5633
rect 9725 5632 9762 5702
rect 9787 5722 9874 5729
rect 9787 5719 9845 5722
rect 9787 5699 9792 5719
rect 9813 5702 9845 5719
rect 9865 5702 9874 5722
rect 9813 5699 9874 5702
rect 9787 5692 9874 5699
rect 9933 5722 9970 5732
rect 9933 5702 9941 5722
rect 9961 5702 9970 5722
rect 9787 5691 9818 5692
rect 9089 5612 9098 5632
rect 9118 5612 9127 5632
rect 9421 5631 9762 5632
rect 9089 5603 9127 5612
rect 9346 5626 9762 5631
rect 9346 5606 9349 5626
rect 9369 5606 9762 5626
rect 9933 5631 9970 5702
rect 10000 5731 10031 5784
rect 10338 5782 10348 5800
rect 10366 5782 10377 5800
rect 10862 5832 11416 5850
rect 11922 5841 12040 5861
rect 12060 5841 12071 5861
rect 11922 5833 12071 5841
rect 12138 5865 12497 5869
rect 12138 5860 12460 5865
rect 12138 5836 12251 5860
rect 12275 5841 12460 5860
rect 12484 5841 12497 5865
rect 12275 5836 12497 5841
rect 12138 5833 12497 5836
rect 12559 5833 12594 5870
rect 12662 5867 12762 5870
rect 12662 5863 12729 5867
rect 12662 5837 12674 5863
rect 12700 5841 12729 5863
rect 12755 5841 12762 5867
rect 12700 5837 12762 5841
rect 12662 5833 12762 5837
rect 10338 5773 10375 5782
rect 10782 5773 10819 5779
rect 10862 5773 10888 5832
rect 11395 5813 11416 5832
rect 10782 5770 10888 5773
rect 10782 5752 10791 5770
rect 10809 5756 10888 5770
rect 10973 5788 11223 5812
rect 10809 5754 10885 5756
rect 10809 5752 10819 5754
rect 10782 5742 10819 5752
rect 10050 5731 10087 5732
rect 10000 5722 10087 5731
rect 10000 5702 10058 5722
rect 10078 5702 10087 5722
rect 10000 5692 10087 5702
rect 10146 5722 10183 5732
rect 10146 5702 10154 5722
rect 10174 5702 10183 5722
rect 10341 5707 10378 5711
rect 10000 5691 10031 5692
rect 10146 5631 10183 5702
rect 9933 5607 10183 5631
rect 10339 5701 10378 5707
rect 10339 5683 10350 5701
rect 10368 5683 10378 5701
rect 10339 5674 10378 5683
rect 10787 5677 10818 5742
rect 10973 5717 11010 5788
rect 11125 5727 11156 5728
rect 10973 5697 10982 5717
rect 11002 5697 11010 5717
rect 10973 5687 11010 5697
rect 11069 5717 11156 5727
rect 11069 5697 11078 5717
rect 11098 5697 11156 5717
rect 11069 5688 11156 5697
rect 11069 5687 11106 5688
rect 9089 5602 9126 5603
rect 8512 5581 8548 5602
rect 8938 5581 8969 5602
rect 9725 5583 9762 5606
rect 10339 5596 10374 5674
rect 10786 5668 10823 5677
rect 10786 5650 10796 5668
rect 10814 5650 10823 5668
rect 10786 5640 10823 5650
rect 11125 5635 11156 5688
rect 11186 5717 11223 5788
rect 11394 5793 11787 5813
rect 11807 5793 11810 5813
rect 12138 5812 12169 5833
rect 12559 5812 12595 5833
rect 11981 5811 12018 5812
rect 11394 5788 11810 5793
rect 11980 5802 12018 5811
rect 11394 5787 11735 5788
rect 11338 5727 11369 5728
rect 11186 5697 11195 5717
rect 11215 5697 11223 5717
rect 11186 5687 11223 5697
rect 11282 5720 11369 5727
rect 11282 5717 11343 5720
rect 11282 5697 11291 5717
rect 11311 5700 11343 5717
rect 11364 5700 11369 5720
rect 11311 5697 11369 5700
rect 11282 5690 11369 5697
rect 11394 5717 11431 5787
rect 11697 5786 11734 5787
rect 11980 5782 11989 5802
rect 12009 5782 12018 5802
rect 11980 5774 12018 5782
rect 12084 5806 12169 5812
rect 12194 5811 12231 5812
rect 12084 5786 12092 5806
rect 12112 5786 12169 5806
rect 12084 5778 12169 5786
rect 12193 5802 12231 5811
rect 12193 5782 12202 5802
rect 12222 5782 12231 5802
rect 12084 5777 12120 5778
rect 12193 5774 12231 5782
rect 12297 5806 12382 5812
rect 12402 5811 12439 5812
rect 12297 5786 12305 5806
rect 12325 5805 12382 5806
rect 12325 5786 12354 5805
rect 12297 5785 12354 5786
rect 12375 5785 12382 5805
rect 12297 5778 12382 5785
rect 12401 5802 12439 5811
rect 12401 5782 12410 5802
rect 12430 5782 12439 5802
rect 12297 5777 12333 5778
rect 12401 5774 12439 5782
rect 12505 5806 12649 5812
rect 12505 5786 12513 5806
rect 12533 5786 12565 5806
rect 12589 5786 12621 5806
rect 12641 5786 12649 5806
rect 12505 5778 12649 5786
rect 12505 5777 12541 5778
rect 12613 5777 12649 5778
rect 12715 5811 12752 5812
rect 12715 5810 12753 5811
rect 12715 5802 12779 5810
rect 12715 5782 12724 5802
rect 12744 5788 12779 5802
rect 12799 5788 12802 5808
rect 12744 5783 12802 5788
rect 12744 5782 12779 5783
rect 11981 5745 12018 5774
rect 11982 5743 12018 5745
rect 12194 5743 12231 5774
rect 11546 5727 11582 5728
rect 11394 5697 11403 5717
rect 11423 5697 11431 5717
rect 11282 5688 11338 5690
rect 11282 5687 11319 5688
rect 11394 5687 11431 5697
rect 11490 5717 11638 5727
rect 11738 5724 11834 5726
rect 11490 5697 11499 5717
rect 11519 5697 11609 5717
rect 11629 5697 11638 5717
rect 11490 5688 11638 5697
rect 11696 5717 11834 5724
rect 11982 5721 12231 5743
rect 12402 5742 12439 5774
rect 12715 5770 12779 5782
rect 12819 5744 12846 5922
rect 12678 5742 12846 5744
rect 12402 5738 12846 5742
rect 11696 5697 11705 5717
rect 11725 5697 11834 5717
rect 12402 5719 12451 5738
rect 12471 5719 12846 5738
rect 12402 5716 12846 5719
rect 12678 5715 12846 5716
rect 11696 5688 11834 5697
rect 11490 5687 11527 5688
rect 11546 5636 11582 5688
rect 11601 5687 11638 5688
rect 11697 5687 11734 5688
rect 11017 5634 11058 5635
rect 10909 5627 11058 5634
rect 10909 5607 11027 5627
rect 11047 5607 11058 5627
rect 10909 5599 11058 5607
rect 11125 5631 11484 5635
rect 11125 5626 11447 5631
rect 11125 5602 11238 5626
rect 11262 5607 11447 5626
rect 11471 5607 11484 5631
rect 11262 5602 11484 5607
rect 11125 5599 11484 5602
rect 11546 5599 11581 5636
rect 11649 5633 11749 5636
rect 11649 5629 11716 5633
rect 11649 5603 11661 5629
rect 11687 5607 11716 5629
rect 11742 5607 11749 5633
rect 11687 5603 11749 5607
rect 11649 5599 11749 5603
rect 10336 5586 10374 5596
rect 9725 5582 9895 5583
rect 10336 5582 10346 5586
rect 8345 5577 8445 5581
rect 8345 5573 8407 5577
rect 8345 5547 8352 5573
rect 8378 5551 8407 5573
rect 8433 5551 8445 5577
rect 8378 5547 8445 5551
rect 8345 5544 8445 5547
rect 8513 5544 8548 5581
rect 8610 5578 8969 5581
rect 8610 5573 8832 5578
rect 8610 5549 8623 5573
rect 8647 5554 8832 5573
rect 8856 5554 8969 5578
rect 8647 5549 8969 5554
rect 8610 5545 8969 5549
rect 9036 5573 9185 5581
rect 9036 5553 9047 5573
rect 9067 5553 9185 5573
rect 9725 5568 10346 5582
rect 10364 5568 10374 5586
rect 11125 5578 11156 5599
rect 11546 5578 11582 5599
rect 9725 5562 10374 5568
rect 10789 5569 10826 5578
rect 10968 5577 11005 5578
rect 9725 5561 10373 5562
rect 10336 5559 10373 5561
rect 9036 5546 9185 5553
rect 10789 5551 10798 5569
rect 10816 5551 10826 5569
rect 9036 5545 9077 5546
rect 8360 5492 8397 5493
rect 8456 5492 8493 5493
rect 8512 5492 8548 5544
rect 8567 5492 8604 5493
rect 8260 5483 8398 5492
rect 8260 5463 8369 5483
rect 8389 5463 8398 5483
rect 8260 5456 8398 5463
rect 8456 5483 8604 5492
rect 8456 5463 8465 5483
rect 8485 5463 8575 5483
rect 8595 5463 8604 5483
rect 8260 5454 8356 5456
rect 8456 5453 8604 5463
rect 8663 5483 8700 5493
rect 8775 5492 8812 5493
rect 8756 5490 8812 5492
rect 8663 5463 8671 5483
rect 8691 5463 8700 5483
rect 8512 5452 8548 5453
rect 8360 5393 8397 5394
rect 8663 5393 8700 5463
rect 8725 5483 8812 5490
rect 8725 5480 8783 5483
rect 8725 5460 8730 5480
rect 8751 5463 8783 5480
rect 8803 5463 8812 5483
rect 8751 5460 8812 5463
rect 8725 5453 8812 5460
rect 8871 5483 8908 5493
rect 8871 5463 8879 5483
rect 8899 5463 8908 5483
rect 8725 5452 8756 5453
rect 8359 5392 8700 5393
rect 8284 5387 8700 5392
rect 8284 5367 8287 5387
rect 8307 5367 8700 5387
rect 8871 5392 8908 5463
rect 8938 5492 8969 5545
rect 10789 5541 10826 5551
rect 10790 5506 10826 5541
rect 10967 5568 11005 5577
rect 10967 5548 10976 5568
rect 10996 5548 11005 5568
rect 10967 5540 11005 5548
rect 11071 5572 11156 5578
rect 11181 5577 11218 5578
rect 11071 5552 11079 5572
rect 11099 5552 11156 5572
rect 11071 5544 11156 5552
rect 11180 5568 11218 5577
rect 11180 5548 11189 5568
rect 11209 5548 11218 5568
rect 11071 5543 11107 5544
rect 11180 5540 11218 5548
rect 11284 5572 11369 5578
rect 11389 5577 11426 5578
rect 11284 5552 11292 5572
rect 11312 5571 11369 5572
rect 11312 5552 11341 5571
rect 11284 5551 11341 5552
rect 11362 5551 11369 5571
rect 11284 5544 11369 5551
rect 11388 5568 11426 5577
rect 11388 5548 11397 5568
rect 11417 5548 11426 5568
rect 11284 5543 11320 5544
rect 11388 5540 11426 5548
rect 11492 5572 11636 5578
rect 11492 5552 11500 5572
rect 11520 5571 11608 5572
rect 11520 5552 11548 5571
rect 11492 5550 11548 5552
rect 11570 5552 11608 5571
rect 11628 5552 11636 5572
rect 11570 5550 11636 5552
rect 11492 5544 11636 5550
rect 11492 5543 11528 5544
rect 11600 5543 11636 5544
rect 11702 5577 11739 5578
rect 11702 5576 11740 5577
rect 11702 5568 11766 5576
rect 11702 5548 11711 5568
rect 11731 5554 11766 5568
rect 11786 5554 11789 5574
rect 11731 5549 11789 5554
rect 11731 5548 11766 5549
rect 10968 5511 11005 5540
rect 8988 5492 9025 5493
rect 8938 5483 9025 5492
rect 8938 5463 8996 5483
rect 9016 5463 9025 5483
rect 8938 5453 9025 5463
rect 9084 5483 9121 5493
rect 9084 5463 9092 5483
rect 9112 5463 9121 5483
rect 8938 5452 8969 5453
rect 9084 5392 9121 5463
rect 10339 5487 10376 5497
rect 10339 5469 10348 5487
rect 10366 5469 10376 5487
rect 10339 5460 10376 5469
rect 10788 5465 10826 5506
rect 10969 5509 11005 5511
rect 11181 5509 11218 5540
rect 10969 5487 11218 5509
rect 11389 5508 11426 5540
rect 11702 5536 11766 5548
rect 11806 5510 11833 5688
rect 11665 5508 11833 5510
rect 11389 5482 11833 5508
rect 11390 5465 11414 5482
rect 11665 5481 11833 5482
rect 10339 5436 10374 5460
rect 10337 5412 10374 5436
rect 10336 5406 10374 5412
rect 8871 5368 9121 5392
rect 9747 5388 10374 5406
rect 10788 5447 11415 5465
rect 12041 5461 12291 5485
rect 10788 5441 10826 5447
rect 10788 5417 10825 5441
rect 10788 5393 10823 5417
rect 9329 5371 9497 5372
rect 9748 5371 9772 5388
rect 9329 5345 9773 5371
rect 9329 5343 9497 5345
rect 9329 5165 9356 5343
rect 9396 5305 9460 5317
rect 9736 5313 9773 5345
rect 9944 5344 10193 5366
rect 9944 5313 9981 5344
rect 10157 5342 10193 5344
rect 10336 5347 10374 5388
rect 10786 5384 10823 5393
rect 10786 5366 10796 5384
rect 10814 5366 10823 5384
rect 10786 5356 10823 5366
rect 12041 5390 12078 5461
rect 12193 5400 12224 5401
rect 12041 5370 12050 5390
rect 12070 5370 12078 5390
rect 12041 5360 12078 5370
rect 12137 5390 12224 5400
rect 12137 5370 12146 5390
rect 12166 5370 12224 5390
rect 12137 5361 12224 5370
rect 12137 5360 12174 5361
rect 10157 5313 10194 5342
rect 9396 5304 9431 5305
rect 9373 5299 9431 5304
rect 9373 5279 9376 5299
rect 9396 5285 9431 5299
rect 9451 5285 9460 5305
rect 9396 5277 9460 5285
rect 9422 5276 9460 5277
rect 9423 5275 9460 5276
rect 9526 5309 9562 5310
rect 9634 5309 9670 5310
rect 9526 5303 9670 5309
rect 9526 5301 9592 5303
rect 9526 5281 9534 5301
rect 9554 5282 9592 5301
rect 9614 5301 9670 5303
rect 9614 5282 9642 5301
rect 9554 5281 9642 5282
rect 9662 5281 9670 5301
rect 9526 5275 9670 5281
rect 9736 5305 9774 5313
rect 9842 5309 9878 5310
rect 9736 5285 9745 5305
rect 9765 5285 9774 5305
rect 9736 5276 9774 5285
rect 9793 5302 9878 5309
rect 9793 5282 9800 5302
rect 9821 5301 9878 5302
rect 9821 5282 9850 5301
rect 9793 5281 9850 5282
rect 9870 5281 9878 5301
rect 9736 5275 9773 5276
rect 9793 5275 9878 5281
rect 9944 5305 9982 5313
rect 10055 5309 10091 5310
rect 9944 5285 9953 5305
rect 9973 5285 9982 5305
rect 9944 5276 9982 5285
rect 10006 5301 10091 5309
rect 10006 5281 10063 5301
rect 10083 5281 10091 5301
rect 9944 5275 9981 5276
rect 10006 5275 10091 5281
rect 10157 5305 10195 5313
rect 10157 5285 10166 5305
rect 10186 5285 10195 5305
rect 10157 5276 10195 5285
rect 10336 5312 10372 5347
rect 10336 5302 10373 5312
rect 12193 5308 12224 5361
rect 12254 5390 12291 5461
rect 12462 5466 12855 5486
rect 12875 5466 12878 5486
rect 12462 5461 12878 5466
rect 12462 5460 12803 5461
rect 12406 5400 12437 5401
rect 12254 5370 12263 5390
rect 12283 5370 12291 5390
rect 12254 5360 12291 5370
rect 12350 5393 12437 5400
rect 12350 5390 12411 5393
rect 12350 5370 12359 5390
rect 12379 5373 12411 5390
rect 12432 5373 12437 5393
rect 12379 5370 12437 5373
rect 12350 5363 12437 5370
rect 12462 5390 12499 5460
rect 12765 5459 12802 5460
rect 12614 5400 12650 5401
rect 12462 5370 12471 5390
rect 12491 5370 12499 5390
rect 12350 5361 12406 5363
rect 12350 5360 12387 5361
rect 12462 5360 12499 5370
rect 12558 5390 12706 5400
rect 12806 5397 12902 5399
rect 12558 5370 12567 5390
rect 12587 5370 12677 5390
rect 12697 5370 12706 5390
rect 12558 5361 12706 5370
rect 12764 5390 12902 5397
rect 12764 5370 12773 5390
rect 12793 5370 12902 5390
rect 12764 5361 12902 5370
rect 12558 5360 12595 5361
rect 12614 5309 12650 5361
rect 12669 5360 12706 5361
rect 12765 5360 12802 5361
rect 12085 5307 12126 5308
rect 10336 5284 10346 5302
rect 10364 5284 10373 5302
rect 11977 5300 12126 5307
rect 10789 5292 10826 5294
rect 10789 5291 11437 5292
rect 10157 5275 10194 5276
rect 10336 5275 10373 5284
rect 10788 5285 11437 5291
rect 9580 5254 9616 5275
rect 10006 5254 10037 5275
rect 10788 5267 10798 5285
rect 10816 5271 11437 5285
rect 11977 5280 12095 5300
rect 12115 5280 12126 5300
rect 11977 5272 12126 5280
rect 12193 5304 12552 5308
rect 12193 5299 12515 5304
rect 12193 5275 12306 5299
rect 12330 5280 12515 5299
rect 12539 5280 12552 5304
rect 12330 5275 12552 5280
rect 12193 5272 12552 5275
rect 12614 5272 12649 5309
rect 12717 5306 12817 5309
rect 12717 5302 12784 5306
rect 12717 5276 12729 5302
rect 12755 5280 12784 5302
rect 12810 5280 12817 5306
rect 12755 5276 12817 5280
rect 12717 5272 12817 5276
rect 10816 5267 10826 5271
rect 11267 5270 11437 5271
rect 10788 5257 10826 5267
rect 9413 5250 9513 5254
rect 9413 5246 9475 5250
rect 9413 5220 9420 5246
rect 9446 5224 9475 5246
rect 9501 5224 9513 5250
rect 9446 5220 9513 5224
rect 9413 5217 9513 5220
rect 9581 5217 9616 5254
rect 9678 5251 10037 5254
rect 9678 5246 9900 5251
rect 9678 5222 9691 5246
rect 9715 5227 9900 5246
rect 9924 5227 10037 5251
rect 9715 5222 10037 5227
rect 9678 5218 10037 5222
rect 10104 5246 10253 5254
rect 10104 5226 10115 5246
rect 10135 5226 10253 5246
rect 10104 5219 10253 5226
rect 10104 5218 10145 5219
rect 9428 5165 9465 5166
rect 9524 5165 9561 5166
rect 9580 5165 9616 5217
rect 9635 5165 9672 5166
rect 9328 5156 9466 5165
rect 8316 5137 8484 5138
rect 8316 5134 8760 5137
rect 8316 5115 8691 5134
rect 8711 5115 8760 5134
rect 9328 5136 9437 5156
rect 9457 5136 9466 5156
rect 8316 5111 8760 5115
rect 8316 5109 8484 5111
rect 8316 4931 8343 5109
rect 8383 5071 8447 5083
rect 8723 5079 8760 5111
rect 8931 5110 9180 5132
rect 9328 5129 9466 5136
rect 9524 5156 9672 5165
rect 9524 5136 9533 5156
rect 9553 5136 9643 5156
rect 9663 5136 9672 5156
rect 9328 5127 9424 5129
rect 9524 5126 9672 5136
rect 9731 5156 9768 5166
rect 9843 5165 9880 5166
rect 9824 5163 9880 5165
rect 9731 5136 9739 5156
rect 9759 5136 9768 5156
rect 9580 5125 9616 5126
rect 8931 5079 8968 5110
rect 9144 5108 9180 5110
rect 9144 5079 9181 5108
rect 8383 5070 8418 5071
rect 8360 5065 8418 5070
rect 8360 5045 8363 5065
rect 8383 5051 8418 5065
rect 8438 5051 8447 5071
rect 8383 5043 8447 5051
rect 8409 5042 8447 5043
rect 8410 5041 8447 5042
rect 8513 5075 8549 5076
rect 8621 5075 8657 5076
rect 8513 5067 8657 5075
rect 8513 5047 8521 5067
rect 8541 5047 8573 5067
rect 8597 5047 8629 5067
rect 8649 5047 8657 5067
rect 8513 5041 8657 5047
rect 8723 5071 8761 5079
rect 8829 5075 8865 5076
rect 8723 5051 8732 5071
rect 8752 5051 8761 5071
rect 8723 5042 8761 5051
rect 8780 5068 8865 5075
rect 8780 5048 8787 5068
rect 8808 5067 8865 5068
rect 8808 5048 8837 5067
rect 8780 5047 8837 5048
rect 8857 5047 8865 5067
rect 8723 5041 8760 5042
rect 8780 5041 8865 5047
rect 8931 5071 8969 5079
rect 9042 5075 9078 5076
rect 8931 5051 8940 5071
rect 8960 5051 8969 5071
rect 8931 5042 8969 5051
rect 8993 5067 9078 5075
rect 8993 5047 9050 5067
rect 9070 5047 9078 5067
rect 8931 5041 8968 5042
rect 8993 5041 9078 5047
rect 9144 5071 9182 5079
rect 9144 5051 9153 5071
rect 9173 5051 9182 5071
rect 9428 5066 9465 5067
rect 9731 5066 9768 5136
rect 9793 5156 9880 5163
rect 9793 5153 9851 5156
rect 9793 5133 9798 5153
rect 9819 5136 9851 5153
rect 9871 5136 9880 5156
rect 9819 5133 9880 5136
rect 9793 5126 9880 5133
rect 9939 5156 9976 5166
rect 9939 5136 9947 5156
rect 9967 5136 9976 5156
rect 9793 5125 9824 5126
rect 9427 5065 9768 5066
rect 9144 5042 9182 5051
rect 9352 5060 9768 5065
rect 9144 5041 9181 5042
rect 8567 5020 8603 5041
rect 8993 5020 9024 5041
rect 9352 5040 9355 5060
rect 9375 5040 9768 5060
rect 9939 5065 9976 5136
rect 10006 5165 10037 5218
rect 10339 5203 10376 5213
rect 10339 5185 10348 5203
rect 10366 5185 10376 5203
rect 10339 5176 10376 5185
rect 10788 5179 10823 5257
rect 11400 5247 11437 5270
rect 12193 5251 12224 5272
rect 12614 5251 12650 5272
rect 12036 5250 12073 5251
rect 10056 5165 10093 5166
rect 10006 5156 10093 5165
rect 10006 5136 10064 5156
rect 10084 5136 10093 5156
rect 10006 5126 10093 5136
rect 10152 5156 10189 5166
rect 10152 5136 10160 5156
rect 10180 5136 10189 5156
rect 10006 5125 10037 5126
rect 10152 5065 10189 5136
rect 10344 5111 10375 5176
rect 10784 5170 10823 5179
rect 10784 5152 10794 5170
rect 10812 5152 10823 5170
rect 10784 5146 10823 5152
rect 10979 5222 11229 5246
rect 10979 5151 11016 5222
rect 11131 5161 11162 5162
rect 10784 5142 10821 5146
rect 10979 5131 10988 5151
rect 11008 5131 11016 5151
rect 10979 5121 11016 5131
rect 11075 5151 11162 5161
rect 11075 5131 11084 5151
rect 11104 5131 11162 5151
rect 11075 5122 11162 5131
rect 11075 5121 11112 5122
rect 10343 5101 10380 5111
rect 10343 5099 10353 5101
rect 10277 5097 10353 5099
rect 9939 5041 10189 5065
rect 10274 5083 10353 5097
rect 10371 5083 10380 5101
rect 10274 5080 10380 5083
rect 9746 5021 9767 5040
rect 10274 5021 10300 5080
rect 10343 5074 10380 5080
rect 10787 5071 10824 5080
rect 8400 5016 8500 5020
rect 8400 5012 8462 5016
rect 8400 4986 8407 5012
rect 8433 4990 8462 5012
rect 8488 4990 8500 5016
rect 8433 4986 8500 4990
rect 8400 4983 8500 4986
rect 8568 4983 8603 5020
rect 8665 5017 9024 5020
rect 8665 5012 8887 5017
rect 8665 4988 8678 5012
rect 8702 4993 8887 5012
rect 8911 4993 9024 5017
rect 8702 4988 9024 4993
rect 8665 4984 9024 4988
rect 9091 5012 9240 5020
rect 9091 4992 9102 5012
rect 9122 4992 9240 5012
rect 9746 5003 10300 5021
rect 10785 5053 10796 5071
rect 10814 5053 10824 5071
rect 11131 5069 11162 5122
rect 11192 5151 11229 5222
rect 11400 5227 11793 5247
rect 11813 5227 11816 5247
rect 11400 5222 11816 5227
rect 12035 5241 12073 5250
rect 11400 5221 11741 5222
rect 12035 5221 12044 5241
rect 12064 5221 12073 5241
rect 11344 5161 11375 5162
rect 11192 5131 11201 5151
rect 11221 5131 11229 5151
rect 11192 5121 11229 5131
rect 11288 5154 11375 5161
rect 11288 5151 11349 5154
rect 11288 5131 11297 5151
rect 11317 5134 11349 5151
rect 11370 5134 11375 5154
rect 11317 5131 11375 5134
rect 11288 5124 11375 5131
rect 11400 5151 11437 5221
rect 11703 5220 11740 5221
rect 12035 5213 12073 5221
rect 12139 5245 12224 5251
rect 12249 5250 12286 5251
rect 12139 5225 12147 5245
rect 12167 5225 12224 5245
rect 12139 5217 12224 5225
rect 12248 5241 12286 5250
rect 12248 5221 12257 5241
rect 12277 5221 12286 5241
rect 12139 5216 12175 5217
rect 12248 5213 12286 5221
rect 12352 5245 12437 5251
rect 12457 5250 12494 5251
rect 12352 5225 12360 5245
rect 12380 5244 12437 5245
rect 12380 5225 12409 5244
rect 12352 5224 12409 5225
rect 12430 5224 12437 5244
rect 12352 5217 12437 5224
rect 12456 5241 12494 5250
rect 12456 5221 12465 5241
rect 12485 5221 12494 5241
rect 12352 5216 12388 5217
rect 12456 5213 12494 5221
rect 12560 5245 12704 5251
rect 12560 5225 12568 5245
rect 12588 5244 12676 5245
rect 12588 5225 12621 5244
rect 12644 5225 12676 5244
rect 12696 5225 12704 5245
rect 12560 5217 12704 5225
rect 12560 5216 12596 5217
rect 12668 5216 12704 5217
rect 12770 5250 12807 5251
rect 12770 5249 12808 5250
rect 12770 5241 12834 5249
rect 12770 5221 12779 5241
rect 12799 5227 12834 5241
rect 12854 5227 12857 5247
rect 12799 5222 12857 5227
rect 12799 5221 12834 5222
rect 12036 5184 12073 5213
rect 12037 5182 12073 5184
rect 12249 5182 12286 5213
rect 11552 5161 11588 5162
rect 11400 5131 11409 5151
rect 11429 5131 11437 5151
rect 11288 5122 11344 5124
rect 11288 5121 11325 5122
rect 11400 5121 11437 5131
rect 11496 5151 11644 5161
rect 12037 5160 12286 5182
rect 12457 5181 12494 5213
rect 12770 5209 12834 5221
rect 12874 5183 12901 5361
rect 12733 5181 12901 5183
rect 12457 5170 12901 5181
rect 12964 5181 12994 6182
rect 12964 5176 12996 5181
rect 11744 5158 11840 5160
rect 11496 5131 11505 5151
rect 11525 5131 11615 5151
rect 11635 5131 11644 5151
rect 11496 5122 11644 5131
rect 11702 5151 11840 5158
rect 12457 5155 12903 5170
rect 12733 5154 12903 5155
rect 11702 5131 11711 5151
rect 11731 5131 11840 5151
rect 11702 5122 11840 5131
rect 11496 5121 11533 5122
rect 11552 5070 11588 5122
rect 11607 5121 11644 5122
rect 11703 5121 11740 5122
rect 11023 5068 11064 5069
rect 10346 5010 10383 5012
rect 10274 5002 10300 5003
rect 10343 5002 10383 5010
rect 9091 4985 9240 4992
rect 10343 4990 10355 5002
rect 10334 4985 10355 4990
rect 9091 4984 9132 4985
rect 9750 4984 10355 4985
rect 10373 4984 10383 5002
rect 8415 4931 8452 4932
rect 8511 4931 8548 4932
rect 8567 4931 8603 4983
rect 8622 4931 8659 4932
rect 8315 4922 8453 4931
rect 8315 4902 8424 4922
rect 8444 4902 8453 4922
rect 8315 4895 8453 4902
rect 8511 4922 8659 4931
rect 8511 4902 8520 4922
rect 8540 4902 8630 4922
rect 8650 4902 8659 4922
rect 8315 4893 8411 4895
rect 8511 4892 8659 4902
rect 8718 4922 8755 4932
rect 8830 4931 8867 4932
rect 8811 4929 8867 4931
rect 8718 4902 8726 4922
rect 8746 4902 8755 4922
rect 8567 4891 8603 4892
rect 8415 4832 8452 4833
rect 8718 4832 8755 4902
rect 8780 4922 8867 4929
rect 8780 4919 8838 4922
rect 8780 4899 8785 4919
rect 8806 4902 8838 4919
rect 8858 4902 8867 4922
rect 8806 4899 8867 4902
rect 8780 4892 8867 4899
rect 8926 4922 8963 4932
rect 8926 4902 8934 4922
rect 8954 4902 8963 4922
rect 8780 4891 8811 4892
rect 8414 4831 8755 4832
rect 8339 4826 8755 4831
rect 8339 4806 8342 4826
rect 8362 4806 8755 4826
rect 8926 4831 8963 4902
rect 8993 4931 9024 4984
rect 9750 4975 10383 4984
rect 9750 4968 10382 4975
rect 9750 4966 9812 4968
rect 9328 4956 9496 4957
rect 9750 4956 9772 4966
rect 9043 4931 9080 4932
rect 8993 4922 9080 4931
rect 8993 4902 9051 4922
rect 9071 4902 9080 4922
rect 8993 4892 9080 4902
rect 9139 4922 9176 4932
rect 9139 4902 9147 4922
rect 9167 4902 9176 4922
rect 8993 4891 9024 4892
rect 9139 4831 9176 4902
rect 8926 4807 9176 4831
rect 9328 4930 9772 4956
rect 9328 4928 9496 4930
rect 9328 4750 9355 4928
rect 9395 4890 9459 4902
rect 9735 4898 9772 4930
rect 9943 4929 10192 4951
rect 9943 4898 9980 4929
rect 10156 4927 10192 4929
rect 10156 4898 10193 4927
rect 9395 4889 9430 4890
rect 9372 4884 9430 4889
rect 9372 4864 9375 4884
rect 9395 4870 9430 4884
rect 9450 4870 9459 4890
rect 9395 4862 9459 4870
rect 9421 4861 9459 4862
rect 9422 4860 9459 4861
rect 9525 4894 9561 4895
rect 9633 4894 9669 4895
rect 9525 4886 9669 4894
rect 9525 4866 9533 4886
rect 9553 4866 9582 4886
rect 9525 4865 9582 4866
rect 9604 4866 9641 4886
rect 9661 4866 9669 4886
rect 9604 4865 9669 4866
rect 9525 4860 9669 4865
rect 9735 4890 9773 4898
rect 9841 4894 9877 4895
rect 9735 4870 9744 4890
rect 9764 4870 9773 4890
rect 9735 4861 9773 4870
rect 9792 4887 9877 4894
rect 9792 4867 9799 4887
rect 9820 4886 9877 4887
rect 9820 4867 9849 4886
rect 9792 4866 9849 4867
rect 9869 4866 9877 4886
rect 9735 4860 9772 4861
rect 9792 4860 9877 4866
rect 9943 4890 9981 4898
rect 10054 4894 10090 4895
rect 9943 4870 9952 4890
rect 9972 4870 9981 4890
rect 9943 4861 9981 4870
rect 10005 4886 10090 4894
rect 10005 4866 10062 4886
rect 10082 4866 10090 4886
rect 9943 4860 9980 4861
rect 10005 4860 10090 4866
rect 10156 4890 10194 4898
rect 10156 4870 10165 4890
rect 10185 4870 10194 4890
rect 10156 4861 10194 4870
rect 10156 4860 10193 4861
rect 9579 4839 9615 4860
rect 10005 4839 10036 4860
rect 9412 4835 9512 4839
rect 9412 4831 9474 4835
rect 9412 4805 9419 4831
rect 9445 4809 9474 4831
rect 9500 4809 9512 4835
rect 9445 4805 9512 4809
rect 9412 4802 9512 4805
rect 9580 4802 9615 4839
rect 9677 4836 10036 4839
rect 9677 4831 9899 4836
rect 9677 4807 9690 4831
rect 9714 4812 9899 4831
rect 9923 4812 10036 4836
rect 9714 4807 10036 4812
rect 9677 4803 10036 4807
rect 10103 4831 10252 4839
rect 10103 4811 10114 4831
rect 10134 4811 10252 4831
rect 10103 4804 10252 4811
rect 10343 4819 10382 4968
rect 10785 4904 10824 5053
rect 10915 5061 11064 5068
rect 10915 5041 11033 5061
rect 11053 5041 11064 5061
rect 10915 5033 11064 5041
rect 11131 5065 11490 5069
rect 11131 5060 11453 5065
rect 11131 5036 11244 5060
rect 11268 5041 11453 5060
rect 11477 5041 11490 5065
rect 11268 5036 11490 5041
rect 11131 5033 11490 5036
rect 11552 5033 11587 5070
rect 11655 5067 11755 5070
rect 11655 5063 11722 5067
rect 11655 5037 11667 5063
rect 11693 5041 11722 5063
rect 11748 5041 11755 5067
rect 11693 5037 11755 5041
rect 11655 5033 11755 5037
rect 11131 5012 11162 5033
rect 11552 5012 11588 5033
rect 10974 5011 11011 5012
rect 10973 5002 11011 5011
rect 10973 4982 10982 5002
rect 11002 4982 11011 5002
rect 10973 4974 11011 4982
rect 11077 5006 11162 5012
rect 11187 5011 11224 5012
rect 11077 4986 11085 5006
rect 11105 4986 11162 5006
rect 11077 4978 11162 4986
rect 11186 5002 11224 5011
rect 11186 4982 11195 5002
rect 11215 4982 11224 5002
rect 11077 4977 11113 4978
rect 11186 4974 11224 4982
rect 11290 5006 11375 5012
rect 11395 5011 11432 5012
rect 11290 4986 11298 5006
rect 11318 5005 11375 5006
rect 11318 4986 11347 5005
rect 11290 4985 11347 4986
rect 11368 4985 11375 5005
rect 11290 4978 11375 4985
rect 11394 5002 11432 5011
rect 11394 4982 11403 5002
rect 11423 4982 11432 5002
rect 11290 4977 11326 4978
rect 11394 4974 11432 4982
rect 11498 5007 11642 5012
rect 11498 5006 11563 5007
rect 11498 4986 11506 5006
rect 11526 4986 11563 5006
rect 11585 5006 11642 5007
rect 11585 4986 11614 5006
rect 11634 4986 11642 5006
rect 11498 4978 11642 4986
rect 11498 4977 11534 4978
rect 11606 4977 11642 4978
rect 11708 5011 11745 5012
rect 11708 5010 11746 5011
rect 11708 5002 11772 5010
rect 11708 4982 11717 5002
rect 11737 4988 11772 5002
rect 11792 4988 11795 5008
rect 11737 4983 11795 4988
rect 11737 4982 11772 4983
rect 10974 4945 11011 4974
rect 10975 4943 11011 4945
rect 11187 4943 11224 4974
rect 10975 4921 11224 4943
rect 11395 4942 11432 4974
rect 11708 4970 11772 4982
rect 11812 4944 11839 5122
rect 11671 4942 11839 4944
rect 11395 4916 11839 4942
rect 11991 5041 12241 5065
rect 11991 4970 12028 5041
rect 12143 4980 12174 4981
rect 11991 4950 12000 4970
rect 12020 4950 12028 4970
rect 11991 4940 12028 4950
rect 12087 4970 12174 4980
rect 12087 4950 12096 4970
rect 12116 4950 12174 4970
rect 12087 4941 12174 4950
rect 12087 4940 12124 4941
rect 11395 4906 11417 4916
rect 11671 4915 11839 4916
rect 11355 4904 11417 4906
rect 10785 4897 11417 4904
rect 10784 4888 11417 4897
rect 12143 4888 12174 4941
rect 12204 4970 12241 5041
rect 12412 5046 12805 5066
rect 12825 5046 12828 5066
rect 12412 5041 12828 5046
rect 12412 5040 12753 5041
rect 12356 4980 12387 4981
rect 12204 4950 12213 4970
rect 12233 4950 12241 4970
rect 12204 4940 12241 4950
rect 12300 4973 12387 4980
rect 12300 4970 12361 4973
rect 12300 4950 12309 4970
rect 12329 4953 12361 4970
rect 12382 4953 12387 4973
rect 12329 4950 12387 4953
rect 12300 4943 12387 4950
rect 12412 4970 12449 5040
rect 12715 5039 12752 5040
rect 12564 4980 12600 4981
rect 12412 4950 12421 4970
rect 12441 4950 12449 4970
rect 12300 4941 12356 4943
rect 12300 4940 12337 4941
rect 12412 4940 12449 4950
rect 12508 4970 12656 4980
rect 12756 4977 12852 4979
rect 12508 4950 12517 4970
rect 12537 4950 12627 4970
rect 12647 4950 12656 4970
rect 12508 4941 12656 4950
rect 12714 4970 12852 4977
rect 12714 4950 12723 4970
rect 12743 4950 12852 4970
rect 12714 4941 12852 4950
rect 12508 4940 12545 4941
rect 12564 4889 12600 4941
rect 12619 4940 12656 4941
rect 12715 4940 12752 4941
rect 10784 4870 10794 4888
rect 10812 4887 11417 4888
rect 12035 4887 12076 4888
rect 10812 4882 10833 4887
rect 10812 4870 10824 4882
rect 11927 4880 12076 4887
rect 10784 4862 10824 4870
rect 10867 4869 10893 4870
rect 10784 4860 10821 4862
rect 10103 4803 10144 4804
rect 9427 4750 9464 4751
rect 9523 4750 9560 4751
rect 9579 4750 9615 4802
rect 9634 4750 9671 4751
rect 9327 4741 9465 4750
rect 9327 4721 9436 4741
rect 9456 4721 9465 4741
rect 9327 4714 9465 4721
rect 9523 4741 9671 4750
rect 9523 4721 9532 4741
rect 9552 4721 9642 4741
rect 9662 4721 9671 4741
rect 9327 4712 9423 4714
rect 9523 4711 9671 4721
rect 9730 4741 9767 4751
rect 9842 4750 9879 4751
rect 9823 4748 9879 4750
rect 9730 4721 9738 4741
rect 9758 4721 9767 4741
rect 9579 4710 9615 4711
rect 7492 4702 7523 4705
rect 8021 4705 8189 4706
rect 6321 4678 6459 4687
rect 8021 4679 8465 4705
rect 6115 4677 6152 4678
rect 6171 4626 6207 4678
rect 6226 4677 6263 4678
rect 6322 4677 6359 4678
rect 5642 4624 5683 4625
rect 4449 4602 5098 4608
rect 5534 4617 5683 4624
rect 4449 4601 5097 4602
rect 3515 4581 3526 4601
rect 3546 4581 3664 4601
rect 5060 4599 5097 4601
rect 5534 4597 5652 4617
rect 5672 4597 5683 4617
rect 5534 4589 5683 4597
rect 5750 4621 6109 4625
rect 5750 4616 6072 4621
rect 5750 4592 5863 4616
rect 5887 4597 6072 4616
rect 6096 4597 6109 4621
rect 5887 4592 6109 4597
rect 5750 4589 6109 4592
rect 6171 4589 6206 4626
rect 6274 4623 6374 4626
rect 6274 4619 6341 4623
rect 6274 4593 6286 4619
rect 6312 4597 6341 4619
rect 6367 4597 6374 4623
rect 6312 4593 6374 4597
rect 6274 4589 6374 4593
rect 3515 4574 3664 4581
rect 3515 4573 3556 4574
rect 2839 4520 2876 4521
rect 2935 4520 2972 4521
rect 2991 4520 3027 4572
rect 3046 4520 3083 4521
rect 733 4493 1177 4519
rect 734 4476 758 4493
rect 1009 4492 1177 4493
rect 1628 4489 1878 4513
rect 132 4458 759 4476
rect 132 4457 170 4458
rect 130 4452 170 4457
rect 130 4409 165 4452
rect 128 4400 165 4409
rect 128 4382 138 4400
rect 156 4382 165 4400
rect 1628 4418 1665 4489
rect 1780 4428 1811 4429
rect 1628 4398 1637 4418
rect 1657 4398 1665 4418
rect 1628 4388 1665 4398
rect 1724 4418 1811 4428
rect 1724 4398 1733 4418
rect 1753 4398 1811 4418
rect 1724 4389 1811 4398
rect 1724 4388 1761 4389
rect 128 4372 165 4382
rect 1780 4336 1811 4389
rect 1841 4418 1878 4489
rect 2049 4494 2442 4514
rect 2462 4494 2465 4514
rect 2049 4489 2465 4494
rect 2739 4511 2877 4520
rect 2739 4491 2848 4511
rect 2868 4491 2877 4511
rect 2049 4488 2390 4489
rect 1993 4428 2024 4429
rect 1841 4398 1850 4418
rect 1870 4398 1878 4418
rect 1841 4388 1878 4398
rect 1937 4421 2024 4428
rect 1937 4418 1998 4421
rect 1937 4398 1946 4418
rect 1966 4401 1998 4418
rect 2019 4401 2024 4421
rect 1966 4398 2024 4401
rect 1937 4391 2024 4398
rect 2049 4418 2086 4488
rect 2352 4487 2389 4488
rect 2739 4484 2877 4491
rect 2935 4511 3083 4520
rect 2935 4491 2944 4511
rect 2964 4491 3054 4511
rect 3074 4491 3083 4511
rect 2739 4482 2835 4484
rect 2935 4481 3083 4491
rect 3142 4511 3179 4521
rect 3254 4520 3291 4521
rect 3235 4518 3291 4520
rect 3142 4491 3150 4511
rect 3170 4491 3179 4511
rect 2991 4480 3027 4481
rect 2201 4428 2237 4429
rect 2049 4398 2058 4418
rect 2078 4398 2086 4418
rect 1937 4389 1993 4391
rect 1937 4388 1974 4389
rect 2049 4388 2086 4398
rect 2145 4418 2293 4428
rect 2393 4425 2489 4427
rect 2145 4398 2154 4418
rect 2174 4398 2264 4418
rect 2284 4398 2293 4418
rect 2145 4389 2293 4398
rect 2351 4418 2489 4425
rect 2839 4421 2876 4422
rect 3142 4421 3179 4491
rect 3204 4511 3291 4518
rect 3204 4508 3262 4511
rect 3204 4488 3209 4508
rect 3230 4491 3262 4508
rect 3282 4491 3291 4511
rect 3230 4488 3291 4491
rect 3204 4481 3291 4488
rect 3350 4511 3387 4521
rect 3350 4491 3358 4511
rect 3378 4491 3387 4511
rect 3204 4480 3235 4481
rect 2838 4420 3179 4421
rect 2351 4398 2360 4418
rect 2380 4398 2489 4418
rect 2351 4389 2489 4398
rect 2763 4415 3179 4420
rect 2763 4395 2766 4415
rect 2786 4395 3179 4415
rect 3350 4420 3387 4491
rect 3417 4520 3448 4573
rect 5750 4568 5781 4589
rect 6171 4568 6207 4589
rect 5414 4559 5451 4568
rect 5593 4567 5630 4568
rect 5414 4541 5423 4559
rect 5441 4541 5451 4559
rect 5063 4527 5100 4537
rect 5414 4531 5451 4541
rect 3467 4520 3504 4521
rect 3417 4511 3504 4520
rect 3417 4491 3475 4511
rect 3495 4491 3504 4511
rect 3417 4481 3504 4491
rect 3563 4511 3600 4521
rect 3563 4491 3571 4511
rect 3591 4491 3600 4511
rect 3417 4480 3448 4481
rect 3563 4420 3600 4491
rect 5063 4509 5072 4527
rect 5090 4509 5100 4527
rect 5063 4500 5100 4509
rect 5063 4457 5098 4500
rect 5415 4496 5451 4531
rect 5592 4558 5630 4567
rect 5592 4538 5601 4558
rect 5621 4538 5630 4558
rect 5592 4530 5630 4538
rect 5696 4562 5781 4568
rect 5806 4567 5843 4568
rect 5696 4542 5704 4562
rect 5724 4542 5781 4562
rect 5696 4534 5781 4542
rect 5805 4558 5843 4567
rect 5805 4538 5814 4558
rect 5834 4538 5843 4558
rect 5696 4533 5732 4534
rect 5805 4530 5843 4538
rect 5909 4562 5994 4568
rect 6014 4567 6051 4568
rect 5909 4542 5917 4562
rect 5937 4561 5994 4562
rect 5937 4542 5966 4561
rect 5909 4541 5966 4542
rect 5987 4541 5994 4561
rect 5909 4534 5994 4541
rect 6013 4558 6051 4567
rect 6013 4538 6022 4558
rect 6042 4538 6051 4558
rect 5909 4533 5945 4534
rect 6013 4530 6051 4538
rect 6117 4562 6261 4568
rect 6117 4542 6125 4562
rect 6145 4561 6233 4562
rect 6145 4542 6173 4561
rect 6117 4540 6173 4542
rect 6195 4542 6233 4561
rect 6253 4542 6261 4562
rect 6195 4540 6261 4542
rect 6117 4534 6261 4540
rect 6117 4533 6153 4534
rect 6225 4533 6261 4534
rect 6327 4567 6364 4568
rect 6327 4566 6365 4567
rect 6327 4558 6391 4566
rect 6327 4538 6336 4558
rect 6356 4544 6391 4558
rect 6411 4544 6414 4564
rect 6356 4539 6414 4544
rect 6356 4538 6391 4539
rect 5593 4501 5630 4530
rect 5058 4452 5098 4457
rect 5413 4455 5451 4496
rect 5594 4499 5630 4501
rect 5806 4499 5843 4530
rect 5594 4477 5843 4499
rect 6014 4498 6051 4530
rect 6327 4526 6391 4538
rect 6431 4500 6458 4678
rect 6290 4498 6458 4500
rect 8021 4677 8189 4679
rect 8021 4674 8068 4677
rect 8021 4499 8048 4674
rect 8088 4639 8152 4651
rect 8428 4647 8465 4679
rect 8636 4678 8885 4700
rect 8636 4647 8673 4678
rect 8849 4676 8885 4678
rect 8849 4647 8886 4676
rect 9427 4651 9464 4652
rect 9730 4651 9767 4721
rect 9792 4741 9879 4748
rect 9792 4738 9850 4741
rect 9792 4718 9797 4738
rect 9818 4721 9850 4738
rect 9870 4721 9879 4741
rect 9818 4718 9879 4721
rect 9792 4711 9879 4718
rect 9938 4741 9975 4751
rect 9938 4721 9946 4741
rect 9966 4721 9975 4741
rect 9792 4710 9823 4711
rect 9426 4650 9767 4651
rect 8088 4638 8123 4639
rect 8065 4633 8123 4638
rect 8065 4613 8068 4633
rect 8088 4619 8123 4633
rect 8143 4619 8152 4639
rect 8088 4611 8152 4619
rect 8114 4610 8152 4611
rect 8115 4609 8152 4610
rect 8218 4643 8254 4644
rect 8326 4643 8362 4644
rect 8218 4635 8362 4643
rect 8218 4615 8226 4635
rect 8246 4633 8334 4635
rect 8246 4615 8272 4633
rect 8218 4614 8272 4615
rect 8298 4615 8334 4633
rect 8354 4615 8362 4635
rect 8298 4614 8362 4615
rect 8218 4609 8362 4614
rect 8428 4639 8466 4647
rect 8534 4643 8570 4644
rect 8428 4619 8437 4639
rect 8457 4619 8466 4639
rect 8428 4610 8466 4619
rect 8485 4636 8570 4643
rect 8485 4616 8492 4636
rect 8513 4635 8570 4636
rect 8513 4616 8542 4635
rect 8485 4615 8542 4616
rect 8562 4615 8570 4635
rect 8428 4609 8465 4610
rect 8485 4609 8570 4615
rect 8636 4639 8674 4647
rect 8747 4643 8783 4644
rect 8636 4619 8645 4639
rect 8665 4619 8674 4639
rect 8636 4610 8674 4619
rect 8698 4635 8783 4643
rect 8698 4615 8755 4635
rect 8775 4615 8783 4635
rect 8636 4609 8673 4610
rect 8698 4609 8783 4615
rect 8849 4639 8887 4647
rect 8849 4619 8858 4639
rect 8878 4619 8887 4639
rect 9351 4645 9767 4650
rect 9351 4625 9354 4645
rect 9374 4625 9767 4645
rect 9938 4650 9975 4721
rect 10005 4750 10036 4803
rect 10343 4801 10353 4819
rect 10371 4801 10382 4819
rect 10867 4851 11421 4869
rect 11927 4860 12045 4880
rect 12065 4860 12076 4880
rect 11927 4852 12076 4860
rect 12143 4884 12502 4888
rect 12143 4879 12465 4884
rect 12143 4855 12256 4879
rect 12280 4860 12465 4879
rect 12489 4860 12502 4884
rect 12280 4855 12502 4860
rect 12143 4852 12502 4855
rect 12564 4852 12599 4889
rect 12667 4886 12767 4889
rect 12667 4882 12734 4886
rect 12667 4856 12679 4882
rect 12705 4860 12734 4882
rect 12760 4860 12767 4886
rect 12705 4856 12767 4860
rect 12667 4852 12767 4856
rect 10343 4792 10380 4801
rect 10787 4792 10824 4798
rect 10867 4792 10893 4851
rect 11400 4832 11421 4851
rect 10787 4789 10893 4792
rect 10787 4771 10796 4789
rect 10814 4775 10893 4789
rect 10978 4807 11228 4831
rect 10814 4773 10890 4775
rect 10814 4771 10824 4773
rect 10787 4761 10824 4771
rect 10055 4750 10092 4751
rect 10005 4741 10092 4750
rect 10005 4721 10063 4741
rect 10083 4721 10092 4741
rect 10005 4711 10092 4721
rect 10151 4741 10188 4751
rect 10151 4721 10159 4741
rect 10179 4721 10188 4741
rect 10346 4726 10383 4730
rect 10005 4710 10036 4711
rect 10151 4650 10188 4721
rect 9938 4626 10188 4650
rect 10344 4720 10383 4726
rect 10344 4702 10355 4720
rect 10373 4702 10383 4720
rect 10344 4693 10383 4702
rect 10792 4696 10823 4761
rect 10978 4736 11015 4807
rect 11130 4746 11161 4747
rect 10978 4716 10987 4736
rect 11007 4716 11015 4736
rect 10978 4706 11015 4716
rect 11074 4736 11161 4746
rect 11074 4716 11083 4736
rect 11103 4716 11161 4736
rect 11074 4707 11161 4716
rect 11074 4706 11111 4707
rect 8849 4610 8887 4619
rect 8849 4609 8886 4610
rect 8272 4588 8308 4609
rect 8698 4588 8729 4609
rect 9730 4602 9767 4625
rect 10344 4615 10379 4693
rect 10791 4687 10828 4696
rect 10791 4669 10801 4687
rect 10819 4669 10828 4687
rect 10791 4659 10828 4669
rect 11130 4654 11161 4707
rect 11191 4736 11228 4807
rect 11399 4812 11792 4832
rect 11812 4812 11815 4832
rect 12143 4831 12174 4852
rect 12564 4831 12600 4852
rect 11986 4830 12023 4831
rect 11399 4807 11815 4812
rect 11985 4821 12023 4830
rect 11399 4806 11740 4807
rect 11343 4746 11374 4747
rect 11191 4716 11200 4736
rect 11220 4716 11228 4736
rect 11191 4706 11228 4716
rect 11287 4739 11374 4746
rect 11287 4736 11348 4739
rect 11287 4716 11296 4736
rect 11316 4719 11348 4736
rect 11369 4719 11374 4739
rect 11316 4716 11374 4719
rect 11287 4709 11374 4716
rect 11399 4736 11436 4806
rect 11702 4805 11739 4806
rect 11985 4801 11994 4821
rect 12014 4801 12023 4821
rect 11985 4793 12023 4801
rect 12089 4825 12174 4831
rect 12199 4830 12236 4831
rect 12089 4805 12097 4825
rect 12117 4805 12174 4825
rect 12089 4797 12174 4805
rect 12198 4821 12236 4830
rect 12198 4801 12207 4821
rect 12227 4801 12236 4821
rect 12089 4796 12125 4797
rect 12198 4793 12236 4801
rect 12302 4825 12387 4831
rect 12407 4830 12444 4831
rect 12302 4805 12310 4825
rect 12330 4824 12387 4825
rect 12330 4805 12359 4824
rect 12302 4804 12359 4805
rect 12380 4804 12387 4824
rect 12302 4797 12387 4804
rect 12406 4821 12444 4830
rect 12406 4801 12415 4821
rect 12435 4801 12444 4821
rect 12302 4796 12338 4797
rect 12406 4793 12444 4801
rect 12510 4826 12654 4831
rect 12510 4825 12569 4826
rect 12510 4805 12518 4825
rect 12538 4806 12569 4825
rect 12593 4825 12654 4826
rect 12593 4806 12626 4825
rect 12538 4805 12626 4806
rect 12646 4805 12654 4825
rect 12510 4797 12654 4805
rect 12510 4796 12546 4797
rect 12618 4796 12654 4797
rect 12720 4830 12757 4831
rect 12720 4829 12758 4830
rect 12720 4821 12784 4829
rect 12720 4801 12729 4821
rect 12749 4807 12784 4821
rect 12804 4807 12807 4827
rect 12749 4802 12807 4807
rect 12749 4801 12784 4802
rect 11986 4764 12023 4793
rect 11987 4762 12023 4764
rect 12199 4762 12236 4793
rect 11551 4746 11587 4747
rect 11399 4716 11408 4736
rect 11428 4716 11436 4736
rect 11287 4707 11343 4709
rect 11287 4706 11324 4707
rect 11399 4706 11436 4716
rect 11495 4736 11643 4746
rect 11743 4743 11839 4745
rect 11495 4716 11504 4736
rect 11524 4716 11614 4736
rect 11634 4716 11643 4736
rect 11495 4707 11643 4716
rect 11701 4736 11839 4743
rect 11987 4740 12236 4762
rect 12407 4761 12444 4793
rect 12720 4789 12784 4801
rect 12824 4763 12851 4941
rect 12683 4761 12851 4763
rect 12407 4757 12851 4761
rect 11701 4716 11710 4736
rect 11730 4716 11839 4736
rect 12407 4738 12456 4757
rect 12476 4738 12851 4757
rect 12407 4735 12851 4738
rect 12683 4734 12851 4735
rect 12872 4760 12903 5154
rect 12964 5158 12969 5176
rect 12989 5158 12996 5176
rect 12964 5153 12996 5158
rect 12967 5151 12996 5153
rect 12872 4734 12877 4760
rect 12896 4734 12903 4760
rect 13410 4735 13448 6566
rect 13476 6453 13503 6631
rect 13543 6593 13607 6605
rect 13883 6601 13920 6633
rect 14091 6632 14340 6654
rect 14795 6640 14832 6641
rect 15098 6640 15135 6710
rect 15160 6730 15247 6737
rect 15160 6727 15218 6730
rect 15160 6707 15165 6727
rect 15186 6710 15218 6727
rect 15238 6710 15247 6730
rect 15186 6707 15247 6710
rect 15160 6700 15247 6707
rect 15306 6730 15343 6740
rect 15306 6710 15314 6730
rect 15334 6710 15343 6730
rect 15160 6699 15191 6700
rect 14794 6639 15135 6640
rect 14091 6601 14128 6632
rect 14304 6630 14340 6632
rect 14719 6634 15135 6639
rect 14304 6601 14341 6630
rect 14719 6614 14722 6634
rect 14742 6614 15135 6634
rect 15306 6639 15343 6710
rect 15373 6739 15404 6792
rect 15711 6790 15721 6808
rect 15739 6790 15750 6808
rect 16053 6827 16686 6836
rect 17412 6827 17443 6880
rect 17473 6909 17510 6980
rect 17681 6985 18074 7005
rect 18094 6985 18097 7005
rect 17681 6980 18097 6985
rect 17681 6979 18022 6980
rect 17625 6919 17656 6920
rect 17473 6889 17482 6909
rect 17502 6889 17510 6909
rect 17473 6879 17510 6889
rect 17569 6912 17656 6919
rect 17569 6909 17630 6912
rect 17569 6889 17578 6909
rect 17598 6892 17630 6909
rect 17651 6892 17656 6912
rect 17598 6889 17656 6892
rect 17569 6882 17656 6889
rect 17681 6909 17718 6979
rect 17984 6978 18021 6979
rect 17833 6919 17869 6920
rect 17681 6889 17690 6909
rect 17710 6889 17718 6909
rect 17569 6880 17625 6882
rect 17569 6879 17606 6880
rect 17681 6879 17718 6889
rect 17777 6909 17925 6919
rect 18025 6916 18121 6918
rect 17777 6889 17786 6909
rect 17806 6889 17896 6909
rect 17916 6889 17925 6909
rect 17777 6880 17925 6889
rect 17983 6909 18121 6916
rect 17983 6889 17992 6909
rect 18012 6889 18121 6909
rect 17983 6880 18121 6889
rect 17777 6879 17814 6880
rect 17833 6828 17869 6880
rect 17888 6879 17925 6880
rect 17984 6879 18021 6880
rect 16053 6809 16063 6827
rect 16081 6826 16686 6827
rect 17304 6826 17345 6827
rect 16081 6821 16102 6826
rect 16081 6809 16093 6821
rect 17196 6819 17345 6826
rect 16053 6801 16093 6809
rect 16136 6808 16162 6809
rect 16053 6799 16090 6801
rect 16136 6790 16690 6808
rect 17196 6799 17314 6819
rect 17334 6799 17345 6819
rect 17196 6791 17345 6799
rect 17412 6823 17771 6827
rect 17412 6818 17734 6823
rect 17412 6794 17525 6818
rect 17549 6799 17734 6818
rect 17758 6799 17771 6823
rect 17549 6794 17771 6799
rect 17412 6791 17771 6794
rect 17833 6791 17868 6828
rect 17936 6825 18036 6828
rect 17936 6821 18003 6825
rect 17936 6795 17948 6821
rect 17974 6799 18003 6821
rect 18029 6799 18036 6825
rect 17974 6795 18036 6799
rect 17936 6791 18036 6795
rect 15711 6781 15748 6790
rect 15423 6739 15460 6740
rect 15373 6730 15460 6739
rect 15373 6710 15431 6730
rect 15451 6710 15460 6730
rect 15373 6700 15460 6710
rect 15519 6730 15556 6740
rect 15519 6710 15527 6730
rect 15547 6710 15556 6730
rect 16056 6731 16093 6737
rect 16136 6731 16162 6790
rect 16669 6771 16690 6790
rect 16056 6728 16162 6731
rect 15714 6715 15751 6719
rect 15373 6699 15404 6700
rect 15519 6639 15556 6710
rect 15306 6615 15556 6639
rect 15712 6709 15751 6715
rect 15712 6691 15723 6709
rect 15741 6691 15751 6709
rect 16056 6710 16065 6728
rect 16083 6714 16162 6728
rect 16247 6746 16497 6770
rect 16083 6712 16159 6714
rect 16083 6710 16093 6712
rect 16056 6700 16093 6710
rect 15712 6682 15751 6691
rect 13543 6592 13578 6593
rect 13520 6587 13578 6592
rect 13520 6567 13523 6587
rect 13543 6573 13578 6587
rect 13598 6573 13607 6593
rect 13543 6565 13607 6573
rect 13569 6564 13607 6565
rect 13570 6563 13607 6564
rect 13673 6597 13709 6598
rect 13781 6597 13817 6598
rect 13673 6589 13817 6597
rect 13673 6569 13681 6589
rect 13701 6588 13789 6589
rect 13701 6569 13730 6588
rect 13753 6569 13789 6588
rect 13809 6569 13817 6589
rect 13673 6563 13817 6569
rect 13883 6593 13921 6601
rect 13989 6597 14025 6598
rect 13883 6573 13892 6593
rect 13912 6573 13921 6593
rect 13883 6564 13921 6573
rect 13940 6590 14025 6597
rect 13940 6570 13947 6590
rect 13968 6589 14025 6590
rect 13968 6570 13997 6589
rect 13940 6569 13997 6570
rect 14017 6569 14025 6589
rect 13883 6563 13920 6564
rect 13940 6563 14025 6569
rect 14091 6593 14129 6601
rect 14202 6597 14238 6598
rect 14091 6573 14100 6593
rect 14120 6573 14129 6593
rect 14091 6564 14129 6573
rect 14153 6589 14238 6597
rect 14153 6569 14210 6589
rect 14230 6569 14238 6589
rect 14091 6563 14128 6564
rect 14153 6563 14238 6569
rect 14304 6593 14342 6601
rect 14304 6573 14313 6593
rect 14333 6573 14342 6593
rect 14304 6564 14342 6573
rect 15098 6591 15135 6614
rect 15712 6604 15747 6682
rect 16061 6635 16092 6700
rect 16247 6675 16284 6746
rect 16399 6685 16430 6686
rect 16247 6655 16256 6675
rect 16276 6655 16284 6675
rect 16247 6645 16284 6655
rect 16343 6675 16430 6685
rect 16343 6655 16352 6675
rect 16372 6655 16430 6675
rect 16343 6646 16430 6655
rect 16343 6645 16380 6646
rect 15709 6594 15747 6604
rect 16060 6626 16097 6635
rect 16060 6608 16070 6626
rect 16088 6608 16097 6626
rect 16060 6598 16097 6608
rect 15098 6590 15268 6591
rect 15709 6590 15719 6594
rect 15098 6576 15719 6590
rect 15737 6576 15747 6594
rect 16399 6593 16430 6646
rect 16460 6675 16497 6746
rect 16668 6751 17061 6771
rect 17081 6751 17084 6771
rect 17412 6770 17443 6791
rect 17833 6770 17869 6791
rect 17255 6769 17292 6770
rect 16668 6746 17084 6751
rect 17254 6760 17292 6769
rect 16668 6745 17009 6746
rect 16612 6685 16643 6686
rect 16460 6655 16469 6675
rect 16489 6655 16497 6675
rect 16460 6645 16497 6655
rect 16556 6678 16643 6685
rect 16556 6675 16617 6678
rect 16556 6655 16565 6675
rect 16585 6658 16617 6675
rect 16638 6658 16643 6678
rect 16585 6655 16643 6658
rect 16556 6648 16643 6655
rect 16668 6675 16705 6745
rect 16971 6744 17008 6745
rect 17254 6740 17263 6760
rect 17283 6740 17292 6760
rect 17254 6732 17292 6740
rect 17358 6764 17443 6770
rect 17468 6769 17505 6770
rect 17358 6744 17366 6764
rect 17386 6744 17443 6764
rect 17358 6736 17443 6744
rect 17467 6760 17505 6769
rect 17467 6740 17476 6760
rect 17496 6740 17505 6760
rect 17358 6735 17394 6736
rect 17467 6732 17505 6740
rect 17571 6764 17656 6770
rect 17676 6769 17713 6770
rect 17571 6744 17579 6764
rect 17599 6763 17656 6764
rect 17599 6744 17628 6763
rect 17571 6743 17628 6744
rect 17649 6743 17656 6763
rect 17571 6736 17656 6743
rect 17675 6760 17713 6769
rect 17675 6740 17684 6760
rect 17704 6740 17713 6760
rect 17571 6735 17607 6736
rect 17675 6732 17713 6740
rect 17779 6765 17923 6770
rect 17779 6764 17838 6765
rect 17779 6744 17787 6764
rect 17807 6745 17838 6764
rect 17862 6764 17923 6765
rect 17862 6745 17895 6764
rect 17807 6744 17895 6745
rect 17915 6744 17923 6764
rect 17779 6736 17923 6744
rect 17779 6735 17815 6736
rect 17887 6735 17923 6736
rect 17989 6769 18026 6770
rect 17989 6768 18027 6769
rect 17989 6760 18053 6768
rect 17989 6740 17998 6760
rect 18018 6746 18053 6760
rect 18073 6746 18076 6766
rect 18018 6741 18076 6746
rect 18018 6740 18053 6741
rect 17255 6703 17292 6732
rect 17256 6701 17292 6703
rect 17468 6701 17505 6732
rect 16820 6685 16856 6686
rect 16668 6655 16677 6675
rect 16697 6655 16705 6675
rect 16556 6646 16612 6648
rect 16556 6645 16593 6646
rect 16668 6645 16705 6655
rect 16764 6675 16912 6685
rect 17012 6682 17108 6684
rect 16764 6655 16773 6675
rect 16793 6655 16883 6675
rect 16903 6655 16912 6675
rect 16764 6646 16912 6655
rect 16970 6675 17108 6682
rect 17256 6679 17505 6701
rect 17676 6700 17713 6732
rect 17989 6728 18053 6740
rect 18093 6702 18120 6880
rect 17952 6700 18120 6702
rect 17676 6696 18120 6700
rect 16970 6655 16979 6675
rect 16999 6655 17108 6675
rect 17676 6677 17725 6696
rect 17745 6677 18120 6696
rect 17676 6674 18120 6677
rect 17952 6673 18120 6674
rect 18141 6699 18172 7093
rect 18141 6673 18146 6699
rect 18165 6673 18172 6699
rect 18141 6670 18172 6673
rect 16970 6646 17108 6655
rect 16764 6645 16801 6646
rect 16820 6594 16856 6646
rect 16875 6645 16912 6646
rect 16971 6645 17008 6646
rect 16291 6592 16332 6593
rect 15098 6570 15747 6576
rect 16183 6585 16332 6592
rect 15098 6569 15746 6570
rect 15709 6567 15746 6569
rect 16183 6565 16301 6585
rect 16321 6565 16332 6585
rect 14304 6563 14341 6564
rect 13727 6542 13763 6563
rect 14153 6542 14184 6563
rect 16183 6557 16332 6565
rect 16399 6589 16758 6593
rect 16399 6584 16721 6589
rect 16399 6560 16512 6584
rect 16536 6565 16721 6584
rect 16745 6565 16758 6589
rect 16536 6560 16758 6565
rect 16399 6557 16758 6560
rect 16820 6557 16855 6594
rect 16923 6591 17023 6594
rect 16923 6587 16990 6591
rect 16923 6561 16935 6587
rect 16961 6565 16990 6587
rect 17016 6565 17023 6591
rect 16961 6561 17023 6565
rect 16923 6557 17023 6561
rect 13560 6538 13660 6542
rect 13560 6534 13622 6538
rect 13560 6508 13567 6534
rect 13593 6512 13622 6534
rect 13648 6512 13660 6538
rect 13593 6508 13660 6512
rect 13560 6505 13660 6508
rect 13728 6505 13763 6542
rect 13825 6539 14184 6542
rect 13825 6534 14047 6539
rect 13825 6510 13838 6534
rect 13862 6515 14047 6534
rect 14071 6515 14184 6539
rect 13862 6510 14184 6515
rect 13825 6506 14184 6510
rect 14251 6534 14400 6542
rect 16399 6536 16430 6557
rect 16820 6536 16856 6557
rect 14251 6514 14262 6534
rect 14282 6514 14400 6534
rect 14251 6507 14400 6514
rect 16063 6527 16100 6536
rect 16242 6535 16279 6536
rect 16063 6509 16072 6527
rect 16090 6509 16100 6527
rect 14251 6506 14292 6507
rect 13575 6453 13612 6454
rect 13671 6453 13708 6454
rect 13727 6453 13763 6505
rect 13782 6453 13819 6454
rect 13475 6444 13613 6453
rect 13475 6424 13584 6444
rect 13604 6424 13613 6444
rect 13475 6417 13613 6424
rect 13671 6444 13819 6453
rect 13671 6424 13680 6444
rect 13700 6424 13790 6444
rect 13810 6424 13819 6444
rect 13475 6415 13571 6417
rect 13671 6414 13819 6424
rect 13878 6444 13915 6454
rect 13990 6453 14027 6454
rect 13971 6451 14027 6453
rect 13878 6424 13886 6444
rect 13906 6424 13915 6444
rect 13727 6413 13763 6414
rect 13575 6354 13612 6355
rect 13878 6354 13915 6424
rect 13940 6444 14027 6451
rect 13940 6441 13998 6444
rect 13940 6421 13945 6441
rect 13966 6424 13998 6441
rect 14018 6424 14027 6444
rect 13966 6421 14027 6424
rect 13940 6414 14027 6421
rect 14086 6444 14123 6454
rect 14086 6424 14094 6444
rect 14114 6424 14123 6444
rect 13940 6413 13971 6414
rect 13574 6353 13915 6354
rect 13499 6348 13915 6353
rect 13499 6328 13502 6348
rect 13522 6328 13915 6348
rect 14086 6353 14123 6424
rect 14153 6453 14184 6506
rect 15712 6495 15749 6505
rect 16063 6499 16100 6509
rect 15712 6477 15721 6495
rect 15739 6477 15749 6495
rect 15712 6468 15749 6477
rect 14203 6453 14240 6454
rect 14153 6444 14240 6453
rect 14153 6424 14211 6444
rect 14231 6424 14240 6444
rect 14153 6414 14240 6424
rect 14299 6444 14336 6454
rect 14299 6424 14307 6444
rect 14327 6424 14336 6444
rect 14153 6413 14184 6414
rect 14299 6353 14336 6424
rect 15712 6422 15747 6468
rect 16064 6464 16100 6499
rect 16241 6526 16279 6535
rect 16241 6506 16250 6526
rect 16270 6506 16279 6526
rect 16241 6498 16279 6506
rect 16345 6530 16430 6536
rect 16455 6535 16492 6536
rect 16345 6510 16353 6530
rect 16373 6510 16430 6530
rect 16345 6502 16430 6510
rect 16454 6526 16492 6535
rect 16454 6506 16463 6526
rect 16483 6506 16492 6526
rect 16345 6501 16381 6502
rect 16454 6498 16492 6506
rect 16558 6530 16643 6536
rect 16663 6535 16700 6536
rect 16558 6510 16566 6530
rect 16586 6529 16643 6530
rect 16586 6510 16615 6529
rect 16558 6509 16615 6510
rect 16636 6509 16643 6529
rect 16558 6502 16643 6509
rect 16662 6526 16700 6535
rect 16662 6506 16671 6526
rect 16691 6506 16700 6526
rect 16558 6501 16594 6502
rect 16662 6498 16700 6506
rect 16766 6530 16910 6536
rect 16766 6510 16774 6530
rect 16794 6529 16882 6530
rect 16794 6510 16822 6529
rect 16766 6508 16822 6510
rect 16844 6510 16882 6529
rect 16902 6510 16910 6530
rect 16844 6508 16910 6510
rect 16766 6502 16910 6508
rect 16766 6501 16802 6502
rect 16874 6501 16910 6502
rect 16976 6535 17013 6536
rect 16976 6534 17014 6535
rect 16976 6526 17040 6534
rect 16976 6506 16985 6526
rect 17005 6512 17040 6526
rect 17060 6512 17063 6532
rect 17005 6507 17063 6512
rect 17005 6506 17040 6507
rect 16242 6469 16279 6498
rect 16062 6423 16100 6464
rect 16243 6467 16279 6469
rect 16455 6467 16492 6498
rect 16243 6445 16492 6467
rect 16663 6466 16700 6498
rect 16976 6494 17040 6506
rect 17080 6468 17107 6646
rect 18691 6635 18728 6646
rect 18817 6639 18847 7640
rect 18910 7640 19354 7651
rect 18910 7638 19078 7640
rect 18910 7460 18937 7638
rect 18977 7600 19041 7612
rect 19317 7608 19354 7640
rect 19525 7639 19774 7661
rect 20167 7660 20315 7670
rect 20374 7690 20411 7700
rect 20486 7699 20523 7700
rect 20467 7697 20523 7699
rect 20374 7670 20382 7690
rect 20402 7670 20411 7690
rect 20223 7659 20259 7660
rect 19525 7608 19562 7639
rect 19738 7637 19774 7639
rect 19738 7608 19775 7637
rect 18977 7599 19012 7600
rect 18954 7594 19012 7599
rect 18954 7574 18957 7594
rect 18977 7580 19012 7594
rect 19032 7580 19041 7600
rect 18977 7572 19041 7580
rect 19003 7571 19041 7572
rect 19004 7570 19041 7571
rect 19107 7604 19143 7605
rect 19215 7604 19251 7605
rect 19107 7596 19251 7604
rect 19107 7576 19115 7596
rect 19135 7577 19167 7596
rect 19190 7577 19223 7596
rect 19135 7576 19223 7577
rect 19243 7576 19251 7596
rect 19107 7570 19251 7576
rect 19317 7600 19355 7608
rect 19423 7604 19459 7605
rect 19317 7580 19326 7600
rect 19346 7580 19355 7600
rect 19317 7571 19355 7580
rect 19374 7597 19459 7604
rect 19374 7577 19381 7597
rect 19402 7596 19459 7597
rect 19402 7577 19431 7596
rect 19374 7576 19431 7577
rect 19451 7576 19459 7596
rect 19317 7570 19354 7571
rect 19374 7570 19459 7576
rect 19525 7600 19563 7608
rect 19636 7604 19672 7605
rect 19525 7580 19534 7600
rect 19554 7580 19563 7600
rect 19525 7571 19563 7580
rect 19587 7596 19672 7604
rect 19587 7576 19644 7596
rect 19664 7576 19672 7596
rect 19525 7570 19562 7571
rect 19587 7570 19672 7576
rect 19738 7600 19776 7608
rect 20071 7600 20108 7601
rect 20374 7600 20411 7670
rect 20436 7690 20523 7697
rect 20436 7687 20494 7690
rect 20436 7667 20441 7687
rect 20462 7670 20494 7687
rect 20514 7670 20523 7690
rect 20462 7667 20523 7670
rect 20436 7660 20523 7667
rect 20582 7690 20619 7700
rect 20582 7670 20590 7690
rect 20610 7670 20619 7690
rect 20436 7659 20467 7660
rect 19738 7580 19747 7600
rect 19767 7580 19776 7600
rect 20070 7599 20411 7600
rect 19738 7571 19776 7580
rect 19995 7594 20411 7599
rect 19995 7574 19998 7594
rect 20018 7574 20411 7594
rect 20582 7599 20619 7670
rect 20649 7699 20680 7752
rect 20987 7750 20997 7768
rect 21015 7750 21026 7768
rect 20987 7741 21024 7750
rect 20699 7699 20736 7700
rect 20649 7690 20736 7699
rect 20649 7670 20707 7690
rect 20727 7670 20736 7690
rect 20649 7660 20736 7670
rect 20795 7690 20832 7700
rect 20795 7670 20803 7690
rect 20823 7670 20832 7690
rect 20990 7675 21027 7679
rect 20649 7659 20680 7660
rect 20795 7599 20832 7670
rect 20582 7575 20832 7599
rect 20988 7669 21027 7675
rect 20988 7651 20999 7669
rect 21017 7651 21027 7669
rect 20988 7642 21027 7651
rect 19738 7570 19775 7571
rect 19161 7549 19197 7570
rect 19587 7549 19618 7570
rect 20374 7551 20411 7574
rect 20988 7564 21023 7642
rect 20985 7554 21023 7564
rect 20374 7550 20544 7551
rect 20985 7550 20995 7554
rect 18994 7545 19094 7549
rect 18994 7541 19056 7545
rect 18994 7515 19001 7541
rect 19027 7519 19056 7541
rect 19082 7519 19094 7545
rect 19027 7515 19094 7519
rect 18994 7512 19094 7515
rect 19162 7512 19197 7549
rect 19259 7546 19618 7549
rect 19259 7541 19481 7546
rect 19259 7517 19272 7541
rect 19296 7522 19481 7541
rect 19505 7522 19618 7546
rect 19296 7517 19618 7522
rect 19259 7513 19618 7517
rect 19685 7541 19834 7549
rect 19685 7521 19696 7541
rect 19716 7521 19834 7541
rect 20374 7536 20995 7550
rect 21013 7536 21023 7554
rect 20374 7530 21023 7536
rect 20374 7529 21022 7530
rect 20985 7527 21022 7529
rect 19685 7514 19834 7521
rect 19685 7513 19726 7514
rect 19009 7460 19046 7461
rect 19105 7460 19142 7461
rect 19161 7460 19197 7512
rect 19216 7460 19253 7461
rect 18909 7451 19047 7460
rect 18909 7431 19018 7451
rect 19038 7431 19047 7451
rect 18909 7424 19047 7431
rect 19105 7451 19253 7460
rect 19105 7431 19114 7451
rect 19134 7431 19224 7451
rect 19244 7431 19253 7451
rect 18909 7422 19005 7424
rect 19105 7421 19253 7431
rect 19312 7451 19349 7461
rect 19424 7460 19461 7461
rect 19405 7458 19461 7460
rect 19312 7431 19320 7451
rect 19340 7431 19349 7451
rect 19161 7420 19197 7421
rect 19009 7361 19046 7362
rect 19312 7361 19349 7431
rect 19374 7451 19461 7458
rect 19374 7448 19432 7451
rect 19374 7428 19379 7448
rect 19400 7431 19432 7448
rect 19452 7431 19461 7451
rect 19400 7428 19461 7431
rect 19374 7421 19461 7428
rect 19520 7451 19557 7461
rect 19520 7431 19528 7451
rect 19548 7431 19557 7451
rect 19374 7420 19405 7421
rect 19008 7360 19349 7361
rect 18933 7355 19349 7360
rect 18933 7335 18936 7355
rect 18956 7335 19349 7355
rect 19520 7360 19557 7431
rect 19587 7460 19618 7513
rect 19637 7460 19674 7461
rect 19587 7451 19674 7460
rect 19587 7431 19645 7451
rect 19665 7431 19674 7451
rect 19587 7421 19674 7431
rect 19733 7451 19770 7461
rect 19733 7431 19741 7451
rect 19761 7431 19770 7451
rect 19587 7420 19618 7421
rect 19733 7360 19770 7431
rect 20988 7455 21025 7465
rect 20988 7437 20997 7455
rect 21015 7437 21025 7455
rect 20988 7428 21025 7437
rect 20988 7404 21023 7428
rect 20986 7380 21023 7404
rect 20985 7374 21023 7380
rect 19520 7336 19770 7360
rect 20396 7356 21023 7374
rect 19978 7339 20146 7340
rect 20397 7339 20421 7356
rect 19978 7313 20422 7339
rect 19978 7311 20146 7313
rect 19978 7133 20005 7311
rect 20045 7273 20109 7285
rect 20385 7281 20422 7313
rect 20593 7312 20842 7334
rect 20593 7281 20630 7312
rect 20806 7310 20842 7312
rect 20985 7315 21023 7356
rect 20806 7281 20843 7310
rect 20045 7272 20080 7273
rect 20022 7267 20080 7272
rect 20022 7247 20025 7267
rect 20045 7253 20080 7267
rect 20100 7253 20109 7273
rect 20045 7245 20109 7253
rect 20071 7244 20109 7245
rect 20072 7243 20109 7244
rect 20175 7277 20211 7278
rect 20283 7277 20319 7278
rect 20175 7271 20319 7277
rect 20175 7269 20241 7271
rect 20175 7249 20183 7269
rect 20203 7250 20241 7269
rect 20263 7269 20319 7271
rect 20263 7250 20291 7269
rect 20203 7249 20291 7250
rect 20311 7249 20319 7269
rect 20175 7243 20319 7249
rect 20385 7273 20423 7281
rect 20491 7277 20527 7278
rect 20385 7253 20394 7273
rect 20414 7253 20423 7273
rect 20385 7244 20423 7253
rect 20442 7270 20527 7277
rect 20442 7250 20449 7270
rect 20470 7269 20527 7270
rect 20470 7250 20499 7269
rect 20442 7249 20499 7250
rect 20519 7249 20527 7269
rect 20385 7243 20422 7244
rect 20442 7243 20527 7249
rect 20593 7273 20631 7281
rect 20704 7277 20740 7278
rect 20593 7253 20602 7273
rect 20622 7253 20631 7273
rect 20593 7244 20631 7253
rect 20655 7269 20740 7277
rect 20655 7249 20712 7269
rect 20732 7249 20740 7269
rect 20593 7243 20630 7244
rect 20655 7243 20740 7249
rect 20806 7273 20844 7281
rect 20806 7253 20815 7273
rect 20835 7253 20844 7273
rect 20806 7244 20844 7253
rect 20985 7280 21021 7315
rect 20985 7270 21022 7280
rect 20985 7252 20995 7270
rect 21013 7252 21022 7270
rect 20806 7243 20843 7244
rect 20985 7243 21022 7252
rect 20229 7222 20265 7243
rect 20655 7222 20686 7243
rect 20062 7218 20162 7222
rect 20062 7214 20124 7218
rect 20062 7188 20069 7214
rect 20095 7192 20124 7214
rect 20150 7192 20162 7218
rect 20095 7188 20162 7192
rect 20062 7185 20162 7188
rect 20230 7185 20265 7222
rect 20327 7219 20686 7222
rect 20327 7214 20549 7219
rect 20327 7190 20340 7214
rect 20364 7195 20549 7214
rect 20573 7195 20686 7219
rect 20364 7190 20686 7195
rect 20327 7186 20686 7190
rect 20753 7214 20902 7222
rect 20753 7194 20764 7214
rect 20784 7194 20902 7214
rect 20753 7187 20902 7194
rect 20753 7186 20794 7187
rect 20077 7133 20114 7134
rect 20173 7133 20210 7134
rect 20229 7133 20265 7185
rect 20284 7133 20321 7134
rect 19977 7124 20115 7133
rect 18965 7105 19133 7106
rect 18965 7102 19409 7105
rect 18965 7083 19340 7102
rect 19360 7083 19409 7102
rect 19977 7104 20086 7124
rect 20106 7104 20115 7124
rect 18965 7079 19409 7083
rect 18965 7077 19133 7079
rect 18965 6899 18992 7077
rect 19032 7039 19096 7051
rect 19372 7047 19409 7079
rect 19580 7078 19829 7100
rect 19977 7097 20115 7104
rect 20173 7124 20321 7133
rect 20173 7104 20182 7124
rect 20202 7104 20292 7124
rect 20312 7104 20321 7124
rect 19977 7095 20073 7097
rect 20173 7094 20321 7104
rect 20380 7124 20417 7134
rect 20492 7133 20529 7134
rect 20473 7131 20529 7133
rect 20380 7104 20388 7124
rect 20408 7104 20417 7124
rect 20229 7093 20265 7094
rect 19580 7047 19617 7078
rect 19793 7076 19829 7078
rect 19793 7047 19830 7076
rect 19032 7038 19067 7039
rect 19009 7033 19067 7038
rect 19009 7013 19012 7033
rect 19032 7019 19067 7033
rect 19087 7019 19096 7039
rect 19032 7011 19096 7019
rect 19058 7010 19096 7011
rect 19059 7009 19096 7010
rect 19162 7043 19198 7044
rect 19270 7043 19306 7044
rect 19162 7035 19306 7043
rect 19162 7015 19170 7035
rect 19190 7015 19222 7035
rect 19246 7015 19278 7035
rect 19298 7015 19306 7035
rect 19162 7009 19306 7015
rect 19372 7039 19410 7047
rect 19478 7043 19514 7044
rect 19372 7019 19381 7039
rect 19401 7019 19410 7039
rect 19372 7010 19410 7019
rect 19429 7036 19514 7043
rect 19429 7016 19436 7036
rect 19457 7035 19514 7036
rect 19457 7016 19486 7035
rect 19429 7015 19486 7016
rect 19506 7015 19514 7035
rect 19372 7009 19409 7010
rect 19429 7009 19514 7015
rect 19580 7039 19618 7047
rect 19691 7043 19727 7044
rect 19580 7019 19589 7039
rect 19609 7019 19618 7039
rect 19580 7010 19618 7019
rect 19642 7035 19727 7043
rect 19642 7015 19699 7035
rect 19719 7015 19727 7035
rect 19580 7009 19617 7010
rect 19642 7009 19727 7015
rect 19793 7039 19831 7047
rect 19793 7019 19802 7039
rect 19822 7019 19831 7039
rect 20077 7034 20114 7035
rect 20380 7034 20417 7104
rect 20442 7124 20529 7131
rect 20442 7121 20500 7124
rect 20442 7101 20447 7121
rect 20468 7104 20500 7121
rect 20520 7104 20529 7124
rect 20468 7101 20529 7104
rect 20442 7094 20529 7101
rect 20588 7124 20625 7134
rect 20588 7104 20596 7124
rect 20616 7104 20625 7124
rect 20442 7093 20473 7094
rect 20076 7033 20417 7034
rect 19793 7010 19831 7019
rect 20001 7028 20417 7033
rect 19793 7009 19830 7010
rect 19216 6988 19252 7009
rect 19642 6988 19673 7009
rect 20001 7008 20004 7028
rect 20024 7008 20417 7028
rect 20588 7033 20625 7104
rect 20655 7133 20686 7186
rect 20988 7171 21025 7181
rect 20988 7153 20997 7171
rect 21015 7153 21025 7171
rect 20988 7144 21025 7153
rect 20705 7133 20742 7134
rect 20655 7124 20742 7133
rect 20655 7104 20713 7124
rect 20733 7104 20742 7124
rect 20655 7094 20742 7104
rect 20801 7124 20838 7134
rect 20801 7104 20809 7124
rect 20829 7104 20838 7124
rect 20655 7093 20686 7094
rect 20801 7033 20838 7104
rect 20993 7079 21024 7144
rect 20992 7069 21029 7079
rect 20992 7067 21002 7069
rect 20926 7065 21002 7067
rect 20588 7009 20838 7033
rect 20923 7051 21002 7065
rect 21020 7051 21029 7069
rect 20923 7048 21029 7051
rect 20395 6989 20416 7008
rect 20923 6989 20949 7048
rect 20992 7042 21029 7048
rect 19049 6984 19149 6988
rect 19049 6980 19111 6984
rect 19049 6954 19056 6980
rect 19082 6958 19111 6980
rect 19137 6958 19149 6984
rect 19082 6954 19149 6958
rect 19049 6951 19149 6954
rect 19217 6951 19252 6988
rect 19314 6985 19673 6988
rect 19314 6980 19536 6985
rect 19314 6956 19327 6980
rect 19351 6961 19536 6980
rect 19560 6961 19673 6985
rect 19351 6956 19673 6961
rect 19314 6952 19673 6956
rect 19740 6980 19889 6988
rect 19740 6960 19751 6980
rect 19771 6960 19889 6980
rect 20395 6971 20949 6989
rect 20995 6978 21032 6980
rect 20923 6970 20949 6971
rect 20992 6970 21032 6978
rect 19740 6953 19889 6960
rect 20992 6958 21004 6970
rect 20983 6953 21004 6958
rect 19740 6952 19781 6953
rect 20399 6952 21004 6953
rect 21022 6952 21032 6970
rect 19064 6899 19101 6900
rect 19160 6899 19197 6900
rect 19216 6899 19252 6951
rect 19271 6899 19308 6900
rect 18964 6890 19102 6899
rect 18964 6870 19073 6890
rect 19093 6870 19102 6890
rect 18964 6863 19102 6870
rect 19160 6890 19308 6899
rect 19160 6870 19169 6890
rect 19189 6870 19279 6890
rect 19299 6870 19308 6890
rect 18964 6861 19060 6863
rect 19160 6860 19308 6870
rect 19367 6890 19404 6900
rect 19479 6899 19516 6900
rect 19460 6897 19516 6899
rect 19367 6870 19375 6890
rect 19395 6870 19404 6890
rect 19216 6859 19252 6860
rect 19064 6800 19101 6801
rect 19367 6800 19404 6870
rect 19429 6890 19516 6897
rect 19429 6887 19487 6890
rect 19429 6867 19434 6887
rect 19455 6870 19487 6887
rect 19507 6870 19516 6890
rect 19455 6867 19516 6870
rect 19429 6860 19516 6867
rect 19575 6890 19612 6900
rect 19575 6870 19583 6890
rect 19603 6870 19612 6890
rect 19429 6859 19460 6860
rect 19063 6799 19404 6800
rect 18988 6794 19404 6799
rect 18988 6774 18991 6794
rect 19011 6774 19404 6794
rect 19575 6799 19612 6870
rect 19642 6899 19673 6952
rect 20399 6943 21032 6952
rect 20399 6936 21031 6943
rect 20399 6934 20461 6936
rect 19977 6924 20145 6925
rect 20399 6924 20421 6934
rect 19692 6899 19729 6900
rect 19642 6890 19729 6899
rect 19642 6870 19700 6890
rect 19720 6870 19729 6890
rect 19642 6860 19729 6870
rect 19788 6890 19825 6900
rect 19788 6870 19796 6890
rect 19816 6870 19825 6890
rect 19642 6859 19673 6860
rect 19788 6799 19825 6870
rect 19575 6775 19825 6799
rect 19977 6898 20421 6924
rect 19977 6896 20145 6898
rect 19977 6718 20004 6896
rect 20044 6858 20108 6870
rect 20384 6866 20421 6898
rect 20592 6897 20841 6919
rect 20592 6866 20629 6897
rect 20805 6895 20841 6897
rect 20805 6866 20842 6895
rect 20044 6857 20079 6858
rect 20021 6852 20079 6857
rect 20021 6832 20024 6852
rect 20044 6838 20079 6852
rect 20099 6838 20108 6858
rect 20044 6830 20108 6838
rect 20070 6829 20108 6830
rect 20071 6828 20108 6829
rect 20174 6862 20210 6863
rect 20282 6862 20318 6863
rect 20174 6854 20318 6862
rect 20174 6834 20182 6854
rect 20202 6834 20231 6854
rect 20174 6833 20231 6834
rect 20253 6834 20290 6854
rect 20310 6834 20318 6854
rect 20253 6833 20318 6834
rect 20174 6828 20318 6833
rect 20384 6858 20422 6866
rect 20490 6862 20526 6863
rect 20384 6838 20393 6858
rect 20413 6838 20422 6858
rect 20384 6829 20422 6838
rect 20441 6855 20526 6862
rect 20441 6835 20448 6855
rect 20469 6854 20526 6855
rect 20469 6835 20498 6854
rect 20441 6834 20498 6835
rect 20518 6834 20526 6854
rect 20384 6828 20421 6829
rect 20441 6828 20526 6834
rect 20592 6858 20630 6866
rect 20703 6862 20739 6863
rect 20592 6838 20601 6858
rect 20621 6838 20630 6858
rect 20592 6829 20630 6838
rect 20654 6854 20739 6862
rect 20654 6834 20711 6854
rect 20731 6834 20739 6854
rect 20592 6828 20629 6829
rect 20654 6828 20739 6834
rect 20805 6858 20843 6866
rect 20805 6838 20814 6858
rect 20834 6838 20843 6858
rect 20805 6829 20843 6838
rect 20805 6828 20842 6829
rect 20228 6807 20264 6828
rect 20654 6807 20685 6828
rect 20061 6803 20161 6807
rect 20061 6799 20123 6803
rect 20061 6773 20068 6799
rect 20094 6777 20123 6799
rect 20149 6777 20161 6803
rect 20094 6773 20161 6777
rect 20061 6770 20161 6773
rect 20229 6770 20264 6807
rect 20326 6804 20685 6807
rect 20326 6799 20548 6804
rect 20326 6775 20339 6799
rect 20363 6780 20548 6799
rect 20572 6780 20685 6804
rect 20363 6775 20685 6780
rect 20326 6771 20685 6775
rect 20752 6799 20901 6807
rect 20752 6779 20763 6799
rect 20783 6779 20901 6799
rect 20752 6772 20901 6779
rect 20992 6787 21031 6936
rect 20752 6771 20793 6772
rect 20076 6718 20113 6719
rect 20172 6718 20209 6719
rect 20228 6718 20264 6770
rect 20283 6718 20320 6719
rect 19976 6709 20114 6718
rect 19976 6689 20085 6709
rect 20105 6689 20114 6709
rect 19976 6682 20114 6689
rect 20172 6709 20320 6718
rect 20172 6689 20181 6709
rect 20201 6689 20291 6709
rect 20311 6689 20320 6709
rect 19976 6680 20072 6682
rect 20172 6679 20320 6689
rect 20379 6709 20416 6719
rect 20491 6718 20528 6719
rect 20472 6716 20528 6718
rect 20379 6689 20387 6709
rect 20407 6689 20416 6709
rect 20228 6678 20264 6679
rect 18691 6616 18699 6635
rect 18722 6616 18728 6635
rect 18691 6605 18728 6616
rect 18757 6638 18925 6639
rect 18757 6612 19201 6638
rect 18757 6610 18925 6612
rect 18694 6545 18727 6605
rect 16939 6466 17107 6468
rect 16663 6440 17107 6466
rect 16664 6423 16688 6440
rect 16939 6439 17107 6440
rect 17475 6468 17725 6492
rect 15711 6416 15749 6422
rect 15122 6398 15749 6416
rect 16062 6405 16689 6423
rect 16062 6399 16100 6405
rect 14086 6329 14336 6353
rect 14704 6381 14872 6382
rect 15123 6381 15147 6398
rect 14704 6355 15148 6381
rect 14704 6353 14872 6355
rect 14704 6175 14731 6353
rect 14771 6315 14835 6327
rect 15111 6323 15148 6355
rect 15319 6354 15568 6376
rect 15319 6323 15356 6354
rect 15532 6352 15568 6354
rect 15711 6357 15749 6398
rect 15532 6323 15569 6352
rect 14771 6314 14806 6315
rect 14748 6309 14806 6314
rect 14748 6289 14751 6309
rect 14771 6295 14806 6309
rect 14826 6295 14835 6315
rect 14771 6287 14835 6295
rect 14797 6286 14835 6287
rect 14798 6285 14835 6286
rect 14901 6319 14937 6320
rect 15009 6319 15045 6320
rect 14901 6313 15045 6319
rect 14901 6311 14967 6313
rect 14901 6291 14909 6311
rect 14929 6292 14967 6311
rect 14989 6311 15045 6313
rect 14989 6292 15017 6311
rect 14929 6291 15017 6292
rect 15037 6291 15045 6311
rect 14901 6285 15045 6291
rect 15111 6315 15149 6323
rect 15217 6319 15253 6320
rect 15111 6295 15120 6315
rect 15140 6295 15149 6315
rect 15111 6286 15149 6295
rect 15168 6312 15253 6319
rect 15168 6292 15175 6312
rect 15196 6311 15253 6312
rect 15196 6292 15225 6311
rect 15168 6291 15225 6292
rect 15245 6291 15253 6311
rect 15111 6285 15148 6286
rect 15168 6285 15253 6291
rect 15319 6315 15357 6323
rect 15430 6319 15466 6320
rect 15319 6295 15328 6315
rect 15348 6295 15357 6315
rect 15319 6286 15357 6295
rect 15381 6311 15466 6319
rect 15381 6291 15438 6311
rect 15458 6291 15466 6311
rect 15319 6285 15356 6286
rect 15381 6285 15466 6291
rect 15532 6315 15570 6323
rect 15532 6295 15541 6315
rect 15561 6295 15570 6315
rect 15532 6286 15570 6295
rect 15711 6322 15747 6357
rect 16064 6353 16099 6399
rect 17475 6397 17512 6468
rect 17627 6407 17658 6408
rect 17475 6377 17484 6397
rect 17504 6377 17512 6397
rect 17475 6367 17512 6377
rect 17571 6397 17658 6407
rect 17571 6377 17580 6397
rect 17600 6377 17658 6397
rect 17571 6368 17658 6377
rect 17571 6367 17608 6368
rect 16062 6344 16099 6353
rect 16062 6326 16072 6344
rect 16090 6326 16099 6344
rect 15711 6312 15748 6322
rect 16062 6316 16099 6326
rect 17627 6315 17658 6368
rect 17688 6397 17725 6468
rect 17896 6473 18289 6493
rect 18309 6473 18312 6493
rect 17896 6468 18312 6473
rect 17896 6467 18237 6468
rect 17840 6407 17871 6408
rect 17688 6377 17697 6397
rect 17717 6377 17725 6397
rect 17688 6367 17725 6377
rect 17784 6400 17871 6407
rect 17784 6397 17845 6400
rect 17784 6377 17793 6397
rect 17813 6380 17845 6397
rect 17866 6380 17871 6400
rect 17813 6377 17871 6380
rect 17784 6370 17871 6377
rect 17896 6397 17933 6467
rect 18199 6466 18236 6467
rect 18048 6407 18084 6408
rect 17896 6377 17905 6397
rect 17925 6377 17933 6397
rect 17784 6368 17840 6370
rect 17784 6367 17821 6368
rect 17896 6367 17933 6377
rect 17992 6397 18140 6407
rect 18240 6404 18336 6406
rect 17992 6377 18001 6397
rect 18021 6377 18111 6397
rect 18131 6377 18140 6397
rect 17992 6368 18140 6377
rect 18198 6397 18336 6404
rect 18198 6377 18207 6397
rect 18227 6377 18336 6397
rect 18198 6368 18336 6377
rect 17992 6367 18029 6368
rect 18048 6316 18084 6368
rect 18103 6367 18140 6368
rect 18199 6367 18236 6368
rect 17519 6314 17560 6315
rect 15711 6294 15721 6312
rect 15739 6294 15748 6312
rect 15532 6285 15569 6286
rect 15711 6285 15748 6294
rect 17411 6307 17560 6314
rect 17411 6287 17529 6307
rect 17549 6287 17560 6307
rect 14955 6264 14991 6285
rect 15381 6264 15412 6285
rect 17411 6279 17560 6287
rect 17627 6311 17986 6315
rect 17627 6306 17949 6311
rect 17627 6282 17740 6306
rect 17764 6287 17949 6306
rect 17973 6287 17986 6311
rect 17764 6282 17986 6287
rect 17627 6279 17986 6282
rect 18048 6279 18083 6316
rect 18151 6313 18251 6316
rect 18151 6309 18218 6313
rect 18151 6283 18163 6309
rect 18189 6287 18218 6309
rect 18244 6287 18251 6313
rect 18189 6283 18251 6287
rect 18151 6279 18251 6283
rect 14788 6260 14888 6264
rect 14788 6256 14850 6260
rect 14788 6230 14795 6256
rect 14821 6234 14850 6256
rect 14876 6234 14888 6260
rect 14821 6230 14888 6234
rect 14788 6227 14888 6230
rect 14956 6227 14991 6264
rect 15053 6261 15412 6264
rect 15053 6256 15275 6261
rect 15053 6232 15066 6256
rect 15090 6237 15275 6256
rect 15299 6237 15412 6261
rect 15090 6232 15412 6237
rect 15053 6228 15412 6232
rect 15479 6256 15628 6264
rect 17627 6258 17658 6279
rect 18048 6258 18084 6279
rect 17470 6257 17507 6258
rect 15479 6236 15490 6256
rect 15510 6236 15628 6256
rect 16065 6252 16102 6254
rect 16065 6251 16713 6252
rect 15479 6229 15628 6236
rect 16064 6245 16713 6251
rect 15479 6228 15520 6229
rect 14803 6175 14840 6176
rect 14899 6175 14936 6176
rect 14955 6175 14991 6227
rect 15010 6175 15047 6176
rect 14703 6166 14841 6175
rect 13639 6148 13670 6151
rect 13639 6122 13646 6148
rect 13665 6122 13670 6148
rect 13639 5728 13670 6122
rect 13691 6147 13859 6148
rect 13691 6144 14135 6147
rect 13691 6125 14066 6144
rect 14086 6125 14135 6144
rect 14703 6146 14812 6166
rect 14832 6146 14841 6166
rect 13691 6121 14135 6125
rect 13691 6119 13859 6121
rect 13691 5941 13718 6119
rect 13758 6081 13822 6093
rect 14098 6089 14135 6121
rect 14306 6120 14555 6142
rect 14703 6139 14841 6146
rect 14899 6166 15047 6175
rect 14899 6146 14908 6166
rect 14928 6146 15018 6166
rect 15038 6146 15047 6166
rect 14703 6137 14799 6139
rect 14899 6136 15047 6146
rect 15106 6166 15143 6176
rect 15218 6175 15255 6176
rect 15199 6173 15255 6175
rect 15106 6146 15114 6166
rect 15134 6146 15143 6166
rect 14955 6135 14991 6136
rect 14306 6089 14343 6120
rect 14519 6118 14555 6120
rect 14519 6089 14556 6118
rect 13758 6080 13793 6081
rect 13735 6075 13793 6080
rect 13735 6055 13738 6075
rect 13758 6061 13793 6075
rect 13813 6061 13822 6081
rect 13758 6053 13822 6061
rect 13784 6052 13822 6053
rect 13785 6051 13822 6052
rect 13888 6085 13924 6086
rect 13996 6085 14032 6086
rect 13888 6077 14032 6085
rect 13888 6057 13896 6077
rect 13916 6076 14004 6077
rect 13916 6057 13949 6076
rect 13888 6056 13949 6057
rect 13973 6057 14004 6076
rect 14024 6057 14032 6077
rect 13973 6056 14032 6057
rect 13888 6051 14032 6056
rect 14098 6081 14136 6089
rect 14204 6085 14240 6086
rect 14098 6061 14107 6081
rect 14127 6061 14136 6081
rect 14098 6052 14136 6061
rect 14155 6078 14240 6085
rect 14155 6058 14162 6078
rect 14183 6077 14240 6078
rect 14183 6058 14212 6077
rect 14155 6057 14212 6058
rect 14232 6057 14240 6077
rect 14098 6051 14135 6052
rect 14155 6051 14240 6057
rect 14306 6081 14344 6089
rect 14417 6085 14453 6086
rect 14306 6061 14315 6081
rect 14335 6061 14344 6081
rect 14306 6052 14344 6061
rect 14368 6077 14453 6085
rect 14368 6057 14425 6077
rect 14445 6057 14453 6077
rect 14306 6051 14343 6052
rect 14368 6051 14453 6057
rect 14519 6081 14557 6089
rect 14519 6061 14528 6081
rect 14548 6061 14557 6081
rect 14803 6076 14840 6077
rect 15106 6076 15143 6146
rect 15168 6166 15255 6173
rect 15168 6163 15226 6166
rect 15168 6143 15173 6163
rect 15194 6146 15226 6163
rect 15246 6146 15255 6166
rect 15194 6143 15255 6146
rect 15168 6136 15255 6143
rect 15314 6166 15351 6176
rect 15314 6146 15322 6166
rect 15342 6146 15351 6166
rect 15168 6135 15199 6136
rect 14802 6075 15143 6076
rect 14519 6052 14557 6061
rect 14727 6070 15143 6075
rect 14519 6051 14556 6052
rect 13942 6030 13978 6051
rect 14368 6030 14399 6051
rect 14727 6050 14730 6070
rect 14750 6050 15143 6070
rect 15314 6075 15351 6146
rect 15381 6175 15412 6228
rect 16064 6227 16074 6245
rect 16092 6231 16713 6245
rect 16092 6227 16102 6231
rect 16543 6230 16713 6231
rect 15714 6213 15751 6223
rect 15714 6195 15723 6213
rect 15741 6195 15751 6213
rect 15714 6186 15751 6195
rect 16064 6217 16102 6227
rect 15431 6175 15468 6176
rect 15381 6166 15468 6175
rect 15381 6146 15439 6166
rect 15459 6146 15468 6166
rect 15381 6136 15468 6146
rect 15527 6166 15564 6176
rect 15527 6146 15535 6166
rect 15555 6146 15564 6166
rect 15381 6135 15412 6136
rect 15527 6075 15564 6146
rect 15719 6121 15750 6186
rect 16064 6139 16099 6217
rect 16676 6207 16713 6230
rect 17469 6248 17507 6257
rect 17469 6228 17478 6248
rect 17498 6228 17507 6248
rect 17469 6220 17507 6228
rect 17573 6252 17658 6258
rect 17683 6257 17720 6258
rect 17573 6232 17581 6252
rect 17601 6232 17658 6252
rect 17573 6224 17658 6232
rect 17682 6248 17720 6257
rect 17682 6228 17691 6248
rect 17711 6228 17720 6248
rect 17573 6223 17609 6224
rect 17682 6220 17720 6228
rect 17786 6252 17871 6258
rect 17891 6257 17928 6258
rect 17786 6232 17794 6252
rect 17814 6251 17871 6252
rect 17814 6232 17843 6251
rect 17786 6231 17843 6232
rect 17864 6231 17871 6251
rect 17786 6224 17871 6231
rect 17890 6248 17928 6257
rect 17890 6228 17899 6248
rect 17919 6228 17928 6248
rect 17786 6223 17822 6224
rect 17890 6220 17928 6228
rect 17994 6256 18138 6258
rect 17994 6252 18052 6256
rect 17994 6232 18002 6252
rect 18022 6232 18052 6252
rect 17994 6230 18052 6232
rect 18077 6252 18138 6256
rect 18077 6232 18110 6252
rect 18130 6232 18138 6252
rect 18077 6230 18138 6232
rect 17994 6224 18138 6230
rect 17994 6223 18030 6224
rect 18102 6223 18138 6224
rect 18204 6257 18241 6258
rect 18204 6256 18242 6257
rect 18204 6248 18268 6256
rect 18204 6228 18213 6248
rect 18233 6234 18268 6248
rect 18288 6234 18291 6254
rect 18233 6229 18291 6234
rect 18233 6228 18268 6229
rect 16060 6130 16099 6139
rect 15718 6111 15755 6121
rect 15718 6109 15728 6111
rect 15652 6107 15728 6109
rect 15314 6051 15564 6075
rect 15649 6093 15728 6107
rect 15746 6093 15755 6111
rect 16060 6112 16070 6130
rect 16088 6112 16099 6130
rect 16060 6106 16099 6112
rect 16255 6182 16505 6206
rect 16255 6111 16292 6182
rect 16407 6121 16438 6122
rect 16060 6102 16097 6106
rect 15649 6090 15755 6093
rect 15121 6031 15142 6050
rect 15649 6031 15675 6090
rect 15718 6084 15755 6090
rect 16255 6091 16264 6111
rect 16284 6091 16292 6111
rect 16255 6081 16292 6091
rect 16351 6111 16438 6121
rect 16351 6091 16360 6111
rect 16380 6091 16438 6111
rect 16351 6082 16438 6091
rect 16351 6081 16388 6082
rect 16063 6031 16100 6040
rect 13775 6026 13875 6030
rect 13775 6022 13837 6026
rect 13775 5996 13782 6022
rect 13808 6000 13837 6022
rect 13863 6000 13875 6026
rect 13808 5996 13875 6000
rect 13775 5993 13875 5996
rect 13943 5993 13978 6030
rect 14040 6027 14399 6030
rect 14040 6022 14262 6027
rect 14040 5998 14053 6022
rect 14077 6003 14262 6022
rect 14286 6003 14399 6027
rect 14077 5998 14399 6003
rect 14040 5994 14399 5998
rect 14466 6022 14615 6030
rect 14466 6002 14477 6022
rect 14497 6002 14615 6022
rect 15121 6013 15675 6031
rect 15721 6020 15758 6022
rect 15649 6012 15675 6013
rect 15718 6012 15758 6020
rect 14466 5995 14615 6002
rect 15718 6000 15730 6012
rect 15709 5995 15730 6000
rect 14466 5994 14507 5995
rect 15125 5994 15730 5995
rect 15748 5994 15758 6012
rect 13790 5941 13827 5942
rect 13886 5941 13923 5942
rect 13942 5941 13978 5993
rect 13997 5941 14034 5942
rect 13690 5932 13828 5941
rect 13690 5912 13799 5932
rect 13819 5912 13828 5932
rect 13690 5905 13828 5912
rect 13886 5932 14034 5941
rect 13886 5912 13895 5932
rect 13915 5912 14005 5932
rect 14025 5912 14034 5932
rect 13690 5903 13786 5905
rect 13886 5902 14034 5912
rect 14093 5932 14130 5942
rect 14205 5941 14242 5942
rect 14186 5939 14242 5941
rect 14093 5912 14101 5932
rect 14121 5912 14130 5932
rect 13942 5901 13978 5902
rect 13790 5842 13827 5843
rect 14093 5842 14130 5912
rect 14155 5932 14242 5939
rect 14155 5929 14213 5932
rect 14155 5909 14160 5929
rect 14181 5912 14213 5929
rect 14233 5912 14242 5932
rect 14181 5909 14242 5912
rect 14155 5902 14242 5909
rect 14301 5932 14338 5942
rect 14301 5912 14309 5932
rect 14329 5912 14338 5932
rect 14155 5901 14186 5902
rect 13789 5841 14130 5842
rect 13714 5836 14130 5841
rect 13714 5816 13717 5836
rect 13737 5816 14130 5836
rect 14301 5841 14338 5912
rect 14368 5941 14399 5994
rect 15125 5985 15758 5994
rect 16061 6013 16072 6031
rect 16090 6013 16100 6031
rect 16407 6029 16438 6082
rect 16468 6111 16505 6182
rect 16676 6187 17069 6207
rect 17089 6187 17092 6207
rect 17470 6191 17507 6220
rect 16676 6182 17092 6187
rect 17471 6189 17507 6191
rect 17683 6189 17720 6220
rect 16676 6181 17017 6182
rect 16620 6121 16651 6122
rect 16468 6091 16477 6111
rect 16497 6091 16505 6111
rect 16468 6081 16505 6091
rect 16564 6114 16651 6121
rect 16564 6111 16625 6114
rect 16564 6091 16573 6111
rect 16593 6094 16625 6111
rect 16646 6094 16651 6114
rect 16593 6091 16651 6094
rect 16564 6084 16651 6091
rect 16676 6111 16713 6181
rect 16979 6180 17016 6181
rect 17471 6167 17720 6189
rect 17891 6188 17928 6220
rect 18204 6216 18268 6228
rect 18308 6190 18335 6368
rect 18167 6188 18335 6190
rect 17891 6162 18335 6188
rect 18167 6161 18335 6162
rect 16828 6121 16864 6122
rect 16676 6091 16685 6111
rect 16705 6091 16713 6111
rect 16564 6082 16620 6084
rect 16564 6081 16601 6082
rect 16676 6081 16713 6091
rect 16772 6111 16920 6121
rect 17020 6118 17116 6120
rect 16772 6091 16781 6111
rect 16801 6091 16891 6111
rect 16911 6091 16920 6111
rect 16772 6082 16920 6091
rect 16978 6111 17116 6118
rect 16978 6091 16987 6111
rect 17007 6091 17116 6111
rect 16978 6082 17116 6091
rect 16772 6081 16809 6082
rect 16828 6030 16864 6082
rect 16883 6081 16920 6082
rect 16979 6081 17016 6082
rect 16299 6028 16340 6029
rect 15125 5978 15757 5985
rect 15125 5976 15187 5978
rect 14703 5966 14871 5967
rect 15125 5966 15147 5976
rect 14418 5941 14455 5942
rect 14368 5932 14455 5941
rect 14368 5912 14426 5932
rect 14446 5912 14455 5932
rect 14368 5902 14455 5912
rect 14514 5932 14551 5942
rect 14514 5912 14522 5932
rect 14542 5912 14551 5932
rect 14368 5901 14399 5902
rect 14514 5841 14551 5912
rect 14301 5817 14551 5841
rect 14703 5940 15147 5966
rect 14703 5938 14871 5940
rect 14703 5760 14730 5938
rect 14770 5900 14834 5912
rect 15110 5908 15147 5940
rect 15318 5939 15567 5961
rect 15318 5908 15355 5939
rect 15531 5937 15567 5939
rect 15531 5908 15568 5937
rect 14770 5899 14805 5900
rect 14747 5894 14805 5899
rect 14747 5874 14750 5894
rect 14770 5880 14805 5894
rect 14825 5880 14834 5900
rect 14770 5872 14834 5880
rect 14796 5871 14834 5872
rect 14797 5870 14834 5871
rect 14900 5904 14936 5905
rect 15008 5904 15044 5905
rect 14900 5896 15044 5904
rect 14900 5876 14908 5896
rect 14928 5876 14957 5896
rect 14900 5875 14957 5876
rect 14979 5876 15016 5896
rect 15036 5876 15044 5896
rect 14979 5875 15044 5876
rect 14900 5870 15044 5875
rect 15110 5900 15148 5908
rect 15216 5904 15252 5905
rect 15110 5880 15119 5900
rect 15139 5880 15148 5900
rect 15110 5871 15148 5880
rect 15167 5897 15252 5904
rect 15167 5877 15174 5897
rect 15195 5896 15252 5897
rect 15195 5877 15224 5896
rect 15167 5876 15224 5877
rect 15244 5876 15252 5896
rect 15110 5870 15147 5871
rect 15167 5870 15252 5876
rect 15318 5900 15356 5908
rect 15429 5904 15465 5905
rect 15318 5880 15327 5900
rect 15347 5880 15356 5900
rect 15318 5871 15356 5880
rect 15380 5896 15465 5904
rect 15380 5876 15437 5896
rect 15457 5876 15465 5896
rect 15318 5870 15355 5871
rect 15380 5870 15465 5876
rect 15531 5900 15569 5908
rect 15531 5880 15540 5900
rect 15560 5880 15569 5900
rect 15531 5871 15569 5880
rect 15531 5870 15568 5871
rect 14954 5849 14990 5870
rect 15380 5849 15411 5870
rect 14787 5845 14887 5849
rect 14787 5841 14849 5845
rect 14787 5815 14794 5841
rect 14820 5819 14849 5841
rect 14875 5819 14887 5845
rect 14820 5815 14887 5819
rect 14787 5812 14887 5815
rect 14955 5812 14990 5849
rect 15052 5846 15411 5849
rect 15052 5841 15274 5846
rect 15052 5817 15065 5841
rect 15089 5822 15274 5841
rect 15298 5822 15411 5846
rect 15089 5817 15411 5822
rect 15052 5813 15411 5817
rect 15478 5841 15627 5849
rect 15478 5821 15489 5841
rect 15509 5821 15627 5841
rect 15478 5814 15627 5821
rect 15718 5829 15757 5978
rect 16061 5864 16100 6013
rect 16191 6021 16340 6028
rect 16191 6001 16309 6021
rect 16329 6001 16340 6021
rect 16191 5993 16340 6001
rect 16407 6025 16766 6029
rect 16407 6020 16729 6025
rect 16407 5996 16520 6020
rect 16544 6001 16729 6020
rect 16753 6001 16766 6025
rect 16544 5996 16766 6001
rect 16407 5993 16766 5996
rect 16828 5993 16863 6030
rect 16931 6027 17031 6030
rect 16931 6023 16998 6027
rect 16931 5997 16943 6023
rect 16969 6001 16998 6023
rect 17024 6001 17031 6027
rect 16969 5997 17031 6001
rect 16931 5993 17031 5997
rect 16407 5972 16438 5993
rect 16828 5972 16864 5993
rect 16250 5971 16287 5972
rect 16249 5962 16287 5971
rect 16249 5942 16258 5962
rect 16278 5942 16287 5962
rect 16249 5934 16287 5942
rect 16353 5966 16438 5972
rect 16463 5971 16500 5972
rect 16353 5946 16361 5966
rect 16381 5946 16438 5966
rect 16353 5938 16438 5946
rect 16462 5962 16500 5971
rect 16462 5942 16471 5962
rect 16491 5942 16500 5962
rect 16353 5937 16389 5938
rect 16462 5934 16500 5942
rect 16566 5966 16651 5972
rect 16671 5971 16708 5972
rect 16566 5946 16574 5966
rect 16594 5965 16651 5966
rect 16594 5946 16623 5965
rect 16566 5945 16623 5946
rect 16644 5945 16651 5965
rect 16566 5938 16651 5945
rect 16670 5962 16708 5971
rect 16670 5942 16679 5962
rect 16699 5942 16708 5962
rect 16566 5937 16602 5938
rect 16670 5934 16708 5942
rect 16774 5967 16918 5972
rect 16774 5966 16839 5967
rect 16774 5946 16782 5966
rect 16802 5946 16839 5966
rect 16861 5966 16918 5967
rect 16861 5946 16890 5966
rect 16910 5946 16918 5966
rect 16774 5938 16918 5946
rect 16774 5937 16810 5938
rect 16882 5937 16918 5938
rect 16984 5971 17021 5972
rect 16984 5970 17022 5971
rect 16984 5962 17048 5970
rect 16984 5942 16993 5962
rect 17013 5948 17048 5962
rect 17068 5948 17071 5968
rect 17013 5943 17071 5948
rect 17013 5942 17048 5943
rect 16250 5905 16287 5934
rect 16251 5903 16287 5905
rect 16463 5903 16500 5934
rect 16251 5881 16500 5903
rect 16671 5902 16708 5934
rect 16984 5930 17048 5942
rect 17088 5904 17115 6082
rect 16947 5902 17115 5904
rect 16671 5876 17115 5902
rect 17267 6001 17517 6025
rect 17267 5930 17304 6001
rect 17419 5940 17450 5941
rect 17267 5910 17276 5930
rect 17296 5910 17304 5930
rect 17267 5900 17304 5910
rect 17363 5930 17450 5940
rect 17363 5910 17372 5930
rect 17392 5910 17450 5930
rect 17363 5901 17450 5910
rect 17363 5900 17400 5901
rect 16671 5866 16693 5876
rect 16947 5875 17115 5876
rect 16631 5864 16693 5866
rect 16061 5857 16693 5864
rect 15478 5813 15519 5814
rect 14802 5760 14839 5761
rect 14898 5760 14935 5761
rect 14954 5760 14990 5812
rect 15009 5760 15046 5761
rect 14702 5751 14840 5760
rect 14702 5731 14811 5751
rect 14831 5731 14840 5751
rect 13639 5727 13809 5728
rect 13639 5712 14085 5727
rect 14702 5724 14840 5731
rect 14898 5751 15046 5760
rect 14898 5731 14907 5751
rect 14927 5731 15017 5751
rect 15037 5731 15046 5751
rect 14702 5722 14798 5724
rect 13641 5701 14085 5712
rect 13641 5699 13809 5701
rect 13641 5521 13668 5699
rect 13708 5661 13772 5673
rect 14048 5669 14085 5701
rect 14256 5700 14505 5722
rect 14898 5721 15046 5731
rect 15105 5751 15142 5761
rect 15217 5760 15254 5761
rect 15198 5758 15254 5760
rect 15105 5731 15113 5751
rect 15133 5731 15142 5751
rect 14954 5720 14990 5721
rect 14256 5669 14293 5700
rect 14469 5698 14505 5700
rect 14469 5669 14506 5698
rect 13708 5660 13743 5661
rect 13685 5655 13743 5660
rect 13685 5635 13688 5655
rect 13708 5641 13743 5655
rect 13763 5641 13772 5661
rect 13708 5633 13772 5641
rect 13734 5632 13772 5633
rect 13735 5631 13772 5632
rect 13838 5665 13874 5666
rect 13946 5665 13982 5666
rect 13838 5657 13982 5665
rect 13838 5637 13846 5657
rect 13866 5656 13954 5657
rect 13866 5639 13894 5656
rect 13918 5639 13954 5656
rect 13866 5637 13954 5639
rect 13974 5637 13982 5657
rect 13838 5631 13982 5637
rect 14048 5661 14086 5669
rect 14154 5665 14190 5666
rect 14048 5641 14057 5661
rect 14077 5641 14086 5661
rect 14048 5632 14086 5641
rect 14105 5658 14190 5665
rect 14105 5638 14112 5658
rect 14133 5657 14190 5658
rect 14133 5638 14162 5657
rect 14105 5637 14162 5638
rect 14182 5637 14190 5657
rect 14048 5631 14085 5632
rect 14105 5631 14190 5637
rect 14256 5661 14294 5669
rect 14367 5665 14403 5666
rect 14256 5641 14265 5661
rect 14285 5641 14294 5661
rect 14256 5632 14294 5641
rect 14318 5657 14403 5665
rect 14318 5637 14375 5657
rect 14395 5637 14403 5657
rect 14256 5631 14293 5632
rect 14318 5631 14403 5637
rect 14469 5661 14507 5669
rect 14802 5661 14839 5662
rect 15105 5661 15142 5731
rect 15167 5751 15254 5758
rect 15167 5748 15225 5751
rect 15167 5728 15172 5748
rect 15193 5731 15225 5748
rect 15245 5731 15254 5751
rect 15193 5728 15254 5731
rect 15167 5721 15254 5728
rect 15313 5751 15350 5761
rect 15313 5731 15321 5751
rect 15341 5731 15350 5751
rect 15167 5720 15198 5721
rect 14469 5641 14478 5661
rect 14498 5641 14507 5661
rect 14801 5660 15142 5661
rect 14469 5632 14507 5641
rect 14726 5655 15142 5660
rect 14726 5635 14729 5655
rect 14749 5635 15142 5655
rect 15313 5660 15350 5731
rect 15380 5760 15411 5813
rect 15718 5811 15728 5829
rect 15746 5811 15757 5829
rect 16060 5848 16693 5857
rect 17419 5848 17450 5901
rect 17480 5930 17517 6001
rect 17688 6006 18081 6026
rect 18101 6006 18104 6026
rect 17688 6001 18104 6006
rect 17688 6000 18029 6001
rect 17632 5940 17663 5941
rect 17480 5910 17489 5930
rect 17509 5910 17517 5930
rect 17480 5900 17517 5910
rect 17576 5933 17663 5940
rect 17576 5930 17637 5933
rect 17576 5910 17585 5930
rect 17605 5913 17637 5930
rect 17658 5913 17663 5933
rect 17605 5910 17663 5913
rect 17576 5903 17663 5910
rect 17688 5930 17725 6000
rect 17991 5999 18028 6000
rect 17840 5940 17876 5941
rect 17688 5910 17697 5930
rect 17717 5910 17725 5930
rect 17576 5901 17632 5903
rect 17576 5900 17613 5901
rect 17688 5900 17725 5910
rect 17784 5930 17932 5940
rect 18032 5937 18128 5939
rect 17784 5910 17793 5930
rect 17813 5910 17903 5930
rect 17923 5910 17932 5930
rect 17784 5901 17932 5910
rect 17990 5930 18128 5937
rect 17990 5910 17999 5930
rect 18019 5910 18128 5930
rect 17990 5901 18128 5910
rect 17784 5900 17821 5901
rect 17840 5849 17876 5901
rect 17895 5900 17932 5901
rect 17991 5900 18028 5901
rect 16060 5830 16070 5848
rect 16088 5847 16693 5848
rect 17311 5847 17352 5848
rect 16088 5842 16109 5847
rect 16088 5830 16100 5842
rect 17203 5840 17352 5847
rect 16060 5822 16100 5830
rect 16143 5829 16169 5830
rect 16060 5820 16097 5822
rect 16143 5811 16697 5829
rect 17203 5820 17321 5840
rect 17341 5820 17352 5840
rect 17203 5812 17352 5820
rect 17419 5844 17778 5848
rect 17419 5839 17741 5844
rect 17419 5815 17532 5839
rect 17556 5820 17741 5839
rect 17765 5820 17778 5844
rect 17556 5815 17778 5820
rect 17419 5812 17778 5815
rect 17840 5812 17875 5849
rect 17943 5846 18043 5849
rect 17943 5842 18010 5846
rect 17943 5816 17955 5842
rect 17981 5820 18010 5842
rect 18036 5820 18043 5846
rect 17981 5816 18043 5820
rect 17943 5812 18043 5816
rect 15718 5802 15755 5811
rect 15430 5760 15467 5761
rect 15380 5751 15467 5760
rect 15380 5731 15438 5751
rect 15458 5731 15467 5751
rect 15380 5721 15467 5731
rect 15526 5751 15563 5761
rect 15526 5731 15534 5751
rect 15554 5731 15563 5751
rect 16063 5752 16100 5758
rect 16143 5752 16169 5811
rect 16676 5792 16697 5811
rect 16063 5749 16169 5752
rect 15721 5736 15758 5740
rect 15380 5720 15411 5721
rect 15526 5660 15563 5731
rect 15313 5636 15563 5660
rect 15719 5730 15758 5736
rect 15719 5712 15730 5730
rect 15748 5712 15758 5730
rect 16063 5731 16072 5749
rect 16090 5735 16169 5749
rect 16254 5767 16504 5791
rect 16090 5733 16166 5735
rect 16090 5731 16100 5733
rect 16063 5721 16100 5731
rect 15719 5703 15758 5712
rect 14469 5631 14506 5632
rect 13892 5610 13928 5631
rect 14318 5610 14349 5631
rect 15105 5612 15142 5635
rect 15719 5625 15754 5703
rect 16068 5656 16099 5721
rect 16254 5696 16291 5767
rect 16406 5706 16437 5707
rect 16254 5676 16263 5696
rect 16283 5676 16291 5696
rect 16254 5666 16291 5676
rect 16350 5696 16437 5706
rect 16350 5676 16359 5696
rect 16379 5676 16437 5696
rect 16350 5667 16437 5676
rect 16350 5666 16387 5667
rect 15716 5615 15754 5625
rect 16067 5647 16104 5656
rect 16067 5629 16077 5647
rect 16095 5629 16104 5647
rect 16067 5619 16104 5629
rect 15105 5611 15275 5612
rect 15716 5611 15726 5615
rect 13725 5606 13825 5610
rect 13725 5602 13787 5606
rect 13725 5576 13732 5602
rect 13758 5580 13787 5602
rect 13813 5580 13825 5606
rect 13758 5576 13825 5580
rect 13725 5573 13825 5576
rect 13893 5573 13928 5610
rect 13990 5607 14349 5610
rect 13990 5602 14212 5607
rect 13990 5578 14003 5602
rect 14027 5583 14212 5602
rect 14236 5583 14349 5607
rect 14027 5578 14349 5583
rect 13990 5574 14349 5578
rect 14416 5602 14565 5610
rect 14416 5582 14427 5602
rect 14447 5582 14565 5602
rect 15105 5597 15726 5611
rect 15744 5597 15754 5615
rect 16406 5614 16437 5667
rect 16467 5696 16504 5767
rect 16675 5772 17068 5792
rect 17088 5772 17091 5792
rect 17419 5791 17450 5812
rect 17840 5791 17876 5812
rect 17262 5790 17299 5791
rect 16675 5767 17091 5772
rect 17261 5781 17299 5790
rect 16675 5766 17016 5767
rect 16619 5706 16650 5707
rect 16467 5676 16476 5696
rect 16496 5676 16504 5696
rect 16467 5666 16504 5676
rect 16563 5699 16650 5706
rect 16563 5696 16624 5699
rect 16563 5676 16572 5696
rect 16592 5679 16624 5696
rect 16645 5679 16650 5699
rect 16592 5676 16650 5679
rect 16563 5669 16650 5676
rect 16675 5696 16712 5766
rect 16978 5765 17015 5766
rect 17261 5761 17270 5781
rect 17290 5761 17299 5781
rect 17261 5753 17299 5761
rect 17365 5785 17450 5791
rect 17475 5790 17512 5791
rect 17365 5765 17373 5785
rect 17393 5765 17450 5785
rect 17365 5757 17450 5765
rect 17474 5781 17512 5790
rect 17474 5761 17483 5781
rect 17503 5761 17512 5781
rect 17365 5756 17401 5757
rect 17474 5753 17512 5761
rect 17578 5785 17663 5791
rect 17683 5790 17720 5791
rect 17578 5765 17586 5785
rect 17606 5784 17663 5785
rect 17606 5765 17635 5784
rect 17578 5764 17635 5765
rect 17656 5764 17663 5784
rect 17578 5757 17663 5764
rect 17682 5781 17720 5790
rect 17682 5761 17691 5781
rect 17711 5761 17720 5781
rect 17578 5756 17614 5757
rect 17682 5753 17720 5761
rect 17786 5785 17930 5791
rect 17786 5765 17794 5785
rect 17814 5765 17846 5785
rect 17870 5765 17902 5785
rect 17922 5765 17930 5785
rect 17786 5757 17930 5765
rect 17786 5756 17822 5757
rect 17894 5756 17930 5757
rect 17996 5790 18033 5791
rect 17996 5789 18034 5790
rect 17996 5781 18060 5789
rect 17996 5761 18005 5781
rect 18025 5767 18060 5781
rect 18080 5767 18083 5787
rect 18025 5762 18083 5767
rect 18025 5761 18060 5762
rect 17262 5724 17299 5753
rect 17263 5722 17299 5724
rect 17475 5722 17512 5753
rect 16827 5706 16863 5707
rect 16675 5676 16684 5696
rect 16704 5676 16712 5696
rect 16563 5667 16619 5669
rect 16563 5666 16600 5667
rect 16675 5666 16712 5676
rect 16771 5696 16919 5706
rect 17019 5703 17115 5705
rect 16771 5676 16780 5696
rect 16800 5676 16890 5696
rect 16910 5676 16919 5696
rect 16771 5667 16919 5676
rect 16977 5696 17115 5703
rect 17263 5700 17512 5722
rect 17683 5721 17720 5753
rect 17996 5749 18060 5761
rect 18100 5723 18127 5901
rect 17959 5721 18127 5723
rect 17683 5717 18127 5721
rect 16977 5676 16986 5696
rect 17006 5676 17115 5696
rect 17683 5698 17732 5717
rect 17752 5698 18127 5717
rect 17683 5695 18127 5698
rect 17959 5694 18127 5695
rect 16977 5667 17115 5676
rect 16771 5666 16808 5667
rect 16827 5615 16863 5667
rect 16882 5666 16919 5667
rect 16978 5666 17015 5667
rect 16298 5613 16339 5614
rect 15105 5591 15754 5597
rect 16190 5606 16339 5613
rect 15105 5590 15753 5591
rect 15716 5588 15753 5590
rect 14416 5575 14565 5582
rect 16190 5586 16308 5606
rect 16328 5586 16339 5606
rect 16190 5578 16339 5586
rect 16406 5610 16765 5614
rect 16406 5605 16728 5610
rect 16406 5581 16519 5605
rect 16543 5586 16728 5605
rect 16752 5586 16765 5610
rect 16543 5581 16765 5586
rect 16406 5578 16765 5581
rect 16827 5578 16862 5615
rect 16930 5612 17030 5615
rect 16930 5608 16997 5612
rect 16930 5582 16942 5608
rect 16968 5586 16997 5608
rect 17023 5586 17030 5612
rect 16968 5582 17030 5586
rect 16930 5578 17030 5582
rect 14416 5574 14457 5575
rect 13740 5521 13777 5522
rect 13836 5521 13873 5522
rect 13892 5521 13928 5573
rect 13947 5521 13984 5522
rect 13640 5512 13778 5521
rect 13640 5492 13749 5512
rect 13769 5492 13778 5512
rect 13640 5485 13778 5492
rect 13836 5512 13984 5521
rect 13836 5492 13845 5512
rect 13865 5492 13955 5512
rect 13975 5492 13984 5512
rect 13640 5483 13736 5485
rect 13836 5482 13984 5492
rect 14043 5512 14080 5522
rect 14155 5521 14192 5522
rect 14136 5519 14192 5521
rect 14043 5492 14051 5512
rect 14071 5492 14080 5512
rect 13892 5481 13928 5482
rect 13740 5422 13777 5423
rect 14043 5422 14080 5492
rect 14105 5512 14192 5519
rect 14105 5509 14163 5512
rect 14105 5489 14110 5509
rect 14131 5492 14163 5509
rect 14183 5492 14192 5512
rect 14131 5489 14192 5492
rect 14105 5482 14192 5489
rect 14251 5512 14288 5522
rect 14251 5492 14259 5512
rect 14279 5492 14288 5512
rect 14105 5481 14136 5482
rect 13739 5421 14080 5422
rect 13664 5416 14080 5421
rect 13664 5396 13667 5416
rect 13687 5396 14080 5416
rect 14251 5421 14288 5492
rect 14318 5521 14349 5574
rect 16406 5557 16437 5578
rect 16827 5557 16863 5578
rect 16070 5548 16107 5557
rect 16249 5556 16286 5557
rect 16070 5530 16079 5548
rect 16097 5530 16107 5548
rect 14368 5521 14405 5522
rect 14318 5512 14405 5521
rect 14318 5492 14376 5512
rect 14396 5492 14405 5512
rect 14318 5482 14405 5492
rect 14464 5512 14501 5522
rect 14464 5492 14472 5512
rect 14492 5492 14501 5512
rect 14318 5481 14349 5482
rect 14464 5421 14501 5492
rect 15719 5516 15756 5526
rect 16070 5520 16107 5530
rect 15719 5498 15728 5516
rect 15746 5498 15756 5516
rect 15719 5489 15756 5498
rect 15719 5465 15754 5489
rect 16071 5485 16107 5520
rect 16248 5547 16286 5556
rect 16248 5527 16257 5547
rect 16277 5527 16286 5547
rect 16248 5519 16286 5527
rect 16352 5551 16437 5557
rect 16462 5556 16499 5557
rect 16352 5531 16360 5551
rect 16380 5531 16437 5551
rect 16352 5523 16437 5531
rect 16461 5547 16499 5556
rect 16461 5527 16470 5547
rect 16490 5527 16499 5547
rect 16352 5522 16388 5523
rect 16461 5519 16499 5527
rect 16565 5551 16650 5557
rect 16670 5556 16707 5557
rect 16565 5531 16573 5551
rect 16593 5550 16650 5551
rect 16593 5531 16622 5550
rect 16565 5530 16622 5531
rect 16643 5530 16650 5550
rect 16565 5523 16650 5530
rect 16669 5547 16707 5556
rect 16669 5527 16678 5547
rect 16698 5527 16707 5547
rect 16565 5522 16601 5523
rect 16669 5519 16707 5527
rect 16773 5551 16917 5557
rect 16773 5531 16781 5551
rect 16801 5550 16889 5551
rect 16801 5531 16829 5550
rect 16773 5529 16829 5531
rect 16851 5531 16889 5550
rect 16909 5531 16917 5551
rect 16851 5529 16917 5531
rect 16773 5523 16917 5529
rect 16773 5522 16809 5523
rect 16881 5522 16917 5523
rect 16983 5556 17020 5557
rect 16983 5555 17021 5556
rect 16983 5547 17047 5555
rect 16983 5527 16992 5547
rect 17012 5533 17047 5547
rect 17067 5533 17070 5553
rect 17012 5528 17070 5533
rect 17012 5527 17047 5528
rect 16249 5490 16286 5519
rect 15717 5441 15754 5465
rect 15716 5435 15754 5441
rect 14251 5397 14501 5421
rect 15127 5417 15754 5435
rect 14709 5400 14877 5401
rect 15128 5400 15152 5417
rect 14709 5374 15153 5400
rect 14709 5372 14877 5374
rect 14709 5194 14736 5372
rect 14776 5334 14840 5346
rect 15116 5342 15153 5374
rect 15324 5373 15573 5395
rect 15324 5342 15361 5373
rect 15537 5371 15573 5373
rect 15716 5376 15754 5417
rect 16069 5444 16107 5485
rect 16250 5488 16286 5490
rect 16462 5488 16499 5519
rect 16250 5466 16499 5488
rect 16670 5487 16707 5519
rect 16983 5515 17047 5527
rect 17087 5489 17114 5667
rect 16946 5487 17114 5489
rect 16670 5461 17114 5487
rect 16671 5444 16695 5461
rect 16946 5460 17114 5461
rect 16069 5426 16696 5444
rect 17322 5440 17572 5464
rect 16069 5420 16107 5426
rect 16069 5396 16106 5420
rect 15537 5342 15574 5371
rect 14776 5333 14811 5334
rect 14753 5328 14811 5333
rect 14753 5308 14756 5328
rect 14776 5314 14811 5328
rect 14831 5314 14840 5334
rect 14776 5306 14840 5314
rect 14802 5305 14840 5306
rect 14803 5304 14840 5305
rect 14906 5338 14942 5339
rect 15014 5338 15050 5339
rect 14906 5332 15050 5338
rect 14906 5330 14972 5332
rect 14906 5310 14914 5330
rect 14934 5311 14972 5330
rect 14994 5330 15050 5332
rect 14994 5311 15022 5330
rect 14934 5310 15022 5311
rect 15042 5310 15050 5330
rect 14906 5304 15050 5310
rect 15116 5334 15154 5342
rect 15222 5338 15258 5339
rect 15116 5314 15125 5334
rect 15145 5314 15154 5334
rect 15116 5305 15154 5314
rect 15173 5331 15258 5338
rect 15173 5311 15180 5331
rect 15201 5330 15258 5331
rect 15201 5311 15230 5330
rect 15173 5310 15230 5311
rect 15250 5310 15258 5330
rect 15116 5304 15153 5305
rect 15173 5304 15258 5310
rect 15324 5334 15362 5342
rect 15435 5338 15471 5339
rect 15324 5314 15333 5334
rect 15353 5314 15362 5334
rect 15324 5305 15362 5314
rect 15386 5330 15471 5338
rect 15386 5310 15443 5330
rect 15463 5310 15471 5330
rect 15324 5304 15361 5305
rect 15386 5304 15471 5310
rect 15537 5334 15575 5342
rect 15537 5314 15546 5334
rect 15566 5314 15575 5334
rect 15537 5305 15575 5314
rect 15716 5341 15752 5376
rect 16069 5372 16104 5396
rect 16067 5363 16104 5372
rect 16067 5345 16077 5363
rect 16095 5345 16104 5363
rect 15716 5331 15753 5341
rect 16067 5335 16104 5345
rect 17322 5369 17359 5440
rect 17474 5379 17505 5380
rect 17322 5349 17331 5369
rect 17351 5349 17359 5369
rect 17322 5339 17359 5349
rect 17418 5369 17505 5379
rect 17418 5349 17427 5369
rect 17447 5349 17505 5369
rect 17418 5340 17505 5349
rect 17418 5339 17455 5340
rect 15716 5313 15726 5331
rect 15744 5313 15753 5331
rect 15537 5304 15574 5305
rect 15716 5304 15753 5313
rect 14960 5283 14996 5304
rect 15386 5283 15417 5304
rect 17474 5287 17505 5340
rect 17535 5369 17572 5440
rect 17743 5445 18136 5465
rect 18156 5445 18159 5465
rect 17743 5440 18159 5445
rect 17743 5439 18084 5440
rect 17687 5379 17718 5380
rect 17535 5349 17544 5369
rect 17564 5349 17572 5369
rect 17535 5339 17572 5349
rect 17631 5372 17718 5379
rect 17631 5369 17692 5372
rect 17631 5349 17640 5369
rect 17660 5352 17692 5369
rect 17713 5352 17718 5372
rect 17660 5349 17718 5352
rect 17631 5342 17718 5349
rect 17743 5369 17780 5439
rect 18046 5438 18083 5439
rect 17895 5379 17931 5380
rect 17743 5349 17752 5369
rect 17772 5349 17780 5369
rect 17631 5340 17687 5342
rect 17631 5339 17668 5340
rect 17743 5339 17780 5349
rect 17839 5369 17987 5379
rect 18087 5376 18183 5378
rect 17839 5349 17848 5369
rect 17868 5349 17958 5369
rect 17978 5349 17987 5369
rect 17839 5340 17987 5349
rect 18045 5369 18183 5376
rect 18045 5349 18054 5369
rect 18074 5349 18183 5369
rect 18045 5340 18183 5349
rect 17839 5339 17876 5340
rect 17895 5288 17931 5340
rect 17950 5339 17987 5340
rect 18046 5339 18083 5340
rect 17366 5286 17407 5287
rect 14793 5279 14893 5283
rect 14793 5275 14855 5279
rect 14793 5249 14800 5275
rect 14826 5253 14855 5275
rect 14881 5253 14893 5279
rect 14826 5249 14893 5253
rect 14793 5246 14893 5249
rect 14961 5246 14996 5283
rect 15058 5280 15417 5283
rect 15058 5275 15280 5280
rect 15058 5251 15071 5275
rect 15095 5256 15280 5275
rect 15304 5256 15417 5280
rect 15095 5251 15417 5256
rect 15058 5247 15417 5251
rect 15484 5275 15633 5283
rect 15484 5255 15495 5275
rect 15515 5255 15633 5275
rect 17258 5279 17407 5286
rect 16070 5271 16107 5273
rect 16070 5270 16718 5271
rect 15484 5248 15633 5255
rect 16069 5264 16718 5270
rect 15484 5247 15525 5248
rect 14808 5194 14845 5195
rect 14904 5194 14941 5195
rect 14960 5194 14996 5246
rect 15015 5194 15052 5195
rect 14708 5185 14846 5194
rect 13696 5166 13864 5167
rect 13696 5163 14140 5166
rect 13696 5144 14071 5163
rect 14091 5144 14140 5163
rect 14708 5165 14817 5185
rect 14837 5165 14846 5185
rect 13696 5140 14140 5144
rect 13696 5138 13864 5140
rect 13696 4960 13723 5138
rect 13763 5100 13827 5112
rect 14103 5108 14140 5140
rect 14311 5139 14560 5161
rect 14708 5158 14846 5165
rect 14904 5185 15052 5194
rect 14904 5165 14913 5185
rect 14933 5165 15023 5185
rect 15043 5165 15052 5185
rect 14708 5156 14804 5158
rect 14904 5155 15052 5165
rect 15111 5185 15148 5195
rect 15223 5194 15260 5195
rect 15204 5192 15260 5194
rect 15111 5165 15119 5185
rect 15139 5165 15148 5185
rect 14960 5154 14996 5155
rect 14311 5108 14348 5139
rect 14524 5137 14560 5139
rect 14524 5108 14561 5137
rect 13763 5099 13798 5100
rect 13740 5094 13798 5099
rect 13740 5074 13743 5094
rect 13763 5080 13798 5094
rect 13818 5080 13827 5100
rect 13763 5072 13827 5080
rect 13789 5071 13827 5072
rect 13790 5070 13827 5071
rect 13893 5104 13929 5105
rect 14001 5104 14037 5105
rect 13893 5096 14037 5104
rect 13893 5076 13901 5096
rect 13921 5076 13953 5096
rect 13977 5076 14009 5096
rect 14029 5076 14037 5096
rect 13893 5070 14037 5076
rect 14103 5100 14141 5108
rect 14209 5104 14245 5105
rect 14103 5080 14112 5100
rect 14132 5080 14141 5100
rect 14103 5071 14141 5080
rect 14160 5097 14245 5104
rect 14160 5077 14167 5097
rect 14188 5096 14245 5097
rect 14188 5077 14217 5096
rect 14160 5076 14217 5077
rect 14237 5076 14245 5096
rect 14103 5070 14140 5071
rect 14160 5070 14245 5076
rect 14311 5100 14349 5108
rect 14422 5104 14458 5105
rect 14311 5080 14320 5100
rect 14340 5080 14349 5100
rect 14311 5071 14349 5080
rect 14373 5096 14458 5104
rect 14373 5076 14430 5096
rect 14450 5076 14458 5096
rect 14311 5070 14348 5071
rect 14373 5070 14458 5076
rect 14524 5100 14562 5108
rect 14524 5080 14533 5100
rect 14553 5080 14562 5100
rect 14808 5095 14845 5096
rect 15111 5095 15148 5165
rect 15173 5185 15260 5192
rect 15173 5182 15231 5185
rect 15173 5162 15178 5182
rect 15199 5165 15231 5182
rect 15251 5165 15260 5185
rect 15199 5162 15260 5165
rect 15173 5155 15260 5162
rect 15319 5185 15356 5195
rect 15319 5165 15327 5185
rect 15347 5165 15356 5185
rect 15173 5154 15204 5155
rect 14807 5094 15148 5095
rect 14524 5071 14562 5080
rect 14732 5089 15148 5094
rect 14524 5070 14561 5071
rect 13947 5049 13983 5070
rect 14373 5049 14404 5070
rect 14732 5069 14735 5089
rect 14755 5069 15148 5089
rect 15319 5094 15356 5165
rect 15386 5194 15417 5247
rect 16069 5246 16079 5264
rect 16097 5250 16718 5264
rect 17258 5259 17376 5279
rect 17396 5259 17407 5279
rect 17258 5251 17407 5259
rect 17474 5283 17833 5287
rect 17474 5278 17796 5283
rect 17474 5254 17587 5278
rect 17611 5259 17796 5278
rect 17820 5259 17833 5283
rect 17611 5254 17833 5259
rect 17474 5251 17833 5254
rect 17895 5251 17930 5288
rect 17998 5285 18098 5288
rect 17998 5281 18065 5285
rect 17998 5255 18010 5281
rect 18036 5259 18065 5281
rect 18091 5259 18098 5285
rect 18036 5255 18098 5259
rect 17998 5251 18098 5255
rect 16097 5246 16107 5250
rect 16548 5249 16718 5250
rect 15719 5232 15756 5242
rect 15719 5214 15728 5232
rect 15746 5214 15756 5232
rect 15719 5205 15756 5214
rect 16069 5236 16107 5246
rect 15436 5194 15473 5195
rect 15386 5185 15473 5194
rect 15386 5165 15444 5185
rect 15464 5165 15473 5185
rect 15386 5155 15473 5165
rect 15532 5185 15569 5195
rect 15532 5165 15540 5185
rect 15560 5165 15569 5185
rect 15386 5154 15417 5155
rect 15532 5094 15569 5165
rect 15724 5140 15755 5205
rect 16069 5158 16104 5236
rect 16681 5226 16718 5249
rect 17474 5230 17505 5251
rect 17895 5230 17931 5251
rect 17317 5229 17354 5230
rect 16065 5149 16104 5158
rect 15723 5130 15760 5140
rect 15723 5128 15733 5130
rect 15657 5126 15733 5128
rect 15319 5070 15569 5094
rect 15654 5112 15733 5126
rect 15751 5112 15760 5130
rect 16065 5131 16075 5149
rect 16093 5131 16104 5149
rect 16065 5125 16104 5131
rect 16260 5201 16510 5225
rect 16260 5130 16297 5201
rect 16412 5140 16443 5141
rect 16065 5121 16102 5125
rect 15654 5109 15760 5112
rect 15126 5050 15147 5069
rect 15654 5050 15680 5109
rect 15723 5103 15760 5109
rect 16260 5110 16269 5130
rect 16289 5110 16297 5130
rect 16260 5100 16297 5110
rect 16356 5130 16443 5140
rect 16356 5110 16365 5130
rect 16385 5110 16443 5130
rect 16356 5101 16443 5110
rect 16356 5100 16393 5101
rect 16068 5050 16105 5059
rect 13780 5045 13880 5049
rect 13780 5041 13842 5045
rect 13780 5015 13787 5041
rect 13813 5019 13842 5041
rect 13868 5019 13880 5045
rect 13813 5015 13880 5019
rect 13780 5012 13880 5015
rect 13948 5012 13983 5049
rect 14045 5046 14404 5049
rect 14045 5041 14267 5046
rect 14045 5017 14058 5041
rect 14082 5022 14267 5041
rect 14291 5022 14404 5046
rect 14082 5017 14404 5022
rect 14045 5013 14404 5017
rect 14471 5041 14620 5049
rect 14471 5021 14482 5041
rect 14502 5021 14620 5041
rect 15126 5032 15680 5050
rect 15726 5039 15763 5041
rect 15654 5031 15680 5032
rect 15723 5031 15763 5039
rect 14471 5014 14620 5021
rect 15723 5019 15735 5031
rect 15714 5014 15735 5019
rect 14471 5013 14512 5014
rect 15130 5013 15735 5014
rect 15753 5013 15763 5031
rect 13795 4960 13832 4961
rect 13891 4960 13928 4961
rect 13947 4960 13983 5012
rect 14002 4960 14039 4961
rect 13695 4951 13833 4960
rect 13695 4931 13804 4951
rect 13824 4931 13833 4951
rect 13695 4924 13833 4931
rect 13891 4951 14039 4960
rect 13891 4931 13900 4951
rect 13920 4931 14010 4951
rect 14030 4931 14039 4951
rect 13695 4922 13791 4924
rect 13891 4921 14039 4931
rect 14098 4951 14135 4961
rect 14210 4960 14247 4961
rect 14191 4958 14247 4960
rect 14098 4931 14106 4951
rect 14126 4931 14135 4951
rect 13947 4920 13983 4921
rect 13795 4861 13832 4862
rect 14098 4861 14135 4931
rect 14160 4951 14247 4958
rect 14160 4948 14218 4951
rect 14160 4928 14165 4948
rect 14186 4931 14218 4948
rect 14238 4931 14247 4951
rect 14186 4928 14247 4931
rect 14160 4921 14247 4928
rect 14306 4951 14343 4961
rect 14306 4931 14314 4951
rect 14334 4931 14343 4951
rect 14160 4920 14191 4921
rect 13794 4860 14135 4861
rect 13719 4855 14135 4860
rect 13719 4835 13722 4855
rect 13742 4835 14135 4855
rect 14306 4860 14343 4931
rect 14373 4960 14404 5013
rect 15130 5004 15763 5013
rect 16066 5032 16077 5050
rect 16095 5032 16105 5050
rect 16412 5048 16443 5101
rect 16473 5130 16510 5201
rect 16681 5206 17074 5226
rect 17094 5206 17097 5226
rect 16681 5201 17097 5206
rect 17316 5220 17354 5229
rect 16681 5200 17022 5201
rect 17316 5200 17325 5220
rect 17345 5200 17354 5220
rect 16625 5140 16656 5141
rect 16473 5110 16482 5130
rect 16502 5110 16510 5130
rect 16473 5100 16510 5110
rect 16569 5133 16656 5140
rect 16569 5130 16630 5133
rect 16569 5110 16578 5130
rect 16598 5113 16630 5130
rect 16651 5113 16656 5133
rect 16598 5110 16656 5113
rect 16569 5103 16656 5110
rect 16681 5130 16718 5200
rect 16984 5199 17021 5200
rect 17316 5192 17354 5200
rect 17420 5224 17505 5230
rect 17530 5229 17567 5230
rect 17420 5204 17428 5224
rect 17448 5204 17505 5224
rect 17420 5196 17505 5204
rect 17529 5220 17567 5229
rect 17529 5200 17538 5220
rect 17558 5200 17567 5220
rect 17420 5195 17456 5196
rect 17529 5192 17567 5200
rect 17633 5224 17718 5230
rect 17738 5229 17775 5230
rect 17633 5204 17641 5224
rect 17661 5223 17718 5224
rect 17661 5204 17690 5223
rect 17633 5203 17690 5204
rect 17711 5203 17718 5223
rect 17633 5196 17718 5203
rect 17737 5220 17775 5229
rect 17737 5200 17746 5220
rect 17766 5200 17775 5220
rect 17633 5195 17669 5196
rect 17737 5192 17775 5200
rect 17841 5224 17985 5230
rect 17841 5204 17849 5224
rect 17869 5223 17957 5224
rect 17869 5204 17902 5223
rect 17925 5204 17957 5223
rect 17977 5204 17985 5224
rect 17841 5196 17985 5204
rect 17841 5195 17877 5196
rect 17949 5195 17985 5196
rect 18051 5229 18088 5230
rect 18051 5228 18089 5229
rect 18051 5220 18115 5228
rect 18051 5200 18060 5220
rect 18080 5206 18115 5220
rect 18135 5206 18138 5226
rect 18080 5201 18138 5206
rect 18080 5200 18115 5201
rect 17317 5163 17354 5192
rect 17318 5161 17354 5163
rect 17530 5161 17567 5192
rect 16833 5140 16869 5141
rect 16681 5110 16690 5130
rect 16710 5110 16718 5130
rect 16569 5101 16625 5103
rect 16569 5100 16606 5101
rect 16681 5100 16718 5110
rect 16777 5130 16925 5140
rect 17318 5139 17567 5161
rect 17738 5160 17775 5192
rect 18051 5188 18115 5200
rect 18155 5162 18182 5340
rect 18014 5160 18182 5162
rect 17738 5149 18182 5160
rect 18245 5160 18275 6161
rect 18245 5155 18277 5160
rect 17025 5137 17121 5139
rect 16777 5110 16786 5130
rect 16806 5110 16896 5130
rect 16916 5110 16925 5130
rect 16777 5101 16925 5110
rect 16983 5130 17121 5137
rect 17738 5134 18184 5149
rect 18014 5133 18184 5134
rect 16983 5110 16992 5130
rect 17012 5110 17121 5130
rect 16983 5101 17121 5110
rect 16777 5100 16814 5101
rect 16833 5049 16869 5101
rect 16888 5100 16925 5101
rect 16984 5100 17021 5101
rect 16304 5047 16345 5048
rect 15130 4997 15762 5004
rect 15130 4995 15192 4997
rect 14708 4985 14876 4986
rect 15130 4985 15152 4995
rect 14423 4960 14460 4961
rect 14373 4951 14460 4960
rect 14373 4931 14431 4951
rect 14451 4931 14460 4951
rect 14373 4921 14460 4931
rect 14519 4951 14556 4961
rect 14519 4931 14527 4951
rect 14547 4931 14556 4951
rect 14373 4920 14404 4921
rect 14519 4860 14556 4931
rect 14306 4836 14556 4860
rect 14708 4959 15152 4985
rect 14708 4957 14876 4959
rect 14708 4779 14735 4957
rect 14775 4919 14839 4931
rect 15115 4927 15152 4959
rect 15323 4958 15572 4980
rect 15323 4927 15360 4958
rect 15536 4956 15572 4958
rect 15536 4927 15573 4956
rect 14775 4918 14810 4919
rect 14752 4913 14810 4918
rect 14752 4893 14755 4913
rect 14775 4899 14810 4913
rect 14830 4899 14839 4919
rect 14775 4891 14839 4899
rect 14801 4890 14839 4891
rect 14802 4889 14839 4890
rect 14905 4923 14941 4924
rect 15013 4923 15049 4924
rect 14905 4915 15049 4923
rect 14905 4895 14913 4915
rect 14933 4895 14962 4915
rect 14905 4894 14962 4895
rect 14984 4895 15021 4915
rect 15041 4895 15049 4915
rect 14984 4894 15049 4895
rect 14905 4889 15049 4894
rect 15115 4919 15153 4927
rect 15221 4923 15257 4924
rect 15115 4899 15124 4919
rect 15144 4899 15153 4919
rect 15115 4890 15153 4899
rect 15172 4916 15257 4923
rect 15172 4896 15179 4916
rect 15200 4915 15257 4916
rect 15200 4896 15229 4915
rect 15172 4895 15229 4896
rect 15249 4895 15257 4915
rect 15115 4889 15152 4890
rect 15172 4889 15257 4895
rect 15323 4919 15361 4927
rect 15434 4923 15470 4924
rect 15323 4899 15332 4919
rect 15352 4899 15361 4919
rect 15323 4890 15361 4899
rect 15385 4915 15470 4923
rect 15385 4895 15442 4915
rect 15462 4895 15470 4915
rect 15323 4889 15360 4890
rect 15385 4889 15470 4895
rect 15536 4919 15574 4927
rect 15536 4899 15545 4919
rect 15565 4899 15574 4919
rect 15536 4890 15574 4899
rect 15536 4889 15573 4890
rect 14959 4868 14995 4889
rect 15385 4868 15416 4889
rect 14792 4864 14892 4868
rect 14792 4860 14854 4864
rect 14792 4834 14799 4860
rect 14825 4838 14854 4860
rect 14880 4838 14892 4864
rect 14825 4834 14892 4838
rect 14792 4831 14892 4834
rect 14960 4831 14995 4868
rect 15057 4865 15416 4868
rect 15057 4860 15279 4865
rect 15057 4836 15070 4860
rect 15094 4841 15279 4860
rect 15303 4841 15416 4865
rect 15094 4836 15416 4841
rect 15057 4832 15416 4836
rect 15483 4860 15632 4868
rect 15483 4840 15494 4860
rect 15514 4840 15632 4860
rect 15483 4833 15632 4840
rect 15723 4848 15762 4997
rect 16066 4883 16105 5032
rect 16196 5040 16345 5047
rect 16196 5020 16314 5040
rect 16334 5020 16345 5040
rect 16196 5012 16345 5020
rect 16412 5044 16771 5048
rect 16412 5039 16734 5044
rect 16412 5015 16525 5039
rect 16549 5020 16734 5039
rect 16758 5020 16771 5044
rect 16549 5015 16771 5020
rect 16412 5012 16771 5015
rect 16833 5012 16868 5049
rect 16936 5046 17036 5049
rect 16936 5042 17003 5046
rect 16936 5016 16948 5042
rect 16974 5020 17003 5042
rect 17029 5020 17036 5046
rect 16974 5016 17036 5020
rect 16936 5012 17036 5016
rect 16412 4991 16443 5012
rect 16833 4991 16869 5012
rect 16255 4990 16292 4991
rect 16254 4981 16292 4990
rect 16254 4961 16263 4981
rect 16283 4961 16292 4981
rect 16254 4953 16292 4961
rect 16358 4985 16443 4991
rect 16468 4990 16505 4991
rect 16358 4965 16366 4985
rect 16386 4965 16443 4985
rect 16358 4957 16443 4965
rect 16467 4981 16505 4990
rect 16467 4961 16476 4981
rect 16496 4961 16505 4981
rect 16358 4956 16394 4957
rect 16467 4953 16505 4961
rect 16571 4985 16656 4991
rect 16676 4990 16713 4991
rect 16571 4965 16579 4985
rect 16599 4984 16656 4985
rect 16599 4965 16628 4984
rect 16571 4964 16628 4965
rect 16649 4964 16656 4984
rect 16571 4957 16656 4964
rect 16675 4981 16713 4990
rect 16675 4961 16684 4981
rect 16704 4961 16713 4981
rect 16571 4956 16607 4957
rect 16675 4953 16713 4961
rect 16779 4986 16923 4991
rect 16779 4985 16844 4986
rect 16779 4965 16787 4985
rect 16807 4965 16844 4985
rect 16866 4985 16923 4986
rect 16866 4965 16895 4985
rect 16915 4965 16923 4985
rect 16779 4957 16923 4965
rect 16779 4956 16815 4957
rect 16887 4956 16923 4957
rect 16989 4990 17026 4991
rect 16989 4989 17027 4990
rect 16989 4981 17053 4989
rect 16989 4961 16998 4981
rect 17018 4967 17053 4981
rect 17073 4967 17076 4987
rect 17018 4962 17076 4967
rect 17018 4961 17053 4962
rect 16255 4924 16292 4953
rect 16256 4922 16292 4924
rect 16468 4922 16505 4953
rect 16256 4900 16505 4922
rect 16676 4921 16713 4953
rect 16989 4949 17053 4961
rect 17093 4923 17120 5101
rect 16952 4921 17120 4923
rect 16676 4895 17120 4921
rect 17272 5020 17522 5044
rect 17272 4949 17309 5020
rect 17424 4959 17455 4960
rect 17272 4929 17281 4949
rect 17301 4929 17309 4949
rect 17272 4919 17309 4929
rect 17368 4949 17455 4959
rect 17368 4929 17377 4949
rect 17397 4929 17455 4949
rect 17368 4920 17455 4929
rect 17368 4919 17405 4920
rect 16676 4885 16698 4895
rect 16952 4894 17120 4895
rect 16636 4883 16698 4885
rect 16066 4876 16698 4883
rect 15483 4832 15524 4833
rect 14807 4779 14844 4780
rect 14903 4779 14940 4780
rect 14959 4779 14995 4831
rect 15014 4779 15051 4780
rect 14707 4770 14845 4779
rect 14707 4750 14816 4770
rect 14836 4750 14845 4770
rect 14707 4743 14845 4750
rect 14903 4770 15051 4779
rect 14903 4750 14912 4770
rect 14932 4750 15022 4770
rect 15042 4750 15051 4770
rect 14707 4741 14803 4743
rect 14903 4740 15051 4750
rect 15110 4770 15147 4780
rect 15222 4779 15259 4780
rect 15203 4777 15259 4779
rect 15110 4750 15118 4770
rect 15138 4750 15147 4770
rect 14959 4739 14995 4740
rect 12872 4731 12903 4734
rect 13401 4734 13569 4735
rect 11701 4707 11839 4716
rect 13401 4708 13845 4734
rect 11495 4706 11532 4707
rect 11551 4655 11587 4707
rect 11606 4706 11643 4707
rect 11702 4706 11739 4707
rect 11022 4653 11063 4654
rect 10914 4646 11063 4653
rect 10914 4626 11032 4646
rect 11052 4626 11063 4646
rect 10914 4618 11063 4626
rect 11130 4650 11489 4654
rect 11130 4645 11452 4650
rect 11130 4621 11243 4645
rect 11267 4626 11452 4645
rect 11476 4626 11489 4650
rect 11267 4621 11489 4626
rect 11130 4618 11489 4621
rect 11551 4618 11586 4655
rect 11654 4652 11754 4655
rect 11654 4648 11721 4652
rect 11654 4622 11666 4648
rect 11692 4626 11721 4648
rect 11747 4626 11754 4652
rect 11692 4622 11754 4626
rect 11654 4618 11754 4622
rect 10341 4605 10379 4615
rect 9730 4601 9900 4602
rect 10341 4601 10351 4605
rect 8105 4584 8205 4588
rect 8105 4580 8167 4584
rect 8105 4554 8112 4580
rect 8138 4558 8167 4580
rect 8193 4558 8205 4584
rect 8138 4554 8205 4558
rect 8105 4551 8205 4554
rect 8273 4551 8308 4588
rect 8370 4585 8729 4588
rect 8370 4580 8592 4585
rect 8370 4556 8383 4580
rect 8407 4561 8592 4580
rect 8616 4561 8729 4585
rect 8407 4556 8729 4561
rect 8370 4552 8729 4556
rect 8796 4580 8945 4588
rect 9730 4587 10351 4601
rect 10369 4587 10379 4605
rect 11130 4597 11161 4618
rect 11551 4597 11587 4618
rect 9730 4581 10379 4587
rect 10794 4588 10831 4597
rect 10973 4596 11010 4597
rect 9730 4580 10378 4581
rect 8796 4560 8807 4580
rect 8827 4560 8945 4580
rect 10341 4578 10378 4580
rect 10794 4570 10803 4588
rect 10821 4570 10831 4588
rect 10794 4560 10831 4570
rect 8796 4553 8945 4560
rect 8796 4552 8837 4553
rect 8120 4499 8157 4500
rect 8216 4499 8253 4500
rect 8272 4499 8308 4551
rect 8327 4499 8364 4500
rect 6014 4472 6458 4498
rect 6015 4455 6039 4472
rect 6290 4471 6458 4472
rect 6909 4468 7159 4492
rect 5058 4451 5096 4452
rect 4469 4433 5096 4451
rect 5413 4437 6040 4455
rect 5413 4436 5451 4437
rect 3350 4396 3600 4420
rect 4051 4416 4219 4417
rect 4470 4416 4494 4433
rect 4051 4390 4495 4416
rect 2145 4388 2182 4389
rect 2201 4337 2237 4389
rect 2256 4388 2293 4389
rect 2352 4388 2389 4389
rect 1672 4335 1713 4336
rect 1564 4328 1713 4335
rect 131 4308 168 4310
rect 1564 4308 1682 4328
rect 1702 4308 1713 4328
rect 131 4307 779 4308
rect 130 4301 779 4307
rect 130 4283 140 4301
rect 158 4287 779 4301
rect 1564 4300 1713 4308
rect 1780 4332 2139 4336
rect 1780 4327 2102 4332
rect 1780 4303 1893 4327
rect 1917 4308 2102 4327
rect 2126 4308 2139 4332
rect 1917 4303 2139 4308
rect 1780 4300 2139 4303
rect 2201 4300 2236 4337
rect 2304 4334 2404 4337
rect 2304 4330 2371 4334
rect 2304 4304 2316 4330
rect 2342 4308 2371 4330
rect 2397 4308 2404 4334
rect 2342 4304 2404 4308
rect 2304 4300 2404 4304
rect 158 4283 168 4287
rect 609 4286 779 4287
rect 130 4273 168 4283
rect 130 4195 165 4273
rect 742 4263 779 4286
rect 1780 4279 1811 4300
rect 2201 4279 2237 4300
rect 1623 4278 1660 4279
rect 1622 4269 1660 4278
rect 126 4186 165 4195
rect 126 4168 136 4186
rect 154 4168 165 4186
rect 126 4162 165 4168
rect 321 4238 571 4262
rect 321 4167 358 4238
rect 473 4177 504 4178
rect 126 4158 163 4162
rect 321 4147 330 4167
rect 350 4147 358 4167
rect 321 4137 358 4147
rect 417 4167 504 4177
rect 417 4147 426 4167
rect 446 4147 504 4167
rect 417 4138 504 4147
rect 417 4137 454 4138
rect 129 4087 166 4096
rect 127 4069 138 4087
rect 156 4069 166 4087
rect 473 4085 504 4138
rect 534 4167 571 4238
rect 742 4243 1135 4263
rect 1155 4243 1158 4263
rect 742 4238 1158 4243
rect 1622 4249 1631 4269
rect 1651 4249 1660 4269
rect 1622 4241 1660 4249
rect 1726 4273 1811 4279
rect 1836 4278 1873 4279
rect 1726 4253 1734 4273
rect 1754 4253 1811 4273
rect 1726 4245 1811 4253
rect 1835 4269 1873 4278
rect 1835 4249 1844 4269
rect 1864 4249 1873 4269
rect 1726 4244 1762 4245
rect 1835 4241 1873 4249
rect 1939 4273 2024 4279
rect 2044 4278 2081 4279
rect 1939 4253 1947 4273
rect 1967 4272 2024 4273
rect 1967 4253 1996 4272
rect 1939 4252 1996 4253
rect 2017 4252 2024 4272
rect 1939 4245 2024 4252
rect 2043 4269 2081 4278
rect 2043 4249 2052 4269
rect 2072 4249 2081 4269
rect 1939 4244 1975 4245
rect 2043 4241 2081 4249
rect 2147 4274 2291 4279
rect 2147 4273 2211 4274
rect 2147 4253 2155 4273
rect 2175 4255 2211 4273
rect 2237 4273 2291 4274
rect 2237 4255 2263 4273
rect 2175 4253 2263 4255
rect 2283 4253 2291 4273
rect 2147 4245 2291 4253
rect 2147 4244 2183 4245
rect 2255 4244 2291 4245
rect 2357 4278 2394 4279
rect 2357 4277 2395 4278
rect 2357 4269 2421 4277
rect 2357 4249 2366 4269
rect 2386 4255 2421 4269
rect 2441 4255 2444 4275
rect 2386 4250 2444 4255
rect 2386 4249 2421 4250
rect 742 4237 1083 4238
rect 686 4177 717 4178
rect 534 4147 543 4167
rect 563 4147 571 4167
rect 534 4137 571 4147
rect 630 4170 717 4177
rect 630 4167 691 4170
rect 630 4147 639 4167
rect 659 4150 691 4167
rect 712 4150 717 4170
rect 659 4147 717 4150
rect 630 4140 717 4147
rect 742 4167 779 4237
rect 1045 4236 1082 4237
rect 1623 4212 1660 4241
rect 1624 4210 1660 4212
rect 1836 4210 1873 4241
rect 1624 4188 1873 4210
rect 2044 4209 2081 4241
rect 2357 4237 2421 4249
rect 2461 4214 2488 4389
rect 2441 4211 2488 4214
rect 2320 4209 2488 4211
rect 4051 4388 4219 4390
rect 4051 4210 4078 4388
rect 4118 4350 4182 4362
rect 4458 4358 4495 4390
rect 4666 4389 4915 4411
rect 4666 4358 4703 4389
rect 4879 4387 4915 4389
rect 5058 4392 5096 4433
rect 5411 4431 5451 4436
rect 4879 4358 4916 4387
rect 4118 4349 4153 4350
rect 4095 4344 4153 4349
rect 4095 4324 4098 4344
rect 4118 4330 4153 4344
rect 4173 4330 4182 4350
rect 4118 4322 4182 4330
rect 4144 4321 4182 4322
rect 4145 4320 4182 4321
rect 4248 4354 4284 4355
rect 4356 4354 4392 4355
rect 4248 4348 4392 4354
rect 4248 4346 4314 4348
rect 4248 4326 4256 4346
rect 4276 4327 4314 4346
rect 4336 4346 4392 4348
rect 4336 4327 4364 4346
rect 4276 4326 4364 4327
rect 4384 4326 4392 4346
rect 4248 4320 4392 4326
rect 4458 4350 4496 4358
rect 4564 4354 4600 4355
rect 4458 4330 4467 4350
rect 4487 4330 4496 4350
rect 4458 4321 4496 4330
rect 4515 4347 4600 4354
rect 4515 4327 4522 4347
rect 4543 4346 4600 4347
rect 4543 4327 4572 4346
rect 4515 4326 4572 4327
rect 4592 4326 4600 4346
rect 4458 4320 4495 4321
rect 4515 4320 4600 4326
rect 4666 4350 4704 4358
rect 4777 4354 4813 4355
rect 4666 4330 4675 4350
rect 4695 4330 4704 4350
rect 4666 4321 4704 4330
rect 4728 4346 4813 4354
rect 4728 4326 4785 4346
rect 4805 4326 4813 4346
rect 4666 4320 4703 4321
rect 4728 4320 4813 4326
rect 4879 4350 4917 4358
rect 4879 4330 4888 4350
rect 4908 4330 4917 4350
rect 4879 4321 4917 4330
rect 5058 4357 5094 4392
rect 5411 4388 5446 4431
rect 5409 4379 5446 4388
rect 5409 4361 5419 4379
rect 5437 4361 5446 4379
rect 6909 4397 6946 4468
rect 7061 4407 7092 4408
rect 6909 4377 6918 4397
rect 6938 4377 6946 4397
rect 6909 4367 6946 4377
rect 7005 4397 7092 4407
rect 7005 4377 7014 4397
rect 7034 4377 7092 4397
rect 7005 4368 7092 4377
rect 7005 4367 7042 4368
rect 5058 4347 5095 4357
rect 5409 4351 5446 4361
rect 5058 4329 5068 4347
rect 5086 4329 5095 4347
rect 4879 4320 4916 4321
rect 5058 4320 5095 4329
rect 4302 4299 4338 4320
rect 4728 4299 4759 4320
rect 7061 4315 7092 4368
rect 7122 4397 7159 4468
rect 7330 4473 7723 4493
rect 7743 4473 7746 4493
rect 7330 4468 7746 4473
rect 8020 4490 8158 4499
rect 8020 4470 8129 4490
rect 8149 4470 8158 4490
rect 7330 4467 7671 4468
rect 7274 4407 7305 4408
rect 7122 4377 7131 4397
rect 7151 4377 7159 4397
rect 7122 4367 7159 4377
rect 7218 4400 7305 4407
rect 7218 4397 7279 4400
rect 7218 4377 7227 4397
rect 7247 4380 7279 4397
rect 7300 4380 7305 4400
rect 7247 4377 7305 4380
rect 7218 4370 7305 4377
rect 7330 4397 7367 4467
rect 7633 4466 7670 4467
rect 8020 4463 8158 4470
rect 8216 4490 8364 4499
rect 8216 4470 8225 4490
rect 8245 4470 8335 4490
rect 8355 4470 8364 4490
rect 8020 4461 8116 4463
rect 8216 4460 8364 4470
rect 8423 4490 8460 4500
rect 8535 4499 8572 4500
rect 8516 4497 8572 4499
rect 8423 4470 8431 4490
rect 8451 4470 8460 4490
rect 8272 4459 8308 4460
rect 7482 4407 7518 4408
rect 7330 4377 7339 4397
rect 7359 4377 7367 4397
rect 7218 4368 7274 4370
rect 7218 4367 7255 4368
rect 7330 4367 7367 4377
rect 7426 4397 7574 4407
rect 7674 4404 7770 4406
rect 7426 4377 7435 4397
rect 7455 4377 7545 4397
rect 7565 4377 7574 4397
rect 7426 4368 7574 4377
rect 7632 4397 7770 4404
rect 8120 4400 8157 4401
rect 8423 4400 8460 4470
rect 8485 4490 8572 4497
rect 8485 4487 8543 4490
rect 8485 4467 8490 4487
rect 8511 4470 8543 4487
rect 8563 4470 8572 4490
rect 8511 4467 8572 4470
rect 8485 4460 8572 4467
rect 8631 4490 8668 4500
rect 8631 4470 8639 4490
rect 8659 4470 8668 4490
rect 8485 4459 8516 4460
rect 8119 4399 8460 4400
rect 7632 4377 7641 4397
rect 7661 4377 7770 4397
rect 7632 4368 7770 4377
rect 8044 4394 8460 4399
rect 8044 4374 8047 4394
rect 8067 4374 8460 4394
rect 8631 4399 8668 4470
rect 8698 4499 8729 4552
rect 10795 4525 10831 4560
rect 10972 4587 11010 4596
rect 10972 4567 10981 4587
rect 11001 4567 11010 4587
rect 10972 4559 11010 4567
rect 11076 4591 11161 4597
rect 11186 4596 11223 4597
rect 11076 4571 11084 4591
rect 11104 4571 11161 4591
rect 11076 4563 11161 4571
rect 11185 4587 11223 4596
rect 11185 4567 11194 4587
rect 11214 4567 11223 4587
rect 11076 4562 11112 4563
rect 11185 4559 11223 4567
rect 11289 4591 11374 4597
rect 11394 4596 11431 4597
rect 11289 4571 11297 4591
rect 11317 4590 11374 4591
rect 11317 4571 11346 4590
rect 11289 4570 11346 4571
rect 11367 4570 11374 4590
rect 11289 4563 11374 4570
rect 11393 4587 11431 4596
rect 11393 4567 11402 4587
rect 11422 4567 11431 4587
rect 11289 4562 11325 4563
rect 11393 4559 11431 4567
rect 11497 4591 11641 4597
rect 11497 4571 11505 4591
rect 11525 4590 11613 4591
rect 11525 4571 11553 4590
rect 11497 4569 11553 4571
rect 11575 4571 11613 4590
rect 11633 4571 11641 4591
rect 11575 4569 11641 4571
rect 11497 4563 11641 4569
rect 11497 4562 11533 4563
rect 11605 4562 11641 4563
rect 11707 4596 11744 4597
rect 11707 4595 11745 4596
rect 11707 4587 11771 4595
rect 11707 4567 11716 4587
rect 11736 4573 11771 4587
rect 11791 4573 11794 4593
rect 11736 4568 11794 4573
rect 11736 4567 11771 4568
rect 10973 4530 11010 4559
rect 10344 4506 10381 4516
rect 8748 4499 8785 4500
rect 8698 4490 8785 4499
rect 8698 4470 8756 4490
rect 8776 4470 8785 4490
rect 8698 4460 8785 4470
rect 8844 4490 8881 4500
rect 8844 4470 8852 4490
rect 8872 4470 8881 4490
rect 8698 4459 8729 4460
rect 8844 4399 8881 4470
rect 10344 4488 10353 4506
rect 10371 4488 10381 4506
rect 10344 4479 10381 4488
rect 10793 4484 10831 4525
rect 10974 4528 11010 4530
rect 11186 4528 11223 4559
rect 10974 4506 11223 4528
rect 11394 4527 11431 4559
rect 11707 4555 11771 4567
rect 11811 4529 11838 4707
rect 11670 4527 11838 4529
rect 13401 4706 13569 4708
rect 13401 4703 13448 4706
rect 13401 4528 13428 4703
rect 13468 4668 13532 4680
rect 13808 4676 13845 4708
rect 14016 4707 14265 4729
rect 14016 4676 14053 4707
rect 14229 4705 14265 4707
rect 14229 4676 14266 4705
rect 14807 4680 14844 4681
rect 15110 4680 15147 4750
rect 15172 4770 15259 4777
rect 15172 4767 15230 4770
rect 15172 4747 15177 4767
rect 15198 4750 15230 4767
rect 15250 4750 15259 4770
rect 15198 4747 15259 4750
rect 15172 4740 15259 4747
rect 15318 4770 15355 4780
rect 15318 4750 15326 4770
rect 15346 4750 15355 4770
rect 15172 4739 15203 4740
rect 14806 4679 15147 4680
rect 13468 4667 13503 4668
rect 13445 4662 13503 4667
rect 13445 4642 13448 4662
rect 13468 4648 13503 4662
rect 13523 4648 13532 4668
rect 13468 4640 13532 4648
rect 13494 4639 13532 4640
rect 13495 4638 13532 4639
rect 13598 4672 13634 4673
rect 13706 4672 13742 4673
rect 13598 4664 13742 4672
rect 13598 4644 13606 4664
rect 13626 4662 13714 4664
rect 13626 4644 13652 4662
rect 13598 4643 13652 4644
rect 13678 4644 13714 4662
rect 13734 4644 13742 4664
rect 13678 4643 13742 4644
rect 13598 4638 13742 4643
rect 13808 4668 13846 4676
rect 13914 4672 13950 4673
rect 13808 4648 13817 4668
rect 13837 4648 13846 4668
rect 13808 4639 13846 4648
rect 13865 4665 13950 4672
rect 13865 4645 13872 4665
rect 13893 4664 13950 4665
rect 13893 4645 13922 4664
rect 13865 4644 13922 4645
rect 13942 4644 13950 4664
rect 13808 4638 13845 4639
rect 13865 4638 13950 4644
rect 14016 4668 14054 4676
rect 14127 4672 14163 4673
rect 14016 4648 14025 4668
rect 14045 4648 14054 4668
rect 14016 4639 14054 4648
rect 14078 4664 14163 4672
rect 14078 4644 14135 4664
rect 14155 4644 14163 4664
rect 14016 4638 14053 4639
rect 14078 4638 14163 4644
rect 14229 4668 14267 4676
rect 14229 4648 14238 4668
rect 14258 4648 14267 4668
rect 14731 4674 15147 4679
rect 14731 4654 14734 4674
rect 14754 4654 15147 4674
rect 15318 4679 15355 4750
rect 15385 4779 15416 4832
rect 15723 4830 15733 4848
rect 15751 4830 15762 4848
rect 16065 4867 16698 4876
rect 17424 4867 17455 4920
rect 17485 4949 17522 5020
rect 17693 5025 18086 5045
rect 18106 5025 18109 5045
rect 17693 5020 18109 5025
rect 17693 5019 18034 5020
rect 17637 4959 17668 4960
rect 17485 4929 17494 4949
rect 17514 4929 17522 4949
rect 17485 4919 17522 4929
rect 17581 4952 17668 4959
rect 17581 4949 17642 4952
rect 17581 4929 17590 4949
rect 17610 4932 17642 4949
rect 17663 4932 17668 4952
rect 17610 4929 17668 4932
rect 17581 4922 17668 4929
rect 17693 4949 17730 5019
rect 17996 5018 18033 5019
rect 17845 4959 17881 4960
rect 17693 4929 17702 4949
rect 17722 4929 17730 4949
rect 17581 4920 17637 4922
rect 17581 4919 17618 4920
rect 17693 4919 17730 4929
rect 17789 4949 17937 4959
rect 18037 4956 18133 4958
rect 17789 4929 17798 4949
rect 17818 4929 17908 4949
rect 17928 4929 17937 4949
rect 17789 4920 17937 4929
rect 17995 4949 18133 4956
rect 17995 4929 18004 4949
rect 18024 4929 18133 4949
rect 17995 4920 18133 4929
rect 17789 4919 17826 4920
rect 17845 4868 17881 4920
rect 17900 4919 17937 4920
rect 17996 4919 18033 4920
rect 16065 4849 16075 4867
rect 16093 4866 16698 4867
rect 17316 4866 17357 4867
rect 16093 4861 16114 4866
rect 16093 4849 16105 4861
rect 17208 4859 17357 4866
rect 16065 4841 16105 4849
rect 16148 4848 16174 4849
rect 16065 4839 16102 4841
rect 16148 4830 16702 4848
rect 17208 4839 17326 4859
rect 17346 4839 17357 4859
rect 17208 4831 17357 4839
rect 17424 4863 17783 4867
rect 17424 4858 17746 4863
rect 17424 4834 17537 4858
rect 17561 4839 17746 4858
rect 17770 4839 17783 4863
rect 17561 4834 17783 4839
rect 17424 4831 17783 4834
rect 17845 4831 17880 4868
rect 17948 4865 18048 4868
rect 17948 4861 18015 4865
rect 17948 4835 17960 4861
rect 17986 4839 18015 4861
rect 18041 4839 18048 4865
rect 17986 4835 18048 4839
rect 17948 4831 18048 4835
rect 15723 4821 15760 4830
rect 15435 4779 15472 4780
rect 15385 4770 15472 4779
rect 15385 4750 15443 4770
rect 15463 4750 15472 4770
rect 15385 4740 15472 4750
rect 15531 4770 15568 4780
rect 15531 4750 15539 4770
rect 15559 4750 15568 4770
rect 16068 4771 16105 4777
rect 16148 4771 16174 4830
rect 16681 4811 16702 4830
rect 16068 4768 16174 4771
rect 15726 4755 15763 4759
rect 15385 4739 15416 4740
rect 15531 4679 15568 4750
rect 15318 4655 15568 4679
rect 15724 4749 15763 4755
rect 15724 4731 15735 4749
rect 15753 4731 15763 4749
rect 16068 4750 16077 4768
rect 16095 4754 16174 4768
rect 16259 4786 16509 4810
rect 16095 4752 16171 4754
rect 16095 4750 16105 4752
rect 16068 4740 16105 4750
rect 15724 4722 15763 4731
rect 14229 4639 14267 4648
rect 14229 4638 14266 4639
rect 13652 4617 13688 4638
rect 14078 4617 14109 4638
rect 15110 4631 15147 4654
rect 15724 4644 15759 4722
rect 16073 4675 16104 4740
rect 16259 4715 16296 4786
rect 16411 4725 16442 4726
rect 16259 4695 16268 4715
rect 16288 4695 16296 4715
rect 16259 4685 16296 4695
rect 16355 4715 16442 4725
rect 16355 4695 16364 4715
rect 16384 4695 16442 4715
rect 16355 4686 16442 4695
rect 16355 4685 16392 4686
rect 15721 4634 15759 4644
rect 16072 4666 16109 4675
rect 16072 4648 16082 4666
rect 16100 4648 16109 4666
rect 16072 4638 16109 4648
rect 15110 4630 15280 4631
rect 15721 4630 15731 4634
rect 13485 4613 13585 4617
rect 13485 4609 13547 4613
rect 13485 4583 13492 4609
rect 13518 4587 13547 4609
rect 13573 4587 13585 4613
rect 13518 4583 13585 4587
rect 13485 4580 13585 4583
rect 13653 4580 13688 4617
rect 13750 4614 14109 4617
rect 13750 4609 13972 4614
rect 13750 4585 13763 4609
rect 13787 4590 13972 4609
rect 13996 4590 14109 4614
rect 13787 4585 14109 4590
rect 13750 4581 14109 4585
rect 14176 4609 14325 4617
rect 15110 4616 15731 4630
rect 15749 4616 15759 4634
rect 16411 4633 16442 4686
rect 16472 4715 16509 4786
rect 16680 4791 17073 4811
rect 17093 4791 17096 4811
rect 17424 4810 17455 4831
rect 17845 4810 17881 4831
rect 17267 4809 17304 4810
rect 16680 4786 17096 4791
rect 17266 4800 17304 4809
rect 16680 4785 17021 4786
rect 16624 4725 16655 4726
rect 16472 4695 16481 4715
rect 16501 4695 16509 4715
rect 16472 4685 16509 4695
rect 16568 4718 16655 4725
rect 16568 4715 16629 4718
rect 16568 4695 16577 4715
rect 16597 4698 16629 4715
rect 16650 4698 16655 4718
rect 16597 4695 16655 4698
rect 16568 4688 16655 4695
rect 16680 4715 16717 4785
rect 16983 4784 17020 4785
rect 17266 4780 17275 4800
rect 17295 4780 17304 4800
rect 17266 4772 17304 4780
rect 17370 4804 17455 4810
rect 17480 4809 17517 4810
rect 17370 4784 17378 4804
rect 17398 4784 17455 4804
rect 17370 4776 17455 4784
rect 17479 4800 17517 4809
rect 17479 4780 17488 4800
rect 17508 4780 17517 4800
rect 17370 4775 17406 4776
rect 17479 4772 17517 4780
rect 17583 4804 17668 4810
rect 17688 4809 17725 4810
rect 17583 4784 17591 4804
rect 17611 4803 17668 4804
rect 17611 4784 17640 4803
rect 17583 4783 17640 4784
rect 17661 4783 17668 4803
rect 17583 4776 17668 4783
rect 17687 4800 17725 4809
rect 17687 4780 17696 4800
rect 17716 4780 17725 4800
rect 17583 4775 17619 4776
rect 17687 4772 17725 4780
rect 17791 4805 17935 4810
rect 17791 4804 17850 4805
rect 17791 4784 17799 4804
rect 17819 4785 17850 4804
rect 17874 4804 17935 4805
rect 17874 4785 17907 4804
rect 17819 4784 17907 4785
rect 17927 4784 17935 4804
rect 17791 4776 17935 4784
rect 17791 4775 17827 4776
rect 17899 4775 17935 4776
rect 18001 4809 18038 4810
rect 18001 4808 18039 4809
rect 18001 4800 18065 4808
rect 18001 4780 18010 4800
rect 18030 4786 18065 4800
rect 18085 4786 18088 4806
rect 18030 4781 18088 4786
rect 18030 4780 18065 4781
rect 17267 4743 17304 4772
rect 17268 4741 17304 4743
rect 17480 4741 17517 4772
rect 16832 4725 16868 4726
rect 16680 4695 16689 4715
rect 16709 4695 16717 4715
rect 16568 4686 16624 4688
rect 16568 4685 16605 4686
rect 16680 4685 16717 4695
rect 16776 4715 16924 4725
rect 17024 4722 17120 4724
rect 16776 4695 16785 4715
rect 16805 4695 16895 4715
rect 16915 4695 16924 4715
rect 16776 4686 16924 4695
rect 16982 4715 17120 4722
rect 17268 4719 17517 4741
rect 17688 4740 17725 4772
rect 18001 4768 18065 4780
rect 18105 4742 18132 4920
rect 17964 4740 18132 4742
rect 17688 4736 18132 4740
rect 16982 4695 16991 4715
rect 17011 4695 17120 4715
rect 17688 4717 17737 4736
rect 17757 4717 18132 4736
rect 17688 4714 18132 4717
rect 17964 4713 18132 4714
rect 18153 4739 18184 5133
rect 18245 5137 18250 5155
rect 18270 5137 18277 5155
rect 18245 5132 18277 5137
rect 18248 5130 18277 5132
rect 18153 4713 18158 4739
rect 18177 4713 18184 4739
rect 18691 4714 18729 6545
rect 18757 6432 18784 6610
rect 18824 6572 18888 6584
rect 19164 6580 19201 6612
rect 19372 6611 19621 6633
rect 20076 6619 20113 6620
rect 20379 6619 20416 6689
rect 20441 6709 20528 6716
rect 20441 6706 20499 6709
rect 20441 6686 20446 6706
rect 20467 6689 20499 6706
rect 20519 6689 20528 6709
rect 20467 6686 20528 6689
rect 20441 6679 20528 6686
rect 20587 6709 20624 6719
rect 20587 6689 20595 6709
rect 20615 6689 20624 6709
rect 20441 6678 20472 6679
rect 20075 6618 20416 6619
rect 19372 6580 19409 6611
rect 19585 6609 19621 6611
rect 20000 6613 20416 6618
rect 19585 6580 19622 6609
rect 20000 6593 20003 6613
rect 20023 6593 20416 6613
rect 20587 6618 20624 6689
rect 20654 6718 20685 6771
rect 20992 6769 21002 6787
rect 21020 6769 21031 6787
rect 20992 6760 21029 6769
rect 20704 6718 20741 6719
rect 20654 6709 20741 6718
rect 20654 6689 20712 6709
rect 20732 6689 20741 6709
rect 20654 6679 20741 6689
rect 20800 6709 20837 6719
rect 20800 6689 20808 6709
rect 20828 6689 20837 6709
rect 20995 6694 21032 6698
rect 20654 6678 20685 6679
rect 20800 6618 20837 6689
rect 20587 6594 20837 6618
rect 20993 6688 21032 6694
rect 20993 6670 21004 6688
rect 21022 6670 21032 6688
rect 20993 6661 21032 6670
rect 18824 6571 18859 6572
rect 18801 6566 18859 6571
rect 18801 6546 18804 6566
rect 18824 6552 18859 6566
rect 18879 6552 18888 6572
rect 18824 6544 18888 6552
rect 18850 6543 18888 6544
rect 18851 6542 18888 6543
rect 18954 6576 18990 6577
rect 19062 6576 19098 6577
rect 18954 6568 19098 6576
rect 18954 6548 18962 6568
rect 18982 6567 19070 6568
rect 18982 6548 19011 6567
rect 19034 6548 19070 6567
rect 19090 6548 19098 6568
rect 18954 6542 19098 6548
rect 19164 6572 19202 6580
rect 19270 6576 19306 6577
rect 19164 6552 19173 6572
rect 19193 6552 19202 6572
rect 19164 6543 19202 6552
rect 19221 6569 19306 6576
rect 19221 6549 19228 6569
rect 19249 6568 19306 6569
rect 19249 6549 19278 6568
rect 19221 6548 19278 6549
rect 19298 6548 19306 6568
rect 19164 6542 19201 6543
rect 19221 6542 19306 6548
rect 19372 6572 19410 6580
rect 19483 6576 19519 6577
rect 19372 6552 19381 6572
rect 19401 6552 19410 6572
rect 19372 6543 19410 6552
rect 19434 6568 19519 6576
rect 19434 6548 19491 6568
rect 19511 6548 19519 6568
rect 19372 6542 19409 6543
rect 19434 6542 19519 6548
rect 19585 6572 19623 6580
rect 19585 6552 19594 6572
rect 19614 6552 19623 6572
rect 19585 6543 19623 6552
rect 20379 6570 20416 6593
rect 20993 6583 21028 6661
rect 20990 6573 21028 6583
rect 20379 6569 20549 6570
rect 20990 6569 21000 6573
rect 20379 6555 21000 6569
rect 21018 6555 21028 6573
rect 20379 6549 21028 6555
rect 20379 6548 21027 6549
rect 20990 6546 21027 6548
rect 19585 6542 19622 6543
rect 19008 6521 19044 6542
rect 19434 6521 19465 6542
rect 18841 6517 18941 6521
rect 18841 6513 18903 6517
rect 18841 6487 18848 6513
rect 18874 6491 18903 6513
rect 18929 6491 18941 6517
rect 18874 6487 18941 6491
rect 18841 6484 18941 6487
rect 19009 6484 19044 6521
rect 19106 6518 19465 6521
rect 19106 6513 19328 6518
rect 19106 6489 19119 6513
rect 19143 6494 19328 6513
rect 19352 6494 19465 6518
rect 19143 6489 19465 6494
rect 19106 6485 19465 6489
rect 19532 6513 19681 6521
rect 19532 6493 19543 6513
rect 19563 6493 19681 6513
rect 19532 6486 19681 6493
rect 19532 6485 19573 6486
rect 18856 6432 18893 6433
rect 18952 6432 18989 6433
rect 19008 6432 19044 6484
rect 19063 6432 19100 6433
rect 18756 6423 18894 6432
rect 18756 6403 18865 6423
rect 18885 6403 18894 6423
rect 18756 6396 18894 6403
rect 18952 6423 19100 6432
rect 18952 6403 18961 6423
rect 18981 6403 19071 6423
rect 19091 6403 19100 6423
rect 18756 6394 18852 6396
rect 18952 6393 19100 6403
rect 19159 6423 19196 6433
rect 19271 6432 19308 6433
rect 19252 6430 19308 6432
rect 19159 6403 19167 6423
rect 19187 6403 19196 6423
rect 19008 6392 19044 6393
rect 18856 6333 18893 6334
rect 19159 6333 19196 6403
rect 19221 6423 19308 6430
rect 19221 6420 19279 6423
rect 19221 6400 19226 6420
rect 19247 6403 19279 6420
rect 19299 6403 19308 6423
rect 19247 6400 19308 6403
rect 19221 6393 19308 6400
rect 19367 6423 19404 6433
rect 19367 6403 19375 6423
rect 19395 6403 19404 6423
rect 19221 6392 19252 6393
rect 18855 6332 19196 6333
rect 18780 6327 19196 6332
rect 18780 6307 18783 6327
rect 18803 6307 19196 6327
rect 19367 6332 19404 6403
rect 19434 6432 19465 6485
rect 20993 6474 21030 6484
rect 20993 6456 21002 6474
rect 21020 6456 21030 6474
rect 20993 6447 21030 6456
rect 19484 6432 19521 6433
rect 19434 6423 19521 6432
rect 19434 6403 19492 6423
rect 19512 6403 19521 6423
rect 19434 6393 19521 6403
rect 19580 6423 19617 6433
rect 19580 6403 19588 6423
rect 19608 6403 19617 6423
rect 19434 6392 19465 6393
rect 19580 6332 19617 6403
rect 20993 6401 21028 6447
rect 20992 6395 21030 6401
rect 20403 6377 21030 6395
rect 19367 6308 19617 6332
rect 19985 6360 20153 6361
rect 20404 6360 20428 6377
rect 19985 6334 20429 6360
rect 19985 6332 20153 6334
rect 19985 6154 20012 6332
rect 20052 6294 20116 6306
rect 20392 6302 20429 6334
rect 20600 6333 20849 6355
rect 20600 6302 20637 6333
rect 20813 6331 20849 6333
rect 20992 6336 21030 6377
rect 20813 6302 20850 6331
rect 20052 6293 20087 6294
rect 20029 6288 20087 6293
rect 20029 6268 20032 6288
rect 20052 6274 20087 6288
rect 20107 6274 20116 6294
rect 20052 6266 20116 6274
rect 20078 6265 20116 6266
rect 20079 6264 20116 6265
rect 20182 6298 20218 6299
rect 20290 6298 20326 6299
rect 20182 6292 20326 6298
rect 20182 6290 20248 6292
rect 20182 6270 20190 6290
rect 20210 6271 20248 6290
rect 20270 6290 20326 6292
rect 20270 6271 20298 6290
rect 20210 6270 20298 6271
rect 20318 6270 20326 6290
rect 20182 6264 20326 6270
rect 20392 6294 20430 6302
rect 20498 6298 20534 6299
rect 20392 6274 20401 6294
rect 20421 6274 20430 6294
rect 20392 6265 20430 6274
rect 20449 6291 20534 6298
rect 20449 6271 20456 6291
rect 20477 6290 20534 6291
rect 20477 6271 20506 6290
rect 20449 6270 20506 6271
rect 20526 6270 20534 6290
rect 20392 6264 20429 6265
rect 20449 6264 20534 6270
rect 20600 6294 20638 6302
rect 20711 6298 20747 6299
rect 20600 6274 20609 6294
rect 20629 6274 20638 6294
rect 20600 6265 20638 6274
rect 20662 6290 20747 6298
rect 20662 6270 20719 6290
rect 20739 6270 20747 6290
rect 20600 6264 20637 6265
rect 20662 6264 20747 6270
rect 20813 6294 20851 6302
rect 20813 6274 20822 6294
rect 20842 6274 20851 6294
rect 20813 6265 20851 6274
rect 20992 6301 21028 6336
rect 20992 6291 21029 6301
rect 20992 6273 21002 6291
rect 21020 6273 21029 6291
rect 20813 6264 20850 6265
rect 20992 6264 21029 6273
rect 20236 6243 20272 6264
rect 20662 6243 20693 6264
rect 20069 6239 20169 6243
rect 20069 6235 20131 6239
rect 20069 6209 20076 6235
rect 20102 6213 20131 6235
rect 20157 6213 20169 6239
rect 20102 6209 20169 6213
rect 20069 6206 20169 6209
rect 20237 6206 20272 6243
rect 20334 6240 20693 6243
rect 20334 6235 20556 6240
rect 20334 6211 20347 6235
rect 20371 6216 20556 6235
rect 20580 6216 20693 6240
rect 20371 6211 20693 6216
rect 20334 6207 20693 6211
rect 20760 6235 20909 6243
rect 20760 6215 20771 6235
rect 20791 6215 20909 6235
rect 20760 6208 20909 6215
rect 20760 6207 20801 6208
rect 20084 6154 20121 6155
rect 20180 6154 20217 6155
rect 20236 6154 20272 6206
rect 20291 6154 20328 6155
rect 19984 6145 20122 6154
rect 18920 6127 18951 6130
rect 18920 6101 18927 6127
rect 18946 6101 18951 6127
rect 18920 5707 18951 6101
rect 18972 6126 19140 6127
rect 18972 6123 19416 6126
rect 18972 6104 19347 6123
rect 19367 6104 19416 6123
rect 19984 6125 20093 6145
rect 20113 6125 20122 6145
rect 18972 6100 19416 6104
rect 18972 6098 19140 6100
rect 18972 5920 18999 6098
rect 19039 6060 19103 6072
rect 19379 6068 19416 6100
rect 19587 6099 19836 6121
rect 19984 6118 20122 6125
rect 20180 6145 20328 6154
rect 20180 6125 20189 6145
rect 20209 6125 20299 6145
rect 20319 6125 20328 6145
rect 19984 6116 20080 6118
rect 20180 6115 20328 6125
rect 20387 6145 20424 6155
rect 20499 6154 20536 6155
rect 20480 6152 20536 6154
rect 20387 6125 20395 6145
rect 20415 6125 20424 6145
rect 20236 6114 20272 6115
rect 19587 6068 19624 6099
rect 19800 6097 19836 6099
rect 19800 6068 19837 6097
rect 19039 6059 19074 6060
rect 19016 6054 19074 6059
rect 19016 6034 19019 6054
rect 19039 6040 19074 6054
rect 19094 6040 19103 6060
rect 19039 6032 19103 6040
rect 19065 6031 19103 6032
rect 19066 6030 19103 6031
rect 19169 6064 19205 6065
rect 19277 6064 19313 6065
rect 19169 6056 19313 6064
rect 19169 6036 19177 6056
rect 19197 6055 19285 6056
rect 19197 6036 19230 6055
rect 19169 6035 19230 6036
rect 19254 6036 19285 6055
rect 19305 6036 19313 6056
rect 19254 6035 19313 6036
rect 19169 6030 19313 6035
rect 19379 6060 19417 6068
rect 19485 6064 19521 6065
rect 19379 6040 19388 6060
rect 19408 6040 19417 6060
rect 19379 6031 19417 6040
rect 19436 6057 19521 6064
rect 19436 6037 19443 6057
rect 19464 6056 19521 6057
rect 19464 6037 19493 6056
rect 19436 6036 19493 6037
rect 19513 6036 19521 6056
rect 19379 6030 19416 6031
rect 19436 6030 19521 6036
rect 19587 6060 19625 6068
rect 19698 6064 19734 6065
rect 19587 6040 19596 6060
rect 19616 6040 19625 6060
rect 19587 6031 19625 6040
rect 19649 6056 19734 6064
rect 19649 6036 19706 6056
rect 19726 6036 19734 6056
rect 19587 6030 19624 6031
rect 19649 6030 19734 6036
rect 19800 6060 19838 6068
rect 19800 6040 19809 6060
rect 19829 6040 19838 6060
rect 20084 6055 20121 6056
rect 20387 6055 20424 6125
rect 20449 6145 20536 6152
rect 20449 6142 20507 6145
rect 20449 6122 20454 6142
rect 20475 6125 20507 6142
rect 20527 6125 20536 6145
rect 20475 6122 20536 6125
rect 20449 6115 20536 6122
rect 20595 6145 20632 6155
rect 20595 6125 20603 6145
rect 20623 6125 20632 6145
rect 20449 6114 20480 6115
rect 20083 6054 20424 6055
rect 19800 6031 19838 6040
rect 20008 6049 20424 6054
rect 19800 6030 19837 6031
rect 19223 6009 19259 6030
rect 19649 6009 19680 6030
rect 20008 6029 20011 6049
rect 20031 6029 20424 6049
rect 20595 6054 20632 6125
rect 20662 6154 20693 6207
rect 20995 6192 21032 6202
rect 20995 6174 21004 6192
rect 21022 6174 21032 6192
rect 20995 6165 21032 6174
rect 20712 6154 20749 6155
rect 20662 6145 20749 6154
rect 20662 6125 20720 6145
rect 20740 6125 20749 6145
rect 20662 6115 20749 6125
rect 20808 6145 20845 6155
rect 20808 6125 20816 6145
rect 20836 6125 20845 6145
rect 20662 6114 20693 6115
rect 20808 6054 20845 6125
rect 21000 6100 21031 6165
rect 20999 6090 21036 6100
rect 20999 6088 21009 6090
rect 20933 6086 21009 6088
rect 20595 6030 20845 6054
rect 20930 6072 21009 6086
rect 21027 6072 21036 6090
rect 20930 6069 21036 6072
rect 20402 6010 20423 6029
rect 20930 6010 20956 6069
rect 20999 6063 21036 6069
rect 19056 6005 19156 6009
rect 19056 6001 19118 6005
rect 19056 5975 19063 6001
rect 19089 5979 19118 6001
rect 19144 5979 19156 6005
rect 19089 5975 19156 5979
rect 19056 5972 19156 5975
rect 19224 5972 19259 6009
rect 19321 6006 19680 6009
rect 19321 6001 19543 6006
rect 19321 5977 19334 6001
rect 19358 5982 19543 6001
rect 19567 5982 19680 6006
rect 19358 5977 19680 5982
rect 19321 5973 19680 5977
rect 19747 6001 19896 6009
rect 19747 5981 19758 6001
rect 19778 5981 19896 6001
rect 20402 5992 20956 6010
rect 21002 5999 21039 6001
rect 20930 5991 20956 5992
rect 20999 5991 21039 5999
rect 19747 5974 19896 5981
rect 20999 5979 21011 5991
rect 20990 5974 21011 5979
rect 19747 5973 19788 5974
rect 20406 5973 21011 5974
rect 21029 5973 21039 5991
rect 19071 5920 19108 5921
rect 19167 5920 19204 5921
rect 19223 5920 19259 5972
rect 19278 5920 19315 5921
rect 18971 5911 19109 5920
rect 18971 5891 19080 5911
rect 19100 5891 19109 5911
rect 18971 5884 19109 5891
rect 19167 5911 19315 5920
rect 19167 5891 19176 5911
rect 19196 5891 19286 5911
rect 19306 5891 19315 5911
rect 18971 5882 19067 5884
rect 19167 5881 19315 5891
rect 19374 5911 19411 5921
rect 19486 5920 19523 5921
rect 19467 5918 19523 5920
rect 19374 5891 19382 5911
rect 19402 5891 19411 5911
rect 19223 5880 19259 5881
rect 19071 5821 19108 5822
rect 19374 5821 19411 5891
rect 19436 5911 19523 5918
rect 19436 5908 19494 5911
rect 19436 5888 19441 5908
rect 19462 5891 19494 5908
rect 19514 5891 19523 5911
rect 19462 5888 19523 5891
rect 19436 5881 19523 5888
rect 19582 5911 19619 5921
rect 19582 5891 19590 5911
rect 19610 5891 19619 5911
rect 19436 5880 19467 5881
rect 19070 5820 19411 5821
rect 18995 5815 19411 5820
rect 18995 5795 18998 5815
rect 19018 5795 19411 5815
rect 19582 5820 19619 5891
rect 19649 5920 19680 5973
rect 20406 5964 21039 5973
rect 20406 5957 21038 5964
rect 20406 5955 20468 5957
rect 19984 5945 20152 5946
rect 20406 5945 20428 5955
rect 19699 5920 19736 5921
rect 19649 5911 19736 5920
rect 19649 5891 19707 5911
rect 19727 5891 19736 5911
rect 19649 5881 19736 5891
rect 19795 5911 19832 5921
rect 19795 5891 19803 5911
rect 19823 5891 19832 5911
rect 19649 5880 19680 5881
rect 19795 5820 19832 5891
rect 19582 5796 19832 5820
rect 19984 5919 20428 5945
rect 19984 5917 20152 5919
rect 19984 5739 20011 5917
rect 20051 5879 20115 5891
rect 20391 5887 20428 5919
rect 20599 5918 20848 5940
rect 20599 5887 20636 5918
rect 20812 5916 20848 5918
rect 20812 5887 20849 5916
rect 20051 5878 20086 5879
rect 20028 5873 20086 5878
rect 20028 5853 20031 5873
rect 20051 5859 20086 5873
rect 20106 5859 20115 5879
rect 20051 5851 20115 5859
rect 20077 5850 20115 5851
rect 20078 5849 20115 5850
rect 20181 5883 20217 5884
rect 20289 5883 20325 5884
rect 20181 5875 20325 5883
rect 20181 5855 20189 5875
rect 20209 5855 20238 5875
rect 20181 5854 20238 5855
rect 20260 5855 20297 5875
rect 20317 5855 20325 5875
rect 20260 5854 20325 5855
rect 20181 5849 20325 5854
rect 20391 5879 20429 5887
rect 20497 5883 20533 5884
rect 20391 5859 20400 5879
rect 20420 5859 20429 5879
rect 20391 5850 20429 5859
rect 20448 5876 20533 5883
rect 20448 5856 20455 5876
rect 20476 5875 20533 5876
rect 20476 5856 20505 5875
rect 20448 5855 20505 5856
rect 20525 5855 20533 5875
rect 20391 5849 20428 5850
rect 20448 5849 20533 5855
rect 20599 5879 20637 5887
rect 20710 5883 20746 5884
rect 20599 5859 20608 5879
rect 20628 5859 20637 5879
rect 20599 5850 20637 5859
rect 20661 5875 20746 5883
rect 20661 5855 20718 5875
rect 20738 5855 20746 5875
rect 20599 5849 20636 5850
rect 20661 5849 20746 5855
rect 20812 5879 20850 5887
rect 20812 5859 20821 5879
rect 20841 5859 20850 5879
rect 20812 5850 20850 5859
rect 20812 5849 20849 5850
rect 20235 5828 20271 5849
rect 20661 5828 20692 5849
rect 20068 5824 20168 5828
rect 20068 5820 20130 5824
rect 20068 5794 20075 5820
rect 20101 5798 20130 5820
rect 20156 5798 20168 5824
rect 20101 5794 20168 5798
rect 20068 5791 20168 5794
rect 20236 5791 20271 5828
rect 20333 5825 20692 5828
rect 20333 5820 20555 5825
rect 20333 5796 20346 5820
rect 20370 5801 20555 5820
rect 20579 5801 20692 5825
rect 20370 5796 20692 5801
rect 20333 5792 20692 5796
rect 20759 5820 20908 5828
rect 20759 5800 20770 5820
rect 20790 5800 20908 5820
rect 20759 5793 20908 5800
rect 20999 5808 21038 5957
rect 20759 5792 20800 5793
rect 20083 5739 20120 5740
rect 20179 5739 20216 5740
rect 20235 5739 20271 5791
rect 20290 5739 20327 5740
rect 19983 5730 20121 5739
rect 19983 5710 20092 5730
rect 20112 5710 20121 5730
rect 18920 5706 19090 5707
rect 18920 5691 19366 5706
rect 19983 5703 20121 5710
rect 20179 5730 20327 5739
rect 20179 5710 20188 5730
rect 20208 5710 20298 5730
rect 20318 5710 20327 5730
rect 19983 5701 20079 5703
rect 18922 5680 19366 5691
rect 18922 5678 19090 5680
rect 18922 5500 18949 5678
rect 18989 5640 19053 5652
rect 19329 5648 19366 5680
rect 19537 5679 19786 5701
rect 20179 5700 20327 5710
rect 20386 5730 20423 5740
rect 20498 5739 20535 5740
rect 20479 5737 20535 5739
rect 20386 5710 20394 5730
rect 20414 5710 20423 5730
rect 20235 5699 20271 5700
rect 19537 5648 19574 5679
rect 19750 5677 19786 5679
rect 19750 5648 19787 5677
rect 18989 5639 19024 5640
rect 18966 5634 19024 5639
rect 18966 5614 18969 5634
rect 18989 5620 19024 5634
rect 19044 5620 19053 5640
rect 18989 5612 19053 5620
rect 19015 5611 19053 5612
rect 19016 5610 19053 5611
rect 19119 5644 19155 5645
rect 19227 5644 19263 5645
rect 19119 5636 19263 5644
rect 19119 5616 19127 5636
rect 19147 5635 19235 5636
rect 19147 5618 19175 5635
rect 19199 5618 19235 5635
rect 19147 5616 19235 5618
rect 19255 5616 19263 5636
rect 19119 5610 19263 5616
rect 19329 5640 19367 5648
rect 19435 5644 19471 5645
rect 19329 5620 19338 5640
rect 19358 5620 19367 5640
rect 19329 5611 19367 5620
rect 19386 5637 19471 5644
rect 19386 5617 19393 5637
rect 19414 5636 19471 5637
rect 19414 5617 19443 5636
rect 19386 5616 19443 5617
rect 19463 5616 19471 5636
rect 19329 5610 19366 5611
rect 19386 5610 19471 5616
rect 19537 5640 19575 5648
rect 19648 5644 19684 5645
rect 19537 5620 19546 5640
rect 19566 5620 19575 5640
rect 19537 5611 19575 5620
rect 19599 5636 19684 5644
rect 19599 5616 19656 5636
rect 19676 5616 19684 5636
rect 19537 5610 19574 5611
rect 19599 5610 19684 5616
rect 19750 5640 19788 5648
rect 20083 5640 20120 5641
rect 20386 5640 20423 5710
rect 20448 5730 20535 5737
rect 20448 5727 20506 5730
rect 20448 5707 20453 5727
rect 20474 5710 20506 5727
rect 20526 5710 20535 5730
rect 20474 5707 20535 5710
rect 20448 5700 20535 5707
rect 20594 5730 20631 5740
rect 20594 5710 20602 5730
rect 20622 5710 20631 5730
rect 20448 5699 20479 5700
rect 19750 5620 19759 5640
rect 19779 5620 19788 5640
rect 20082 5639 20423 5640
rect 19750 5611 19788 5620
rect 20007 5634 20423 5639
rect 20007 5614 20010 5634
rect 20030 5614 20423 5634
rect 20594 5639 20631 5710
rect 20661 5739 20692 5792
rect 20999 5790 21009 5808
rect 21027 5790 21038 5808
rect 20999 5781 21036 5790
rect 20711 5739 20748 5740
rect 20661 5730 20748 5739
rect 20661 5710 20719 5730
rect 20739 5710 20748 5730
rect 20661 5700 20748 5710
rect 20807 5730 20844 5740
rect 20807 5710 20815 5730
rect 20835 5710 20844 5730
rect 21002 5715 21039 5719
rect 20661 5699 20692 5700
rect 20807 5639 20844 5710
rect 20594 5615 20844 5639
rect 21000 5709 21039 5715
rect 21000 5691 21011 5709
rect 21029 5691 21039 5709
rect 21000 5682 21039 5691
rect 19750 5610 19787 5611
rect 19173 5589 19209 5610
rect 19599 5589 19630 5610
rect 20386 5591 20423 5614
rect 21000 5604 21035 5682
rect 20997 5594 21035 5604
rect 20386 5590 20556 5591
rect 20997 5590 21007 5594
rect 19006 5585 19106 5589
rect 19006 5581 19068 5585
rect 19006 5555 19013 5581
rect 19039 5559 19068 5581
rect 19094 5559 19106 5585
rect 19039 5555 19106 5559
rect 19006 5552 19106 5555
rect 19174 5552 19209 5589
rect 19271 5586 19630 5589
rect 19271 5581 19493 5586
rect 19271 5557 19284 5581
rect 19308 5562 19493 5581
rect 19517 5562 19630 5586
rect 19308 5557 19630 5562
rect 19271 5553 19630 5557
rect 19697 5581 19846 5589
rect 19697 5561 19708 5581
rect 19728 5561 19846 5581
rect 20386 5576 21007 5590
rect 21025 5576 21035 5594
rect 20386 5570 21035 5576
rect 20386 5569 21034 5570
rect 20997 5567 21034 5569
rect 19697 5554 19846 5561
rect 19697 5553 19738 5554
rect 19021 5500 19058 5501
rect 19117 5500 19154 5501
rect 19173 5500 19209 5552
rect 19228 5500 19265 5501
rect 18921 5491 19059 5500
rect 18921 5471 19030 5491
rect 19050 5471 19059 5491
rect 18921 5464 19059 5471
rect 19117 5491 19265 5500
rect 19117 5471 19126 5491
rect 19146 5471 19236 5491
rect 19256 5471 19265 5491
rect 18921 5462 19017 5464
rect 19117 5461 19265 5471
rect 19324 5491 19361 5501
rect 19436 5500 19473 5501
rect 19417 5498 19473 5500
rect 19324 5471 19332 5491
rect 19352 5471 19361 5491
rect 19173 5460 19209 5461
rect 19021 5401 19058 5402
rect 19324 5401 19361 5471
rect 19386 5491 19473 5498
rect 19386 5488 19444 5491
rect 19386 5468 19391 5488
rect 19412 5471 19444 5488
rect 19464 5471 19473 5491
rect 19412 5468 19473 5471
rect 19386 5461 19473 5468
rect 19532 5491 19569 5501
rect 19532 5471 19540 5491
rect 19560 5471 19569 5491
rect 19386 5460 19417 5461
rect 19020 5400 19361 5401
rect 18945 5395 19361 5400
rect 18945 5375 18948 5395
rect 18968 5375 19361 5395
rect 19532 5400 19569 5471
rect 19599 5500 19630 5553
rect 19649 5500 19686 5501
rect 19599 5491 19686 5500
rect 19599 5471 19657 5491
rect 19677 5471 19686 5491
rect 19599 5461 19686 5471
rect 19745 5491 19782 5501
rect 19745 5471 19753 5491
rect 19773 5471 19782 5491
rect 19599 5460 19630 5461
rect 19745 5400 19782 5471
rect 21000 5495 21037 5505
rect 21000 5477 21009 5495
rect 21027 5477 21037 5495
rect 21000 5468 21037 5477
rect 21000 5444 21035 5468
rect 20998 5420 21035 5444
rect 20997 5414 21035 5420
rect 19532 5376 19782 5400
rect 20408 5396 21035 5414
rect 19990 5379 20158 5380
rect 20409 5379 20433 5396
rect 19990 5353 20434 5379
rect 19990 5351 20158 5353
rect 19990 5173 20017 5351
rect 20057 5313 20121 5325
rect 20397 5321 20434 5353
rect 20605 5352 20854 5374
rect 20605 5321 20642 5352
rect 20818 5350 20854 5352
rect 20997 5355 21035 5396
rect 20818 5321 20855 5350
rect 20057 5312 20092 5313
rect 20034 5307 20092 5312
rect 20034 5287 20037 5307
rect 20057 5293 20092 5307
rect 20112 5293 20121 5313
rect 20057 5285 20121 5293
rect 20083 5284 20121 5285
rect 20084 5283 20121 5284
rect 20187 5317 20223 5318
rect 20295 5317 20331 5318
rect 20187 5311 20331 5317
rect 20187 5309 20253 5311
rect 20187 5289 20195 5309
rect 20215 5290 20253 5309
rect 20275 5309 20331 5311
rect 20275 5290 20303 5309
rect 20215 5289 20303 5290
rect 20323 5289 20331 5309
rect 20187 5283 20331 5289
rect 20397 5313 20435 5321
rect 20503 5317 20539 5318
rect 20397 5293 20406 5313
rect 20426 5293 20435 5313
rect 20397 5284 20435 5293
rect 20454 5310 20539 5317
rect 20454 5290 20461 5310
rect 20482 5309 20539 5310
rect 20482 5290 20511 5309
rect 20454 5289 20511 5290
rect 20531 5289 20539 5309
rect 20397 5283 20434 5284
rect 20454 5283 20539 5289
rect 20605 5313 20643 5321
rect 20716 5317 20752 5318
rect 20605 5293 20614 5313
rect 20634 5293 20643 5313
rect 20605 5284 20643 5293
rect 20667 5309 20752 5317
rect 20667 5289 20724 5309
rect 20744 5289 20752 5309
rect 20605 5283 20642 5284
rect 20667 5283 20752 5289
rect 20818 5313 20856 5321
rect 20818 5293 20827 5313
rect 20847 5293 20856 5313
rect 20818 5284 20856 5293
rect 20997 5320 21033 5355
rect 20997 5310 21034 5320
rect 20997 5292 21007 5310
rect 21025 5292 21034 5310
rect 20818 5283 20855 5284
rect 20997 5283 21034 5292
rect 20241 5262 20277 5283
rect 20667 5262 20698 5283
rect 20074 5258 20174 5262
rect 20074 5254 20136 5258
rect 20074 5228 20081 5254
rect 20107 5232 20136 5254
rect 20162 5232 20174 5258
rect 20107 5228 20174 5232
rect 20074 5225 20174 5228
rect 20242 5225 20277 5262
rect 20339 5259 20698 5262
rect 20339 5254 20561 5259
rect 20339 5230 20352 5254
rect 20376 5235 20561 5254
rect 20585 5235 20698 5259
rect 20376 5230 20698 5235
rect 20339 5226 20698 5230
rect 20765 5254 20914 5262
rect 20765 5234 20776 5254
rect 20796 5234 20914 5254
rect 20765 5227 20914 5234
rect 20765 5226 20806 5227
rect 20089 5173 20126 5174
rect 20185 5173 20222 5174
rect 20241 5173 20277 5225
rect 20296 5173 20333 5174
rect 19989 5164 20127 5173
rect 18977 5145 19145 5146
rect 18977 5142 19421 5145
rect 18977 5123 19352 5142
rect 19372 5123 19421 5142
rect 19989 5144 20098 5164
rect 20118 5144 20127 5164
rect 18977 5119 19421 5123
rect 18977 5117 19145 5119
rect 18977 4939 19004 5117
rect 19044 5079 19108 5091
rect 19384 5087 19421 5119
rect 19592 5118 19841 5140
rect 19989 5137 20127 5144
rect 20185 5164 20333 5173
rect 20185 5144 20194 5164
rect 20214 5144 20304 5164
rect 20324 5144 20333 5164
rect 19989 5135 20085 5137
rect 20185 5134 20333 5144
rect 20392 5164 20429 5174
rect 20504 5173 20541 5174
rect 20485 5171 20541 5173
rect 20392 5144 20400 5164
rect 20420 5144 20429 5164
rect 20241 5133 20277 5134
rect 19592 5087 19629 5118
rect 19805 5116 19841 5118
rect 19805 5087 19842 5116
rect 19044 5078 19079 5079
rect 19021 5073 19079 5078
rect 19021 5053 19024 5073
rect 19044 5059 19079 5073
rect 19099 5059 19108 5079
rect 19044 5051 19108 5059
rect 19070 5050 19108 5051
rect 19071 5049 19108 5050
rect 19174 5083 19210 5084
rect 19282 5083 19318 5084
rect 19174 5075 19318 5083
rect 19174 5055 19182 5075
rect 19202 5055 19234 5075
rect 19258 5055 19290 5075
rect 19310 5055 19318 5075
rect 19174 5049 19318 5055
rect 19384 5079 19422 5087
rect 19490 5083 19526 5084
rect 19384 5059 19393 5079
rect 19413 5059 19422 5079
rect 19384 5050 19422 5059
rect 19441 5076 19526 5083
rect 19441 5056 19448 5076
rect 19469 5075 19526 5076
rect 19469 5056 19498 5075
rect 19441 5055 19498 5056
rect 19518 5055 19526 5075
rect 19384 5049 19421 5050
rect 19441 5049 19526 5055
rect 19592 5079 19630 5087
rect 19703 5083 19739 5084
rect 19592 5059 19601 5079
rect 19621 5059 19630 5079
rect 19592 5050 19630 5059
rect 19654 5075 19739 5083
rect 19654 5055 19711 5075
rect 19731 5055 19739 5075
rect 19592 5049 19629 5050
rect 19654 5049 19739 5055
rect 19805 5079 19843 5087
rect 19805 5059 19814 5079
rect 19834 5059 19843 5079
rect 20089 5074 20126 5075
rect 20392 5074 20429 5144
rect 20454 5164 20541 5171
rect 20454 5161 20512 5164
rect 20454 5141 20459 5161
rect 20480 5144 20512 5161
rect 20532 5144 20541 5164
rect 20480 5141 20541 5144
rect 20454 5134 20541 5141
rect 20600 5164 20637 5174
rect 20600 5144 20608 5164
rect 20628 5144 20637 5164
rect 20454 5133 20485 5134
rect 20088 5073 20429 5074
rect 19805 5050 19843 5059
rect 20013 5068 20429 5073
rect 19805 5049 19842 5050
rect 19228 5028 19264 5049
rect 19654 5028 19685 5049
rect 20013 5048 20016 5068
rect 20036 5048 20429 5068
rect 20600 5073 20637 5144
rect 20667 5173 20698 5226
rect 21000 5211 21037 5221
rect 21000 5193 21009 5211
rect 21027 5193 21037 5211
rect 21000 5184 21037 5193
rect 20717 5173 20754 5174
rect 20667 5164 20754 5173
rect 20667 5144 20725 5164
rect 20745 5144 20754 5164
rect 20667 5134 20754 5144
rect 20813 5164 20850 5174
rect 20813 5144 20821 5164
rect 20841 5144 20850 5164
rect 20667 5133 20698 5134
rect 20813 5073 20850 5144
rect 21005 5119 21036 5184
rect 21004 5109 21041 5119
rect 21004 5107 21014 5109
rect 20938 5105 21014 5107
rect 20600 5049 20850 5073
rect 20935 5091 21014 5105
rect 21032 5091 21041 5109
rect 20935 5088 21041 5091
rect 20407 5029 20428 5048
rect 20935 5029 20961 5088
rect 21004 5082 21041 5088
rect 19061 5024 19161 5028
rect 19061 5020 19123 5024
rect 19061 4994 19068 5020
rect 19094 4998 19123 5020
rect 19149 4998 19161 5024
rect 19094 4994 19161 4998
rect 19061 4991 19161 4994
rect 19229 4991 19264 5028
rect 19326 5025 19685 5028
rect 19326 5020 19548 5025
rect 19326 4996 19339 5020
rect 19363 5001 19548 5020
rect 19572 5001 19685 5025
rect 19363 4996 19685 5001
rect 19326 4992 19685 4996
rect 19752 5020 19901 5028
rect 19752 5000 19763 5020
rect 19783 5000 19901 5020
rect 20407 5011 20961 5029
rect 21007 5018 21044 5020
rect 20935 5010 20961 5011
rect 21004 5010 21044 5018
rect 19752 4993 19901 5000
rect 21004 4998 21016 5010
rect 20995 4993 21016 4998
rect 19752 4992 19793 4993
rect 20411 4992 21016 4993
rect 21034 4992 21044 5010
rect 19076 4939 19113 4940
rect 19172 4939 19209 4940
rect 19228 4939 19264 4991
rect 19283 4939 19320 4940
rect 18976 4930 19114 4939
rect 18976 4910 19085 4930
rect 19105 4910 19114 4930
rect 18976 4903 19114 4910
rect 19172 4930 19320 4939
rect 19172 4910 19181 4930
rect 19201 4910 19291 4930
rect 19311 4910 19320 4930
rect 18976 4901 19072 4903
rect 19172 4900 19320 4910
rect 19379 4930 19416 4940
rect 19491 4939 19528 4940
rect 19472 4937 19528 4939
rect 19379 4910 19387 4930
rect 19407 4910 19416 4930
rect 19228 4899 19264 4900
rect 19076 4840 19113 4841
rect 19379 4840 19416 4910
rect 19441 4930 19528 4937
rect 19441 4927 19499 4930
rect 19441 4907 19446 4927
rect 19467 4910 19499 4927
rect 19519 4910 19528 4930
rect 19467 4907 19528 4910
rect 19441 4900 19528 4907
rect 19587 4930 19624 4940
rect 19587 4910 19595 4930
rect 19615 4910 19624 4930
rect 19441 4899 19472 4900
rect 19075 4839 19416 4840
rect 19000 4834 19416 4839
rect 19000 4814 19003 4834
rect 19023 4814 19416 4834
rect 19587 4839 19624 4910
rect 19654 4939 19685 4992
rect 20411 4983 21044 4992
rect 20411 4976 21043 4983
rect 20411 4974 20473 4976
rect 19989 4964 20157 4965
rect 20411 4964 20433 4974
rect 19704 4939 19741 4940
rect 19654 4930 19741 4939
rect 19654 4910 19712 4930
rect 19732 4910 19741 4930
rect 19654 4900 19741 4910
rect 19800 4930 19837 4940
rect 19800 4910 19808 4930
rect 19828 4910 19837 4930
rect 19654 4899 19685 4900
rect 19800 4839 19837 4910
rect 19587 4815 19837 4839
rect 19989 4938 20433 4964
rect 19989 4936 20157 4938
rect 19989 4758 20016 4936
rect 20056 4898 20120 4910
rect 20396 4906 20433 4938
rect 20604 4937 20853 4959
rect 20604 4906 20641 4937
rect 20817 4935 20853 4937
rect 20817 4906 20854 4935
rect 20056 4897 20091 4898
rect 20033 4892 20091 4897
rect 20033 4872 20036 4892
rect 20056 4878 20091 4892
rect 20111 4878 20120 4898
rect 20056 4870 20120 4878
rect 20082 4869 20120 4870
rect 20083 4868 20120 4869
rect 20186 4902 20222 4903
rect 20294 4902 20330 4903
rect 20186 4894 20330 4902
rect 20186 4874 20194 4894
rect 20214 4874 20243 4894
rect 20186 4873 20243 4874
rect 20265 4874 20302 4894
rect 20322 4874 20330 4894
rect 20265 4873 20330 4874
rect 20186 4868 20330 4873
rect 20396 4898 20434 4906
rect 20502 4902 20538 4903
rect 20396 4878 20405 4898
rect 20425 4878 20434 4898
rect 20396 4869 20434 4878
rect 20453 4895 20538 4902
rect 20453 4875 20460 4895
rect 20481 4894 20538 4895
rect 20481 4875 20510 4894
rect 20453 4874 20510 4875
rect 20530 4874 20538 4894
rect 20396 4868 20433 4869
rect 20453 4868 20538 4874
rect 20604 4898 20642 4906
rect 20715 4902 20751 4903
rect 20604 4878 20613 4898
rect 20633 4878 20642 4898
rect 20604 4869 20642 4878
rect 20666 4894 20751 4902
rect 20666 4874 20723 4894
rect 20743 4874 20751 4894
rect 20604 4868 20641 4869
rect 20666 4868 20751 4874
rect 20817 4898 20855 4906
rect 20817 4878 20826 4898
rect 20846 4878 20855 4898
rect 20817 4869 20855 4878
rect 20817 4868 20854 4869
rect 20240 4847 20276 4868
rect 20666 4847 20697 4868
rect 20073 4843 20173 4847
rect 20073 4839 20135 4843
rect 20073 4813 20080 4839
rect 20106 4817 20135 4839
rect 20161 4817 20173 4843
rect 20106 4813 20173 4817
rect 20073 4810 20173 4813
rect 20241 4810 20276 4847
rect 20338 4844 20697 4847
rect 20338 4839 20560 4844
rect 20338 4815 20351 4839
rect 20375 4820 20560 4839
rect 20584 4820 20697 4844
rect 20375 4815 20697 4820
rect 20338 4811 20697 4815
rect 20764 4839 20913 4847
rect 20764 4819 20775 4839
rect 20795 4819 20913 4839
rect 20764 4812 20913 4819
rect 21004 4827 21043 4976
rect 20764 4811 20805 4812
rect 20088 4758 20125 4759
rect 20184 4758 20221 4759
rect 20240 4758 20276 4810
rect 20295 4758 20332 4759
rect 19988 4749 20126 4758
rect 19988 4729 20097 4749
rect 20117 4729 20126 4749
rect 19988 4722 20126 4729
rect 20184 4749 20332 4758
rect 20184 4729 20193 4749
rect 20213 4729 20303 4749
rect 20323 4729 20332 4749
rect 19988 4720 20084 4722
rect 20184 4719 20332 4729
rect 20391 4749 20428 4759
rect 20503 4758 20540 4759
rect 20484 4756 20540 4758
rect 20391 4729 20399 4749
rect 20419 4729 20428 4749
rect 20240 4718 20276 4719
rect 18153 4710 18184 4713
rect 18682 4713 18850 4714
rect 16982 4686 17120 4695
rect 18682 4687 19126 4713
rect 16776 4685 16813 4686
rect 16832 4634 16868 4686
rect 16887 4685 16924 4686
rect 16983 4685 17020 4686
rect 16303 4632 16344 4633
rect 15110 4610 15759 4616
rect 16195 4625 16344 4632
rect 15110 4609 15758 4610
rect 14176 4589 14187 4609
rect 14207 4589 14325 4609
rect 15721 4607 15758 4609
rect 16195 4605 16313 4625
rect 16333 4605 16344 4625
rect 16195 4597 16344 4605
rect 16411 4629 16770 4633
rect 16411 4624 16733 4629
rect 16411 4600 16524 4624
rect 16548 4605 16733 4624
rect 16757 4605 16770 4629
rect 16548 4600 16770 4605
rect 16411 4597 16770 4600
rect 16832 4597 16867 4634
rect 16935 4631 17035 4634
rect 16935 4627 17002 4631
rect 16935 4601 16947 4627
rect 16973 4605 17002 4627
rect 17028 4605 17035 4631
rect 16973 4601 17035 4605
rect 16935 4597 17035 4601
rect 14176 4582 14325 4589
rect 14176 4581 14217 4582
rect 13500 4528 13537 4529
rect 13596 4528 13633 4529
rect 13652 4528 13688 4580
rect 13707 4528 13744 4529
rect 11394 4501 11838 4527
rect 11395 4484 11419 4501
rect 11670 4500 11838 4501
rect 12289 4497 12539 4521
rect 10344 4436 10379 4479
rect 10793 4466 11420 4484
rect 10793 4465 10831 4466
rect 10339 4431 10379 4436
rect 10791 4460 10831 4465
rect 10339 4430 10377 4431
rect 9750 4412 10377 4430
rect 10791 4417 10826 4460
rect 8631 4375 8881 4399
rect 9332 4395 9500 4396
rect 9751 4395 9775 4412
rect 9332 4369 9776 4395
rect 7426 4367 7463 4368
rect 7482 4316 7518 4368
rect 7537 4367 7574 4368
rect 7633 4367 7670 4368
rect 6953 4314 6994 4315
rect 6845 4307 6994 4314
rect 4135 4295 4235 4299
rect 4135 4291 4197 4295
rect 4135 4265 4142 4291
rect 4168 4269 4197 4291
rect 4223 4269 4235 4295
rect 4168 4265 4235 4269
rect 4135 4262 4235 4265
rect 4303 4262 4338 4299
rect 4400 4296 4759 4299
rect 4400 4291 4622 4296
rect 4400 4267 4413 4291
rect 4437 4272 4622 4291
rect 4646 4272 4759 4296
rect 4437 4267 4759 4272
rect 4400 4263 4759 4267
rect 4826 4291 4975 4299
rect 4826 4271 4837 4291
rect 4857 4271 4975 4291
rect 5412 4287 5449 4289
rect 6845 4287 6963 4307
rect 6983 4287 6994 4307
rect 5412 4286 6060 4287
rect 4826 4264 4975 4271
rect 5411 4280 6060 4286
rect 4826 4263 4867 4264
rect 4150 4210 4187 4211
rect 4246 4210 4283 4211
rect 4302 4210 4338 4262
rect 4357 4210 4394 4211
rect 2044 4183 2488 4209
rect 4050 4201 4188 4210
rect 2320 4182 2488 4183
rect 2986 4183 3017 4186
rect 894 4177 930 4178
rect 742 4147 751 4167
rect 771 4147 779 4167
rect 630 4138 686 4140
rect 630 4137 667 4138
rect 742 4137 779 4147
rect 838 4167 986 4177
rect 1086 4174 1182 4176
rect 838 4147 847 4167
rect 867 4147 957 4167
rect 977 4147 986 4167
rect 838 4138 986 4147
rect 1044 4167 1182 4174
rect 1044 4147 1053 4167
rect 1073 4147 1182 4167
rect 1044 4138 1182 4147
rect 838 4137 875 4138
rect 894 4086 930 4138
rect 949 4137 986 4138
rect 1045 4137 1082 4138
rect 365 4084 406 4085
rect 127 3920 166 4069
rect 257 4077 406 4084
rect 257 4057 375 4077
rect 395 4057 406 4077
rect 257 4049 406 4057
rect 473 4081 832 4085
rect 473 4076 795 4081
rect 473 4052 586 4076
rect 610 4057 795 4076
rect 819 4057 832 4081
rect 610 4052 832 4057
rect 473 4049 832 4052
rect 894 4049 929 4086
rect 997 4083 1097 4086
rect 997 4079 1064 4083
rect 997 4053 1009 4079
rect 1035 4057 1064 4079
rect 1090 4057 1097 4083
rect 1035 4053 1097 4057
rect 997 4049 1097 4053
rect 473 4028 504 4049
rect 894 4028 930 4049
rect 316 4027 353 4028
rect 315 4018 353 4027
rect 315 3998 324 4018
rect 344 3998 353 4018
rect 315 3990 353 3998
rect 419 4022 504 4028
rect 529 4027 566 4028
rect 419 4002 427 4022
rect 447 4002 504 4022
rect 419 3994 504 4002
rect 528 4018 566 4027
rect 528 3998 537 4018
rect 557 3998 566 4018
rect 419 3993 455 3994
rect 528 3990 566 3998
rect 632 4022 717 4028
rect 737 4027 774 4028
rect 632 4002 640 4022
rect 660 4021 717 4022
rect 660 4002 689 4021
rect 632 4001 689 4002
rect 710 4001 717 4021
rect 632 3994 717 4001
rect 736 4018 774 4027
rect 736 3998 745 4018
rect 765 3998 774 4018
rect 632 3993 668 3994
rect 736 3990 774 3998
rect 840 4023 984 4028
rect 840 4022 905 4023
rect 840 4002 848 4022
rect 868 4002 905 4022
rect 927 4022 984 4023
rect 927 4002 956 4022
rect 976 4002 984 4022
rect 840 3994 984 4002
rect 840 3993 876 3994
rect 948 3993 984 3994
rect 1050 4027 1087 4028
rect 1050 4026 1088 4027
rect 1050 4018 1114 4026
rect 1050 3998 1059 4018
rect 1079 4004 1114 4018
rect 1134 4004 1137 4024
rect 1079 3999 1137 4004
rect 1079 3998 1114 3999
rect 316 3961 353 3990
rect 317 3959 353 3961
rect 529 3959 566 3990
rect 317 3937 566 3959
rect 737 3958 774 3990
rect 1050 3986 1114 3998
rect 1154 3960 1181 4138
rect 1013 3958 1181 3960
rect 737 3932 1181 3958
rect 1333 4057 1583 4081
rect 1333 3986 1370 4057
rect 1485 3996 1516 3997
rect 1333 3966 1342 3986
rect 1362 3966 1370 3986
rect 1333 3956 1370 3966
rect 1429 3986 1516 3996
rect 1429 3966 1438 3986
rect 1458 3966 1516 3986
rect 1429 3957 1516 3966
rect 1429 3956 1466 3957
rect 737 3922 759 3932
rect 1013 3931 1181 3932
rect 697 3920 759 3922
rect 127 3913 759 3920
rect 126 3904 759 3913
rect 1485 3904 1516 3957
rect 1546 3986 1583 4057
rect 1754 4062 2147 4082
rect 2167 4062 2170 4082
rect 1754 4057 2170 4062
rect 1754 4056 2095 4057
rect 1698 3996 1729 3997
rect 1546 3966 1555 3986
rect 1575 3966 1583 3986
rect 1546 3956 1583 3966
rect 1642 3989 1729 3996
rect 1642 3986 1703 3989
rect 1642 3966 1651 3986
rect 1671 3969 1703 3986
rect 1724 3969 1729 3989
rect 1671 3966 1729 3969
rect 1642 3959 1729 3966
rect 1754 3986 1791 4056
rect 2057 4055 2094 4056
rect 1906 3996 1942 3997
rect 1754 3966 1763 3986
rect 1783 3966 1791 3986
rect 1642 3957 1698 3959
rect 1642 3956 1679 3957
rect 1754 3956 1791 3966
rect 1850 3986 1998 3996
rect 2098 3993 2194 3995
rect 1850 3966 1859 3986
rect 1879 3966 1969 3986
rect 1989 3966 1998 3986
rect 1850 3957 1998 3966
rect 2056 3986 2194 3993
rect 2056 3966 2065 3986
rect 2085 3966 2194 3986
rect 2056 3957 2194 3966
rect 1850 3956 1887 3957
rect 1906 3905 1942 3957
rect 1961 3956 1998 3957
rect 2057 3956 2094 3957
rect 126 3886 136 3904
rect 154 3903 759 3904
rect 1377 3903 1418 3904
rect 154 3898 175 3903
rect 154 3886 166 3898
rect 1269 3896 1418 3903
rect 126 3878 166 3886
rect 209 3885 235 3886
rect 126 3876 163 3878
rect 209 3867 763 3885
rect 1269 3876 1387 3896
rect 1407 3876 1418 3896
rect 1269 3868 1418 3876
rect 1485 3900 1844 3904
rect 1485 3895 1807 3900
rect 1485 3871 1598 3895
rect 1622 3876 1807 3895
rect 1831 3876 1844 3900
rect 1622 3871 1844 3876
rect 1485 3868 1844 3871
rect 1906 3868 1941 3905
rect 2009 3902 2109 3905
rect 2009 3898 2076 3902
rect 2009 3872 2021 3898
rect 2047 3876 2076 3898
rect 2102 3876 2109 3902
rect 2047 3872 2109 3876
rect 2009 3868 2109 3872
rect 129 3808 166 3814
rect 209 3808 235 3867
rect 742 3848 763 3867
rect 129 3805 235 3808
rect 129 3787 138 3805
rect 156 3791 235 3805
rect 320 3823 570 3847
rect 156 3789 232 3791
rect 156 3787 166 3789
rect 129 3777 166 3787
rect 134 3712 165 3777
rect 320 3752 357 3823
rect 472 3762 503 3763
rect 320 3732 329 3752
rect 349 3732 357 3752
rect 320 3722 357 3732
rect 416 3752 503 3762
rect 416 3732 425 3752
rect 445 3732 503 3752
rect 416 3723 503 3732
rect 416 3722 453 3723
rect 133 3703 170 3712
rect 133 3685 143 3703
rect 161 3685 170 3703
rect 133 3675 170 3685
rect 472 3670 503 3723
rect 533 3752 570 3823
rect 741 3828 1134 3848
rect 1154 3828 1157 3848
rect 1485 3847 1516 3868
rect 1906 3847 1942 3868
rect 1328 3846 1365 3847
rect 741 3823 1157 3828
rect 1327 3837 1365 3846
rect 741 3822 1082 3823
rect 685 3762 716 3763
rect 533 3732 542 3752
rect 562 3732 570 3752
rect 533 3722 570 3732
rect 629 3755 716 3762
rect 629 3752 690 3755
rect 629 3732 638 3752
rect 658 3735 690 3752
rect 711 3735 716 3755
rect 658 3732 716 3735
rect 629 3725 716 3732
rect 741 3752 778 3822
rect 1044 3821 1081 3822
rect 1327 3817 1336 3837
rect 1356 3817 1365 3837
rect 1327 3809 1365 3817
rect 1431 3841 1516 3847
rect 1541 3846 1578 3847
rect 1431 3821 1439 3841
rect 1459 3821 1516 3841
rect 1431 3813 1516 3821
rect 1540 3837 1578 3846
rect 1540 3817 1549 3837
rect 1569 3817 1578 3837
rect 1431 3812 1467 3813
rect 1540 3809 1578 3817
rect 1644 3841 1729 3847
rect 1749 3846 1786 3847
rect 1644 3821 1652 3841
rect 1672 3840 1729 3841
rect 1672 3821 1701 3840
rect 1644 3820 1701 3821
rect 1722 3820 1729 3840
rect 1644 3813 1729 3820
rect 1748 3837 1786 3846
rect 1748 3817 1757 3837
rect 1777 3817 1786 3837
rect 1644 3812 1680 3813
rect 1748 3809 1786 3817
rect 1852 3841 1996 3847
rect 1852 3821 1860 3841
rect 1880 3821 1912 3841
rect 1936 3821 1968 3841
rect 1988 3821 1996 3841
rect 1852 3813 1996 3821
rect 1852 3812 1888 3813
rect 1960 3812 1996 3813
rect 2062 3846 2099 3847
rect 2062 3845 2100 3846
rect 2062 3837 2126 3845
rect 2062 3817 2071 3837
rect 2091 3823 2126 3837
rect 2146 3823 2149 3843
rect 2091 3818 2149 3823
rect 2091 3817 2126 3818
rect 1328 3780 1365 3809
rect 1329 3778 1365 3780
rect 1541 3778 1578 3809
rect 893 3762 929 3763
rect 741 3732 750 3752
rect 770 3732 778 3752
rect 629 3723 685 3725
rect 629 3722 666 3723
rect 741 3722 778 3732
rect 837 3752 985 3762
rect 1085 3759 1181 3761
rect 837 3732 846 3752
rect 866 3732 956 3752
rect 976 3732 985 3752
rect 837 3723 985 3732
rect 1043 3752 1181 3759
rect 1329 3756 1578 3778
rect 1749 3777 1786 3809
rect 2062 3805 2126 3817
rect 2166 3779 2193 3957
rect 2025 3777 2193 3779
rect 1749 3773 2193 3777
rect 1043 3732 1052 3752
rect 1072 3732 1181 3752
rect 1749 3754 1798 3773
rect 1818 3754 2193 3773
rect 1749 3751 2193 3754
rect 2025 3750 2193 3751
rect 1043 3723 1181 3732
rect 837 3722 874 3723
rect 893 3671 929 3723
rect 948 3722 985 3723
rect 1044 3722 1081 3723
rect 364 3669 405 3670
rect 256 3662 405 3669
rect 256 3642 374 3662
rect 394 3642 405 3662
rect 256 3634 405 3642
rect 472 3666 831 3670
rect 472 3661 794 3666
rect 472 3637 585 3661
rect 609 3642 794 3661
rect 818 3642 831 3666
rect 609 3637 831 3642
rect 472 3634 831 3637
rect 893 3634 928 3671
rect 996 3668 1096 3671
rect 996 3664 1063 3668
rect 996 3638 1008 3664
rect 1034 3642 1063 3664
rect 1089 3642 1096 3668
rect 1034 3638 1096 3642
rect 996 3634 1096 3638
rect 472 3613 503 3634
rect 893 3613 929 3634
rect 136 3604 173 3613
rect 315 3612 352 3613
rect 136 3586 145 3604
rect 163 3586 173 3604
rect 136 3576 173 3586
rect 137 3541 173 3576
rect 314 3603 352 3612
rect 314 3583 323 3603
rect 343 3583 352 3603
rect 314 3575 352 3583
rect 418 3607 503 3613
rect 528 3612 565 3613
rect 418 3587 426 3607
rect 446 3587 503 3607
rect 418 3579 503 3587
rect 527 3603 565 3612
rect 527 3583 536 3603
rect 556 3583 565 3603
rect 418 3578 454 3579
rect 527 3575 565 3583
rect 631 3607 716 3613
rect 736 3612 773 3613
rect 631 3587 639 3607
rect 659 3606 716 3607
rect 659 3587 688 3606
rect 631 3586 688 3587
rect 709 3586 716 3606
rect 631 3579 716 3586
rect 735 3603 773 3612
rect 735 3583 744 3603
rect 764 3583 773 3603
rect 631 3578 667 3579
rect 735 3575 773 3583
rect 839 3607 983 3613
rect 839 3587 847 3607
rect 867 3606 955 3607
rect 867 3587 895 3606
rect 839 3585 895 3587
rect 917 3587 955 3606
rect 975 3587 983 3607
rect 917 3585 983 3587
rect 839 3579 983 3585
rect 839 3578 875 3579
rect 947 3578 983 3579
rect 1049 3612 1086 3613
rect 1049 3611 1087 3612
rect 1049 3603 1113 3611
rect 1049 3583 1058 3603
rect 1078 3589 1113 3603
rect 1133 3589 1136 3609
rect 1078 3584 1136 3589
rect 1078 3583 1113 3584
rect 315 3546 352 3575
rect 135 3500 173 3541
rect 316 3544 352 3546
rect 528 3544 565 3575
rect 316 3522 565 3544
rect 736 3543 773 3575
rect 1049 3571 1113 3583
rect 1153 3545 1180 3723
rect 1012 3543 1180 3545
rect 736 3517 1180 3543
rect 737 3500 761 3517
rect 1012 3516 1180 3517
rect 135 3482 762 3500
rect 1388 3496 1638 3520
rect 135 3476 173 3482
rect 135 3452 172 3476
rect 135 3428 170 3452
rect 133 3419 170 3428
rect 133 3401 143 3419
rect 161 3401 170 3419
rect 133 3391 170 3401
rect 1388 3425 1425 3496
rect 1540 3435 1571 3436
rect 1388 3405 1397 3425
rect 1417 3405 1425 3425
rect 1388 3395 1425 3405
rect 1484 3425 1571 3435
rect 1484 3405 1493 3425
rect 1513 3405 1571 3425
rect 1484 3396 1571 3405
rect 1484 3395 1521 3396
rect 1540 3343 1571 3396
rect 1601 3425 1638 3496
rect 1809 3501 2202 3521
rect 2222 3501 2225 3521
rect 1809 3496 2225 3501
rect 1809 3495 2150 3496
rect 1753 3435 1784 3436
rect 1601 3405 1610 3425
rect 1630 3405 1638 3425
rect 1601 3395 1638 3405
rect 1697 3428 1784 3435
rect 1697 3425 1758 3428
rect 1697 3405 1706 3425
rect 1726 3408 1758 3425
rect 1779 3408 1784 3428
rect 1726 3405 1784 3408
rect 1697 3398 1784 3405
rect 1809 3425 1846 3495
rect 2112 3494 2149 3495
rect 1961 3435 1997 3436
rect 1809 3405 1818 3425
rect 1838 3405 1846 3425
rect 1697 3396 1753 3398
rect 1697 3395 1734 3396
rect 1809 3395 1846 3405
rect 1905 3425 2053 3435
rect 2153 3432 2249 3434
rect 1905 3405 1914 3425
rect 1934 3405 2024 3425
rect 2044 3405 2053 3425
rect 1905 3396 2053 3405
rect 2111 3425 2249 3432
rect 2111 3405 2120 3425
rect 2140 3405 2249 3425
rect 2111 3396 2249 3405
rect 1905 3395 1942 3396
rect 1961 3344 1997 3396
rect 2016 3395 2053 3396
rect 2112 3395 2149 3396
rect 1432 3342 1473 3343
rect 1324 3335 1473 3342
rect 136 3327 173 3329
rect 136 3326 784 3327
rect 135 3320 784 3326
rect 135 3302 145 3320
rect 163 3306 784 3320
rect 1324 3315 1442 3335
rect 1462 3315 1473 3335
rect 1324 3307 1473 3315
rect 1540 3339 1899 3343
rect 1540 3334 1862 3339
rect 1540 3310 1653 3334
rect 1677 3315 1862 3334
rect 1886 3315 1899 3339
rect 1677 3310 1899 3315
rect 1540 3307 1899 3310
rect 1961 3307 1996 3344
rect 2064 3341 2164 3344
rect 2064 3337 2131 3341
rect 2064 3311 2076 3337
rect 2102 3315 2131 3337
rect 2157 3315 2164 3341
rect 2102 3311 2164 3315
rect 2064 3307 2164 3311
rect 163 3302 173 3306
rect 614 3305 784 3306
rect 135 3292 173 3302
rect 135 3214 170 3292
rect 747 3282 784 3305
rect 1540 3286 1571 3307
rect 1961 3286 1997 3307
rect 1383 3285 1420 3286
rect 131 3205 170 3214
rect 131 3187 141 3205
rect 159 3187 170 3205
rect 131 3181 170 3187
rect 326 3257 576 3281
rect 326 3186 363 3257
rect 478 3196 509 3197
rect 131 3177 168 3181
rect 326 3166 335 3186
rect 355 3166 363 3186
rect 326 3156 363 3166
rect 422 3186 509 3196
rect 422 3166 431 3186
rect 451 3166 509 3186
rect 422 3157 509 3166
rect 422 3156 459 3157
rect 134 3106 171 3115
rect 132 3088 143 3106
rect 161 3088 171 3106
rect 478 3104 509 3157
rect 539 3186 576 3257
rect 747 3262 1140 3282
rect 1160 3262 1163 3282
rect 747 3257 1163 3262
rect 1382 3276 1420 3285
rect 747 3256 1088 3257
rect 1382 3256 1391 3276
rect 1411 3256 1420 3276
rect 691 3196 722 3197
rect 539 3166 548 3186
rect 568 3166 576 3186
rect 539 3156 576 3166
rect 635 3189 722 3196
rect 635 3186 696 3189
rect 635 3166 644 3186
rect 664 3169 696 3186
rect 717 3169 722 3189
rect 664 3166 722 3169
rect 635 3159 722 3166
rect 747 3186 784 3256
rect 1050 3255 1087 3256
rect 1382 3248 1420 3256
rect 1486 3280 1571 3286
rect 1596 3285 1633 3286
rect 1486 3260 1494 3280
rect 1514 3260 1571 3280
rect 1486 3252 1571 3260
rect 1595 3276 1633 3285
rect 1595 3256 1604 3276
rect 1624 3256 1633 3276
rect 1486 3251 1522 3252
rect 1595 3248 1633 3256
rect 1699 3280 1784 3286
rect 1804 3285 1841 3286
rect 1699 3260 1707 3280
rect 1727 3279 1784 3280
rect 1727 3260 1756 3279
rect 1699 3259 1756 3260
rect 1777 3259 1784 3279
rect 1699 3252 1784 3259
rect 1803 3276 1841 3285
rect 1803 3256 1812 3276
rect 1832 3256 1841 3276
rect 1699 3251 1735 3252
rect 1803 3248 1841 3256
rect 1907 3280 2051 3286
rect 1907 3260 1915 3280
rect 1935 3278 2023 3280
rect 1935 3261 1971 3278
rect 1995 3261 2023 3278
rect 1935 3260 2023 3261
rect 2043 3260 2051 3280
rect 1907 3252 2051 3260
rect 1907 3251 1943 3252
rect 2015 3251 2051 3252
rect 2117 3285 2154 3286
rect 2117 3284 2155 3285
rect 2117 3276 2181 3284
rect 2117 3256 2126 3276
rect 2146 3262 2181 3276
rect 2201 3262 2204 3282
rect 2146 3257 2204 3262
rect 2146 3256 2181 3257
rect 1383 3219 1420 3248
rect 1384 3217 1420 3219
rect 1596 3217 1633 3248
rect 899 3196 935 3197
rect 747 3166 756 3186
rect 776 3166 784 3186
rect 635 3157 691 3159
rect 635 3156 672 3157
rect 747 3156 784 3166
rect 843 3186 991 3196
rect 1384 3195 1633 3217
rect 1804 3216 1841 3248
rect 2117 3244 2181 3256
rect 2221 3218 2248 3396
rect 2080 3216 2248 3218
rect 1804 3205 2248 3216
rect 1091 3193 1187 3195
rect 843 3166 852 3186
rect 872 3166 962 3186
rect 982 3166 991 3186
rect 843 3157 991 3166
rect 1049 3186 1187 3193
rect 1804 3190 2250 3205
rect 2080 3189 2250 3190
rect 1049 3166 1058 3186
rect 1078 3166 1187 3186
rect 1049 3157 1187 3166
rect 843 3156 880 3157
rect 899 3105 935 3157
rect 954 3156 991 3157
rect 1050 3156 1087 3157
rect 370 3103 411 3104
rect 132 2939 171 3088
rect 262 3096 411 3103
rect 262 3076 380 3096
rect 400 3076 411 3096
rect 262 3068 411 3076
rect 478 3100 837 3104
rect 478 3095 800 3100
rect 478 3071 591 3095
rect 615 3076 800 3095
rect 824 3076 837 3100
rect 615 3071 837 3076
rect 478 3068 837 3071
rect 899 3068 934 3105
rect 1002 3102 1102 3105
rect 1002 3098 1069 3102
rect 1002 3072 1014 3098
rect 1040 3076 1069 3098
rect 1095 3076 1102 3102
rect 1040 3072 1102 3076
rect 1002 3068 1102 3072
rect 478 3047 509 3068
rect 899 3047 935 3068
rect 321 3046 358 3047
rect 320 3037 358 3046
rect 320 3017 329 3037
rect 349 3017 358 3037
rect 320 3009 358 3017
rect 424 3041 509 3047
rect 534 3046 571 3047
rect 424 3021 432 3041
rect 452 3021 509 3041
rect 424 3013 509 3021
rect 533 3037 571 3046
rect 533 3017 542 3037
rect 562 3017 571 3037
rect 424 3012 460 3013
rect 533 3009 571 3017
rect 637 3041 722 3047
rect 742 3046 779 3047
rect 637 3021 645 3041
rect 665 3040 722 3041
rect 665 3021 694 3040
rect 637 3020 694 3021
rect 715 3020 722 3040
rect 637 3013 722 3020
rect 741 3037 779 3046
rect 741 3017 750 3037
rect 770 3017 779 3037
rect 637 3012 673 3013
rect 741 3009 779 3017
rect 845 3042 989 3047
rect 845 3041 910 3042
rect 845 3021 853 3041
rect 873 3021 910 3041
rect 932 3041 989 3042
rect 932 3021 961 3041
rect 981 3021 989 3041
rect 845 3013 989 3021
rect 845 3012 881 3013
rect 953 3012 989 3013
rect 1055 3046 1092 3047
rect 1055 3045 1093 3046
rect 1055 3037 1119 3045
rect 1055 3017 1064 3037
rect 1084 3023 1119 3037
rect 1139 3023 1142 3043
rect 1084 3018 1142 3023
rect 1084 3017 1119 3018
rect 321 2980 358 3009
rect 322 2978 358 2980
rect 534 2978 571 3009
rect 322 2956 571 2978
rect 742 2977 779 3009
rect 1055 3005 1119 3017
rect 1159 2979 1186 3157
rect 1018 2977 1186 2979
rect 742 2951 1186 2977
rect 1338 3076 1588 3100
rect 1338 3005 1375 3076
rect 1490 3015 1521 3016
rect 1338 2985 1347 3005
rect 1367 2985 1375 3005
rect 1338 2975 1375 2985
rect 1434 3005 1521 3015
rect 1434 2985 1443 3005
rect 1463 2985 1521 3005
rect 1434 2976 1521 2985
rect 1434 2975 1471 2976
rect 742 2941 764 2951
rect 1018 2950 1186 2951
rect 702 2939 764 2941
rect 132 2932 764 2939
rect 131 2923 764 2932
rect 1490 2923 1521 2976
rect 1551 3005 1588 3076
rect 1759 3081 2152 3101
rect 2172 3081 2175 3101
rect 1759 3076 2175 3081
rect 1759 3075 2100 3076
rect 1703 3015 1734 3016
rect 1551 2985 1560 3005
rect 1580 2985 1588 3005
rect 1551 2975 1588 2985
rect 1647 3008 1734 3015
rect 1647 3005 1708 3008
rect 1647 2985 1656 3005
rect 1676 2988 1708 3005
rect 1729 2988 1734 3008
rect 1676 2985 1734 2988
rect 1647 2978 1734 2985
rect 1759 3005 1796 3075
rect 2062 3074 2099 3075
rect 1911 3015 1947 3016
rect 1759 2985 1768 3005
rect 1788 2985 1796 3005
rect 1647 2976 1703 2978
rect 1647 2975 1684 2976
rect 1759 2975 1796 2985
rect 1855 3005 2003 3015
rect 2103 3012 2199 3014
rect 1855 2985 1864 3005
rect 1884 2985 1974 3005
rect 1994 2985 2003 3005
rect 1855 2976 2003 2985
rect 2061 3005 2199 3012
rect 2061 2985 2070 3005
rect 2090 2985 2199 3005
rect 2061 2976 2199 2985
rect 1855 2975 1892 2976
rect 1911 2924 1947 2976
rect 1966 2975 2003 2976
rect 2062 2975 2099 2976
rect 131 2905 141 2923
rect 159 2922 764 2923
rect 1382 2922 1423 2923
rect 159 2917 180 2922
rect 159 2905 171 2917
rect 1274 2915 1423 2922
rect 131 2897 171 2905
rect 214 2904 240 2905
rect 131 2895 168 2897
rect 214 2886 768 2904
rect 1274 2895 1392 2915
rect 1412 2895 1423 2915
rect 1274 2887 1423 2895
rect 1490 2919 1849 2923
rect 1490 2914 1812 2919
rect 1490 2890 1603 2914
rect 1627 2895 1812 2914
rect 1836 2895 1849 2919
rect 1627 2890 1849 2895
rect 1490 2887 1849 2890
rect 1911 2887 1946 2924
rect 2014 2921 2114 2924
rect 2014 2917 2081 2921
rect 2014 2891 2026 2917
rect 2052 2895 2081 2917
rect 2107 2895 2114 2921
rect 2052 2891 2114 2895
rect 2014 2887 2114 2891
rect 134 2827 171 2833
rect 214 2827 240 2886
rect 747 2867 768 2886
rect 134 2824 240 2827
rect 134 2806 143 2824
rect 161 2810 240 2824
rect 325 2842 575 2866
rect 161 2808 237 2810
rect 161 2806 171 2808
rect 134 2796 171 2806
rect 139 2731 170 2796
rect 325 2771 362 2842
rect 477 2781 508 2782
rect 325 2751 334 2771
rect 354 2751 362 2771
rect 325 2741 362 2751
rect 421 2771 508 2781
rect 421 2751 430 2771
rect 450 2751 508 2771
rect 421 2742 508 2751
rect 421 2741 458 2742
rect 138 2722 175 2731
rect 138 2704 148 2722
rect 166 2704 175 2722
rect 138 2694 175 2704
rect 477 2689 508 2742
rect 538 2771 575 2842
rect 746 2847 1139 2867
rect 1159 2847 1162 2867
rect 1490 2866 1521 2887
rect 1911 2866 1947 2887
rect 1333 2865 1370 2866
rect 746 2842 1162 2847
rect 1332 2856 1370 2865
rect 746 2841 1087 2842
rect 690 2781 721 2782
rect 538 2751 547 2771
rect 567 2751 575 2771
rect 538 2741 575 2751
rect 634 2774 721 2781
rect 634 2771 695 2774
rect 634 2751 643 2771
rect 663 2754 695 2771
rect 716 2754 721 2774
rect 663 2751 721 2754
rect 634 2744 721 2751
rect 746 2771 783 2841
rect 1049 2840 1086 2841
rect 1332 2836 1341 2856
rect 1361 2836 1370 2856
rect 1332 2828 1370 2836
rect 1436 2860 1521 2866
rect 1546 2865 1583 2866
rect 1436 2840 1444 2860
rect 1464 2840 1521 2860
rect 1436 2832 1521 2840
rect 1545 2856 1583 2865
rect 1545 2836 1554 2856
rect 1574 2836 1583 2856
rect 1436 2831 1472 2832
rect 1545 2828 1583 2836
rect 1649 2860 1734 2866
rect 1754 2865 1791 2866
rect 1649 2840 1657 2860
rect 1677 2859 1734 2860
rect 1677 2840 1706 2859
rect 1649 2839 1706 2840
rect 1727 2839 1734 2859
rect 1649 2832 1734 2839
rect 1753 2856 1791 2865
rect 1753 2836 1762 2856
rect 1782 2836 1791 2856
rect 1649 2831 1685 2832
rect 1753 2828 1791 2836
rect 1857 2861 2001 2866
rect 1857 2860 1916 2861
rect 1857 2840 1865 2860
rect 1885 2841 1916 2860
rect 1940 2860 2001 2861
rect 1940 2841 1973 2860
rect 1885 2840 1973 2841
rect 1993 2840 2001 2860
rect 1857 2832 2001 2840
rect 1857 2831 1893 2832
rect 1965 2831 2001 2832
rect 2067 2865 2104 2866
rect 2067 2864 2105 2865
rect 2067 2856 2131 2864
rect 2067 2836 2076 2856
rect 2096 2842 2131 2856
rect 2151 2842 2154 2862
rect 2096 2837 2154 2842
rect 2096 2836 2131 2837
rect 1333 2799 1370 2828
rect 1334 2797 1370 2799
rect 1546 2797 1583 2828
rect 898 2781 934 2782
rect 746 2751 755 2771
rect 775 2751 783 2771
rect 634 2742 690 2744
rect 634 2741 671 2742
rect 746 2741 783 2751
rect 842 2771 990 2781
rect 1090 2778 1186 2780
rect 842 2751 851 2771
rect 871 2751 961 2771
rect 981 2751 990 2771
rect 842 2742 990 2751
rect 1048 2771 1186 2778
rect 1334 2775 1583 2797
rect 1754 2796 1791 2828
rect 2067 2824 2131 2836
rect 2171 2798 2198 2976
rect 2030 2796 2198 2798
rect 1754 2792 2198 2796
rect 1048 2751 1057 2771
rect 1077 2751 1186 2771
rect 1754 2773 1803 2792
rect 1823 2773 2198 2792
rect 1754 2770 2198 2773
rect 2030 2769 2198 2770
rect 2219 2795 2250 3189
rect 2219 2769 2224 2795
rect 2243 2769 2250 2795
rect 2219 2766 2250 2769
rect 1048 2742 1186 2751
rect 842 2741 879 2742
rect 898 2690 934 2742
rect 953 2741 990 2742
rect 1049 2741 1086 2742
rect 369 2688 410 2689
rect 261 2681 410 2688
rect 261 2661 379 2681
rect 399 2661 410 2681
rect 261 2653 410 2661
rect 477 2685 836 2689
rect 477 2680 799 2685
rect 477 2656 590 2680
rect 614 2661 799 2680
rect 823 2661 836 2685
rect 614 2656 836 2661
rect 477 2653 836 2656
rect 898 2653 933 2690
rect 1001 2687 1101 2690
rect 1001 2683 1068 2687
rect 1001 2657 1013 2683
rect 1039 2661 1068 2683
rect 1094 2661 1101 2687
rect 1039 2657 1101 2661
rect 1001 2653 1101 2657
rect 477 2632 508 2653
rect 898 2632 934 2653
rect 141 2623 178 2632
rect 320 2631 357 2632
rect 141 2605 150 2623
rect 168 2605 178 2623
rect 141 2595 178 2605
rect 142 2560 178 2595
rect 319 2622 357 2631
rect 319 2602 328 2622
rect 348 2602 357 2622
rect 319 2594 357 2602
rect 423 2626 508 2632
rect 533 2631 570 2632
rect 423 2606 431 2626
rect 451 2606 508 2626
rect 423 2598 508 2606
rect 532 2622 570 2631
rect 532 2602 541 2622
rect 561 2602 570 2622
rect 423 2597 459 2598
rect 532 2594 570 2602
rect 636 2626 721 2632
rect 741 2631 778 2632
rect 636 2606 644 2626
rect 664 2625 721 2626
rect 664 2606 693 2625
rect 636 2605 693 2606
rect 714 2605 721 2625
rect 636 2598 721 2605
rect 740 2622 778 2631
rect 740 2602 749 2622
rect 769 2602 778 2622
rect 636 2597 672 2598
rect 740 2594 778 2602
rect 844 2626 988 2632
rect 844 2606 852 2626
rect 872 2625 960 2626
rect 872 2606 900 2625
rect 844 2604 900 2606
rect 922 2606 960 2625
rect 980 2606 988 2626
rect 922 2604 988 2606
rect 844 2598 988 2604
rect 844 2597 880 2598
rect 952 2597 988 2598
rect 1054 2631 1091 2632
rect 1054 2630 1092 2631
rect 1054 2622 1118 2630
rect 1054 2602 1063 2622
rect 1083 2608 1118 2622
rect 1138 2608 1141 2628
rect 1083 2603 1141 2608
rect 1083 2602 1118 2603
rect 320 2565 357 2594
rect 140 2519 178 2560
rect 321 2563 357 2565
rect 533 2563 570 2594
rect 321 2541 570 2563
rect 741 2562 778 2594
rect 1054 2590 1118 2602
rect 1158 2564 1185 2742
rect 1017 2562 1185 2564
rect 741 2536 1185 2562
rect 742 2519 766 2536
rect 1017 2535 1185 2536
rect 1553 2564 1803 2588
rect 140 2501 767 2519
rect 140 2495 178 2501
rect 142 2449 177 2495
rect 1553 2493 1590 2564
rect 1705 2503 1736 2504
rect 1553 2473 1562 2493
rect 1582 2473 1590 2493
rect 1553 2463 1590 2473
rect 1649 2493 1736 2503
rect 1649 2473 1658 2493
rect 1678 2473 1736 2493
rect 1649 2464 1736 2473
rect 1649 2463 1686 2464
rect 140 2440 177 2449
rect 140 2422 150 2440
rect 168 2422 177 2440
rect 140 2412 177 2422
rect 1705 2411 1736 2464
rect 1766 2493 1803 2564
rect 1974 2569 2367 2589
rect 2387 2569 2390 2589
rect 1974 2564 2390 2569
rect 1974 2563 2315 2564
rect 1918 2503 1949 2504
rect 1766 2473 1775 2493
rect 1795 2473 1803 2493
rect 1766 2463 1803 2473
rect 1862 2496 1949 2503
rect 1862 2493 1923 2496
rect 1862 2473 1871 2493
rect 1891 2476 1923 2493
rect 1944 2476 1949 2496
rect 1891 2473 1949 2476
rect 1862 2466 1949 2473
rect 1974 2493 2011 2563
rect 2277 2562 2314 2563
rect 2126 2503 2162 2504
rect 1974 2473 1983 2493
rect 2003 2473 2011 2493
rect 1862 2464 1918 2466
rect 1862 2463 1899 2464
rect 1974 2463 2011 2473
rect 2070 2493 2218 2503
rect 2318 2500 2414 2502
rect 2070 2473 2079 2493
rect 2099 2473 2189 2493
rect 2209 2473 2218 2493
rect 2070 2464 2218 2473
rect 2276 2493 2414 2500
rect 2276 2473 2285 2493
rect 2305 2473 2414 2493
rect 2276 2464 2414 2473
rect 2070 2463 2107 2464
rect 2126 2412 2162 2464
rect 2181 2463 2218 2464
rect 2277 2463 2314 2464
rect 1597 2410 1638 2411
rect 1489 2403 1638 2410
rect 1489 2383 1607 2403
rect 1627 2383 1638 2403
rect 1489 2375 1638 2383
rect 1705 2407 2064 2411
rect 1705 2402 2027 2407
rect 1705 2378 1818 2402
rect 1842 2383 2027 2402
rect 2051 2383 2064 2407
rect 1842 2378 2064 2383
rect 1705 2375 2064 2378
rect 2126 2375 2161 2412
rect 2229 2409 2329 2412
rect 2229 2405 2296 2409
rect 2229 2379 2241 2405
rect 2267 2383 2296 2405
rect 2322 2383 2329 2409
rect 2267 2379 2329 2383
rect 2229 2375 2329 2379
rect 1705 2354 1736 2375
rect 2126 2354 2162 2375
rect 1548 2353 1585 2354
rect 143 2348 180 2350
rect 143 2347 791 2348
rect 142 2341 791 2347
rect 142 2323 152 2341
rect 170 2327 791 2341
rect 170 2323 180 2327
rect 621 2326 791 2327
rect 142 2313 180 2323
rect 142 2235 177 2313
rect 754 2303 791 2326
rect 1547 2344 1585 2353
rect 1547 2324 1556 2344
rect 1576 2324 1585 2344
rect 1547 2316 1585 2324
rect 1651 2348 1736 2354
rect 1761 2353 1798 2354
rect 1651 2328 1659 2348
rect 1679 2328 1736 2348
rect 1651 2320 1736 2328
rect 1760 2344 1798 2353
rect 1760 2324 1769 2344
rect 1789 2324 1798 2344
rect 1651 2319 1687 2320
rect 1760 2316 1798 2324
rect 1864 2348 1949 2354
rect 1969 2353 2006 2354
rect 1864 2328 1872 2348
rect 1892 2347 1949 2348
rect 1892 2328 1921 2347
rect 1864 2327 1921 2328
rect 1942 2327 1949 2347
rect 1864 2320 1949 2327
rect 1968 2344 2006 2353
rect 1968 2324 1977 2344
rect 1997 2324 2006 2344
rect 1864 2319 1900 2320
rect 1968 2316 2006 2324
rect 2072 2348 2216 2354
rect 2072 2328 2080 2348
rect 2100 2329 2136 2348
rect 2159 2329 2188 2348
rect 2100 2328 2188 2329
rect 2208 2328 2216 2348
rect 2072 2320 2216 2328
rect 2072 2319 2108 2320
rect 2180 2319 2216 2320
rect 2282 2353 2319 2354
rect 2282 2352 2320 2353
rect 2282 2344 2346 2352
rect 2282 2324 2291 2344
rect 2311 2330 2346 2344
rect 2366 2330 2369 2350
rect 2311 2325 2369 2330
rect 2311 2324 2346 2325
rect 138 2226 177 2235
rect 138 2208 148 2226
rect 166 2208 177 2226
rect 138 2202 177 2208
rect 333 2278 583 2302
rect 333 2207 370 2278
rect 485 2217 516 2218
rect 138 2198 175 2202
rect 333 2187 342 2207
rect 362 2187 370 2207
rect 333 2177 370 2187
rect 429 2207 516 2217
rect 429 2187 438 2207
rect 458 2187 516 2207
rect 429 2178 516 2187
rect 429 2177 466 2178
rect 141 2127 178 2136
rect 139 2109 150 2127
rect 168 2109 178 2127
rect 485 2125 516 2178
rect 546 2207 583 2278
rect 754 2283 1147 2303
rect 1167 2283 1170 2303
rect 1548 2287 1585 2316
rect 754 2278 1170 2283
rect 1549 2285 1585 2287
rect 1761 2285 1798 2316
rect 754 2277 1095 2278
rect 698 2217 729 2218
rect 546 2187 555 2207
rect 575 2187 583 2207
rect 546 2177 583 2187
rect 642 2210 729 2217
rect 642 2207 703 2210
rect 642 2187 651 2207
rect 671 2190 703 2207
rect 724 2190 729 2210
rect 671 2187 729 2190
rect 642 2180 729 2187
rect 754 2207 791 2277
rect 1057 2276 1094 2277
rect 1549 2263 1798 2285
rect 1969 2284 2006 2316
rect 2282 2312 2346 2324
rect 2386 2286 2413 2464
rect 2441 2351 2479 4182
rect 2986 4157 2993 4183
rect 3012 4157 3017 4183
rect 2893 3764 2922 3766
rect 2893 3759 2925 3764
rect 2893 3741 2900 3759
rect 2920 3741 2925 3759
rect 2986 3763 3017 4157
rect 3038 4182 3206 4183
rect 3038 4179 3482 4182
rect 3038 4160 3413 4179
rect 3433 4160 3482 4179
rect 4050 4181 4159 4201
rect 4179 4181 4188 4201
rect 3038 4156 3482 4160
rect 3038 4154 3206 4156
rect 3038 3976 3065 4154
rect 3105 4116 3169 4128
rect 3445 4124 3482 4156
rect 3653 4155 3902 4177
rect 4050 4174 4188 4181
rect 4246 4201 4394 4210
rect 4246 4181 4255 4201
rect 4275 4181 4365 4201
rect 4385 4181 4394 4201
rect 4050 4172 4146 4174
rect 4246 4171 4394 4181
rect 4453 4201 4490 4211
rect 4565 4210 4602 4211
rect 4546 4208 4602 4210
rect 4453 4181 4461 4201
rect 4481 4181 4490 4201
rect 4302 4170 4338 4171
rect 3653 4124 3690 4155
rect 3866 4153 3902 4155
rect 3866 4124 3903 4153
rect 3105 4115 3140 4116
rect 3082 4110 3140 4115
rect 3082 4090 3085 4110
rect 3105 4096 3140 4110
rect 3160 4096 3169 4116
rect 3105 4088 3169 4096
rect 3131 4087 3169 4088
rect 3132 4086 3169 4087
rect 3235 4120 3271 4121
rect 3343 4120 3379 4121
rect 3235 4112 3379 4120
rect 3235 4092 3243 4112
rect 3263 4111 3351 4112
rect 3263 4092 3296 4111
rect 3235 4091 3296 4092
rect 3320 4092 3351 4111
rect 3371 4092 3379 4112
rect 3320 4091 3379 4092
rect 3235 4086 3379 4091
rect 3445 4116 3483 4124
rect 3551 4120 3587 4121
rect 3445 4096 3454 4116
rect 3474 4096 3483 4116
rect 3445 4087 3483 4096
rect 3502 4113 3587 4120
rect 3502 4093 3509 4113
rect 3530 4112 3587 4113
rect 3530 4093 3559 4112
rect 3502 4092 3559 4093
rect 3579 4092 3587 4112
rect 3445 4086 3482 4087
rect 3502 4086 3587 4092
rect 3653 4116 3691 4124
rect 3764 4120 3800 4121
rect 3653 4096 3662 4116
rect 3682 4096 3691 4116
rect 3653 4087 3691 4096
rect 3715 4112 3800 4120
rect 3715 4092 3772 4112
rect 3792 4092 3800 4112
rect 3653 4086 3690 4087
rect 3715 4086 3800 4092
rect 3866 4116 3904 4124
rect 3866 4096 3875 4116
rect 3895 4096 3904 4116
rect 4150 4111 4187 4112
rect 4453 4111 4490 4181
rect 4515 4201 4602 4208
rect 4515 4198 4573 4201
rect 4515 4178 4520 4198
rect 4541 4181 4573 4198
rect 4593 4181 4602 4201
rect 4541 4178 4602 4181
rect 4515 4171 4602 4178
rect 4661 4201 4698 4211
rect 4661 4181 4669 4201
rect 4689 4181 4698 4201
rect 4515 4170 4546 4171
rect 4149 4110 4490 4111
rect 3866 4087 3904 4096
rect 4074 4105 4490 4110
rect 3866 4086 3903 4087
rect 3289 4065 3325 4086
rect 3715 4065 3746 4086
rect 4074 4085 4077 4105
rect 4097 4085 4490 4105
rect 4661 4110 4698 4181
rect 4728 4210 4759 4263
rect 5411 4262 5421 4280
rect 5439 4266 6060 4280
rect 6845 4279 6994 4287
rect 7061 4311 7420 4315
rect 7061 4306 7383 4311
rect 7061 4282 7174 4306
rect 7198 4287 7383 4306
rect 7407 4287 7420 4311
rect 7198 4282 7420 4287
rect 7061 4279 7420 4282
rect 7482 4279 7517 4316
rect 7585 4313 7685 4316
rect 7585 4309 7652 4313
rect 7585 4283 7597 4309
rect 7623 4287 7652 4309
rect 7678 4287 7685 4313
rect 7623 4283 7685 4287
rect 7585 4279 7685 4283
rect 5439 4262 5449 4266
rect 5890 4265 6060 4266
rect 5061 4248 5098 4258
rect 5061 4230 5070 4248
rect 5088 4230 5098 4248
rect 5061 4221 5098 4230
rect 5411 4252 5449 4262
rect 4778 4210 4815 4211
rect 4728 4201 4815 4210
rect 4728 4181 4786 4201
rect 4806 4181 4815 4201
rect 4728 4171 4815 4181
rect 4874 4201 4911 4211
rect 4874 4181 4882 4201
rect 4902 4181 4911 4201
rect 4728 4170 4759 4171
rect 4874 4110 4911 4181
rect 5066 4156 5097 4221
rect 5411 4174 5446 4252
rect 6023 4242 6060 4265
rect 7061 4258 7092 4279
rect 7482 4258 7518 4279
rect 6904 4257 6941 4258
rect 6903 4248 6941 4257
rect 5407 4165 5446 4174
rect 5065 4146 5102 4156
rect 5065 4144 5075 4146
rect 4999 4142 5075 4144
rect 4661 4086 4911 4110
rect 4996 4128 5075 4142
rect 5093 4128 5102 4146
rect 5407 4147 5417 4165
rect 5435 4147 5446 4165
rect 5407 4141 5446 4147
rect 5602 4217 5852 4241
rect 5602 4146 5639 4217
rect 5754 4156 5785 4157
rect 5407 4137 5444 4141
rect 4996 4125 5102 4128
rect 4468 4066 4489 4085
rect 4996 4066 5022 4125
rect 5065 4119 5102 4125
rect 5602 4126 5611 4146
rect 5631 4126 5639 4146
rect 5602 4116 5639 4126
rect 5698 4146 5785 4156
rect 5698 4126 5707 4146
rect 5727 4126 5785 4146
rect 5698 4117 5785 4126
rect 5698 4116 5735 4117
rect 5410 4066 5447 4075
rect 3122 4061 3222 4065
rect 3122 4057 3184 4061
rect 3122 4031 3129 4057
rect 3155 4035 3184 4057
rect 3210 4035 3222 4061
rect 3155 4031 3222 4035
rect 3122 4028 3222 4031
rect 3290 4028 3325 4065
rect 3387 4062 3746 4065
rect 3387 4057 3609 4062
rect 3387 4033 3400 4057
rect 3424 4038 3609 4057
rect 3633 4038 3746 4062
rect 3424 4033 3746 4038
rect 3387 4029 3746 4033
rect 3813 4057 3962 4065
rect 3813 4037 3824 4057
rect 3844 4037 3962 4057
rect 4468 4048 5022 4066
rect 5068 4055 5105 4057
rect 4996 4047 5022 4048
rect 5065 4047 5105 4055
rect 3813 4030 3962 4037
rect 5065 4035 5077 4047
rect 5056 4030 5077 4035
rect 3813 4029 3854 4030
rect 4472 4029 5077 4030
rect 5095 4029 5105 4047
rect 3137 3976 3174 3977
rect 3233 3976 3270 3977
rect 3289 3976 3325 4028
rect 3344 3976 3381 3977
rect 3037 3967 3175 3976
rect 3037 3947 3146 3967
rect 3166 3947 3175 3967
rect 3037 3940 3175 3947
rect 3233 3967 3381 3976
rect 3233 3947 3242 3967
rect 3262 3947 3352 3967
rect 3372 3947 3381 3967
rect 3037 3938 3133 3940
rect 3233 3937 3381 3947
rect 3440 3967 3477 3977
rect 3552 3976 3589 3977
rect 3533 3974 3589 3976
rect 3440 3947 3448 3967
rect 3468 3947 3477 3967
rect 3289 3936 3325 3937
rect 3137 3877 3174 3878
rect 3440 3877 3477 3947
rect 3502 3967 3589 3974
rect 3502 3964 3560 3967
rect 3502 3944 3507 3964
rect 3528 3947 3560 3964
rect 3580 3947 3589 3967
rect 3528 3944 3589 3947
rect 3502 3937 3589 3944
rect 3648 3967 3685 3977
rect 3648 3947 3656 3967
rect 3676 3947 3685 3967
rect 3502 3936 3533 3937
rect 3136 3876 3477 3877
rect 3061 3871 3477 3876
rect 3061 3851 3064 3871
rect 3084 3851 3477 3871
rect 3648 3876 3685 3947
rect 3715 3976 3746 4029
rect 4472 4020 5105 4029
rect 5408 4048 5419 4066
rect 5437 4048 5447 4066
rect 5754 4064 5785 4117
rect 5815 4146 5852 4217
rect 6023 4222 6416 4242
rect 6436 4222 6439 4242
rect 6023 4217 6439 4222
rect 6903 4228 6912 4248
rect 6932 4228 6941 4248
rect 6903 4220 6941 4228
rect 7007 4252 7092 4258
rect 7117 4257 7154 4258
rect 7007 4232 7015 4252
rect 7035 4232 7092 4252
rect 7007 4224 7092 4232
rect 7116 4248 7154 4257
rect 7116 4228 7125 4248
rect 7145 4228 7154 4248
rect 7007 4223 7043 4224
rect 7116 4220 7154 4228
rect 7220 4252 7305 4258
rect 7325 4257 7362 4258
rect 7220 4232 7228 4252
rect 7248 4251 7305 4252
rect 7248 4232 7277 4251
rect 7220 4231 7277 4232
rect 7298 4231 7305 4251
rect 7220 4224 7305 4231
rect 7324 4248 7362 4257
rect 7324 4228 7333 4248
rect 7353 4228 7362 4248
rect 7220 4223 7256 4224
rect 7324 4220 7362 4228
rect 7428 4253 7572 4258
rect 7428 4252 7492 4253
rect 7428 4232 7436 4252
rect 7456 4234 7492 4252
rect 7518 4252 7572 4253
rect 7518 4234 7544 4252
rect 7456 4232 7544 4234
rect 7564 4232 7572 4252
rect 7428 4224 7572 4232
rect 7428 4223 7464 4224
rect 7536 4223 7572 4224
rect 7638 4257 7675 4258
rect 7638 4256 7676 4257
rect 7638 4248 7702 4256
rect 7638 4228 7647 4248
rect 7667 4234 7702 4248
rect 7722 4234 7725 4254
rect 7667 4229 7725 4234
rect 7667 4228 7702 4229
rect 6023 4216 6364 4217
rect 5967 4156 5998 4157
rect 5815 4126 5824 4146
rect 5844 4126 5852 4146
rect 5815 4116 5852 4126
rect 5911 4149 5998 4156
rect 5911 4146 5972 4149
rect 5911 4126 5920 4146
rect 5940 4129 5972 4146
rect 5993 4129 5998 4149
rect 5940 4126 5998 4129
rect 5911 4119 5998 4126
rect 6023 4146 6060 4216
rect 6326 4215 6363 4216
rect 6904 4191 6941 4220
rect 6905 4189 6941 4191
rect 7117 4189 7154 4220
rect 6905 4167 7154 4189
rect 7325 4188 7362 4220
rect 7638 4216 7702 4228
rect 7742 4193 7769 4368
rect 7722 4190 7769 4193
rect 7601 4188 7769 4190
rect 9332 4367 9500 4369
rect 9332 4189 9359 4367
rect 9399 4329 9463 4341
rect 9739 4337 9776 4369
rect 9947 4368 10196 4390
rect 9947 4337 9984 4368
rect 10160 4366 10196 4368
rect 10339 4371 10377 4412
rect 10789 4408 10826 4417
rect 10789 4390 10799 4408
rect 10817 4390 10826 4408
rect 12289 4426 12326 4497
rect 12441 4436 12472 4437
rect 12289 4406 12298 4426
rect 12318 4406 12326 4426
rect 12289 4396 12326 4406
rect 12385 4426 12472 4436
rect 12385 4406 12394 4426
rect 12414 4406 12472 4426
rect 12385 4397 12472 4406
rect 12385 4396 12422 4397
rect 10789 4380 10826 4390
rect 10160 4337 10197 4366
rect 9399 4328 9434 4329
rect 9376 4323 9434 4328
rect 9376 4303 9379 4323
rect 9399 4309 9434 4323
rect 9454 4309 9463 4329
rect 9399 4301 9463 4309
rect 9425 4300 9463 4301
rect 9426 4299 9463 4300
rect 9529 4333 9565 4334
rect 9637 4333 9673 4334
rect 9529 4327 9673 4333
rect 9529 4325 9595 4327
rect 9529 4305 9537 4325
rect 9557 4306 9595 4325
rect 9617 4325 9673 4327
rect 9617 4306 9645 4325
rect 9557 4305 9645 4306
rect 9665 4305 9673 4325
rect 9529 4299 9673 4305
rect 9739 4329 9777 4337
rect 9845 4333 9881 4334
rect 9739 4309 9748 4329
rect 9768 4309 9777 4329
rect 9739 4300 9777 4309
rect 9796 4326 9881 4333
rect 9796 4306 9803 4326
rect 9824 4325 9881 4326
rect 9824 4306 9853 4325
rect 9796 4305 9853 4306
rect 9873 4305 9881 4325
rect 9739 4299 9776 4300
rect 9796 4299 9881 4305
rect 9947 4329 9985 4337
rect 10058 4333 10094 4334
rect 9947 4309 9956 4329
rect 9976 4309 9985 4329
rect 9947 4300 9985 4309
rect 10009 4325 10094 4333
rect 10009 4305 10066 4325
rect 10086 4305 10094 4325
rect 9947 4299 9984 4300
rect 10009 4299 10094 4305
rect 10160 4329 10198 4337
rect 10160 4309 10169 4329
rect 10189 4309 10198 4329
rect 10160 4300 10198 4309
rect 10339 4336 10375 4371
rect 12441 4344 12472 4397
rect 12502 4426 12539 4497
rect 12710 4502 13103 4522
rect 13123 4502 13126 4522
rect 12710 4497 13126 4502
rect 13400 4519 13538 4528
rect 13400 4499 13509 4519
rect 13529 4499 13538 4519
rect 12710 4496 13051 4497
rect 12654 4436 12685 4437
rect 12502 4406 12511 4426
rect 12531 4406 12539 4426
rect 12502 4396 12539 4406
rect 12598 4429 12685 4436
rect 12598 4426 12659 4429
rect 12598 4406 12607 4426
rect 12627 4409 12659 4426
rect 12680 4409 12685 4429
rect 12627 4406 12685 4409
rect 12598 4399 12685 4406
rect 12710 4426 12747 4496
rect 13013 4495 13050 4496
rect 13400 4492 13538 4499
rect 13596 4519 13744 4528
rect 13596 4499 13605 4519
rect 13625 4499 13715 4519
rect 13735 4499 13744 4519
rect 13400 4490 13496 4492
rect 13596 4489 13744 4499
rect 13803 4519 13840 4529
rect 13915 4528 13952 4529
rect 13896 4526 13952 4528
rect 13803 4499 13811 4519
rect 13831 4499 13840 4519
rect 13652 4488 13688 4489
rect 12862 4436 12898 4437
rect 12710 4406 12719 4426
rect 12739 4406 12747 4426
rect 12598 4397 12654 4399
rect 12598 4396 12635 4397
rect 12710 4396 12747 4406
rect 12806 4426 12954 4436
rect 13054 4433 13150 4435
rect 12806 4406 12815 4426
rect 12835 4406 12925 4426
rect 12945 4406 12954 4426
rect 12806 4397 12954 4406
rect 13012 4426 13150 4433
rect 13500 4429 13537 4430
rect 13803 4429 13840 4499
rect 13865 4519 13952 4526
rect 13865 4516 13923 4519
rect 13865 4496 13870 4516
rect 13891 4499 13923 4516
rect 13943 4499 13952 4519
rect 13891 4496 13952 4499
rect 13865 4489 13952 4496
rect 14011 4519 14048 4529
rect 14011 4499 14019 4519
rect 14039 4499 14048 4519
rect 13865 4488 13896 4489
rect 13499 4428 13840 4429
rect 13012 4406 13021 4426
rect 13041 4406 13150 4426
rect 13012 4397 13150 4406
rect 13424 4423 13840 4428
rect 13424 4403 13427 4423
rect 13447 4403 13840 4423
rect 14011 4428 14048 4499
rect 14078 4528 14109 4581
rect 16411 4576 16442 4597
rect 16832 4576 16868 4597
rect 16075 4567 16112 4576
rect 16254 4575 16291 4576
rect 16075 4549 16084 4567
rect 16102 4549 16112 4567
rect 15724 4535 15761 4545
rect 16075 4539 16112 4549
rect 14128 4528 14165 4529
rect 14078 4519 14165 4528
rect 14078 4499 14136 4519
rect 14156 4499 14165 4519
rect 14078 4489 14165 4499
rect 14224 4519 14261 4529
rect 14224 4499 14232 4519
rect 14252 4499 14261 4519
rect 14078 4488 14109 4489
rect 14224 4428 14261 4499
rect 15724 4517 15733 4535
rect 15751 4517 15761 4535
rect 15724 4508 15761 4517
rect 15724 4465 15759 4508
rect 16076 4504 16112 4539
rect 16253 4566 16291 4575
rect 16253 4546 16262 4566
rect 16282 4546 16291 4566
rect 16253 4538 16291 4546
rect 16357 4570 16442 4576
rect 16467 4575 16504 4576
rect 16357 4550 16365 4570
rect 16385 4550 16442 4570
rect 16357 4542 16442 4550
rect 16466 4566 16504 4575
rect 16466 4546 16475 4566
rect 16495 4546 16504 4566
rect 16357 4541 16393 4542
rect 16466 4538 16504 4546
rect 16570 4570 16655 4576
rect 16675 4575 16712 4576
rect 16570 4550 16578 4570
rect 16598 4569 16655 4570
rect 16598 4550 16627 4569
rect 16570 4549 16627 4550
rect 16648 4549 16655 4569
rect 16570 4542 16655 4549
rect 16674 4566 16712 4575
rect 16674 4546 16683 4566
rect 16703 4546 16712 4566
rect 16570 4541 16606 4542
rect 16674 4538 16712 4546
rect 16778 4570 16922 4576
rect 16778 4550 16786 4570
rect 16806 4569 16894 4570
rect 16806 4550 16834 4569
rect 16778 4548 16834 4550
rect 16856 4550 16894 4569
rect 16914 4550 16922 4570
rect 16856 4548 16922 4550
rect 16778 4542 16922 4548
rect 16778 4541 16814 4542
rect 16886 4541 16922 4542
rect 16988 4575 17025 4576
rect 16988 4574 17026 4575
rect 16988 4566 17052 4574
rect 16988 4546 16997 4566
rect 17017 4552 17052 4566
rect 17072 4552 17075 4572
rect 17017 4547 17075 4552
rect 17017 4546 17052 4547
rect 16254 4509 16291 4538
rect 15719 4460 15759 4465
rect 16074 4463 16112 4504
rect 16255 4507 16291 4509
rect 16467 4507 16504 4538
rect 16255 4485 16504 4507
rect 16675 4506 16712 4538
rect 16988 4534 17052 4546
rect 17092 4508 17119 4686
rect 16951 4506 17119 4508
rect 18682 4685 18850 4687
rect 18682 4682 18729 4685
rect 18682 4507 18709 4682
rect 18749 4647 18813 4659
rect 19089 4655 19126 4687
rect 19297 4686 19546 4708
rect 19297 4655 19334 4686
rect 19510 4684 19546 4686
rect 19510 4655 19547 4684
rect 20088 4659 20125 4660
rect 20391 4659 20428 4729
rect 20453 4749 20540 4756
rect 20453 4746 20511 4749
rect 20453 4726 20458 4746
rect 20479 4729 20511 4746
rect 20531 4729 20540 4749
rect 20479 4726 20540 4729
rect 20453 4719 20540 4726
rect 20599 4749 20636 4759
rect 20599 4729 20607 4749
rect 20627 4729 20636 4749
rect 20453 4718 20484 4719
rect 20087 4658 20428 4659
rect 18749 4646 18784 4647
rect 18726 4641 18784 4646
rect 18726 4621 18729 4641
rect 18749 4627 18784 4641
rect 18804 4627 18813 4647
rect 18749 4619 18813 4627
rect 18775 4618 18813 4619
rect 18776 4617 18813 4618
rect 18879 4651 18915 4652
rect 18987 4651 19023 4652
rect 18879 4643 19023 4651
rect 18879 4623 18887 4643
rect 18907 4641 18995 4643
rect 18907 4623 18933 4641
rect 18879 4622 18933 4623
rect 18959 4623 18995 4641
rect 19015 4623 19023 4643
rect 18959 4622 19023 4623
rect 18879 4617 19023 4622
rect 19089 4647 19127 4655
rect 19195 4651 19231 4652
rect 19089 4627 19098 4647
rect 19118 4627 19127 4647
rect 19089 4618 19127 4627
rect 19146 4644 19231 4651
rect 19146 4624 19153 4644
rect 19174 4643 19231 4644
rect 19174 4624 19203 4643
rect 19146 4623 19203 4624
rect 19223 4623 19231 4643
rect 19089 4617 19126 4618
rect 19146 4617 19231 4623
rect 19297 4647 19335 4655
rect 19408 4651 19444 4652
rect 19297 4627 19306 4647
rect 19326 4627 19335 4647
rect 19297 4618 19335 4627
rect 19359 4643 19444 4651
rect 19359 4623 19416 4643
rect 19436 4623 19444 4643
rect 19297 4617 19334 4618
rect 19359 4617 19444 4623
rect 19510 4647 19548 4655
rect 19510 4627 19519 4647
rect 19539 4627 19548 4647
rect 20012 4653 20428 4658
rect 20012 4633 20015 4653
rect 20035 4633 20428 4653
rect 20599 4658 20636 4729
rect 20666 4758 20697 4811
rect 21004 4809 21014 4827
rect 21032 4809 21043 4827
rect 21004 4800 21041 4809
rect 20716 4758 20753 4759
rect 20666 4749 20753 4758
rect 20666 4729 20724 4749
rect 20744 4729 20753 4749
rect 20666 4719 20753 4729
rect 20812 4749 20849 4759
rect 20812 4729 20820 4749
rect 20840 4729 20849 4749
rect 21007 4734 21044 4738
rect 20666 4718 20697 4719
rect 20812 4658 20849 4729
rect 20599 4634 20849 4658
rect 21005 4728 21044 4734
rect 21005 4710 21016 4728
rect 21034 4710 21044 4728
rect 21005 4701 21044 4710
rect 19510 4618 19548 4627
rect 19510 4617 19547 4618
rect 18933 4596 18969 4617
rect 19359 4596 19390 4617
rect 20391 4610 20428 4633
rect 21005 4623 21040 4701
rect 21002 4613 21040 4623
rect 20391 4609 20561 4610
rect 21002 4609 21012 4613
rect 18766 4592 18866 4596
rect 18766 4588 18828 4592
rect 18766 4562 18773 4588
rect 18799 4566 18828 4588
rect 18854 4566 18866 4592
rect 18799 4562 18866 4566
rect 18766 4559 18866 4562
rect 18934 4559 18969 4596
rect 19031 4593 19390 4596
rect 19031 4588 19253 4593
rect 19031 4564 19044 4588
rect 19068 4569 19253 4588
rect 19277 4569 19390 4593
rect 19068 4564 19390 4569
rect 19031 4560 19390 4564
rect 19457 4588 19606 4596
rect 20391 4595 21012 4609
rect 21030 4595 21040 4613
rect 20391 4589 21040 4595
rect 20391 4588 21039 4589
rect 19457 4568 19468 4588
rect 19488 4568 19606 4588
rect 21002 4586 21039 4588
rect 19457 4561 19606 4568
rect 19457 4560 19498 4561
rect 18781 4507 18818 4508
rect 18877 4507 18914 4508
rect 18933 4507 18969 4559
rect 18988 4507 19025 4508
rect 16675 4480 17119 4506
rect 16676 4463 16700 4480
rect 16951 4479 17119 4480
rect 17570 4476 17820 4500
rect 15719 4459 15757 4460
rect 15130 4441 15757 4459
rect 16074 4445 16701 4463
rect 16074 4444 16112 4445
rect 14011 4404 14261 4428
rect 14712 4424 14880 4425
rect 15131 4424 15155 4441
rect 14712 4398 15156 4424
rect 12806 4396 12843 4397
rect 12862 4345 12898 4397
rect 12917 4396 12954 4397
rect 13013 4396 13050 4397
rect 12333 4343 12374 4344
rect 12225 4336 12374 4343
rect 10339 4326 10376 4336
rect 10339 4308 10349 4326
rect 10367 4308 10376 4326
rect 10792 4316 10829 4318
rect 12225 4316 12343 4336
rect 12363 4316 12374 4336
rect 10792 4315 11440 4316
rect 10160 4299 10197 4300
rect 10339 4299 10376 4308
rect 10791 4309 11440 4315
rect 9583 4278 9619 4299
rect 10009 4278 10040 4299
rect 10791 4291 10801 4309
rect 10819 4295 11440 4309
rect 12225 4308 12374 4316
rect 12441 4340 12800 4344
rect 12441 4335 12763 4340
rect 12441 4311 12554 4335
rect 12578 4316 12763 4335
rect 12787 4316 12800 4340
rect 12578 4311 12800 4316
rect 12441 4308 12800 4311
rect 12862 4308 12897 4345
rect 12965 4342 13065 4345
rect 12965 4338 13032 4342
rect 12965 4312 12977 4338
rect 13003 4316 13032 4338
rect 13058 4316 13065 4342
rect 13003 4312 13065 4316
rect 12965 4308 13065 4312
rect 10819 4291 10829 4295
rect 11270 4294 11440 4295
rect 10791 4281 10829 4291
rect 9416 4274 9516 4278
rect 9416 4270 9478 4274
rect 9416 4244 9423 4270
rect 9449 4248 9478 4270
rect 9504 4248 9516 4274
rect 9449 4244 9516 4248
rect 9416 4241 9516 4244
rect 9584 4241 9619 4278
rect 9681 4275 10040 4278
rect 9681 4270 9903 4275
rect 9681 4246 9694 4270
rect 9718 4251 9903 4270
rect 9927 4251 10040 4275
rect 9718 4246 10040 4251
rect 9681 4242 10040 4246
rect 10107 4270 10256 4278
rect 10107 4250 10118 4270
rect 10138 4250 10256 4270
rect 10107 4243 10256 4250
rect 10107 4242 10148 4243
rect 9431 4189 9468 4190
rect 9527 4189 9564 4190
rect 9583 4189 9619 4241
rect 9638 4189 9675 4190
rect 7325 4162 7769 4188
rect 9331 4180 9469 4189
rect 7601 4161 7769 4162
rect 8267 4162 8298 4165
rect 6175 4156 6211 4157
rect 6023 4126 6032 4146
rect 6052 4126 6060 4146
rect 5911 4117 5967 4119
rect 5911 4116 5948 4117
rect 6023 4116 6060 4126
rect 6119 4146 6267 4156
rect 6367 4153 6463 4155
rect 6119 4126 6128 4146
rect 6148 4126 6238 4146
rect 6258 4126 6267 4146
rect 6119 4117 6267 4126
rect 6325 4146 6463 4153
rect 6325 4126 6334 4146
rect 6354 4126 6463 4146
rect 6325 4117 6463 4126
rect 6119 4116 6156 4117
rect 6175 4065 6211 4117
rect 6230 4116 6267 4117
rect 6326 4116 6363 4117
rect 5646 4063 5687 4064
rect 4472 4013 5104 4020
rect 4472 4011 4534 4013
rect 4050 4001 4218 4002
rect 4472 4001 4494 4011
rect 3765 3976 3802 3977
rect 3715 3967 3802 3976
rect 3715 3947 3773 3967
rect 3793 3947 3802 3967
rect 3715 3937 3802 3947
rect 3861 3967 3898 3977
rect 3861 3947 3869 3967
rect 3889 3947 3898 3967
rect 3715 3936 3746 3937
rect 3861 3876 3898 3947
rect 3648 3852 3898 3876
rect 4050 3975 4494 4001
rect 4050 3973 4218 3975
rect 4050 3795 4077 3973
rect 4117 3935 4181 3947
rect 4457 3943 4494 3975
rect 4665 3974 4914 3996
rect 4665 3943 4702 3974
rect 4878 3972 4914 3974
rect 4878 3943 4915 3972
rect 4117 3934 4152 3935
rect 4094 3929 4152 3934
rect 4094 3909 4097 3929
rect 4117 3915 4152 3929
rect 4172 3915 4181 3935
rect 4117 3907 4181 3915
rect 4143 3906 4181 3907
rect 4144 3905 4181 3906
rect 4247 3939 4283 3940
rect 4355 3939 4391 3940
rect 4247 3931 4391 3939
rect 4247 3911 4255 3931
rect 4275 3911 4304 3931
rect 4247 3910 4304 3911
rect 4326 3911 4363 3931
rect 4383 3911 4391 3931
rect 4326 3910 4391 3911
rect 4247 3905 4391 3910
rect 4457 3935 4495 3943
rect 4563 3939 4599 3940
rect 4457 3915 4466 3935
rect 4486 3915 4495 3935
rect 4457 3906 4495 3915
rect 4514 3932 4599 3939
rect 4514 3912 4521 3932
rect 4542 3931 4599 3932
rect 4542 3912 4571 3931
rect 4514 3911 4571 3912
rect 4591 3911 4599 3931
rect 4457 3905 4494 3906
rect 4514 3905 4599 3911
rect 4665 3935 4703 3943
rect 4776 3939 4812 3940
rect 4665 3915 4674 3935
rect 4694 3915 4703 3935
rect 4665 3906 4703 3915
rect 4727 3931 4812 3939
rect 4727 3911 4784 3931
rect 4804 3911 4812 3931
rect 4665 3905 4702 3906
rect 4727 3905 4812 3911
rect 4878 3935 4916 3943
rect 4878 3915 4887 3935
rect 4907 3915 4916 3935
rect 4878 3906 4916 3915
rect 4878 3905 4915 3906
rect 4301 3884 4337 3905
rect 4727 3884 4758 3905
rect 4134 3880 4234 3884
rect 4134 3876 4196 3880
rect 4134 3850 4141 3876
rect 4167 3854 4196 3876
rect 4222 3854 4234 3880
rect 4167 3850 4234 3854
rect 4134 3847 4234 3850
rect 4302 3847 4337 3884
rect 4399 3881 4758 3884
rect 4399 3876 4621 3881
rect 4399 3852 4412 3876
rect 4436 3857 4621 3876
rect 4645 3857 4758 3881
rect 4436 3852 4758 3857
rect 4399 3848 4758 3852
rect 4825 3876 4974 3884
rect 4825 3856 4836 3876
rect 4856 3856 4974 3876
rect 4825 3849 4974 3856
rect 5065 3864 5104 4013
rect 5408 3899 5447 4048
rect 5538 4056 5687 4063
rect 5538 4036 5656 4056
rect 5676 4036 5687 4056
rect 5538 4028 5687 4036
rect 5754 4060 6113 4064
rect 5754 4055 6076 4060
rect 5754 4031 5867 4055
rect 5891 4036 6076 4055
rect 6100 4036 6113 4060
rect 5891 4031 6113 4036
rect 5754 4028 6113 4031
rect 6175 4028 6210 4065
rect 6278 4062 6378 4065
rect 6278 4058 6345 4062
rect 6278 4032 6290 4058
rect 6316 4036 6345 4058
rect 6371 4036 6378 4062
rect 6316 4032 6378 4036
rect 6278 4028 6378 4032
rect 5754 4007 5785 4028
rect 6175 4007 6211 4028
rect 5597 4006 5634 4007
rect 5596 3997 5634 4006
rect 5596 3977 5605 3997
rect 5625 3977 5634 3997
rect 5596 3969 5634 3977
rect 5700 4001 5785 4007
rect 5810 4006 5847 4007
rect 5700 3981 5708 4001
rect 5728 3981 5785 4001
rect 5700 3973 5785 3981
rect 5809 3997 5847 4006
rect 5809 3977 5818 3997
rect 5838 3977 5847 3997
rect 5700 3972 5736 3973
rect 5809 3969 5847 3977
rect 5913 4001 5998 4007
rect 6018 4006 6055 4007
rect 5913 3981 5921 4001
rect 5941 4000 5998 4001
rect 5941 3981 5970 4000
rect 5913 3980 5970 3981
rect 5991 3980 5998 4000
rect 5913 3973 5998 3980
rect 6017 3997 6055 4006
rect 6017 3977 6026 3997
rect 6046 3977 6055 3997
rect 5913 3972 5949 3973
rect 6017 3969 6055 3977
rect 6121 4002 6265 4007
rect 6121 4001 6186 4002
rect 6121 3981 6129 4001
rect 6149 3981 6186 4001
rect 6208 4001 6265 4002
rect 6208 3981 6237 4001
rect 6257 3981 6265 4001
rect 6121 3973 6265 3981
rect 6121 3972 6157 3973
rect 6229 3972 6265 3973
rect 6331 4006 6368 4007
rect 6331 4005 6369 4006
rect 6331 3997 6395 4005
rect 6331 3977 6340 3997
rect 6360 3983 6395 3997
rect 6415 3983 6418 4003
rect 6360 3978 6418 3983
rect 6360 3977 6395 3978
rect 5597 3940 5634 3969
rect 5598 3938 5634 3940
rect 5810 3938 5847 3969
rect 5598 3916 5847 3938
rect 6018 3937 6055 3969
rect 6331 3965 6395 3977
rect 6435 3939 6462 4117
rect 6294 3937 6462 3939
rect 6018 3911 6462 3937
rect 6614 4036 6864 4060
rect 6614 3965 6651 4036
rect 6766 3975 6797 3976
rect 6614 3945 6623 3965
rect 6643 3945 6651 3965
rect 6614 3935 6651 3945
rect 6710 3965 6797 3975
rect 6710 3945 6719 3965
rect 6739 3945 6797 3965
rect 6710 3936 6797 3945
rect 6710 3935 6747 3936
rect 6018 3901 6040 3911
rect 6294 3910 6462 3911
rect 5978 3899 6040 3901
rect 5408 3892 6040 3899
rect 4825 3848 4866 3849
rect 4149 3795 4186 3796
rect 4245 3795 4282 3796
rect 4301 3795 4337 3847
rect 4356 3795 4393 3796
rect 4049 3786 4187 3795
rect 4049 3766 4158 3786
rect 4178 3766 4187 3786
rect 2986 3762 3156 3763
rect 2986 3747 3432 3762
rect 4049 3759 4187 3766
rect 4245 3786 4393 3795
rect 4245 3766 4254 3786
rect 4274 3766 4364 3786
rect 4384 3766 4393 3786
rect 4049 3757 4145 3759
rect 2893 3736 2925 3741
rect 2895 2735 2925 3736
rect 2988 3736 3432 3747
rect 2988 3734 3156 3736
rect 2988 3556 3015 3734
rect 3055 3696 3119 3708
rect 3395 3704 3432 3736
rect 3603 3735 3852 3757
rect 4245 3756 4393 3766
rect 4452 3786 4489 3796
rect 4564 3795 4601 3796
rect 4545 3793 4601 3795
rect 4452 3766 4460 3786
rect 4480 3766 4489 3786
rect 4301 3755 4337 3756
rect 3603 3704 3640 3735
rect 3816 3733 3852 3735
rect 3816 3704 3853 3733
rect 3055 3695 3090 3696
rect 3032 3690 3090 3695
rect 3032 3670 3035 3690
rect 3055 3676 3090 3690
rect 3110 3676 3119 3696
rect 3055 3668 3119 3676
rect 3081 3667 3119 3668
rect 3082 3666 3119 3667
rect 3185 3700 3221 3701
rect 3293 3700 3329 3701
rect 3185 3692 3329 3700
rect 3185 3672 3193 3692
rect 3213 3673 3245 3692
rect 3268 3673 3301 3692
rect 3213 3672 3301 3673
rect 3321 3672 3329 3692
rect 3185 3666 3329 3672
rect 3395 3696 3433 3704
rect 3501 3700 3537 3701
rect 3395 3676 3404 3696
rect 3424 3676 3433 3696
rect 3395 3667 3433 3676
rect 3452 3693 3537 3700
rect 3452 3673 3459 3693
rect 3480 3692 3537 3693
rect 3480 3673 3509 3692
rect 3452 3672 3509 3673
rect 3529 3672 3537 3692
rect 3395 3666 3432 3667
rect 3452 3666 3537 3672
rect 3603 3696 3641 3704
rect 3714 3700 3750 3701
rect 3603 3676 3612 3696
rect 3632 3676 3641 3696
rect 3603 3667 3641 3676
rect 3665 3692 3750 3700
rect 3665 3672 3722 3692
rect 3742 3672 3750 3692
rect 3603 3666 3640 3667
rect 3665 3666 3750 3672
rect 3816 3696 3854 3704
rect 4149 3696 4186 3697
rect 4452 3696 4489 3766
rect 4514 3786 4601 3793
rect 4514 3783 4572 3786
rect 4514 3763 4519 3783
rect 4540 3766 4572 3783
rect 4592 3766 4601 3786
rect 4540 3763 4601 3766
rect 4514 3756 4601 3763
rect 4660 3786 4697 3796
rect 4660 3766 4668 3786
rect 4688 3766 4697 3786
rect 4514 3755 4545 3756
rect 3816 3676 3825 3696
rect 3845 3676 3854 3696
rect 4148 3695 4489 3696
rect 3816 3667 3854 3676
rect 4073 3690 4489 3695
rect 4073 3670 4076 3690
rect 4096 3670 4489 3690
rect 4660 3695 4697 3766
rect 4727 3795 4758 3848
rect 5065 3846 5075 3864
rect 5093 3846 5104 3864
rect 5407 3883 6040 3892
rect 6766 3883 6797 3936
rect 6827 3965 6864 4036
rect 7035 4041 7428 4061
rect 7448 4041 7451 4061
rect 7035 4036 7451 4041
rect 7035 4035 7376 4036
rect 6979 3975 7010 3976
rect 6827 3945 6836 3965
rect 6856 3945 6864 3965
rect 6827 3935 6864 3945
rect 6923 3968 7010 3975
rect 6923 3965 6984 3968
rect 6923 3945 6932 3965
rect 6952 3948 6984 3965
rect 7005 3948 7010 3968
rect 6952 3945 7010 3948
rect 6923 3938 7010 3945
rect 7035 3965 7072 4035
rect 7338 4034 7375 4035
rect 7187 3975 7223 3976
rect 7035 3945 7044 3965
rect 7064 3945 7072 3965
rect 6923 3936 6979 3938
rect 6923 3935 6960 3936
rect 7035 3935 7072 3945
rect 7131 3965 7279 3975
rect 7379 3972 7475 3974
rect 7131 3945 7140 3965
rect 7160 3945 7250 3965
rect 7270 3945 7279 3965
rect 7131 3936 7279 3945
rect 7337 3965 7475 3972
rect 7337 3945 7346 3965
rect 7366 3945 7475 3965
rect 7337 3936 7475 3945
rect 7131 3935 7168 3936
rect 7187 3884 7223 3936
rect 7242 3935 7279 3936
rect 7338 3935 7375 3936
rect 5407 3865 5417 3883
rect 5435 3882 6040 3883
rect 6658 3882 6699 3883
rect 5435 3877 5456 3882
rect 5435 3865 5447 3877
rect 6550 3875 6699 3882
rect 5407 3857 5447 3865
rect 5490 3864 5516 3865
rect 5407 3855 5444 3857
rect 5490 3846 6044 3864
rect 6550 3855 6668 3875
rect 6688 3855 6699 3875
rect 6550 3847 6699 3855
rect 6766 3879 7125 3883
rect 6766 3874 7088 3879
rect 6766 3850 6879 3874
rect 6903 3855 7088 3874
rect 7112 3855 7125 3879
rect 6903 3850 7125 3855
rect 6766 3847 7125 3850
rect 7187 3847 7222 3884
rect 7290 3881 7390 3884
rect 7290 3877 7357 3881
rect 7290 3851 7302 3877
rect 7328 3855 7357 3877
rect 7383 3855 7390 3881
rect 7328 3851 7390 3855
rect 7290 3847 7390 3851
rect 5065 3837 5102 3846
rect 4777 3795 4814 3796
rect 4727 3786 4814 3795
rect 4727 3766 4785 3786
rect 4805 3766 4814 3786
rect 4727 3756 4814 3766
rect 4873 3786 4910 3796
rect 4873 3766 4881 3786
rect 4901 3766 4910 3786
rect 5410 3787 5447 3793
rect 5490 3787 5516 3846
rect 6023 3827 6044 3846
rect 5410 3784 5516 3787
rect 5068 3771 5105 3775
rect 4727 3755 4758 3756
rect 4873 3695 4910 3766
rect 4660 3671 4910 3695
rect 5066 3765 5105 3771
rect 5066 3747 5077 3765
rect 5095 3747 5105 3765
rect 5410 3766 5419 3784
rect 5437 3770 5516 3784
rect 5601 3802 5851 3826
rect 5437 3768 5513 3770
rect 5437 3766 5447 3768
rect 5410 3756 5447 3766
rect 5066 3738 5105 3747
rect 3816 3666 3853 3667
rect 3239 3645 3275 3666
rect 3665 3645 3696 3666
rect 4452 3647 4489 3670
rect 5066 3660 5101 3738
rect 5415 3691 5446 3756
rect 5601 3731 5638 3802
rect 5753 3741 5784 3742
rect 5601 3711 5610 3731
rect 5630 3711 5638 3731
rect 5601 3701 5638 3711
rect 5697 3731 5784 3741
rect 5697 3711 5706 3731
rect 5726 3711 5784 3731
rect 5697 3702 5784 3711
rect 5697 3701 5734 3702
rect 5063 3650 5101 3660
rect 5414 3682 5451 3691
rect 5414 3664 5424 3682
rect 5442 3664 5451 3682
rect 5414 3654 5451 3664
rect 4452 3646 4622 3647
rect 5063 3646 5073 3650
rect 3072 3641 3172 3645
rect 3072 3637 3134 3641
rect 3072 3611 3079 3637
rect 3105 3615 3134 3637
rect 3160 3615 3172 3641
rect 3105 3611 3172 3615
rect 3072 3608 3172 3611
rect 3240 3608 3275 3645
rect 3337 3642 3696 3645
rect 3337 3637 3559 3642
rect 3337 3613 3350 3637
rect 3374 3618 3559 3637
rect 3583 3618 3696 3642
rect 3374 3613 3696 3618
rect 3337 3609 3696 3613
rect 3763 3637 3912 3645
rect 3763 3617 3774 3637
rect 3794 3617 3912 3637
rect 4452 3632 5073 3646
rect 5091 3632 5101 3650
rect 5753 3649 5784 3702
rect 5814 3731 5851 3802
rect 6022 3807 6415 3827
rect 6435 3807 6438 3827
rect 6766 3826 6797 3847
rect 7187 3826 7223 3847
rect 6609 3825 6646 3826
rect 6022 3802 6438 3807
rect 6608 3816 6646 3825
rect 6022 3801 6363 3802
rect 5966 3741 5997 3742
rect 5814 3711 5823 3731
rect 5843 3711 5851 3731
rect 5814 3701 5851 3711
rect 5910 3734 5997 3741
rect 5910 3731 5971 3734
rect 5910 3711 5919 3731
rect 5939 3714 5971 3731
rect 5992 3714 5997 3734
rect 5939 3711 5997 3714
rect 5910 3704 5997 3711
rect 6022 3731 6059 3801
rect 6325 3800 6362 3801
rect 6608 3796 6617 3816
rect 6637 3796 6646 3816
rect 6608 3788 6646 3796
rect 6712 3820 6797 3826
rect 6822 3825 6859 3826
rect 6712 3800 6720 3820
rect 6740 3800 6797 3820
rect 6712 3792 6797 3800
rect 6821 3816 6859 3825
rect 6821 3796 6830 3816
rect 6850 3796 6859 3816
rect 6712 3791 6748 3792
rect 6821 3788 6859 3796
rect 6925 3820 7010 3826
rect 7030 3825 7067 3826
rect 6925 3800 6933 3820
rect 6953 3819 7010 3820
rect 6953 3800 6982 3819
rect 6925 3799 6982 3800
rect 7003 3799 7010 3819
rect 6925 3792 7010 3799
rect 7029 3816 7067 3825
rect 7029 3796 7038 3816
rect 7058 3796 7067 3816
rect 6925 3791 6961 3792
rect 7029 3788 7067 3796
rect 7133 3820 7277 3826
rect 7133 3800 7141 3820
rect 7161 3800 7193 3820
rect 7217 3800 7249 3820
rect 7269 3800 7277 3820
rect 7133 3792 7277 3800
rect 7133 3791 7169 3792
rect 7241 3791 7277 3792
rect 7343 3825 7380 3826
rect 7343 3824 7381 3825
rect 7343 3816 7407 3824
rect 7343 3796 7352 3816
rect 7372 3802 7407 3816
rect 7427 3802 7430 3822
rect 7372 3797 7430 3802
rect 7372 3796 7407 3797
rect 6609 3759 6646 3788
rect 6610 3757 6646 3759
rect 6822 3757 6859 3788
rect 6174 3741 6210 3742
rect 6022 3711 6031 3731
rect 6051 3711 6059 3731
rect 5910 3702 5966 3704
rect 5910 3701 5947 3702
rect 6022 3701 6059 3711
rect 6118 3731 6266 3741
rect 6366 3738 6462 3740
rect 6118 3711 6127 3731
rect 6147 3711 6237 3731
rect 6257 3711 6266 3731
rect 6118 3702 6266 3711
rect 6324 3731 6462 3738
rect 6610 3735 6859 3757
rect 7030 3756 7067 3788
rect 7343 3784 7407 3796
rect 7447 3758 7474 3936
rect 7306 3756 7474 3758
rect 7030 3752 7474 3756
rect 6324 3711 6333 3731
rect 6353 3711 6462 3731
rect 7030 3733 7079 3752
rect 7099 3733 7474 3752
rect 7030 3730 7474 3733
rect 7306 3729 7474 3730
rect 6324 3702 6462 3711
rect 6118 3701 6155 3702
rect 6174 3650 6210 3702
rect 6229 3701 6266 3702
rect 6325 3701 6362 3702
rect 5645 3648 5686 3649
rect 4452 3626 5101 3632
rect 5537 3641 5686 3648
rect 4452 3625 5100 3626
rect 5063 3623 5100 3625
rect 3763 3610 3912 3617
rect 5537 3621 5655 3641
rect 5675 3621 5686 3641
rect 5537 3613 5686 3621
rect 5753 3645 6112 3649
rect 5753 3640 6075 3645
rect 5753 3616 5866 3640
rect 5890 3621 6075 3640
rect 6099 3621 6112 3645
rect 5890 3616 6112 3621
rect 5753 3613 6112 3616
rect 6174 3613 6209 3650
rect 6277 3647 6377 3650
rect 6277 3643 6344 3647
rect 6277 3617 6289 3643
rect 6315 3621 6344 3643
rect 6370 3621 6377 3647
rect 6315 3617 6377 3621
rect 6277 3613 6377 3617
rect 3763 3609 3804 3610
rect 3087 3556 3124 3557
rect 3183 3556 3220 3557
rect 3239 3556 3275 3608
rect 3294 3556 3331 3557
rect 2987 3547 3125 3556
rect 2987 3527 3096 3547
rect 3116 3527 3125 3547
rect 2987 3520 3125 3527
rect 3183 3547 3331 3556
rect 3183 3527 3192 3547
rect 3212 3527 3302 3547
rect 3322 3527 3331 3547
rect 2987 3518 3083 3520
rect 3183 3517 3331 3527
rect 3390 3547 3427 3557
rect 3502 3556 3539 3557
rect 3483 3554 3539 3556
rect 3390 3527 3398 3547
rect 3418 3527 3427 3547
rect 3239 3516 3275 3517
rect 3087 3457 3124 3458
rect 3390 3457 3427 3527
rect 3452 3547 3539 3554
rect 3452 3544 3510 3547
rect 3452 3524 3457 3544
rect 3478 3527 3510 3544
rect 3530 3527 3539 3547
rect 3478 3524 3539 3527
rect 3452 3517 3539 3524
rect 3598 3547 3635 3557
rect 3598 3527 3606 3547
rect 3626 3527 3635 3547
rect 3452 3516 3483 3517
rect 3086 3456 3427 3457
rect 3011 3451 3427 3456
rect 3011 3431 3014 3451
rect 3034 3431 3427 3451
rect 3598 3456 3635 3527
rect 3665 3556 3696 3609
rect 5753 3592 5784 3613
rect 6174 3592 6210 3613
rect 5417 3583 5454 3592
rect 5596 3591 5633 3592
rect 5417 3565 5426 3583
rect 5444 3565 5454 3583
rect 3715 3556 3752 3557
rect 3665 3547 3752 3556
rect 3665 3527 3723 3547
rect 3743 3527 3752 3547
rect 3665 3517 3752 3527
rect 3811 3547 3848 3557
rect 3811 3527 3819 3547
rect 3839 3527 3848 3547
rect 3665 3516 3696 3517
rect 3811 3456 3848 3527
rect 5066 3551 5103 3561
rect 5417 3555 5454 3565
rect 5066 3533 5075 3551
rect 5093 3533 5103 3551
rect 5066 3524 5103 3533
rect 5066 3500 5101 3524
rect 5418 3520 5454 3555
rect 5595 3582 5633 3591
rect 5595 3562 5604 3582
rect 5624 3562 5633 3582
rect 5595 3554 5633 3562
rect 5699 3586 5784 3592
rect 5809 3591 5846 3592
rect 5699 3566 5707 3586
rect 5727 3566 5784 3586
rect 5699 3558 5784 3566
rect 5808 3582 5846 3591
rect 5808 3562 5817 3582
rect 5837 3562 5846 3582
rect 5699 3557 5735 3558
rect 5808 3554 5846 3562
rect 5912 3586 5997 3592
rect 6017 3591 6054 3592
rect 5912 3566 5920 3586
rect 5940 3585 5997 3586
rect 5940 3566 5969 3585
rect 5912 3565 5969 3566
rect 5990 3565 5997 3585
rect 5912 3558 5997 3565
rect 6016 3582 6054 3591
rect 6016 3562 6025 3582
rect 6045 3562 6054 3582
rect 5912 3557 5948 3558
rect 6016 3554 6054 3562
rect 6120 3586 6264 3592
rect 6120 3566 6128 3586
rect 6148 3585 6236 3586
rect 6148 3566 6176 3585
rect 6120 3564 6176 3566
rect 6198 3566 6236 3585
rect 6256 3566 6264 3586
rect 6198 3564 6264 3566
rect 6120 3558 6264 3564
rect 6120 3557 6156 3558
rect 6228 3557 6264 3558
rect 6330 3591 6367 3592
rect 6330 3590 6368 3591
rect 6330 3582 6394 3590
rect 6330 3562 6339 3582
rect 6359 3568 6394 3582
rect 6414 3568 6417 3588
rect 6359 3563 6417 3568
rect 6359 3562 6394 3563
rect 5596 3525 5633 3554
rect 5064 3476 5101 3500
rect 5063 3470 5101 3476
rect 3598 3432 3848 3456
rect 4474 3452 5101 3470
rect 4056 3435 4224 3436
rect 4475 3435 4499 3452
rect 4056 3409 4500 3435
rect 4056 3407 4224 3409
rect 4056 3229 4083 3407
rect 4123 3369 4187 3381
rect 4463 3377 4500 3409
rect 4671 3408 4920 3430
rect 4671 3377 4708 3408
rect 4884 3406 4920 3408
rect 5063 3411 5101 3452
rect 5416 3479 5454 3520
rect 5597 3523 5633 3525
rect 5809 3523 5846 3554
rect 5597 3501 5846 3523
rect 6017 3522 6054 3554
rect 6330 3550 6394 3562
rect 6434 3524 6461 3702
rect 6293 3522 6461 3524
rect 6017 3496 6461 3522
rect 6018 3479 6042 3496
rect 6293 3495 6461 3496
rect 5416 3461 6043 3479
rect 6669 3475 6919 3499
rect 5416 3455 5454 3461
rect 5416 3431 5453 3455
rect 4884 3377 4921 3406
rect 4123 3368 4158 3369
rect 4100 3363 4158 3368
rect 4100 3343 4103 3363
rect 4123 3349 4158 3363
rect 4178 3349 4187 3369
rect 4123 3341 4187 3349
rect 4149 3340 4187 3341
rect 4150 3339 4187 3340
rect 4253 3373 4289 3374
rect 4361 3373 4397 3374
rect 4253 3367 4397 3373
rect 4253 3365 4319 3367
rect 4253 3345 4261 3365
rect 4281 3346 4319 3365
rect 4341 3365 4397 3367
rect 4341 3346 4369 3365
rect 4281 3345 4369 3346
rect 4389 3345 4397 3365
rect 4253 3339 4397 3345
rect 4463 3369 4501 3377
rect 4569 3373 4605 3374
rect 4463 3349 4472 3369
rect 4492 3349 4501 3369
rect 4463 3340 4501 3349
rect 4520 3366 4605 3373
rect 4520 3346 4527 3366
rect 4548 3365 4605 3366
rect 4548 3346 4577 3365
rect 4520 3345 4577 3346
rect 4597 3345 4605 3365
rect 4463 3339 4500 3340
rect 4520 3339 4605 3345
rect 4671 3369 4709 3377
rect 4782 3373 4818 3374
rect 4671 3349 4680 3369
rect 4700 3349 4709 3369
rect 4671 3340 4709 3349
rect 4733 3365 4818 3373
rect 4733 3345 4790 3365
rect 4810 3345 4818 3365
rect 4671 3339 4708 3340
rect 4733 3339 4818 3345
rect 4884 3369 4922 3377
rect 4884 3349 4893 3369
rect 4913 3349 4922 3369
rect 4884 3340 4922 3349
rect 5063 3376 5099 3411
rect 5416 3407 5451 3431
rect 5414 3398 5451 3407
rect 5414 3380 5424 3398
rect 5442 3380 5451 3398
rect 5063 3366 5100 3376
rect 5414 3370 5451 3380
rect 6669 3404 6706 3475
rect 6821 3414 6852 3415
rect 6669 3384 6678 3404
rect 6698 3384 6706 3404
rect 6669 3374 6706 3384
rect 6765 3404 6852 3414
rect 6765 3384 6774 3404
rect 6794 3384 6852 3404
rect 6765 3375 6852 3384
rect 6765 3374 6802 3375
rect 5063 3348 5073 3366
rect 5091 3348 5100 3366
rect 4884 3339 4921 3340
rect 5063 3339 5100 3348
rect 4307 3318 4343 3339
rect 4733 3318 4764 3339
rect 6821 3322 6852 3375
rect 6882 3404 6919 3475
rect 7090 3480 7483 3500
rect 7503 3480 7506 3500
rect 7090 3475 7506 3480
rect 7090 3474 7431 3475
rect 7034 3414 7065 3415
rect 6882 3384 6891 3404
rect 6911 3384 6919 3404
rect 6882 3374 6919 3384
rect 6978 3407 7065 3414
rect 6978 3404 7039 3407
rect 6978 3384 6987 3404
rect 7007 3387 7039 3404
rect 7060 3387 7065 3407
rect 7007 3384 7065 3387
rect 6978 3377 7065 3384
rect 7090 3404 7127 3474
rect 7393 3473 7430 3474
rect 7242 3414 7278 3415
rect 7090 3384 7099 3404
rect 7119 3384 7127 3404
rect 6978 3375 7034 3377
rect 6978 3374 7015 3375
rect 7090 3374 7127 3384
rect 7186 3404 7334 3414
rect 7434 3411 7530 3413
rect 7186 3384 7195 3404
rect 7215 3384 7305 3404
rect 7325 3384 7334 3404
rect 7186 3375 7334 3384
rect 7392 3404 7530 3411
rect 7392 3384 7401 3404
rect 7421 3384 7530 3404
rect 7392 3375 7530 3384
rect 7186 3374 7223 3375
rect 7242 3323 7278 3375
rect 7297 3374 7334 3375
rect 7393 3374 7430 3375
rect 6713 3321 6754 3322
rect 4140 3314 4240 3318
rect 4140 3310 4202 3314
rect 4140 3284 4147 3310
rect 4173 3288 4202 3310
rect 4228 3288 4240 3314
rect 4173 3284 4240 3288
rect 4140 3281 4240 3284
rect 4308 3281 4343 3318
rect 4405 3315 4764 3318
rect 4405 3310 4627 3315
rect 4405 3286 4418 3310
rect 4442 3291 4627 3310
rect 4651 3291 4764 3315
rect 4442 3286 4764 3291
rect 4405 3282 4764 3286
rect 4831 3310 4980 3318
rect 4831 3290 4842 3310
rect 4862 3290 4980 3310
rect 6605 3314 6754 3321
rect 5417 3306 5454 3308
rect 5417 3305 6065 3306
rect 4831 3283 4980 3290
rect 5416 3299 6065 3305
rect 4831 3282 4872 3283
rect 4155 3229 4192 3230
rect 4251 3229 4288 3230
rect 4307 3229 4343 3281
rect 4362 3229 4399 3230
rect 4055 3220 4193 3229
rect 3043 3201 3211 3202
rect 3043 3198 3487 3201
rect 3043 3179 3418 3198
rect 3438 3179 3487 3198
rect 4055 3200 4164 3220
rect 4184 3200 4193 3220
rect 3043 3175 3487 3179
rect 3043 3173 3211 3175
rect 3043 2995 3070 3173
rect 3110 3135 3174 3147
rect 3450 3143 3487 3175
rect 3658 3174 3907 3196
rect 4055 3193 4193 3200
rect 4251 3220 4399 3229
rect 4251 3200 4260 3220
rect 4280 3200 4370 3220
rect 4390 3200 4399 3220
rect 4055 3191 4151 3193
rect 4251 3190 4399 3200
rect 4458 3220 4495 3230
rect 4570 3229 4607 3230
rect 4551 3227 4607 3229
rect 4458 3200 4466 3220
rect 4486 3200 4495 3220
rect 4307 3189 4343 3190
rect 3658 3143 3695 3174
rect 3871 3172 3907 3174
rect 3871 3143 3908 3172
rect 3110 3134 3145 3135
rect 3087 3129 3145 3134
rect 3087 3109 3090 3129
rect 3110 3115 3145 3129
rect 3165 3115 3174 3135
rect 3110 3107 3174 3115
rect 3136 3106 3174 3107
rect 3137 3105 3174 3106
rect 3240 3139 3276 3140
rect 3348 3139 3384 3140
rect 3240 3131 3384 3139
rect 3240 3111 3248 3131
rect 3268 3111 3300 3131
rect 3324 3111 3356 3131
rect 3376 3111 3384 3131
rect 3240 3105 3384 3111
rect 3450 3135 3488 3143
rect 3556 3139 3592 3140
rect 3450 3115 3459 3135
rect 3479 3115 3488 3135
rect 3450 3106 3488 3115
rect 3507 3132 3592 3139
rect 3507 3112 3514 3132
rect 3535 3131 3592 3132
rect 3535 3112 3564 3131
rect 3507 3111 3564 3112
rect 3584 3111 3592 3131
rect 3450 3105 3487 3106
rect 3507 3105 3592 3111
rect 3658 3135 3696 3143
rect 3769 3139 3805 3140
rect 3658 3115 3667 3135
rect 3687 3115 3696 3135
rect 3658 3106 3696 3115
rect 3720 3131 3805 3139
rect 3720 3111 3777 3131
rect 3797 3111 3805 3131
rect 3658 3105 3695 3106
rect 3720 3105 3805 3111
rect 3871 3135 3909 3143
rect 3871 3115 3880 3135
rect 3900 3115 3909 3135
rect 4155 3130 4192 3131
rect 4458 3130 4495 3200
rect 4520 3220 4607 3227
rect 4520 3217 4578 3220
rect 4520 3197 4525 3217
rect 4546 3200 4578 3217
rect 4598 3200 4607 3220
rect 4546 3197 4607 3200
rect 4520 3190 4607 3197
rect 4666 3220 4703 3230
rect 4666 3200 4674 3220
rect 4694 3200 4703 3220
rect 4520 3189 4551 3190
rect 4154 3129 4495 3130
rect 3871 3106 3909 3115
rect 4079 3124 4495 3129
rect 3871 3105 3908 3106
rect 3294 3084 3330 3105
rect 3720 3084 3751 3105
rect 4079 3104 4082 3124
rect 4102 3104 4495 3124
rect 4666 3129 4703 3200
rect 4733 3229 4764 3282
rect 5416 3281 5426 3299
rect 5444 3285 6065 3299
rect 6605 3294 6723 3314
rect 6743 3294 6754 3314
rect 6605 3286 6754 3294
rect 6821 3318 7180 3322
rect 6821 3313 7143 3318
rect 6821 3289 6934 3313
rect 6958 3294 7143 3313
rect 7167 3294 7180 3318
rect 6958 3289 7180 3294
rect 6821 3286 7180 3289
rect 7242 3286 7277 3323
rect 7345 3320 7445 3323
rect 7345 3316 7412 3320
rect 7345 3290 7357 3316
rect 7383 3294 7412 3316
rect 7438 3294 7445 3320
rect 7383 3290 7445 3294
rect 7345 3286 7445 3290
rect 5444 3281 5454 3285
rect 5895 3284 6065 3285
rect 5066 3267 5103 3277
rect 5066 3249 5075 3267
rect 5093 3249 5103 3267
rect 5066 3240 5103 3249
rect 5416 3271 5454 3281
rect 4783 3229 4820 3230
rect 4733 3220 4820 3229
rect 4733 3200 4791 3220
rect 4811 3200 4820 3220
rect 4733 3190 4820 3200
rect 4879 3220 4916 3230
rect 4879 3200 4887 3220
rect 4907 3200 4916 3220
rect 4733 3189 4764 3190
rect 4879 3129 4916 3200
rect 5071 3175 5102 3240
rect 5416 3193 5451 3271
rect 6028 3261 6065 3284
rect 6821 3265 6852 3286
rect 7242 3265 7278 3286
rect 6664 3264 6701 3265
rect 5412 3184 5451 3193
rect 5070 3165 5107 3175
rect 5070 3163 5080 3165
rect 5004 3161 5080 3163
rect 4666 3105 4916 3129
rect 5001 3147 5080 3161
rect 5098 3147 5107 3165
rect 5412 3166 5422 3184
rect 5440 3166 5451 3184
rect 5412 3160 5451 3166
rect 5607 3236 5857 3260
rect 5607 3165 5644 3236
rect 5759 3175 5790 3176
rect 5412 3156 5449 3160
rect 5001 3144 5107 3147
rect 4473 3085 4494 3104
rect 5001 3085 5027 3144
rect 5070 3138 5107 3144
rect 5607 3145 5616 3165
rect 5636 3145 5644 3165
rect 5607 3135 5644 3145
rect 5703 3165 5790 3175
rect 5703 3145 5712 3165
rect 5732 3145 5790 3165
rect 5703 3136 5790 3145
rect 5703 3135 5740 3136
rect 5415 3085 5452 3094
rect 3127 3080 3227 3084
rect 3127 3076 3189 3080
rect 3127 3050 3134 3076
rect 3160 3054 3189 3076
rect 3215 3054 3227 3080
rect 3160 3050 3227 3054
rect 3127 3047 3227 3050
rect 3295 3047 3330 3084
rect 3392 3081 3751 3084
rect 3392 3076 3614 3081
rect 3392 3052 3405 3076
rect 3429 3057 3614 3076
rect 3638 3057 3751 3081
rect 3429 3052 3751 3057
rect 3392 3048 3751 3052
rect 3818 3076 3967 3084
rect 3818 3056 3829 3076
rect 3849 3056 3967 3076
rect 4473 3067 5027 3085
rect 5073 3074 5110 3076
rect 5001 3066 5027 3067
rect 5070 3066 5110 3074
rect 3818 3049 3967 3056
rect 5070 3054 5082 3066
rect 5061 3049 5082 3054
rect 3818 3048 3859 3049
rect 4477 3048 5082 3049
rect 5100 3048 5110 3066
rect 3142 2995 3179 2996
rect 3238 2995 3275 2996
rect 3294 2995 3330 3047
rect 3349 2995 3386 2996
rect 3042 2986 3180 2995
rect 3042 2966 3151 2986
rect 3171 2966 3180 2986
rect 3042 2959 3180 2966
rect 3238 2986 3386 2995
rect 3238 2966 3247 2986
rect 3267 2966 3357 2986
rect 3377 2966 3386 2986
rect 3042 2957 3138 2959
rect 3238 2956 3386 2966
rect 3445 2986 3482 2996
rect 3557 2995 3594 2996
rect 3538 2993 3594 2995
rect 3445 2966 3453 2986
rect 3473 2966 3482 2986
rect 3294 2955 3330 2956
rect 3142 2896 3179 2897
rect 3445 2896 3482 2966
rect 3507 2986 3594 2993
rect 3507 2983 3565 2986
rect 3507 2963 3512 2983
rect 3533 2966 3565 2983
rect 3585 2966 3594 2986
rect 3533 2963 3594 2966
rect 3507 2956 3594 2963
rect 3653 2986 3690 2996
rect 3653 2966 3661 2986
rect 3681 2966 3690 2986
rect 3507 2955 3538 2956
rect 3141 2895 3482 2896
rect 3066 2890 3482 2895
rect 3066 2870 3069 2890
rect 3089 2870 3482 2890
rect 3653 2895 3690 2966
rect 3720 2995 3751 3048
rect 4477 3039 5110 3048
rect 5413 3067 5424 3085
rect 5442 3067 5452 3085
rect 5759 3083 5790 3136
rect 5820 3165 5857 3236
rect 6028 3241 6421 3261
rect 6441 3241 6444 3261
rect 6028 3236 6444 3241
rect 6663 3255 6701 3264
rect 6028 3235 6369 3236
rect 6663 3235 6672 3255
rect 6692 3235 6701 3255
rect 5972 3175 6003 3176
rect 5820 3145 5829 3165
rect 5849 3145 5857 3165
rect 5820 3135 5857 3145
rect 5916 3168 6003 3175
rect 5916 3165 5977 3168
rect 5916 3145 5925 3165
rect 5945 3148 5977 3165
rect 5998 3148 6003 3168
rect 5945 3145 6003 3148
rect 5916 3138 6003 3145
rect 6028 3165 6065 3235
rect 6331 3234 6368 3235
rect 6663 3227 6701 3235
rect 6767 3259 6852 3265
rect 6877 3264 6914 3265
rect 6767 3239 6775 3259
rect 6795 3239 6852 3259
rect 6767 3231 6852 3239
rect 6876 3255 6914 3264
rect 6876 3235 6885 3255
rect 6905 3235 6914 3255
rect 6767 3230 6803 3231
rect 6876 3227 6914 3235
rect 6980 3259 7065 3265
rect 7085 3264 7122 3265
rect 6980 3239 6988 3259
rect 7008 3258 7065 3259
rect 7008 3239 7037 3258
rect 6980 3238 7037 3239
rect 7058 3238 7065 3258
rect 6980 3231 7065 3238
rect 7084 3255 7122 3264
rect 7084 3235 7093 3255
rect 7113 3235 7122 3255
rect 6980 3230 7016 3231
rect 7084 3227 7122 3235
rect 7188 3259 7332 3265
rect 7188 3239 7196 3259
rect 7216 3257 7304 3259
rect 7216 3240 7252 3257
rect 7276 3240 7304 3257
rect 7216 3239 7304 3240
rect 7324 3239 7332 3259
rect 7188 3231 7332 3239
rect 7188 3230 7224 3231
rect 7296 3230 7332 3231
rect 7398 3264 7435 3265
rect 7398 3263 7436 3264
rect 7398 3255 7462 3263
rect 7398 3235 7407 3255
rect 7427 3241 7462 3255
rect 7482 3241 7485 3261
rect 7427 3236 7485 3241
rect 7427 3235 7462 3236
rect 6664 3198 6701 3227
rect 6665 3196 6701 3198
rect 6877 3196 6914 3227
rect 6180 3175 6216 3176
rect 6028 3145 6037 3165
rect 6057 3145 6065 3165
rect 5916 3136 5972 3138
rect 5916 3135 5953 3136
rect 6028 3135 6065 3145
rect 6124 3165 6272 3175
rect 6665 3174 6914 3196
rect 7085 3195 7122 3227
rect 7398 3223 7462 3235
rect 7502 3197 7529 3375
rect 7361 3195 7529 3197
rect 7085 3184 7529 3195
rect 6372 3172 6468 3174
rect 6124 3145 6133 3165
rect 6153 3145 6243 3165
rect 6263 3145 6272 3165
rect 6124 3136 6272 3145
rect 6330 3165 6468 3172
rect 7085 3169 7531 3184
rect 7361 3168 7531 3169
rect 6330 3145 6339 3165
rect 6359 3145 6468 3165
rect 6330 3136 6468 3145
rect 6124 3135 6161 3136
rect 6180 3084 6216 3136
rect 6235 3135 6272 3136
rect 6331 3135 6368 3136
rect 5651 3082 5692 3083
rect 4477 3032 5109 3039
rect 4477 3030 4539 3032
rect 4055 3020 4223 3021
rect 4477 3020 4499 3030
rect 3770 2995 3807 2996
rect 3720 2986 3807 2995
rect 3720 2966 3778 2986
rect 3798 2966 3807 2986
rect 3720 2956 3807 2966
rect 3866 2986 3903 2996
rect 3866 2966 3874 2986
rect 3894 2966 3903 2986
rect 3720 2955 3751 2956
rect 3866 2895 3903 2966
rect 3653 2871 3903 2895
rect 4055 2994 4499 3020
rect 4055 2992 4223 2994
rect 4055 2814 4082 2992
rect 4122 2954 4186 2966
rect 4462 2962 4499 2994
rect 4670 2993 4919 3015
rect 4670 2962 4707 2993
rect 4883 2991 4919 2993
rect 4883 2962 4920 2991
rect 4122 2953 4157 2954
rect 4099 2948 4157 2953
rect 4099 2928 4102 2948
rect 4122 2934 4157 2948
rect 4177 2934 4186 2954
rect 4122 2926 4186 2934
rect 4148 2925 4186 2926
rect 4149 2924 4186 2925
rect 4252 2958 4288 2959
rect 4360 2958 4396 2959
rect 4252 2950 4396 2958
rect 4252 2930 4260 2950
rect 4280 2930 4309 2950
rect 4252 2929 4309 2930
rect 4331 2930 4368 2950
rect 4388 2930 4396 2950
rect 4331 2929 4396 2930
rect 4252 2924 4396 2929
rect 4462 2954 4500 2962
rect 4568 2958 4604 2959
rect 4462 2934 4471 2954
rect 4491 2934 4500 2954
rect 4462 2925 4500 2934
rect 4519 2951 4604 2958
rect 4519 2931 4526 2951
rect 4547 2950 4604 2951
rect 4547 2931 4576 2950
rect 4519 2930 4576 2931
rect 4596 2930 4604 2950
rect 4462 2924 4499 2925
rect 4519 2924 4604 2930
rect 4670 2954 4708 2962
rect 4781 2958 4817 2959
rect 4670 2934 4679 2954
rect 4699 2934 4708 2954
rect 4670 2925 4708 2934
rect 4732 2950 4817 2958
rect 4732 2930 4789 2950
rect 4809 2930 4817 2950
rect 4670 2924 4707 2925
rect 4732 2924 4817 2930
rect 4883 2954 4921 2962
rect 4883 2934 4892 2954
rect 4912 2934 4921 2954
rect 4883 2925 4921 2934
rect 4883 2924 4920 2925
rect 4306 2903 4342 2924
rect 4732 2903 4763 2924
rect 4139 2899 4239 2903
rect 4139 2895 4201 2899
rect 4139 2869 4146 2895
rect 4172 2873 4201 2895
rect 4227 2873 4239 2899
rect 4172 2869 4239 2873
rect 4139 2866 4239 2869
rect 4307 2866 4342 2903
rect 4404 2900 4763 2903
rect 4404 2895 4626 2900
rect 4404 2871 4417 2895
rect 4441 2876 4626 2895
rect 4650 2876 4763 2900
rect 4441 2871 4763 2876
rect 4404 2867 4763 2871
rect 4830 2895 4979 2903
rect 4830 2875 4841 2895
rect 4861 2875 4979 2895
rect 4830 2868 4979 2875
rect 5070 2883 5109 3032
rect 5413 2918 5452 3067
rect 5543 3075 5692 3082
rect 5543 3055 5661 3075
rect 5681 3055 5692 3075
rect 5543 3047 5692 3055
rect 5759 3079 6118 3083
rect 5759 3074 6081 3079
rect 5759 3050 5872 3074
rect 5896 3055 6081 3074
rect 6105 3055 6118 3079
rect 5896 3050 6118 3055
rect 5759 3047 6118 3050
rect 6180 3047 6215 3084
rect 6283 3081 6383 3084
rect 6283 3077 6350 3081
rect 6283 3051 6295 3077
rect 6321 3055 6350 3077
rect 6376 3055 6383 3081
rect 6321 3051 6383 3055
rect 6283 3047 6383 3051
rect 5759 3026 5790 3047
rect 6180 3026 6216 3047
rect 5602 3025 5639 3026
rect 5601 3016 5639 3025
rect 5601 2996 5610 3016
rect 5630 2996 5639 3016
rect 5601 2988 5639 2996
rect 5705 3020 5790 3026
rect 5815 3025 5852 3026
rect 5705 3000 5713 3020
rect 5733 3000 5790 3020
rect 5705 2992 5790 3000
rect 5814 3016 5852 3025
rect 5814 2996 5823 3016
rect 5843 2996 5852 3016
rect 5705 2991 5741 2992
rect 5814 2988 5852 2996
rect 5918 3020 6003 3026
rect 6023 3025 6060 3026
rect 5918 3000 5926 3020
rect 5946 3019 6003 3020
rect 5946 3000 5975 3019
rect 5918 2999 5975 3000
rect 5996 2999 6003 3019
rect 5918 2992 6003 2999
rect 6022 3016 6060 3025
rect 6022 2996 6031 3016
rect 6051 2996 6060 3016
rect 5918 2991 5954 2992
rect 6022 2988 6060 2996
rect 6126 3021 6270 3026
rect 6126 3020 6191 3021
rect 6126 3000 6134 3020
rect 6154 3000 6191 3020
rect 6213 3020 6270 3021
rect 6213 3000 6242 3020
rect 6262 3000 6270 3020
rect 6126 2992 6270 3000
rect 6126 2991 6162 2992
rect 6234 2991 6270 2992
rect 6336 3025 6373 3026
rect 6336 3024 6374 3025
rect 6336 3016 6400 3024
rect 6336 2996 6345 3016
rect 6365 3002 6400 3016
rect 6420 3002 6423 3022
rect 6365 2997 6423 3002
rect 6365 2996 6400 2997
rect 5602 2959 5639 2988
rect 5603 2957 5639 2959
rect 5815 2957 5852 2988
rect 5603 2935 5852 2957
rect 6023 2956 6060 2988
rect 6336 2984 6400 2996
rect 6440 2958 6467 3136
rect 6299 2956 6467 2958
rect 6023 2930 6467 2956
rect 6619 3055 6869 3079
rect 6619 2984 6656 3055
rect 6771 2994 6802 2995
rect 6619 2964 6628 2984
rect 6648 2964 6656 2984
rect 6619 2954 6656 2964
rect 6715 2984 6802 2994
rect 6715 2964 6724 2984
rect 6744 2964 6802 2984
rect 6715 2955 6802 2964
rect 6715 2954 6752 2955
rect 6023 2920 6045 2930
rect 6299 2929 6467 2930
rect 5983 2918 6045 2920
rect 5413 2911 6045 2918
rect 4830 2867 4871 2868
rect 4154 2814 4191 2815
rect 4250 2814 4287 2815
rect 4306 2814 4342 2866
rect 4361 2814 4398 2815
rect 4054 2805 4192 2814
rect 4054 2785 4163 2805
rect 4183 2785 4192 2805
rect 4054 2778 4192 2785
rect 4250 2805 4398 2814
rect 4250 2785 4259 2805
rect 4279 2785 4369 2805
rect 4389 2785 4398 2805
rect 4054 2776 4150 2778
rect 4250 2775 4398 2785
rect 4457 2805 4494 2815
rect 4569 2814 4606 2815
rect 4550 2812 4606 2814
rect 4457 2785 4465 2805
rect 4485 2785 4494 2805
rect 4306 2774 4342 2775
rect 2835 2734 3003 2735
rect 2835 2708 3279 2734
rect 2835 2706 3003 2708
rect 2835 2528 2862 2706
rect 2902 2668 2966 2680
rect 3242 2676 3279 2708
rect 3450 2707 3699 2729
rect 4154 2715 4191 2716
rect 4457 2715 4494 2785
rect 4519 2805 4606 2812
rect 4519 2802 4577 2805
rect 4519 2782 4524 2802
rect 4545 2785 4577 2802
rect 4597 2785 4606 2805
rect 4545 2782 4606 2785
rect 4519 2775 4606 2782
rect 4665 2805 4702 2815
rect 4665 2785 4673 2805
rect 4693 2785 4702 2805
rect 4519 2774 4550 2775
rect 4153 2714 4494 2715
rect 3450 2676 3487 2707
rect 3663 2705 3699 2707
rect 4078 2709 4494 2714
rect 3663 2676 3700 2705
rect 4078 2689 4081 2709
rect 4101 2689 4494 2709
rect 4665 2714 4702 2785
rect 4732 2814 4763 2867
rect 5070 2865 5080 2883
rect 5098 2865 5109 2883
rect 5412 2902 6045 2911
rect 6771 2902 6802 2955
rect 6832 2984 6869 3055
rect 7040 3060 7433 3080
rect 7453 3060 7456 3080
rect 7040 3055 7456 3060
rect 7040 3054 7381 3055
rect 6984 2994 7015 2995
rect 6832 2964 6841 2984
rect 6861 2964 6869 2984
rect 6832 2954 6869 2964
rect 6928 2987 7015 2994
rect 6928 2984 6989 2987
rect 6928 2964 6937 2984
rect 6957 2967 6989 2984
rect 7010 2967 7015 2987
rect 6957 2964 7015 2967
rect 6928 2957 7015 2964
rect 7040 2984 7077 3054
rect 7343 3053 7380 3054
rect 7192 2994 7228 2995
rect 7040 2964 7049 2984
rect 7069 2964 7077 2984
rect 6928 2955 6984 2957
rect 6928 2954 6965 2955
rect 7040 2954 7077 2964
rect 7136 2984 7284 2994
rect 7384 2991 7480 2993
rect 7136 2964 7145 2984
rect 7165 2964 7255 2984
rect 7275 2964 7284 2984
rect 7136 2955 7284 2964
rect 7342 2984 7480 2991
rect 7342 2964 7351 2984
rect 7371 2964 7480 2984
rect 7342 2955 7480 2964
rect 7136 2954 7173 2955
rect 7192 2903 7228 2955
rect 7247 2954 7284 2955
rect 7343 2954 7380 2955
rect 5412 2884 5422 2902
rect 5440 2901 6045 2902
rect 6663 2901 6704 2902
rect 5440 2896 5461 2901
rect 5440 2884 5452 2896
rect 6555 2894 6704 2901
rect 5412 2876 5452 2884
rect 5495 2883 5521 2884
rect 5412 2874 5449 2876
rect 5495 2865 6049 2883
rect 6555 2874 6673 2894
rect 6693 2874 6704 2894
rect 6555 2866 6704 2874
rect 6771 2898 7130 2902
rect 6771 2893 7093 2898
rect 6771 2869 6884 2893
rect 6908 2874 7093 2893
rect 7117 2874 7130 2898
rect 6908 2869 7130 2874
rect 6771 2866 7130 2869
rect 7192 2866 7227 2903
rect 7295 2900 7395 2903
rect 7295 2896 7362 2900
rect 7295 2870 7307 2896
rect 7333 2874 7362 2896
rect 7388 2874 7395 2900
rect 7333 2870 7395 2874
rect 7295 2866 7395 2870
rect 5070 2856 5107 2865
rect 4782 2814 4819 2815
rect 4732 2805 4819 2814
rect 4732 2785 4790 2805
rect 4810 2785 4819 2805
rect 4732 2775 4819 2785
rect 4878 2805 4915 2815
rect 4878 2785 4886 2805
rect 4906 2785 4915 2805
rect 5415 2806 5452 2812
rect 5495 2806 5521 2865
rect 6028 2846 6049 2865
rect 5415 2803 5521 2806
rect 5073 2790 5110 2794
rect 4732 2774 4763 2775
rect 4878 2714 4915 2785
rect 4665 2690 4915 2714
rect 5071 2784 5110 2790
rect 5071 2766 5082 2784
rect 5100 2766 5110 2784
rect 5415 2785 5424 2803
rect 5442 2789 5521 2803
rect 5606 2821 5856 2845
rect 5442 2787 5518 2789
rect 5442 2785 5452 2787
rect 5415 2775 5452 2785
rect 5071 2757 5110 2766
rect 2902 2667 2937 2668
rect 2879 2662 2937 2667
rect 2879 2642 2882 2662
rect 2902 2648 2937 2662
rect 2957 2648 2966 2668
rect 2902 2640 2966 2648
rect 2928 2639 2966 2640
rect 2929 2638 2966 2639
rect 3032 2672 3068 2673
rect 3140 2672 3176 2673
rect 3032 2666 3176 2672
rect 3032 2664 3093 2666
rect 3032 2644 3040 2664
rect 3060 2644 3093 2664
rect 3032 2640 3093 2644
rect 3118 2664 3176 2666
rect 3118 2644 3148 2664
rect 3168 2644 3176 2664
rect 3118 2640 3176 2644
rect 3032 2638 3176 2640
rect 3242 2668 3280 2676
rect 3348 2672 3384 2673
rect 3242 2648 3251 2668
rect 3271 2648 3280 2668
rect 3242 2639 3280 2648
rect 3299 2665 3384 2672
rect 3299 2645 3306 2665
rect 3327 2664 3384 2665
rect 3327 2645 3356 2664
rect 3299 2644 3356 2645
rect 3376 2644 3384 2664
rect 3242 2638 3279 2639
rect 3299 2638 3384 2644
rect 3450 2668 3488 2676
rect 3561 2672 3597 2673
rect 3450 2648 3459 2668
rect 3479 2648 3488 2668
rect 3450 2639 3488 2648
rect 3512 2664 3597 2672
rect 3512 2644 3569 2664
rect 3589 2644 3597 2664
rect 3450 2638 3487 2639
rect 3512 2638 3597 2644
rect 3663 2668 3701 2676
rect 3663 2648 3672 2668
rect 3692 2648 3701 2668
rect 3663 2639 3701 2648
rect 4457 2666 4494 2689
rect 5071 2679 5106 2757
rect 5420 2710 5451 2775
rect 5606 2750 5643 2821
rect 5758 2760 5789 2761
rect 5606 2730 5615 2750
rect 5635 2730 5643 2750
rect 5606 2720 5643 2730
rect 5702 2750 5789 2760
rect 5702 2730 5711 2750
rect 5731 2730 5789 2750
rect 5702 2721 5789 2730
rect 5702 2720 5739 2721
rect 5068 2669 5106 2679
rect 5419 2701 5456 2710
rect 5419 2683 5429 2701
rect 5447 2683 5456 2701
rect 5419 2673 5456 2683
rect 4457 2665 4627 2666
rect 5068 2665 5078 2669
rect 4457 2651 5078 2665
rect 5096 2651 5106 2669
rect 5758 2668 5789 2721
rect 5819 2750 5856 2821
rect 6027 2826 6420 2846
rect 6440 2826 6443 2846
rect 6771 2845 6802 2866
rect 7192 2845 7228 2866
rect 6614 2844 6651 2845
rect 6027 2821 6443 2826
rect 6613 2835 6651 2844
rect 6027 2820 6368 2821
rect 5971 2760 6002 2761
rect 5819 2730 5828 2750
rect 5848 2730 5856 2750
rect 5819 2720 5856 2730
rect 5915 2753 6002 2760
rect 5915 2750 5976 2753
rect 5915 2730 5924 2750
rect 5944 2733 5976 2750
rect 5997 2733 6002 2753
rect 5944 2730 6002 2733
rect 5915 2723 6002 2730
rect 6027 2750 6064 2820
rect 6330 2819 6367 2820
rect 6613 2815 6622 2835
rect 6642 2815 6651 2835
rect 6613 2807 6651 2815
rect 6717 2839 6802 2845
rect 6827 2844 6864 2845
rect 6717 2819 6725 2839
rect 6745 2819 6802 2839
rect 6717 2811 6802 2819
rect 6826 2835 6864 2844
rect 6826 2815 6835 2835
rect 6855 2815 6864 2835
rect 6717 2810 6753 2811
rect 6826 2807 6864 2815
rect 6930 2839 7015 2845
rect 7035 2844 7072 2845
rect 6930 2819 6938 2839
rect 6958 2838 7015 2839
rect 6958 2819 6987 2838
rect 6930 2818 6987 2819
rect 7008 2818 7015 2838
rect 6930 2811 7015 2818
rect 7034 2835 7072 2844
rect 7034 2815 7043 2835
rect 7063 2815 7072 2835
rect 6930 2810 6966 2811
rect 7034 2807 7072 2815
rect 7138 2840 7282 2845
rect 7138 2839 7197 2840
rect 7138 2819 7146 2839
rect 7166 2820 7197 2839
rect 7221 2839 7282 2840
rect 7221 2820 7254 2839
rect 7166 2819 7254 2820
rect 7274 2819 7282 2839
rect 7138 2811 7282 2819
rect 7138 2810 7174 2811
rect 7246 2810 7282 2811
rect 7348 2844 7385 2845
rect 7348 2843 7386 2844
rect 7348 2835 7412 2843
rect 7348 2815 7357 2835
rect 7377 2821 7412 2835
rect 7432 2821 7435 2841
rect 7377 2816 7435 2821
rect 7377 2815 7412 2816
rect 6614 2778 6651 2807
rect 6615 2776 6651 2778
rect 6827 2776 6864 2807
rect 6179 2760 6215 2761
rect 6027 2730 6036 2750
rect 6056 2730 6064 2750
rect 5915 2721 5971 2723
rect 5915 2720 5952 2721
rect 6027 2720 6064 2730
rect 6123 2750 6271 2760
rect 6371 2757 6467 2759
rect 6123 2730 6132 2750
rect 6152 2730 6242 2750
rect 6262 2730 6271 2750
rect 6123 2721 6271 2730
rect 6329 2750 6467 2757
rect 6615 2754 6864 2776
rect 7035 2775 7072 2807
rect 7348 2803 7412 2815
rect 7452 2777 7479 2955
rect 7311 2775 7479 2777
rect 7035 2771 7479 2775
rect 6329 2730 6338 2750
rect 6358 2730 6467 2750
rect 7035 2752 7084 2771
rect 7104 2752 7479 2771
rect 7035 2749 7479 2752
rect 7311 2748 7479 2749
rect 7500 2774 7531 3168
rect 7500 2748 7505 2774
rect 7524 2748 7531 2774
rect 7500 2745 7531 2748
rect 6329 2721 6467 2730
rect 6123 2720 6160 2721
rect 6179 2669 6215 2721
rect 6234 2720 6271 2721
rect 6330 2720 6367 2721
rect 5650 2667 5691 2668
rect 4457 2645 5106 2651
rect 5542 2660 5691 2667
rect 4457 2644 5105 2645
rect 5068 2642 5105 2644
rect 5542 2640 5660 2660
rect 5680 2640 5691 2660
rect 3663 2638 3700 2639
rect 3086 2617 3122 2638
rect 3512 2617 3543 2638
rect 5542 2632 5691 2640
rect 5758 2664 6117 2668
rect 5758 2659 6080 2664
rect 5758 2635 5871 2659
rect 5895 2640 6080 2659
rect 6104 2640 6117 2664
rect 5895 2635 6117 2640
rect 5758 2632 6117 2635
rect 6179 2632 6214 2669
rect 6282 2666 6382 2669
rect 6282 2662 6349 2666
rect 6282 2636 6294 2662
rect 6320 2640 6349 2662
rect 6375 2640 6382 2666
rect 6320 2636 6382 2640
rect 6282 2632 6382 2636
rect 2919 2613 3019 2617
rect 2919 2609 2981 2613
rect 2919 2583 2926 2609
rect 2952 2587 2981 2609
rect 3007 2587 3019 2613
rect 2952 2583 3019 2587
rect 2919 2580 3019 2583
rect 3087 2580 3122 2617
rect 3184 2614 3543 2617
rect 3184 2609 3406 2614
rect 3184 2585 3197 2609
rect 3221 2590 3406 2609
rect 3430 2590 3543 2614
rect 3221 2585 3543 2590
rect 3184 2581 3543 2585
rect 3610 2609 3759 2617
rect 5758 2611 5789 2632
rect 6179 2611 6215 2632
rect 3610 2589 3621 2609
rect 3641 2589 3759 2609
rect 3610 2582 3759 2589
rect 5422 2602 5459 2611
rect 5601 2610 5638 2611
rect 5422 2584 5431 2602
rect 5449 2584 5459 2602
rect 3610 2581 3651 2582
rect 2934 2528 2971 2529
rect 3030 2528 3067 2529
rect 3086 2528 3122 2580
rect 3141 2528 3178 2529
rect 2834 2519 2972 2528
rect 2834 2499 2943 2519
rect 2963 2499 2972 2519
rect 2834 2492 2972 2499
rect 3030 2519 3178 2528
rect 3030 2499 3039 2519
rect 3059 2499 3149 2519
rect 3169 2499 3178 2519
rect 2834 2490 2930 2492
rect 3030 2489 3178 2499
rect 3237 2519 3274 2529
rect 3349 2528 3386 2529
rect 3330 2526 3386 2528
rect 3237 2499 3245 2519
rect 3265 2499 3274 2519
rect 3086 2488 3122 2489
rect 2934 2429 2971 2430
rect 3237 2429 3274 2499
rect 3299 2519 3386 2526
rect 3299 2516 3357 2519
rect 3299 2496 3304 2516
rect 3325 2499 3357 2516
rect 3377 2499 3386 2519
rect 3325 2496 3386 2499
rect 3299 2489 3386 2496
rect 3445 2519 3482 2529
rect 3445 2499 3453 2519
rect 3473 2499 3482 2519
rect 3299 2488 3330 2489
rect 2933 2428 3274 2429
rect 2858 2423 3274 2428
rect 2858 2403 2861 2423
rect 2881 2403 3274 2423
rect 3445 2428 3482 2499
rect 3512 2528 3543 2581
rect 5071 2570 5108 2580
rect 5422 2574 5459 2584
rect 5071 2552 5080 2570
rect 5098 2552 5108 2570
rect 5071 2543 5108 2552
rect 3562 2528 3599 2529
rect 3512 2519 3599 2528
rect 3512 2499 3570 2519
rect 3590 2499 3599 2519
rect 3512 2489 3599 2499
rect 3658 2519 3695 2529
rect 3658 2499 3666 2519
rect 3686 2499 3695 2519
rect 3512 2488 3543 2489
rect 3658 2428 3695 2499
rect 5071 2497 5106 2543
rect 5423 2539 5459 2574
rect 5600 2601 5638 2610
rect 5600 2581 5609 2601
rect 5629 2581 5638 2601
rect 5600 2573 5638 2581
rect 5704 2605 5789 2611
rect 5814 2610 5851 2611
rect 5704 2585 5712 2605
rect 5732 2585 5789 2605
rect 5704 2577 5789 2585
rect 5813 2601 5851 2610
rect 5813 2581 5822 2601
rect 5842 2581 5851 2601
rect 5704 2576 5740 2577
rect 5813 2573 5851 2581
rect 5917 2605 6002 2611
rect 6022 2610 6059 2611
rect 5917 2585 5925 2605
rect 5945 2604 6002 2605
rect 5945 2585 5974 2604
rect 5917 2584 5974 2585
rect 5995 2584 6002 2604
rect 5917 2577 6002 2584
rect 6021 2601 6059 2610
rect 6021 2581 6030 2601
rect 6050 2581 6059 2601
rect 5917 2576 5953 2577
rect 6021 2573 6059 2581
rect 6125 2605 6269 2611
rect 6125 2585 6133 2605
rect 6153 2604 6241 2605
rect 6153 2585 6181 2604
rect 6125 2583 6181 2585
rect 6203 2585 6241 2604
rect 6261 2585 6269 2605
rect 6203 2583 6269 2585
rect 6125 2577 6269 2583
rect 6125 2576 6161 2577
rect 6233 2576 6269 2577
rect 6335 2610 6372 2611
rect 6335 2609 6373 2610
rect 6335 2601 6399 2609
rect 6335 2581 6344 2601
rect 6364 2587 6399 2601
rect 6419 2587 6422 2607
rect 6364 2582 6422 2587
rect 6364 2581 6399 2582
rect 5601 2544 5638 2573
rect 5421 2498 5459 2539
rect 5602 2542 5638 2544
rect 5814 2542 5851 2573
rect 5602 2520 5851 2542
rect 6022 2541 6059 2573
rect 6335 2569 6399 2581
rect 6439 2543 6466 2721
rect 6298 2541 6466 2543
rect 6022 2515 6466 2541
rect 6023 2498 6047 2515
rect 6298 2514 6466 2515
rect 6834 2543 7084 2567
rect 5070 2491 5108 2497
rect 4481 2473 5108 2491
rect 5421 2480 6048 2498
rect 5421 2474 5459 2480
rect 3445 2404 3695 2428
rect 4063 2456 4231 2457
rect 4482 2456 4506 2473
rect 4063 2430 4507 2456
rect 4063 2428 4231 2430
rect 2443 2291 2476 2351
rect 2245 2284 2413 2286
rect 1969 2258 2413 2284
rect 2245 2257 2413 2258
rect 2442 2280 2479 2291
rect 2442 2261 2448 2280
rect 2471 2261 2479 2280
rect 906 2217 942 2218
rect 754 2187 763 2207
rect 783 2187 791 2207
rect 642 2178 698 2180
rect 642 2177 679 2178
rect 754 2177 791 2187
rect 850 2207 998 2217
rect 1098 2214 1194 2216
rect 850 2187 859 2207
rect 879 2187 969 2207
rect 989 2187 998 2207
rect 850 2178 998 2187
rect 1056 2207 1194 2214
rect 1056 2187 1065 2207
rect 1085 2187 1194 2207
rect 1056 2178 1194 2187
rect 850 2177 887 2178
rect 906 2126 942 2178
rect 961 2177 998 2178
rect 1057 2177 1094 2178
rect 377 2124 418 2125
rect 139 1960 178 2109
rect 269 2117 418 2124
rect 269 2097 387 2117
rect 407 2097 418 2117
rect 269 2089 418 2097
rect 485 2121 844 2125
rect 485 2116 807 2121
rect 485 2092 598 2116
rect 622 2097 807 2116
rect 831 2097 844 2121
rect 622 2092 844 2097
rect 485 2089 844 2092
rect 906 2089 941 2126
rect 1009 2123 1109 2126
rect 1009 2119 1076 2123
rect 1009 2093 1021 2119
rect 1047 2097 1076 2119
rect 1102 2097 1109 2123
rect 1047 2093 1109 2097
rect 1009 2089 1109 2093
rect 485 2068 516 2089
rect 906 2068 942 2089
rect 328 2067 365 2068
rect 327 2058 365 2067
rect 327 2038 336 2058
rect 356 2038 365 2058
rect 327 2030 365 2038
rect 431 2062 516 2068
rect 541 2067 578 2068
rect 431 2042 439 2062
rect 459 2042 516 2062
rect 431 2034 516 2042
rect 540 2058 578 2067
rect 540 2038 549 2058
rect 569 2038 578 2058
rect 431 2033 467 2034
rect 540 2030 578 2038
rect 644 2062 729 2068
rect 749 2067 786 2068
rect 644 2042 652 2062
rect 672 2061 729 2062
rect 672 2042 701 2061
rect 644 2041 701 2042
rect 722 2041 729 2061
rect 644 2034 729 2041
rect 748 2058 786 2067
rect 748 2038 757 2058
rect 777 2038 786 2058
rect 644 2033 680 2034
rect 748 2030 786 2038
rect 852 2063 996 2068
rect 852 2062 917 2063
rect 852 2042 860 2062
rect 880 2042 917 2062
rect 939 2062 996 2063
rect 939 2042 968 2062
rect 988 2042 996 2062
rect 852 2034 996 2042
rect 852 2033 888 2034
rect 960 2033 996 2034
rect 1062 2067 1099 2068
rect 1062 2066 1100 2067
rect 1062 2058 1126 2066
rect 1062 2038 1071 2058
rect 1091 2044 1126 2058
rect 1146 2044 1149 2064
rect 1091 2039 1149 2044
rect 1091 2038 1126 2039
rect 328 2001 365 2030
rect 329 1999 365 2001
rect 541 1999 578 2030
rect 329 1977 578 1999
rect 749 1998 786 2030
rect 1062 2026 1126 2038
rect 1166 2000 1193 2178
rect 1025 1998 1193 2000
rect 749 1972 1193 1998
rect 1345 2097 1595 2121
rect 1345 2026 1382 2097
rect 1497 2036 1528 2037
rect 1345 2006 1354 2026
rect 1374 2006 1382 2026
rect 1345 1996 1382 2006
rect 1441 2026 1528 2036
rect 1441 2006 1450 2026
rect 1470 2006 1528 2026
rect 1441 1997 1528 2006
rect 1441 1996 1478 1997
rect 749 1962 771 1972
rect 1025 1971 1193 1972
rect 709 1960 771 1962
rect 139 1953 771 1960
rect 138 1944 771 1953
rect 1497 1944 1528 1997
rect 1558 2026 1595 2097
rect 1766 2102 2159 2122
rect 2179 2102 2182 2122
rect 1766 2097 2182 2102
rect 1766 2096 2107 2097
rect 1710 2036 1741 2037
rect 1558 2006 1567 2026
rect 1587 2006 1595 2026
rect 1558 1996 1595 2006
rect 1654 2029 1741 2036
rect 1654 2026 1715 2029
rect 1654 2006 1663 2026
rect 1683 2009 1715 2026
rect 1736 2009 1741 2029
rect 1683 2006 1741 2009
rect 1654 1999 1741 2006
rect 1766 2026 1803 2096
rect 2069 2095 2106 2096
rect 1918 2036 1954 2037
rect 1766 2006 1775 2026
rect 1795 2006 1803 2026
rect 1654 1997 1710 1999
rect 1654 1996 1691 1997
rect 1766 1996 1803 2006
rect 1862 2026 2010 2036
rect 2110 2033 2206 2035
rect 1862 2006 1871 2026
rect 1891 2006 1981 2026
rect 2001 2006 2010 2026
rect 1862 1997 2010 2006
rect 2068 2026 2206 2033
rect 2068 2006 2077 2026
rect 2097 2006 2206 2026
rect 2068 1997 2206 2006
rect 1862 1996 1899 1997
rect 1918 1945 1954 1997
rect 1973 1996 2010 1997
rect 2069 1996 2106 1997
rect 138 1926 148 1944
rect 166 1943 771 1944
rect 1389 1943 1430 1944
rect 166 1938 187 1943
rect 166 1926 178 1938
rect 1281 1936 1430 1943
rect 138 1918 178 1926
rect 221 1925 247 1926
rect 138 1916 175 1918
rect 221 1907 775 1925
rect 1281 1916 1399 1936
rect 1419 1916 1430 1936
rect 1281 1908 1430 1916
rect 1497 1940 1856 1944
rect 1497 1935 1819 1940
rect 1497 1911 1610 1935
rect 1634 1916 1819 1935
rect 1843 1916 1856 1940
rect 1634 1911 1856 1916
rect 1497 1908 1856 1911
rect 1918 1908 1953 1945
rect 2021 1942 2121 1945
rect 2021 1938 2088 1942
rect 2021 1912 2033 1938
rect 2059 1916 2088 1938
rect 2114 1916 2121 1942
rect 2059 1912 2121 1916
rect 2021 1908 2121 1912
rect 141 1848 178 1854
rect 221 1848 247 1907
rect 754 1888 775 1907
rect 141 1845 247 1848
rect 141 1827 150 1845
rect 168 1831 247 1845
rect 332 1863 582 1887
rect 168 1829 244 1831
rect 168 1827 178 1829
rect 141 1817 178 1827
rect 146 1752 177 1817
rect 332 1792 369 1863
rect 484 1802 515 1803
rect 332 1772 341 1792
rect 361 1772 369 1792
rect 332 1762 369 1772
rect 428 1792 515 1802
rect 428 1772 437 1792
rect 457 1772 515 1792
rect 428 1763 515 1772
rect 428 1762 465 1763
rect 145 1743 182 1752
rect 145 1725 155 1743
rect 173 1725 182 1743
rect 145 1715 182 1725
rect 484 1710 515 1763
rect 545 1792 582 1863
rect 753 1868 1146 1888
rect 1166 1868 1169 1888
rect 1497 1887 1528 1908
rect 1918 1887 1954 1908
rect 1340 1886 1377 1887
rect 753 1863 1169 1868
rect 1339 1877 1377 1886
rect 753 1862 1094 1863
rect 697 1802 728 1803
rect 545 1772 554 1792
rect 574 1772 582 1792
rect 545 1762 582 1772
rect 641 1795 728 1802
rect 641 1792 702 1795
rect 641 1772 650 1792
rect 670 1775 702 1792
rect 723 1775 728 1795
rect 670 1772 728 1775
rect 641 1765 728 1772
rect 753 1792 790 1862
rect 1056 1861 1093 1862
rect 1339 1857 1348 1877
rect 1368 1857 1377 1877
rect 1339 1849 1377 1857
rect 1443 1881 1528 1887
rect 1553 1886 1590 1887
rect 1443 1861 1451 1881
rect 1471 1861 1528 1881
rect 1443 1853 1528 1861
rect 1552 1877 1590 1886
rect 1552 1857 1561 1877
rect 1581 1857 1590 1877
rect 1443 1852 1479 1853
rect 1552 1849 1590 1857
rect 1656 1881 1741 1887
rect 1761 1886 1798 1887
rect 1656 1861 1664 1881
rect 1684 1880 1741 1881
rect 1684 1861 1713 1880
rect 1656 1860 1713 1861
rect 1734 1860 1741 1880
rect 1656 1853 1741 1860
rect 1760 1877 1798 1886
rect 1760 1857 1769 1877
rect 1789 1857 1798 1877
rect 1656 1852 1692 1853
rect 1760 1849 1798 1857
rect 1864 1881 2008 1887
rect 1864 1861 1872 1881
rect 1892 1861 1924 1881
rect 1948 1861 1980 1881
rect 2000 1861 2008 1881
rect 1864 1853 2008 1861
rect 1864 1852 1900 1853
rect 1972 1852 2008 1853
rect 2074 1886 2111 1887
rect 2074 1885 2112 1886
rect 2074 1877 2138 1885
rect 2074 1857 2083 1877
rect 2103 1863 2138 1877
rect 2158 1863 2161 1883
rect 2103 1858 2161 1863
rect 2103 1857 2138 1858
rect 1340 1820 1377 1849
rect 1341 1818 1377 1820
rect 1553 1818 1590 1849
rect 905 1802 941 1803
rect 753 1772 762 1792
rect 782 1772 790 1792
rect 641 1763 697 1765
rect 641 1762 678 1763
rect 753 1762 790 1772
rect 849 1792 997 1802
rect 1097 1799 1193 1801
rect 849 1772 858 1792
rect 878 1772 968 1792
rect 988 1772 997 1792
rect 849 1763 997 1772
rect 1055 1792 1193 1799
rect 1341 1796 1590 1818
rect 1761 1817 1798 1849
rect 2074 1845 2138 1857
rect 2178 1819 2205 1997
rect 2037 1817 2205 1819
rect 1761 1813 2205 1817
rect 1055 1772 1064 1792
rect 1084 1772 1193 1792
rect 1761 1794 1810 1813
rect 1830 1794 2205 1813
rect 1761 1791 2205 1794
rect 2037 1790 2205 1791
rect 1055 1763 1193 1772
rect 849 1762 886 1763
rect 905 1711 941 1763
rect 960 1762 997 1763
rect 1056 1762 1093 1763
rect 376 1709 417 1710
rect 268 1702 417 1709
rect 268 1682 386 1702
rect 406 1682 417 1702
rect 268 1674 417 1682
rect 484 1706 843 1710
rect 484 1701 806 1706
rect 484 1677 597 1701
rect 621 1682 806 1701
rect 830 1682 843 1706
rect 621 1677 843 1682
rect 484 1674 843 1677
rect 905 1674 940 1711
rect 1008 1708 1108 1711
rect 1008 1704 1075 1708
rect 1008 1678 1020 1704
rect 1046 1682 1075 1704
rect 1101 1682 1108 1708
rect 1046 1678 1108 1682
rect 1008 1674 1108 1678
rect 484 1653 515 1674
rect 905 1653 941 1674
rect 148 1644 185 1653
rect 327 1652 364 1653
rect 148 1626 157 1644
rect 175 1626 185 1644
rect 148 1616 185 1626
rect 149 1581 185 1616
rect 326 1643 364 1652
rect 326 1623 335 1643
rect 355 1623 364 1643
rect 326 1615 364 1623
rect 430 1647 515 1653
rect 540 1652 577 1653
rect 430 1627 438 1647
rect 458 1627 515 1647
rect 430 1619 515 1627
rect 539 1643 577 1652
rect 539 1623 548 1643
rect 568 1623 577 1643
rect 430 1618 466 1619
rect 539 1615 577 1623
rect 643 1647 728 1653
rect 748 1652 785 1653
rect 643 1627 651 1647
rect 671 1646 728 1647
rect 671 1627 700 1646
rect 643 1626 700 1627
rect 721 1626 728 1646
rect 643 1619 728 1626
rect 747 1643 785 1652
rect 747 1623 756 1643
rect 776 1623 785 1643
rect 643 1618 679 1619
rect 747 1615 785 1623
rect 851 1647 995 1653
rect 851 1627 859 1647
rect 879 1646 967 1647
rect 879 1627 907 1646
rect 851 1625 907 1627
rect 929 1627 967 1646
rect 987 1627 995 1647
rect 929 1625 995 1627
rect 851 1619 995 1625
rect 851 1618 887 1619
rect 959 1618 995 1619
rect 1061 1652 1098 1653
rect 1061 1651 1099 1652
rect 1061 1643 1125 1651
rect 1061 1623 1070 1643
rect 1090 1629 1125 1643
rect 1145 1629 1148 1649
rect 1090 1624 1148 1629
rect 1090 1623 1125 1624
rect 327 1586 364 1615
rect 147 1540 185 1581
rect 328 1584 364 1586
rect 540 1584 577 1615
rect 328 1562 577 1584
rect 748 1583 785 1615
rect 1061 1611 1125 1623
rect 1165 1585 1192 1763
rect 1024 1583 1192 1585
rect 748 1557 1192 1583
rect 749 1540 773 1557
rect 1024 1556 1192 1557
rect 147 1522 774 1540
rect 1400 1536 1650 1560
rect 147 1516 185 1522
rect 147 1492 184 1516
rect 147 1468 182 1492
rect 145 1459 182 1468
rect 145 1441 155 1459
rect 173 1441 182 1459
rect 145 1431 182 1441
rect 1400 1465 1437 1536
rect 1552 1475 1583 1476
rect 1400 1445 1409 1465
rect 1429 1445 1437 1465
rect 1400 1435 1437 1445
rect 1496 1465 1583 1475
rect 1496 1445 1505 1465
rect 1525 1445 1583 1465
rect 1496 1436 1583 1445
rect 1496 1435 1533 1436
rect 1552 1383 1583 1436
rect 1613 1465 1650 1536
rect 1821 1541 2214 1561
rect 2234 1541 2237 1561
rect 1821 1536 2237 1541
rect 1821 1535 2162 1536
rect 1765 1475 1796 1476
rect 1613 1445 1622 1465
rect 1642 1445 1650 1465
rect 1613 1435 1650 1445
rect 1709 1468 1796 1475
rect 1709 1465 1770 1468
rect 1709 1445 1718 1465
rect 1738 1448 1770 1465
rect 1791 1448 1796 1468
rect 1738 1445 1796 1448
rect 1709 1438 1796 1445
rect 1821 1465 1858 1535
rect 2124 1534 2161 1535
rect 1973 1475 2009 1476
rect 1821 1445 1830 1465
rect 1850 1445 1858 1465
rect 1709 1436 1765 1438
rect 1709 1435 1746 1436
rect 1821 1435 1858 1445
rect 1917 1465 2065 1475
rect 2165 1472 2261 1474
rect 1917 1445 1926 1465
rect 1946 1445 2036 1465
rect 2056 1445 2065 1465
rect 1917 1436 2065 1445
rect 2123 1465 2261 1472
rect 2123 1445 2132 1465
rect 2152 1445 2261 1465
rect 2123 1436 2261 1445
rect 1917 1435 1954 1436
rect 1973 1384 2009 1436
rect 2028 1435 2065 1436
rect 2124 1435 2161 1436
rect 1444 1382 1485 1383
rect 1336 1375 1485 1382
rect 148 1367 185 1369
rect 148 1366 796 1367
rect 147 1360 796 1366
rect 147 1342 157 1360
rect 175 1346 796 1360
rect 1336 1355 1454 1375
rect 1474 1355 1485 1375
rect 1336 1347 1485 1355
rect 1552 1379 1911 1383
rect 1552 1374 1874 1379
rect 1552 1350 1665 1374
rect 1689 1355 1874 1374
rect 1898 1355 1911 1379
rect 1689 1350 1911 1355
rect 1552 1347 1911 1350
rect 1973 1347 2008 1384
rect 2076 1381 2176 1384
rect 2076 1377 2143 1381
rect 2076 1351 2088 1377
rect 2114 1355 2143 1377
rect 2169 1355 2176 1381
rect 2114 1351 2176 1355
rect 2076 1347 2176 1351
rect 175 1342 185 1346
rect 626 1345 796 1346
rect 147 1332 185 1342
rect 147 1254 182 1332
rect 759 1322 796 1345
rect 1552 1326 1583 1347
rect 1973 1326 2009 1347
rect 1395 1325 1432 1326
rect 143 1245 182 1254
rect 143 1227 153 1245
rect 171 1227 182 1245
rect 143 1221 182 1227
rect 338 1297 588 1321
rect 338 1226 375 1297
rect 490 1236 521 1237
rect 143 1217 180 1221
rect 338 1206 347 1226
rect 367 1206 375 1226
rect 338 1196 375 1206
rect 434 1226 521 1236
rect 434 1206 443 1226
rect 463 1206 521 1226
rect 434 1197 521 1206
rect 434 1196 471 1197
rect 146 1146 183 1155
rect 144 1128 155 1146
rect 173 1128 183 1146
rect 490 1144 521 1197
rect 551 1226 588 1297
rect 759 1302 1152 1322
rect 1172 1302 1175 1322
rect 759 1297 1175 1302
rect 1394 1316 1432 1325
rect 759 1296 1100 1297
rect 1394 1296 1403 1316
rect 1423 1296 1432 1316
rect 703 1236 734 1237
rect 551 1206 560 1226
rect 580 1206 588 1226
rect 551 1196 588 1206
rect 647 1229 734 1236
rect 647 1226 708 1229
rect 647 1206 656 1226
rect 676 1209 708 1226
rect 729 1209 734 1229
rect 676 1206 734 1209
rect 647 1199 734 1206
rect 759 1226 796 1296
rect 1062 1295 1099 1296
rect 1394 1288 1432 1296
rect 1498 1320 1583 1326
rect 1608 1325 1645 1326
rect 1498 1300 1506 1320
rect 1526 1300 1583 1320
rect 1498 1292 1583 1300
rect 1607 1316 1645 1325
rect 1607 1296 1616 1316
rect 1636 1296 1645 1316
rect 1498 1291 1534 1292
rect 1607 1288 1645 1296
rect 1711 1320 1796 1326
rect 1816 1325 1853 1326
rect 1711 1300 1719 1320
rect 1739 1319 1796 1320
rect 1739 1300 1768 1319
rect 1711 1299 1768 1300
rect 1789 1299 1796 1319
rect 1711 1292 1796 1299
rect 1815 1316 1853 1325
rect 1815 1296 1824 1316
rect 1844 1296 1853 1316
rect 1711 1291 1747 1292
rect 1815 1288 1853 1296
rect 1919 1320 2063 1326
rect 1919 1300 1927 1320
rect 1947 1319 2035 1320
rect 1947 1300 1980 1319
rect 2003 1300 2035 1319
rect 2055 1300 2063 1320
rect 1919 1292 2063 1300
rect 1919 1291 1955 1292
rect 2027 1291 2063 1292
rect 2129 1325 2166 1326
rect 2129 1324 2167 1325
rect 2129 1316 2193 1324
rect 2129 1296 2138 1316
rect 2158 1302 2193 1316
rect 2213 1302 2216 1322
rect 2158 1297 2216 1302
rect 2158 1296 2193 1297
rect 1395 1259 1432 1288
rect 1396 1257 1432 1259
rect 1608 1257 1645 1288
rect 911 1236 947 1237
rect 759 1206 768 1226
rect 788 1206 796 1226
rect 647 1197 703 1199
rect 647 1196 684 1197
rect 759 1196 796 1206
rect 855 1226 1003 1236
rect 1396 1235 1645 1257
rect 1816 1256 1853 1288
rect 2129 1284 2193 1296
rect 2233 1258 2260 1436
rect 2092 1256 2260 1258
rect 1816 1245 2260 1256
rect 2323 1256 2353 2257
rect 2442 2250 2479 2261
rect 4063 2250 4090 2428
rect 4130 2390 4194 2402
rect 4470 2398 4507 2430
rect 4678 2429 4927 2451
rect 4678 2398 4715 2429
rect 4891 2427 4927 2429
rect 5070 2432 5108 2473
rect 4891 2398 4928 2427
rect 4130 2389 4165 2390
rect 4107 2384 4165 2389
rect 4107 2364 4110 2384
rect 4130 2370 4165 2384
rect 4185 2370 4194 2390
rect 4130 2362 4194 2370
rect 4156 2361 4194 2362
rect 4157 2360 4194 2361
rect 4260 2394 4296 2395
rect 4368 2394 4404 2395
rect 4260 2388 4404 2394
rect 4260 2386 4326 2388
rect 4260 2366 4268 2386
rect 4288 2367 4326 2386
rect 4348 2386 4404 2388
rect 4348 2367 4376 2386
rect 4288 2366 4376 2367
rect 4396 2366 4404 2386
rect 4260 2360 4404 2366
rect 4470 2390 4508 2398
rect 4576 2394 4612 2395
rect 4470 2370 4479 2390
rect 4499 2370 4508 2390
rect 4470 2361 4508 2370
rect 4527 2387 4612 2394
rect 4527 2367 4534 2387
rect 4555 2386 4612 2387
rect 4555 2367 4584 2386
rect 4527 2366 4584 2367
rect 4604 2366 4612 2386
rect 4470 2360 4507 2361
rect 4527 2360 4612 2366
rect 4678 2390 4716 2398
rect 4789 2394 4825 2395
rect 4678 2370 4687 2390
rect 4707 2370 4716 2390
rect 4678 2361 4716 2370
rect 4740 2386 4825 2394
rect 4740 2366 4797 2386
rect 4817 2366 4825 2386
rect 4678 2360 4715 2361
rect 4740 2360 4825 2366
rect 4891 2390 4929 2398
rect 4891 2370 4900 2390
rect 4920 2370 4929 2390
rect 4891 2361 4929 2370
rect 5070 2397 5106 2432
rect 5423 2428 5458 2474
rect 6834 2472 6871 2543
rect 6986 2482 7017 2483
rect 6834 2452 6843 2472
rect 6863 2452 6871 2472
rect 6834 2442 6871 2452
rect 6930 2472 7017 2482
rect 6930 2452 6939 2472
rect 6959 2452 7017 2472
rect 6930 2443 7017 2452
rect 6930 2442 6967 2443
rect 5421 2419 5458 2428
rect 5421 2401 5431 2419
rect 5449 2401 5458 2419
rect 5070 2387 5107 2397
rect 5421 2391 5458 2401
rect 6986 2390 7017 2443
rect 7047 2472 7084 2543
rect 7255 2548 7648 2568
rect 7668 2548 7671 2568
rect 7255 2543 7671 2548
rect 7255 2542 7596 2543
rect 7199 2482 7230 2483
rect 7047 2452 7056 2472
rect 7076 2452 7084 2472
rect 7047 2442 7084 2452
rect 7143 2475 7230 2482
rect 7143 2472 7204 2475
rect 7143 2452 7152 2472
rect 7172 2455 7204 2472
rect 7225 2455 7230 2475
rect 7172 2452 7230 2455
rect 7143 2445 7230 2452
rect 7255 2472 7292 2542
rect 7558 2541 7595 2542
rect 7407 2482 7443 2483
rect 7255 2452 7264 2472
rect 7284 2452 7292 2472
rect 7143 2443 7199 2445
rect 7143 2442 7180 2443
rect 7255 2442 7292 2452
rect 7351 2472 7499 2482
rect 7599 2479 7695 2481
rect 7351 2452 7360 2472
rect 7380 2452 7470 2472
rect 7490 2452 7499 2472
rect 7351 2443 7499 2452
rect 7557 2472 7695 2479
rect 7557 2452 7566 2472
rect 7586 2452 7695 2472
rect 7557 2443 7695 2452
rect 7351 2442 7388 2443
rect 7407 2391 7443 2443
rect 7462 2442 7499 2443
rect 7558 2442 7595 2443
rect 6878 2389 6919 2390
rect 5070 2369 5080 2387
rect 5098 2369 5107 2387
rect 4891 2360 4928 2361
rect 5070 2360 5107 2369
rect 6770 2382 6919 2389
rect 6770 2362 6888 2382
rect 6908 2362 6919 2382
rect 4314 2339 4350 2360
rect 4740 2339 4771 2360
rect 6770 2354 6919 2362
rect 6986 2386 7345 2390
rect 6986 2381 7308 2386
rect 6986 2357 7099 2381
rect 7123 2362 7308 2381
rect 7332 2362 7345 2386
rect 7123 2357 7345 2362
rect 6986 2354 7345 2357
rect 7407 2354 7442 2391
rect 7510 2388 7610 2391
rect 7510 2384 7577 2388
rect 7510 2358 7522 2384
rect 7548 2362 7577 2384
rect 7603 2362 7610 2388
rect 7548 2358 7610 2362
rect 7510 2354 7610 2358
rect 4147 2335 4247 2339
rect 4147 2331 4209 2335
rect 4147 2305 4154 2331
rect 4180 2309 4209 2331
rect 4235 2309 4247 2335
rect 4180 2305 4247 2309
rect 4147 2302 4247 2305
rect 4315 2302 4350 2339
rect 4412 2336 4771 2339
rect 4412 2331 4634 2336
rect 4412 2307 4425 2331
rect 4449 2312 4634 2331
rect 4658 2312 4771 2336
rect 4449 2307 4771 2312
rect 4412 2303 4771 2307
rect 4838 2331 4987 2339
rect 6986 2333 7017 2354
rect 7407 2333 7443 2354
rect 6829 2332 6866 2333
rect 4838 2311 4849 2331
rect 4869 2311 4987 2331
rect 5424 2327 5461 2329
rect 5424 2326 6072 2327
rect 4838 2304 4987 2311
rect 5423 2320 6072 2326
rect 4838 2303 4879 2304
rect 4162 2250 4199 2251
rect 4258 2250 4295 2251
rect 4314 2250 4350 2302
rect 4369 2250 4406 2251
rect 4062 2241 4200 2250
rect 2998 2223 3029 2226
rect 2998 2197 3005 2223
rect 3024 2197 3029 2223
rect 2998 1803 3029 2197
rect 3050 2222 3218 2223
rect 3050 2219 3494 2222
rect 3050 2200 3425 2219
rect 3445 2200 3494 2219
rect 4062 2221 4171 2241
rect 4191 2221 4200 2241
rect 3050 2196 3494 2200
rect 3050 2194 3218 2196
rect 3050 2016 3077 2194
rect 3117 2156 3181 2168
rect 3457 2164 3494 2196
rect 3665 2195 3914 2217
rect 4062 2214 4200 2221
rect 4258 2241 4406 2250
rect 4258 2221 4267 2241
rect 4287 2221 4377 2241
rect 4397 2221 4406 2241
rect 4062 2212 4158 2214
rect 4258 2211 4406 2221
rect 4465 2241 4502 2251
rect 4577 2250 4614 2251
rect 4558 2248 4614 2250
rect 4465 2221 4473 2241
rect 4493 2221 4502 2241
rect 4314 2210 4350 2211
rect 3665 2164 3702 2195
rect 3878 2193 3914 2195
rect 3878 2164 3915 2193
rect 3117 2155 3152 2156
rect 3094 2150 3152 2155
rect 3094 2130 3097 2150
rect 3117 2136 3152 2150
rect 3172 2136 3181 2156
rect 3117 2128 3181 2136
rect 3143 2127 3181 2128
rect 3144 2126 3181 2127
rect 3247 2160 3283 2161
rect 3355 2160 3391 2161
rect 3247 2152 3391 2160
rect 3247 2132 3255 2152
rect 3275 2151 3363 2152
rect 3275 2132 3308 2151
rect 3247 2131 3308 2132
rect 3332 2132 3363 2151
rect 3383 2132 3391 2152
rect 3332 2131 3391 2132
rect 3247 2126 3391 2131
rect 3457 2156 3495 2164
rect 3563 2160 3599 2161
rect 3457 2136 3466 2156
rect 3486 2136 3495 2156
rect 3457 2127 3495 2136
rect 3514 2153 3599 2160
rect 3514 2133 3521 2153
rect 3542 2152 3599 2153
rect 3542 2133 3571 2152
rect 3514 2132 3571 2133
rect 3591 2132 3599 2152
rect 3457 2126 3494 2127
rect 3514 2126 3599 2132
rect 3665 2156 3703 2164
rect 3776 2160 3812 2161
rect 3665 2136 3674 2156
rect 3694 2136 3703 2156
rect 3665 2127 3703 2136
rect 3727 2152 3812 2160
rect 3727 2132 3784 2152
rect 3804 2132 3812 2152
rect 3665 2126 3702 2127
rect 3727 2126 3812 2132
rect 3878 2156 3916 2164
rect 3878 2136 3887 2156
rect 3907 2136 3916 2156
rect 4162 2151 4199 2152
rect 4465 2151 4502 2221
rect 4527 2241 4614 2248
rect 4527 2238 4585 2241
rect 4527 2218 4532 2238
rect 4553 2221 4585 2238
rect 4605 2221 4614 2241
rect 4553 2218 4614 2221
rect 4527 2211 4614 2218
rect 4673 2241 4710 2251
rect 4673 2221 4681 2241
rect 4701 2221 4710 2241
rect 4527 2210 4558 2211
rect 4161 2150 4502 2151
rect 3878 2127 3916 2136
rect 4086 2145 4502 2150
rect 3878 2126 3915 2127
rect 3301 2105 3337 2126
rect 3727 2105 3758 2126
rect 4086 2125 4089 2145
rect 4109 2125 4502 2145
rect 4673 2150 4710 2221
rect 4740 2250 4771 2303
rect 5423 2302 5433 2320
rect 5451 2306 6072 2320
rect 5451 2302 5461 2306
rect 5902 2305 6072 2306
rect 5073 2288 5110 2298
rect 5073 2270 5082 2288
rect 5100 2270 5110 2288
rect 5073 2261 5110 2270
rect 5423 2292 5461 2302
rect 4790 2250 4827 2251
rect 4740 2241 4827 2250
rect 4740 2221 4798 2241
rect 4818 2221 4827 2241
rect 4740 2211 4827 2221
rect 4886 2241 4923 2251
rect 4886 2221 4894 2241
rect 4914 2221 4923 2241
rect 4740 2210 4771 2211
rect 4886 2150 4923 2221
rect 5078 2196 5109 2261
rect 5423 2214 5458 2292
rect 6035 2282 6072 2305
rect 6828 2323 6866 2332
rect 6828 2303 6837 2323
rect 6857 2303 6866 2323
rect 6828 2295 6866 2303
rect 6932 2327 7017 2333
rect 7042 2332 7079 2333
rect 6932 2307 6940 2327
rect 6960 2307 7017 2327
rect 6932 2299 7017 2307
rect 7041 2323 7079 2332
rect 7041 2303 7050 2323
rect 7070 2303 7079 2323
rect 6932 2298 6968 2299
rect 7041 2295 7079 2303
rect 7145 2327 7230 2333
rect 7250 2332 7287 2333
rect 7145 2307 7153 2327
rect 7173 2326 7230 2327
rect 7173 2307 7202 2326
rect 7145 2306 7202 2307
rect 7223 2306 7230 2326
rect 7145 2299 7230 2306
rect 7249 2323 7287 2332
rect 7249 2303 7258 2323
rect 7278 2303 7287 2323
rect 7145 2298 7181 2299
rect 7249 2295 7287 2303
rect 7353 2327 7497 2333
rect 7353 2307 7361 2327
rect 7381 2308 7417 2327
rect 7440 2308 7469 2327
rect 7381 2307 7469 2308
rect 7489 2307 7497 2327
rect 7353 2299 7497 2307
rect 7353 2298 7389 2299
rect 7461 2298 7497 2299
rect 7563 2332 7600 2333
rect 7563 2331 7601 2332
rect 7563 2323 7627 2331
rect 7563 2303 7572 2323
rect 7592 2309 7627 2323
rect 7647 2309 7650 2329
rect 7592 2304 7650 2309
rect 7592 2303 7627 2304
rect 5419 2205 5458 2214
rect 5077 2186 5114 2196
rect 5077 2184 5087 2186
rect 5011 2182 5087 2184
rect 4673 2126 4923 2150
rect 5008 2168 5087 2182
rect 5105 2168 5114 2186
rect 5419 2187 5429 2205
rect 5447 2187 5458 2205
rect 5419 2181 5458 2187
rect 5614 2257 5864 2281
rect 5614 2186 5651 2257
rect 5766 2196 5797 2197
rect 5419 2177 5456 2181
rect 5008 2165 5114 2168
rect 4480 2106 4501 2125
rect 5008 2106 5034 2165
rect 5077 2159 5114 2165
rect 5614 2166 5623 2186
rect 5643 2166 5651 2186
rect 5614 2156 5651 2166
rect 5710 2186 5797 2196
rect 5710 2166 5719 2186
rect 5739 2166 5797 2186
rect 5710 2157 5797 2166
rect 5710 2156 5747 2157
rect 5422 2106 5459 2115
rect 3134 2101 3234 2105
rect 3134 2097 3196 2101
rect 3134 2071 3141 2097
rect 3167 2075 3196 2097
rect 3222 2075 3234 2101
rect 3167 2071 3234 2075
rect 3134 2068 3234 2071
rect 3302 2068 3337 2105
rect 3399 2102 3758 2105
rect 3399 2097 3621 2102
rect 3399 2073 3412 2097
rect 3436 2078 3621 2097
rect 3645 2078 3758 2102
rect 3436 2073 3758 2078
rect 3399 2069 3758 2073
rect 3825 2097 3974 2105
rect 3825 2077 3836 2097
rect 3856 2077 3974 2097
rect 4480 2088 5034 2106
rect 5080 2095 5117 2097
rect 5008 2087 5034 2088
rect 5077 2087 5117 2095
rect 3825 2070 3974 2077
rect 5077 2075 5089 2087
rect 5068 2070 5089 2075
rect 3825 2069 3866 2070
rect 4484 2069 5089 2070
rect 5107 2069 5117 2087
rect 3149 2016 3186 2017
rect 3245 2016 3282 2017
rect 3301 2016 3337 2068
rect 3356 2016 3393 2017
rect 3049 2007 3187 2016
rect 3049 1987 3158 2007
rect 3178 1987 3187 2007
rect 3049 1980 3187 1987
rect 3245 2007 3393 2016
rect 3245 1987 3254 2007
rect 3274 1987 3364 2007
rect 3384 1987 3393 2007
rect 3049 1978 3145 1980
rect 3245 1977 3393 1987
rect 3452 2007 3489 2017
rect 3564 2016 3601 2017
rect 3545 2014 3601 2016
rect 3452 1987 3460 2007
rect 3480 1987 3489 2007
rect 3301 1976 3337 1977
rect 3149 1917 3186 1918
rect 3452 1917 3489 1987
rect 3514 2007 3601 2014
rect 3514 2004 3572 2007
rect 3514 1984 3519 2004
rect 3540 1987 3572 2004
rect 3592 1987 3601 2007
rect 3540 1984 3601 1987
rect 3514 1977 3601 1984
rect 3660 2007 3697 2017
rect 3660 1987 3668 2007
rect 3688 1987 3697 2007
rect 3514 1976 3545 1977
rect 3148 1916 3489 1917
rect 3073 1911 3489 1916
rect 3073 1891 3076 1911
rect 3096 1891 3489 1911
rect 3660 1916 3697 1987
rect 3727 2016 3758 2069
rect 4484 2060 5117 2069
rect 5420 2088 5431 2106
rect 5449 2088 5459 2106
rect 5766 2104 5797 2157
rect 5827 2186 5864 2257
rect 6035 2262 6428 2282
rect 6448 2262 6451 2282
rect 6829 2266 6866 2295
rect 6035 2257 6451 2262
rect 6830 2264 6866 2266
rect 7042 2264 7079 2295
rect 6035 2256 6376 2257
rect 5979 2196 6010 2197
rect 5827 2166 5836 2186
rect 5856 2166 5864 2186
rect 5827 2156 5864 2166
rect 5923 2189 6010 2196
rect 5923 2186 5984 2189
rect 5923 2166 5932 2186
rect 5952 2169 5984 2186
rect 6005 2169 6010 2189
rect 5952 2166 6010 2169
rect 5923 2159 6010 2166
rect 6035 2186 6072 2256
rect 6338 2255 6375 2256
rect 6830 2242 7079 2264
rect 7250 2263 7287 2295
rect 7563 2291 7627 2303
rect 7667 2265 7694 2443
rect 7722 2330 7760 4161
rect 8267 4136 8274 4162
rect 8293 4136 8298 4162
rect 8174 3743 8203 3745
rect 8174 3738 8206 3743
rect 8174 3720 8181 3738
rect 8201 3720 8206 3738
rect 8267 3742 8298 4136
rect 8319 4161 8487 4162
rect 8319 4158 8763 4161
rect 8319 4139 8694 4158
rect 8714 4139 8763 4158
rect 9331 4160 9440 4180
rect 9460 4160 9469 4180
rect 8319 4135 8763 4139
rect 8319 4133 8487 4135
rect 8319 3955 8346 4133
rect 8386 4095 8450 4107
rect 8726 4103 8763 4135
rect 8934 4134 9183 4156
rect 9331 4153 9469 4160
rect 9527 4180 9675 4189
rect 9527 4160 9536 4180
rect 9556 4160 9646 4180
rect 9666 4160 9675 4180
rect 9331 4151 9427 4153
rect 9527 4150 9675 4160
rect 9734 4180 9771 4190
rect 9846 4189 9883 4190
rect 9827 4187 9883 4189
rect 9734 4160 9742 4180
rect 9762 4160 9771 4180
rect 9583 4149 9619 4150
rect 8934 4103 8971 4134
rect 9147 4132 9183 4134
rect 9147 4103 9184 4132
rect 8386 4094 8421 4095
rect 8363 4089 8421 4094
rect 8363 4069 8366 4089
rect 8386 4075 8421 4089
rect 8441 4075 8450 4095
rect 8386 4067 8450 4075
rect 8412 4066 8450 4067
rect 8413 4065 8450 4066
rect 8516 4099 8552 4100
rect 8624 4099 8660 4100
rect 8516 4091 8660 4099
rect 8516 4071 8524 4091
rect 8544 4090 8632 4091
rect 8544 4071 8577 4090
rect 8516 4070 8577 4071
rect 8601 4071 8632 4090
rect 8652 4071 8660 4091
rect 8601 4070 8660 4071
rect 8516 4065 8660 4070
rect 8726 4095 8764 4103
rect 8832 4099 8868 4100
rect 8726 4075 8735 4095
rect 8755 4075 8764 4095
rect 8726 4066 8764 4075
rect 8783 4092 8868 4099
rect 8783 4072 8790 4092
rect 8811 4091 8868 4092
rect 8811 4072 8840 4091
rect 8783 4071 8840 4072
rect 8860 4071 8868 4091
rect 8726 4065 8763 4066
rect 8783 4065 8868 4071
rect 8934 4095 8972 4103
rect 9045 4099 9081 4100
rect 8934 4075 8943 4095
rect 8963 4075 8972 4095
rect 8934 4066 8972 4075
rect 8996 4091 9081 4099
rect 8996 4071 9053 4091
rect 9073 4071 9081 4091
rect 8934 4065 8971 4066
rect 8996 4065 9081 4071
rect 9147 4095 9185 4103
rect 9147 4075 9156 4095
rect 9176 4075 9185 4095
rect 9431 4090 9468 4091
rect 9734 4090 9771 4160
rect 9796 4180 9883 4187
rect 9796 4177 9854 4180
rect 9796 4157 9801 4177
rect 9822 4160 9854 4177
rect 9874 4160 9883 4180
rect 9822 4157 9883 4160
rect 9796 4150 9883 4157
rect 9942 4180 9979 4190
rect 9942 4160 9950 4180
rect 9970 4160 9979 4180
rect 9796 4149 9827 4150
rect 9430 4089 9771 4090
rect 9147 4066 9185 4075
rect 9355 4084 9771 4089
rect 9147 4065 9184 4066
rect 8570 4044 8606 4065
rect 8996 4044 9027 4065
rect 9355 4064 9358 4084
rect 9378 4064 9771 4084
rect 9942 4089 9979 4160
rect 10009 4189 10040 4242
rect 10342 4227 10379 4237
rect 10342 4209 10351 4227
rect 10369 4209 10379 4227
rect 10342 4200 10379 4209
rect 10791 4203 10826 4281
rect 11403 4271 11440 4294
rect 12441 4287 12472 4308
rect 12862 4287 12898 4308
rect 12284 4286 12321 4287
rect 12283 4277 12321 4286
rect 10059 4189 10096 4190
rect 10009 4180 10096 4189
rect 10009 4160 10067 4180
rect 10087 4160 10096 4180
rect 10009 4150 10096 4160
rect 10155 4180 10192 4190
rect 10155 4160 10163 4180
rect 10183 4160 10192 4180
rect 10009 4149 10040 4150
rect 10155 4089 10192 4160
rect 10347 4135 10378 4200
rect 10787 4194 10826 4203
rect 10787 4176 10797 4194
rect 10815 4176 10826 4194
rect 10787 4170 10826 4176
rect 10982 4246 11232 4270
rect 10982 4175 11019 4246
rect 11134 4185 11165 4186
rect 10787 4166 10824 4170
rect 10982 4155 10991 4175
rect 11011 4155 11019 4175
rect 10982 4145 11019 4155
rect 11078 4175 11165 4185
rect 11078 4155 11087 4175
rect 11107 4155 11165 4175
rect 11078 4146 11165 4155
rect 11078 4145 11115 4146
rect 10346 4125 10383 4135
rect 10346 4123 10356 4125
rect 10280 4121 10356 4123
rect 9942 4065 10192 4089
rect 10277 4107 10356 4121
rect 10374 4107 10383 4125
rect 10277 4104 10383 4107
rect 9749 4045 9770 4064
rect 10277 4045 10303 4104
rect 10346 4098 10383 4104
rect 10790 4095 10827 4104
rect 8403 4040 8503 4044
rect 8403 4036 8465 4040
rect 8403 4010 8410 4036
rect 8436 4014 8465 4036
rect 8491 4014 8503 4040
rect 8436 4010 8503 4014
rect 8403 4007 8503 4010
rect 8571 4007 8606 4044
rect 8668 4041 9027 4044
rect 8668 4036 8890 4041
rect 8668 4012 8681 4036
rect 8705 4017 8890 4036
rect 8914 4017 9027 4041
rect 8705 4012 9027 4017
rect 8668 4008 9027 4012
rect 9094 4036 9243 4044
rect 9094 4016 9105 4036
rect 9125 4016 9243 4036
rect 9749 4027 10303 4045
rect 10788 4077 10799 4095
rect 10817 4077 10827 4095
rect 11134 4093 11165 4146
rect 11195 4175 11232 4246
rect 11403 4251 11796 4271
rect 11816 4251 11819 4271
rect 11403 4246 11819 4251
rect 12283 4257 12292 4277
rect 12312 4257 12321 4277
rect 12283 4249 12321 4257
rect 12387 4281 12472 4287
rect 12497 4286 12534 4287
rect 12387 4261 12395 4281
rect 12415 4261 12472 4281
rect 12387 4253 12472 4261
rect 12496 4277 12534 4286
rect 12496 4257 12505 4277
rect 12525 4257 12534 4277
rect 12387 4252 12423 4253
rect 12496 4249 12534 4257
rect 12600 4281 12685 4287
rect 12705 4286 12742 4287
rect 12600 4261 12608 4281
rect 12628 4280 12685 4281
rect 12628 4261 12657 4280
rect 12600 4260 12657 4261
rect 12678 4260 12685 4280
rect 12600 4253 12685 4260
rect 12704 4277 12742 4286
rect 12704 4257 12713 4277
rect 12733 4257 12742 4277
rect 12600 4252 12636 4253
rect 12704 4249 12742 4257
rect 12808 4282 12952 4287
rect 12808 4281 12872 4282
rect 12808 4261 12816 4281
rect 12836 4263 12872 4281
rect 12898 4281 12952 4282
rect 12898 4263 12924 4281
rect 12836 4261 12924 4263
rect 12944 4261 12952 4281
rect 12808 4253 12952 4261
rect 12808 4252 12844 4253
rect 12916 4252 12952 4253
rect 13018 4286 13055 4287
rect 13018 4285 13056 4286
rect 13018 4277 13082 4285
rect 13018 4257 13027 4277
rect 13047 4263 13082 4277
rect 13102 4263 13105 4283
rect 13047 4258 13105 4263
rect 13047 4257 13082 4258
rect 11403 4245 11744 4246
rect 11347 4185 11378 4186
rect 11195 4155 11204 4175
rect 11224 4155 11232 4175
rect 11195 4145 11232 4155
rect 11291 4178 11378 4185
rect 11291 4175 11352 4178
rect 11291 4155 11300 4175
rect 11320 4158 11352 4175
rect 11373 4158 11378 4178
rect 11320 4155 11378 4158
rect 11291 4148 11378 4155
rect 11403 4175 11440 4245
rect 11706 4244 11743 4245
rect 12284 4220 12321 4249
rect 12285 4218 12321 4220
rect 12497 4218 12534 4249
rect 12285 4196 12534 4218
rect 12705 4217 12742 4249
rect 13018 4245 13082 4257
rect 13122 4222 13149 4397
rect 13102 4219 13149 4222
rect 12981 4217 13149 4219
rect 14712 4396 14880 4398
rect 14712 4218 14739 4396
rect 14779 4358 14843 4370
rect 15119 4366 15156 4398
rect 15327 4397 15576 4419
rect 15327 4366 15364 4397
rect 15540 4395 15576 4397
rect 15719 4400 15757 4441
rect 16072 4439 16112 4444
rect 15540 4366 15577 4395
rect 14779 4357 14814 4358
rect 14756 4352 14814 4357
rect 14756 4332 14759 4352
rect 14779 4338 14814 4352
rect 14834 4338 14843 4358
rect 14779 4330 14843 4338
rect 14805 4329 14843 4330
rect 14806 4328 14843 4329
rect 14909 4362 14945 4363
rect 15017 4362 15053 4363
rect 14909 4356 15053 4362
rect 14909 4354 14975 4356
rect 14909 4334 14917 4354
rect 14937 4335 14975 4354
rect 14997 4354 15053 4356
rect 14997 4335 15025 4354
rect 14937 4334 15025 4335
rect 15045 4334 15053 4354
rect 14909 4328 15053 4334
rect 15119 4358 15157 4366
rect 15225 4362 15261 4363
rect 15119 4338 15128 4358
rect 15148 4338 15157 4358
rect 15119 4329 15157 4338
rect 15176 4355 15261 4362
rect 15176 4335 15183 4355
rect 15204 4354 15261 4355
rect 15204 4335 15233 4354
rect 15176 4334 15233 4335
rect 15253 4334 15261 4354
rect 15119 4328 15156 4329
rect 15176 4328 15261 4334
rect 15327 4358 15365 4366
rect 15438 4362 15474 4363
rect 15327 4338 15336 4358
rect 15356 4338 15365 4358
rect 15327 4329 15365 4338
rect 15389 4354 15474 4362
rect 15389 4334 15446 4354
rect 15466 4334 15474 4354
rect 15327 4328 15364 4329
rect 15389 4328 15474 4334
rect 15540 4358 15578 4366
rect 15540 4338 15549 4358
rect 15569 4338 15578 4358
rect 15540 4329 15578 4338
rect 15719 4365 15755 4400
rect 16072 4396 16107 4439
rect 16070 4387 16107 4396
rect 16070 4369 16080 4387
rect 16098 4369 16107 4387
rect 17570 4405 17607 4476
rect 17722 4415 17753 4416
rect 17570 4385 17579 4405
rect 17599 4385 17607 4405
rect 17570 4375 17607 4385
rect 17666 4405 17753 4415
rect 17666 4385 17675 4405
rect 17695 4385 17753 4405
rect 17666 4376 17753 4385
rect 17666 4375 17703 4376
rect 15719 4355 15756 4365
rect 16070 4359 16107 4369
rect 15719 4337 15729 4355
rect 15747 4337 15756 4355
rect 15540 4328 15577 4329
rect 15719 4328 15756 4337
rect 14963 4307 14999 4328
rect 15389 4307 15420 4328
rect 17722 4323 17753 4376
rect 17783 4405 17820 4476
rect 17991 4481 18384 4501
rect 18404 4481 18407 4501
rect 17991 4476 18407 4481
rect 18681 4498 18819 4507
rect 18681 4478 18790 4498
rect 18810 4478 18819 4498
rect 17991 4475 18332 4476
rect 17935 4415 17966 4416
rect 17783 4385 17792 4405
rect 17812 4385 17820 4405
rect 17783 4375 17820 4385
rect 17879 4408 17966 4415
rect 17879 4405 17940 4408
rect 17879 4385 17888 4405
rect 17908 4388 17940 4405
rect 17961 4388 17966 4408
rect 17908 4385 17966 4388
rect 17879 4378 17966 4385
rect 17991 4405 18028 4475
rect 18294 4474 18331 4475
rect 18681 4471 18819 4478
rect 18877 4498 19025 4507
rect 18877 4478 18886 4498
rect 18906 4478 18996 4498
rect 19016 4478 19025 4498
rect 18681 4469 18777 4471
rect 18877 4468 19025 4478
rect 19084 4498 19121 4508
rect 19196 4507 19233 4508
rect 19177 4505 19233 4507
rect 19084 4478 19092 4498
rect 19112 4478 19121 4498
rect 18933 4467 18969 4468
rect 18143 4415 18179 4416
rect 17991 4385 18000 4405
rect 18020 4385 18028 4405
rect 17879 4376 17935 4378
rect 17879 4375 17916 4376
rect 17991 4375 18028 4385
rect 18087 4405 18235 4415
rect 18335 4412 18431 4414
rect 18087 4385 18096 4405
rect 18116 4385 18206 4405
rect 18226 4385 18235 4405
rect 18087 4376 18235 4385
rect 18293 4405 18431 4412
rect 18781 4408 18818 4409
rect 19084 4408 19121 4478
rect 19146 4498 19233 4505
rect 19146 4495 19204 4498
rect 19146 4475 19151 4495
rect 19172 4478 19204 4495
rect 19224 4478 19233 4498
rect 19172 4475 19233 4478
rect 19146 4468 19233 4475
rect 19292 4498 19329 4508
rect 19292 4478 19300 4498
rect 19320 4478 19329 4498
rect 19146 4467 19177 4468
rect 18780 4407 19121 4408
rect 18293 4385 18302 4405
rect 18322 4385 18431 4405
rect 18293 4376 18431 4385
rect 18705 4402 19121 4407
rect 18705 4382 18708 4402
rect 18728 4382 19121 4402
rect 19292 4407 19329 4478
rect 19359 4507 19390 4560
rect 21005 4514 21042 4524
rect 19409 4507 19446 4508
rect 19359 4498 19446 4507
rect 19359 4478 19417 4498
rect 19437 4478 19446 4498
rect 19359 4468 19446 4478
rect 19505 4498 19542 4508
rect 19505 4478 19513 4498
rect 19533 4478 19542 4498
rect 19359 4467 19390 4468
rect 19505 4407 19542 4478
rect 21005 4496 21014 4514
rect 21032 4496 21042 4514
rect 21005 4487 21042 4496
rect 21005 4444 21040 4487
rect 21000 4439 21040 4444
rect 21000 4438 21038 4439
rect 20411 4420 21038 4438
rect 19292 4383 19542 4407
rect 19993 4403 20161 4404
rect 20412 4403 20436 4420
rect 19993 4377 20437 4403
rect 18087 4375 18124 4376
rect 18143 4324 18179 4376
rect 18198 4375 18235 4376
rect 18294 4375 18331 4376
rect 17614 4322 17655 4323
rect 17506 4315 17655 4322
rect 14796 4303 14896 4307
rect 14796 4299 14858 4303
rect 14796 4273 14803 4299
rect 14829 4277 14858 4299
rect 14884 4277 14896 4303
rect 14829 4273 14896 4277
rect 14796 4270 14896 4273
rect 14964 4270 14999 4307
rect 15061 4304 15420 4307
rect 15061 4299 15283 4304
rect 15061 4275 15074 4299
rect 15098 4280 15283 4299
rect 15307 4280 15420 4304
rect 15098 4275 15420 4280
rect 15061 4271 15420 4275
rect 15487 4299 15636 4307
rect 15487 4279 15498 4299
rect 15518 4279 15636 4299
rect 16073 4295 16110 4297
rect 17506 4295 17624 4315
rect 17644 4295 17655 4315
rect 16073 4294 16721 4295
rect 15487 4272 15636 4279
rect 16072 4288 16721 4294
rect 15487 4271 15528 4272
rect 14811 4218 14848 4219
rect 14907 4218 14944 4219
rect 14963 4218 14999 4270
rect 15018 4218 15055 4219
rect 12705 4191 13149 4217
rect 14711 4209 14849 4218
rect 12981 4190 13149 4191
rect 13647 4191 13678 4194
rect 11555 4185 11591 4186
rect 11403 4155 11412 4175
rect 11432 4155 11440 4175
rect 11291 4146 11347 4148
rect 11291 4145 11328 4146
rect 11403 4145 11440 4155
rect 11499 4175 11647 4185
rect 11747 4182 11843 4184
rect 11499 4155 11508 4175
rect 11528 4155 11618 4175
rect 11638 4155 11647 4175
rect 11499 4146 11647 4155
rect 11705 4175 11843 4182
rect 11705 4155 11714 4175
rect 11734 4155 11843 4175
rect 11705 4146 11843 4155
rect 11499 4145 11536 4146
rect 11555 4094 11591 4146
rect 11610 4145 11647 4146
rect 11706 4145 11743 4146
rect 11026 4092 11067 4093
rect 10349 4034 10386 4036
rect 10277 4026 10303 4027
rect 10346 4026 10386 4034
rect 9094 4009 9243 4016
rect 10346 4014 10358 4026
rect 10337 4009 10358 4014
rect 9094 4008 9135 4009
rect 9753 4008 10358 4009
rect 10376 4008 10386 4026
rect 8418 3955 8455 3956
rect 8514 3955 8551 3956
rect 8570 3955 8606 4007
rect 8625 3955 8662 3956
rect 8318 3946 8456 3955
rect 8318 3926 8427 3946
rect 8447 3926 8456 3946
rect 8318 3919 8456 3926
rect 8514 3946 8662 3955
rect 8514 3926 8523 3946
rect 8543 3926 8633 3946
rect 8653 3926 8662 3946
rect 8318 3917 8414 3919
rect 8514 3916 8662 3926
rect 8721 3946 8758 3956
rect 8833 3955 8870 3956
rect 8814 3953 8870 3955
rect 8721 3926 8729 3946
rect 8749 3926 8758 3946
rect 8570 3915 8606 3916
rect 8418 3856 8455 3857
rect 8721 3856 8758 3926
rect 8783 3946 8870 3953
rect 8783 3943 8841 3946
rect 8783 3923 8788 3943
rect 8809 3926 8841 3943
rect 8861 3926 8870 3946
rect 8809 3923 8870 3926
rect 8783 3916 8870 3923
rect 8929 3946 8966 3956
rect 8929 3926 8937 3946
rect 8957 3926 8966 3946
rect 8783 3915 8814 3916
rect 8417 3855 8758 3856
rect 8342 3850 8758 3855
rect 8342 3830 8345 3850
rect 8365 3830 8758 3850
rect 8929 3855 8966 3926
rect 8996 3955 9027 4008
rect 9753 3999 10386 4008
rect 9753 3992 10385 3999
rect 9753 3990 9815 3992
rect 9331 3980 9499 3981
rect 9753 3980 9775 3990
rect 9046 3955 9083 3956
rect 8996 3946 9083 3955
rect 8996 3926 9054 3946
rect 9074 3926 9083 3946
rect 8996 3916 9083 3926
rect 9142 3946 9179 3956
rect 9142 3926 9150 3946
rect 9170 3926 9179 3946
rect 8996 3915 9027 3916
rect 9142 3855 9179 3926
rect 8929 3831 9179 3855
rect 9331 3954 9775 3980
rect 9331 3952 9499 3954
rect 9331 3774 9358 3952
rect 9398 3914 9462 3926
rect 9738 3922 9775 3954
rect 9946 3953 10195 3975
rect 9946 3922 9983 3953
rect 10159 3951 10195 3953
rect 10159 3922 10196 3951
rect 9398 3913 9433 3914
rect 9375 3908 9433 3913
rect 9375 3888 9378 3908
rect 9398 3894 9433 3908
rect 9453 3894 9462 3914
rect 9398 3886 9462 3894
rect 9424 3885 9462 3886
rect 9425 3884 9462 3885
rect 9528 3918 9564 3919
rect 9636 3918 9672 3919
rect 9528 3910 9672 3918
rect 9528 3890 9536 3910
rect 9556 3890 9585 3910
rect 9528 3889 9585 3890
rect 9607 3890 9644 3910
rect 9664 3890 9672 3910
rect 9607 3889 9672 3890
rect 9528 3884 9672 3889
rect 9738 3914 9776 3922
rect 9844 3918 9880 3919
rect 9738 3894 9747 3914
rect 9767 3894 9776 3914
rect 9738 3885 9776 3894
rect 9795 3911 9880 3918
rect 9795 3891 9802 3911
rect 9823 3910 9880 3911
rect 9823 3891 9852 3910
rect 9795 3890 9852 3891
rect 9872 3890 9880 3910
rect 9738 3884 9775 3885
rect 9795 3884 9880 3890
rect 9946 3914 9984 3922
rect 10057 3918 10093 3919
rect 9946 3894 9955 3914
rect 9975 3894 9984 3914
rect 9946 3885 9984 3894
rect 10008 3910 10093 3918
rect 10008 3890 10065 3910
rect 10085 3890 10093 3910
rect 9946 3884 9983 3885
rect 10008 3884 10093 3890
rect 10159 3914 10197 3922
rect 10159 3894 10168 3914
rect 10188 3894 10197 3914
rect 10159 3885 10197 3894
rect 10159 3884 10196 3885
rect 9582 3863 9618 3884
rect 10008 3863 10039 3884
rect 9415 3859 9515 3863
rect 9415 3855 9477 3859
rect 9415 3829 9422 3855
rect 9448 3833 9477 3855
rect 9503 3833 9515 3859
rect 9448 3829 9515 3833
rect 9415 3826 9515 3829
rect 9583 3826 9618 3863
rect 9680 3860 10039 3863
rect 9680 3855 9902 3860
rect 9680 3831 9693 3855
rect 9717 3836 9902 3855
rect 9926 3836 10039 3860
rect 9717 3831 10039 3836
rect 9680 3827 10039 3831
rect 10106 3855 10255 3863
rect 10106 3835 10117 3855
rect 10137 3835 10255 3855
rect 10106 3828 10255 3835
rect 10346 3843 10385 3992
rect 10788 3928 10827 4077
rect 10918 4085 11067 4092
rect 10918 4065 11036 4085
rect 11056 4065 11067 4085
rect 10918 4057 11067 4065
rect 11134 4089 11493 4093
rect 11134 4084 11456 4089
rect 11134 4060 11247 4084
rect 11271 4065 11456 4084
rect 11480 4065 11493 4089
rect 11271 4060 11493 4065
rect 11134 4057 11493 4060
rect 11555 4057 11590 4094
rect 11658 4091 11758 4094
rect 11658 4087 11725 4091
rect 11658 4061 11670 4087
rect 11696 4065 11725 4087
rect 11751 4065 11758 4091
rect 11696 4061 11758 4065
rect 11658 4057 11758 4061
rect 11134 4036 11165 4057
rect 11555 4036 11591 4057
rect 10977 4035 11014 4036
rect 10976 4026 11014 4035
rect 10976 4006 10985 4026
rect 11005 4006 11014 4026
rect 10976 3998 11014 4006
rect 11080 4030 11165 4036
rect 11190 4035 11227 4036
rect 11080 4010 11088 4030
rect 11108 4010 11165 4030
rect 11080 4002 11165 4010
rect 11189 4026 11227 4035
rect 11189 4006 11198 4026
rect 11218 4006 11227 4026
rect 11080 4001 11116 4002
rect 11189 3998 11227 4006
rect 11293 4030 11378 4036
rect 11398 4035 11435 4036
rect 11293 4010 11301 4030
rect 11321 4029 11378 4030
rect 11321 4010 11350 4029
rect 11293 4009 11350 4010
rect 11371 4009 11378 4029
rect 11293 4002 11378 4009
rect 11397 4026 11435 4035
rect 11397 4006 11406 4026
rect 11426 4006 11435 4026
rect 11293 4001 11329 4002
rect 11397 3998 11435 4006
rect 11501 4031 11645 4036
rect 11501 4030 11566 4031
rect 11501 4010 11509 4030
rect 11529 4010 11566 4030
rect 11588 4030 11645 4031
rect 11588 4010 11617 4030
rect 11637 4010 11645 4030
rect 11501 4002 11645 4010
rect 11501 4001 11537 4002
rect 11609 4001 11645 4002
rect 11711 4035 11748 4036
rect 11711 4034 11749 4035
rect 11711 4026 11775 4034
rect 11711 4006 11720 4026
rect 11740 4012 11775 4026
rect 11795 4012 11798 4032
rect 11740 4007 11798 4012
rect 11740 4006 11775 4007
rect 10977 3969 11014 3998
rect 10978 3967 11014 3969
rect 11190 3967 11227 3998
rect 10978 3945 11227 3967
rect 11398 3966 11435 3998
rect 11711 3994 11775 4006
rect 11815 3968 11842 4146
rect 11674 3966 11842 3968
rect 11398 3940 11842 3966
rect 11994 4065 12244 4089
rect 11994 3994 12031 4065
rect 12146 4004 12177 4005
rect 11994 3974 12003 3994
rect 12023 3974 12031 3994
rect 11994 3964 12031 3974
rect 12090 3994 12177 4004
rect 12090 3974 12099 3994
rect 12119 3974 12177 3994
rect 12090 3965 12177 3974
rect 12090 3964 12127 3965
rect 11398 3930 11420 3940
rect 11674 3939 11842 3940
rect 11358 3928 11420 3930
rect 10788 3921 11420 3928
rect 10787 3912 11420 3921
rect 12146 3912 12177 3965
rect 12207 3994 12244 4065
rect 12415 4070 12808 4090
rect 12828 4070 12831 4090
rect 12415 4065 12831 4070
rect 12415 4064 12756 4065
rect 12359 4004 12390 4005
rect 12207 3974 12216 3994
rect 12236 3974 12244 3994
rect 12207 3964 12244 3974
rect 12303 3997 12390 4004
rect 12303 3994 12364 3997
rect 12303 3974 12312 3994
rect 12332 3977 12364 3994
rect 12385 3977 12390 3997
rect 12332 3974 12390 3977
rect 12303 3967 12390 3974
rect 12415 3994 12452 4064
rect 12718 4063 12755 4064
rect 12567 4004 12603 4005
rect 12415 3974 12424 3994
rect 12444 3974 12452 3994
rect 12303 3965 12359 3967
rect 12303 3964 12340 3965
rect 12415 3964 12452 3974
rect 12511 3994 12659 4004
rect 12759 4001 12855 4003
rect 12511 3974 12520 3994
rect 12540 3974 12630 3994
rect 12650 3974 12659 3994
rect 12511 3965 12659 3974
rect 12717 3994 12855 4001
rect 12717 3974 12726 3994
rect 12746 3974 12855 3994
rect 12717 3965 12855 3974
rect 12511 3964 12548 3965
rect 12567 3913 12603 3965
rect 12622 3964 12659 3965
rect 12718 3964 12755 3965
rect 10787 3894 10797 3912
rect 10815 3911 11420 3912
rect 12038 3911 12079 3912
rect 10815 3906 10836 3911
rect 10815 3894 10827 3906
rect 11930 3904 12079 3911
rect 10787 3886 10827 3894
rect 10870 3893 10896 3894
rect 10787 3884 10824 3886
rect 10106 3827 10147 3828
rect 9430 3774 9467 3775
rect 9526 3774 9563 3775
rect 9582 3774 9618 3826
rect 9637 3774 9674 3775
rect 9330 3765 9468 3774
rect 9330 3745 9439 3765
rect 9459 3745 9468 3765
rect 8267 3741 8437 3742
rect 8267 3726 8713 3741
rect 9330 3738 9468 3745
rect 9526 3765 9674 3774
rect 9526 3745 9535 3765
rect 9555 3745 9645 3765
rect 9665 3745 9674 3765
rect 9330 3736 9426 3738
rect 8174 3715 8206 3720
rect 8176 2714 8206 3715
rect 8269 3715 8713 3726
rect 8269 3713 8437 3715
rect 8269 3535 8296 3713
rect 8336 3675 8400 3687
rect 8676 3683 8713 3715
rect 8884 3714 9133 3736
rect 9526 3735 9674 3745
rect 9733 3765 9770 3775
rect 9845 3774 9882 3775
rect 9826 3772 9882 3774
rect 9733 3745 9741 3765
rect 9761 3745 9770 3765
rect 9582 3734 9618 3735
rect 8884 3683 8921 3714
rect 9097 3712 9133 3714
rect 9097 3683 9134 3712
rect 8336 3674 8371 3675
rect 8313 3669 8371 3674
rect 8313 3649 8316 3669
rect 8336 3655 8371 3669
rect 8391 3655 8400 3675
rect 8336 3647 8400 3655
rect 8362 3646 8400 3647
rect 8363 3645 8400 3646
rect 8466 3679 8502 3680
rect 8574 3679 8610 3680
rect 8466 3671 8610 3679
rect 8466 3651 8474 3671
rect 8494 3652 8526 3671
rect 8549 3652 8582 3671
rect 8494 3651 8582 3652
rect 8602 3651 8610 3671
rect 8466 3645 8610 3651
rect 8676 3675 8714 3683
rect 8782 3679 8818 3680
rect 8676 3655 8685 3675
rect 8705 3655 8714 3675
rect 8676 3646 8714 3655
rect 8733 3672 8818 3679
rect 8733 3652 8740 3672
rect 8761 3671 8818 3672
rect 8761 3652 8790 3671
rect 8733 3651 8790 3652
rect 8810 3651 8818 3671
rect 8676 3645 8713 3646
rect 8733 3645 8818 3651
rect 8884 3675 8922 3683
rect 8995 3679 9031 3680
rect 8884 3655 8893 3675
rect 8913 3655 8922 3675
rect 8884 3646 8922 3655
rect 8946 3671 9031 3679
rect 8946 3651 9003 3671
rect 9023 3651 9031 3671
rect 8884 3645 8921 3646
rect 8946 3645 9031 3651
rect 9097 3675 9135 3683
rect 9430 3675 9467 3676
rect 9733 3675 9770 3745
rect 9795 3765 9882 3772
rect 9795 3762 9853 3765
rect 9795 3742 9800 3762
rect 9821 3745 9853 3762
rect 9873 3745 9882 3765
rect 9821 3742 9882 3745
rect 9795 3735 9882 3742
rect 9941 3765 9978 3775
rect 9941 3745 9949 3765
rect 9969 3745 9978 3765
rect 9795 3734 9826 3735
rect 9097 3655 9106 3675
rect 9126 3655 9135 3675
rect 9429 3674 9770 3675
rect 9097 3646 9135 3655
rect 9354 3669 9770 3674
rect 9354 3649 9357 3669
rect 9377 3649 9770 3669
rect 9941 3674 9978 3745
rect 10008 3774 10039 3827
rect 10346 3825 10356 3843
rect 10374 3825 10385 3843
rect 10870 3875 11424 3893
rect 11930 3884 12048 3904
rect 12068 3884 12079 3904
rect 11930 3876 12079 3884
rect 12146 3908 12505 3912
rect 12146 3903 12468 3908
rect 12146 3879 12259 3903
rect 12283 3884 12468 3903
rect 12492 3884 12505 3908
rect 12283 3879 12505 3884
rect 12146 3876 12505 3879
rect 12567 3876 12602 3913
rect 12670 3910 12770 3913
rect 12670 3906 12737 3910
rect 12670 3880 12682 3906
rect 12708 3884 12737 3906
rect 12763 3884 12770 3910
rect 12708 3880 12770 3884
rect 12670 3876 12770 3880
rect 10346 3816 10383 3825
rect 10790 3816 10827 3822
rect 10870 3816 10896 3875
rect 11403 3856 11424 3875
rect 10790 3813 10896 3816
rect 10790 3795 10799 3813
rect 10817 3799 10896 3813
rect 10981 3831 11231 3855
rect 10817 3797 10893 3799
rect 10817 3795 10827 3797
rect 10790 3785 10827 3795
rect 10058 3774 10095 3775
rect 10008 3765 10095 3774
rect 10008 3745 10066 3765
rect 10086 3745 10095 3765
rect 10008 3735 10095 3745
rect 10154 3765 10191 3775
rect 10154 3745 10162 3765
rect 10182 3745 10191 3765
rect 10349 3750 10386 3754
rect 10008 3734 10039 3735
rect 10154 3674 10191 3745
rect 9941 3650 10191 3674
rect 10347 3744 10386 3750
rect 10347 3726 10358 3744
rect 10376 3726 10386 3744
rect 10347 3717 10386 3726
rect 10795 3720 10826 3785
rect 10981 3760 11018 3831
rect 11133 3770 11164 3771
rect 10981 3740 10990 3760
rect 11010 3740 11018 3760
rect 10981 3730 11018 3740
rect 11077 3760 11164 3770
rect 11077 3740 11086 3760
rect 11106 3740 11164 3760
rect 11077 3731 11164 3740
rect 11077 3730 11114 3731
rect 9097 3645 9134 3646
rect 8520 3624 8556 3645
rect 8946 3624 8977 3645
rect 9733 3626 9770 3649
rect 10347 3639 10382 3717
rect 10794 3711 10831 3720
rect 10794 3693 10804 3711
rect 10822 3693 10831 3711
rect 10794 3683 10831 3693
rect 11133 3678 11164 3731
rect 11194 3760 11231 3831
rect 11402 3836 11795 3856
rect 11815 3836 11818 3856
rect 12146 3855 12177 3876
rect 12567 3855 12603 3876
rect 11989 3854 12026 3855
rect 11402 3831 11818 3836
rect 11988 3845 12026 3854
rect 11402 3830 11743 3831
rect 11346 3770 11377 3771
rect 11194 3740 11203 3760
rect 11223 3740 11231 3760
rect 11194 3730 11231 3740
rect 11290 3763 11377 3770
rect 11290 3760 11351 3763
rect 11290 3740 11299 3760
rect 11319 3743 11351 3760
rect 11372 3743 11377 3763
rect 11319 3740 11377 3743
rect 11290 3733 11377 3740
rect 11402 3760 11439 3830
rect 11705 3829 11742 3830
rect 11988 3825 11997 3845
rect 12017 3825 12026 3845
rect 11988 3817 12026 3825
rect 12092 3849 12177 3855
rect 12202 3854 12239 3855
rect 12092 3829 12100 3849
rect 12120 3829 12177 3849
rect 12092 3821 12177 3829
rect 12201 3845 12239 3854
rect 12201 3825 12210 3845
rect 12230 3825 12239 3845
rect 12092 3820 12128 3821
rect 12201 3817 12239 3825
rect 12305 3849 12390 3855
rect 12410 3854 12447 3855
rect 12305 3829 12313 3849
rect 12333 3848 12390 3849
rect 12333 3829 12362 3848
rect 12305 3828 12362 3829
rect 12383 3828 12390 3848
rect 12305 3821 12390 3828
rect 12409 3845 12447 3854
rect 12409 3825 12418 3845
rect 12438 3825 12447 3845
rect 12305 3820 12341 3821
rect 12409 3817 12447 3825
rect 12513 3849 12657 3855
rect 12513 3829 12521 3849
rect 12541 3829 12573 3849
rect 12597 3829 12629 3849
rect 12649 3829 12657 3849
rect 12513 3821 12657 3829
rect 12513 3820 12549 3821
rect 12621 3820 12657 3821
rect 12723 3854 12760 3855
rect 12723 3853 12761 3854
rect 12723 3845 12787 3853
rect 12723 3825 12732 3845
rect 12752 3831 12787 3845
rect 12807 3831 12810 3851
rect 12752 3826 12810 3831
rect 12752 3825 12787 3826
rect 11989 3788 12026 3817
rect 11990 3786 12026 3788
rect 12202 3786 12239 3817
rect 11554 3770 11590 3771
rect 11402 3740 11411 3760
rect 11431 3740 11439 3760
rect 11290 3731 11346 3733
rect 11290 3730 11327 3731
rect 11402 3730 11439 3740
rect 11498 3760 11646 3770
rect 11746 3767 11842 3769
rect 11498 3740 11507 3760
rect 11527 3740 11617 3760
rect 11637 3740 11646 3760
rect 11498 3731 11646 3740
rect 11704 3760 11842 3767
rect 11990 3764 12239 3786
rect 12410 3785 12447 3817
rect 12723 3813 12787 3825
rect 12827 3787 12854 3965
rect 12686 3785 12854 3787
rect 12410 3781 12854 3785
rect 11704 3740 11713 3760
rect 11733 3740 11842 3760
rect 12410 3762 12459 3781
rect 12479 3762 12854 3781
rect 12410 3759 12854 3762
rect 12686 3758 12854 3759
rect 11704 3731 11842 3740
rect 11498 3730 11535 3731
rect 11554 3679 11590 3731
rect 11609 3730 11646 3731
rect 11705 3730 11742 3731
rect 11025 3677 11066 3678
rect 10917 3670 11066 3677
rect 10917 3650 11035 3670
rect 11055 3650 11066 3670
rect 10917 3642 11066 3650
rect 11133 3674 11492 3678
rect 11133 3669 11455 3674
rect 11133 3645 11246 3669
rect 11270 3650 11455 3669
rect 11479 3650 11492 3674
rect 11270 3645 11492 3650
rect 11133 3642 11492 3645
rect 11554 3642 11589 3679
rect 11657 3676 11757 3679
rect 11657 3672 11724 3676
rect 11657 3646 11669 3672
rect 11695 3650 11724 3672
rect 11750 3650 11757 3676
rect 11695 3646 11757 3650
rect 11657 3642 11757 3646
rect 10344 3629 10382 3639
rect 9733 3625 9903 3626
rect 10344 3625 10354 3629
rect 8353 3620 8453 3624
rect 8353 3616 8415 3620
rect 8353 3590 8360 3616
rect 8386 3594 8415 3616
rect 8441 3594 8453 3620
rect 8386 3590 8453 3594
rect 8353 3587 8453 3590
rect 8521 3587 8556 3624
rect 8618 3621 8977 3624
rect 8618 3616 8840 3621
rect 8618 3592 8631 3616
rect 8655 3597 8840 3616
rect 8864 3597 8977 3621
rect 8655 3592 8977 3597
rect 8618 3588 8977 3592
rect 9044 3616 9193 3624
rect 9044 3596 9055 3616
rect 9075 3596 9193 3616
rect 9733 3611 10354 3625
rect 10372 3611 10382 3629
rect 11133 3621 11164 3642
rect 11554 3621 11590 3642
rect 9733 3605 10382 3611
rect 10797 3612 10834 3621
rect 10976 3620 11013 3621
rect 9733 3604 10381 3605
rect 10344 3602 10381 3604
rect 9044 3589 9193 3596
rect 10797 3594 10806 3612
rect 10824 3594 10834 3612
rect 9044 3588 9085 3589
rect 8368 3535 8405 3536
rect 8464 3535 8501 3536
rect 8520 3535 8556 3587
rect 8575 3535 8612 3536
rect 8268 3526 8406 3535
rect 8268 3506 8377 3526
rect 8397 3506 8406 3526
rect 8268 3499 8406 3506
rect 8464 3526 8612 3535
rect 8464 3506 8473 3526
rect 8493 3506 8583 3526
rect 8603 3506 8612 3526
rect 8268 3497 8364 3499
rect 8464 3496 8612 3506
rect 8671 3526 8708 3536
rect 8783 3535 8820 3536
rect 8764 3533 8820 3535
rect 8671 3506 8679 3526
rect 8699 3506 8708 3526
rect 8520 3495 8556 3496
rect 8368 3436 8405 3437
rect 8671 3436 8708 3506
rect 8733 3526 8820 3533
rect 8733 3523 8791 3526
rect 8733 3503 8738 3523
rect 8759 3506 8791 3523
rect 8811 3506 8820 3526
rect 8759 3503 8820 3506
rect 8733 3496 8820 3503
rect 8879 3526 8916 3536
rect 8879 3506 8887 3526
rect 8907 3506 8916 3526
rect 8733 3495 8764 3496
rect 8367 3435 8708 3436
rect 8292 3430 8708 3435
rect 8292 3410 8295 3430
rect 8315 3410 8708 3430
rect 8879 3435 8916 3506
rect 8946 3535 8977 3588
rect 10797 3584 10834 3594
rect 10798 3549 10834 3584
rect 10975 3611 11013 3620
rect 10975 3591 10984 3611
rect 11004 3591 11013 3611
rect 10975 3583 11013 3591
rect 11079 3615 11164 3621
rect 11189 3620 11226 3621
rect 11079 3595 11087 3615
rect 11107 3595 11164 3615
rect 11079 3587 11164 3595
rect 11188 3611 11226 3620
rect 11188 3591 11197 3611
rect 11217 3591 11226 3611
rect 11079 3586 11115 3587
rect 11188 3583 11226 3591
rect 11292 3615 11377 3621
rect 11397 3620 11434 3621
rect 11292 3595 11300 3615
rect 11320 3614 11377 3615
rect 11320 3595 11349 3614
rect 11292 3594 11349 3595
rect 11370 3594 11377 3614
rect 11292 3587 11377 3594
rect 11396 3611 11434 3620
rect 11396 3591 11405 3611
rect 11425 3591 11434 3611
rect 11292 3586 11328 3587
rect 11396 3583 11434 3591
rect 11500 3615 11644 3621
rect 11500 3595 11508 3615
rect 11528 3614 11616 3615
rect 11528 3595 11556 3614
rect 11500 3593 11556 3595
rect 11578 3595 11616 3614
rect 11636 3595 11644 3615
rect 11578 3593 11644 3595
rect 11500 3587 11644 3593
rect 11500 3586 11536 3587
rect 11608 3586 11644 3587
rect 11710 3620 11747 3621
rect 11710 3619 11748 3620
rect 11710 3611 11774 3619
rect 11710 3591 11719 3611
rect 11739 3597 11774 3611
rect 11794 3597 11797 3617
rect 11739 3592 11797 3597
rect 11739 3591 11774 3592
rect 10976 3554 11013 3583
rect 8996 3535 9033 3536
rect 8946 3526 9033 3535
rect 8946 3506 9004 3526
rect 9024 3506 9033 3526
rect 8946 3496 9033 3506
rect 9092 3526 9129 3536
rect 9092 3506 9100 3526
rect 9120 3506 9129 3526
rect 8946 3495 8977 3496
rect 9092 3435 9129 3506
rect 10347 3530 10384 3540
rect 10347 3512 10356 3530
rect 10374 3512 10384 3530
rect 10347 3503 10384 3512
rect 10796 3508 10834 3549
rect 10977 3552 11013 3554
rect 11189 3552 11226 3583
rect 10977 3530 11226 3552
rect 11397 3551 11434 3583
rect 11710 3579 11774 3591
rect 11814 3553 11841 3731
rect 11673 3551 11841 3553
rect 11397 3525 11841 3551
rect 11398 3508 11422 3525
rect 11673 3524 11841 3525
rect 10347 3479 10382 3503
rect 10345 3455 10382 3479
rect 10344 3449 10382 3455
rect 8879 3411 9129 3435
rect 9755 3431 10382 3449
rect 10796 3490 11423 3508
rect 12049 3504 12299 3528
rect 10796 3484 10834 3490
rect 10796 3460 10833 3484
rect 10796 3436 10831 3460
rect 9337 3414 9505 3415
rect 9756 3414 9780 3431
rect 9337 3388 9781 3414
rect 9337 3386 9505 3388
rect 9337 3208 9364 3386
rect 9404 3348 9468 3360
rect 9744 3356 9781 3388
rect 9952 3387 10201 3409
rect 9952 3356 9989 3387
rect 10165 3385 10201 3387
rect 10344 3390 10382 3431
rect 10794 3427 10831 3436
rect 10794 3409 10804 3427
rect 10822 3409 10831 3427
rect 10794 3399 10831 3409
rect 12049 3433 12086 3504
rect 12201 3443 12232 3444
rect 12049 3413 12058 3433
rect 12078 3413 12086 3433
rect 12049 3403 12086 3413
rect 12145 3433 12232 3443
rect 12145 3413 12154 3433
rect 12174 3413 12232 3433
rect 12145 3404 12232 3413
rect 12145 3403 12182 3404
rect 10165 3356 10202 3385
rect 9404 3347 9439 3348
rect 9381 3342 9439 3347
rect 9381 3322 9384 3342
rect 9404 3328 9439 3342
rect 9459 3328 9468 3348
rect 9404 3320 9468 3328
rect 9430 3319 9468 3320
rect 9431 3318 9468 3319
rect 9534 3352 9570 3353
rect 9642 3352 9678 3353
rect 9534 3346 9678 3352
rect 9534 3344 9600 3346
rect 9534 3324 9542 3344
rect 9562 3325 9600 3344
rect 9622 3344 9678 3346
rect 9622 3325 9650 3344
rect 9562 3324 9650 3325
rect 9670 3324 9678 3344
rect 9534 3318 9678 3324
rect 9744 3348 9782 3356
rect 9850 3352 9886 3353
rect 9744 3328 9753 3348
rect 9773 3328 9782 3348
rect 9744 3319 9782 3328
rect 9801 3345 9886 3352
rect 9801 3325 9808 3345
rect 9829 3344 9886 3345
rect 9829 3325 9858 3344
rect 9801 3324 9858 3325
rect 9878 3324 9886 3344
rect 9744 3318 9781 3319
rect 9801 3318 9886 3324
rect 9952 3348 9990 3356
rect 10063 3352 10099 3353
rect 9952 3328 9961 3348
rect 9981 3328 9990 3348
rect 9952 3319 9990 3328
rect 10014 3344 10099 3352
rect 10014 3324 10071 3344
rect 10091 3324 10099 3344
rect 9952 3318 9989 3319
rect 10014 3318 10099 3324
rect 10165 3348 10203 3356
rect 10165 3328 10174 3348
rect 10194 3328 10203 3348
rect 10165 3319 10203 3328
rect 10344 3355 10380 3390
rect 10344 3345 10381 3355
rect 12201 3351 12232 3404
rect 12262 3433 12299 3504
rect 12470 3509 12863 3529
rect 12883 3509 12886 3529
rect 12470 3504 12886 3509
rect 12470 3503 12811 3504
rect 12414 3443 12445 3444
rect 12262 3413 12271 3433
rect 12291 3413 12299 3433
rect 12262 3403 12299 3413
rect 12358 3436 12445 3443
rect 12358 3433 12419 3436
rect 12358 3413 12367 3433
rect 12387 3416 12419 3433
rect 12440 3416 12445 3436
rect 12387 3413 12445 3416
rect 12358 3406 12445 3413
rect 12470 3433 12507 3503
rect 12773 3502 12810 3503
rect 12622 3443 12658 3444
rect 12470 3413 12479 3433
rect 12499 3413 12507 3433
rect 12358 3404 12414 3406
rect 12358 3403 12395 3404
rect 12470 3403 12507 3413
rect 12566 3433 12714 3443
rect 12814 3440 12910 3442
rect 12566 3413 12575 3433
rect 12595 3413 12685 3433
rect 12705 3413 12714 3433
rect 12566 3404 12714 3413
rect 12772 3433 12910 3440
rect 12772 3413 12781 3433
rect 12801 3413 12910 3433
rect 12772 3404 12910 3413
rect 12566 3403 12603 3404
rect 12622 3352 12658 3404
rect 12677 3403 12714 3404
rect 12773 3403 12810 3404
rect 12093 3350 12134 3351
rect 10344 3327 10354 3345
rect 10372 3327 10381 3345
rect 11985 3343 12134 3350
rect 10797 3335 10834 3337
rect 10797 3334 11445 3335
rect 10165 3318 10202 3319
rect 10344 3318 10381 3327
rect 10796 3328 11445 3334
rect 9588 3297 9624 3318
rect 10014 3297 10045 3318
rect 10796 3310 10806 3328
rect 10824 3314 11445 3328
rect 11985 3323 12103 3343
rect 12123 3323 12134 3343
rect 11985 3315 12134 3323
rect 12201 3347 12560 3351
rect 12201 3342 12523 3347
rect 12201 3318 12314 3342
rect 12338 3323 12523 3342
rect 12547 3323 12560 3347
rect 12338 3318 12560 3323
rect 12201 3315 12560 3318
rect 12622 3315 12657 3352
rect 12725 3349 12825 3352
rect 12725 3345 12792 3349
rect 12725 3319 12737 3345
rect 12763 3323 12792 3345
rect 12818 3323 12825 3349
rect 12763 3319 12825 3323
rect 12725 3315 12825 3319
rect 10824 3310 10834 3314
rect 11275 3313 11445 3314
rect 10796 3300 10834 3310
rect 9421 3293 9521 3297
rect 9421 3289 9483 3293
rect 9421 3263 9428 3289
rect 9454 3267 9483 3289
rect 9509 3267 9521 3293
rect 9454 3263 9521 3267
rect 9421 3260 9521 3263
rect 9589 3260 9624 3297
rect 9686 3294 10045 3297
rect 9686 3289 9908 3294
rect 9686 3265 9699 3289
rect 9723 3270 9908 3289
rect 9932 3270 10045 3294
rect 9723 3265 10045 3270
rect 9686 3261 10045 3265
rect 10112 3289 10261 3297
rect 10112 3269 10123 3289
rect 10143 3269 10261 3289
rect 10112 3262 10261 3269
rect 10112 3261 10153 3262
rect 9436 3208 9473 3209
rect 9532 3208 9569 3209
rect 9588 3208 9624 3260
rect 9643 3208 9680 3209
rect 9336 3199 9474 3208
rect 8324 3180 8492 3181
rect 8324 3177 8768 3180
rect 8324 3158 8699 3177
rect 8719 3158 8768 3177
rect 9336 3179 9445 3199
rect 9465 3179 9474 3199
rect 8324 3154 8768 3158
rect 8324 3152 8492 3154
rect 8324 2974 8351 3152
rect 8391 3114 8455 3126
rect 8731 3122 8768 3154
rect 8939 3153 9188 3175
rect 9336 3172 9474 3179
rect 9532 3199 9680 3208
rect 9532 3179 9541 3199
rect 9561 3179 9651 3199
rect 9671 3179 9680 3199
rect 9336 3170 9432 3172
rect 9532 3169 9680 3179
rect 9739 3199 9776 3209
rect 9851 3208 9888 3209
rect 9832 3206 9888 3208
rect 9739 3179 9747 3199
rect 9767 3179 9776 3199
rect 9588 3168 9624 3169
rect 8939 3122 8976 3153
rect 9152 3151 9188 3153
rect 9152 3122 9189 3151
rect 8391 3113 8426 3114
rect 8368 3108 8426 3113
rect 8368 3088 8371 3108
rect 8391 3094 8426 3108
rect 8446 3094 8455 3114
rect 8391 3086 8455 3094
rect 8417 3085 8455 3086
rect 8418 3084 8455 3085
rect 8521 3118 8557 3119
rect 8629 3118 8665 3119
rect 8521 3110 8665 3118
rect 8521 3090 8529 3110
rect 8549 3090 8581 3110
rect 8605 3090 8637 3110
rect 8657 3090 8665 3110
rect 8521 3084 8665 3090
rect 8731 3114 8769 3122
rect 8837 3118 8873 3119
rect 8731 3094 8740 3114
rect 8760 3094 8769 3114
rect 8731 3085 8769 3094
rect 8788 3111 8873 3118
rect 8788 3091 8795 3111
rect 8816 3110 8873 3111
rect 8816 3091 8845 3110
rect 8788 3090 8845 3091
rect 8865 3090 8873 3110
rect 8731 3084 8768 3085
rect 8788 3084 8873 3090
rect 8939 3114 8977 3122
rect 9050 3118 9086 3119
rect 8939 3094 8948 3114
rect 8968 3094 8977 3114
rect 8939 3085 8977 3094
rect 9001 3110 9086 3118
rect 9001 3090 9058 3110
rect 9078 3090 9086 3110
rect 8939 3084 8976 3085
rect 9001 3084 9086 3090
rect 9152 3114 9190 3122
rect 9152 3094 9161 3114
rect 9181 3094 9190 3114
rect 9436 3109 9473 3110
rect 9739 3109 9776 3179
rect 9801 3199 9888 3206
rect 9801 3196 9859 3199
rect 9801 3176 9806 3196
rect 9827 3179 9859 3196
rect 9879 3179 9888 3199
rect 9827 3176 9888 3179
rect 9801 3169 9888 3176
rect 9947 3199 9984 3209
rect 9947 3179 9955 3199
rect 9975 3179 9984 3199
rect 9801 3168 9832 3169
rect 9435 3108 9776 3109
rect 9152 3085 9190 3094
rect 9360 3103 9776 3108
rect 9152 3084 9189 3085
rect 8575 3063 8611 3084
rect 9001 3063 9032 3084
rect 9360 3083 9363 3103
rect 9383 3083 9776 3103
rect 9947 3108 9984 3179
rect 10014 3208 10045 3261
rect 10347 3246 10384 3256
rect 10347 3228 10356 3246
rect 10374 3228 10384 3246
rect 10347 3219 10384 3228
rect 10796 3222 10831 3300
rect 11408 3290 11445 3313
rect 12201 3294 12232 3315
rect 12622 3294 12658 3315
rect 12044 3293 12081 3294
rect 10064 3208 10101 3209
rect 10014 3199 10101 3208
rect 10014 3179 10072 3199
rect 10092 3179 10101 3199
rect 10014 3169 10101 3179
rect 10160 3199 10197 3209
rect 10160 3179 10168 3199
rect 10188 3179 10197 3199
rect 10014 3168 10045 3169
rect 10160 3108 10197 3179
rect 10352 3154 10383 3219
rect 10792 3213 10831 3222
rect 10792 3195 10802 3213
rect 10820 3195 10831 3213
rect 10792 3189 10831 3195
rect 10987 3265 11237 3289
rect 10987 3194 11024 3265
rect 11139 3204 11170 3205
rect 10792 3185 10829 3189
rect 10987 3174 10996 3194
rect 11016 3174 11024 3194
rect 10987 3164 11024 3174
rect 11083 3194 11170 3204
rect 11083 3174 11092 3194
rect 11112 3174 11170 3194
rect 11083 3165 11170 3174
rect 11083 3164 11120 3165
rect 10351 3144 10388 3154
rect 10351 3142 10361 3144
rect 10285 3140 10361 3142
rect 9947 3084 10197 3108
rect 10282 3126 10361 3140
rect 10379 3126 10388 3144
rect 10282 3123 10388 3126
rect 9754 3064 9775 3083
rect 10282 3064 10308 3123
rect 10351 3117 10388 3123
rect 10795 3114 10832 3123
rect 8408 3059 8508 3063
rect 8408 3055 8470 3059
rect 8408 3029 8415 3055
rect 8441 3033 8470 3055
rect 8496 3033 8508 3059
rect 8441 3029 8508 3033
rect 8408 3026 8508 3029
rect 8576 3026 8611 3063
rect 8673 3060 9032 3063
rect 8673 3055 8895 3060
rect 8673 3031 8686 3055
rect 8710 3036 8895 3055
rect 8919 3036 9032 3060
rect 8710 3031 9032 3036
rect 8673 3027 9032 3031
rect 9099 3055 9248 3063
rect 9099 3035 9110 3055
rect 9130 3035 9248 3055
rect 9754 3046 10308 3064
rect 10793 3096 10804 3114
rect 10822 3096 10832 3114
rect 11139 3112 11170 3165
rect 11200 3194 11237 3265
rect 11408 3270 11801 3290
rect 11821 3270 11824 3290
rect 11408 3265 11824 3270
rect 12043 3284 12081 3293
rect 11408 3264 11749 3265
rect 12043 3264 12052 3284
rect 12072 3264 12081 3284
rect 11352 3204 11383 3205
rect 11200 3174 11209 3194
rect 11229 3174 11237 3194
rect 11200 3164 11237 3174
rect 11296 3197 11383 3204
rect 11296 3194 11357 3197
rect 11296 3174 11305 3194
rect 11325 3177 11357 3194
rect 11378 3177 11383 3197
rect 11325 3174 11383 3177
rect 11296 3167 11383 3174
rect 11408 3194 11445 3264
rect 11711 3263 11748 3264
rect 12043 3256 12081 3264
rect 12147 3288 12232 3294
rect 12257 3293 12294 3294
rect 12147 3268 12155 3288
rect 12175 3268 12232 3288
rect 12147 3260 12232 3268
rect 12256 3284 12294 3293
rect 12256 3264 12265 3284
rect 12285 3264 12294 3284
rect 12147 3259 12183 3260
rect 12256 3256 12294 3264
rect 12360 3288 12445 3294
rect 12465 3293 12502 3294
rect 12360 3268 12368 3288
rect 12388 3287 12445 3288
rect 12388 3268 12417 3287
rect 12360 3267 12417 3268
rect 12438 3267 12445 3287
rect 12360 3260 12445 3267
rect 12464 3284 12502 3293
rect 12464 3264 12473 3284
rect 12493 3264 12502 3284
rect 12360 3259 12396 3260
rect 12464 3256 12502 3264
rect 12568 3288 12712 3294
rect 12568 3268 12576 3288
rect 12596 3286 12684 3288
rect 12596 3269 12632 3286
rect 12656 3269 12684 3286
rect 12596 3268 12684 3269
rect 12704 3268 12712 3288
rect 12568 3260 12712 3268
rect 12568 3259 12604 3260
rect 12676 3259 12712 3260
rect 12778 3293 12815 3294
rect 12778 3292 12816 3293
rect 12778 3284 12842 3292
rect 12778 3264 12787 3284
rect 12807 3270 12842 3284
rect 12862 3270 12865 3290
rect 12807 3265 12865 3270
rect 12807 3264 12842 3265
rect 12044 3227 12081 3256
rect 12045 3225 12081 3227
rect 12257 3225 12294 3256
rect 11560 3204 11596 3205
rect 11408 3174 11417 3194
rect 11437 3174 11445 3194
rect 11296 3165 11352 3167
rect 11296 3164 11333 3165
rect 11408 3164 11445 3174
rect 11504 3194 11652 3204
rect 12045 3203 12294 3225
rect 12465 3224 12502 3256
rect 12778 3252 12842 3264
rect 12882 3226 12909 3404
rect 12741 3224 12909 3226
rect 12465 3213 12909 3224
rect 11752 3201 11848 3203
rect 11504 3174 11513 3194
rect 11533 3174 11623 3194
rect 11643 3174 11652 3194
rect 11504 3165 11652 3174
rect 11710 3194 11848 3201
rect 12465 3198 12911 3213
rect 12741 3197 12911 3198
rect 11710 3174 11719 3194
rect 11739 3174 11848 3194
rect 11710 3165 11848 3174
rect 11504 3164 11541 3165
rect 11560 3113 11596 3165
rect 11615 3164 11652 3165
rect 11711 3164 11748 3165
rect 11031 3111 11072 3112
rect 10354 3053 10391 3055
rect 10282 3045 10308 3046
rect 10351 3045 10391 3053
rect 9099 3028 9248 3035
rect 10351 3033 10363 3045
rect 10342 3028 10363 3033
rect 9099 3027 9140 3028
rect 9758 3027 10363 3028
rect 10381 3027 10391 3045
rect 8423 2974 8460 2975
rect 8519 2974 8556 2975
rect 8575 2974 8611 3026
rect 8630 2974 8667 2975
rect 8323 2965 8461 2974
rect 8323 2945 8432 2965
rect 8452 2945 8461 2965
rect 8323 2938 8461 2945
rect 8519 2965 8667 2974
rect 8519 2945 8528 2965
rect 8548 2945 8638 2965
rect 8658 2945 8667 2965
rect 8323 2936 8419 2938
rect 8519 2935 8667 2945
rect 8726 2965 8763 2975
rect 8838 2974 8875 2975
rect 8819 2972 8875 2974
rect 8726 2945 8734 2965
rect 8754 2945 8763 2965
rect 8575 2934 8611 2935
rect 8423 2875 8460 2876
rect 8726 2875 8763 2945
rect 8788 2965 8875 2972
rect 8788 2962 8846 2965
rect 8788 2942 8793 2962
rect 8814 2945 8846 2962
rect 8866 2945 8875 2965
rect 8814 2942 8875 2945
rect 8788 2935 8875 2942
rect 8934 2965 8971 2975
rect 8934 2945 8942 2965
rect 8962 2945 8971 2965
rect 8788 2934 8819 2935
rect 8422 2874 8763 2875
rect 8347 2869 8763 2874
rect 8347 2849 8350 2869
rect 8370 2849 8763 2869
rect 8934 2874 8971 2945
rect 9001 2974 9032 3027
rect 9758 3018 10391 3027
rect 9758 3011 10390 3018
rect 9758 3009 9820 3011
rect 9336 2999 9504 3000
rect 9758 2999 9780 3009
rect 9051 2974 9088 2975
rect 9001 2965 9088 2974
rect 9001 2945 9059 2965
rect 9079 2945 9088 2965
rect 9001 2935 9088 2945
rect 9147 2965 9184 2975
rect 9147 2945 9155 2965
rect 9175 2945 9184 2965
rect 9001 2934 9032 2935
rect 9147 2874 9184 2945
rect 8934 2850 9184 2874
rect 9336 2973 9780 2999
rect 9336 2971 9504 2973
rect 9336 2793 9363 2971
rect 9403 2933 9467 2945
rect 9743 2941 9780 2973
rect 9951 2972 10200 2994
rect 9951 2941 9988 2972
rect 10164 2970 10200 2972
rect 10164 2941 10201 2970
rect 9403 2932 9438 2933
rect 9380 2927 9438 2932
rect 9380 2907 9383 2927
rect 9403 2913 9438 2927
rect 9458 2913 9467 2933
rect 9403 2905 9467 2913
rect 9429 2904 9467 2905
rect 9430 2903 9467 2904
rect 9533 2937 9569 2938
rect 9641 2937 9677 2938
rect 9533 2929 9677 2937
rect 9533 2909 9541 2929
rect 9561 2909 9590 2929
rect 9533 2908 9590 2909
rect 9612 2909 9649 2929
rect 9669 2909 9677 2929
rect 9612 2908 9677 2909
rect 9533 2903 9677 2908
rect 9743 2933 9781 2941
rect 9849 2937 9885 2938
rect 9743 2913 9752 2933
rect 9772 2913 9781 2933
rect 9743 2904 9781 2913
rect 9800 2930 9885 2937
rect 9800 2910 9807 2930
rect 9828 2929 9885 2930
rect 9828 2910 9857 2929
rect 9800 2909 9857 2910
rect 9877 2909 9885 2929
rect 9743 2903 9780 2904
rect 9800 2903 9885 2909
rect 9951 2933 9989 2941
rect 10062 2937 10098 2938
rect 9951 2913 9960 2933
rect 9980 2913 9989 2933
rect 9951 2904 9989 2913
rect 10013 2929 10098 2937
rect 10013 2909 10070 2929
rect 10090 2909 10098 2929
rect 9951 2903 9988 2904
rect 10013 2903 10098 2909
rect 10164 2933 10202 2941
rect 10164 2913 10173 2933
rect 10193 2913 10202 2933
rect 10164 2904 10202 2913
rect 10164 2903 10201 2904
rect 9587 2882 9623 2903
rect 10013 2882 10044 2903
rect 9420 2878 9520 2882
rect 9420 2874 9482 2878
rect 9420 2848 9427 2874
rect 9453 2852 9482 2874
rect 9508 2852 9520 2878
rect 9453 2848 9520 2852
rect 9420 2845 9520 2848
rect 9588 2845 9623 2882
rect 9685 2879 10044 2882
rect 9685 2874 9907 2879
rect 9685 2850 9698 2874
rect 9722 2855 9907 2874
rect 9931 2855 10044 2879
rect 9722 2850 10044 2855
rect 9685 2846 10044 2850
rect 10111 2874 10260 2882
rect 10111 2854 10122 2874
rect 10142 2854 10260 2874
rect 10111 2847 10260 2854
rect 10351 2862 10390 3011
rect 10793 2947 10832 3096
rect 10923 3104 11072 3111
rect 10923 3084 11041 3104
rect 11061 3084 11072 3104
rect 10923 3076 11072 3084
rect 11139 3108 11498 3112
rect 11139 3103 11461 3108
rect 11139 3079 11252 3103
rect 11276 3084 11461 3103
rect 11485 3084 11498 3108
rect 11276 3079 11498 3084
rect 11139 3076 11498 3079
rect 11560 3076 11595 3113
rect 11663 3110 11763 3113
rect 11663 3106 11730 3110
rect 11663 3080 11675 3106
rect 11701 3084 11730 3106
rect 11756 3084 11763 3110
rect 11701 3080 11763 3084
rect 11663 3076 11763 3080
rect 11139 3055 11170 3076
rect 11560 3055 11596 3076
rect 10982 3054 11019 3055
rect 10981 3045 11019 3054
rect 10981 3025 10990 3045
rect 11010 3025 11019 3045
rect 10981 3017 11019 3025
rect 11085 3049 11170 3055
rect 11195 3054 11232 3055
rect 11085 3029 11093 3049
rect 11113 3029 11170 3049
rect 11085 3021 11170 3029
rect 11194 3045 11232 3054
rect 11194 3025 11203 3045
rect 11223 3025 11232 3045
rect 11085 3020 11121 3021
rect 11194 3017 11232 3025
rect 11298 3049 11383 3055
rect 11403 3054 11440 3055
rect 11298 3029 11306 3049
rect 11326 3048 11383 3049
rect 11326 3029 11355 3048
rect 11298 3028 11355 3029
rect 11376 3028 11383 3048
rect 11298 3021 11383 3028
rect 11402 3045 11440 3054
rect 11402 3025 11411 3045
rect 11431 3025 11440 3045
rect 11298 3020 11334 3021
rect 11402 3017 11440 3025
rect 11506 3050 11650 3055
rect 11506 3049 11571 3050
rect 11506 3029 11514 3049
rect 11534 3029 11571 3049
rect 11593 3049 11650 3050
rect 11593 3029 11622 3049
rect 11642 3029 11650 3049
rect 11506 3021 11650 3029
rect 11506 3020 11542 3021
rect 11614 3020 11650 3021
rect 11716 3054 11753 3055
rect 11716 3053 11754 3054
rect 11716 3045 11780 3053
rect 11716 3025 11725 3045
rect 11745 3031 11780 3045
rect 11800 3031 11803 3051
rect 11745 3026 11803 3031
rect 11745 3025 11780 3026
rect 10982 2988 11019 3017
rect 10983 2986 11019 2988
rect 11195 2986 11232 3017
rect 10983 2964 11232 2986
rect 11403 2985 11440 3017
rect 11716 3013 11780 3025
rect 11820 2987 11847 3165
rect 11679 2985 11847 2987
rect 11403 2959 11847 2985
rect 11999 3084 12249 3108
rect 11999 3013 12036 3084
rect 12151 3023 12182 3024
rect 11999 2993 12008 3013
rect 12028 2993 12036 3013
rect 11999 2983 12036 2993
rect 12095 3013 12182 3023
rect 12095 2993 12104 3013
rect 12124 2993 12182 3013
rect 12095 2984 12182 2993
rect 12095 2983 12132 2984
rect 11403 2949 11425 2959
rect 11679 2958 11847 2959
rect 11363 2947 11425 2949
rect 10793 2940 11425 2947
rect 10792 2931 11425 2940
rect 12151 2931 12182 2984
rect 12212 3013 12249 3084
rect 12420 3089 12813 3109
rect 12833 3089 12836 3109
rect 12420 3084 12836 3089
rect 12420 3083 12761 3084
rect 12364 3023 12395 3024
rect 12212 2993 12221 3013
rect 12241 2993 12249 3013
rect 12212 2983 12249 2993
rect 12308 3016 12395 3023
rect 12308 3013 12369 3016
rect 12308 2993 12317 3013
rect 12337 2996 12369 3013
rect 12390 2996 12395 3016
rect 12337 2993 12395 2996
rect 12308 2986 12395 2993
rect 12420 3013 12457 3083
rect 12723 3082 12760 3083
rect 12572 3023 12608 3024
rect 12420 2993 12429 3013
rect 12449 2993 12457 3013
rect 12308 2984 12364 2986
rect 12308 2983 12345 2984
rect 12420 2983 12457 2993
rect 12516 3013 12664 3023
rect 12764 3020 12860 3022
rect 12516 2993 12525 3013
rect 12545 2993 12635 3013
rect 12655 2993 12664 3013
rect 12516 2984 12664 2993
rect 12722 3013 12860 3020
rect 12722 2993 12731 3013
rect 12751 2993 12860 3013
rect 12722 2984 12860 2993
rect 12516 2983 12553 2984
rect 12572 2932 12608 2984
rect 12627 2983 12664 2984
rect 12723 2983 12760 2984
rect 10792 2913 10802 2931
rect 10820 2930 11425 2931
rect 12043 2930 12084 2931
rect 10820 2925 10841 2930
rect 10820 2913 10832 2925
rect 11935 2923 12084 2930
rect 10792 2905 10832 2913
rect 10875 2912 10901 2913
rect 10792 2903 10829 2905
rect 10111 2846 10152 2847
rect 9435 2793 9472 2794
rect 9531 2793 9568 2794
rect 9587 2793 9623 2845
rect 9642 2793 9679 2794
rect 9335 2784 9473 2793
rect 9335 2764 9444 2784
rect 9464 2764 9473 2784
rect 9335 2757 9473 2764
rect 9531 2784 9679 2793
rect 9531 2764 9540 2784
rect 9560 2764 9650 2784
rect 9670 2764 9679 2784
rect 9335 2755 9431 2757
rect 9531 2754 9679 2764
rect 9738 2784 9775 2794
rect 9850 2793 9887 2794
rect 9831 2791 9887 2793
rect 9738 2764 9746 2784
rect 9766 2764 9775 2784
rect 9587 2753 9623 2754
rect 8116 2713 8284 2714
rect 8116 2687 8560 2713
rect 8116 2685 8284 2687
rect 8116 2507 8143 2685
rect 8183 2647 8247 2659
rect 8523 2655 8560 2687
rect 8731 2686 8980 2708
rect 9435 2694 9472 2695
rect 9738 2694 9775 2764
rect 9800 2784 9887 2791
rect 9800 2781 9858 2784
rect 9800 2761 9805 2781
rect 9826 2764 9858 2781
rect 9878 2764 9887 2784
rect 9826 2761 9887 2764
rect 9800 2754 9887 2761
rect 9946 2784 9983 2794
rect 9946 2764 9954 2784
rect 9974 2764 9983 2784
rect 9800 2753 9831 2754
rect 9434 2693 9775 2694
rect 8731 2655 8768 2686
rect 8944 2684 8980 2686
rect 9359 2688 9775 2693
rect 8944 2655 8981 2684
rect 9359 2668 9362 2688
rect 9382 2668 9775 2688
rect 9946 2693 9983 2764
rect 10013 2793 10044 2846
rect 10351 2844 10361 2862
rect 10379 2844 10390 2862
rect 10875 2894 11429 2912
rect 11935 2903 12053 2923
rect 12073 2903 12084 2923
rect 11935 2895 12084 2903
rect 12151 2927 12510 2931
rect 12151 2922 12473 2927
rect 12151 2898 12264 2922
rect 12288 2903 12473 2922
rect 12497 2903 12510 2927
rect 12288 2898 12510 2903
rect 12151 2895 12510 2898
rect 12572 2895 12607 2932
rect 12675 2929 12775 2932
rect 12675 2925 12742 2929
rect 12675 2899 12687 2925
rect 12713 2903 12742 2925
rect 12768 2903 12775 2929
rect 12713 2899 12775 2903
rect 12675 2895 12775 2899
rect 10351 2835 10388 2844
rect 10795 2835 10832 2841
rect 10875 2835 10901 2894
rect 11408 2875 11429 2894
rect 10795 2832 10901 2835
rect 10795 2814 10804 2832
rect 10822 2818 10901 2832
rect 10986 2850 11236 2874
rect 10822 2816 10898 2818
rect 10822 2814 10832 2816
rect 10795 2804 10832 2814
rect 10063 2793 10100 2794
rect 10013 2784 10100 2793
rect 10013 2764 10071 2784
rect 10091 2764 10100 2784
rect 10013 2754 10100 2764
rect 10159 2784 10196 2794
rect 10159 2764 10167 2784
rect 10187 2764 10196 2784
rect 10354 2769 10391 2773
rect 10013 2753 10044 2754
rect 10159 2693 10196 2764
rect 9946 2669 10196 2693
rect 10352 2763 10391 2769
rect 10352 2745 10363 2763
rect 10381 2745 10391 2763
rect 10352 2736 10391 2745
rect 10800 2739 10831 2804
rect 10986 2779 11023 2850
rect 11138 2789 11169 2790
rect 10986 2759 10995 2779
rect 11015 2759 11023 2779
rect 10986 2749 11023 2759
rect 11082 2779 11169 2789
rect 11082 2759 11091 2779
rect 11111 2759 11169 2779
rect 11082 2750 11169 2759
rect 11082 2749 11119 2750
rect 8183 2646 8218 2647
rect 8160 2641 8218 2646
rect 8160 2621 8163 2641
rect 8183 2627 8218 2641
rect 8238 2627 8247 2647
rect 8183 2619 8247 2627
rect 8209 2618 8247 2619
rect 8210 2617 8247 2618
rect 8313 2651 8349 2652
rect 8421 2651 8457 2652
rect 8313 2645 8457 2651
rect 8313 2643 8374 2645
rect 8313 2623 8321 2643
rect 8341 2623 8374 2643
rect 8313 2619 8374 2623
rect 8399 2643 8457 2645
rect 8399 2623 8429 2643
rect 8449 2623 8457 2643
rect 8399 2619 8457 2623
rect 8313 2617 8457 2619
rect 8523 2647 8561 2655
rect 8629 2651 8665 2652
rect 8523 2627 8532 2647
rect 8552 2627 8561 2647
rect 8523 2618 8561 2627
rect 8580 2644 8665 2651
rect 8580 2624 8587 2644
rect 8608 2643 8665 2644
rect 8608 2624 8637 2643
rect 8580 2623 8637 2624
rect 8657 2623 8665 2643
rect 8523 2617 8560 2618
rect 8580 2617 8665 2623
rect 8731 2647 8769 2655
rect 8842 2651 8878 2652
rect 8731 2627 8740 2647
rect 8760 2627 8769 2647
rect 8731 2618 8769 2627
rect 8793 2643 8878 2651
rect 8793 2623 8850 2643
rect 8870 2623 8878 2643
rect 8731 2617 8768 2618
rect 8793 2617 8878 2623
rect 8944 2647 8982 2655
rect 8944 2627 8953 2647
rect 8973 2627 8982 2647
rect 8944 2618 8982 2627
rect 9738 2645 9775 2668
rect 10352 2658 10387 2736
rect 10799 2730 10836 2739
rect 10799 2712 10809 2730
rect 10827 2712 10836 2730
rect 10799 2702 10836 2712
rect 11138 2697 11169 2750
rect 11199 2779 11236 2850
rect 11407 2855 11800 2875
rect 11820 2855 11823 2875
rect 12151 2874 12182 2895
rect 12572 2874 12608 2895
rect 11994 2873 12031 2874
rect 11407 2850 11823 2855
rect 11993 2864 12031 2873
rect 11407 2849 11748 2850
rect 11351 2789 11382 2790
rect 11199 2759 11208 2779
rect 11228 2759 11236 2779
rect 11199 2749 11236 2759
rect 11295 2782 11382 2789
rect 11295 2779 11356 2782
rect 11295 2759 11304 2779
rect 11324 2762 11356 2779
rect 11377 2762 11382 2782
rect 11324 2759 11382 2762
rect 11295 2752 11382 2759
rect 11407 2779 11444 2849
rect 11710 2848 11747 2849
rect 11993 2844 12002 2864
rect 12022 2844 12031 2864
rect 11993 2836 12031 2844
rect 12097 2868 12182 2874
rect 12207 2873 12244 2874
rect 12097 2848 12105 2868
rect 12125 2848 12182 2868
rect 12097 2840 12182 2848
rect 12206 2864 12244 2873
rect 12206 2844 12215 2864
rect 12235 2844 12244 2864
rect 12097 2839 12133 2840
rect 12206 2836 12244 2844
rect 12310 2868 12395 2874
rect 12415 2873 12452 2874
rect 12310 2848 12318 2868
rect 12338 2867 12395 2868
rect 12338 2848 12367 2867
rect 12310 2847 12367 2848
rect 12388 2847 12395 2867
rect 12310 2840 12395 2847
rect 12414 2864 12452 2873
rect 12414 2844 12423 2864
rect 12443 2844 12452 2864
rect 12310 2839 12346 2840
rect 12414 2836 12452 2844
rect 12518 2869 12662 2874
rect 12518 2868 12577 2869
rect 12518 2848 12526 2868
rect 12546 2849 12577 2868
rect 12601 2868 12662 2869
rect 12601 2849 12634 2868
rect 12546 2848 12634 2849
rect 12654 2848 12662 2868
rect 12518 2840 12662 2848
rect 12518 2839 12554 2840
rect 12626 2839 12662 2840
rect 12728 2873 12765 2874
rect 12728 2872 12766 2873
rect 12728 2864 12792 2872
rect 12728 2844 12737 2864
rect 12757 2850 12792 2864
rect 12812 2850 12815 2870
rect 12757 2845 12815 2850
rect 12757 2844 12792 2845
rect 11994 2807 12031 2836
rect 11995 2805 12031 2807
rect 12207 2805 12244 2836
rect 11559 2789 11595 2790
rect 11407 2759 11416 2779
rect 11436 2759 11444 2779
rect 11295 2750 11351 2752
rect 11295 2749 11332 2750
rect 11407 2749 11444 2759
rect 11503 2779 11651 2789
rect 11751 2786 11847 2788
rect 11503 2759 11512 2779
rect 11532 2759 11622 2779
rect 11642 2759 11651 2779
rect 11503 2750 11651 2759
rect 11709 2779 11847 2786
rect 11995 2783 12244 2805
rect 12415 2804 12452 2836
rect 12728 2832 12792 2844
rect 12832 2806 12859 2984
rect 12691 2804 12859 2806
rect 12415 2800 12859 2804
rect 11709 2759 11718 2779
rect 11738 2759 11847 2779
rect 12415 2781 12464 2800
rect 12484 2781 12859 2800
rect 12415 2778 12859 2781
rect 12691 2777 12859 2778
rect 12880 2803 12911 3197
rect 12880 2777 12885 2803
rect 12904 2777 12911 2803
rect 12880 2774 12911 2777
rect 11709 2750 11847 2759
rect 11503 2749 11540 2750
rect 11559 2698 11595 2750
rect 11614 2749 11651 2750
rect 11710 2749 11747 2750
rect 11030 2696 11071 2697
rect 10922 2689 11071 2696
rect 10922 2669 11040 2689
rect 11060 2669 11071 2689
rect 10922 2661 11071 2669
rect 11138 2693 11497 2697
rect 11138 2688 11460 2693
rect 11138 2664 11251 2688
rect 11275 2669 11460 2688
rect 11484 2669 11497 2693
rect 11275 2664 11497 2669
rect 11138 2661 11497 2664
rect 11559 2661 11594 2698
rect 11662 2695 11762 2698
rect 11662 2691 11729 2695
rect 11662 2665 11674 2691
rect 11700 2669 11729 2691
rect 11755 2669 11762 2695
rect 11700 2665 11762 2669
rect 11662 2661 11762 2665
rect 10349 2648 10387 2658
rect 9738 2644 9908 2645
rect 10349 2644 10359 2648
rect 9738 2630 10359 2644
rect 10377 2630 10387 2648
rect 11138 2640 11169 2661
rect 11559 2640 11595 2661
rect 9738 2624 10387 2630
rect 10802 2631 10839 2640
rect 10981 2639 11018 2640
rect 9738 2623 10386 2624
rect 10349 2621 10386 2623
rect 8944 2617 8981 2618
rect 8367 2596 8403 2617
rect 8793 2596 8824 2617
rect 10802 2613 10811 2631
rect 10829 2613 10839 2631
rect 10802 2603 10839 2613
rect 8200 2592 8300 2596
rect 8200 2588 8262 2592
rect 8200 2562 8207 2588
rect 8233 2566 8262 2588
rect 8288 2566 8300 2592
rect 8233 2562 8300 2566
rect 8200 2559 8300 2562
rect 8368 2559 8403 2596
rect 8465 2593 8824 2596
rect 8465 2588 8687 2593
rect 8465 2564 8478 2588
rect 8502 2569 8687 2588
rect 8711 2569 8824 2593
rect 8502 2564 8824 2569
rect 8465 2560 8824 2564
rect 8891 2588 9040 2596
rect 8891 2568 8902 2588
rect 8922 2568 9040 2588
rect 10803 2568 10839 2603
rect 10980 2630 11018 2639
rect 10980 2610 10989 2630
rect 11009 2610 11018 2630
rect 10980 2602 11018 2610
rect 11084 2634 11169 2640
rect 11194 2639 11231 2640
rect 11084 2614 11092 2634
rect 11112 2614 11169 2634
rect 11084 2606 11169 2614
rect 11193 2630 11231 2639
rect 11193 2610 11202 2630
rect 11222 2610 11231 2630
rect 11084 2605 11120 2606
rect 11193 2602 11231 2610
rect 11297 2634 11382 2640
rect 11402 2639 11439 2640
rect 11297 2614 11305 2634
rect 11325 2633 11382 2634
rect 11325 2614 11354 2633
rect 11297 2613 11354 2614
rect 11375 2613 11382 2633
rect 11297 2606 11382 2613
rect 11401 2630 11439 2639
rect 11401 2610 11410 2630
rect 11430 2610 11439 2630
rect 11297 2605 11333 2606
rect 11401 2602 11439 2610
rect 11505 2634 11649 2640
rect 11505 2614 11513 2634
rect 11533 2633 11621 2634
rect 11533 2614 11561 2633
rect 11505 2612 11561 2614
rect 11583 2614 11621 2633
rect 11641 2614 11649 2634
rect 11583 2612 11649 2614
rect 11505 2606 11649 2612
rect 11505 2605 11541 2606
rect 11613 2605 11649 2606
rect 11715 2639 11752 2640
rect 11715 2638 11753 2639
rect 11715 2630 11779 2638
rect 11715 2610 11724 2630
rect 11744 2616 11779 2630
rect 11799 2616 11802 2636
rect 11744 2611 11802 2616
rect 11744 2610 11779 2611
rect 10981 2573 11018 2602
rect 8891 2561 9040 2568
rect 8891 2560 8932 2561
rect 8215 2507 8252 2508
rect 8311 2507 8348 2508
rect 8367 2507 8403 2559
rect 8422 2507 8459 2508
rect 8115 2498 8253 2507
rect 8115 2478 8224 2498
rect 8244 2478 8253 2498
rect 8115 2471 8253 2478
rect 8311 2498 8459 2507
rect 8311 2478 8320 2498
rect 8340 2478 8430 2498
rect 8450 2478 8459 2498
rect 8115 2469 8211 2471
rect 8311 2468 8459 2478
rect 8518 2498 8555 2508
rect 8630 2507 8667 2508
rect 8611 2505 8667 2507
rect 8518 2478 8526 2498
rect 8546 2478 8555 2498
rect 8367 2467 8403 2468
rect 8215 2408 8252 2409
rect 8518 2408 8555 2478
rect 8580 2498 8667 2505
rect 8580 2495 8638 2498
rect 8580 2475 8585 2495
rect 8606 2478 8638 2495
rect 8658 2478 8667 2498
rect 8606 2475 8667 2478
rect 8580 2468 8667 2475
rect 8726 2498 8763 2508
rect 8726 2478 8734 2498
rect 8754 2478 8763 2498
rect 8580 2467 8611 2468
rect 8214 2407 8555 2408
rect 8139 2402 8555 2407
rect 8139 2382 8142 2402
rect 8162 2382 8555 2402
rect 8726 2407 8763 2478
rect 8793 2507 8824 2560
rect 10352 2549 10389 2559
rect 10352 2531 10361 2549
rect 10379 2531 10389 2549
rect 10352 2522 10389 2531
rect 10801 2527 10839 2568
rect 10982 2571 11018 2573
rect 11194 2571 11231 2602
rect 10982 2549 11231 2571
rect 11402 2570 11439 2602
rect 11715 2598 11779 2610
rect 11819 2572 11846 2750
rect 11678 2570 11846 2572
rect 11402 2544 11846 2570
rect 11403 2527 11427 2544
rect 11678 2543 11846 2544
rect 12214 2572 12464 2596
rect 8843 2507 8880 2508
rect 8793 2498 8880 2507
rect 8793 2478 8851 2498
rect 8871 2478 8880 2498
rect 8793 2468 8880 2478
rect 8939 2498 8976 2508
rect 8939 2478 8947 2498
rect 8967 2478 8976 2498
rect 8793 2467 8824 2468
rect 8939 2407 8976 2478
rect 10352 2476 10387 2522
rect 10801 2509 11428 2527
rect 10801 2503 10839 2509
rect 10351 2470 10389 2476
rect 9762 2452 10389 2470
rect 10803 2457 10838 2503
rect 12214 2501 12251 2572
rect 12366 2511 12397 2512
rect 12214 2481 12223 2501
rect 12243 2481 12251 2501
rect 12214 2471 12251 2481
rect 12310 2501 12397 2511
rect 12310 2481 12319 2501
rect 12339 2481 12397 2501
rect 12310 2472 12397 2481
rect 12310 2471 12347 2472
rect 8726 2383 8976 2407
rect 9344 2435 9512 2436
rect 9763 2435 9787 2452
rect 9344 2409 9788 2435
rect 9344 2407 9512 2409
rect 7724 2270 7757 2330
rect 7526 2263 7694 2265
rect 7250 2237 7694 2263
rect 7526 2236 7694 2237
rect 7723 2259 7760 2270
rect 7723 2240 7729 2259
rect 7752 2240 7760 2259
rect 6187 2196 6223 2197
rect 6035 2166 6044 2186
rect 6064 2166 6072 2186
rect 5923 2157 5979 2159
rect 5923 2156 5960 2157
rect 6035 2156 6072 2166
rect 6131 2186 6279 2196
rect 6379 2193 6475 2195
rect 6131 2166 6140 2186
rect 6160 2166 6250 2186
rect 6270 2166 6279 2186
rect 6131 2157 6279 2166
rect 6337 2186 6475 2193
rect 6337 2166 6346 2186
rect 6366 2166 6475 2186
rect 6337 2157 6475 2166
rect 6131 2156 6168 2157
rect 6187 2105 6223 2157
rect 6242 2156 6279 2157
rect 6338 2156 6375 2157
rect 5658 2103 5699 2104
rect 4484 2053 5116 2060
rect 4484 2051 4546 2053
rect 4062 2041 4230 2042
rect 4484 2041 4506 2051
rect 3777 2016 3814 2017
rect 3727 2007 3814 2016
rect 3727 1987 3785 2007
rect 3805 1987 3814 2007
rect 3727 1977 3814 1987
rect 3873 2007 3910 2017
rect 3873 1987 3881 2007
rect 3901 1987 3910 2007
rect 3727 1976 3758 1977
rect 3873 1916 3910 1987
rect 3660 1892 3910 1916
rect 4062 2015 4506 2041
rect 4062 2013 4230 2015
rect 4062 1835 4089 2013
rect 4129 1975 4193 1987
rect 4469 1983 4506 2015
rect 4677 2014 4926 2036
rect 4677 1983 4714 2014
rect 4890 2012 4926 2014
rect 4890 1983 4927 2012
rect 4129 1974 4164 1975
rect 4106 1969 4164 1974
rect 4106 1949 4109 1969
rect 4129 1955 4164 1969
rect 4184 1955 4193 1975
rect 4129 1947 4193 1955
rect 4155 1946 4193 1947
rect 4156 1945 4193 1946
rect 4259 1979 4295 1980
rect 4367 1979 4403 1980
rect 4259 1971 4403 1979
rect 4259 1951 4267 1971
rect 4287 1951 4316 1971
rect 4259 1950 4316 1951
rect 4338 1951 4375 1971
rect 4395 1951 4403 1971
rect 4338 1950 4403 1951
rect 4259 1945 4403 1950
rect 4469 1975 4507 1983
rect 4575 1979 4611 1980
rect 4469 1955 4478 1975
rect 4498 1955 4507 1975
rect 4469 1946 4507 1955
rect 4526 1972 4611 1979
rect 4526 1952 4533 1972
rect 4554 1971 4611 1972
rect 4554 1952 4583 1971
rect 4526 1951 4583 1952
rect 4603 1951 4611 1971
rect 4469 1945 4506 1946
rect 4526 1945 4611 1951
rect 4677 1975 4715 1983
rect 4788 1979 4824 1980
rect 4677 1955 4686 1975
rect 4706 1955 4715 1975
rect 4677 1946 4715 1955
rect 4739 1971 4824 1979
rect 4739 1951 4796 1971
rect 4816 1951 4824 1971
rect 4677 1945 4714 1946
rect 4739 1945 4824 1951
rect 4890 1975 4928 1983
rect 4890 1955 4899 1975
rect 4919 1955 4928 1975
rect 4890 1946 4928 1955
rect 4890 1945 4927 1946
rect 4313 1924 4349 1945
rect 4739 1924 4770 1945
rect 4146 1920 4246 1924
rect 4146 1916 4208 1920
rect 4146 1890 4153 1916
rect 4179 1894 4208 1916
rect 4234 1894 4246 1920
rect 4179 1890 4246 1894
rect 4146 1887 4246 1890
rect 4314 1887 4349 1924
rect 4411 1921 4770 1924
rect 4411 1916 4633 1921
rect 4411 1892 4424 1916
rect 4448 1897 4633 1916
rect 4657 1897 4770 1921
rect 4448 1892 4770 1897
rect 4411 1888 4770 1892
rect 4837 1916 4986 1924
rect 4837 1896 4848 1916
rect 4868 1896 4986 1916
rect 4837 1889 4986 1896
rect 5077 1904 5116 2053
rect 5420 1939 5459 2088
rect 5550 2096 5699 2103
rect 5550 2076 5668 2096
rect 5688 2076 5699 2096
rect 5550 2068 5699 2076
rect 5766 2100 6125 2104
rect 5766 2095 6088 2100
rect 5766 2071 5879 2095
rect 5903 2076 6088 2095
rect 6112 2076 6125 2100
rect 5903 2071 6125 2076
rect 5766 2068 6125 2071
rect 6187 2068 6222 2105
rect 6290 2102 6390 2105
rect 6290 2098 6357 2102
rect 6290 2072 6302 2098
rect 6328 2076 6357 2098
rect 6383 2076 6390 2102
rect 6328 2072 6390 2076
rect 6290 2068 6390 2072
rect 5766 2047 5797 2068
rect 6187 2047 6223 2068
rect 5609 2046 5646 2047
rect 5608 2037 5646 2046
rect 5608 2017 5617 2037
rect 5637 2017 5646 2037
rect 5608 2009 5646 2017
rect 5712 2041 5797 2047
rect 5822 2046 5859 2047
rect 5712 2021 5720 2041
rect 5740 2021 5797 2041
rect 5712 2013 5797 2021
rect 5821 2037 5859 2046
rect 5821 2017 5830 2037
rect 5850 2017 5859 2037
rect 5712 2012 5748 2013
rect 5821 2009 5859 2017
rect 5925 2041 6010 2047
rect 6030 2046 6067 2047
rect 5925 2021 5933 2041
rect 5953 2040 6010 2041
rect 5953 2021 5982 2040
rect 5925 2020 5982 2021
rect 6003 2020 6010 2040
rect 5925 2013 6010 2020
rect 6029 2037 6067 2046
rect 6029 2017 6038 2037
rect 6058 2017 6067 2037
rect 5925 2012 5961 2013
rect 6029 2009 6067 2017
rect 6133 2042 6277 2047
rect 6133 2041 6198 2042
rect 6133 2021 6141 2041
rect 6161 2021 6198 2041
rect 6220 2041 6277 2042
rect 6220 2021 6249 2041
rect 6269 2021 6277 2041
rect 6133 2013 6277 2021
rect 6133 2012 6169 2013
rect 6241 2012 6277 2013
rect 6343 2046 6380 2047
rect 6343 2045 6381 2046
rect 6343 2037 6407 2045
rect 6343 2017 6352 2037
rect 6372 2023 6407 2037
rect 6427 2023 6430 2043
rect 6372 2018 6430 2023
rect 6372 2017 6407 2018
rect 5609 1980 5646 2009
rect 5610 1978 5646 1980
rect 5822 1978 5859 2009
rect 5610 1956 5859 1978
rect 6030 1977 6067 2009
rect 6343 2005 6407 2017
rect 6447 1979 6474 2157
rect 6306 1977 6474 1979
rect 6030 1951 6474 1977
rect 6626 2076 6876 2100
rect 6626 2005 6663 2076
rect 6778 2015 6809 2016
rect 6626 1985 6635 2005
rect 6655 1985 6663 2005
rect 6626 1975 6663 1985
rect 6722 2005 6809 2015
rect 6722 1985 6731 2005
rect 6751 1985 6809 2005
rect 6722 1976 6809 1985
rect 6722 1975 6759 1976
rect 6030 1941 6052 1951
rect 6306 1950 6474 1951
rect 5990 1939 6052 1941
rect 5420 1932 6052 1939
rect 4837 1888 4878 1889
rect 4161 1835 4198 1836
rect 4257 1835 4294 1836
rect 4313 1835 4349 1887
rect 4368 1835 4405 1836
rect 4061 1826 4199 1835
rect 4061 1806 4170 1826
rect 4190 1806 4199 1826
rect 2998 1802 3168 1803
rect 2998 1787 3444 1802
rect 4061 1799 4199 1806
rect 4257 1826 4405 1835
rect 4257 1806 4266 1826
rect 4286 1806 4376 1826
rect 4396 1806 4405 1826
rect 4061 1797 4157 1799
rect 3000 1776 3444 1787
rect 3000 1774 3168 1776
rect 3000 1596 3027 1774
rect 3067 1736 3131 1748
rect 3407 1744 3444 1776
rect 3615 1775 3864 1797
rect 4257 1796 4405 1806
rect 4464 1826 4501 1836
rect 4576 1835 4613 1836
rect 4557 1833 4613 1835
rect 4464 1806 4472 1826
rect 4492 1806 4501 1826
rect 4313 1795 4349 1796
rect 3615 1744 3652 1775
rect 3828 1773 3864 1775
rect 3828 1744 3865 1773
rect 3067 1735 3102 1736
rect 3044 1730 3102 1735
rect 3044 1710 3047 1730
rect 3067 1716 3102 1730
rect 3122 1716 3131 1736
rect 3067 1708 3131 1716
rect 3093 1707 3131 1708
rect 3094 1706 3131 1707
rect 3197 1740 3233 1741
rect 3305 1740 3341 1741
rect 3197 1732 3341 1740
rect 3197 1712 3205 1732
rect 3225 1731 3313 1732
rect 3225 1714 3253 1731
rect 3277 1714 3313 1731
rect 3225 1712 3313 1714
rect 3333 1712 3341 1732
rect 3197 1706 3341 1712
rect 3407 1736 3445 1744
rect 3513 1740 3549 1741
rect 3407 1716 3416 1736
rect 3436 1716 3445 1736
rect 3407 1707 3445 1716
rect 3464 1733 3549 1740
rect 3464 1713 3471 1733
rect 3492 1732 3549 1733
rect 3492 1713 3521 1732
rect 3464 1712 3521 1713
rect 3541 1712 3549 1732
rect 3407 1706 3444 1707
rect 3464 1706 3549 1712
rect 3615 1736 3653 1744
rect 3726 1740 3762 1741
rect 3615 1716 3624 1736
rect 3644 1716 3653 1736
rect 3615 1707 3653 1716
rect 3677 1732 3762 1740
rect 3677 1712 3734 1732
rect 3754 1712 3762 1732
rect 3615 1706 3652 1707
rect 3677 1706 3762 1712
rect 3828 1736 3866 1744
rect 4161 1736 4198 1737
rect 4464 1736 4501 1806
rect 4526 1826 4613 1833
rect 4526 1823 4584 1826
rect 4526 1803 4531 1823
rect 4552 1806 4584 1823
rect 4604 1806 4613 1826
rect 4552 1803 4613 1806
rect 4526 1796 4613 1803
rect 4672 1826 4709 1836
rect 4672 1806 4680 1826
rect 4700 1806 4709 1826
rect 4526 1795 4557 1796
rect 3828 1716 3837 1736
rect 3857 1716 3866 1736
rect 4160 1735 4501 1736
rect 3828 1707 3866 1716
rect 4085 1730 4501 1735
rect 4085 1710 4088 1730
rect 4108 1710 4501 1730
rect 4672 1735 4709 1806
rect 4739 1835 4770 1888
rect 5077 1886 5087 1904
rect 5105 1886 5116 1904
rect 5419 1923 6052 1932
rect 6778 1923 6809 1976
rect 6839 2005 6876 2076
rect 7047 2081 7440 2101
rect 7460 2081 7463 2101
rect 7047 2076 7463 2081
rect 7047 2075 7388 2076
rect 6991 2015 7022 2016
rect 6839 1985 6848 2005
rect 6868 1985 6876 2005
rect 6839 1975 6876 1985
rect 6935 2008 7022 2015
rect 6935 2005 6996 2008
rect 6935 1985 6944 2005
rect 6964 1988 6996 2005
rect 7017 1988 7022 2008
rect 6964 1985 7022 1988
rect 6935 1978 7022 1985
rect 7047 2005 7084 2075
rect 7350 2074 7387 2075
rect 7199 2015 7235 2016
rect 7047 1985 7056 2005
rect 7076 1985 7084 2005
rect 6935 1976 6991 1978
rect 6935 1975 6972 1976
rect 7047 1975 7084 1985
rect 7143 2005 7291 2015
rect 7391 2012 7487 2014
rect 7143 1985 7152 2005
rect 7172 1985 7262 2005
rect 7282 1985 7291 2005
rect 7143 1976 7291 1985
rect 7349 2005 7487 2012
rect 7349 1985 7358 2005
rect 7378 1985 7487 2005
rect 7349 1976 7487 1985
rect 7143 1975 7180 1976
rect 7199 1924 7235 1976
rect 7254 1975 7291 1976
rect 7350 1975 7387 1976
rect 5419 1905 5429 1923
rect 5447 1922 6052 1923
rect 6670 1922 6711 1923
rect 5447 1917 5468 1922
rect 5447 1905 5459 1917
rect 6562 1915 6711 1922
rect 5419 1897 5459 1905
rect 5502 1904 5528 1905
rect 5419 1895 5456 1897
rect 5502 1886 6056 1904
rect 6562 1895 6680 1915
rect 6700 1895 6711 1915
rect 6562 1887 6711 1895
rect 6778 1919 7137 1923
rect 6778 1914 7100 1919
rect 6778 1890 6891 1914
rect 6915 1895 7100 1914
rect 7124 1895 7137 1919
rect 6915 1890 7137 1895
rect 6778 1887 7137 1890
rect 7199 1887 7234 1924
rect 7302 1921 7402 1924
rect 7302 1917 7369 1921
rect 7302 1891 7314 1917
rect 7340 1895 7369 1917
rect 7395 1895 7402 1921
rect 7340 1891 7402 1895
rect 7302 1887 7402 1891
rect 5077 1877 5114 1886
rect 4789 1835 4826 1836
rect 4739 1826 4826 1835
rect 4739 1806 4797 1826
rect 4817 1806 4826 1826
rect 4739 1796 4826 1806
rect 4885 1826 4922 1836
rect 4885 1806 4893 1826
rect 4913 1806 4922 1826
rect 5422 1827 5459 1833
rect 5502 1827 5528 1886
rect 6035 1867 6056 1886
rect 5422 1824 5528 1827
rect 5080 1811 5117 1815
rect 4739 1795 4770 1796
rect 4885 1735 4922 1806
rect 4672 1711 4922 1735
rect 5078 1805 5117 1811
rect 5078 1787 5089 1805
rect 5107 1787 5117 1805
rect 5422 1806 5431 1824
rect 5449 1810 5528 1824
rect 5613 1842 5863 1866
rect 5449 1808 5525 1810
rect 5449 1806 5459 1808
rect 5422 1796 5459 1806
rect 5078 1778 5117 1787
rect 3828 1706 3865 1707
rect 3251 1685 3287 1706
rect 3677 1685 3708 1706
rect 4464 1687 4501 1710
rect 5078 1700 5113 1778
rect 5427 1731 5458 1796
rect 5613 1771 5650 1842
rect 5765 1781 5796 1782
rect 5613 1751 5622 1771
rect 5642 1751 5650 1771
rect 5613 1741 5650 1751
rect 5709 1771 5796 1781
rect 5709 1751 5718 1771
rect 5738 1751 5796 1771
rect 5709 1742 5796 1751
rect 5709 1741 5746 1742
rect 5075 1690 5113 1700
rect 5426 1722 5463 1731
rect 5426 1704 5436 1722
rect 5454 1704 5463 1722
rect 5426 1694 5463 1704
rect 4464 1686 4634 1687
rect 5075 1686 5085 1690
rect 3084 1681 3184 1685
rect 3084 1677 3146 1681
rect 3084 1651 3091 1677
rect 3117 1655 3146 1677
rect 3172 1655 3184 1681
rect 3117 1651 3184 1655
rect 3084 1648 3184 1651
rect 3252 1648 3287 1685
rect 3349 1682 3708 1685
rect 3349 1677 3571 1682
rect 3349 1653 3362 1677
rect 3386 1658 3571 1677
rect 3595 1658 3708 1682
rect 3386 1653 3708 1658
rect 3349 1649 3708 1653
rect 3775 1677 3924 1685
rect 3775 1657 3786 1677
rect 3806 1657 3924 1677
rect 4464 1672 5085 1686
rect 5103 1672 5113 1690
rect 5765 1689 5796 1742
rect 5826 1771 5863 1842
rect 6034 1847 6427 1867
rect 6447 1847 6450 1867
rect 6778 1866 6809 1887
rect 7199 1866 7235 1887
rect 6621 1865 6658 1866
rect 6034 1842 6450 1847
rect 6620 1856 6658 1865
rect 6034 1841 6375 1842
rect 5978 1781 6009 1782
rect 5826 1751 5835 1771
rect 5855 1751 5863 1771
rect 5826 1741 5863 1751
rect 5922 1774 6009 1781
rect 5922 1771 5983 1774
rect 5922 1751 5931 1771
rect 5951 1754 5983 1771
rect 6004 1754 6009 1774
rect 5951 1751 6009 1754
rect 5922 1744 6009 1751
rect 6034 1771 6071 1841
rect 6337 1840 6374 1841
rect 6620 1836 6629 1856
rect 6649 1836 6658 1856
rect 6620 1828 6658 1836
rect 6724 1860 6809 1866
rect 6834 1865 6871 1866
rect 6724 1840 6732 1860
rect 6752 1840 6809 1860
rect 6724 1832 6809 1840
rect 6833 1856 6871 1865
rect 6833 1836 6842 1856
rect 6862 1836 6871 1856
rect 6724 1831 6760 1832
rect 6833 1828 6871 1836
rect 6937 1860 7022 1866
rect 7042 1865 7079 1866
rect 6937 1840 6945 1860
rect 6965 1859 7022 1860
rect 6965 1840 6994 1859
rect 6937 1839 6994 1840
rect 7015 1839 7022 1859
rect 6937 1832 7022 1839
rect 7041 1856 7079 1865
rect 7041 1836 7050 1856
rect 7070 1836 7079 1856
rect 6937 1831 6973 1832
rect 7041 1828 7079 1836
rect 7145 1860 7289 1866
rect 7145 1840 7153 1860
rect 7173 1840 7205 1860
rect 7229 1840 7261 1860
rect 7281 1840 7289 1860
rect 7145 1832 7289 1840
rect 7145 1831 7181 1832
rect 7253 1831 7289 1832
rect 7355 1865 7392 1866
rect 7355 1864 7393 1865
rect 7355 1856 7419 1864
rect 7355 1836 7364 1856
rect 7384 1842 7419 1856
rect 7439 1842 7442 1862
rect 7384 1837 7442 1842
rect 7384 1836 7419 1837
rect 6621 1799 6658 1828
rect 6622 1797 6658 1799
rect 6834 1797 6871 1828
rect 6186 1781 6222 1782
rect 6034 1751 6043 1771
rect 6063 1751 6071 1771
rect 5922 1742 5978 1744
rect 5922 1741 5959 1742
rect 6034 1741 6071 1751
rect 6130 1771 6278 1781
rect 6378 1778 6474 1780
rect 6130 1751 6139 1771
rect 6159 1751 6249 1771
rect 6269 1751 6278 1771
rect 6130 1742 6278 1751
rect 6336 1771 6474 1778
rect 6622 1775 6871 1797
rect 7042 1796 7079 1828
rect 7355 1824 7419 1836
rect 7459 1798 7486 1976
rect 7318 1796 7486 1798
rect 7042 1792 7486 1796
rect 6336 1751 6345 1771
rect 6365 1751 6474 1771
rect 7042 1773 7091 1792
rect 7111 1773 7486 1792
rect 7042 1770 7486 1773
rect 7318 1769 7486 1770
rect 6336 1742 6474 1751
rect 6130 1741 6167 1742
rect 6186 1690 6222 1742
rect 6241 1741 6278 1742
rect 6337 1741 6374 1742
rect 5657 1688 5698 1689
rect 4464 1666 5113 1672
rect 5549 1681 5698 1688
rect 4464 1665 5112 1666
rect 5075 1663 5112 1665
rect 3775 1650 3924 1657
rect 5549 1661 5667 1681
rect 5687 1661 5698 1681
rect 5549 1653 5698 1661
rect 5765 1685 6124 1689
rect 5765 1680 6087 1685
rect 5765 1656 5878 1680
rect 5902 1661 6087 1680
rect 6111 1661 6124 1685
rect 5902 1656 6124 1661
rect 5765 1653 6124 1656
rect 6186 1653 6221 1690
rect 6289 1687 6389 1690
rect 6289 1683 6356 1687
rect 6289 1657 6301 1683
rect 6327 1661 6356 1683
rect 6382 1661 6389 1687
rect 6327 1657 6389 1661
rect 6289 1653 6389 1657
rect 3775 1649 3816 1650
rect 3099 1596 3136 1597
rect 3195 1596 3232 1597
rect 3251 1596 3287 1648
rect 3306 1596 3343 1597
rect 2999 1587 3137 1596
rect 2999 1567 3108 1587
rect 3128 1567 3137 1587
rect 2999 1560 3137 1567
rect 3195 1587 3343 1596
rect 3195 1567 3204 1587
rect 3224 1567 3314 1587
rect 3334 1567 3343 1587
rect 2999 1558 3095 1560
rect 3195 1557 3343 1567
rect 3402 1587 3439 1597
rect 3514 1596 3551 1597
rect 3495 1594 3551 1596
rect 3402 1567 3410 1587
rect 3430 1567 3439 1587
rect 3251 1556 3287 1557
rect 3099 1497 3136 1498
rect 3402 1497 3439 1567
rect 3464 1587 3551 1594
rect 3464 1584 3522 1587
rect 3464 1564 3469 1584
rect 3490 1567 3522 1584
rect 3542 1567 3551 1587
rect 3490 1564 3551 1567
rect 3464 1557 3551 1564
rect 3610 1587 3647 1597
rect 3610 1567 3618 1587
rect 3638 1567 3647 1587
rect 3464 1556 3495 1557
rect 3098 1496 3439 1497
rect 3023 1491 3439 1496
rect 3023 1471 3026 1491
rect 3046 1471 3439 1491
rect 3610 1496 3647 1567
rect 3677 1596 3708 1649
rect 5765 1632 5796 1653
rect 6186 1632 6222 1653
rect 5429 1623 5466 1632
rect 5608 1631 5645 1632
rect 5429 1605 5438 1623
rect 5456 1605 5466 1623
rect 3727 1596 3764 1597
rect 3677 1587 3764 1596
rect 3677 1567 3735 1587
rect 3755 1567 3764 1587
rect 3677 1557 3764 1567
rect 3823 1587 3860 1597
rect 3823 1567 3831 1587
rect 3851 1567 3860 1587
rect 3677 1556 3708 1557
rect 3823 1496 3860 1567
rect 5078 1591 5115 1601
rect 5429 1595 5466 1605
rect 5078 1573 5087 1591
rect 5105 1573 5115 1591
rect 5078 1564 5115 1573
rect 5078 1540 5113 1564
rect 5430 1560 5466 1595
rect 5607 1622 5645 1631
rect 5607 1602 5616 1622
rect 5636 1602 5645 1622
rect 5607 1594 5645 1602
rect 5711 1626 5796 1632
rect 5821 1631 5858 1632
rect 5711 1606 5719 1626
rect 5739 1606 5796 1626
rect 5711 1598 5796 1606
rect 5820 1622 5858 1631
rect 5820 1602 5829 1622
rect 5849 1602 5858 1622
rect 5711 1597 5747 1598
rect 5820 1594 5858 1602
rect 5924 1626 6009 1632
rect 6029 1631 6066 1632
rect 5924 1606 5932 1626
rect 5952 1625 6009 1626
rect 5952 1606 5981 1625
rect 5924 1605 5981 1606
rect 6002 1605 6009 1625
rect 5924 1598 6009 1605
rect 6028 1622 6066 1631
rect 6028 1602 6037 1622
rect 6057 1602 6066 1622
rect 5924 1597 5960 1598
rect 6028 1594 6066 1602
rect 6132 1626 6276 1632
rect 6132 1606 6140 1626
rect 6160 1625 6248 1626
rect 6160 1606 6188 1625
rect 6132 1604 6188 1606
rect 6210 1606 6248 1625
rect 6268 1606 6276 1626
rect 6210 1604 6276 1606
rect 6132 1598 6276 1604
rect 6132 1597 6168 1598
rect 6240 1597 6276 1598
rect 6342 1631 6379 1632
rect 6342 1630 6380 1631
rect 6342 1622 6406 1630
rect 6342 1602 6351 1622
rect 6371 1608 6406 1622
rect 6426 1608 6429 1628
rect 6371 1603 6429 1608
rect 6371 1602 6406 1603
rect 5608 1565 5645 1594
rect 5076 1516 5113 1540
rect 5075 1510 5113 1516
rect 3610 1472 3860 1496
rect 4486 1492 5113 1510
rect 4068 1475 4236 1476
rect 4487 1475 4511 1492
rect 4068 1449 4512 1475
rect 4068 1447 4236 1449
rect 4068 1269 4095 1447
rect 4135 1409 4199 1421
rect 4475 1417 4512 1449
rect 4683 1448 4932 1470
rect 4683 1417 4720 1448
rect 4896 1446 4932 1448
rect 5075 1451 5113 1492
rect 5428 1519 5466 1560
rect 5609 1563 5645 1565
rect 5821 1563 5858 1594
rect 5609 1541 5858 1563
rect 6029 1562 6066 1594
rect 6342 1590 6406 1602
rect 6446 1564 6473 1742
rect 6305 1562 6473 1564
rect 6029 1536 6473 1562
rect 6030 1519 6054 1536
rect 6305 1535 6473 1536
rect 5428 1501 6055 1519
rect 6681 1515 6931 1539
rect 5428 1495 5466 1501
rect 5428 1471 5465 1495
rect 4896 1417 4933 1446
rect 4135 1408 4170 1409
rect 4112 1403 4170 1408
rect 4112 1383 4115 1403
rect 4135 1389 4170 1403
rect 4190 1389 4199 1409
rect 4135 1381 4199 1389
rect 4161 1380 4199 1381
rect 4162 1379 4199 1380
rect 4265 1413 4301 1414
rect 4373 1413 4409 1414
rect 4265 1407 4409 1413
rect 4265 1405 4331 1407
rect 4265 1385 4273 1405
rect 4293 1386 4331 1405
rect 4353 1405 4409 1407
rect 4353 1386 4381 1405
rect 4293 1385 4381 1386
rect 4401 1385 4409 1405
rect 4265 1379 4409 1385
rect 4475 1409 4513 1417
rect 4581 1413 4617 1414
rect 4475 1389 4484 1409
rect 4504 1389 4513 1409
rect 4475 1380 4513 1389
rect 4532 1406 4617 1413
rect 4532 1386 4539 1406
rect 4560 1405 4617 1406
rect 4560 1386 4589 1405
rect 4532 1385 4589 1386
rect 4609 1385 4617 1405
rect 4475 1379 4512 1380
rect 4532 1379 4617 1385
rect 4683 1409 4721 1417
rect 4794 1413 4830 1414
rect 4683 1389 4692 1409
rect 4712 1389 4721 1409
rect 4683 1380 4721 1389
rect 4745 1405 4830 1413
rect 4745 1385 4802 1405
rect 4822 1385 4830 1405
rect 4683 1379 4720 1380
rect 4745 1379 4830 1385
rect 4896 1409 4934 1417
rect 4896 1389 4905 1409
rect 4925 1389 4934 1409
rect 4896 1380 4934 1389
rect 5075 1416 5111 1451
rect 5428 1447 5463 1471
rect 5426 1438 5463 1447
rect 5426 1420 5436 1438
rect 5454 1420 5463 1438
rect 5075 1406 5112 1416
rect 5426 1410 5463 1420
rect 6681 1444 6718 1515
rect 6833 1454 6864 1455
rect 6681 1424 6690 1444
rect 6710 1424 6718 1444
rect 6681 1414 6718 1424
rect 6777 1444 6864 1454
rect 6777 1424 6786 1444
rect 6806 1424 6864 1444
rect 6777 1415 6864 1424
rect 6777 1414 6814 1415
rect 5075 1388 5085 1406
rect 5103 1388 5112 1406
rect 4896 1379 4933 1380
rect 5075 1379 5112 1388
rect 4319 1358 4355 1379
rect 4745 1358 4776 1379
rect 6833 1362 6864 1415
rect 6894 1444 6931 1515
rect 7102 1520 7495 1540
rect 7515 1520 7518 1540
rect 7102 1515 7518 1520
rect 7102 1514 7443 1515
rect 7046 1454 7077 1455
rect 6894 1424 6903 1444
rect 6923 1424 6931 1444
rect 6894 1414 6931 1424
rect 6990 1447 7077 1454
rect 6990 1444 7051 1447
rect 6990 1424 6999 1444
rect 7019 1427 7051 1444
rect 7072 1427 7077 1447
rect 7019 1424 7077 1427
rect 6990 1417 7077 1424
rect 7102 1444 7139 1514
rect 7405 1513 7442 1514
rect 7254 1454 7290 1455
rect 7102 1424 7111 1444
rect 7131 1424 7139 1444
rect 6990 1415 7046 1417
rect 6990 1414 7027 1415
rect 7102 1414 7139 1424
rect 7198 1444 7346 1454
rect 7446 1451 7542 1453
rect 7198 1424 7207 1444
rect 7227 1424 7317 1444
rect 7337 1424 7346 1444
rect 7198 1415 7346 1424
rect 7404 1444 7542 1451
rect 7404 1424 7413 1444
rect 7433 1424 7542 1444
rect 7404 1415 7542 1424
rect 7198 1414 7235 1415
rect 7254 1363 7290 1415
rect 7309 1414 7346 1415
rect 7405 1414 7442 1415
rect 6725 1361 6766 1362
rect 4152 1354 4252 1358
rect 4152 1350 4214 1354
rect 4152 1324 4159 1350
rect 4185 1328 4214 1350
rect 4240 1328 4252 1354
rect 4185 1324 4252 1328
rect 4152 1321 4252 1324
rect 4320 1321 4355 1358
rect 4417 1355 4776 1358
rect 4417 1350 4639 1355
rect 4417 1326 4430 1350
rect 4454 1331 4639 1350
rect 4663 1331 4776 1355
rect 4454 1326 4776 1331
rect 4417 1322 4776 1326
rect 4843 1350 4992 1358
rect 4843 1330 4854 1350
rect 4874 1330 4992 1350
rect 6617 1354 6766 1361
rect 5429 1346 5466 1348
rect 5429 1345 6077 1346
rect 4843 1323 4992 1330
rect 5428 1339 6077 1345
rect 4843 1322 4884 1323
rect 4167 1269 4204 1270
rect 4263 1269 4300 1270
rect 4319 1269 4355 1321
rect 4374 1269 4411 1270
rect 4067 1260 4205 1269
rect 2323 1251 2355 1256
rect 1103 1233 1199 1235
rect 855 1206 864 1226
rect 884 1206 974 1226
rect 994 1206 1003 1226
rect 855 1197 1003 1206
rect 1061 1226 1199 1233
rect 1816 1230 2262 1245
rect 2092 1229 2262 1230
rect 1061 1206 1070 1226
rect 1090 1206 1199 1226
rect 1061 1197 1199 1206
rect 855 1196 892 1197
rect 911 1145 947 1197
rect 966 1196 1003 1197
rect 1062 1196 1099 1197
rect 382 1143 423 1144
rect 144 979 183 1128
rect 274 1136 423 1143
rect 274 1116 392 1136
rect 412 1116 423 1136
rect 274 1108 423 1116
rect 490 1140 849 1144
rect 490 1135 812 1140
rect 490 1111 603 1135
rect 627 1116 812 1135
rect 836 1116 849 1140
rect 627 1111 849 1116
rect 490 1108 849 1111
rect 911 1108 946 1145
rect 1014 1142 1114 1145
rect 1014 1138 1081 1142
rect 1014 1112 1026 1138
rect 1052 1116 1081 1138
rect 1107 1116 1114 1142
rect 1052 1112 1114 1116
rect 1014 1108 1114 1112
rect 490 1087 521 1108
rect 911 1087 947 1108
rect 333 1086 370 1087
rect 332 1077 370 1086
rect 332 1057 341 1077
rect 361 1057 370 1077
rect 332 1049 370 1057
rect 436 1081 521 1087
rect 546 1086 583 1087
rect 436 1061 444 1081
rect 464 1061 521 1081
rect 436 1053 521 1061
rect 545 1077 583 1086
rect 545 1057 554 1077
rect 574 1057 583 1077
rect 436 1052 472 1053
rect 545 1049 583 1057
rect 649 1081 734 1087
rect 754 1086 791 1087
rect 649 1061 657 1081
rect 677 1080 734 1081
rect 677 1061 706 1080
rect 649 1060 706 1061
rect 727 1060 734 1080
rect 649 1053 734 1060
rect 753 1077 791 1086
rect 753 1057 762 1077
rect 782 1057 791 1077
rect 649 1052 685 1053
rect 753 1049 791 1057
rect 857 1082 1001 1087
rect 857 1081 922 1082
rect 857 1061 865 1081
rect 885 1061 922 1081
rect 944 1081 1001 1082
rect 944 1061 973 1081
rect 993 1061 1001 1081
rect 857 1053 1001 1061
rect 857 1052 893 1053
rect 965 1052 1001 1053
rect 1067 1086 1104 1087
rect 1067 1085 1105 1086
rect 1067 1077 1131 1085
rect 1067 1057 1076 1077
rect 1096 1063 1131 1077
rect 1151 1063 1154 1083
rect 1096 1058 1154 1063
rect 1096 1057 1131 1058
rect 333 1020 370 1049
rect 334 1018 370 1020
rect 546 1018 583 1049
rect 334 996 583 1018
rect 754 1017 791 1049
rect 1067 1045 1131 1057
rect 1171 1019 1198 1197
rect 1030 1017 1198 1019
rect 754 991 1198 1017
rect 1350 1116 1600 1140
rect 1350 1045 1387 1116
rect 1502 1055 1533 1056
rect 1350 1025 1359 1045
rect 1379 1025 1387 1045
rect 1350 1015 1387 1025
rect 1446 1045 1533 1055
rect 1446 1025 1455 1045
rect 1475 1025 1533 1045
rect 1446 1016 1533 1025
rect 1446 1015 1483 1016
rect 754 981 776 991
rect 1030 990 1198 991
rect 714 979 776 981
rect 144 972 776 979
rect 143 963 776 972
rect 1502 963 1533 1016
rect 1563 1045 1600 1116
rect 1771 1121 2164 1141
rect 2184 1121 2187 1141
rect 1771 1116 2187 1121
rect 1771 1115 2112 1116
rect 1715 1055 1746 1056
rect 1563 1025 1572 1045
rect 1592 1025 1600 1045
rect 1563 1015 1600 1025
rect 1659 1048 1746 1055
rect 1659 1045 1720 1048
rect 1659 1025 1668 1045
rect 1688 1028 1720 1045
rect 1741 1028 1746 1048
rect 1688 1025 1746 1028
rect 1659 1018 1746 1025
rect 1771 1045 1808 1115
rect 2074 1114 2111 1115
rect 1923 1055 1959 1056
rect 1771 1025 1780 1045
rect 1800 1025 1808 1045
rect 1659 1016 1715 1018
rect 1659 1015 1696 1016
rect 1771 1015 1808 1025
rect 1867 1045 2015 1055
rect 2115 1052 2211 1054
rect 1867 1025 1876 1045
rect 1896 1025 1986 1045
rect 2006 1025 2015 1045
rect 1867 1016 2015 1025
rect 2073 1045 2211 1052
rect 2073 1025 2082 1045
rect 2102 1025 2211 1045
rect 2073 1016 2211 1025
rect 1867 1015 1904 1016
rect 1923 964 1959 1016
rect 1978 1015 2015 1016
rect 2074 1015 2111 1016
rect 143 945 153 963
rect 171 962 776 963
rect 1394 962 1435 963
rect 171 957 192 962
rect 171 945 183 957
rect 1286 955 1435 962
rect 143 937 183 945
rect 226 944 252 945
rect 143 935 180 937
rect 226 926 780 944
rect 1286 935 1404 955
rect 1424 935 1435 955
rect 1286 927 1435 935
rect 1502 959 1861 963
rect 1502 954 1824 959
rect 1502 930 1615 954
rect 1639 935 1824 954
rect 1848 935 1861 959
rect 1639 930 1861 935
rect 1502 927 1861 930
rect 1923 927 1958 964
rect 2026 961 2126 964
rect 2026 957 2093 961
rect 2026 931 2038 957
rect 2064 935 2093 957
rect 2119 935 2126 961
rect 2064 931 2126 935
rect 2026 927 2126 931
rect 146 867 183 873
rect 226 867 252 926
rect 759 907 780 926
rect 146 864 252 867
rect 146 846 155 864
rect 173 850 252 864
rect 337 882 587 906
rect 173 848 249 850
rect 173 846 183 848
rect 146 836 183 846
rect 151 771 182 836
rect 337 811 374 882
rect 489 821 520 822
rect 337 791 346 811
rect 366 791 374 811
rect 337 781 374 791
rect 433 811 520 821
rect 433 791 442 811
rect 462 791 520 811
rect 433 782 520 791
rect 433 781 470 782
rect 150 762 187 771
rect 150 744 160 762
rect 178 744 187 762
rect 150 734 187 744
rect 489 729 520 782
rect 550 811 587 882
rect 758 887 1151 907
rect 1171 887 1174 907
rect 1502 906 1533 927
rect 1923 906 1959 927
rect 1345 905 1382 906
rect 758 882 1174 887
rect 1344 896 1382 905
rect 758 881 1099 882
rect 702 821 733 822
rect 550 791 559 811
rect 579 791 587 811
rect 550 781 587 791
rect 646 814 733 821
rect 646 811 707 814
rect 646 791 655 811
rect 675 794 707 811
rect 728 794 733 814
rect 675 791 733 794
rect 646 784 733 791
rect 758 811 795 881
rect 1061 880 1098 881
rect 1344 876 1353 896
rect 1373 876 1382 896
rect 1344 868 1382 876
rect 1448 900 1533 906
rect 1558 905 1595 906
rect 1448 880 1456 900
rect 1476 880 1533 900
rect 1448 872 1533 880
rect 1557 896 1595 905
rect 1557 876 1566 896
rect 1586 876 1595 896
rect 1448 871 1484 872
rect 1557 868 1595 876
rect 1661 900 1746 906
rect 1766 905 1803 906
rect 1661 880 1669 900
rect 1689 899 1746 900
rect 1689 880 1718 899
rect 1661 879 1718 880
rect 1739 879 1746 899
rect 1661 872 1746 879
rect 1765 896 1803 905
rect 1765 876 1774 896
rect 1794 876 1803 896
rect 1661 871 1697 872
rect 1765 868 1803 876
rect 1869 901 2013 906
rect 1869 900 1928 901
rect 1869 880 1877 900
rect 1897 881 1928 900
rect 1952 900 2013 901
rect 1952 881 1985 900
rect 1897 880 1985 881
rect 2005 880 2013 900
rect 1869 872 2013 880
rect 1869 871 1905 872
rect 1977 871 2013 872
rect 2079 905 2116 906
rect 2079 904 2117 905
rect 2079 896 2143 904
rect 2079 876 2088 896
rect 2108 882 2143 896
rect 2163 882 2166 902
rect 2108 877 2166 882
rect 2108 876 2143 877
rect 1345 839 1382 868
rect 1346 837 1382 839
rect 1558 837 1595 868
rect 910 821 946 822
rect 758 791 767 811
rect 787 791 795 811
rect 646 782 702 784
rect 646 781 683 782
rect 758 781 795 791
rect 854 811 1002 821
rect 1102 818 1198 820
rect 854 791 863 811
rect 883 791 973 811
rect 993 791 1002 811
rect 854 782 1002 791
rect 1060 811 1198 818
rect 1346 815 1595 837
rect 1766 836 1803 868
rect 2079 864 2143 876
rect 2183 838 2210 1016
rect 2042 836 2210 838
rect 1766 832 2210 836
rect 1060 791 1069 811
rect 1089 791 1198 811
rect 1766 813 1815 832
rect 1835 813 2210 832
rect 1766 810 2210 813
rect 2042 809 2210 810
rect 2231 835 2262 1229
rect 2323 1233 2328 1251
rect 2348 1233 2355 1251
rect 2323 1228 2355 1233
rect 2326 1226 2355 1228
rect 3055 1241 3223 1242
rect 3055 1238 3499 1241
rect 3055 1219 3430 1238
rect 3450 1219 3499 1238
rect 4067 1240 4176 1260
rect 4196 1240 4205 1260
rect 3055 1215 3499 1219
rect 3055 1213 3223 1215
rect 3055 1035 3082 1213
rect 3122 1175 3186 1187
rect 3462 1183 3499 1215
rect 3670 1214 3919 1236
rect 4067 1233 4205 1240
rect 4263 1260 4411 1269
rect 4263 1240 4272 1260
rect 4292 1240 4382 1260
rect 4402 1240 4411 1260
rect 4067 1231 4163 1233
rect 4263 1230 4411 1240
rect 4470 1260 4507 1270
rect 4582 1269 4619 1270
rect 4563 1267 4619 1269
rect 4470 1240 4478 1260
rect 4498 1240 4507 1260
rect 4319 1229 4355 1230
rect 3670 1183 3707 1214
rect 3883 1212 3919 1214
rect 3883 1183 3920 1212
rect 3122 1174 3157 1175
rect 3099 1169 3157 1174
rect 3099 1149 3102 1169
rect 3122 1155 3157 1169
rect 3177 1155 3186 1175
rect 3122 1147 3186 1155
rect 3148 1146 3186 1147
rect 3149 1145 3186 1146
rect 3252 1179 3288 1180
rect 3360 1179 3396 1180
rect 3252 1171 3396 1179
rect 3252 1151 3260 1171
rect 3280 1151 3312 1171
rect 3336 1151 3368 1171
rect 3388 1151 3396 1171
rect 3252 1145 3396 1151
rect 3462 1175 3500 1183
rect 3568 1179 3604 1180
rect 3462 1155 3471 1175
rect 3491 1155 3500 1175
rect 3462 1146 3500 1155
rect 3519 1172 3604 1179
rect 3519 1152 3526 1172
rect 3547 1171 3604 1172
rect 3547 1152 3576 1171
rect 3519 1151 3576 1152
rect 3596 1151 3604 1171
rect 3462 1145 3499 1146
rect 3519 1145 3604 1151
rect 3670 1175 3708 1183
rect 3781 1179 3817 1180
rect 3670 1155 3679 1175
rect 3699 1155 3708 1175
rect 3670 1146 3708 1155
rect 3732 1171 3817 1179
rect 3732 1151 3789 1171
rect 3809 1151 3817 1171
rect 3670 1145 3707 1146
rect 3732 1145 3817 1151
rect 3883 1175 3921 1183
rect 3883 1155 3892 1175
rect 3912 1155 3921 1175
rect 4167 1170 4204 1171
rect 4470 1170 4507 1240
rect 4532 1260 4619 1267
rect 4532 1257 4590 1260
rect 4532 1237 4537 1257
rect 4558 1240 4590 1257
rect 4610 1240 4619 1260
rect 4558 1237 4619 1240
rect 4532 1230 4619 1237
rect 4678 1260 4715 1270
rect 4678 1240 4686 1260
rect 4706 1240 4715 1260
rect 4532 1229 4563 1230
rect 4166 1169 4507 1170
rect 3883 1146 3921 1155
rect 4091 1164 4507 1169
rect 3883 1145 3920 1146
rect 3306 1124 3342 1145
rect 3732 1124 3763 1145
rect 4091 1144 4094 1164
rect 4114 1144 4507 1164
rect 4678 1169 4715 1240
rect 4745 1269 4776 1322
rect 5428 1321 5438 1339
rect 5456 1325 6077 1339
rect 6617 1334 6735 1354
rect 6755 1334 6766 1354
rect 6617 1326 6766 1334
rect 6833 1358 7192 1362
rect 6833 1353 7155 1358
rect 6833 1329 6946 1353
rect 6970 1334 7155 1353
rect 7179 1334 7192 1358
rect 6970 1329 7192 1334
rect 6833 1326 7192 1329
rect 7254 1326 7289 1363
rect 7357 1360 7457 1363
rect 7357 1356 7424 1360
rect 7357 1330 7369 1356
rect 7395 1334 7424 1356
rect 7450 1334 7457 1360
rect 7395 1330 7457 1334
rect 7357 1326 7457 1330
rect 5456 1321 5466 1325
rect 5907 1324 6077 1325
rect 5078 1307 5115 1317
rect 5078 1289 5087 1307
rect 5105 1289 5115 1307
rect 5078 1280 5115 1289
rect 5428 1311 5466 1321
rect 4795 1269 4832 1270
rect 4745 1260 4832 1269
rect 4745 1240 4803 1260
rect 4823 1240 4832 1260
rect 4745 1230 4832 1240
rect 4891 1260 4928 1270
rect 4891 1240 4899 1260
rect 4919 1240 4928 1260
rect 4745 1229 4776 1230
rect 4891 1169 4928 1240
rect 5083 1215 5114 1280
rect 5428 1233 5463 1311
rect 6040 1301 6077 1324
rect 6833 1305 6864 1326
rect 7254 1305 7290 1326
rect 6676 1304 6713 1305
rect 5424 1224 5463 1233
rect 5082 1205 5119 1215
rect 5082 1203 5092 1205
rect 5016 1201 5092 1203
rect 4678 1145 4928 1169
rect 5013 1187 5092 1201
rect 5110 1187 5119 1205
rect 5424 1206 5434 1224
rect 5452 1206 5463 1224
rect 5424 1200 5463 1206
rect 5619 1276 5869 1300
rect 5619 1205 5656 1276
rect 5771 1215 5802 1216
rect 5424 1196 5461 1200
rect 5013 1184 5119 1187
rect 4485 1125 4506 1144
rect 5013 1125 5039 1184
rect 5082 1178 5119 1184
rect 5619 1185 5628 1205
rect 5648 1185 5656 1205
rect 5619 1175 5656 1185
rect 5715 1205 5802 1215
rect 5715 1185 5724 1205
rect 5744 1185 5802 1205
rect 5715 1176 5802 1185
rect 5715 1175 5752 1176
rect 5427 1125 5464 1134
rect 3139 1120 3239 1124
rect 3139 1116 3201 1120
rect 3139 1090 3146 1116
rect 3172 1094 3201 1116
rect 3227 1094 3239 1120
rect 3172 1090 3239 1094
rect 3139 1087 3239 1090
rect 3307 1087 3342 1124
rect 3404 1121 3763 1124
rect 3404 1116 3626 1121
rect 3404 1092 3417 1116
rect 3441 1097 3626 1116
rect 3650 1097 3763 1121
rect 3441 1092 3763 1097
rect 3404 1088 3763 1092
rect 3830 1116 3979 1124
rect 3830 1096 3841 1116
rect 3861 1096 3979 1116
rect 4485 1107 5039 1125
rect 5085 1114 5122 1116
rect 5013 1106 5039 1107
rect 5082 1106 5122 1114
rect 3830 1089 3979 1096
rect 5082 1094 5094 1106
rect 5073 1089 5094 1094
rect 3830 1088 3871 1089
rect 4489 1088 5094 1089
rect 5112 1088 5122 1106
rect 3154 1035 3191 1036
rect 3250 1035 3287 1036
rect 3306 1035 3342 1087
rect 3361 1035 3398 1036
rect 3054 1026 3192 1035
rect 3054 1006 3163 1026
rect 3183 1006 3192 1026
rect 3054 999 3192 1006
rect 3250 1026 3398 1035
rect 3250 1006 3259 1026
rect 3279 1006 3369 1026
rect 3389 1006 3398 1026
rect 3054 997 3150 999
rect 3250 996 3398 1006
rect 3457 1026 3494 1036
rect 3569 1035 3606 1036
rect 3550 1033 3606 1035
rect 3457 1006 3465 1026
rect 3485 1006 3494 1026
rect 3306 995 3342 996
rect 3154 936 3191 937
rect 3457 936 3494 1006
rect 3519 1026 3606 1033
rect 3519 1023 3577 1026
rect 3519 1003 3524 1023
rect 3545 1006 3577 1023
rect 3597 1006 3606 1026
rect 3545 1003 3606 1006
rect 3519 996 3606 1003
rect 3665 1026 3702 1036
rect 3665 1006 3673 1026
rect 3693 1006 3702 1026
rect 3519 995 3550 996
rect 3153 935 3494 936
rect 3078 930 3494 935
rect 3078 910 3081 930
rect 3101 910 3494 930
rect 3665 935 3702 1006
rect 3732 1035 3763 1088
rect 4489 1079 5122 1088
rect 5425 1107 5436 1125
rect 5454 1107 5464 1125
rect 5771 1123 5802 1176
rect 5832 1205 5869 1276
rect 6040 1281 6433 1301
rect 6453 1281 6456 1301
rect 6040 1276 6456 1281
rect 6675 1295 6713 1304
rect 6040 1275 6381 1276
rect 6675 1275 6684 1295
rect 6704 1275 6713 1295
rect 5984 1215 6015 1216
rect 5832 1185 5841 1205
rect 5861 1185 5869 1205
rect 5832 1175 5869 1185
rect 5928 1208 6015 1215
rect 5928 1205 5989 1208
rect 5928 1185 5937 1205
rect 5957 1188 5989 1205
rect 6010 1188 6015 1208
rect 5957 1185 6015 1188
rect 5928 1178 6015 1185
rect 6040 1205 6077 1275
rect 6343 1274 6380 1275
rect 6675 1267 6713 1275
rect 6779 1299 6864 1305
rect 6889 1304 6926 1305
rect 6779 1279 6787 1299
rect 6807 1279 6864 1299
rect 6779 1271 6864 1279
rect 6888 1295 6926 1304
rect 6888 1275 6897 1295
rect 6917 1275 6926 1295
rect 6779 1270 6815 1271
rect 6888 1267 6926 1275
rect 6992 1299 7077 1305
rect 7097 1304 7134 1305
rect 6992 1279 7000 1299
rect 7020 1298 7077 1299
rect 7020 1279 7049 1298
rect 6992 1278 7049 1279
rect 7070 1278 7077 1298
rect 6992 1271 7077 1278
rect 7096 1295 7134 1304
rect 7096 1275 7105 1295
rect 7125 1275 7134 1295
rect 6992 1270 7028 1271
rect 7096 1267 7134 1275
rect 7200 1299 7344 1305
rect 7200 1279 7208 1299
rect 7228 1298 7316 1299
rect 7228 1279 7261 1298
rect 7284 1279 7316 1298
rect 7336 1279 7344 1299
rect 7200 1271 7344 1279
rect 7200 1270 7236 1271
rect 7308 1270 7344 1271
rect 7410 1304 7447 1305
rect 7410 1303 7448 1304
rect 7410 1295 7474 1303
rect 7410 1275 7419 1295
rect 7439 1281 7474 1295
rect 7494 1281 7497 1301
rect 7439 1276 7497 1281
rect 7439 1275 7474 1276
rect 6676 1238 6713 1267
rect 6677 1236 6713 1238
rect 6889 1236 6926 1267
rect 6192 1215 6228 1216
rect 6040 1185 6049 1205
rect 6069 1185 6077 1205
rect 5928 1176 5984 1178
rect 5928 1175 5965 1176
rect 6040 1175 6077 1185
rect 6136 1205 6284 1215
rect 6677 1214 6926 1236
rect 7097 1235 7134 1267
rect 7410 1263 7474 1275
rect 7514 1237 7541 1415
rect 7373 1235 7541 1237
rect 7097 1224 7541 1235
rect 7604 1235 7634 2236
rect 7723 2229 7760 2240
rect 9344 2229 9371 2407
rect 9411 2369 9475 2381
rect 9751 2377 9788 2409
rect 9959 2408 10208 2430
rect 9959 2377 9996 2408
rect 10172 2406 10208 2408
rect 10351 2411 10389 2452
rect 10801 2448 10838 2457
rect 10801 2430 10811 2448
rect 10829 2430 10838 2448
rect 10801 2420 10838 2430
rect 12366 2419 12397 2472
rect 12427 2501 12464 2572
rect 12635 2577 13028 2597
rect 13048 2577 13051 2597
rect 12635 2572 13051 2577
rect 12635 2571 12976 2572
rect 12579 2511 12610 2512
rect 12427 2481 12436 2501
rect 12456 2481 12464 2501
rect 12427 2471 12464 2481
rect 12523 2504 12610 2511
rect 12523 2501 12584 2504
rect 12523 2481 12532 2501
rect 12552 2484 12584 2501
rect 12605 2484 12610 2504
rect 12552 2481 12610 2484
rect 12523 2474 12610 2481
rect 12635 2501 12672 2571
rect 12938 2570 12975 2571
rect 12787 2511 12823 2512
rect 12635 2481 12644 2501
rect 12664 2481 12672 2501
rect 12523 2472 12579 2474
rect 12523 2471 12560 2472
rect 12635 2471 12672 2481
rect 12731 2501 12879 2511
rect 12979 2508 13075 2510
rect 12731 2481 12740 2501
rect 12760 2481 12850 2501
rect 12870 2481 12879 2501
rect 12731 2472 12879 2481
rect 12937 2501 13075 2508
rect 12937 2481 12946 2501
rect 12966 2481 13075 2501
rect 12937 2472 13075 2481
rect 12731 2471 12768 2472
rect 12787 2420 12823 2472
rect 12842 2471 12879 2472
rect 12938 2471 12975 2472
rect 12258 2418 12299 2419
rect 12150 2411 12299 2418
rect 10172 2377 10209 2406
rect 9411 2368 9446 2369
rect 9388 2363 9446 2368
rect 9388 2343 9391 2363
rect 9411 2349 9446 2363
rect 9466 2349 9475 2369
rect 9411 2341 9475 2349
rect 9437 2340 9475 2341
rect 9438 2339 9475 2340
rect 9541 2373 9577 2374
rect 9649 2373 9685 2374
rect 9541 2367 9685 2373
rect 9541 2365 9607 2367
rect 9541 2345 9549 2365
rect 9569 2346 9607 2365
rect 9629 2365 9685 2367
rect 9629 2346 9657 2365
rect 9569 2345 9657 2346
rect 9677 2345 9685 2365
rect 9541 2339 9685 2345
rect 9751 2369 9789 2377
rect 9857 2373 9893 2374
rect 9751 2349 9760 2369
rect 9780 2349 9789 2369
rect 9751 2340 9789 2349
rect 9808 2366 9893 2373
rect 9808 2346 9815 2366
rect 9836 2365 9893 2366
rect 9836 2346 9865 2365
rect 9808 2345 9865 2346
rect 9885 2345 9893 2365
rect 9751 2339 9788 2340
rect 9808 2339 9893 2345
rect 9959 2369 9997 2377
rect 10070 2373 10106 2374
rect 9959 2349 9968 2369
rect 9988 2349 9997 2369
rect 9959 2340 9997 2349
rect 10021 2365 10106 2373
rect 10021 2345 10078 2365
rect 10098 2345 10106 2365
rect 9959 2339 9996 2340
rect 10021 2339 10106 2345
rect 10172 2369 10210 2377
rect 10172 2349 10181 2369
rect 10201 2349 10210 2369
rect 10172 2340 10210 2349
rect 10351 2376 10387 2411
rect 12150 2391 12268 2411
rect 12288 2391 12299 2411
rect 12150 2383 12299 2391
rect 12366 2415 12725 2419
rect 12366 2410 12688 2415
rect 12366 2386 12479 2410
rect 12503 2391 12688 2410
rect 12712 2391 12725 2415
rect 12503 2386 12725 2391
rect 12366 2383 12725 2386
rect 12787 2383 12822 2420
rect 12890 2417 12990 2420
rect 12890 2413 12957 2417
rect 12890 2387 12902 2413
rect 12928 2391 12957 2413
rect 12983 2391 12990 2417
rect 12928 2387 12990 2391
rect 12890 2383 12990 2387
rect 10351 2366 10388 2376
rect 10351 2348 10361 2366
rect 10379 2348 10388 2366
rect 12366 2362 12397 2383
rect 12787 2362 12823 2383
rect 12209 2361 12246 2362
rect 10804 2356 10841 2358
rect 10804 2355 11452 2356
rect 10172 2339 10209 2340
rect 10351 2339 10388 2348
rect 10803 2349 11452 2355
rect 9595 2318 9631 2339
rect 10021 2318 10052 2339
rect 10803 2331 10813 2349
rect 10831 2335 11452 2349
rect 10831 2331 10841 2335
rect 11282 2334 11452 2335
rect 10803 2321 10841 2331
rect 9428 2314 9528 2318
rect 9428 2310 9490 2314
rect 9428 2284 9435 2310
rect 9461 2288 9490 2310
rect 9516 2288 9528 2314
rect 9461 2284 9528 2288
rect 9428 2281 9528 2284
rect 9596 2281 9631 2318
rect 9693 2315 10052 2318
rect 9693 2310 9915 2315
rect 9693 2286 9706 2310
rect 9730 2291 9915 2310
rect 9939 2291 10052 2315
rect 9730 2286 10052 2291
rect 9693 2282 10052 2286
rect 10119 2310 10268 2318
rect 10119 2290 10130 2310
rect 10150 2290 10268 2310
rect 10119 2283 10268 2290
rect 10119 2282 10160 2283
rect 9443 2229 9480 2230
rect 9539 2229 9576 2230
rect 9595 2229 9631 2281
rect 9650 2229 9687 2230
rect 9343 2220 9481 2229
rect 8279 2202 8310 2205
rect 8279 2176 8286 2202
rect 8305 2176 8310 2202
rect 8279 1782 8310 2176
rect 8331 2201 8499 2202
rect 8331 2198 8775 2201
rect 8331 2179 8706 2198
rect 8726 2179 8775 2198
rect 9343 2200 9452 2220
rect 9472 2200 9481 2220
rect 8331 2175 8775 2179
rect 8331 2173 8499 2175
rect 8331 1995 8358 2173
rect 8398 2135 8462 2147
rect 8738 2143 8775 2175
rect 8946 2174 9195 2196
rect 9343 2193 9481 2200
rect 9539 2220 9687 2229
rect 9539 2200 9548 2220
rect 9568 2200 9658 2220
rect 9678 2200 9687 2220
rect 9343 2191 9439 2193
rect 9539 2190 9687 2200
rect 9746 2220 9783 2230
rect 9858 2229 9895 2230
rect 9839 2227 9895 2229
rect 9746 2200 9754 2220
rect 9774 2200 9783 2220
rect 9595 2189 9631 2190
rect 8946 2143 8983 2174
rect 9159 2172 9195 2174
rect 9159 2143 9196 2172
rect 8398 2134 8433 2135
rect 8375 2129 8433 2134
rect 8375 2109 8378 2129
rect 8398 2115 8433 2129
rect 8453 2115 8462 2135
rect 8398 2107 8462 2115
rect 8424 2106 8462 2107
rect 8425 2105 8462 2106
rect 8528 2139 8564 2140
rect 8636 2139 8672 2140
rect 8528 2131 8672 2139
rect 8528 2111 8536 2131
rect 8556 2130 8644 2131
rect 8556 2111 8589 2130
rect 8528 2110 8589 2111
rect 8613 2111 8644 2130
rect 8664 2111 8672 2131
rect 8613 2110 8672 2111
rect 8528 2105 8672 2110
rect 8738 2135 8776 2143
rect 8844 2139 8880 2140
rect 8738 2115 8747 2135
rect 8767 2115 8776 2135
rect 8738 2106 8776 2115
rect 8795 2132 8880 2139
rect 8795 2112 8802 2132
rect 8823 2131 8880 2132
rect 8823 2112 8852 2131
rect 8795 2111 8852 2112
rect 8872 2111 8880 2131
rect 8738 2105 8775 2106
rect 8795 2105 8880 2111
rect 8946 2135 8984 2143
rect 9057 2139 9093 2140
rect 8946 2115 8955 2135
rect 8975 2115 8984 2135
rect 8946 2106 8984 2115
rect 9008 2131 9093 2139
rect 9008 2111 9065 2131
rect 9085 2111 9093 2131
rect 8946 2105 8983 2106
rect 9008 2105 9093 2111
rect 9159 2135 9197 2143
rect 9159 2115 9168 2135
rect 9188 2115 9197 2135
rect 9443 2130 9480 2131
rect 9746 2130 9783 2200
rect 9808 2220 9895 2227
rect 9808 2217 9866 2220
rect 9808 2197 9813 2217
rect 9834 2200 9866 2217
rect 9886 2200 9895 2220
rect 9834 2197 9895 2200
rect 9808 2190 9895 2197
rect 9954 2220 9991 2230
rect 9954 2200 9962 2220
rect 9982 2200 9991 2220
rect 9808 2189 9839 2190
rect 9442 2129 9783 2130
rect 9159 2106 9197 2115
rect 9367 2124 9783 2129
rect 9159 2105 9196 2106
rect 8582 2084 8618 2105
rect 9008 2084 9039 2105
rect 9367 2104 9370 2124
rect 9390 2104 9783 2124
rect 9954 2129 9991 2200
rect 10021 2229 10052 2282
rect 10354 2267 10391 2277
rect 10354 2249 10363 2267
rect 10381 2249 10391 2267
rect 10354 2240 10391 2249
rect 10803 2243 10838 2321
rect 11415 2311 11452 2334
rect 12208 2352 12246 2361
rect 12208 2332 12217 2352
rect 12237 2332 12246 2352
rect 12208 2324 12246 2332
rect 12312 2356 12397 2362
rect 12422 2361 12459 2362
rect 12312 2336 12320 2356
rect 12340 2336 12397 2356
rect 12312 2328 12397 2336
rect 12421 2352 12459 2361
rect 12421 2332 12430 2352
rect 12450 2332 12459 2352
rect 12312 2327 12348 2328
rect 12421 2324 12459 2332
rect 12525 2356 12610 2362
rect 12630 2361 12667 2362
rect 12525 2336 12533 2356
rect 12553 2355 12610 2356
rect 12553 2336 12582 2355
rect 12525 2335 12582 2336
rect 12603 2335 12610 2355
rect 12525 2328 12610 2335
rect 12629 2352 12667 2361
rect 12629 2332 12638 2352
rect 12658 2332 12667 2352
rect 12525 2327 12561 2328
rect 12629 2324 12667 2332
rect 12733 2356 12877 2362
rect 12733 2336 12741 2356
rect 12761 2337 12797 2356
rect 12820 2337 12849 2356
rect 12761 2336 12849 2337
rect 12869 2336 12877 2356
rect 12733 2328 12877 2336
rect 12733 2327 12769 2328
rect 12841 2327 12877 2328
rect 12943 2361 12980 2362
rect 12943 2360 12981 2361
rect 12943 2352 13007 2360
rect 12943 2332 12952 2352
rect 12972 2338 13007 2352
rect 13027 2338 13030 2358
rect 12972 2333 13030 2338
rect 12972 2332 13007 2333
rect 10071 2229 10108 2230
rect 10021 2220 10108 2229
rect 10021 2200 10079 2220
rect 10099 2200 10108 2220
rect 10021 2190 10108 2200
rect 10167 2220 10204 2230
rect 10167 2200 10175 2220
rect 10195 2200 10204 2220
rect 10021 2189 10052 2190
rect 10167 2129 10204 2200
rect 10359 2175 10390 2240
rect 10799 2234 10838 2243
rect 10799 2216 10809 2234
rect 10827 2216 10838 2234
rect 10799 2210 10838 2216
rect 10994 2286 11244 2310
rect 10994 2215 11031 2286
rect 11146 2225 11177 2226
rect 10799 2206 10836 2210
rect 10994 2195 11003 2215
rect 11023 2195 11031 2215
rect 10994 2185 11031 2195
rect 11090 2215 11177 2225
rect 11090 2195 11099 2215
rect 11119 2195 11177 2215
rect 11090 2186 11177 2195
rect 11090 2185 11127 2186
rect 10358 2165 10395 2175
rect 10358 2163 10368 2165
rect 10292 2161 10368 2163
rect 9954 2105 10204 2129
rect 10289 2147 10368 2161
rect 10386 2147 10395 2165
rect 10289 2144 10395 2147
rect 9761 2085 9782 2104
rect 10289 2085 10315 2144
rect 10358 2138 10395 2144
rect 10802 2135 10839 2144
rect 8415 2080 8515 2084
rect 8415 2076 8477 2080
rect 8415 2050 8422 2076
rect 8448 2054 8477 2076
rect 8503 2054 8515 2080
rect 8448 2050 8515 2054
rect 8415 2047 8515 2050
rect 8583 2047 8618 2084
rect 8680 2081 9039 2084
rect 8680 2076 8902 2081
rect 8680 2052 8693 2076
rect 8717 2057 8902 2076
rect 8926 2057 9039 2081
rect 8717 2052 9039 2057
rect 8680 2048 9039 2052
rect 9106 2076 9255 2084
rect 9106 2056 9117 2076
rect 9137 2056 9255 2076
rect 9761 2067 10315 2085
rect 10800 2117 10811 2135
rect 10829 2117 10839 2135
rect 11146 2133 11177 2186
rect 11207 2215 11244 2286
rect 11415 2291 11808 2311
rect 11828 2291 11831 2311
rect 12209 2295 12246 2324
rect 11415 2286 11831 2291
rect 12210 2293 12246 2295
rect 12422 2293 12459 2324
rect 11415 2285 11756 2286
rect 11359 2225 11390 2226
rect 11207 2195 11216 2215
rect 11236 2195 11244 2215
rect 11207 2185 11244 2195
rect 11303 2218 11390 2225
rect 11303 2215 11364 2218
rect 11303 2195 11312 2215
rect 11332 2198 11364 2215
rect 11385 2198 11390 2218
rect 11332 2195 11390 2198
rect 11303 2188 11390 2195
rect 11415 2215 11452 2285
rect 11718 2284 11755 2285
rect 12210 2271 12459 2293
rect 12630 2292 12667 2324
rect 12943 2320 13007 2332
rect 13047 2294 13074 2472
rect 13102 2359 13140 4190
rect 13647 4165 13654 4191
rect 13673 4165 13678 4191
rect 13554 3772 13583 3774
rect 13554 3767 13586 3772
rect 13554 3749 13561 3767
rect 13581 3749 13586 3767
rect 13647 3771 13678 4165
rect 13699 4190 13867 4191
rect 13699 4187 14143 4190
rect 13699 4168 14074 4187
rect 14094 4168 14143 4187
rect 14711 4189 14820 4209
rect 14840 4189 14849 4209
rect 13699 4164 14143 4168
rect 13699 4162 13867 4164
rect 13699 3984 13726 4162
rect 13766 4124 13830 4136
rect 14106 4132 14143 4164
rect 14314 4163 14563 4185
rect 14711 4182 14849 4189
rect 14907 4209 15055 4218
rect 14907 4189 14916 4209
rect 14936 4189 15026 4209
rect 15046 4189 15055 4209
rect 14711 4180 14807 4182
rect 14907 4179 15055 4189
rect 15114 4209 15151 4219
rect 15226 4218 15263 4219
rect 15207 4216 15263 4218
rect 15114 4189 15122 4209
rect 15142 4189 15151 4209
rect 14963 4178 14999 4179
rect 14314 4132 14351 4163
rect 14527 4161 14563 4163
rect 14527 4132 14564 4161
rect 13766 4123 13801 4124
rect 13743 4118 13801 4123
rect 13743 4098 13746 4118
rect 13766 4104 13801 4118
rect 13821 4104 13830 4124
rect 13766 4096 13830 4104
rect 13792 4095 13830 4096
rect 13793 4094 13830 4095
rect 13896 4128 13932 4129
rect 14004 4128 14040 4129
rect 13896 4120 14040 4128
rect 13896 4100 13904 4120
rect 13924 4119 14012 4120
rect 13924 4100 13957 4119
rect 13896 4099 13957 4100
rect 13981 4100 14012 4119
rect 14032 4100 14040 4120
rect 13981 4099 14040 4100
rect 13896 4094 14040 4099
rect 14106 4124 14144 4132
rect 14212 4128 14248 4129
rect 14106 4104 14115 4124
rect 14135 4104 14144 4124
rect 14106 4095 14144 4104
rect 14163 4121 14248 4128
rect 14163 4101 14170 4121
rect 14191 4120 14248 4121
rect 14191 4101 14220 4120
rect 14163 4100 14220 4101
rect 14240 4100 14248 4120
rect 14106 4094 14143 4095
rect 14163 4094 14248 4100
rect 14314 4124 14352 4132
rect 14425 4128 14461 4129
rect 14314 4104 14323 4124
rect 14343 4104 14352 4124
rect 14314 4095 14352 4104
rect 14376 4120 14461 4128
rect 14376 4100 14433 4120
rect 14453 4100 14461 4120
rect 14314 4094 14351 4095
rect 14376 4094 14461 4100
rect 14527 4124 14565 4132
rect 14527 4104 14536 4124
rect 14556 4104 14565 4124
rect 14811 4119 14848 4120
rect 15114 4119 15151 4189
rect 15176 4209 15263 4216
rect 15176 4206 15234 4209
rect 15176 4186 15181 4206
rect 15202 4189 15234 4206
rect 15254 4189 15263 4209
rect 15202 4186 15263 4189
rect 15176 4179 15263 4186
rect 15322 4209 15359 4219
rect 15322 4189 15330 4209
rect 15350 4189 15359 4209
rect 15176 4178 15207 4179
rect 14810 4118 15151 4119
rect 14527 4095 14565 4104
rect 14735 4113 15151 4118
rect 14527 4094 14564 4095
rect 13950 4073 13986 4094
rect 14376 4073 14407 4094
rect 14735 4093 14738 4113
rect 14758 4093 15151 4113
rect 15322 4118 15359 4189
rect 15389 4218 15420 4271
rect 16072 4270 16082 4288
rect 16100 4274 16721 4288
rect 17506 4287 17655 4295
rect 17722 4319 18081 4323
rect 17722 4314 18044 4319
rect 17722 4290 17835 4314
rect 17859 4295 18044 4314
rect 18068 4295 18081 4319
rect 17859 4290 18081 4295
rect 17722 4287 18081 4290
rect 18143 4287 18178 4324
rect 18246 4321 18346 4324
rect 18246 4317 18313 4321
rect 18246 4291 18258 4317
rect 18284 4295 18313 4317
rect 18339 4295 18346 4321
rect 18284 4291 18346 4295
rect 18246 4287 18346 4291
rect 16100 4270 16110 4274
rect 16551 4273 16721 4274
rect 15722 4256 15759 4266
rect 15722 4238 15731 4256
rect 15749 4238 15759 4256
rect 15722 4229 15759 4238
rect 16072 4260 16110 4270
rect 15439 4218 15476 4219
rect 15389 4209 15476 4218
rect 15389 4189 15447 4209
rect 15467 4189 15476 4209
rect 15389 4179 15476 4189
rect 15535 4209 15572 4219
rect 15535 4189 15543 4209
rect 15563 4189 15572 4209
rect 15389 4178 15420 4179
rect 15535 4118 15572 4189
rect 15727 4164 15758 4229
rect 16072 4182 16107 4260
rect 16684 4250 16721 4273
rect 17722 4266 17753 4287
rect 18143 4266 18179 4287
rect 17565 4265 17602 4266
rect 17564 4256 17602 4265
rect 16068 4173 16107 4182
rect 15726 4154 15763 4164
rect 15726 4152 15736 4154
rect 15660 4150 15736 4152
rect 15322 4094 15572 4118
rect 15657 4136 15736 4150
rect 15754 4136 15763 4154
rect 16068 4155 16078 4173
rect 16096 4155 16107 4173
rect 16068 4149 16107 4155
rect 16263 4225 16513 4249
rect 16263 4154 16300 4225
rect 16415 4164 16446 4165
rect 16068 4145 16105 4149
rect 15657 4133 15763 4136
rect 15129 4074 15150 4093
rect 15657 4074 15683 4133
rect 15726 4127 15763 4133
rect 16263 4134 16272 4154
rect 16292 4134 16300 4154
rect 16263 4124 16300 4134
rect 16359 4154 16446 4164
rect 16359 4134 16368 4154
rect 16388 4134 16446 4154
rect 16359 4125 16446 4134
rect 16359 4124 16396 4125
rect 16071 4074 16108 4083
rect 13783 4069 13883 4073
rect 13783 4065 13845 4069
rect 13783 4039 13790 4065
rect 13816 4043 13845 4065
rect 13871 4043 13883 4069
rect 13816 4039 13883 4043
rect 13783 4036 13883 4039
rect 13951 4036 13986 4073
rect 14048 4070 14407 4073
rect 14048 4065 14270 4070
rect 14048 4041 14061 4065
rect 14085 4046 14270 4065
rect 14294 4046 14407 4070
rect 14085 4041 14407 4046
rect 14048 4037 14407 4041
rect 14474 4065 14623 4073
rect 14474 4045 14485 4065
rect 14505 4045 14623 4065
rect 15129 4056 15683 4074
rect 15729 4063 15766 4065
rect 15657 4055 15683 4056
rect 15726 4055 15766 4063
rect 14474 4038 14623 4045
rect 15726 4043 15738 4055
rect 15717 4038 15738 4043
rect 14474 4037 14515 4038
rect 15133 4037 15738 4038
rect 15756 4037 15766 4055
rect 13798 3984 13835 3985
rect 13894 3984 13931 3985
rect 13950 3984 13986 4036
rect 14005 3984 14042 3985
rect 13698 3975 13836 3984
rect 13698 3955 13807 3975
rect 13827 3955 13836 3975
rect 13698 3948 13836 3955
rect 13894 3975 14042 3984
rect 13894 3955 13903 3975
rect 13923 3955 14013 3975
rect 14033 3955 14042 3975
rect 13698 3946 13794 3948
rect 13894 3945 14042 3955
rect 14101 3975 14138 3985
rect 14213 3984 14250 3985
rect 14194 3982 14250 3984
rect 14101 3955 14109 3975
rect 14129 3955 14138 3975
rect 13950 3944 13986 3945
rect 13798 3885 13835 3886
rect 14101 3885 14138 3955
rect 14163 3975 14250 3982
rect 14163 3972 14221 3975
rect 14163 3952 14168 3972
rect 14189 3955 14221 3972
rect 14241 3955 14250 3975
rect 14189 3952 14250 3955
rect 14163 3945 14250 3952
rect 14309 3975 14346 3985
rect 14309 3955 14317 3975
rect 14337 3955 14346 3975
rect 14163 3944 14194 3945
rect 13797 3884 14138 3885
rect 13722 3879 14138 3884
rect 13722 3859 13725 3879
rect 13745 3859 14138 3879
rect 14309 3884 14346 3955
rect 14376 3984 14407 4037
rect 15133 4028 15766 4037
rect 16069 4056 16080 4074
rect 16098 4056 16108 4074
rect 16415 4072 16446 4125
rect 16476 4154 16513 4225
rect 16684 4230 17077 4250
rect 17097 4230 17100 4250
rect 16684 4225 17100 4230
rect 17564 4236 17573 4256
rect 17593 4236 17602 4256
rect 17564 4228 17602 4236
rect 17668 4260 17753 4266
rect 17778 4265 17815 4266
rect 17668 4240 17676 4260
rect 17696 4240 17753 4260
rect 17668 4232 17753 4240
rect 17777 4256 17815 4265
rect 17777 4236 17786 4256
rect 17806 4236 17815 4256
rect 17668 4231 17704 4232
rect 17777 4228 17815 4236
rect 17881 4260 17966 4266
rect 17986 4265 18023 4266
rect 17881 4240 17889 4260
rect 17909 4259 17966 4260
rect 17909 4240 17938 4259
rect 17881 4239 17938 4240
rect 17959 4239 17966 4259
rect 17881 4232 17966 4239
rect 17985 4256 18023 4265
rect 17985 4236 17994 4256
rect 18014 4236 18023 4256
rect 17881 4231 17917 4232
rect 17985 4228 18023 4236
rect 18089 4261 18233 4266
rect 18089 4260 18153 4261
rect 18089 4240 18097 4260
rect 18117 4242 18153 4260
rect 18179 4260 18233 4261
rect 18179 4242 18205 4260
rect 18117 4240 18205 4242
rect 18225 4240 18233 4260
rect 18089 4232 18233 4240
rect 18089 4231 18125 4232
rect 18197 4231 18233 4232
rect 18299 4265 18336 4266
rect 18299 4264 18337 4265
rect 18299 4256 18363 4264
rect 18299 4236 18308 4256
rect 18328 4242 18363 4256
rect 18383 4242 18386 4262
rect 18328 4237 18386 4242
rect 18328 4236 18363 4237
rect 16684 4224 17025 4225
rect 16628 4164 16659 4165
rect 16476 4134 16485 4154
rect 16505 4134 16513 4154
rect 16476 4124 16513 4134
rect 16572 4157 16659 4164
rect 16572 4154 16633 4157
rect 16572 4134 16581 4154
rect 16601 4137 16633 4154
rect 16654 4137 16659 4157
rect 16601 4134 16659 4137
rect 16572 4127 16659 4134
rect 16684 4154 16721 4224
rect 16987 4223 17024 4224
rect 17565 4199 17602 4228
rect 17566 4197 17602 4199
rect 17778 4197 17815 4228
rect 17566 4175 17815 4197
rect 17986 4196 18023 4228
rect 18299 4224 18363 4236
rect 18403 4201 18430 4376
rect 18383 4198 18430 4201
rect 18262 4196 18430 4198
rect 19993 4375 20161 4377
rect 19993 4197 20020 4375
rect 20060 4337 20124 4349
rect 20400 4345 20437 4377
rect 20608 4376 20857 4398
rect 20608 4345 20645 4376
rect 20821 4374 20857 4376
rect 21000 4379 21038 4420
rect 20821 4345 20858 4374
rect 20060 4336 20095 4337
rect 20037 4331 20095 4336
rect 20037 4311 20040 4331
rect 20060 4317 20095 4331
rect 20115 4317 20124 4337
rect 20060 4309 20124 4317
rect 20086 4308 20124 4309
rect 20087 4307 20124 4308
rect 20190 4341 20226 4342
rect 20298 4341 20334 4342
rect 20190 4335 20334 4341
rect 20190 4333 20256 4335
rect 20190 4313 20198 4333
rect 20218 4314 20256 4333
rect 20278 4333 20334 4335
rect 20278 4314 20306 4333
rect 20218 4313 20306 4314
rect 20326 4313 20334 4333
rect 20190 4307 20334 4313
rect 20400 4337 20438 4345
rect 20506 4341 20542 4342
rect 20400 4317 20409 4337
rect 20429 4317 20438 4337
rect 20400 4308 20438 4317
rect 20457 4334 20542 4341
rect 20457 4314 20464 4334
rect 20485 4333 20542 4334
rect 20485 4314 20514 4333
rect 20457 4313 20514 4314
rect 20534 4313 20542 4333
rect 20400 4307 20437 4308
rect 20457 4307 20542 4313
rect 20608 4337 20646 4345
rect 20719 4341 20755 4342
rect 20608 4317 20617 4337
rect 20637 4317 20646 4337
rect 20608 4308 20646 4317
rect 20670 4333 20755 4341
rect 20670 4313 20727 4333
rect 20747 4313 20755 4333
rect 20608 4307 20645 4308
rect 20670 4307 20755 4313
rect 20821 4337 20859 4345
rect 20821 4317 20830 4337
rect 20850 4317 20859 4337
rect 20821 4308 20859 4317
rect 21000 4344 21036 4379
rect 21000 4334 21037 4344
rect 21000 4316 21010 4334
rect 21028 4316 21037 4334
rect 20821 4307 20858 4308
rect 21000 4307 21037 4316
rect 20244 4286 20280 4307
rect 20670 4286 20701 4307
rect 20077 4282 20177 4286
rect 20077 4278 20139 4282
rect 20077 4252 20084 4278
rect 20110 4256 20139 4278
rect 20165 4256 20177 4282
rect 20110 4252 20177 4256
rect 20077 4249 20177 4252
rect 20245 4249 20280 4286
rect 20342 4283 20701 4286
rect 20342 4278 20564 4283
rect 20342 4254 20355 4278
rect 20379 4259 20564 4278
rect 20588 4259 20701 4283
rect 20379 4254 20701 4259
rect 20342 4250 20701 4254
rect 20768 4278 20917 4286
rect 20768 4258 20779 4278
rect 20799 4258 20917 4278
rect 20768 4251 20917 4258
rect 20768 4250 20809 4251
rect 20092 4197 20129 4198
rect 20188 4197 20225 4198
rect 20244 4197 20280 4249
rect 20299 4197 20336 4198
rect 17986 4170 18430 4196
rect 19992 4188 20130 4197
rect 18262 4169 18430 4170
rect 18928 4170 18959 4173
rect 16836 4164 16872 4165
rect 16684 4134 16693 4154
rect 16713 4134 16721 4154
rect 16572 4125 16628 4127
rect 16572 4124 16609 4125
rect 16684 4124 16721 4134
rect 16780 4154 16928 4164
rect 17028 4161 17124 4163
rect 16780 4134 16789 4154
rect 16809 4134 16899 4154
rect 16919 4134 16928 4154
rect 16780 4125 16928 4134
rect 16986 4154 17124 4161
rect 16986 4134 16995 4154
rect 17015 4134 17124 4154
rect 16986 4125 17124 4134
rect 16780 4124 16817 4125
rect 16836 4073 16872 4125
rect 16891 4124 16928 4125
rect 16987 4124 17024 4125
rect 16307 4071 16348 4072
rect 15133 4021 15765 4028
rect 15133 4019 15195 4021
rect 14711 4009 14879 4010
rect 15133 4009 15155 4019
rect 14426 3984 14463 3985
rect 14376 3975 14463 3984
rect 14376 3955 14434 3975
rect 14454 3955 14463 3975
rect 14376 3945 14463 3955
rect 14522 3975 14559 3985
rect 14522 3955 14530 3975
rect 14550 3955 14559 3975
rect 14376 3944 14407 3945
rect 14522 3884 14559 3955
rect 14309 3860 14559 3884
rect 14711 3983 15155 4009
rect 14711 3981 14879 3983
rect 14711 3803 14738 3981
rect 14778 3943 14842 3955
rect 15118 3951 15155 3983
rect 15326 3982 15575 4004
rect 15326 3951 15363 3982
rect 15539 3980 15575 3982
rect 15539 3951 15576 3980
rect 14778 3942 14813 3943
rect 14755 3937 14813 3942
rect 14755 3917 14758 3937
rect 14778 3923 14813 3937
rect 14833 3923 14842 3943
rect 14778 3915 14842 3923
rect 14804 3914 14842 3915
rect 14805 3913 14842 3914
rect 14908 3947 14944 3948
rect 15016 3947 15052 3948
rect 14908 3939 15052 3947
rect 14908 3919 14916 3939
rect 14936 3919 14965 3939
rect 14908 3918 14965 3919
rect 14987 3919 15024 3939
rect 15044 3919 15052 3939
rect 14987 3918 15052 3919
rect 14908 3913 15052 3918
rect 15118 3943 15156 3951
rect 15224 3947 15260 3948
rect 15118 3923 15127 3943
rect 15147 3923 15156 3943
rect 15118 3914 15156 3923
rect 15175 3940 15260 3947
rect 15175 3920 15182 3940
rect 15203 3939 15260 3940
rect 15203 3920 15232 3939
rect 15175 3919 15232 3920
rect 15252 3919 15260 3939
rect 15118 3913 15155 3914
rect 15175 3913 15260 3919
rect 15326 3943 15364 3951
rect 15437 3947 15473 3948
rect 15326 3923 15335 3943
rect 15355 3923 15364 3943
rect 15326 3914 15364 3923
rect 15388 3939 15473 3947
rect 15388 3919 15445 3939
rect 15465 3919 15473 3939
rect 15326 3913 15363 3914
rect 15388 3913 15473 3919
rect 15539 3943 15577 3951
rect 15539 3923 15548 3943
rect 15568 3923 15577 3943
rect 15539 3914 15577 3923
rect 15539 3913 15576 3914
rect 14962 3892 14998 3913
rect 15388 3892 15419 3913
rect 14795 3888 14895 3892
rect 14795 3884 14857 3888
rect 14795 3858 14802 3884
rect 14828 3862 14857 3884
rect 14883 3862 14895 3888
rect 14828 3858 14895 3862
rect 14795 3855 14895 3858
rect 14963 3855 14998 3892
rect 15060 3889 15419 3892
rect 15060 3884 15282 3889
rect 15060 3860 15073 3884
rect 15097 3865 15282 3884
rect 15306 3865 15419 3889
rect 15097 3860 15419 3865
rect 15060 3856 15419 3860
rect 15486 3884 15635 3892
rect 15486 3864 15497 3884
rect 15517 3864 15635 3884
rect 15486 3857 15635 3864
rect 15726 3872 15765 4021
rect 16069 3907 16108 4056
rect 16199 4064 16348 4071
rect 16199 4044 16317 4064
rect 16337 4044 16348 4064
rect 16199 4036 16348 4044
rect 16415 4068 16774 4072
rect 16415 4063 16737 4068
rect 16415 4039 16528 4063
rect 16552 4044 16737 4063
rect 16761 4044 16774 4068
rect 16552 4039 16774 4044
rect 16415 4036 16774 4039
rect 16836 4036 16871 4073
rect 16939 4070 17039 4073
rect 16939 4066 17006 4070
rect 16939 4040 16951 4066
rect 16977 4044 17006 4066
rect 17032 4044 17039 4070
rect 16977 4040 17039 4044
rect 16939 4036 17039 4040
rect 16415 4015 16446 4036
rect 16836 4015 16872 4036
rect 16258 4014 16295 4015
rect 16257 4005 16295 4014
rect 16257 3985 16266 4005
rect 16286 3985 16295 4005
rect 16257 3977 16295 3985
rect 16361 4009 16446 4015
rect 16471 4014 16508 4015
rect 16361 3989 16369 4009
rect 16389 3989 16446 4009
rect 16361 3981 16446 3989
rect 16470 4005 16508 4014
rect 16470 3985 16479 4005
rect 16499 3985 16508 4005
rect 16361 3980 16397 3981
rect 16470 3977 16508 3985
rect 16574 4009 16659 4015
rect 16679 4014 16716 4015
rect 16574 3989 16582 4009
rect 16602 4008 16659 4009
rect 16602 3989 16631 4008
rect 16574 3988 16631 3989
rect 16652 3988 16659 4008
rect 16574 3981 16659 3988
rect 16678 4005 16716 4014
rect 16678 3985 16687 4005
rect 16707 3985 16716 4005
rect 16574 3980 16610 3981
rect 16678 3977 16716 3985
rect 16782 4010 16926 4015
rect 16782 4009 16847 4010
rect 16782 3989 16790 4009
rect 16810 3989 16847 4009
rect 16869 4009 16926 4010
rect 16869 3989 16898 4009
rect 16918 3989 16926 4009
rect 16782 3981 16926 3989
rect 16782 3980 16818 3981
rect 16890 3980 16926 3981
rect 16992 4014 17029 4015
rect 16992 4013 17030 4014
rect 16992 4005 17056 4013
rect 16992 3985 17001 4005
rect 17021 3991 17056 4005
rect 17076 3991 17079 4011
rect 17021 3986 17079 3991
rect 17021 3985 17056 3986
rect 16258 3948 16295 3977
rect 16259 3946 16295 3948
rect 16471 3946 16508 3977
rect 16259 3924 16508 3946
rect 16679 3945 16716 3977
rect 16992 3973 17056 3985
rect 17096 3947 17123 4125
rect 16955 3945 17123 3947
rect 16679 3919 17123 3945
rect 17275 4044 17525 4068
rect 17275 3973 17312 4044
rect 17427 3983 17458 3984
rect 17275 3953 17284 3973
rect 17304 3953 17312 3973
rect 17275 3943 17312 3953
rect 17371 3973 17458 3983
rect 17371 3953 17380 3973
rect 17400 3953 17458 3973
rect 17371 3944 17458 3953
rect 17371 3943 17408 3944
rect 16679 3909 16701 3919
rect 16955 3918 17123 3919
rect 16639 3907 16701 3909
rect 16069 3900 16701 3907
rect 15486 3856 15527 3857
rect 14810 3803 14847 3804
rect 14906 3803 14943 3804
rect 14962 3803 14998 3855
rect 15017 3803 15054 3804
rect 14710 3794 14848 3803
rect 14710 3774 14819 3794
rect 14839 3774 14848 3794
rect 13647 3770 13817 3771
rect 13647 3755 14093 3770
rect 14710 3767 14848 3774
rect 14906 3794 15054 3803
rect 14906 3774 14915 3794
rect 14935 3774 15025 3794
rect 15045 3774 15054 3794
rect 14710 3765 14806 3767
rect 13554 3744 13586 3749
rect 13556 2743 13586 3744
rect 13649 3744 14093 3755
rect 13649 3742 13817 3744
rect 13649 3564 13676 3742
rect 13716 3704 13780 3716
rect 14056 3712 14093 3744
rect 14264 3743 14513 3765
rect 14906 3764 15054 3774
rect 15113 3794 15150 3804
rect 15225 3803 15262 3804
rect 15206 3801 15262 3803
rect 15113 3774 15121 3794
rect 15141 3774 15150 3794
rect 14962 3763 14998 3764
rect 14264 3712 14301 3743
rect 14477 3741 14513 3743
rect 14477 3712 14514 3741
rect 13716 3703 13751 3704
rect 13693 3698 13751 3703
rect 13693 3678 13696 3698
rect 13716 3684 13751 3698
rect 13771 3684 13780 3704
rect 13716 3676 13780 3684
rect 13742 3675 13780 3676
rect 13743 3674 13780 3675
rect 13846 3708 13882 3709
rect 13954 3708 13990 3709
rect 13846 3700 13990 3708
rect 13846 3680 13854 3700
rect 13874 3681 13906 3700
rect 13929 3681 13962 3700
rect 13874 3680 13962 3681
rect 13982 3680 13990 3700
rect 13846 3674 13990 3680
rect 14056 3704 14094 3712
rect 14162 3708 14198 3709
rect 14056 3684 14065 3704
rect 14085 3684 14094 3704
rect 14056 3675 14094 3684
rect 14113 3701 14198 3708
rect 14113 3681 14120 3701
rect 14141 3700 14198 3701
rect 14141 3681 14170 3700
rect 14113 3680 14170 3681
rect 14190 3680 14198 3700
rect 14056 3674 14093 3675
rect 14113 3674 14198 3680
rect 14264 3704 14302 3712
rect 14375 3708 14411 3709
rect 14264 3684 14273 3704
rect 14293 3684 14302 3704
rect 14264 3675 14302 3684
rect 14326 3700 14411 3708
rect 14326 3680 14383 3700
rect 14403 3680 14411 3700
rect 14264 3674 14301 3675
rect 14326 3674 14411 3680
rect 14477 3704 14515 3712
rect 14810 3704 14847 3705
rect 15113 3704 15150 3774
rect 15175 3794 15262 3801
rect 15175 3791 15233 3794
rect 15175 3771 15180 3791
rect 15201 3774 15233 3791
rect 15253 3774 15262 3794
rect 15201 3771 15262 3774
rect 15175 3764 15262 3771
rect 15321 3794 15358 3804
rect 15321 3774 15329 3794
rect 15349 3774 15358 3794
rect 15175 3763 15206 3764
rect 14477 3684 14486 3704
rect 14506 3684 14515 3704
rect 14809 3703 15150 3704
rect 14477 3675 14515 3684
rect 14734 3698 15150 3703
rect 14734 3678 14737 3698
rect 14757 3678 15150 3698
rect 15321 3703 15358 3774
rect 15388 3803 15419 3856
rect 15726 3854 15736 3872
rect 15754 3854 15765 3872
rect 16068 3891 16701 3900
rect 17427 3891 17458 3944
rect 17488 3973 17525 4044
rect 17696 4049 18089 4069
rect 18109 4049 18112 4069
rect 17696 4044 18112 4049
rect 17696 4043 18037 4044
rect 17640 3983 17671 3984
rect 17488 3953 17497 3973
rect 17517 3953 17525 3973
rect 17488 3943 17525 3953
rect 17584 3976 17671 3983
rect 17584 3973 17645 3976
rect 17584 3953 17593 3973
rect 17613 3956 17645 3973
rect 17666 3956 17671 3976
rect 17613 3953 17671 3956
rect 17584 3946 17671 3953
rect 17696 3973 17733 4043
rect 17999 4042 18036 4043
rect 17848 3983 17884 3984
rect 17696 3953 17705 3973
rect 17725 3953 17733 3973
rect 17584 3944 17640 3946
rect 17584 3943 17621 3944
rect 17696 3943 17733 3953
rect 17792 3973 17940 3983
rect 18040 3980 18136 3982
rect 17792 3953 17801 3973
rect 17821 3953 17911 3973
rect 17931 3953 17940 3973
rect 17792 3944 17940 3953
rect 17998 3973 18136 3980
rect 17998 3953 18007 3973
rect 18027 3953 18136 3973
rect 17998 3944 18136 3953
rect 17792 3943 17829 3944
rect 17848 3892 17884 3944
rect 17903 3943 17940 3944
rect 17999 3943 18036 3944
rect 16068 3873 16078 3891
rect 16096 3890 16701 3891
rect 17319 3890 17360 3891
rect 16096 3885 16117 3890
rect 16096 3873 16108 3885
rect 17211 3883 17360 3890
rect 16068 3865 16108 3873
rect 16151 3872 16177 3873
rect 16068 3863 16105 3865
rect 16151 3854 16705 3872
rect 17211 3863 17329 3883
rect 17349 3863 17360 3883
rect 17211 3855 17360 3863
rect 17427 3887 17786 3891
rect 17427 3882 17749 3887
rect 17427 3858 17540 3882
rect 17564 3863 17749 3882
rect 17773 3863 17786 3887
rect 17564 3858 17786 3863
rect 17427 3855 17786 3858
rect 17848 3855 17883 3892
rect 17951 3889 18051 3892
rect 17951 3885 18018 3889
rect 17951 3859 17963 3885
rect 17989 3863 18018 3885
rect 18044 3863 18051 3889
rect 17989 3859 18051 3863
rect 17951 3855 18051 3859
rect 15726 3845 15763 3854
rect 15438 3803 15475 3804
rect 15388 3794 15475 3803
rect 15388 3774 15446 3794
rect 15466 3774 15475 3794
rect 15388 3764 15475 3774
rect 15534 3794 15571 3804
rect 15534 3774 15542 3794
rect 15562 3774 15571 3794
rect 16071 3795 16108 3801
rect 16151 3795 16177 3854
rect 16684 3835 16705 3854
rect 16071 3792 16177 3795
rect 15729 3779 15766 3783
rect 15388 3763 15419 3764
rect 15534 3703 15571 3774
rect 15321 3679 15571 3703
rect 15727 3773 15766 3779
rect 15727 3755 15738 3773
rect 15756 3755 15766 3773
rect 16071 3774 16080 3792
rect 16098 3778 16177 3792
rect 16262 3810 16512 3834
rect 16098 3776 16174 3778
rect 16098 3774 16108 3776
rect 16071 3764 16108 3774
rect 15727 3746 15766 3755
rect 14477 3674 14514 3675
rect 13900 3653 13936 3674
rect 14326 3653 14357 3674
rect 15113 3655 15150 3678
rect 15727 3668 15762 3746
rect 16076 3699 16107 3764
rect 16262 3739 16299 3810
rect 16414 3749 16445 3750
rect 16262 3719 16271 3739
rect 16291 3719 16299 3739
rect 16262 3709 16299 3719
rect 16358 3739 16445 3749
rect 16358 3719 16367 3739
rect 16387 3719 16445 3739
rect 16358 3710 16445 3719
rect 16358 3709 16395 3710
rect 15724 3658 15762 3668
rect 16075 3690 16112 3699
rect 16075 3672 16085 3690
rect 16103 3672 16112 3690
rect 16075 3662 16112 3672
rect 15113 3654 15283 3655
rect 15724 3654 15734 3658
rect 13733 3649 13833 3653
rect 13733 3645 13795 3649
rect 13733 3619 13740 3645
rect 13766 3623 13795 3645
rect 13821 3623 13833 3649
rect 13766 3619 13833 3623
rect 13733 3616 13833 3619
rect 13901 3616 13936 3653
rect 13998 3650 14357 3653
rect 13998 3645 14220 3650
rect 13998 3621 14011 3645
rect 14035 3626 14220 3645
rect 14244 3626 14357 3650
rect 14035 3621 14357 3626
rect 13998 3617 14357 3621
rect 14424 3645 14573 3653
rect 14424 3625 14435 3645
rect 14455 3625 14573 3645
rect 15113 3640 15734 3654
rect 15752 3640 15762 3658
rect 16414 3657 16445 3710
rect 16475 3739 16512 3810
rect 16683 3815 17076 3835
rect 17096 3815 17099 3835
rect 17427 3834 17458 3855
rect 17848 3834 17884 3855
rect 17270 3833 17307 3834
rect 16683 3810 17099 3815
rect 17269 3824 17307 3833
rect 16683 3809 17024 3810
rect 16627 3749 16658 3750
rect 16475 3719 16484 3739
rect 16504 3719 16512 3739
rect 16475 3709 16512 3719
rect 16571 3742 16658 3749
rect 16571 3739 16632 3742
rect 16571 3719 16580 3739
rect 16600 3722 16632 3739
rect 16653 3722 16658 3742
rect 16600 3719 16658 3722
rect 16571 3712 16658 3719
rect 16683 3739 16720 3809
rect 16986 3808 17023 3809
rect 17269 3804 17278 3824
rect 17298 3804 17307 3824
rect 17269 3796 17307 3804
rect 17373 3828 17458 3834
rect 17483 3833 17520 3834
rect 17373 3808 17381 3828
rect 17401 3808 17458 3828
rect 17373 3800 17458 3808
rect 17482 3824 17520 3833
rect 17482 3804 17491 3824
rect 17511 3804 17520 3824
rect 17373 3799 17409 3800
rect 17482 3796 17520 3804
rect 17586 3828 17671 3834
rect 17691 3833 17728 3834
rect 17586 3808 17594 3828
rect 17614 3827 17671 3828
rect 17614 3808 17643 3827
rect 17586 3807 17643 3808
rect 17664 3807 17671 3827
rect 17586 3800 17671 3807
rect 17690 3824 17728 3833
rect 17690 3804 17699 3824
rect 17719 3804 17728 3824
rect 17586 3799 17622 3800
rect 17690 3796 17728 3804
rect 17794 3828 17938 3834
rect 17794 3808 17802 3828
rect 17822 3808 17854 3828
rect 17878 3808 17910 3828
rect 17930 3808 17938 3828
rect 17794 3800 17938 3808
rect 17794 3799 17830 3800
rect 17902 3799 17938 3800
rect 18004 3833 18041 3834
rect 18004 3832 18042 3833
rect 18004 3824 18068 3832
rect 18004 3804 18013 3824
rect 18033 3810 18068 3824
rect 18088 3810 18091 3830
rect 18033 3805 18091 3810
rect 18033 3804 18068 3805
rect 17270 3767 17307 3796
rect 17271 3765 17307 3767
rect 17483 3765 17520 3796
rect 16835 3749 16871 3750
rect 16683 3719 16692 3739
rect 16712 3719 16720 3739
rect 16571 3710 16627 3712
rect 16571 3709 16608 3710
rect 16683 3709 16720 3719
rect 16779 3739 16927 3749
rect 17027 3746 17123 3748
rect 16779 3719 16788 3739
rect 16808 3719 16898 3739
rect 16918 3719 16927 3739
rect 16779 3710 16927 3719
rect 16985 3739 17123 3746
rect 17271 3743 17520 3765
rect 17691 3764 17728 3796
rect 18004 3792 18068 3804
rect 18108 3766 18135 3944
rect 17967 3764 18135 3766
rect 17691 3760 18135 3764
rect 16985 3719 16994 3739
rect 17014 3719 17123 3739
rect 17691 3741 17740 3760
rect 17760 3741 18135 3760
rect 17691 3738 18135 3741
rect 17967 3737 18135 3738
rect 16985 3710 17123 3719
rect 16779 3709 16816 3710
rect 16835 3658 16871 3710
rect 16890 3709 16927 3710
rect 16986 3709 17023 3710
rect 16306 3656 16347 3657
rect 15113 3634 15762 3640
rect 16198 3649 16347 3656
rect 15113 3633 15761 3634
rect 15724 3631 15761 3633
rect 14424 3618 14573 3625
rect 16198 3629 16316 3649
rect 16336 3629 16347 3649
rect 16198 3621 16347 3629
rect 16414 3653 16773 3657
rect 16414 3648 16736 3653
rect 16414 3624 16527 3648
rect 16551 3629 16736 3648
rect 16760 3629 16773 3653
rect 16551 3624 16773 3629
rect 16414 3621 16773 3624
rect 16835 3621 16870 3658
rect 16938 3655 17038 3658
rect 16938 3651 17005 3655
rect 16938 3625 16950 3651
rect 16976 3629 17005 3651
rect 17031 3629 17038 3655
rect 16976 3625 17038 3629
rect 16938 3621 17038 3625
rect 14424 3617 14465 3618
rect 13748 3564 13785 3565
rect 13844 3564 13881 3565
rect 13900 3564 13936 3616
rect 13955 3564 13992 3565
rect 13648 3555 13786 3564
rect 13648 3535 13757 3555
rect 13777 3535 13786 3555
rect 13648 3528 13786 3535
rect 13844 3555 13992 3564
rect 13844 3535 13853 3555
rect 13873 3535 13963 3555
rect 13983 3535 13992 3555
rect 13648 3526 13744 3528
rect 13844 3525 13992 3535
rect 14051 3555 14088 3565
rect 14163 3564 14200 3565
rect 14144 3562 14200 3564
rect 14051 3535 14059 3555
rect 14079 3535 14088 3555
rect 13900 3524 13936 3525
rect 13748 3465 13785 3466
rect 14051 3465 14088 3535
rect 14113 3555 14200 3562
rect 14113 3552 14171 3555
rect 14113 3532 14118 3552
rect 14139 3535 14171 3552
rect 14191 3535 14200 3555
rect 14139 3532 14200 3535
rect 14113 3525 14200 3532
rect 14259 3555 14296 3565
rect 14259 3535 14267 3555
rect 14287 3535 14296 3555
rect 14113 3524 14144 3525
rect 13747 3464 14088 3465
rect 13672 3459 14088 3464
rect 13672 3439 13675 3459
rect 13695 3439 14088 3459
rect 14259 3464 14296 3535
rect 14326 3564 14357 3617
rect 16414 3600 16445 3621
rect 16835 3600 16871 3621
rect 16078 3591 16115 3600
rect 16257 3599 16294 3600
rect 16078 3573 16087 3591
rect 16105 3573 16115 3591
rect 14376 3564 14413 3565
rect 14326 3555 14413 3564
rect 14326 3535 14384 3555
rect 14404 3535 14413 3555
rect 14326 3525 14413 3535
rect 14472 3555 14509 3565
rect 14472 3535 14480 3555
rect 14500 3535 14509 3555
rect 14326 3524 14357 3525
rect 14472 3464 14509 3535
rect 15727 3559 15764 3569
rect 16078 3563 16115 3573
rect 15727 3541 15736 3559
rect 15754 3541 15764 3559
rect 15727 3532 15764 3541
rect 15727 3508 15762 3532
rect 16079 3528 16115 3563
rect 16256 3590 16294 3599
rect 16256 3570 16265 3590
rect 16285 3570 16294 3590
rect 16256 3562 16294 3570
rect 16360 3594 16445 3600
rect 16470 3599 16507 3600
rect 16360 3574 16368 3594
rect 16388 3574 16445 3594
rect 16360 3566 16445 3574
rect 16469 3590 16507 3599
rect 16469 3570 16478 3590
rect 16498 3570 16507 3590
rect 16360 3565 16396 3566
rect 16469 3562 16507 3570
rect 16573 3594 16658 3600
rect 16678 3599 16715 3600
rect 16573 3574 16581 3594
rect 16601 3593 16658 3594
rect 16601 3574 16630 3593
rect 16573 3573 16630 3574
rect 16651 3573 16658 3593
rect 16573 3566 16658 3573
rect 16677 3590 16715 3599
rect 16677 3570 16686 3590
rect 16706 3570 16715 3590
rect 16573 3565 16609 3566
rect 16677 3562 16715 3570
rect 16781 3594 16925 3600
rect 16781 3574 16789 3594
rect 16809 3593 16897 3594
rect 16809 3574 16837 3593
rect 16781 3572 16837 3574
rect 16859 3574 16897 3593
rect 16917 3574 16925 3594
rect 16859 3572 16925 3574
rect 16781 3566 16925 3572
rect 16781 3565 16817 3566
rect 16889 3565 16925 3566
rect 16991 3599 17028 3600
rect 16991 3598 17029 3599
rect 16991 3590 17055 3598
rect 16991 3570 17000 3590
rect 17020 3576 17055 3590
rect 17075 3576 17078 3596
rect 17020 3571 17078 3576
rect 17020 3570 17055 3571
rect 16257 3533 16294 3562
rect 15725 3484 15762 3508
rect 15724 3478 15762 3484
rect 14259 3440 14509 3464
rect 15135 3460 15762 3478
rect 14717 3443 14885 3444
rect 15136 3443 15160 3460
rect 14717 3417 15161 3443
rect 14717 3415 14885 3417
rect 14717 3237 14744 3415
rect 14784 3377 14848 3389
rect 15124 3385 15161 3417
rect 15332 3416 15581 3438
rect 15332 3385 15369 3416
rect 15545 3414 15581 3416
rect 15724 3419 15762 3460
rect 16077 3487 16115 3528
rect 16258 3531 16294 3533
rect 16470 3531 16507 3562
rect 16258 3509 16507 3531
rect 16678 3530 16715 3562
rect 16991 3558 17055 3570
rect 17095 3532 17122 3710
rect 16954 3530 17122 3532
rect 16678 3504 17122 3530
rect 16679 3487 16703 3504
rect 16954 3503 17122 3504
rect 16077 3469 16704 3487
rect 17330 3483 17580 3507
rect 16077 3463 16115 3469
rect 16077 3439 16114 3463
rect 15545 3385 15582 3414
rect 14784 3376 14819 3377
rect 14761 3371 14819 3376
rect 14761 3351 14764 3371
rect 14784 3357 14819 3371
rect 14839 3357 14848 3377
rect 14784 3349 14848 3357
rect 14810 3348 14848 3349
rect 14811 3347 14848 3348
rect 14914 3381 14950 3382
rect 15022 3381 15058 3382
rect 14914 3375 15058 3381
rect 14914 3373 14980 3375
rect 14914 3353 14922 3373
rect 14942 3354 14980 3373
rect 15002 3373 15058 3375
rect 15002 3354 15030 3373
rect 14942 3353 15030 3354
rect 15050 3353 15058 3373
rect 14914 3347 15058 3353
rect 15124 3377 15162 3385
rect 15230 3381 15266 3382
rect 15124 3357 15133 3377
rect 15153 3357 15162 3377
rect 15124 3348 15162 3357
rect 15181 3374 15266 3381
rect 15181 3354 15188 3374
rect 15209 3373 15266 3374
rect 15209 3354 15238 3373
rect 15181 3353 15238 3354
rect 15258 3353 15266 3373
rect 15124 3347 15161 3348
rect 15181 3347 15266 3353
rect 15332 3377 15370 3385
rect 15443 3381 15479 3382
rect 15332 3357 15341 3377
rect 15361 3357 15370 3377
rect 15332 3348 15370 3357
rect 15394 3373 15479 3381
rect 15394 3353 15451 3373
rect 15471 3353 15479 3373
rect 15332 3347 15369 3348
rect 15394 3347 15479 3353
rect 15545 3377 15583 3385
rect 15545 3357 15554 3377
rect 15574 3357 15583 3377
rect 15545 3348 15583 3357
rect 15724 3384 15760 3419
rect 16077 3415 16112 3439
rect 16075 3406 16112 3415
rect 16075 3388 16085 3406
rect 16103 3388 16112 3406
rect 15724 3374 15761 3384
rect 16075 3378 16112 3388
rect 17330 3412 17367 3483
rect 17482 3422 17513 3423
rect 17330 3392 17339 3412
rect 17359 3392 17367 3412
rect 17330 3382 17367 3392
rect 17426 3412 17513 3422
rect 17426 3392 17435 3412
rect 17455 3392 17513 3412
rect 17426 3383 17513 3392
rect 17426 3382 17463 3383
rect 15724 3356 15734 3374
rect 15752 3356 15761 3374
rect 15545 3347 15582 3348
rect 15724 3347 15761 3356
rect 14968 3326 15004 3347
rect 15394 3326 15425 3347
rect 17482 3330 17513 3383
rect 17543 3412 17580 3483
rect 17751 3488 18144 3508
rect 18164 3488 18167 3508
rect 17751 3483 18167 3488
rect 17751 3482 18092 3483
rect 17695 3422 17726 3423
rect 17543 3392 17552 3412
rect 17572 3392 17580 3412
rect 17543 3382 17580 3392
rect 17639 3415 17726 3422
rect 17639 3412 17700 3415
rect 17639 3392 17648 3412
rect 17668 3395 17700 3412
rect 17721 3395 17726 3415
rect 17668 3392 17726 3395
rect 17639 3385 17726 3392
rect 17751 3412 17788 3482
rect 18054 3481 18091 3482
rect 17903 3422 17939 3423
rect 17751 3392 17760 3412
rect 17780 3392 17788 3412
rect 17639 3383 17695 3385
rect 17639 3382 17676 3383
rect 17751 3382 17788 3392
rect 17847 3412 17995 3422
rect 18095 3419 18191 3421
rect 17847 3392 17856 3412
rect 17876 3392 17966 3412
rect 17986 3392 17995 3412
rect 17847 3383 17995 3392
rect 18053 3412 18191 3419
rect 18053 3392 18062 3412
rect 18082 3392 18191 3412
rect 18053 3383 18191 3392
rect 17847 3382 17884 3383
rect 17903 3331 17939 3383
rect 17958 3382 17995 3383
rect 18054 3382 18091 3383
rect 17374 3329 17415 3330
rect 14801 3322 14901 3326
rect 14801 3318 14863 3322
rect 14801 3292 14808 3318
rect 14834 3296 14863 3318
rect 14889 3296 14901 3322
rect 14834 3292 14901 3296
rect 14801 3289 14901 3292
rect 14969 3289 15004 3326
rect 15066 3323 15425 3326
rect 15066 3318 15288 3323
rect 15066 3294 15079 3318
rect 15103 3299 15288 3318
rect 15312 3299 15425 3323
rect 15103 3294 15425 3299
rect 15066 3290 15425 3294
rect 15492 3318 15641 3326
rect 15492 3298 15503 3318
rect 15523 3298 15641 3318
rect 17266 3322 17415 3329
rect 16078 3314 16115 3316
rect 16078 3313 16726 3314
rect 15492 3291 15641 3298
rect 16077 3307 16726 3313
rect 15492 3290 15533 3291
rect 14816 3237 14853 3238
rect 14912 3237 14949 3238
rect 14968 3237 15004 3289
rect 15023 3237 15060 3238
rect 14716 3228 14854 3237
rect 13704 3209 13872 3210
rect 13704 3206 14148 3209
rect 13704 3187 14079 3206
rect 14099 3187 14148 3206
rect 14716 3208 14825 3228
rect 14845 3208 14854 3228
rect 13704 3183 14148 3187
rect 13704 3181 13872 3183
rect 13704 3003 13731 3181
rect 13771 3143 13835 3155
rect 14111 3151 14148 3183
rect 14319 3182 14568 3204
rect 14716 3201 14854 3208
rect 14912 3228 15060 3237
rect 14912 3208 14921 3228
rect 14941 3208 15031 3228
rect 15051 3208 15060 3228
rect 14716 3199 14812 3201
rect 14912 3198 15060 3208
rect 15119 3228 15156 3238
rect 15231 3237 15268 3238
rect 15212 3235 15268 3237
rect 15119 3208 15127 3228
rect 15147 3208 15156 3228
rect 14968 3197 15004 3198
rect 14319 3151 14356 3182
rect 14532 3180 14568 3182
rect 14532 3151 14569 3180
rect 13771 3142 13806 3143
rect 13748 3137 13806 3142
rect 13748 3117 13751 3137
rect 13771 3123 13806 3137
rect 13826 3123 13835 3143
rect 13771 3115 13835 3123
rect 13797 3114 13835 3115
rect 13798 3113 13835 3114
rect 13901 3147 13937 3148
rect 14009 3147 14045 3148
rect 13901 3139 14045 3147
rect 13901 3119 13909 3139
rect 13929 3119 13961 3139
rect 13985 3119 14017 3139
rect 14037 3119 14045 3139
rect 13901 3113 14045 3119
rect 14111 3143 14149 3151
rect 14217 3147 14253 3148
rect 14111 3123 14120 3143
rect 14140 3123 14149 3143
rect 14111 3114 14149 3123
rect 14168 3140 14253 3147
rect 14168 3120 14175 3140
rect 14196 3139 14253 3140
rect 14196 3120 14225 3139
rect 14168 3119 14225 3120
rect 14245 3119 14253 3139
rect 14111 3113 14148 3114
rect 14168 3113 14253 3119
rect 14319 3143 14357 3151
rect 14430 3147 14466 3148
rect 14319 3123 14328 3143
rect 14348 3123 14357 3143
rect 14319 3114 14357 3123
rect 14381 3139 14466 3147
rect 14381 3119 14438 3139
rect 14458 3119 14466 3139
rect 14319 3113 14356 3114
rect 14381 3113 14466 3119
rect 14532 3143 14570 3151
rect 14532 3123 14541 3143
rect 14561 3123 14570 3143
rect 14816 3138 14853 3139
rect 15119 3138 15156 3208
rect 15181 3228 15268 3235
rect 15181 3225 15239 3228
rect 15181 3205 15186 3225
rect 15207 3208 15239 3225
rect 15259 3208 15268 3228
rect 15207 3205 15268 3208
rect 15181 3198 15268 3205
rect 15327 3228 15364 3238
rect 15327 3208 15335 3228
rect 15355 3208 15364 3228
rect 15181 3197 15212 3198
rect 14815 3137 15156 3138
rect 14532 3114 14570 3123
rect 14740 3132 15156 3137
rect 14532 3113 14569 3114
rect 13955 3092 13991 3113
rect 14381 3092 14412 3113
rect 14740 3112 14743 3132
rect 14763 3112 15156 3132
rect 15327 3137 15364 3208
rect 15394 3237 15425 3290
rect 16077 3289 16087 3307
rect 16105 3293 16726 3307
rect 17266 3302 17384 3322
rect 17404 3302 17415 3322
rect 17266 3294 17415 3302
rect 17482 3326 17841 3330
rect 17482 3321 17804 3326
rect 17482 3297 17595 3321
rect 17619 3302 17804 3321
rect 17828 3302 17841 3326
rect 17619 3297 17841 3302
rect 17482 3294 17841 3297
rect 17903 3294 17938 3331
rect 18006 3328 18106 3331
rect 18006 3324 18073 3328
rect 18006 3298 18018 3324
rect 18044 3302 18073 3324
rect 18099 3302 18106 3328
rect 18044 3298 18106 3302
rect 18006 3294 18106 3298
rect 16105 3289 16115 3293
rect 16556 3292 16726 3293
rect 15727 3275 15764 3285
rect 15727 3257 15736 3275
rect 15754 3257 15764 3275
rect 15727 3248 15764 3257
rect 16077 3279 16115 3289
rect 15444 3237 15481 3238
rect 15394 3228 15481 3237
rect 15394 3208 15452 3228
rect 15472 3208 15481 3228
rect 15394 3198 15481 3208
rect 15540 3228 15577 3238
rect 15540 3208 15548 3228
rect 15568 3208 15577 3228
rect 15394 3197 15425 3198
rect 15540 3137 15577 3208
rect 15732 3183 15763 3248
rect 16077 3201 16112 3279
rect 16689 3269 16726 3292
rect 17482 3273 17513 3294
rect 17903 3273 17939 3294
rect 17325 3272 17362 3273
rect 16073 3192 16112 3201
rect 15731 3173 15768 3183
rect 15731 3171 15741 3173
rect 15665 3169 15741 3171
rect 15327 3113 15577 3137
rect 15662 3155 15741 3169
rect 15759 3155 15768 3173
rect 16073 3174 16083 3192
rect 16101 3174 16112 3192
rect 16073 3168 16112 3174
rect 16268 3244 16518 3268
rect 16268 3173 16305 3244
rect 16420 3183 16451 3184
rect 16073 3164 16110 3168
rect 15662 3152 15768 3155
rect 15134 3093 15155 3112
rect 15662 3093 15688 3152
rect 15731 3146 15768 3152
rect 16268 3153 16277 3173
rect 16297 3153 16305 3173
rect 16268 3143 16305 3153
rect 16364 3173 16451 3183
rect 16364 3153 16373 3173
rect 16393 3153 16451 3173
rect 16364 3144 16451 3153
rect 16364 3143 16401 3144
rect 16076 3093 16113 3102
rect 13788 3088 13888 3092
rect 13788 3084 13850 3088
rect 13788 3058 13795 3084
rect 13821 3062 13850 3084
rect 13876 3062 13888 3088
rect 13821 3058 13888 3062
rect 13788 3055 13888 3058
rect 13956 3055 13991 3092
rect 14053 3089 14412 3092
rect 14053 3084 14275 3089
rect 14053 3060 14066 3084
rect 14090 3065 14275 3084
rect 14299 3065 14412 3089
rect 14090 3060 14412 3065
rect 14053 3056 14412 3060
rect 14479 3084 14628 3092
rect 14479 3064 14490 3084
rect 14510 3064 14628 3084
rect 15134 3075 15688 3093
rect 15734 3082 15771 3084
rect 15662 3074 15688 3075
rect 15731 3074 15771 3082
rect 14479 3057 14628 3064
rect 15731 3062 15743 3074
rect 15722 3057 15743 3062
rect 14479 3056 14520 3057
rect 15138 3056 15743 3057
rect 15761 3056 15771 3074
rect 13803 3003 13840 3004
rect 13899 3003 13936 3004
rect 13955 3003 13991 3055
rect 14010 3003 14047 3004
rect 13703 2994 13841 3003
rect 13703 2974 13812 2994
rect 13832 2974 13841 2994
rect 13703 2967 13841 2974
rect 13899 2994 14047 3003
rect 13899 2974 13908 2994
rect 13928 2974 14018 2994
rect 14038 2974 14047 2994
rect 13703 2965 13799 2967
rect 13899 2964 14047 2974
rect 14106 2994 14143 3004
rect 14218 3003 14255 3004
rect 14199 3001 14255 3003
rect 14106 2974 14114 2994
rect 14134 2974 14143 2994
rect 13955 2963 13991 2964
rect 13803 2904 13840 2905
rect 14106 2904 14143 2974
rect 14168 2994 14255 3001
rect 14168 2991 14226 2994
rect 14168 2971 14173 2991
rect 14194 2974 14226 2991
rect 14246 2974 14255 2994
rect 14194 2971 14255 2974
rect 14168 2964 14255 2971
rect 14314 2994 14351 3004
rect 14314 2974 14322 2994
rect 14342 2974 14351 2994
rect 14168 2963 14199 2964
rect 13802 2903 14143 2904
rect 13727 2898 14143 2903
rect 13727 2878 13730 2898
rect 13750 2878 14143 2898
rect 14314 2903 14351 2974
rect 14381 3003 14412 3056
rect 15138 3047 15771 3056
rect 16074 3075 16085 3093
rect 16103 3075 16113 3093
rect 16420 3091 16451 3144
rect 16481 3173 16518 3244
rect 16689 3249 17082 3269
rect 17102 3249 17105 3269
rect 16689 3244 17105 3249
rect 17324 3263 17362 3272
rect 16689 3243 17030 3244
rect 17324 3243 17333 3263
rect 17353 3243 17362 3263
rect 16633 3183 16664 3184
rect 16481 3153 16490 3173
rect 16510 3153 16518 3173
rect 16481 3143 16518 3153
rect 16577 3176 16664 3183
rect 16577 3173 16638 3176
rect 16577 3153 16586 3173
rect 16606 3156 16638 3173
rect 16659 3156 16664 3176
rect 16606 3153 16664 3156
rect 16577 3146 16664 3153
rect 16689 3173 16726 3243
rect 16992 3242 17029 3243
rect 17324 3235 17362 3243
rect 17428 3267 17513 3273
rect 17538 3272 17575 3273
rect 17428 3247 17436 3267
rect 17456 3247 17513 3267
rect 17428 3239 17513 3247
rect 17537 3263 17575 3272
rect 17537 3243 17546 3263
rect 17566 3243 17575 3263
rect 17428 3238 17464 3239
rect 17537 3235 17575 3243
rect 17641 3267 17726 3273
rect 17746 3272 17783 3273
rect 17641 3247 17649 3267
rect 17669 3266 17726 3267
rect 17669 3247 17698 3266
rect 17641 3246 17698 3247
rect 17719 3246 17726 3266
rect 17641 3239 17726 3246
rect 17745 3263 17783 3272
rect 17745 3243 17754 3263
rect 17774 3243 17783 3263
rect 17641 3238 17677 3239
rect 17745 3235 17783 3243
rect 17849 3267 17993 3273
rect 17849 3247 17857 3267
rect 17877 3265 17965 3267
rect 17877 3248 17913 3265
rect 17937 3248 17965 3265
rect 17877 3247 17965 3248
rect 17985 3247 17993 3267
rect 17849 3239 17993 3247
rect 17849 3238 17885 3239
rect 17957 3238 17993 3239
rect 18059 3272 18096 3273
rect 18059 3271 18097 3272
rect 18059 3263 18123 3271
rect 18059 3243 18068 3263
rect 18088 3249 18123 3263
rect 18143 3249 18146 3269
rect 18088 3244 18146 3249
rect 18088 3243 18123 3244
rect 17325 3206 17362 3235
rect 17326 3204 17362 3206
rect 17538 3204 17575 3235
rect 16841 3183 16877 3184
rect 16689 3153 16698 3173
rect 16718 3153 16726 3173
rect 16577 3144 16633 3146
rect 16577 3143 16614 3144
rect 16689 3143 16726 3153
rect 16785 3173 16933 3183
rect 17326 3182 17575 3204
rect 17746 3203 17783 3235
rect 18059 3231 18123 3243
rect 18163 3205 18190 3383
rect 18022 3203 18190 3205
rect 17746 3192 18190 3203
rect 17033 3180 17129 3182
rect 16785 3153 16794 3173
rect 16814 3153 16904 3173
rect 16924 3153 16933 3173
rect 16785 3144 16933 3153
rect 16991 3173 17129 3180
rect 17746 3177 18192 3192
rect 18022 3176 18192 3177
rect 16991 3153 17000 3173
rect 17020 3153 17129 3173
rect 16991 3144 17129 3153
rect 16785 3143 16822 3144
rect 16841 3092 16877 3144
rect 16896 3143 16933 3144
rect 16992 3143 17029 3144
rect 16312 3090 16353 3091
rect 15138 3040 15770 3047
rect 15138 3038 15200 3040
rect 14716 3028 14884 3029
rect 15138 3028 15160 3038
rect 14431 3003 14468 3004
rect 14381 2994 14468 3003
rect 14381 2974 14439 2994
rect 14459 2974 14468 2994
rect 14381 2964 14468 2974
rect 14527 2994 14564 3004
rect 14527 2974 14535 2994
rect 14555 2974 14564 2994
rect 14381 2963 14412 2964
rect 14527 2903 14564 2974
rect 14314 2879 14564 2903
rect 14716 3002 15160 3028
rect 14716 3000 14884 3002
rect 14716 2822 14743 3000
rect 14783 2962 14847 2974
rect 15123 2970 15160 3002
rect 15331 3001 15580 3023
rect 15331 2970 15368 3001
rect 15544 2999 15580 3001
rect 15544 2970 15581 2999
rect 14783 2961 14818 2962
rect 14760 2956 14818 2961
rect 14760 2936 14763 2956
rect 14783 2942 14818 2956
rect 14838 2942 14847 2962
rect 14783 2934 14847 2942
rect 14809 2933 14847 2934
rect 14810 2932 14847 2933
rect 14913 2966 14949 2967
rect 15021 2966 15057 2967
rect 14913 2958 15057 2966
rect 14913 2938 14921 2958
rect 14941 2938 14970 2958
rect 14913 2937 14970 2938
rect 14992 2938 15029 2958
rect 15049 2938 15057 2958
rect 14992 2937 15057 2938
rect 14913 2932 15057 2937
rect 15123 2962 15161 2970
rect 15229 2966 15265 2967
rect 15123 2942 15132 2962
rect 15152 2942 15161 2962
rect 15123 2933 15161 2942
rect 15180 2959 15265 2966
rect 15180 2939 15187 2959
rect 15208 2958 15265 2959
rect 15208 2939 15237 2958
rect 15180 2938 15237 2939
rect 15257 2938 15265 2958
rect 15123 2932 15160 2933
rect 15180 2932 15265 2938
rect 15331 2962 15369 2970
rect 15442 2966 15478 2967
rect 15331 2942 15340 2962
rect 15360 2942 15369 2962
rect 15331 2933 15369 2942
rect 15393 2958 15478 2966
rect 15393 2938 15450 2958
rect 15470 2938 15478 2958
rect 15331 2932 15368 2933
rect 15393 2932 15478 2938
rect 15544 2962 15582 2970
rect 15544 2942 15553 2962
rect 15573 2942 15582 2962
rect 15544 2933 15582 2942
rect 15544 2932 15581 2933
rect 14967 2911 15003 2932
rect 15393 2911 15424 2932
rect 14800 2907 14900 2911
rect 14800 2903 14862 2907
rect 14800 2877 14807 2903
rect 14833 2881 14862 2903
rect 14888 2881 14900 2907
rect 14833 2877 14900 2881
rect 14800 2874 14900 2877
rect 14968 2874 15003 2911
rect 15065 2908 15424 2911
rect 15065 2903 15287 2908
rect 15065 2879 15078 2903
rect 15102 2884 15287 2903
rect 15311 2884 15424 2908
rect 15102 2879 15424 2884
rect 15065 2875 15424 2879
rect 15491 2903 15640 2911
rect 15491 2883 15502 2903
rect 15522 2883 15640 2903
rect 15491 2876 15640 2883
rect 15731 2891 15770 3040
rect 16074 2926 16113 3075
rect 16204 3083 16353 3090
rect 16204 3063 16322 3083
rect 16342 3063 16353 3083
rect 16204 3055 16353 3063
rect 16420 3087 16779 3091
rect 16420 3082 16742 3087
rect 16420 3058 16533 3082
rect 16557 3063 16742 3082
rect 16766 3063 16779 3087
rect 16557 3058 16779 3063
rect 16420 3055 16779 3058
rect 16841 3055 16876 3092
rect 16944 3089 17044 3092
rect 16944 3085 17011 3089
rect 16944 3059 16956 3085
rect 16982 3063 17011 3085
rect 17037 3063 17044 3089
rect 16982 3059 17044 3063
rect 16944 3055 17044 3059
rect 16420 3034 16451 3055
rect 16841 3034 16877 3055
rect 16263 3033 16300 3034
rect 16262 3024 16300 3033
rect 16262 3004 16271 3024
rect 16291 3004 16300 3024
rect 16262 2996 16300 3004
rect 16366 3028 16451 3034
rect 16476 3033 16513 3034
rect 16366 3008 16374 3028
rect 16394 3008 16451 3028
rect 16366 3000 16451 3008
rect 16475 3024 16513 3033
rect 16475 3004 16484 3024
rect 16504 3004 16513 3024
rect 16366 2999 16402 3000
rect 16475 2996 16513 3004
rect 16579 3028 16664 3034
rect 16684 3033 16721 3034
rect 16579 3008 16587 3028
rect 16607 3027 16664 3028
rect 16607 3008 16636 3027
rect 16579 3007 16636 3008
rect 16657 3007 16664 3027
rect 16579 3000 16664 3007
rect 16683 3024 16721 3033
rect 16683 3004 16692 3024
rect 16712 3004 16721 3024
rect 16579 2999 16615 3000
rect 16683 2996 16721 3004
rect 16787 3029 16931 3034
rect 16787 3028 16852 3029
rect 16787 3008 16795 3028
rect 16815 3008 16852 3028
rect 16874 3028 16931 3029
rect 16874 3008 16903 3028
rect 16923 3008 16931 3028
rect 16787 3000 16931 3008
rect 16787 2999 16823 3000
rect 16895 2999 16931 3000
rect 16997 3033 17034 3034
rect 16997 3032 17035 3033
rect 16997 3024 17061 3032
rect 16997 3004 17006 3024
rect 17026 3010 17061 3024
rect 17081 3010 17084 3030
rect 17026 3005 17084 3010
rect 17026 3004 17061 3005
rect 16263 2967 16300 2996
rect 16264 2965 16300 2967
rect 16476 2965 16513 2996
rect 16264 2943 16513 2965
rect 16684 2964 16721 2996
rect 16997 2992 17061 3004
rect 17101 2966 17128 3144
rect 16960 2964 17128 2966
rect 16684 2938 17128 2964
rect 17280 3063 17530 3087
rect 17280 2992 17317 3063
rect 17432 3002 17463 3003
rect 17280 2972 17289 2992
rect 17309 2972 17317 2992
rect 17280 2962 17317 2972
rect 17376 2992 17463 3002
rect 17376 2972 17385 2992
rect 17405 2972 17463 2992
rect 17376 2963 17463 2972
rect 17376 2962 17413 2963
rect 16684 2928 16706 2938
rect 16960 2937 17128 2938
rect 16644 2926 16706 2928
rect 16074 2919 16706 2926
rect 15491 2875 15532 2876
rect 14815 2822 14852 2823
rect 14911 2822 14948 2823
rect 14967 2822 15003 2874
rect 15022 2822 15059 2823
rect 14715 2813 14853 2822
rect 14715 2793 14824 2813
rect 14844 2793 14853 2813
rect 14715 2786 14853 2793
rect 14911 2813 15059 2822
rect 14911 2793 14920 2813
rect 14940 2793 15030 2813
rect 15050 2793 15059 2813
rect 14715 2784 14811 2786
rect 14911 2783 15059 2793
rect 15118 2813 15155 2823
rect 15230 2822 15267 2823
rect 15211 2820 15267 2822
rect 15118 2793 15126 2813
rect 15146 2793 15155 2813
rect 14967 2782 15003 2783
rect 13496 2742 13664 2743
rect 13496 2716 13940 2742
rect 13496 2714 13664 2716
rect 13496 2536 13523 2714
rect 13563 2676 13627 2688
rect 13903 2684 13940 2716
rect 14111 2715 14360 2737
rect 14815 2723 14852 2724
rect 15118 2723 15155 2793
rect 15180 2813 15267 2820
rect 15180 2810 15238 2813
rect 15180 2790 15185 2810
rect 15206 2793 15238 2810
rect 15258 2793 15267 2813
rect 15206 2790 15267 2793
rect 15180 2783 15267 2790
rect 15326 2813 15363 2823
rect 15326 2793 15334 2813
rect 15354 2793 15363 2813
rect 15180 2782 15211 2783
rect 14814 2722 15155 2723
rect 14111 2684 14148 2715
rect 14324 2713 14360 2715
rect 14739 2717 15155 2722
rect 14324 2684 14361 2713
rect 14739 2697 14742 2717
rect 14762 2697 15155 2717
rect 15326 2722 15363 2793
rect 15393 2822 15424 2875
rect 15731 2873 15741 2891
rect 15759 2873 15770 2891
rect 16073 2910 16706 2919
rect 17432 2910 17463 2963
rect 17493 2992 17530 3063
rect 17701 3068 18094 3088
rect 18114 3068 18117 3088
rect 17701 3063 18117 3068
rect 17701 3062 18042 3063
rect 17645 3002 17676 3003
rect 17493 2972 17502 2992
rect 17522 2972 17530 2992
rect 17493 2962 17530 2972
rect 17589 2995 17676 3002
rect 17589 2992 17650 2995
rect 17589 2972 17598 2992
rect 17618 2975 17650 2992
rect 17671 2975 17676 2995
rect 17618 2972 17676 2975
rect 17589 2965 17676 2972
rect 17701 2992 17738 3062
rect 18004 3061 18041 3062
rect 17853 3002 17889 3003
rect 17701 2972 17710 2992
rect 17730 2972 17738 2992
rect 17589 2963 17645 2965
rect 17589 2962 17626 2963
rect 17701 2962 17738 2972
rect 17797 2992 17945 3002
rect 18045 2999 18141 3001
rect 17797 2972 17806 2992
rect 17826 2972 17916 2992
rect 17936 2972 17945 2992
rect 17797 2963 17945 2972
rect 18003 2992 18141 2999
rect 18003 2972 18012 2992
rect 18032 2972 18141 2992
rect 18003 2963 18141 2972
rect 17797 2962 17834 2963
rect 17853 2911 17889 2963
rect 17908 2962 17945 2963
rect 18004 2962 18041 2963
rect 16073 2892 16083 2910
rect 16101 2909 16706 2910
rect 17324 2909 17365 2910
rect 16101 2904 16122 2909
rect 16101 2892 16113 2904
rect 17216 2902 17365 2909
rect 16073 2884 16113 2892
rect 16156 2891 16182 2892
rect 16073 2882 16110 2884
rect 16156 2873 16710 2891
rect 17216 2882 17334 2902
rect 17354 2882 17365 2902
rect 17216 2874 17365 2882
rect 17432 2906 17791 2910
rect 17432 2901 17754 2906
rect 17432 2877 17545 2901
rect 17569 2882 17754 2901
rect 17778 2882 17791 2906
rect 17569 2877 17791 2882
rect 17432 2874 17791 2877
rect 17853 2874 17888 2911
rect 17956 2908 18056 2911
rect 17956 2904 18023 2908
rect 17956 2878 17968 2904
rect 17994 2882 18023 2904
rect 18049 2882 18056 2908
rect 17994 2878 18056 2882
rect 17956 2874 18056 2878
rect 15731 2864 15768 2873
rect 15443 2822 15480 2823
rect 15393 2813 15480 2822
rect 15393 2793 15451 2813
rect 15471 2793 15480 2813
rect 15393 2783 15480 2793
rect 15539 2813 15576 2823
rect 15539 2793 15547 2813
rect 15567 2793 15576 2813
rect 16076 2814 16113 2820
rect 16156 2814 16182 2873
rect 16689 2854 16710 2873
rect 16076 2811 16182 2814
rect 15734 2798 15771 2802
rect 15393 2782 15424 2783
rect 15539 2722 15576 2793
rect 15326 2698 15576 2722
rect 15732 2792 15771 2798
rect 15732 2774 15743 2792
rect 15761 2774 15771 2792
rect 16076 2793 16085 2811
rect 16103 2797 16182 2811
rect 16267 2829 16517 2853
rect 16103 2795 16179 2797
rect 16103 2793 16113 2795
rect 16076 2783 16113 2793
rect 15732 2765 15771 2774
rect 13563 2675 13598 2676
rect 13540 2670 13598 2675
rect 13540 2650 13543 2670
rect 13563 2656 13598 2670
rect 13618 2656 13627 2676
rect 13563 2648 13627 2656
rect 13589 2647 13627 2648
rect 13590 2646 13627 2647
rect 13693 2680 13729 2681
rect 13801 2680 13837 2681
rect 13693 2674 13837 2680
rect 13693 2672 13754 2674
rect 13693 2652 13701 2672
rect 13721 2652 13754 2672
rect 13693 2648 13754 2652
rect 13779 2672 13837 2674
rect 13779 2652 13809 2672
rect 13829 2652 13837 2672
rect 13779 2648 13837 2652
rect 13693 2646 13837 2648
rect 13903 2676 13941 2684
rect 14009 2680 14045 2681
rect 13903 2656 13912 2676
rect 13932 2656 13941 2676
rect 13903 2647 13941 2656
rect 13960 2673 14045 2680
rect 13960 2653 13967 2673
rect 13988 2672 14045 2673
rect 13988 2653 14017 2672
rect 13960 2652 14017 2653
rect 14037 2652 14045 2672
rect 13903 2646 13940 2647
rect 13960 2646 14045 2652
rect 14111 2676 14149 2684
rect 14222 2680 14258 2681
rect 14111 2656 14120 2676
rect 14140 2656 14149 2676
rect 14111 2647 14149 2656
rect 14173 2672 14258 2680
rect 14173 2652 14230 2672
rect 14250 2652 14258 2672
rect 14111 2646 14148 2647
rect 14173 2646 14258 2652
rect 14324 2676 14362 2684
rect 14324 2656 14333 2676
rect 14353 2656 14362 2676
rect 14324 2647 14362 2656
rect 15118 2674 15155 2697
rect 15732 2687 15767 2765
rect 16081 2718 16112 2783
rect 16267 2758 16304 2829
rect 16419 2768 16450 2769
rect 16267 2738 16276 2758
rect 16296 2738 16304 2758
rect 16267 2728 16304 2738
rect 16363 2758 16450 2768
rect 16363 2738 16372 2758
rect 16392 2738 16450 2758
rect 16363 2729 16450 2738
rect 16363 2728 16400 2729
rect 15729 2677 15767 2687
rect 16080 2709 16117 2718
rect 16080 2691 16090 2709
rect 16108 2691 16117 2709
rect 16080 2681 16117 2691
rect 15118 2673 15288 2674
rect 15729 2673 15739 2677
rect 15118 2659 15739 2673
rect 15757 2659 15767 2677
rect 16419 2676 16450 2729
rect 16480 2758 16517 2829
rect 16688 2834 17081 2854
rect 17101 2834 17104 2854
rect 17432 2853 17463 2874
rect 17853 2853 17889 2874
rect 17275 2852 17312 2853
rect 16688 2829 17104 2834
rect 17274 2843 17312 2852
rect 16688 2828 17029 2829
rect 16632 2768 16663 2769
rect 16480 2738 16489 2758
rect 16509 2738 16517 2758
rect 16480 2728 16517 2738
rect 16576 2761 16663 2768
rect 16576 2758 16637 2761
rect 16576 2738 16585 2758
rect 16605 2741 16637 2758
rect 16658 2741 16663 2761
rect 16605 2738 16663 2741
rect 16576 2731 16663 2738
rect 16688 2758 16725 2828
rect 16991 2827 17028 2828
rect 17274 2823 17283 2843
rect 17303 2823 17312 2843
rect 17274 2815 17312 2823
rect 17378 2847 17463 2853
rect 17488 2852 17525 2853
rect 17378 2827 17386 2847
rect 17406 2827 17463 2847
rect 17378 2819 17463 2827
rect 17487 2843 17525 2852
rect 17487 2823 17496 2843
rect 17516 2823 17525 2843
rect 17378 2818 17414 2819
rect 17487 2815 17525 2823
rect 17591 2847 17676 2853
rect 17696 2852 17733 2853
rect 17591 2827 17599 2847
rect 17619 2846 17676 2847
rect 17619 2827 17648 2846
rect 17591 2826 17648 2827
rect 17669 2826 17676 2846
rect 17591 2819 17676 2826
rect 17695 2843 17733 2852
rect 17695 2823 17704 2843
rect 17724 2823 17733 2843
rect 17591 2818 17627 2819
rect 17695 2815 17733 2823
rect 17799 2848 17943 2853
rect 17799 2847 17858 2848
rect 17799 2827 17807 2847
rect 17827 2828 17858 2847
rect 17882 2847 17943 2848
rect 17882 2828 17915 2847
rect 17827 2827 17915 2828
rect 17935 2827 17943 2847
rect 17799 2819 17943 2827
rect 17799 2818 17835 2819
rect 17907 2818 17943 2819
rect 18009 2852 18046 2853
rect 18009 2851 18047 2852
rect 18009 2843 18073 2851
rect 18009 2823 18018 2843
rect 18038 2829 18073 2843
rect 18093 2829 18096 2849
rect 18038 2824 18096 2829
rect 18038 2823 18073 2824
rect 17275 2786 17312 2815
rect 17276 2784 17312 2786
rect 17488 2784 17525 2815
rect 16840 2768 16876 2769
rect 16688 2738 16697 2758
rect 16717 2738 16725 2758
rect 16576 2729 16632 2731
rect 16576 2728 16613 2729
rect 16688 2728 16725 2738
rect 16784 2758 16932 2768
rect 17032 2765 17128 2767
rect 16784 2738 16793 2758
rect 16813 2738 16903 2758
rect 16923 2738 16932 2758
rect 16784 2729 16932 2738
rect 16990 2758 17128 2765
rect 17276 2762 17525 2784
rect 17696 2783 17733 2815
rect 18009 2811 18073 2823
rect 18113 2785 18140 2963
rect 17972 2783 18140 2785
rect 17696 2779 18140 2783
rect 16990 2738 16999 2758
rect 17019 2738 17128 2758
rect 17696 2760 17745 2779
rect 17765 2760 18140 2779
rect 17696 2757 18140 2760
rect 17972 2756 18140 2757
rect 18161 2782 18192 3176
rect 18161 2756 18166 2782
rect 18185 2756 18192 2782
rect 18161 2753 18192 2756
rect 16990 2729 17128 2738
rect 16784 2728 16821 2729
rect 16840 2677 16876 2729
rect 16895 2728 16932 2729
rect 16991 2728 17028 2729
rect 16311 2675 16352 2676
rect 15118 2653 15767 2659
rect 16203 2668 16352 2675
rect 15118 2652 15766 2653
rect 15729 2650 15766 2652
rect 16203 2648 16321 2668
rect 16341 2648 16352 2668
rect 14324 2646 14361 2647
rect 13747 2625 13783 2646
rect 14173 2625 14204 2646
rect 16203 2640 16352 2648
rect 16419 2672 16778 2676
rect 16419 2667 16741 2672
rect 16419 2643 16532 2667
rect 16556 2648 16741 2667
rect 16765 2648 16778 2672
rect 16556 2643 16778 2648
rect 16419 2640 16778 2643
rect 16840 2640 16875 2677
rect 16943 2674 17043 2677
rect 16943 2670 17010 2674
rect 16943 2644 16955 2670
rect 16981 2648 17010 2670
rect 17036 2648 17043 2674
rect 16981 2644 17043 2648
rect 16943 2640 17043 2644
rect 13580 2621 13680 2625
rect 13580 2617 13642 2621
rect 13580 2591 13587 2617
rect 13613 2595 13642 2617
rect 13668 2595 13680 2621
rect 13613 2591 13680 2595
rect 13580 2588 13680 2591
rect 13748 2588 13783 2625
rect 13845 2622 14204 2625
rect 13845 2617 14067 2622
rect 13845 2593 13858 2617
rect 13882 2598 14067 2617
rect 14091 2598 14204 2622
rect 13882 2593 14204 2598
rect 13845 2589 14204 2593
rect 14271 2617 14420 2625
rect 16419 2619 16450 2640
rect 16840 2619 16876 2640
rect 14271 2597 14282 2617
rect 14302 2597 14420 2617
rect 14271 2590 14420 2597
rect 16083 2610 16120 2619
rect 16262 2618 16299 2619
rect 16083 2592 16092 2610
rect 16110 2592 16120 2610
rect 14271 2589 14312 2590
rect 13595 2536 13632 2537
rect 13691 2536 13728 2537
rect 13747 2536 13783 2588
rect 13802 2536 13839 2537
rect 13495 2527 13633 2536
rect 13495 2507 13604 2527
rect 13624 2507 13633 2527
rect 13495 2500 13633 2507
rect 13691 2527 13839 2536
rect 13691 2507 13700 2527
rect 13720 2507 13810 2527
rect 13830 2507 13839 2527
rect 13495 2498 13591 2500
rect 13691 2497 13839 2507
rect 13898 2527 13935 2537
rect 14010 2536 14047 2537
rect 13991 2534 14047 2536
rect 13898 2507 13906 2527
rect 13926 2507 13935 2527
rect 13747 2496 13783 2497
rect 13595 2437 13632 2438
rect 13898 2437 13935 2507
rect 13960 2527 14047 2534
rect 13960 2524 14018 2527
rect 13960 2504 13965 2524
rect 13986 2507 14018 2524
rect 14038 2507 14047 2527
rect 13986 2504 14047 2507
rect 13960 2497 14047 2504
rect 14106 2527 14143 2537
rect 14106 2507 14114 2527
rect 14134 2507 14143 2527
rect 13960 2496 13991 2497
rect 13594 2436 13935 2437
rect 13519 2431 13935 2436
rect 13519 2411 13522 2431
rect 13542 2411 13935 2431
rect 14106 2436 14143 2507
rect 14173 2536 14204 2589
rect 15732 2578 15769 2588
rect 16083 2582 16120 2592
rect 15732 2560 15741 2578
rect 15759 2560 15769 2578
rect 15732 2551 15769 2560
rect 14223 2536 14260 2537
rect 14173 2527 14260 2536
rect 14173 2507 14231 2527
rect 14251 2507 14260 2527
rect 14173 2497 14260 2507
rect 14319 2527 14356 2537
rect 14319 2507 14327 2527
rect 14347 2507 14356 2527
rect 14173 2496 14204 2497
rect 14319 2436 14356 2507
rect 15732 2505 15767 2551
rect 16084 2547 16120 2582
rect 16261 2609 16299 2618
rect 16261 2589 16270 2609
rect 16290 2589 16299 2609
rect 16261 2581 16299 2589
rect 16365 2613 16450 2619
rect 16475 2618 16512 2619
rect 16365 2593 16373 2613
rect 16393 2593 16450 2613
rect 16365 2585 16450 2593
rect 16474 2609 16512 2618
rect 16474 2589 16483 2609
rect 16503 2589 16512 2609
rect 16365 2584 16401 2585
rect 16474 2581 16512 2589
rect 16578 2613 16663 2619
rect 16683 2618 16720 2619
rect 16578 2593 16586 2613
rect 16606 2612 16663 2613
rect 16606 2593 16635 2612
rect 16578 2592 16635 2593
rect 16656 2592 16663 2612
rect 16578 2585 16663 2592
rect 16682 2609 16720 2618
rect 16682 2589 16691 2609
rect 16711 2589 16720 2609
rect 16578 2584 16614 2585
rect 16682 2581 16720 2589
rect 16786 2613 16930 2619
rect 16786 2593 16794 2613
rect 16814 2612 16902 2613
rect 16814 2593 16842 2612
rect 16786 2591 16842 2593
rect 16864 2593 16902 2612
rect 16922 2593 16930 2613
rect 16864 2591 16930 2593
rect 16786 2585 16930 2591
rect 16786 2584 16822 2585
rect 16894 2584 16930 2585
rect 16996 2618 17033 2619
rect 16996 2617 17034 2618
rect 16996 2609 17060 2617
rect 16996 2589 17005 2609
rect 17025 2595 17060 2609
rect 17080 2595 17083 2615
rect 17025 2590 17083 2595
rect 17025 2589 17060 2590
rect 16262 2552 16299 2581
rect 16082 2506 16120 2547
rect 16263 2550 16299 2552
rect 16475 2550 16512 2581
rect 16263 2528 16512 2550
rect 16683 2549 16720 2581
rect 16996 2577 17060 2589
rect 17100 2551 17127 2729
rect 16959 2549 17127 2551
rect 16683 2523 17127 2549
rect 16684 2506 16708 2523
rect 16959 2522 17127 2523
rect 17495 2551 17745 2575
rect 15731 2499 15769 2505
rect 15142 2481 15769 2499
rect 16082 2488 16709 2506
rect 16082 2482 16120 2488
rect 14106 2412 14356 2436
rect 14724 2464 14892 2465
rect 15143 2464 15167 2481
rect 14724 2438 15168 2464
rect 14724 2436 14892 2438
rect 13104 2299 13137 2359
rect 12906 2292 13074 2294
rect 12630 2266 13074 2292
rect 12906 2265 13074 2266
rect 13103 2288 13140 2299
rect 13103 2269 13109 2288
rect 13132 2269 13140 2288
rect 11567 2225 11603 2226
rect 11415 2195 11424 2215
rect 11444 2195 11452 2215
rect 11303 2186 11359 2188
rect 11303 2185 11340 2186
rect 11415 2185 11452 2195
rect 11511 2215 11659 2225
rect 11759 2222 11855 2224
rect 11511 2195 11520 2215
rect 11540 2195 11630 2215
rect 11650 2195 11659 2215
rect 11511 2186 11659 2195
rect 11717 2215 11855 2222
rect 11717 2195 11726 2215
rect 11746 2195 11855 2215
rect 11717 2186 11855 2195
rect 11511 2185 11548 2186
rect 11567 2134 11603 2186
rect 11622 2185 11659 2186
rect 11718 2185 11755 2186
rect 11038 2132 11079 2133
rect 10361 2074 10398 2076
rect 10289 2066 10315 2067
rect 10358 2066 10398 2074
rect 9106 2049 9255 2056
rect 10358 2054 10370 2066
rect 10349 2049 10370 2054
rect 9106 2048 9147 2049
rect 9765 2048 10370 2049
rect 10388 2048 10398 2066
rect 8430 1995 8467 1996
rect 8526 1995 8563 1996
rect 8582 1995 8618 2047
rect 8637 1995 8674 1996
rect 8330 1986 8468 1995
rect 8330 1966 8439 1986
rect 8459 1966 8468 1986
rect 8330 1959 8468 1966
rect 8526 1986 8674 1995
rect 8526 1966 8535 1986
rect 8555 1966 8645 1986
rect 8665 1966 8674 1986
rect 8330 1957 8426 1959
rect 8526 1956 8674 1966
rect 8733 1986 8770 1996
rect 8845 1995 8882 1996
rect 8826 1993 8882 1995
rect 8733 1966 8741 1986
rect 8761 1966 8770 1986
rect 8582 1955 8618 1956
rect 8430 1896 8467 1897
rect 8733 1896 8770 1966
rect 8795 1986 8882 1993
rect 8795 1983 8853 1986
rect 8795 1963 8800 1983
rect 8821 1966 8853 1983
rect 8873 1966 8882 1986
rect 8821 1963 8882 1966
rect 8795 1956 8882 1963
rect 8941 1986 8978 1996
rect 8941 1966 8949 1986
rect 8969 1966 8978 1986
rect 8795 1955 8826 1956
rect 8429 1895 8770 1896
rect 8354 1890 8770 1895
rect 8354 1870 8357 1890
rect 8377 1870 8770 1890
rect 8941 1895 8978 1966
rect 9008 1995 9039 2048
rect 9765 2039 10398 2048
rect 9765 2032 10397 2039
rect 9765 2030 9827 2032
rect 9343 2020 9511 2021
rect 9765 2020 9787 2030
rect 9058 1995 9095 1996
rect 9008 1986 9095 1995
rect 9008 1966 9066 1986
rect 9086 1966 9095 1986
rect 9008 1956 9095 1966
rect 9154 1986 9191 1996
rect 9154 1966 9162 1986
rect 9182 1966 9191 1986
rect 9008 1955 9039 1956
rect 9154 1895 9191 1966
rect 8941 1871 9191 1895
rect 9343 1994 9787 2020
rect 9343 1992 9511 1994
rect 9343 1814 9370 1992
rect 9410 1954 9474 1966
rect 9750 1962 9787 1994
rect 9958 1993 10207 2015
rect 9958 1962 9995 1993
rect 10171 1991 10207 1993
rect 10171 1962 10208 1991
rect 9410 1953 9445 1954
rect 9387 1948 9445 1953
rect 9387 1928 9390 1948
rect 9410 1934 9445 1948
rect 9465 1934 9474 1954
rect 9410 1926 9474 1934
rect 9436 1925 9474 1926
rect 9437 1924 9474 1925
rect 9540 1958 9576 1959
rect 9648 1958 9684 1959
rect 9540 1950 9684 1958
rect 9540 1930 9548 1950
rect 9568 1930 9597 1950
rect 9540 1929 9597 1930
rect 9619 1930 9656 1950
rect 9676 1930 9684 1950
rect 9619 1929 9684 1930
rect 9540 1924 9684 1929
rect 9750 1954 9788 1962
rect 9856 1958 9892 1959
rect 9750 1934 9759 1954
rect 9779 1934 9788 1954
rect 9750 1925 9788 1934
rect 9807 1951 9892 1958
rect 9807 1931 9814 1951
rect 9835 1950 9892 1951
rect 9835 1931 9864 1950
rect 9807 1930 9864 1931
rect 9884 1930 9892 1950
rect 9750 1924 9787 1925
rect 9807 1924 9892 1930
rect 9958 1954 9996 1962
rect 10069 1958 10105 1959
rect 9958 1934 9967 1954
rect 9987 1934 9996 1954
rect 9958 1925 9996 1934
rect 10020 1950 10105 1958
rect 10020 1930 10077 1950
rect 10097 1930 10105 1950
rect 9958 1924 9995 1925
rect 10020 1924 10105 1930
rect 10171 1954 10209 1962
rect 10171 1934 10180 1954
rect 10200 1934 10209 1954
rect 10171 1925 10209 1934
rect 10171 1924 10208 1925
rect 9594 1903 9630 1924
rect 10020 1903 10051 1924
rect 9427 1899 9527 1903
rect 9427 1895 9489 1899
rect 9427 1869 9434 1895
rect 9460 1873 9489 1895
rect 9515 1873 9527 1899
rect 9460 1869 9527 1873
rect 9427 1866 9527 1869
rect 9595 1866 9630 1903
rect 9692 1900 10051 1903
rect 9692 1895 9914 1900
rect 9692 1871 9705 1895
rect 9729 1876 9914 1895
rect 9938 1876 10051 1900
rect 9729 1871 10051 1876
rect 9692 1867 10051 1871
rect 10118 1895 10267 1903
rect 10118 1875 10129 1895
rect 10149 1875 10267 1895
rect 10118 1868 10267 1875
rect 10358 1883 10397 2032
rect 10800 1968 10839 2117
rect 10930 2125 11079 2132
rect 10930 2105 11048 2125
rect 11068 2105 11079 2125
rect 10930 2097 11079 2105
rect 11146 2129 11505 2133
rect 11146 2124 11468 2129
rect 11146 2100 11259 2124
rect 11283 2105 11468 2124
rect 11492 2105 11505 2129
rect 11283 2100 11505 2105
rect 11146 2097 11505 2100
rect 11567 2097 11602 2134
rect 11670 2131 11770 2134
rect 11670 2127 11737 2131
rect 11670 2101 11682 2127
rect 11708 2105 11737 2127
rect 11763 2105 11770 2131
rect 11708 2101 11770 2105
rect 11670 2097 11770 2101
rect 11146 2076 11177 2097
rect 11567 2076 11603 2097
rect 10989 2075 11026 2076
rect 10988 2066 11026 2075
rect 10988 2046 10997 2066
rect 11017 2046 11026 2066
rect 10988 2038 11026 2046
rect 11092 2070 11177 2076
rect 11202 2075 11239 2076
rect 11092 2050 11100 2070
rect 11120 2050 11177 2070
rect 11092 2042 11177 2050
rect 11201 2066 11239 2075
rect 11201 2046 11210 2066
rect 11230 2046 11239 2066
rect 11092 2041 11128 2042
rect 11201 2038 11239 2046
rect 11305 2070 11390 2076
rect 11410 2075 11447 2076
rect 11305 2050 11313 2070
rect 11333 2069 11390 2070
rect 11333 2050 11362 2069
rect 11305 2049 11362 2050
rect 11383 2049 11390 2069
rect 11305 2042 11390 2049
rect 11409 2066 11447 2075
rect 11409 2046 11418 2066
rect 11438 2046 11447 2066
rect 11305 2041 11341 2042
rect 11409 2038 11447 2046
rect 11513 2071 11657 2076
rect 11513 2070 11578 2071
rect 11513 2050 11521 2070
rect 11541 2050 11578 2070
rect 11600 2070 11657 2071
rect 11600 2050 11629 2070
rect 11649 2050 11657 2070
rect 11513 2042 11657 2050
rect 11513 2041 11549 2042
rect 11621 2041 11657 2042
rect 11723 2075 11760 2076
rect 11723 2074 11761 2075
rect 11723 2066 11787 2074
rect 11723 2046 11732 2066
rect 11752 2052 11787 2066
rect 11807 2052 11810 2072
rect 11752 2047 11810 2052
rect 11752 2046 11787 2047
rect 10989 2009 11026 2038
rect 10990 2007 11026 2009
rect 11202 2007 11239 2038
rect 10990 1985 11239 2007
rect 11410 2006 11447 2038
rect 11723 2034 11787 2046
rect 11827 2008 11854 2186
rect 11686 2006 11854 2008
rect 11410 1980 11854 2006
rect 12006 2105 12256 2129
rect 12006 2034 12043 2105
rect 12158 2044 12189 2045
rect 12006 2014 12015 2034
rect 12035 2014 12043 2034
rect 12006 2004 12043 2014
rect 12102 2034 12189 2044
rect 12102 2014 12111 2034
rect 12131 2014 12189 2034
rect 12102 2005 12189 2014
rect 12102 2004 12139 2005
rect 11410 1970 11432 1980
rect 11686 1979 11854 1980
rect 11370 1968 11432 1970
rect 10800 1961 11432 1968
rect 10799 1952 11432 1961
rect 12158 1952 12189 2005
rect 12219 2034 12256 2105
rect 12427 2110 12820 2130
rect 12840 2110 12843 2130
rect 12427 2105 12843 2110
rect 12427 2104 12768 2105
rect 12371 2044 12402 2045
rect 12219 2014 12228 2034
rect 12248 2014 12256 2034
rect 12219 2004 12256 2014
rect 12315 2037 12402 2044
rect 12315 2034 12376 2037
rect 12315 2014 12324 2034
rect 12344 2017 12376 2034
rect 12397 2017 12402 2037
rect 12344 2014 12402 2017
rect 12315 2007 12402 2014
rect 12427 2034 12464 2104
rect 12730 2103 12767 2104
rect 12579 2044 12615 2045
rect 12427 2014 12436 2034
rect 12456 2014 12464 2034
rect 12315 2005 12371 2007
rect 12315 2004 12352 2005
rect 12427 2004 12464 2014
rect 12523 2034 12671 2044
rect 12771 2041 12867 2043
rect 12523 2014 12532 2034
rect 12552 2014 12642 2034
rect 12662 2014 12671 2034
rect 12523 2005 12671 2014
rect 12729 2034 12867 2041
rect 12729 2014 12738 2034
rect 12758 2014 12867 2034
rect 12729 2005 12867 2014
rect 12523 2004 12560 2005
rect 12579 1953 12615 2005
rect 12634 2004 12671 2005
rect 12730 2004 12767 2005
rect 10799 1934 10809 1952
rect 10827 1951 11432 1952
rect 12050 1951 12091 1952
rect 10827 1946 10848 1951
rect 10827 1934 10839 1946
rect 11942 1944 12091 1951
rect 10799 1926 10839 1934
rect 10882 1933 10908 1934
rect 10799 1924 10836 1926
rect 10118 1867 10159 1868
rect 9442 1814 9479 1815
rect 9538 1814 9575 1815
rect 9594 1814 9630 1866
rect 9649 1814 9686 1815
rect 9342 1805 9480 1814
rect 9342 1785 9451 1805
rect 9471 1785 9480 1805
rect 8279 1781 8449 1782
rect 8279 1766 8725 1781
rect 9342 1778 9480 1785
rect 9538 1805 9686 1814
rect 9538 1785 9547 1805
rect 9567 1785 9657 1805
rect 9677 1785 9686 1805
rect 9342 1776 9438 1778
rect 8281 1755 8725 1766
rect 8281 1753 8449 1755
rect 8281 1575 8308 1753
rect 8348 1715 8412 1727
rect 8688 1723 8725 1755
rect 8896 1754 9145 1776
rect 9538 1775 9686 1785
rect 9745 1805 9782 1815
rect 9857 1814 9894 1815
rect 9838 1812 9894 1814
rect 9745 1785 9753 1805
rect 9773 1785 9782 1805
rect 9594 1774 9630 1775
rect 8896 1723 8933 1754
rect 9109 1752 9145 1754
rect 9109 1723 9146 1752
rect 8348 1714 8383 1715
rect 8325 1709 8383 1714
rect 8325 1689 8328 1709
rect 8348 1695 8383 1709
rect 8403 1695 8412 1715
rect 8348 1687 8412 1695
rect 8374 1686 8412 1687
rect 8375 1685 8412 1686
rect 8478 1719 8514 1720
rect 8586 1719 8622 1720
rect 8478 1711 8622 1719
rect 8478 1691 8486 1711
rect 8506 1710 8594 1711
rect 8506 1693 8534 1710
rect 8558 1693 8594 1710
rect 8506 1691 8594 1693
rect 8614 1691 8622 1711
rect 8478 1685 8622 1691
rect 8688 1715 8726 1723
rect 8794 1719 8830 1720
rect 8688 1695 8697 1715
rect 8717 1695 8726 1715
rect 8688 1686 8726 1695
rect 8745 1712 8830 1719
rect 8745 1692 8752 1712
rect 8773 1711 8830 1712
rect 8773 1692 8802 1711
rect 8745 1691 8802 1692
rect 8822 1691 8830 1711
rect 8688 1685 8725 1686
rect 8745 1685 8830 1691
rect 8896 1715 8934 1723
rect 9007 1719 9043 1720
rect 8896 1695 8905 1715
rect 8925 1695 8934 1715
rect 8896 1686 8934 1695
rect 8958 1711 9043 1719
rect 8958 1691 9015 1711
rect 9035 1691 9043 1711
rect 8896 1685 8933 1686
rect 8958 1685 9043 1691
rect 9109 1715 9147 1723
rect 9442 1715 9479 1716
rect 9745 1715 9782 1785
rect 9807 1805 9894 1812
rect 9807 1802 9865 1805
rect 9807 1782 9812 1802
rect 9833 1785 9865 1802
rect 9885 1785 9894 1805
rect 9833 1782 9894 1785
rect 9807 1775 9894 1782
rect 9953 1805 9990 1815
rect 9953 1785 9961 1805
rect 9981 1785 9990 1805
rect 9807 1774 9838 1775
rect 9109 1695 9118 1715
rect 9138 1695 9147 1715
rect 9441 1714 9782 1715
rect 9109 1686 9147 1695
rect 9366 1709 9782 1714
rect 9366 1689 9369 1709
rect 9389 1689 9782 1709
rect 9953 1714 9990 1785
rect 10020 1814 10051 1867
rect 10358 1865 10368 1883
rect 10386 1865 10397 1883
rect 10882 1915 11436 1933
rect 11942 1924 12060 1944
rect 12080 1924 12091 1944
rect 11942 1916 12091 1924
rect 12158 1948 12517 1952
rect 12158 1943 12480 1948
rect 12158 1919 12271 1943
rect 12295 1924 12480 1943
rect 12504 1924 12517 1948
rect 12295 1919 12517 1924
rect 12158 1916 12517 1919
rect 12579 1916 12614 1953
rect 12682 1950 12782 1953
rect 12682 1946 12749 1950
rect 12682 1920 12694 1946
rect 12720 1924 12749 1946
rect 12775 1924 12782 1950
rect 12720 1920 12782 1924
rect 12682 1916 12782 1920
rect 10358 1856 10395 1865
rect 10802 1856 10839 1862
rect 10882 1856 10908 1915
rect 11415 1896 11436 1915
rect 10802 1853 10908 1856
rect 10802 1835 10811 1853
rect 10829 1839 10908 1853
rect 10993 1871 11243 1895
rect 10829 1837 10905 1839
rect 10829 1835 10839 1837
rect 10802 1825 10839 1835
rect 10070 1814 10107 1815
rect 10020 1805 10107 1814
rect 10020 1785 10078 1805
rect 10098 1785 10107 1805
rect 10020 1775 10107 1785
rect 10166 1805 10203 1815
rect 10166 1785 10174 1805
rect 10194 1785 10203 1805
rect 10361 1790 10398 1794
rect 10020 1774 10051 1775
rect 10166 1714 10203 1785
rect 9953 1690 10203 1714
rect 10359 1784 10398 1790
rect 10359 1766 10370 1784
rect 10388 1766 10398 1784
rect 10359 1757 10398 1766
rect 10807 1760 10838 1825
rect 10993 1800 11030 1871
rect 11145 1810 11176 1811
rect 10993 1780 11002 1800
rect 11022 1780 11030 1800
rect 10993 1770 11030 1780
rect 11089 1800 11176 1810
rect 11089 1780 11098 1800
rect 11118 1780 11176 1800
rect 11089 1771 11176 1780
rect 11089 1770 11126 1771
rect 9109 1685 9146 1686
rect 8532 1664 8568 1685
rect 8958 1664 8989 1685
rect 9745 1666 9782 1689
rect 10359 1679 10394 1757
rect 10806 1751 10843 1760
rect 10806 1733 10816 1751
rect 10834 1733 10843 1751
rect 10806 1723 10843 1733
rect 11145 1718 11176 1771
rect 11206 1800 11243 1871
rect 11414 1876 11807 1896
rect 11827 1876 11830 1896
rect 12158 1895 12189 1916
rect 12579 1895 12615 1916
rect 12001 1894 12038 1895
rect 11414 1871 11830 1876
rect 12000 1885 12038 1894
rect 11414 1870 11755 1871
rect 11358 1810 11389 1811
rect 11206 1780 11215 1800
rect 11235 1780 11243 1800
rect 11206 1770 11243 1780
rect 11302 1803 11389 1810
rect 11302 1800 11363 1803
rect 11302 1780 11311 1800
rect 11331 1783 11363 1800
rect 11384 1783 11389 1803
rect 11331 1780 11389 1783
rect 11302 1773 11389 1780
rect 11414 1800 11451 1870
rect 11717 1869 11754 1870
rect 12000 1865 12009 1885
rect 12029 1865 12038 1885
rect 12000 1857 12038 1865
rect 12104 1889 12189 1895
rect 12214 1894 12251 1895
rect 12104 1869 12112 1889
rect 12132 1869 12189 1889
rect 12104 1861 12189 1869
rect 12213 1885 12251 1894
rect 12213 1865 12222 1885
rect 12242 1865 12251 1885
rect 12104 1860 12140 1861
rect 12213 1857 12251 1865
rect 12317 1889 12402 1895
rect 12422 1894 12459 1895
rect 12317 1869 12325 1889
rect 12345 1888 12402 1889
rect 12345 1869 12374 1888
rect 12317 1868 12374 1869
rect 12395 1868 12402 1888
rect 12317 1861 12402 1868
rect 12421 1885 12459 1894
rect 12421 1865 12430 1885
rect 12450 1865 12459 1885
rect 12317 1860 12353 1861
rect 12421 1857 12459 1865
rect 12525 1889 12669 1895
rect 12525 1869 12533 1889
rect 12553 1869 12585 1889
rect 12609 1869 12641 1889
rect 12661 1869 12669 1889
rect 12525 1861 12669 1869
rect 12525 1860 12561 1861
rect 12633 1860 12669 1861
rect 12735 1894 12772 1895
rect 12735 1893 12773 1894
rect 12735 1885 12799 1893
rect 12735 1865 12744 1885
rect 12764 1871 12799 1885
rect 12819 1871 12822 1891
rect 12764 1866 12822 1871
rect 12764 1865 12799 1866
rect 12001 1828 12038 1857
rect 12002 1826 12038 1828
rect 12214 1826 12251 1857
rect 11566 1810 11602 1811
rect 11414 1780 11423 1800
rect 11443 1780 11451 1800
rect 11302 1771 11358 1773
rect 11302 1770 11339 1771
rect 11414 1770 11451 1780
rect 11510 1800 11658 1810
rect 11758 1807 11854 1809
rect 11510 1780 11519 1800
rect 11539 1780 11629 1800
rect 11649 1780 11658 1800
rect 11510 1771 11658 1780
rect 11716 1800 11854 1807
rect 12002 1804 12251 1826
rect 12422 1825 12459 1857
rect 12735 1853 12799 1865
rect 12839 1827 12866 2005
rect 12698 1825 12866 1827
rect 12422 1821 12866 1825
rect 11716 1780 11725 1800
rect 11745 1780 11854 1800
rect 12422 1802 12471 1821
rect 12491 1802 12866 1821
rect 12422 1799 12866 1802
rect 12698 1798 12866 1799
rect 11716 1771 11854 1780
rect 11510 1770 11547 1771
rect 11566 1719 11602 1771
rect 11621 1770 11658 1771
rect 11717 1770 11754 1771
rect 11037 1717 11078 1718
rect 10929 1710 11078 1717
rect 10929 1690 11047 1710
rect 11067 1690 11078 1710
rect 10929 1682 11078 1690
rect 11145 1714 11504 1718
rect 11145 1709 11467 1714
rect 11145 1685 11258 1709
rect 11282 1690 11467 1709
rect 11491 1690 11504 1714
rect 11282 1685 11504 1690
rect 11145 1682 11504 1685
rect 11566 1682 11601 1719
rect 11669 1716 11769 1719
rect 11669 1712 11736 1716
rect 11669 1686 11681 1712
rect 11707 1690 11736 1712
rect 11762 1690 11769 1716
rect 11707 1686 11769 1690
rect 11669 1682 11769 1686
rect 10356 1669 10394 1679
rect 9745 1665 9915 1666
rect 10356 1665 10366 1669
rect 8365 1660 8465 1664
rect 8365 1656 8427 1660
rect 8365 1630 8372 1656
rect 8398 1634 8427 1656
rect 8453 1634 8465 1660
rect 8398 1630 8465 1634
rect 8365 1627 8465 1630
rect 8533 1627 8568 1664
rect 8630 1661 8989 1664
rect 8630 1656 8852 1661
rect 8630 1632 8643 1656
rect 8667 1637 8852 1656
rect 8876 1637 8989 1661
rect 8667 1632 8989 1637
rect 8630 1628 8989 1632
rect 9056 1656 9205 1664
rect 9056 1636 9067 1656
rect 9087 1636 9205 1656
rect 9745 1651 10366 1665
rect 10384 1651 10394 1669
rect 11145 1661 11176 1682
rect 11566 1661 11602 1682
rect 9745 1645 10394 1651
rect 10809 1652 10846 1661
rect 10988 1660 11025 1661
rect 9745 1644 10393 1645
rect 10356 1642 10393 1644
rect 9056 1629 9205 1636
rect 10809 1634 10818 1652
rect 10836 1634 10846 1652
rect 9056 1628 9097 1629
rect 8380 1575 8417 1576
rect 8476 1575 8513 1576
rect 8532 1575 8568 1627
rect 8587 1575 8624 1576
rect 8280 1566 8418 1575
rect 8280 1546 8389 1566
rect 8409 1546 8418 1566
rect 8280 1539 8418 1546
rect 8476 1566 8624 1575
rect 8476 1546 8485 1566
rect 8505 1546 8595 1566
rect 8615 1546 8624 1566
rect 8280 1537 8376 1539
rect 8476 1536 8624 1546
rect 8683 1566 8720 1576
rect 8795 1575 8832 1576
rect 8776 1573 8832 1575
rect 8683 1546 8691 1566
rect 8711 1546 8720 1566
rect 8532 1535 8568 1536
rect 8380 1476 8417 1477
rect 8683 1476 8720 1546
rect 8745 1566 8832 1573
rect 8745 1563 8803 1566
rect 8745 1543 8750 1563
rect 8771 1546 8803 1563
rect 8823 1546 8832 1566
rect 8771 1543 8832 1546
rect 8745 1536 8832 1543
rect 8891 1566 8928 1576
rect 8891 1546 8899 1566
rect 8919 1546 8928 1566
rect 8745 1535 8776 1536
rect 8379 1475 8720 1476
rect 8304 1470 8720 1475
rect 8304 1450 8307 1470
rect 8327 1450 8720 1470
rect 8891 1475 8928 1546
rect 8958 1575 8989 1628
rect 10809 1624 10846 1634
rect 10810 1589 10846 1624
rect 10987 1651 11025 1660
rect 10987 1631 10996 1651
rect 11016 1631 11025 1651
rect 10987 1623 11025 1631
rect 11091 1655 11176 1661
rect 11201 1660 11238 1661
rect 11091 1635 11099 1655
rect 11119 1635 11176 1655
rect 11091 1627 11176 1635
rect 11200 1651 11238 1660
rect 11200 1631 11209 1651
rect 11229 1631 11238 1651
rect 11091 1626 11127 1627
rect 11200 1623 11238 1631
rect 11304 1655 11389 1661
rect 11409 1660 11446 1661
rect 11304 1635 11312 1655
rect 11332 1654 11389 1655
rect 11332 1635 11361 1654
rect 11304 1634 11361 1635
rect 11382 1634 11389 1654
rect 11304 1627 11389 1634
rect 11408 1651 11446 1660
rect 11408 1631 11417 1651
rect 11437 1631 11446 1651
rect 11304 1626 11340 1627
rect 11408 1623 11446 1631
rect 11512 1655 11656 1661
rect 11512 1635 11520 1655
rect 11540 1654 11628 1655
rect 11540 1635 11568 1654
rect 11512 1633 11568 1635
rect 11590 1635 11628 1654
rect 11648 1635 11656 1655
rect 11590 1633 11656 1635
rect 11512 1627 11656 1633
rect 11512 1626 11548 1627
rect 11620 1626 11656 1627
rect 11722 1660 11759 1661
rect 11722 1659 11760 1660
rect 11722 1651 11786 1659
rect 11722 1631 11731 1651
rect 11751 1637 11786 1651
rect 11806 1637 11809 1657
rect 11751 1632 11809 1637
rect 11751 1631 11786 1632
rect 10988 1594 11025 1623
rect 9008 1575 9045 1576
rect 8958 1566 9045 1575
rect 8958 1546 9016 1566
rect 9036 1546 9045 1566
rect 8958 1536 9045 1546
rect 9104 1566 9141 1576
rect 9104 1546 9112 1566
rect 9132 1546 9141 1566
rect 8958 1535 8989 1536
rect 9104 1475 9141 1546
rect 10359 1570 10396 1580
rect 10359 1552 10368 1570
rect 10386 1552 10396 1570
rect 10359 1543 10396 1552
rect 10808 1548 10846 1589
rect 10989 1592 11025 1594
rect 11201 1592 11238 1623
rect 10989 1570 11238 1592
rect 11409 1591 11446 1623
rect 11722 1619 11786 1631
rect 11826 1593 11853 1771
rect 11685 1591 11853 1593
rect 11409 1565 11853 1591
rect 11410 1548 11434 1565
rect 11685 1564 11853 1565
rect 10359 1519 10394 1543
rect 10357 1495 10394 1519
rect 10356 1489 10394 1495
rect 8891 1451 9141 1475
rect 9767 1471 10394 1489
rect 10808 1530 11435 1548
rect 12061 1544 12311 1568
rect 10808 1524 10846 1530
rect 10808 1500 10845 1524
rect 10808 1476 10843 1500
rect 9349 1454 9517 1455
rect 9768 1454 9792 1471
rect 9349 1428 9793 1454
rect 9349 1426 9517 1428
rect 9349 1248 9376 1426
rect 9416 1388 9480 1400
rect 9756 1396 9793 1428
rect 9964 1427 10213 1449
rect 9964 1396 10001 1427
rect 10177 1425 10213 1427
rect 10356 1430 10394 1471
rect 10806 1467 10843 1476
rect 10806 1449 10816 1467
rect 10834 1449 10843 1467
rect 10806 1439 10843 1449
rect 12061 1473 12098 1544
rect 12213 1483 12244 1484
rect 12061 1453 12070 1473
rect 12090 1453 12098 1473
rect 12061 1443 12098 1453
rect 12157 1473 12244 1483
rect 12157 1453 12166 1473
rect 12186 1453 12244 1473
rect 12157 1444 12244 1453
rect 12157 1443 12194 1444
rect 10177 1396 10214 1425
rect 9416 1387 9451 1388
rect 9393 1382 9451 1387
rect 9393 1362 9396 1382
rect 9416 1368 9451 1382
rect 9471 1368 9480 1388
rect 9416 1360 9480 1368
rect 9442 1359 9480 1360
rect 9443 1358 9480 1359
rect 9546 1392 9582 1393
rect 9654 1392 9690 1393
rect 9546 1386 9690 1392
rect 9546 1384 9612 1386
rect 9546 1364 9554 1384
rect 9574 1365 9612 1384
rect 9634 1384 9690 1386
rect 9634 1365 9662 1384
rect 9574 1364 9662 1365
rect 9682 1364 9690 1384
rect 9546 1358 9690 1364
rect 9756 1388 9794 1396
rect 9862 1392 9898 1393
rect 9756 1368 9765 1388
rect 9785 1368 9794 1388
rect 9756 1359 9794 1368
rect 9813 1385 9898 1392
rect 9813 1365 9820 1385
rect 9841 1384 9898 1385
rect 9841 1365 9870 1384
rect 9813 1364 9870 1365
rect 9890 1364 9898 1384
rect 9756 1358 9793 1359
rect 9813 1358 9898 1364
rect 9964 1388 10002 1396
rect 10075 1392 10111 1393
rect 9964 1368 9973 1388
rect 9993 1368 10002 1388
rect 9964 1359 10002 1368
rect 10026 1384 10111 1392
rect 10026 1364 10083 1384
rect 10103 1364 10111 1384
rect 9964 1358 10001 1359
rect 10026 1358 10111 1364
rect 10177 1388 10215 1396
rect 10177 1368 10186 1388
rect 10206 1368 10215 1388
rect 10177 1359 10215 1368
rect 10356 1395 10392 1430
rect 10356 1385 10393 1395
rect 12213 1391 12244 1444
rect 12274 1473 12311 1544
rect 12482 1549 12875 1569
rect 12895 1549 12898 1569
rect 12482 1544 12898 1549
rect 12482 1543 12823 1544
rect 12426 1483 12457 1484
rect 12274 1453 12283 1473
rect 12303 1453 12311 1473
rect 12274 1443 12311 1453
rect 12370 1476 12457 1483
rect 12370 1473 12431 1476
rect 12370 1453 12379 1473
rect 12399 1456 12431 1473
rect 12452 1456 12457 1476
rect 12399 1453 12457 1456
rect 12370 1446 12457 1453
rect 12482 1473 12519 1543
rect 12785 1542 12822 1543
rect 12634 1483 12670 1484
rect 12482 1453 12491 1473
rect 12511 1453 12519 1473
rect 12370 1444 12426 1446
rect 12370 1443 12407 1444
rect 12482 1443 12519 1453
rect 12578 1473 12726 1483
rect 12826 1480 12922 1482
rect 12578 1453 12587 1473
rect 12607 1453 12697 1473
rect 12717 1453 12726 1473
rect 12578 1444 12726 1453
rect 12784 1473 12922 1480
rect 12784 1453 12793 1473
rect 12813 1453 12922 1473
rect 12784 1444 12922 1453
rect 12578 1443 12615 1444
rect 12634 1392 12670 1444
rect 12689 1443 12726 1444
rect 12785 1443 12822 1444
rect 12105 1390 12146 1391
rect 10356 1367 10366 1385
rect 10384 1367 10393 1385
rect 11997 1383 12146 1390
rect 10809 1375 10846 1377
rect 10809 1374 11457 1375
rect 10177 1358 10214 1359
rect 10356 1358 10393 1367
rect 10808 1368 11457 1374
rect 9600 1337 9636 1358
rect 10026 1337 10057 1358
rect 10808 1350 10818 1368
rect 10836 1354 11457 1368
rect 11997 1363 12115 1383
rect 12135 1363 12146 1383
rect 11997 1355 12146 1363
rect 12213 1387 12572 1391
rect 12213 1382 12535 1387
rect 12213 1358 12326 1382
rect 12350 1363 12535 1382
rect 12559 1363 12572 1387
rect 12350 1358 12572 1363
rect 12213 1355 12572 1358
rect 12634 1355 12669 1392
rect 12737 1389 12837 1392
rect 12737 1385 12804 1389
rect 12737 1359 12749 1385
rect 12775 1363 12804 1385
rect 12830 1363 12837 1389
rect 12775 1359 12837 1363
rect 12737 1355 12837 1359
rect 10836 1350 10846 1354
rect 11287 1353 11457 1354
rect 10808 1340 10846 1350
rect 9433 1333 9533 1337
rect 9433 1329 9495 1333
rect 9433 1303 9440 1329
rect 9466 1307 9495 1329
rect 9521 1307 9533 1333
rect 9466 1303 9533 1307
rect 9433 1300 9533 1303
rect 9601 1300 9636 1337
rect 9698 1334 10057 1337
rect 9698 1329 9920 1334
rect 9698 1305 9711 1329
rect 9735 1310 9920 1329
rect 9944 1310 10057 1334
rect 9735 1305 10057 1310
rect 9698 1301 10057 1305
rect 10124 1329 10273 1337
rect 10124 1309 10135 1329
rect 10155 1309 10273 1329
rect 10124 1302 10273 1309
rect 10124 1301 10165 1302
rect 9448 1248 9485 1249
rect 9544 1248 9581 1249
rect 9600 1248 9636 1300
rect 9655 1248 9692 1249
rect 9348 1239 9486 1248
rect 7604 1230 7636 1235
rect 6384 1212 6480 1214
rect 6136 1185 6145 1205
rect 6165 1185 6255 1205
rect 6275 1185 6284 1205
rect 6136 1176 6284 1185
rect 6342 1205 6480 1212
rect 7097 1209 7543 1224
rect 7373 1208 7543 1209
rect 6342 1185 6351 1205
rect 6371 1185 6480 1205
rect 6342 1176 6480 1185
rect 6136 1175 6173 1176
rect 6192 1124 6228 1176
rect 6247 1175 6284 1176
rect 6343 1175 6380 1176
rect 5663 1122 5704 1123
rect 4489 1072 5121 1079
rect 4489 1070 4551 1072
rect 4067 1060 4235 1061
rect 4489 1060 4511 1070
rect 3782 1035 3819 1036
rect 3732 1026 3819 1035
rect 3732 1006 3790 1026
rect 3810 1006 3819 1026
rect 3732 996 3819 1006
rect 3878 1026 3915 1036
rect 3878 1006 3886 1026
rect 3906 1006 3915 1026
rect 3732 995 3763 996
rect 3878 935 3915 1006
rect 3665 911 3915 935
rect 4067 1034 4511 1060
rect 4067 1032 4235 1034
rect 4067 854 4094 1032
rect 4134 994 4198 1006
rect 4474 1002 4511 1034
rect 4682 1033 4931 1055
rect 4682 1002 4719 1033
rect 4895 1031 4931 1033
rect 4895 1002 4932 1031
rect 4134 993 4169 994
rect 4111 988 4169 993
rect 4111 968 4114 988
rect 4134 974 4169 988
rect 4189 974 4198 994
rect 4134 966 4198 974
rect 4160 965 4198 966
rect 4161 964 4198 965
rect 4264 998 4300 999
rect 4372 998 4408 999
rect 4264 990 4408 998
rect 4264 970 4272 990
rect 4292 970 4321 990
rect 4264 969 4321 970
rect 4343 970 4380 990
rect 4400 970 4408 990
rect 4343 969 4408 970
rect 4264 964 4408 969
rect 4474 994 4512 1002
rect 4580 998 4616 999
rect 4474 974 4483 994
rect 4503 974 4512 994
rect 4474 965 4512 974
rect 4531 991 4616 998
rect 4531 971 4538 991
rect 4559 990 4616 991
rect 4559 971 4588 990
rect 4531 970 4588 971
rect 4608 970 4616 990
rect 4474 964 4511 965
rect 4531 964 4616 970
rect 4682 994 4720 1002
rect 4793 998 4829 999
rect 4682 974 4691 994
rect 4711 974 4720 994
rect 4682 965 4720 974
rect 4744 990 4829 998
rect 4744 970 4801 990
rect 4821 970 4829 990
rect 4682 964 4719 965
rect 4744 964 4829 970
rect 4895 994 4933 1002
rect 4895 974 4904 994
rect 4924 974 4933 994
rect 4895 965 4933 974
rect 4895 964 4932 965
rect 4318 943 4354 964
rect 4744 943 4775 964
rect 4151 939 4251 943
rect 4151 935 4213 939
rect 4151 909 4158 935
rect 4184 913 4213 935
rect 4239 913 4251 939
rect 4184 909 4251 913
rect 4151 906 4251 909
rect 4319 906 4354 943
rect 4416 940 4775 943
rect 4416 935 4638 940
rect 4416 911 4429 935
rect 4453 916 4638 935
rect 4662 916 4775 940
rect 4453 911 4775 916
rect 4416 907 4775 911
rect 4842 935 4991 943
rect 4842 915 4853 935
rect 4873 915 4991 935
rect 4842 908 4991 915
rect 5082 923 5121 1072
rect 5425 958 5464 1107
rect 5555 1115 5704 1122
rect 5555 1095 5673 1115
rect 5693 1095 5704 1115
rect 5555 1087 5704 1095
rect 5771 1119 6130 1123
rect 5771 1114 6093 1119
rect 5771 1090 5884 1114
rect 5908 1095 6093 1114
rect 6117 1095 6130 1119
rect 5908 1090 6130 1095
rect 5771 1087 6130 1090
rect 6192 1087 6227 1124
rect 6295 1121 6395 1124
rect 6295 1117 6362 1121
rect 6295 1091 6307 1117
rect 6333 1095 6362 1117
rect 6388 1095 6395 1121
rect 6333 1091 6395 1095
rect 6295 1087 6395 1091
rect 5771 1066 5802 1087
rect 6192 1066 6228 1087
rect 5614 1065 5651 1066
rect 5613 1056 5651 1065
rect 5613 1036 5622 1056
rect 5642 1036 5651 1056
rect 5613 1028 5651 1036
rect 5717 1060 5802 1066
rect 5827 1065 5864 1066
rect 5717 1040 5725 1060
rect 5745 1040 5802 1060
rect 5717 1032 5802 1040
rect 5826 1056 5864 1065
rect 5826 1036 5835 1056
rect 5855 1036 5864 1056
rect 5717 1031 5753 1032
rect 5826 1028 5864 1036
rect 5930 1060 6015 1066
rect 6035 1065 6072 1066
rect 5930 1040 5938 1060
rect 5958 1059 6015 1060
rect 5958 1040 5987 1059
rect 5930 1039 5987 1040
rect 6008 1039 6015 1059
rect 5930 1032 6015 1039
rect 6034 1056 6072 1065
rect 6034 1036 6043 1056
rect 6063 1036 6072 1056
rect 5930 1031 5966 1032
rect 6034 1028 6072 1036
rect 6138 1061 6282 1066
rect 6138 1060 6203 1061
rect 6138 1040 6146 1060
rect 6166 1040 6203 1060
rect 6225 1060 6282 1061
rect 6225 1040 6254 1060
rect 6274 1040 6282 1060
rect 6138 1032 6282 1040
rect 6138 1031 6174 1032
rect 6246 1031 6282 1032
rect 6348 1065 6385 1066
rect 6348 1064 6386 1065
rect 6348 1056 6412 1064
rect 6348 1036 6357 1056
rect 6377 1042 6412 1056
rect 6432 1042 6435 1062
rect 6377 1037 6435 1042
rect 6377 1036 6412 1037
rect 5614 999 5651 1028
rect 5615 997 5651 999
rect 5827 997 5864 1028
rect 5615 975 5864 997
rect 6035 996 6072 1028
rect 6348 1024 6412 1036
rect 6452 998 6479 1176
rect 6311 996 6479 998
rect 6035 970 6479 996
rect 6631 1095 6881 1119
rect 6631 1024 6668 1095
rect 6783 1034 6814 1035
rect 6631 1004 6640 1024
rect 6660 1004 6668 1024
rect 6631 994 6668 1004
rect 6727 1024 6814 1034
rect 6727 1004 6736 1024
rect 6756 1004 6814 1024
rect 6727 995 6814 1004
rect 6727 994 6764 995
rect 6035 960 6057 970
rect 6311 969 6479 970
rect 5995 958 6057 960
rect 5425 951 6057 958
rect 4842 907 4883 908
rect 4166 854 4203 855
rect 4262 854 4299 855
rect 4318 854 4354 906
rect 4373 854 4410 855
rect 2231 809 2236 835
rect 2255 809 2262 835
rect 4066 845 4204 854
rect 4066 825 4175 845
rect 4195 825 4204 845
rect 4066 818 4204 825
rect 4262 845 4410 854
rect 4262 825 4271 845
rect 4291 825 4381 845
rect 4401 825 4410 845
rect 4066 816 4162 818
rect 4262 815 4410 825
rect 4469 845 4506 855
rect 4581 854 4618 855
rect 4562 852 4618 854
rect 4469 825 4477 845
rect 4497 825 4506 845
rect 4318 814 4354 815
rect 2231 806 2262 809
rect 1060 782 1198 791
rect 854 781 891 782
rect 910 730 946 782
rect 965 781 1002 782
rect 1061 781 1098 782
rect 381 728 422 729
rect 273 721 422 728
rect 273 701 391 721
rect 411 701 422 721
rect 273 693 422 701
rect 489 725 848 729
rect 489 720 811 725
rect 489 696 602 720
rect 626 701 811 720
rect 835 701 848 725
rect 626 696 848 701
rect 489 693 848 696
rect 910 693 945 730
rect 1013 727 1113 730
rect 1013 723 1080 727
rect 1013 697 1025 723
rect 1051 701 1080 723
rect 1106 701 1113 727
rect 1051 697 1113 701
rect 1013 693 1113 697
rect 489 672 520 693
rect 910 672 946 693
rect 153 663 190 672
rect 332 671 369 672
rect 153 645 162 663
rect 180 645 190 663
rect 153 635 190 645
rect 154 600 190 635
rect 331 662 369 671
rect 331 642 340 662
rect 360 642 369 662
rect 331 634 369 642
rect 435 666 520 672
rect 545 671 582 672
rect 435 646 443 666
rect 463 646 520 666
rect 435 638 520 646
rect 544 662 582 671
rect 544 642 553 662
rect 573 642 582 662
rect 435 637 471 638
rect 544 634 582 642
rect 648 666 733 672
rect 753 671 790 672
rect 648 646 656 666
rect 676 665 733 666
rect 676 646 705 665
rect 648 645 705 646
rect 726 645 733 665
rect 648 638 733 645
rect 752 662 790 671
rect 752 642 761 662
rect 781 642 790 662
rect 648 637 684 638
rect 752 634 790 642
rect 856 666 1000 672
rect 856 646 864 666
rect 884 665 972 666
rect 884 646 912 665
rect 856 644 912 646
rect 934 646 972 665
rect 992 646 1000 666
rect 934 644 1000 646
rect 856 638 1000 644
rect 856 637 892 638
rect 964 637 1000 638
rect 1066 671 1103 672
rect 1066 670 1104 671
rect 1066 662 1130 670
rect 1066 642 1075 662
rect 1095 648 1130 662
rect 1150 648 1153 668
rect 1095 643 1153 648
rect 1095 642 1130 643
rect 332 605 369 634
rect 152 535 190 600
rect 333 603 369 605
rect 545 603 582 634
rect 333 581 582 603
rect 753 602 790 634
rect 1066 630 1130 642
rect 1170 604 1197 782
rect 4166 755 4203 756
rect 4469 755 4506 825
rect 4531 845 4618 852
rect 4531 842 4589 845
rect 4531 822 4536 842
rect 4557 825 4589 842
rect 4609 825 4618 845
rect 4557 822 4618 825
rect 4531 815 4618 822
rect 4677 845 4714 855
rect 4677 825 4685 845
rect 4705 825 4714 845
rect 4531 814 4562 815
rect 4165 754 4506 755
rect 4090 749 4506 754
rect 4090 729 4093 749
rect 4113 729 4506 749
rect 4677 754 4714 825
rect 4744 854 4775 907
rect 5082 905 5092 923
rect 5110 905 5121 923
rect 5424 942 6057 951
rect 6783 942 6814 995
rect 6844 1024 6881 1095
rect 7052 1100 7445 1120
rect 7465 1100 7468 1120
rect 7052 1095 7468 1100
rect 7052 1094 7393 1095
rect 6996 1034 7027 1035
rect 6844 1004 6853 1024
rect 6873 1004 6881 1024
rect 6844 994 6881 1004
rect 6940 1027 7027 1034
rect 6940 1024 7001 1027
rect 6940 1004 6949 1024
rect 6969 1007 7001 1024
rect 7022 1007 7027 1027
rect 6969 1004 7027 1007
rect 6940 997 7027 1004
rect 7052 1024 7089 1094
rect 7355 1093 7392 1094
rect 7204 1034 7240 1035
rect 7052 1004 7061 1024
rect 7081 1004 7089 1024
rect 6940 995 6996 997
rect 6940 994 6977 995
rect 7052 994 7089 1004
rect 7148 1024 7296 1034
rect 7396 1031 7492 1033
rect 7148 1004 7157 1024
rect 7177 1004 7267 1024
rect 7287 1004 7296 1024
rect 7148 995 7296 1004
rect 7354 1024 7492 1031
rect 7354 1004 7363 1024
rect 7383 1004 7492 1024
rect 7354 995 7492 1004
rect 7148 994 7185 995
rect 7204 943 7240 995
rect 7259 994 7296 995
rect 7355 994 7392 995
rect 5424 924 5434 942
rect 5452 941 6057 942
rect 6675 941 6716 942
rect 5452 936 5473 941
rect 5452 924 5464 936
rect 6567 934 6716 941
rect 5424 916 5464 924
rect 5507 923 5533 924
rect 5424 914 5461 916
rect 5507 905 6061 923
rect 6567 914 6685 934
rect 6705 914 6716 934
rect 6567 906 6716 914
rect 6783 938 7142 942
rect 6783 933 7105 938
rect 6783 909 6896 933
rect 6920 914 7105 933
rect 7129 914 7142 938
rect 6920 909 7142 914
rect 6783 906 7142 909
rect 7204 906 7239 943
rect 7307 940 7407 943
rect 7307 936 7374 940
rect 7307 910 7319 936
rect 7345 914 7374 936
rect 7400 914 7407 940
rect 7345 910 7407 914
rect 7307 906 7407 910
rect 5082 896 5119 905
rect 4794 854 4831 855
rect 4744 845 4831 854
rect 4744 825 4802 845
rect 4822 825 4831 845
rect 4744 815 4831 825
rect 4890 845 4927 855
rect 4890 825 4898 845
rect 4918 825 4927 845
rect 5427 846 5464 852
rect 5507 846 5533 905
rect 6040 886 6061 905
rect 5427 843 5533 846
rect 5085 830 5122 834
rect 4744 814 4775 815
rect 4890 754 4927 825
rect 4677 730 4927 754
rect 5083 824 5122 830
rect 5083 806 5094 824
rect 5112 806 5122 824
rect 5427 825 5436 843
rect 5454 829 5533 843
rect 5618 861 5868 885
rect 5454 827 5530 829
rect 5454 825 5464 827
rect 5427 815 5464 825
rect 5083 797 5122 806
rect 4469 706 4506 729
rect 5083 719 5118 797
rect 5432 750 5463 815
rect 5618 790 5655 861
rect 5770 800 5801 801
rect 5618 770 5627 790
rect 5647 770 5655 790
rect 5618 760 5655 770
rect 5714 790 5801 800
rect 5714 770 5723 790
rect 5743 770 5801 790
rect 5714 761 5801 770
rect 5714 760 5751 761
rect 5080 709 5118 719
rect 5431 741 5468 750
rect 5431 723 5441 741
rect 5459 723 5468 741
rect 5431 713 5468 723
rect 4469 705 4639 706
rect 5080 705 5090 709
rect 4469 691 5090 705
rect 5108 691 5118 709
rect 5770 708 5801 761
rect 5831 790 5868 861
rect 6039 866 6432 886
rect 6452 866 6455 886
rect 6783 885 6814 906
rect 7204 885 7240 906
rect 6626 884 6663 885
rect 6039 861 6455 866
rect 6625 875 6663 884
rect 6039 860 6380 861
rect 5983 800 6014 801
rect 5831 770 5840 790
rect 5860 770 5868 790
rect 5831 760 5868 770
rect 5927 793 6014 800
rect 5927 790 5988 793
rect 5927 770 5936 790
rect 5956 773 5988 790
rect 6009 773 6014 793
rect 5956 770 6014 773
rect 5927 763 6014 770
rect 6039 790 6076 860
rect 6342 859 6379 860
rect 6625 855 6634 875
rect 6654 855 6663 875
rect 6625 847 6663 855
rect 6729 879 6814 885
rect 6839 884 6876 885
rect 6729 859 6737 879
rect 6757 859 6814 879
rect 6729 851 6814 859
rect 6838 875 6876 884
rect 6838 855 6847 875
rect 6867 855 6876 875
rect 6729 850 6765 851
rect 6838 847 6876 855
rect 6942 879 7027 885
rect 7047 884 7084 885
rect 6942 859 6950 879
rect 6970 878 7027 879
rect 6970 859 6999 878
rect 6942 858 6999 859
rect 7020 858 7027 878
rect 6942 851 7027 858
rect 7046 875 7084 884
rect 7046 855 7055 875
rect 7075 855 7084 875
rect 6942 850 6978 851
rect 7046 847 7084 855
rect 7150 880 7294 885
rect 7150 879 7209 880
rect 7150 859 7158 879
rect 7178 860 7209 879
rect 7233 879 7294 880
rect 7233 860 7266 879
rect 7178 859 7266 860
rect 7286 859 7294 879
rect 7150 851 7294 859
rect 7150 850 7186 851
rect 7258 850 7294 851
rect 7360 884 7397 885
rect 7360 883 7398 884
rect 7360 875 7424 883
rect 7360 855 7369 875
rect 7389 861 7424 875
rect 7444 861 7447 881
rect 7389 856 7447 861
rect 7389 855 7424 856
rect 6626 818 6663 847
rect 6627 816 6663 818
rect 6839 816 6876 847
rect 6191 800 6227 801
rect 6039 770 6048 790
rect 6068 770 6076 790
rect 5927 761 5983 763
rect 5927 760 5964 761
rect 6039 760 6076 770
rect 6135 790 6283 800
rect 6383 797 6479 799
rect 6135 770 6144 790
rect 6164 770 6254 790
rect 6274 770 6283 790
rect 6135 761 6283 770
rect 6341 790 6479 797
rect 6627 794 6876 816
rect 7047 815 7084 847
rect 7360 843 7424 855
rect 7464 817 7491 995
rect 7323 815 7491 817
rect 7047 811 7491 815
rect 6341 770 6350 790
rect 6370 770 6479 790
rect 7047 792 7096 811
rect 7116 792 7491 811
rect 7047 789 7491 792
rect 7323 788 7491 789
rect 7512 814 7543 1208
rect 7604 1212 7609 1230
rect 7629 1212 7636 1230
rect 7604 1207 7636 1212
rect 7607 1205 7636 1207
rect 8336 1220 8504 1221
rect 8336 1217 8780 1220
rect 8336 1198 8711 1217
rect 8731 1198 8780 1217
rect 9348 1219 9457 1239
rect 9477 1219 9486 1239
rect 8336 1194 8780 1198
rect 8336 1192 8504 1194
rect 8336 1014 8363 1192
rect 8403 1154 8467 1166
rect 8743 1162 8780 1194
rect 8951 1193 9200 1215
rect 9348 1212 9486 1219
rect 9544 1239 9692 1248
rect 9544 1219 9553 1239
rect 9573 1219 9663 1239
rect 9683 1219 9692 1239
rect 9348 1210 9444 1212
rect 9544 1209 9692 1219
rect 9751 1239 9788 1249
rect 9863 1248 9900 1249
rect 9844 1246 9900 1248
rect 9751 1219 9759 1239
rect 9779 1219 9788 1239
rect 9600 1208 9636 1209
rect 8951 1162 8988 1193
rect 9164 1191 9200 1193
rect 9164 1162 9201 1191
rect 8403 1153 8438 1154
rect 8380 1148 8438 1153
rect 8380 1128 8383 1148
rect 8403 1134 8438 1148
rect 8458 1134 8467 1154
rect 8403 1126 8467 1134
rect 8429 1125 8467 1126
rect 8430 1124 8467 1125
rect 8533 1158 8569 1159
rect 8641 1158 8677 1159
rect 8533 1150 8677 1158
rect 8533 1130 8541 1150
rect 8561 1130 8593 1150
rect 8617 1130 8649 1150
rect 8669 1130 8677 1150
rect 8533 1124 8677 1130
rect 8743 1154 8781 1162
rect 8849 1158 8885 1159
rect 8743 1134 8752 1154
rect 8772 1134 8781 1154
rect 8743 1125 8781 1134
rect 8800 1151 8885 1158
rect 8800 1131 8807 1151
rect 8828 1150 8885 1151
rect 8828 1131 8857 1150
rect 8800 1130 8857 1131
rect 8877 1130 8885 1150
rect 8743 1124 8780 1125
rect 8800 1124 8885 1130
rect 8951 1154 8989 1162
rect 9062 1158 9098 1159
rect 8951 1134 8960 1154
rect 8980 1134 8989 1154
rect 8951 1125 8989 1134
rect 9013 1150 9098 1158
rect 9013 1130 9070 1150
rect 9090 1130 9098 1150
rect 8951 1124 8988 1125
rect 9013 1124 9098 1130
rect 9164 1154 9202 1162
rect 9164 1134 9173 1154
rect 9193 1134 9202 1154
rect 9448 1149 9485 1150
rect 9751 1149 9788 1219
rect 9813 1239 9900 1246
rect 9813 1236 9871 1239
rect 9813 1216 9818 1236
rect 9839 1219 9871 1236
rect 9891 1219 9900 1239
rect 9839 1216 9900 1219
rect 9813 1209 9900 1216
rect 9959 1239 9996 1249
rect 9959 1219 9967 1239
rect 9987 1219 9996 1239
rect 9813 1208 9844 1209
rect 9447 1148 9788 1149
rect 9164 1125 9202 1134
rect 9372 1143 9788 1148
rect 9164 1124 9201 1125
rect 8587 1103 8623 1124
rect 9013 1103 9044 1124
rect 9372 1123 9375 1143
rect 9395 1123 9788 1143
rect 9959 1148 9996 1219
rect 10026 1248 10057 1301
rect 10359 1286 10396 1296
rect 10359 1268 10368 1286
rect 10386 1268 10396 1286
rect 10359 1259 10396 1268
rect 10808 1262 10843 1340
rect 11420 1330 11457 1353
rect 12213 1334 12244 1355
rect 12634 1334 12670 1355
rect 12056 1333 12093 1334
rect 10076 1248 10113 1249
rect 10026 1239 10113 1248
rect 10026 1219 10084 1239
rect 10104 1219 10113 1239
rect 10026 1209 10113 1219
rect 10172 1239 10209 1249
rect 10172 1219 10180 1239
rect 10200 1219 10209 1239
rect 10026 1208 10057 1209
rect 10172 1148 10209 1219
rect 10364 1194 10395 1259
rect 10804 1253 10843 1262
rect 10804 1235 10814 1253
rect 10832 1235 10843 1253
rect 10804 1229 10843 1235
rect 10999 1305 11249 1329
rect 10999 1234 11036 1305
rect 11151 1244 11182 1245
rect 10804 1225 10841 1229
rect 10999 1214 11008 1234
rect 11028 1214 11036 1234
rect 10999 1204 11036 1214
rect 11095 1234 11182 1244
rect 11095 1214 11104 1234
rect 11124 1214 11182 1234
rect 11095 1205 11182 1214
rect 11095 1204 11132 1205
rect 10363 1184 10400 1194
rect 10363 1182 10373 1184
rect 10297 1180 10373 1182
rect 9959 1124 10209 1148
rect 10294 1166 10373 1180
rect 10391 1166 10400 1184
rect 10294 1163 10400 1166
rect 9766 1104 9787 1123
rect 10294 1104 10320 1163
rect 10363 1157 10400 1163
rect 10807 1154 10844 1163
rect 8420 1099 8520 1103
rect 8420 1095 8482 1099
rect 8420 1069 8427 1095
rect 8453 1073 8482 1095
rect 8508 1073 8520 1099
rect 8453 1069 8520 1073
rect 8420 1066 8520 1069
rect 8588 1066 8623 1103
rect 8685 1100 9044 1103
rect 8685 1095 8907 1100
rect 8685 1071 8698 1095
rect 8722 1076 8907 1095
rect 8931 1076 9044 1100
rect 8722 1071 9044 1076
rect 8685 1067 9044 1071
rect 9111 1095 9260 1103
rect 9111 1075 9122 1095
rect 9142 1075 9260 1095
rect 9766 1086 10320 1104
rect 10805 1136 10816 1154
rect 10834 1136 10844 1154
rect 11151 1152 11182 1205
rect 11212 1234 11249 1305
rect 11420 1310 11813 1330
rect 11833 1310 11836 1330
rect 11420 1305 11836 1310
rect 12055 1324 12093 1333
rect 11420 1304 11761 1305
rect 12055 1304 12064 1324
rect 12084 1304 12093 1324
rect 11364 1244 11395 1245
rect 11212 1214 11221 1234
rect 11241 1214 11249 1234
rect 11212 1204 11249 1214
rect 11308 1237 11395 1244
rect 11308 1234 11369 1237
rect 11308 1214 11317 1234
rect 11337 1217 11369 1234
rect 11390 1217 11395 1237
rect 11337 1214 11395 1217
rect 11308 1207 11395 1214
rect 11420 1234 11457 1304
rect 11723 1303 11760 1304
rect 12055 1296 12093 1304
rect 12159 1328 12244 1334
rect 12269 1333 12306 1334
rect 12159 1308 12167 1328
rect 12187 1308 12244 1328
rect 12159 1300 12244 1308
rect 12268 1324 12306 1333
rect 12268 1304 12277 1324
rect 12297 1304 12306 1324
rect 12159 1299 12195 1300
rect 12268 1296 12306 1304
rect 12372 1328 12457 1334
rect 12477 1333 12514 1334
rect 12372 1308 12380 1328
rect 12400 1327 12457 1328
rect 12400 1308 12429 1327
rect 12372 1307 12429 1308
rect 12450 1307 12457 1327
rect 12372 1300 12457 1307
rect 12476 1324 12514 1333
rect 12476 1304 12485 1324
rect 12505 1304 12514 1324
rect 12372 1299 12408 1300
rect 12476 1296 12514 1304
rect 12580 1328 12724 1334
rect 12580 1308 12588 1328
rect 12608 1327 12696 1328
rect 12608 1308 12641 1327
rect 12664 1308 12696 1327
rect 12716 1308 12724 1328
rect 12580 1300 12724 1308
rect 12580 1299 12616 1300
rect 12688 1299 12724 1300
rect 12790 1333 12827 1334
rect 12790 1332 12828 1333
rect 12790 1324 12854 1332
rect 12790 1304 12799 1324
rect 12819 1310 12854 1324
rect 12874 1310 12877 1330
rect 12819 1305 12877 1310
rect 12819 1304 12854 1305
rect 12056 1267 12093 1296
rect 12057 1265 12093 1267
rect 12269 1265 12306 1296
rect 11572 1244 11608 1245
rect 11420 1214 11429 1234
rect 11449 1214 11457 1234
rect 11308 1205 11364 1207
rect 11308 1204 11345 1205
rect 11420 1204 11457 1214
rect 11516 1234 11664 1244
rect 12057 1243 12306 1265
rect 12477 1264 12514 1296
rect 12790 1292 12854 1304
rect 12894 1266 12921 1444
rect 12753 1264 12921 1266
rect 12477 1253 12921 1264
rect 12984 1264 13014 2265
rect 13103 2258 13140 2269
rect 14724 2258 14751 2436
rect 14791 2398 14855 2410
rect 15131 2406 15168 2438
rect 15339 2437 15588 2459
rect 15339 2406 15376 2437
rect 15552 2435 15588 2437
rect 15731 2440 15769 2481
rect 15552 2406 15589 2435
rect 14791 2397 14826 2398
rect 14768 2392 14826 2397
rect 14768 2372 14771 2392
rect 14791 2378 14826 2392
rect 14846 2378 14855 2398
rect 14791 2370 14855 2378
rect 14817 2369 14855 2370
rect 14818 2368 14855 2369
rect 14921 2402 14957 2403
rect 15029 2402 15065 2403
rect 14921 2396 15065 2402
rect 14921 2394 14987 2396
rect 14921 2374 14929 2394
rect 14949 2375 14987 2394
rect 15009 2394 15065 2396
rect 15009 2375 15037 2394
rect 14949 2374 15037 2375
rect 15057 2374 15065 2394
rect 14921 2368 15065 2374
rect 15131 2398 15169 2406
rect 15237 2402 15273 2403
rect 15131 2378 15140 2398
rect 15160 2378 15169 2398
rect 15131 2369 15169 2378
rect 15188 2395 15273 2402
rect 15188 2375 15195 2395
rect 15216 2394 15273 2395
rect 15216 2375 15245 2394
rect 15188 2374 15245 2375
rect 15265 2374 15273 2394
rect 15131 2368 15168 2369
rect 15188 2368 15273 2374
rect 15339 2398 15377 2406
rect 15450 2402 15486 2403
rect 15339 2378 15348 2398
rect 15368 2378 15377 2398
rect 15339 2369 15377 2378
rect 15401 2394 15486 2402
rect 15401 2374 15458 2394
rect 15478 2374 15486 2394
rect 15339 2368 15376 2369
rect 15401 2368 15486 2374
rect 15552 2398 15590 2406
rect 15552 2378 15561 2398
rect 15581 2378 15590 2398
rect 15552 2369 15590 2378
rect 15731 2405 15767 2440
rect 16084 2436 16119 2482
rect 17495 2480 17532 2551
rect 17647 2490 17678 2491
rect 17495 2460 17504 2480
rect 17524 2460 17532 2480
rect 17495 2450 17532 2460
rect 17591 2480 17678 2490
rect 17591 2460 17600 2480
rect 17620 2460 17678 2480
rect 17591 2451 17678 2460
rect 17591 2450 17628 2451
rect 16082 2427 16119 2436
rect 16082 2409 16092 2427
rect 16110 2409 16119 2427
rect 15731 2395 15768 2405
rect 16082 2399 16119 2409
rect 17647 2398 17678 2451
rect 17708 2480 17745 2551
rect 17916 2556 18309 2576
rect 18329 2556 18332 2576
rect 17916 2551 18332 2556
rect 17916 2550 18257 2551
rect 17860 2490 17891 2491
rect 17708 2460 17717 2480
rect 17737 2460 17745 2480
rect 17708 2450 17745 2460
rect 17804 2483 17891 2490
rect 17804 2480 17865 2483
rect 17804 2460 17813 2480
rect 17833 2463 17865 2480
rect 17886 2463 17891 2483
rect 17833 2460 17891 2463
rect 17804 2453 17891 2460
rect 17916 2480 17953 2550
rect 18219 2549 18256 2550
rect 18068 2490 18104 2491
rect 17916 2460 17925 2480
rect 17945 2460 17953 2480
rect 17804 2451 17860 2453
rect 17804 2450 17841 2451
rect 17916 2450 17953 2460
rect 18012 2480 18160 2490
rect 18260 2487 18356 2489
rect 18012 2460 18021 2480
rect 18041 2460 18131 2480
rect 18151 2460 18160 2480
rect 18012 2451 18160 2460
rect 18218 2480 18356 2487
rect 18218 2460 18227 2480
rect 18247 2460 18356 2480
rect 18218 2451 18356 2460
rect 18012 2450 18049 2451
rect 18068 2399 18104 2451
rect 18123 2450 18160 2451
rect 18219 2450 18256 2451
rect 17539 2397 17580 2398
rect 15731 2377 15741 2395
rect 15759 2377 15768 2395
rect 15552 2368 15589 2369
rect 15731 2368 15768 2377
rect 17431 2390 17580 2397
rect 17431 2370 17549 2390
rect 17569 2370 17580 2390
rect 14975 2347 15011 2368
rect 15401 2347 15432 2368
rect 17431 2362 17580 2370
rect 17647 2394 18006 2398
rect 17647 2389 17969 2394
rect 17647 2365 17760 2389
rect 17784 2370 17969 2389
rect 17993 2370 18006 2394
rect 17784 2365 18006 2370
rect 17647 2362 18006 2365
rect 18068 2362 18103 2399
rect 18171 2396 18271 2399
rect 18171 2392 18238 2396
rect 18171 2366 18183 2392
rect 18209 2370 18238 2392
rect 18264 2370 18271 2396
rect 18209 2366 18271 2370
rect 18171 2362 18271 2366
rect 14808 2343 14908 2347
rect 14808 2339 14870 2343
rect 14808 2313 14815 2339
rect 14841 2317 14870 2339
rect 14896 2317 14908 2343
rect 14841 2313 14908 2317
rect 14808 2310 14908 2313
rect 14976 2310 15011 2347
rect 15073 2344 15432 2347
rect 15073 2339 15295 2344
rect 15073 2315 15086 2339
rect 15110 2320 15295 2339
rect 15319 2320 15432 2344
rect 15110 2315 15432 2320
rect 15073 2311 15432 2315
rect 15499 2339 15648 2347
rect 17647 2341 17678 2362
rect 18068 2341 18104 2362
rect 17490 2340 17527 2341
rect 15499 2319 15510 2339
rect 15530 2319 15648 2339
rect 16085 2335 16122 2337
rect 16085 2334 16733 2335
rect 15499 2312 15648 2319
rect 16084 2328 16733 2334
rect 15499 2311 15540 2312
rect 14823 2258 14860 2259
rect 14919 2258 14956 2259
rect 14975 2258 15011 2310
rect 15030 2258 15067 2259
rect 14723 2249 14861 2258
rect 13659 2231 13690 2234
rect 13659 2205 13666 2231
rect 13685 2205 13690 2231
rect 13659 1811 13690 2205
rect 13711 2230 13879 2231
rect 13711 2227 14155 2230
rect 13711 2208 14086 2227
rect 14106 2208 14155 2227
rect 14723 2229 14832 2249
rect 14852 2229 14861 2249
rect 13711 2204 14155 2208
rect 13711 2202 13879 2204
rect 13711 2024 13738 2202
rect 13778 2164 13842 2176
rect 14118 2172 14155 2204
rect 14326 2203 14575 2225
rect 14723 2222 14861 2229
rect 14919 2249 15067 2258
rect 14919 2229 14928 2249
rect 14948 2229 15038 2249
rect 15058 2229 15067 2249
rect 14723 2220 14819 2222
rect 14919 2219 15067 2229
rect 15126 2249 15163 2259
rect 15238 2258 15275 2259
rect 15219 2256 15275 2258
rect 15126 2229 15134 2249
rect 15154 2229 15163 2249
rect 14975 2218 15011 2219
rect 14326 2172 14363 2203
rect 14539 2201 14575 2203
rect 14539 2172 14576 2201
rect 13778 2163 13813 2164
rect 13755 2158 13813 2163
rect 13755 2138 13758 2158
rect 13778 2144 13813 2158
rect 13833 2144 13842 2164
rect 13778 2136 13842 2144
rect 13804 2135 13842 2136
rect 13805 2134 13842 2135
rect 13908 2168 13944 2169
rect 14016 2168 14052 2169
rect 13908 2160 14052 2168
rect 13908 2140 13916 2160
rect 13936 2159 14024 2160
rect 13936 2140 13969 2159
rect 13908 2139 13969 2140
rect 13993 2140 14024 2159
rect 14044 2140 14052 2160
rect 13993 2139 14052 2140
rect 13908 2134 14052 2139
rect 14118 2164 14156 2172
rect 14224 2168 14260 2169
rect 14118 2144 14127 2164
rect 14147 2144 14156 2164
rect 14118 2135 14156 2144
rect 14175 2161 14260 2168
rect 14175 2141 14182 2161
rect 14203 2160 14260 2161
rect 14203 2141 14232 2160
rect 14175 2140 14232 2141
rect 14252 2140 14260 2160
rect 14118 2134 14155 2135
rect 14175 2134 14260 2140
rect 14326 2164 14364 2172
rect 14437 2168 14473 2169
rect 14326 2144 14335 2164
rect 14355 2144 14364 2164
rect 14326 2135 14364 2144
rect 14388 2160 14473 2168
rect 14388 2140 14445 2160
rect 14465 2140 14473 2160
rect 14326 2134 14363 2135
rect 14388 2134 14473 2140
rect 14539 2164 14577 2172
rect 14539 2144 14548 2164
rect 14568 2144 14577 2164
rect 14823 2159 14860 2160
rect 15126 2159 15163 2229
rect 15188 2249 15275 2256
rect 15188 2246 15246 2249
rect 15188 2226 15193 2246
rect 15214 2229 15246 2246
rect 15266 2229 15275 2249
rect 15214 2226 15275 2229
rect 15188 2219 15275 2226
rect 15334 2249 15371 2259
rect 15334 2229 15342 2249
rect 15362 2229 15371 2249
rect 15188 2218 15219 2219
rect 14822 2158 15163 2159
rect 14539 2135 14577 2144
rect 14747 2153 15163 2158
rect 14539 2134 14576 2135
rect 13962 2113 13998 2134
rect 14388 2113 14419 2134
rect 14747 2133 14750 2153
rect 14770 2133 15163 2153
rect 15334 2158 15371 2229
rect 15401 2258 15432 2311
rect 16084 2310 16094 2328
rect 16112 2314 16733 2328
rect 16112 2310 16122 2314
rect 16563 2313 16733 2314
rect 15734 2296 15771 2306
rect 15734 2278 15743 2296
rect 15761 2278 15771 2296
rect 15734 2269 15771 2278
rect 16084 2300 16122 2310
rect 15451 2258 15488 2259
rect 15401 2249 15488 2258
rect 15401 2229 15459 2249
rect 15479 2229 15488 2249
rect 15401 2219 15488 2229
rect 15547 2249 15584 2259
rect 15547 2229 15555 2249
rect 15575 2229 15584 2249
rect 15401 2218 15432 2219
rect 15547 2158 15584 2229
rect 15739 2204 15770 2269
rect 16084 2222 16119 2300
rect 16696 2290 16733 2313
rect 17489 2331 17527 2340
rect 17489 2311 17498 2331
rect 17518 2311 17527 2331
rect 17489 2303 17527 2311
rect 17593 2335 17678 2341
rect 17703 2340 17740 2341
rect 17593 2315 17601 2335
rect 17621 2315 17678 2335
rect 17593 2307 17678 2315
rect 17702 2331 17740 2340
rect 17702 2311 17711 2331
rect 17731 2311 17740 2331
rect 17593 2306 17629 2307
rect 17702 2303 17740 2311
rect 17806 2335 17891 2341
rect 17911 2340 17948 2341
rect 17806 2315 17814 2335
rect 17834 2334 17891 2335
rect 17834 2315 17863 2334
rect 17806 2314 17863 2315
rect 17884 2314 17891 2334
rect 17806 2307 17891 2314
rect 17910 2331 17948 2340
rect 17910 2311 17919 2331
rect 17939 2311 17948 2331
rect 17806 2306 17842 2307
rect 17910 2303 17948 2311
rect 18014 2335 18158 2341
rect 18014 2315 18022 2335
rect 18042 2316 18078 2335
rect 18101 2316 18130 2335
rect 18042 2315 18130 2316
rect 18150 2315 18158 2335
rect 18014 2307 18158 2315
rect 18014 2306 18050 2307
rect 18122 2306 18158 2307
rect 18224 2340 18261 2341
rect 18224 2339 18262 2340
rect 18224 2331 18288 2339
rect 18224 2311 18233 2331
rect 18253 2317 18288 2331
rect 18308 2317 18311 2337
rect 18253 2312 18311 2317
rect 18253 2311 18288 2312
rect 16080 2213 16119 2222
rect 15738 2194 15775 2204
rect 15738 2192 15748 2194
rect 15672 2190 15748 2192
rect 15334 2134 15584 2158
rect 15669 2176 15748 2190
rect 15766 2176 15775 2194
rect 16080 2195 16090 2213
rect 16108 2195 16119 2213
rect 16080 2189 16119 2195
rect 16275 2265 16525 2289
rect 16275 2194 16312 2265
rect 16427 2204 16458 2205
rect 16080 2185 16117 2189
rect 15669 2173 15775 2176
rect 15141 2114 15162 2133
rect 15669 2114 15695 2173
rect 15738 2167 15775 2173
rect 16275 2174 16284 2194
rect 16304 2174 16312 2194
rect 16275 2164 16312 2174
rect 16371 2194 16458 2204
rect 16371 2174 16380 2194
rect 16400 2174 16458 2194
rect 16371 2165 16458 2174
rect 16371 2164 16408 2165
rect 16083 2114 16120 2123
rect 13795 2109 13895 2113
rect 13795 2105 13857 2109
rect 13795 2079 13802 2105
rect 13828 2083 13857 2105
rect 13883 2083 13895 2109
rect 13828 2079 13895 2083
rect 13795 2076 13895 2079
rect 13963 2076 13998 2113
rect 14060 2110 14419 2113
rect 14060 2105 14282 2110
rect 14060 2081 14073 2105
rect 14097 2086 14282 2105
rect 14306 2086 14419 2110
rect 14097 2081 14419 2086
rect 14060 2077 14419 2081
rect 14486 2105 14635 2113
rect 14486 2085 14497 2105
rect 14517 2085 14635 2105
rect 15141 2096 15695 2114
rect 15741 2103 15778 2105
rect 15669 2095 15695 2096
rect 15738 2095 15778 2103
rect 14486 2078 14635 2085
rect 15738 2083 15750 2095
rect 15729 2078 15750 2083
rect 14486 2077 14527 2078
rect 15145 2077 15750 2078
rect 15768 2077 15778 2095
rect 13810 2024 13847 2025
rect 13906 2024 13943 2025
rect 13962 2024 13998 2076
rect 14017 2024 14054 2025
rect 13710 2015 13848 2024
rect 13710 1995 13819 2015
rect 13839 1995 13848 2015
rect 13710 1988 13848 1995
rect 13906 2015 14054 2024
rect 13906 1995 13915 2015
rect 13935 1995 14025 2015
rect 14045 1995 14054 2015
rect 13710 1986 13806 1988
rect 13906 1985 14054 1995
rect 14113 2015 14150 2025
rect 14225 2024 14262 2025
rect 14206 2022 14262 2024
rect 14113 1995 14121 2015
rect 14141 1995 14150 2015
rect 13962 1984 13998 1985
rect 13810 1925 13847 1926
rect 14113 1925 14150 1995
rect 14175 2015 14262 2022
rect 14175 2012 14233 2015
rect 14175 1992 14180 2012
rect 14201 1995 14233 2012
rect 14253 1995 14262 2015
rect 14201 1992 14262 1995
rect 14175 1985 14262 1992
rect 14321 2015 14358 2025
rect 14321 1995 14329 2015
rect 14349 1995 14358 2015
rect 14175 1984 14206 1985
rect 13809 1924 14150 1925
rect 13734 1919 14150 1924
rect 13734 1899 13737 1919
rect 13757 1899 14150 1919
rect 14321 1924 14358 1995
rect 14388 2024 14419 2077
rect 15145 2068 15778 2077
rect 16081 2096 16092 2114
rect 16110 2096 16120 2114
rect 16427 2112 16458 2165
rect 16488 2194 16525 2265
rect 16696 2270 17089 2290
rect 17109 2270 17112 2290
rect 17490 2274 17527 2303
rect 16696 2265 17112 2270
rect 17491 2272 17527 2274
rect 17703 2272 17740 2303
rect 16696 2264 17037 2265
rect 16640 2204 16671 2205
rect 16488 2174 16497 2194
rect 16517 2174 16525 2194
rect 16488 2164 16525 2174
rect 16584 2197 16671 2204
rect 16584 2194 16645 2197
rect 16584 2174 16593 2194
rect 16613 2177 16645 2194
rect 16666 2177 16671 2197
rect 16613 2174 16671 2177
rect 16584 2167 16671 2174
rect 16696 2194 16733 2264
rect 16999 2263 17036 2264
rect 17491 2250 17740 2272
rect 17911 2271 17948 2303
rect 18224 2299 18288 2311
rect 18328 2273 18355 2451
rect 18383 2338 18421 4169
rect 18928 4144 18935 4170
rect 18954 4144 18959 4170
rect 18835 3751 18864 3753
rect 18835 3746 18867 3751
rect 18835 3728 18842 3746
rect 18862 3728 18867 3746
rect 18928 3750 18959 4144
rect 18980 4169 19148 4170
rect 18980 4166 19424 4169
rect 18980 4147 19355 4166
rect 19375 4147 19424 4166
rect 19992 4168 20101 4188
rect 20121 4168 20130 4188
rect 18980 4143 19424 4147
rect 18980 4141 19148 4143
rect 18980 3963 19007 4141
rect 19047 4103 19111 4115
rect 19387 4111 19424 4143
rect 19595 4142 19844 4164
rect 19992 4161 20130 4168
rect 20188 4188 20336 4197
rect 20188 4168 20197 4188
rect 20217 4168 20307 4188
rect 20327 4168 20336 4188
rect 19992 4159 20088 4161
rect 20188 4158 20336 4168
rect 20395 4188 20432 4198
rect 20507 4197 20544 4198
rect 20488 4195 20544 4197
rect 20395 4168 20403 4188
rect 20423 4168 20432 4188
rect 20244 4157 20280 4158
rect 19595 4111 19632 4142
rect 19808 4140 19844 4142
rect 19808 4111 19845 4140
rect 19047 4102 19082 4103
rect 19024 4097 19082 4102
rect 19024 4077 19027 4097
rect 19047 4083 19082 4097
rect 19102 4083 19111 4103
rect 19047 4075 19111 4083
rect 19073 4074 19111 4075
rect 19074 4073 19111 4074
rect 19177 4107 19213 4108
rect 19285 4107 19321 4108
rect 19177 4099 19321 4107
rect 19177 4079 19185 4099
rect 19205 4098 19293 4099
rect 19205 4079 19238 4098
rect 19177 4078 19238 4079
rect 19262 4079 19293 4098
rect 19313 4079 19321 4099
rect 19262 4078 19321 4079
rect 19177 4073 19321 4078
rect 19387 4103 19425 4111
rect 19493 4107 19529 4108
rect 19387 4083 19396 4103
rect 19416 4083 19425 4103
rect 19387 4074 19425 4083
rect 19444 4100 19529 4107
rect 19444 4080 19451 4100
rect 19472 4099 19529 4100
rect 19472 4080 19501 4099
rect 19444 4079 19501 4080
rect 19521 4079 19529 4099
rect 19387 4073 19424 4074
rect 19444 4073 19529 4079
rect 19595 4103 19633 4111
rect 19706 4107 19742 4108
rect 19595 4083 19604 4103
rect 19624 4083 19633 4103
rect 19595 4074 19633 4083
rect 19657 4099 19742 4107
rect 19657 4079 19714 4099
rect 19734 4079 19742 4099
rect 19595 4073 19632 4074
rect 19657 4073 19742 4079
rect 19808 4103 19846 4111
rect 19808 4083 19817 4103
rect 19837 4083 19846 4103
rect 20092 4098 20129 4099
rect 20395 4098 20432 4168
rect 20457 4188 20544 4195
rect 20457 4185 20515 4188
rect 20457 4165 20462 4185
rect 20483 4168 20515 4185
rect 20535 4168 20544 4188
rect 20483 4165 20544 4168
rect 20457 4158 20544 4165
rect 20603 4188 20640 4198
rect 20603 4168 20611 4188
rect 20631 4168 20640 4188
rect 20457 4157 20488 4158
rect 20091 4097 20432 4098
rect 19808 4074 19846 4083
rect 20016 4092 20432 4097
rect 19808 4073 19845 4074
rect 19231 4052 19267 4073
rect 19657 4052 19688 4073
rect 20016 4072 20019 4092
rect 20039 4072 20432 4092
rect 20603 4097 20640 4168
rect 20670 4197 20701 4250
rect 21003 4235 21040 4245
rect 21003 4217 21012 4235
rect 21030 4217 21040 4235
rect 21003 4208 21040 4217
rect 20720 4197 20757 4198
rect 20670 4188 20757 4197
rect 20670 4168 20728 4188
rect 20748 4168 20757 4188
rect 20670 4158 20757 4168
rect 20816 4188 20853 4198
rect 20816 4168 20824 4188
rect 20844 4168 20853 4188
rect 20670 4157 20701 4158
rect 20816 4097 20853 4168
rect 21008 4143 21039 4208
rect 21007 4133 21044 4143
rect 21007 4131 21017 4133
rect 20941 4129 21017 4131
rect 20603 4073 20853 4097
rect 20938 4115 21017 4129
rect 21035 4115 21044 4133
rect 20938 4112 21044 4115
rect 20410 4053 20431 4072
rect 20938 4053 20964 4112
rect 21007 4106 21044 4112
rect 19064 4048 19164 4052
rect 19064 4044 19126 4048
rect 19064 4018 19071 4044
rect 19097 4022 19126 4044
rect 19152 4022 19164 4048
rect 19097 4018 19164 4022
rect 19064 4015 19164 4018
rect 19232 4015 19267 4052
rect 19329 4049 19688 4052
rect 19329 4044 19551 4049
rect 19329 4020 19342 4044
rect 19366 4025 19551 4044
rect 19575 4025 19688 4049
rect 19366 4020 19688 4025
rect 19329 4016 19688 4020
rect 19755 4044 19904 4052
rect 19755 4024 19766 4044
rect 19786 4024 19904 4044
rect 20410 4035 20964 4053
rect 21010 4042 21047 4044
rect 20938 4034 20964 4035
rect 21007 4034 21047 4042
rect 19755 4017 19904 4024
rect 21007 4022 21019 4034
rect 20998 4017 21019 4022
rect 19755 4016 19796 4017
rect 20414 4016 21019 4017
rect 21037 4016 21047 4034
rect 19079 3963 19116 3964
rect 19175 3963 19212 3964
rect 19231 3963 19267 4015
rect 19286 3963 19323 3964
rect 18979 3954 19117 3963
rect 18979 3934 19088 3954
rect 19108 3934 19117 3954
rect 18979 3927 19117 3934
rect 19175 3954 19323 3963
rect 19175 3934 19184 3954
rect 19204 3934 19294 3954
rect 19314 3934 19323 3954
rect 18979 3925 19075 3927
rect 19175 3924 19323 3934
rect 19382 3954 19419 3964
rect 19494 3963 19531 3964
rect 19475 3961 19531 3963
rect 19382 3934 19390 3954
rect 19410 3934 19419 3954
rect 19231 3923 19267 3924
rect 19079 3864 19116 3865
rect 19382 3864 19419 3934
rect 19444 3954 19531 3961
rect 19444 3951 19502 3954
rect 19444 3931 19449 3951
rect 19470 3934 19502 3951
rect 19522 3934 19531 3954
rect 19470 3931 19531 3934
rect 19444 3924 19531 3931
rect 19590 3954 19627 3964
rect 19590 3934 19598 3954
rect 19618 3934 19627 3954
rect 19444 3923 19475 3924
rect 19078 3863 19419 3864
rect 19003 3858 19419 3863
rect 19003 3838 19006 3858
rect 19026 3838 19419 3858
rect 19590 3863 19627 3934
rect 19657 3963 19688 4016
rect 20414 4007 21047 4016
rect 20414 4000 21046 4007
rect 20414 3998 20476 4000
rect 19992 3988 20160 3989
rect 20414 3988 20436 3998
rect 19707 3963 19744 3964
rect 19657 3954 19744 3963
rect 19657 3934 19715 3954
rect 19735 3934 19744 3954
rect 19657 3924 19744 3934
rect 19803 3954 19840 3964
rect 19803 3934 19811 3954
rect 19831 3934 19840 3954
rect 19657 3923 19688 3924
rect 19803 3863 19840 3934
rect 19590 3839 19840 3863
rect 19992 3962 20436 3988
rect 19992 3960 20160 3962
rect 19992 3782 20019 3960
rect 20059 3922 20123 3934
rect 20399 3930 20436 3962
rect 20607 3961 20856 3983
rect 20607 3930 20644 3961
rect 20820 3959 20856 3961
rect 20820 3930 20857 3959
rect 20059 3921 20094 3922
rect 20036 3916 20094 3921
rect 20036 3896 20039 3916
rect 20059 3902 20094 3916
rect 20114 3902 20123 3922
rect 20059 3894 20123 3902
rect 20085 3893 20123 3894
rect 20086 3892 20123 3893
rect 20189 3926 20225 3927
rect 20297 3926 20333 3927
rect 20189 3918 20333 3926
rect 20189 3898 20197 3918
rect 20217 3898 20246 3918
rect 20189 3897 20246 3898
rect 20268 3898 20305 3918
rect 20325 3898 20333 3918
rect 20268 3897 20333 3898
rect 20189 3892 20333 3897
rect 20399 3922 20437 3930
rect 20505 3926 20541 3927
rect 20399 3902 20408 3922
rect 20428 3902 20437 3922
rect 20399 3893 20437 3902
rect 20456 3919 20541 3926
rect 20456 3899 20463 3919
rect 20484 3918 20541 3919
rect 20484 3899 20513 3918
rect 20456 3898 20513 3899
rect 20533 3898 20541 3918
rect 20399 3892 20436 3893
rect 20456 3892 20541 3898
rect 20607 3922 20645 3930
rect 20718 3926 20754 3927
rect 20607 3902 20616 3922
rect 20636 3902 20645 3922
rect 20607 3893 20645 3902
rect 20669 3918 20754 3926
rect 20669 3898 20726 3918
rect 20746 3898 20754 3918
rect 20607 3892 20644 3893
rect 20669 3892 20754 3898
rect 20820 3922 20858 3930
rect 20820 3902 20829 3922
rect 20849 3902 20858 3922
rect 20820 3893 20858 3902
rect 20820 3892 20857 3893
rect 20243 3871 20279 3892
rect 20669 3871 20700 3892
rect 20076 3867 20176 3871
rect 20076 3863 20138 3867
rect 20076 3837 20083 3863
rect 20109 3841 20138 3863
rect 20164 3841 20176 3867
rect 20109 3837 20176 3841
rect 20076 3834 20176 3837
rect 20244 3834 20279 3871
rect 20341 3868 20700 3871
rect 20341 3863 20563 3868
rect 20341 3839 20354 3863
rect 20378 3844 20563 3863
rect 20587 3844 20700 3868
rect 20378 3839 20700 3844
rect 20341 3835 20700 3839
rect 20767 3863 20916 3871
rect 20767 3843 20778 3863
rect 20798 3843 20916 3863
rect 20767 3836 20916 3843
rect 21007 3851 21046 4000
rect 20767 3835 20808 3836
rect 20091 3782 20128 3783
rect 20187 3782 20224 3783
rect 20243 3782 20279 3834
rect 20298 3782 20335 3783
rect 19991 3773 20129 3782
rect 19991 3753 20100 3773
rect 20120 3753 20129 3773
rect 18928 3749 19098 3750
rect 18928 3734 19374 3749
rect 19991 3746 20129 3753
rect 20187 3773 20335 3782
rect 20187 3753 20196 3773
rect 20216 3753 20306 3773
rect 20326 3753 20335 3773
rect 19991 3744 20087 3746
rect 18835 3723 18867 3728
rect 18837 2722 18867 3723
rect 18930 3723 19374 3734
rect 18930 3721 19098 3723
rect 18930 3543 18957 3721
rect 18997 3683 19061 3695
rect 19337 3691 19374 3723
rect 19545 3722 19794 3744
rect 20187 3743 20335 3753
rect 20394 3773 20431 3783
rect 20506 3782 20543 3783
rect 20487 3780 20543 3782
rect 20394 3753 20402 3773
rect 20422 3753 20431 3773
rect 20243 3742 20279 3743
rect 19545 3691 19582 3722
rect 19758 3720 19794 3722
rect 19758 3691 19795 3720
rect 18997 3682 19032 3683
rect 18974 3677 19032 3682
rect 18974 3657 18977 3677
rect 18997 3663 19032 3677
rect 19052 3663 19061 3683
rect 18997 3655 19061 3663
rect 19023 3654 19061 3655
rect 19024 3653 19061 3654
rect 19127 3687 19163 3688
rect 19235 3687 19271 3688
rect 19127 3679 19271 3687
rect 19127 3659 19135 3679
rect 19155 3660 19187 3679
rect 19210 3660 19243 3679
rect 19155 3659 19243 3660
rect 19263 3659 19271 3679
rect 19127 3653 19271 3659
rect 19337 3683 19375 3691
rect 19443 3687 19479 3688
rect 19337 3663 19346 3683
rect 19366 3663 19375 3683
rect 19337 3654 19375 3663
rect 19394 3680 19479 3687
rect 19394 3660 19401 3680
rect 19422 3679 19479 3680
rect 19422 3660 19451 3679
rect 19394 3659 19451 3660
rect 19471 3659 19479 3679
rect 19337 3653 19374 3654
rect 19394 3653 19479 3659
rect 19545 3683 19583 3691
rect 19656 3687 19692 3688
rect 19545 3663 19554 3683
rect 19574 3663 19583 3683
rect 19545 3654 19583 3663
rect 19607 3679 19692 3687
rect 19607 3659 19664 3679
rect 19684 3659 19692 3679
rect 19545 3653 19582 3654
rect 19607 3653 19692 3659
rect 19758 3683 19796 3691
rect 20091 3683 20128 3684
rect 20394 3683 20431 3753
rect 20456 3773 20543 3780
rect 20456 3770 20514 3773
rect 20456 3750 20461 3770
rect 20482 3753 20514 3770
rect 20534 3753 20543 3773
rect 20482 3750 20543 3753
rect 20456 3743 20543 3750
rect 20602 3773 20639 3783
rect 20602 3753 20610 3773
rect 20630 3753 20639 3773
rect 20456 3742 20487 3743
rect 19758 3663 19767 3683
rect 19787 3663 19796 3683
rect 20090 3682 20431 3683
rect 19758 3654 19796 3663
rect 20015 3677 20431 3682
rect 20015 3657 20018 3677
rect 20038 3657 20431 3677
rect 20602 3682 20639 3753
rect 20669 3782 20700 3835
rect 21007 3833 21017 3851
rect 21035 3833 21046 3851
rect 21007 3824 21044 3833
rect 20719 3782 20756 3783
rect 20669 3773 20756 3782
rect 20669 3753 20727 3773
rect 20747 3753 20756 3773
rect 20669 3743 20756 3753
rect 20815 3773 20852 3783
rect 20815 3753 20823 3773
rect 20843 3753 20852 3773
rect 21010 3758 21047 3762
rect 20669 3742 20700 3743
rect 20815 3682 20852 3753
rect 20602 3658 20852 3682
rect 21008 3752 21047 3758
rect 21008 3734 21019 3752
rect 21037 3734 21047 3752
rect 21008 3725 21047 3734
rect 19758 3653 19795 3654
rect 19181 3632 19217 3653
rect 19607 3632 19638 3653
rect 20394 3634 20431 3657
rect 21008 3647 21043 3725
rect 21005 3637 21043 3647
rect 20394 3633 20564 3634
rect 21005 3633 21015 3637
rect 19014 3628 19114 3632
rect 19014 3624 19076 3628
rect 19014 3598 19021 3624
rect 19047 3602 19076 3624
rect 19102 3602 19114 3628
rect 19047 3598 19114 3602
rect 19014 3595 19114 3598
rect 19182 3595 19217 3632
rect 19279 3629 19638 3632
rect 19279 3624 19501 3629
rect 19279 3600 19292 3624
rect 19316 3605 19501 3624
rect 19525 3605 19638 3629
rect 19316 3600 19638 3605
rect 19279 3596 19638 3600
rect 19705 3624 19854 3632
rect 19705 3604 19716 3624
rect 19736 3604 19854 3624
rect 20394 3619 21015 3633
rect 21033 3619 21043 3637
rect 20394 3613 21043 3619
rect 20394 3612 21042 3613
rect 21005 3610 21042 3612
rect 19705 3597 19854 3604
rect 19705 3596 19746 3597
rect 19029 3543 19066 3544
rect 19125 3543 19162 3544
rect 19181 3543 19217 3595
rect 19236 3543 19273 3544
rect 18929 3534 19067 3543
rect 18929 3514 19038 3534
rect 19058 3514 19067 3534
rect 18929 3507 19067 3514
rect 19125 3534 19273 3543
rect 19125 3514 19134 3534
rect 19154 3514 19244 3534
rect 19264 3514 19273 3534
rect 18929 3505 19025 3507
rect 19125 3504 19273 3514
rect 19332 3534 19369 3544
rect 19444 3543 19481 3544
rect 19425 3541 19481 3543
rect 19332 3514 19340 3534
rect 19360 3514 19369 3534
rect 19181 3503 19217 3504
rect 19029 3444 19066 3445
rect 19332 3444 19369 3514
rect 19394 3534 19481 3541
rect 19394 3531 19452 3534
rect 19394 3511 19399 3531
rect 19420 3514 19452 3531
rect 19472 3514 19481 3534
rect 19420 3511 19481 3514
rect 19394 3504 19481 3511
rect 19540 3534 19577 3544
rect 19540 3514 19548 3534
rect 19568 3514 19577 3534
rect 19394 3503 19425 3504
rect 19028 3443 19369 3444
rect 18953 3438 19369 3443
rect 18953 3418 18956 3438
rect 18976 3418 19369 3438
rect 19540 3443 19577 3514
rect 19607 3543 19638 3596
rect 19657 3543 19694 3544
rect 19607 3534 19694 3543
rect 19607 3514 19665 3534
rect 19685 3514 19694 3534
rect 19607 3504 19694 3514
rect 19753 3534 19790 3544
rect 19753 3514 19761 3534
rect 19781 3514 19790 3534
rect 19607 3503 19638 3504
rect 19753 3443 19790 3514
rect 21008 3538 21045 3548
rect 21008 3520 21017 3538
rect 21035 3520 21045 3538
rect 21008 3511 21045 3520
rect 21008 3487 21043 3511
rect 21006 3463 21043 3487
rect 21005 3457 21043 3463
rect 19540 3419 19790 3443
rect 20416 3439 21043 3457
rect 19998 3422 20166 3423
rect 20417 3422 20441 3439
rect 19998 3396 20442 3422
rect 19998 3394 20166 3396
rect 19998 3216 20025 3394
rect 20065 3356 20129 3368
rect 20405 3364 20442 3396
rect 20613 3395 20862 3417
rect 20613 3364 20650 3395
rect 20826 3393 20862 3395
rect 21005 3398 21043 3439
rect 20826 3364 20863 3393
rect 20065 3355 20100 3356
rect 20042 3350 20100 3355
rect 20042 3330 20045 3350
rect 20065 3336 20100 3350
rect 20120 3336 20129 3356
rect 20065 3328 20129 3336
rect 20091 3327 20129 3328
rect 20092 3326 20129 3327
rect 20195 3360 20231 3361
rect 20303 3360 20339 3361
rect 20195 3354 20339 3360
rect 20195 3352 20261 3354
rect 20195 3332 20203 3352
rect 20223 3333 20261 3352
rect 20283 3352 20339 3354
rect 20283 3333 20311 3352
rect 20223 3332 20311 3333
rect 20331 3332 20339 3352
rect 20195 3326 20339 3332
rect 20405 3356 20443 3364
rect 20511 3360 20547 3361
rect 20405 3336 20414 3356
rect 20434 3336 20443 3356
rect 20405 3327 20443 3336
rect 20462 3353 20547 3360
rect 20462 3333 20469 3353
rect 20490 3352 20547 3353
rect 20490 3333 20519 3352
rect 20462 3332 20519 3333
rect 20539 3332 20547 3352
rect 20405 3326 20442 3327
rect 20462 3326 20547 3332
rect 20613 3356 20651 3364
rect 20724 3360 20760 3361
rect 20613 3336 20622 3356
rect 20642 3336 20651 3356
rect 20613 3327 20651 3336
rect 20675 3352 20760 3360
rect 20675 3332 20732 3352
rect 20752 3332 20760 3352
rect 20613 3326 20650 3327
rect 20675 3326 20760 3332
rect 20826 3356 20864 3364
rect 20826 3336 20835 3356
rect 20855 3336 20864 3356
rect 20826 3327 20864 3336
rect 21005 3363 21041 3398
rect 21005 3353 21042 3363
rect 21005 3335 21015 3353
rect 21033 3335 21042 3353
rect 20826 3326 20863 3327
rect 21005 3326 21042 3335
rect 20249 3305 20285 3326
rect 20675 3305 20706 3326
rect 20082 3301 20182 3305
rect 20082 3297 20144 3301
rect 20082 3271 20089 3297
rect 20115 3275 20144 3297
rect 20170 3275 20182 3301
rect 20115 3271 20182 3275
rect 20082 3268 20182 3271
rect 20250 3268 20285 3305
rect 20347 3302 20706 3305
rect 20347 3297 20569 3302
rect 20347 3273 20360 3297
rect 20384 3278 20569 3297
rect 20593 3278 20706 3302
rect 20384 3273 20706 3278
rect 20347 3269 20706 3273
rect 20773 3297 20922 3305
rect 20773 3277 20784 3297
rect 20804 3277 20922 3297
rect 20773 3270 20922 3277
rect 20773 3269 20814 3270
rect 20097 3216 20134 3217
rect 20193 3216 20230 3217
rect 20249 3216 20285 3268
rect 20304 3216 20341 3217
rect 19997 3207 20135 3216
rect 18985 3188 19153 3189
rect 18985 3185 19429 3188
rect 18985 3166 19360 3185
rect 19380 3166 19429 3185
rect 19997 3187 20106 3207
rect 20126 3187 20135 3207
rect 18985 3162 19429 3166
rect 18985 3160 19153 3162
rect 18985 2982 19012 3160
rect 19052 3122 19116 3134
rect 19392 3130 19429 3162
rect 19600 3161 19849 3183
rect 19997 3180 20135 3187
rect 20193 3207 20341 3216
rect 20193 3187 20202 3207
rect 20222 3187 20312 3207
rect 20332 3187 20341 3207
rect 19997 3178 20093 3180
rect 20193 3177 20341 3187
rect 20400 3207 20437 3217
rect 20512 3216 20549 3217
rect 20493 3214 20549 3216
rect 20400 3187 20408 3207
rect 20428 3187 20437 3207
rect 20249 3176 20285 3177
rect 19600 3130 19637 3161
rect 19813 3159 19849 3161
rect 19813 3130 19850 3159
rect 19052 3121 19087 3122
rect 19029 3116 19087 3121
rect 19029 3096 19032 3116
rect 19052 3102 19087 3116
rect 19107 3102 19116 3122
rect 19052 3094 19116 3102
rect 19078 3093 19116 3094
rect 19079 3092 19116 3093
rect 19182 3126 19218 3127
rect 19290 3126 19326 3127
rect 19182 3118 19326 3126
rect 19182 3098 19190 3118
rect 19210 3098 19242 3118
rect 19266 3098 19298 3118
rect 19318 3098 19326 3118
rect 19182 3092 19326 3098
rect 19392 3122 19430 3130
rect 19498 3126 19534 3127
rect 19392 3102 19401 3122
rect 19421 3102 19430 3122
rect 19392 3093 19430 3102
rect 19449 3119 19534 3126
rect 19449 3099 19456 3119
rect 19477 3118 19534 3119
rect 19477 3099 19506 3118
rect 19449 3098 19506 3099
rect 19526 3098 19534 3118
rect 19392 3092 19429 3093
rect 19449 3092 19534 3098
rect 19600 3122 19638 3130
rect 19711 3126 19747 3127
rect 19600 3102 19609 3122
rect 19629 3102 19638 3122
rect 19600 3093 19638 3102
rect 19662 3118 19747 3126
rect 19662 3098 19719 3118
rect 19739 3098 19747 3118
rect 19600 3092 19637 3093
rect 19662 3092 19747 3098
rect 19813 3122 19851 3130
rect 19813 3102 19822 3122
rect 19842 3102 19851 3122
rect 20097 3117 20134 3118
rect 20400 3117 20437 3187
rect 20462 3207 20549 3214
rect 20462 3204 20520 3207
rect 20462 3184 20467 3204
rect 20488 3187 20520 3204
rect 20540 3187 20549 3207
rect 20488 3184 20549 3187
rect 20462 3177 20549 3184
rect 20608 3207 20645 3217
rect 20608 3187 20616 3207
rect 20636 3187 20645 3207
rect 20462 3176 20493 3177
rect 20096 3116 20437 3117
rect 19813 3093 19851 3102
rect 20021 3111 20437 3116
rect 19813 3092 19850 3093
rect 19236 3071 19272 3092
rect 19662 3071 19693 3092
rect 20021 3091 20024 3111
rect 20044 3091 20437 3111
rect 20608 3116 20645 3187
rect 20675 3216 20706 3269
rect 21008 3254 21045 3264
rect 21008 3236 21017 3254
rect 21035 3236 21045 3254
rect 21008 3227 21045 3236
rect 20725 3216 20762 3217
rect 20675 3207 20762 3216
rect 20675 3187 20733 3207
rect 20753 3187 20762 3207
rect 20675 3177 20762 3187
rect 20821 3207 20858 3217
rect 20821 3187 20829 3207
rect 20849 3187 20858 3207
rect 20675 3176 20706 3177
rect 20821 3116 20858 3187
rect 21013 3162 21044 3227
rect 21012 3152 21049 3162
rect 21012 3150 21022 3152
rect 20946 3148 21022 3150
rect 20608 3092 20858 3116
rect 20943 3134 21022 3148
rect 21040 3134 21049 3152
rect 20943 3131 21049 3134
rect 20415 3072 20436 3091
rect 20943 3072 20969 3131
rect 21012 3125 21049 3131
rect 19069 3067 19169 3071
rect 19069 3063 19131 3067
rect 19069 3037 19076 3063
rect 19102 3041 19131 3063
rect 19157 3041 19169 3067
rect 19102 3037 19169 3041
rect 19069 3034 19169 3037
rect 19237 3034 19272 3071
rect 19334 3068 19693 3071
rect 19334 3063 19556 3068
rect 19334 3039 19347 3063
rect 19371 3044 19556 3063
rect 19580 3044 19693 3068
rect 19371 3039 19693 3044
rect 19334 3035 19693 3039
rect 19760 3063 19909 3071
rect 19760 3043 19771 3063
rect 19791 3043 19909 3063
rect 20415 3054 20969 3072
rect 21015 3061 21052 3063
rect 20943 3053 20969 3054
rect 21012 3053 21052 3061
rect 19760 3036 19909 3043
rect 21012 3041 21024 3053
rect 21003 3036 21024 3041
rect 19760 3035 19801 3036
rect 20419 3035 21024 3036
rect 21042 3035 21052 3053
rect 19084 2982 19121 2983
rect 19180 2982 19217 2983
rect 19236 2982 19272 3034
rect 19291 2982 19328 2983
rect 18984 2973 19122 2982
rect 18984 2953 19093 2973
rect 19113 2953 19122 2973
rect 18984 2946 19122 2953
rect 19180 2973 19328 2982
rect 19180 2953 19189 2973
rect 19209 2953 19299 2973
rect 19319 2953 19328 2973
rect 18984 2944 19080 2946
rect 19180 2943 19328 2953
rect 19387 2973 19424 2983
rect 19499 2982 19536 2983
rect 19480 2980 19536 2982
rect 19387 2953 19395 2973
rect 19415 2953 19424 2973
rect 19236 2942 19272 2943
rect 19084 2883 19121 2884
rect 19387 2883 19424 2953
rect 19449 2973 19536 2980
rect 19449 2970 19507 2973
rect 19449 2950 19454 2970
rect 19475 2953 19507 2970
rect 19527 2953 19536 2973
rect 19475 2950 19536 2953
rect 19449 2943 19536 2950
rect 19595 2973 19632 2983
rect 19595 2953 19603 2973
rect 19623 2953 19632 2973
rect 19449 2942 19480 2943
rect 19083 2882 19424 2883
rect 19008 2877 19424 2882
rect 19008 2857 19011 2877
rect 19031 2857 19424 2877
rect 19595 2882 19632 2953
rect 19662 2982 19693 3035
rect 20419 3026 21052 3035
rect 20419 3019 21051 3026
rect 20419 3017 20481 3019
rect 19997 3007 20165 3008
rect 20419 3007 20441 3017
rect 19712 2982 19749 2983
rect 19662 2973 19749 2982
rect 19662 2953 19720 2973
rect 19740 2953 19749 2973
rect 19662 2943 19749 2953
rect 19808 2973 19845 2983
rect 19808 2953 19816 2973
rect 19836 2953 19845 2973
rect 19662 2942 19693 2943
rect 19808 2882 19845 2953
rect 19595 2858 19845 2882
rect 19997 2981 20441 3007
rect 19997 2979 20165 2981
rect 19997 2801 20024 2979
rect 20064 2941 20128 2953
rect 20404 2949 20441 2981
rect 20612 2980 20861 3002
rect 20612 2949 20649 2980
rect 20825 2978 20861 2980
rect 20825 2949 20862 2978
rect 20064 2940 20099 2941
rect 20041 2935 20099 2940
rect 20041 2915 20044 2935
rect 20064 2921 20099 2935
rect 20119 2921 20128 2941
rect 20064 2913 20128 2921
rect 20090 2912 20128 2913
rect 20091 2911 20128 2912
rect 20194 2945 20230 2946
rect 20302 2945 20338 2946
rect 20194 2937 20338 2945
rect 20194 2917 20202 2937
rect 20222 2917 20251 2937
rect 20194 2916 20251 2917
rect 20273 2917 20310 2937
rect 20330 2917 20338 2937
rect 20273 2916 20338 2917
rect 20194 2911 20338 2916
rect 20404 2941 20442 2949
rect 20510 2945 20546 2946
rect 20404 2921 20413 2941
rect 20433 2921 20442 2941
rect 20404 2912 20442 2921
rect 20461 2938 20546 2945
rect 20461 2918 20468 2938
rect 20489 2937 20546 2938
rect 20489 2918 20518 2937
rect 20461 2917 20518 2918
rect 20538 2917 20546 2937
rect 20404 2911 20441 2912
rect 20461 2911 20546 2917
rect 20612 2941 20650 2949
rect 20723 2945 20759 2946
rect 20612 2921 20621 2941
rect 20641 2921 20650 2941
rect 20612 2912 20650 2921
rect 20674 2937 20759 2945
rect 20674 2917 20731 2937
rect 20751 2917 20759 2937
rect 20612 2911 20649 2912
rect 20674 2911 20759 2917
rect 20825 2941 20863 2949
rect 20825 2921 20834 2941
rect 20854 2921 20863 2941
rect 20825 2912 20863 2921
rect 20825 2911 20862 2912
rect 20248 2890 20284 2911
rect 20674 2890 20705 2911
rect 20081 2886 20181 2890
rect 20081 2882 20143 2886
rect 20081 2856 20088 2882
rect 20114 2860 20143 2882
rect 20169 2860 20181 2886
rect 20114 2856 20181 2860
rect 20081 2853 20181 2856
rect 20249 2853 20284 2890
rect 20346 2887 20705 2890
rect 20346 2882 20568 2887
rect 20346 2858 20359 2882
rect 20383 2863 20568 2882
rect 20592 2863 20705 2887
rect 20383 2858 20705 2863
rect 20346 2854 20705 2858
rect 20772 2882 20921 2890
rect 20772 2862 20783 2882
rect 20803 2862 20921 2882
rect 20772 2855 20921 2862
rect 21012 2870 21051 3019
rect 20772 2854 20813 2855
rect 20096 2801 20133 2802
rect 20192 2801 20229 2802
rect 20248 2801 20284 2853
rect 20303 2801 20340 2802
rect 19996 2792 20134 2801
rect 19996 2772 20105 2792
rect 20125 2772 20134 2792
rect 19996 2765 20134 2772
rect 20192 2792 20340 2801
rect 20192 2772 20201 2792
rect 20221 2772 20311 2792
rect 20331 2772 20340 2792
rect 19996 2763 20092 2765
rect 20192 2762 20340 2772
rect 20399 2792 20436 2802
rect 20511 2801 20548 2802
rect 20492 2799 20548 2801
rect 20399 2772 20407 2792
rect 20427 2772 20436 2792
rect 20248 2761 20284 2762
rect 18777 2721 18945 2722
rect 18777 2695 19221 2721
rect 18777 2693 18945 2695
rect 18777 2515 18804 2693
rect 18844 2655 18908 2667
rect 19184 2663 19221 2695
rect 19392 2694 19641 2716
rect 20096 2702 20133 2703
rect 20399 2702 20436 2772
rect 20461 2792 20548 2799
rect 20461 2789 20519 2792
rect 20461 2769 20466 2789
rect 20487 2772 20519 2789
rect 20539 2772 20548 2792
rect 20487 2769 20548 2772
rect 20461 2762 20548 2769
rect 20607 2792 20644 2802
rect 20607 2772 20615 2792
rect 20635 2772 20644 2792
rect 20461 2761 20492 2762
rect 20095 2701 20436 2702
rect 19392 2663 19429 2694
rect 19605 2692 19641 2694
rect 20020 2696 20436 2701
rect 19605 2663 19642 2692
rect 20020 2676 20023 2696
rect 20043 2676 20436 2696
rect 20607 2701 20644 2772
rect 20674 2801 20705 2854
rect 21012 2852 21022 2870
rect 21040 2852 21051 2870
rect 21012 2843 21049 2852
rect 20724 2801 20761 2802
rect 20674 2792 20761 2801
rect 20674 2772 20732 2792
rect 20752 2772 20761 2792
rect 20674 2762 20761 2772
rect 20820 2792 20857 2802
rect 20820 2772 20828 2792
rect 20848 2772 20857 2792
rect 21015 2777 21052 2781
rect 20674 2761 20705 2762
rect 20820 2701 20857 2772
rect 20607 2677 20857 2701
rect 21013 2771 21052 2777
rect 21013 2753 21024 2771
rect 21042 2753 21052 2771
rect 21013 2744 21052 2753
rect 18844 2654 18879 2655
rect 18821 2649 18879 2654
rect 18821 2629 18824 2649
rect 18844 2635 18879 2649
rect 18899 2635 18908 2655
rect 18844 2627 18908 2635
rect 18870 2626 18908 2627
rect 18871 2625 18908 2626
rect 18974 2659 19010 2660
rect 19082 2659 19118 2660
rect 18974 2653 19118 2659
rect 18974 2651 19035 2653
rect 18974 2631 18982 2651
rect 19002 2631 19035 2651
rect 18974 2627 19035 2631
rect 19060 2651 19118 2653
rect 19060 2631 19090 2651
rect 19110 2631 19118 2651
rect 19060 2627 19118 2631
rect 18974 2625 19118 2627
rect 19184 2655 19222 2663
rect 19290 2659 19326 2660
rect 19184 2635 19193 2655
rect 19213 2635 19222 2655
rect 19184 2626 19222 2635
rect 19241 2652 19326 2659
rect 19241 2632 19248 2652
rect 19269 2651 19326 2652
rect 19269 2632 19298 2651
rect 19241 2631 19298 2632
rect 19318 2631 19326 2651
rect 19184 2625 19221 2626
rect 19241 2625 19326 2631
rect 19392 2655 19430 2663
rect 19503 2659 19539 2660
rect 19392 2635 19401 2655
rect 19421 2635 19430 2655
rect 19392 2626 19430 2635
rect 19454 2651 19539 2659
rect 19454 2631 19511 2651
rect 19531 2631 19539 2651
rect 19392 2625 19429 2626
rect 19454 2625 19539 2631
rect 19605 2655 19643 2663
rect 19605 2635 19614 2655
rect 19634 2635 19643 2655
rect 19605 2626 19643 2635
rect 20399 2653 20436 2676
rect 21013 2666 21048 2744
rect 21010 2656 21048 2666
rect 20399 2652 20569 2653
rect 21010 2652 21020 2656
rect 20399 2638 21020 2652
rect 21038 2638 21048 2656
rect 20399 2632 21048 2638
rect 20399 2631 21047 2632
rect 21010 2629 21047 2631
rect 19605 2625 19642 2626
rect 19028 2604 19064 2625
rect 19454 2604 19485 2625
rect 18861 2600 18961 2604
rect 18861 2596 18923 2600
rect 18861 2570 18868 2596
rect 18894 2574 18923 2596
rect 18949 2574 18961 2600
rect 18894 2570 18961 2574
rect 18861 2567 18961 2570
rect 19029 2567 19064 2604
rect 19126 2601 19485 2604
rect 19126 2596 19348 2601
rect 19126 2572 19139 2596
rect 19163 2577 19348 2596
rect 19372 2577 19485 2601
rect 19163 2572 19485 2577
rect 19126 2568 19485 2572
rect 19552 2596 19701 2604
rect 19552 2576 19563 2596
rect 19583 2576 19701 2596
rect 19552 2569 19701 2576
rect 19552 2568 19593 2569
rect 18876 2515 18913 2516
rect 18972 2515 19009 2516
rect 19028 2515 19064 2567
rect 19083 2515 19120 2516
rect 18776 2506 18914 2515
rect 18776 2486 18885 2506
rect 18905 2486 18914 2506
rect 18776 2479 18914 2486
rect 18972 2506 19120 2515
rect 18972 2486 18981 2506
rect 19001 2486 19091 2506
rect 19111 2486 19120 2506
rect 18776 2477 18872 2479
rect 18972 2476 19120 2486
rect 19179 2506 19216 2516
rect 19291 2515 19328 2516
rect 19272 2513 19328 2515
rect 19179 2486 19187 2506
rect 19207 2486 19216 2506
rect 19028 2475 19064 2476
rect 18876 2416 18913 2417
rect 19179 2416 19216 2486
rect 19241 2506 19328 2513
rect 19241 2503 19299 2506
rect 19241 2483 19246 2503
rect 19267 2486 19299 2503
rect 19319 2486 19328 2506
rect 19267 2483 19328 2486
rect 19241 2476 19328 2483
rect 19387 2506 19424 2516
rect 19387 2486 19395 2506
rect 19415 2486 19424 2506
rect 19241 2475 19272 2476
rect 18875 2415 19216 2416
rect 18800 2410 19216 2415
rect 18800 2390 18803 2410
rect 18823 2390 19216 2410
rect 19387 2415 19424 2486
rect 19454 2515 19485 2568
rect 21013 2557 21050 2567
rect 21013 2539 21022 2557
rect 21040 2539 21050 2557
rect 21013 2530 21050 2539
rect 19504 2515 19541 2516
rect 19454 2506 19541 2515
rect 19454 2486 19512 2506
rect 19532 2486 19541 2506
rect 19454 2476 19541 2486
rect 19600 2506 19637 2516
rect 19600 2486 19608 2506
rect 19628 2486 19637 2506
rect 19454 2475 19485 2476
rect 19600 2415 19637 2486
rect 21013 2484 21048 2530
rect 21012 2478 21050 2484
rect 20423 2460 21050 2478
rect 19387 2391 19637 2415
rect 20005 2443 20173 2444
rect 20424 2443 20448 2460
rect 20005 2417 20449 2443
rect 20005 2415 20173 2417
rect 18385 2278 18418 2338
rect 18187 2271 18355 2273
rect 17911 2245 18355 2271
rect 18187 2244 18355 2245
rect 18384 2267 18421 2278
rect 18384 2248 18390 2267
rect 18413 2248 18421 2267
rect 16848 2204 16884 2205
rect 16696 2174 16705 2194
rect 16725 2174 16733 2194
rect 16584 2165 16640 2167
rect 16584 2164 16621 2165
rect 16696 2164 16733 2174
rect 16792 2194 16940 2204
rect 17040 2201 17136 2203
rect 16792 2174 16801 2194
rect 16821 2174 16911 2194
rect 16931 2174 16940 2194
rect 16792 2165 16940 2174
rect 16998 2194 17136 2201
rect 16998 2174 17007 2194
rect 17027 2174 17136 2194
rect 16998 2165 17136 2174
rect 16792 2164 16829 2165
rect 16848 2113 16884 2165
rect 16903 2164 16940 2165
rect 16999 2164 17036 2165
rect 16319 2111 16360 2112
rect 15145 2061 15777 2068
rect 15145 2059 15207 2061
rect 14723 2049 14891 2050
rect 15145 2049 15167 2059
rect 14438 2024 14475 2025
rect 14388 2015 14475 2024
rect 14388 1995 14446 2015
rect 14466 1995 14475 2015
rect 14388 1985 14475 1995
rect 14534 2015 14571 2025
rect 14534 1995 14542 2015
rect 14562 1995 14571 2015
rect 14388 1984 14419 1985
rect 14534 1924 14571 1995
rect 14321 1900 14571 1924
rect 14723 2023 15167 2049
rect 14723 2021 14891 2023
rect 14723 1843 14750 2021
rect 14790 1983 14854 1995
rect 15130 1991 15167 2023
rect 15338 2022 15587 2044
rect 15338 1991 15375 2022
rect 15551 2020 15587 2022
rect 15551 1991 15588 2020
rect 14790 1982 14825 1983
rect 14767 1977 14825 1982
rect 14767 1957 14770 1977
rect 14790 1963 14825 1977
rect 14845 1963 14854 1983
rect 14790 1955 14854 1963
rect 14816 1954 14854 1955
rect 14817 1953 14854 1954
rect 14920 1987 14956 1988
rect 15028 1987 15064 1988
rect 14920 1979 15064 1987
rect 14920 1959 14928 1979
rect 14948 1959 14977 1979
rect 14920 1958 14977 1959
rect 14999 1959 15036 1979
rect 15056 1959 15064 1979
rect 14999 1958 15064 1959
rect 14920 1953 15064 1958
rect 15130 1983 15168 1991
rect 15236 1987 15272 1988
rect 15130 1963 15139 1983
rect 15159 1963 15168 1983
rect 15130 1954 15168 1963
rect 15187 1980 15272 1987
rect 15187 1960 15194 1980
rect 15215 1979 15272 1980
rect 15215 1960 15244 1979
rect 15187 1959 15244 1960
rect 15264 1959 15272 1979
rect 15130 1953 15167 1954
rect 15187 1953 15272 1959
rect 15338 1983 15376 1991
rect 15449 1987 15485 1988
rect 15338 1963 15347 1983
rect 15367 1963 15376 1983
rect 15338 1954 15376 1963
rect 15400 1979 15485 1987
rect 15400 1959 15457 1979
rect 15477 1959 15485 1979
rect 15338 1953 15375 1954
rect 15400 1953 15485 1959
rect 15551 1983 15589 1991
rect 15551 1963 15560 1983
rect 15580 1963 15589 1983
rect 15551 1954 15589 1963
rect 15551 1953 15588 1954
rect 14974 1932 15010 1953
rect 15400 1932 15431 1953
rect 14807 1928 14907 1932
rect 14807 1924 14869 1928
rect 14807 1898 14814 1924
rect 14840 1902 14869 1924
rect 14895 1902 14907 1928
rect 14840 1898 14907 1902
rect 14807 1895 14907 1898
rect 14975 1895 15010 1932
rect 15072 1929 15431 1932
rect 15072 1924 15294 1929
rect 15072 1900 15085 1924
rect 15109 1905 15294 1924
rect 15318 1905 15431 1929
rect 15109 1900 15431 1905
rect 15072 1896 15431 1900
rect 15498 1924 15647 1932
rect 15498 1904 15509 1924
rect 15529 1904 15647 1924
rect 15498 1897 15647 1904
rect 15738 1912 15777 2061
rect 16081 1947 16120 2096
rect 16211 2104 16360 2111
rect 16211 2084 16329 2104
rect 16349 2084 16360 2104
rect 16211 2076 16360 2084
rect 16427 2108 16786 2112
rect 16427 2103 16749 2108
rect 16427 2079 16540 2103
rect 16564 2084 16749 2103
rect 16773 2084 16786 2108
rect 16564 2079 16786 2084
rect 16427 2076 16786 2079
rect 16848 2076 16883 2113
rect 16951 2110 17051 2113
rect 16951 2106 17018 2110
rect 16951 2080 16963 2106
rect 16989 2084 17018 2106
rect 17044 2084 17051 2110
rect 16989 2080 17051 2084
rect 16951 2076 17051 2080
rect 16427 2055 16458 2076
rect 16848 2055 16884 2076
rect 16270 2054 16307 2055
rect 16269 2045 16307 2054
rect 16269 2025 16278 2045
rect 16298 2025 16307 2045
rect 16269 2017 16307 2025
rect 16373 2049 16458 2055
rect 16483 2054 16520 2055
rect 16373 2029 16381 2049
rect 16401 2029 16458 2049
rect 16373 2021 16458 2029
rect 16482 2045 16520 2054
rect 16482 2025 16491 2045
rect 16511 2025 16520 2045
rect 16373 2020 16409 2021
rect 16482 2017 16520 2025
rect 16586 2049 16671 2055
rect 16691 2054 16728 2055
rect 16586 2029 16594 2049
rect 16614 2048 16671 2049
rect 16614 2029 16643 2048
rect 16586 2028 16643 2029
rect 16664 2028 16671 2048
rect 16586 2021 16671 2028
rect 16690 2045 16728 2054
rect 16690 2025 16699 2045
rect 16719 2025 16728 2045
rect 16586 2020 16622 2021
rect 16690 2017 16728 2025
rect 16794 2050 16938 2055
rect 16794 2049 16859 2050
rect 16794 2029 16802 2049
rect 16822 2029 16859 2049
rect 16881 2049 16938 2050
rect 16881 2029 16910 2049
rect 16930 2029 16938 2049
rect 16794 2021 16938 2029
rect 16794 2020 16830 2021
rect 16902 2020 16938 2021
rect 17004 2054 17041 2055
rect 17004 2053 17042 2054
rect 17004 2045 17068 2053
rect 17004 2025 17013 2045
rect 17033 2031 17068 2045
rect 17088 2031 17091 2051
rect 17033 2026 17091 2031
rect 17033 2025 17068 2026
rect 16270 1988 16307 2017
rect 16271 1986 16307 1988
rect 16483 1986 16520 2017
rect 16271 1964 16520 1986
rect 16691 1985 16728 2017
rect 17004 2013 17068 2025
rect 17108 1987 17135 2165
rect 16967 1985 17135 1987
rect 16691 1959 17135 1985
rect 17287 2084 17537 2108
rect 17287 2013 17324 2084
rect 17439 2023 17470 2024
rect 17287 1993 17296 2013
rect 17316 1993 17324 2013
rect 17287 1983 17324 1993
rect 17383 2013 17470 2023
rect 17383 1993 17392 2013
rect 17412 1993 17470 2013
rect 17383 1984 17470 1993
rect 17383 1983 17420 1984
rect 16691 1949 16713 1959
rect 16967 1958 17135 1959
rect 16651 1947 16713 1949
rect 16081 1940 16713 1947
rect 15498 1896 15539 1897
rect 14822 1843 14859 1844
rect 14918 1843 14955 1844
rect 14974 1843 15010 1895
rect 15029 1843 15066 1844
rect 14722 1834 14860 1843
rect 14722 1814 14831 1834
rect 14851 1814 14860 1834
rect 13659 1810 13829 1811
rect 13659 1795 14105 1810
rect 14722 1807 14860 1814
rect 14918 1834 15066 1843
rect 14918 1814 14927 1834
rect 14947 1814 15037 1834
rect 15057 1814 15066 1834
rect 14722 1805 14818 1807
rect 13661 1784 14105 1795
rect 13661 1782 13829 1784
rect 13661 1604 13688 1782
rect 13728 1744 13792 1756
rect 14068 1752 14105 1784
rect 14276 1783 14525 1805
rect 14918 1804 15066 1814
rect 15125 1834 15162 1844
rect 15237 1843 15274 1844
rect 15218 1841 15274 1843
rect 15125 1814 15133 1834
rect 15153 1814 15162 1834
rect 14974 1803 15010 1804
rect 14276 1752 14313 1783
rect 14489 1781 14525 1783
rect 14489 1752 14526 1781
rect 13728 1743 13763 1744
rect 13705 1738 13763 1743
rect 13705 1718 13708 1738
rect 13728 1724 13763 1738
rect 13783 1724 13792 1744
rect 13728 1716 13792 1724
rect 13754 1715 13792 1716
rect 13755 1714 13792 1715
rect 13858 1748 13894 1749
rect 13966 1748 14002 1749
rect 13858 1740 14002 1748
rect 13858 1720 13866 1740
rect 13886 1739 13974 1740
rect 13886 1722 13914 1739
rect 13938 1722 13974 1739
rect 13886 1720 13974 1722
rect 13994 1720 14002 1740
rect 13858 1714 14002 1720
rect 14068 1744 14106 1752
rect 14174 1748 14210 1749
rect 14068 1724 14077 1744
rect 14097 1724 14106 1744
rect 14068 1715 14106 1724
rect 14125 1741 14210 1748
rect 14125 1721 14132 1741
rect 14153 1740 14210 1741
rect 14153 1721 14182 1740
rect 14125 1720 14182 1721
rect 14202 1720 14210 1740
rect 14068 1714 14105 1715
rect 14125 1714 14210 1720
rect 14276 1744 14314 1752
rect 14387 1748 14423 1749
rect 14276 1724 14285 1744
rect 14305 1724 14314 1744
rect 14276 1715 14314 1724
rect 14338 1740 14423 1748
rect 14338 1720 14395 1740
rect 14415 1720 14423 1740
rect 14276 1714 14313 1715
rect 14338 1714 14423 1720
rect 14489 1744 14527 1752
rect 14822 1744 14859 1745
rect 15125 1744 15162 1814
rect 15187 1834 15274 1841
rect 15187 1831 15245 1834
rect 15187 1811 15192 1831
rect 15213 1814 15245 1831
rect 15265 1814 15274 1834
rect 15213 1811 15274 1814
rect 15187 1804 15274 1811
rect 15333 1834 15370 1844
rect 15333 1814 15341 1834
rect 15361 1814 15370 1834
rect 15187 1803 15218 1804
rect 14489 1724 14498 1744
rect 14518 1724 14527 1744
rect 14821 1743 15162 1744
rect 14489 1715 14527 1724
rect 14746 1738 15162 1743
rect 14746 1718 14749 1738
rect 14769 1718 15162 1738
rect 15333 1743 15370 1814
rect 15400 1843 15431 1896
rect 15738 1894 15748 1912
rect 15766 1894 15777 1912
rect 16080 1931 16713 1940
rect 17439 1931 17470 1984
rect 17500 2013 17537 2084
rect 17708 2089 18101 2109
rect 18121 2089 18124 2109
rect 17708 2084 18124 2089
rect 17708 2083 18049 2084
rect 17652 2023 17683 2024
rect 17500 1993 17509 2013
rect 17529 1993 17537 2013
rect 17500 1983 17537 1993
rect 17596 2016 17683 2023
rect 17596 2013 17657 2016
rect 17596 1993 17605 2013
rect 17625 1996 17657 2013
rect 17678 1996 17683 2016
rect 17625 1993 17683 1996
rect 17596 1986 17683 1993
rect 17708 2013 17745 2083
rect 18011 2082 18048 2083
rect 17860 2023 17896 2024
rect 17708 1993 17717 2013
rect 17737 1993 17745 2013
rect 17596 1984 17652 1986
rect 17596 1983 17633 1984
rect 17708 1983 17745 1993
rect 17804 2013 17952 2023
rect 18052 2020 18148 2022
rect 17804 1993 17813 2013
rect 17833 1993 17923 2013
rect 17943 1993 17952 2013
rect 17804 1984 17952 1993
rect 18010 2013 18148 2020
rect 18010 1993 18019 2013
rect 18039 1993 18148 2013
rect 18010 1984 18148 1993
rect 17804 1983 17841 1984
rect 17860 1932 17896 1984
rect 17915 1983 17952 1984
rect 18011 1983 18048 1984
rect 16080 1913 16090 1931
rect 16108 1930 16713 1931
rect 17331 1930 17372 1931
rect 16108 1925 16129 1930
rect 16108 1913 16120 1925
rect 17223 1923 17372 1930
rect 16080 1905 16120 1913
rect 16163 1912 16189 1913
rect 16080 1903 16117 1905
rect 16163 1894 16717 1912
rect 17223 1903 17341 1923
rect 17361 1903 17372 1923
rect 17223 1895 17372 1903
rect 17439 1927 17798 1931
rect 17439 1922 17761 1927
rect 17439 1898 17552 1922
rect 17576 1903 17761 1922
rect 17785 1903 17798 1927
rect 17576 1898 17798 1903
rect 17439 1895 17798 1898
rect 17860 1895 17895 1932
rect 17963 1929 18063 1932
rect 17963 1925 18030 1929
rect 17963 1899 17975 1925
rect 18001 1903 18030 1925
rect 18056 1903 18063 1929
rect 18001 1899 18063 1903
rect 17963 1895 18063 1899
rect 15738 1885 15775 1894
rect 15450 1843 15487 1844
rect 15400 1834 15487 1843
rect 15400 1814 15458 1834
rect 15478 1814 15487 1834
rect 15400 1804 15487 1814
rect 15546 1834 15583 1844
rect 15546 1814 15554 1834
rect 15574 1814 15583 1834
rect 16083 1835 16120 1841
rect 16163 1835 16189 1894
rect 16696 1875 16717 1894
rect 16083 1832 16189 1835
rect 15741 1819 15778 1823
rect 15400 1803 15431 1804
rect 15546 1743 15583 1814
rect 15333 1719 15583 1743
rect 15739 1813 15778 1819
rect 15739 1795 15750 1813
rect 15768 1795 15778 1813
rect 16083 1814 16092 1832
rect 16110 1818 16189 1832
rect 16274 1850 16524 1874
rect 16110 1816 16186 1818
rect 16110 1814 16120 1816
rect 16083 1804 16120 1814
rect 15739 1786 15778 1795
rect 14489 1714 14526 1715
rect 13912 1693 13948 1714
rect 14338 1693 14369 1714
rect 15125 1695 15162 1718
rect 15739 1708 15774 1786
rect 16088 1739 16119 1804
rect 16274 1779 16311 1850
rect 16426 1789 16457 1790
rect 16274 1759 16283 1779
rect 16303 1759 16311 1779
rect 16274 1749 16311 1759
rect 16370 1779 16457 1789
rect 16370 1759 16379 1779
rect 16399 1759 16457 1779
rect 16370 1750 16457 1759
rect 16370 1749 16407 1750
rect 15736 1698 15774 1708
rect 16087 1730 16124 1739
rect 16087 1712 16097 1730
rect 16115 1712 16124 1730
rect 16087 1702 16124 1712
rect 15125 1694 15295 1695
rect 15736 1694 15746 1698
rect 13745 1689 13845 1693
rect 13745 1685 13807 1689
rect 13745 1659 13752 1685
rect 13778 1663 13807 1685
rect 13833 1663 13845 1689
rect 13778 1659 13845 1663
rect 13745 1656 13845 1659
rect 13913 1656 13948 1693
rect 14010 1690 14369 1693
rect 14010 1685 14232 1690
rect 14010 1661 14023 1685
rect 14047 1666 14232 1685
rect 14256 1666 14369 1690
rect 14047 1661 14369 1666
rect 14010 1657 14369 1661
rect 14436 1685 14585 1693
rect 14436 1665 14447 1685
rect 14467 1665 14585 1685
rect 15125 1680 15746 1694
rect 15764 1680 15774 1698
rect 16426 1697 16457 1750
rect 16487 1779 16524 1850
rect 16695 1855 17088 1875
rect 17108 1855 17111 1875
rect 17439 1874 17470 1895
rect 17860 1874 17896 1895
rect 17282 1873 17319 1874
rect 16695 1850 17111 1855
rect 17281 1864 17319 1873
rect 16695 1849 17036 1850
rect 16639 1789 16670 1790
rect 16487 1759 16496 1779
rect 16516 1759 16524 1779
rect 16487 1749 16524 1759
rect 16583 1782 16670 1789
rect 16583 1779 16644 1782
rect 16583 1759 16592 1779
rect 16612 1762 16644 1779
rect 16665 1762 16670 1782
rect 16612 1759 16670 1762
rect 16583 1752 16670 1759
rect 16695 1779 16732 1849
rect 16998 1848 17035 1849
rect 17281 1844 17290 1864
rect 17310 1844 17319 1864
rect 17281 1836 17319 1844
rect 17385 1868 17470 1874
rect 17495 1873 17532 1874
rect 17385 1848 17393 1868
rect 17413 1848 17470 1868
rect 17385 1840 17470 1848
rect 17494 1864 17532 1873
rect 17494 1844 17503 1864
rect 17523 1844 17532 1864
rect 17385 1839 17421 1840
rect 17494 1836 17532 1844
rect 17598 1868 17683 1874
rect 17703 1873 17740 1874
rect 17598 1848 17606 1868
rect 17626 1867 17683 1868
rect 17626 1848 17655 1867
rect 17598 1847 17655 1848
rect 17676 1847 17683 1867
rect 17598 1840 17683 1847
rect 17702 1864 17740 1873
rect 17702 1844 17711 1864
rect 17731 1844 17740 1864
rect 17598 1839 17634 1840
rect 17702 1836 17740 1844
rect 17806 1868 17950 1874
rect 17806 1848 17814 1868
rect 17834 1848 17866 1868
rect 17890 1848 17922 1868
rect 17942 1848 17950 1868
rect 17806 1840 17950 1848
rect 17806 1839 17842 1840
rect 17914 1839 17950 1840
rect 18016 1873 18053 1874
rect 18016 1872 18054 1873
rect 18016 1864 18080 1872
rect 18016 1844 18025 1864
rect 18045 1850 18080 1864
rect 18100 1850 18103 1870
rect 18045 1845 18103 1850
rect 18045 1844 18080 1845
rect 17282 1807 17319 1836
rect 17283 1805 17319 1807
rect 17495 1805 17532 1836
rect 16847 1789 16883 1790
rect 16695 1759 16704 1779
rect 16724 1759 16732 1779
rect 16583 1750 16639 1752
rect 16583 1749 16620 1750
rect 16695 1749 16732 1759
rect 16791 1779 16939 1789
rect 17039 1786 17135 1788
rect 16791 1759 16800 1779
rect 16820 1759 16910 1779
rect 16930 1759 16939 1779
rect 16791 1750 16939 1759
rect 16997 1779 17135 1786
rect 17283 1783 17532 1805
rect 17703 1804 17740 1836
rect 18016 1832 18080 1844
rect 18120 1806 18147 1984
rect 17979 1804 18147 1806
rect 17703 1800 18147 1804
rect 16997 1759 17006 1779
rect 17026 1759 17135 1779
rect 17703 1781 17752 1800
rect 17772 1781 18147 1800
rect 17703 1778 18147 1781
rect 17979 1777 18147 1778
rect 16997 1750 17135 1759
rect 16791 1749 16828 1750
rect 16847 1698 16883 1750
rect 16902 1749 16939 1750
rect 16998 1749 17035 1750
rect 16318 1696 16359 1697
rect 15125 1674 15774 1680
rect 16210 1689 16359 1696
rect 15125 1673 15773 1674
rect 15736 1671 15773 1673
rect 14436 1658 14585 1665
rect 16210 1669 16328 1689
rect 16348 1669 16359 1689
rect 16210 1661 16359 1669
rect 16426 1693 16785 1697
rect 16426 1688 16748 1693
rect 16426 1664 16539 1688
rect 16563 1669 16748 1688
rect 16772 1669 16785 1693
rect 16563 1664 16785 1669
rect 16426 1661 16785 1664
rect 16847 1661 16882 1698
rect 16950 1695 17050 1698
rect 16950 1691 17017 1695
rect 16950 1665 16962 1691
rect 16988 1669 17017 1691
rect 17043 1669 17050 1695
rect 16988 1665 17050 1669
rect 16950 1661 17050 1665
rect 14436 1657 14477 1658
rect 13760 1604 13797 1605
rect 13856 1604 13893 1605
rect 13912 1604 13948 1656
rect 13967 1604 14004 1605
rect 13660 1595 13798 1604
rect 13660 1575 13769 1595
rect 13789 1575 13798 1595
rect 13660 1568 13798 1575
rect 13856 1595 14004 1604
rect 13856 1575 13865 1595
rect 13885 1575 13975 1595
rect 13995 1575 14004 1595
rect 13660 1566 13756 1568
rect 13856 1565 14004 1575
rect 14063 1595 14100 1605
rect 14175 1604 14212 1605
rect 14156 1602 14212 1604
rect 14063 1575 14071 1595
rect 14091 1575 14100 1595
rect 13912 1564 13948 1565
rect 13760 1505 13797 1506
rect 14063 1505 14100 1575
rect 14125 1595 14212 1602
rect 14125 1592 14183 1595
rect 14125 1572 14130 1592
rect 14151 1575 14183 1592
rect 14203 1575 14212 1595
rect 14151 1572 14212 1575
rect 14125 1565 14212 1572
rect 14271 1595 14308 1605
rect 14271 1575 14279 1595
rect 14299 1575 14308 1595
rect 14125 1564 14156 1565
rect 13759 1504 14100 1505
rect 13684 1499 14100 1504
rect 13684 1479 13687 1499
rect 13707 1479 14100 1499
rect 14271 1504 14308 1575
rect 14338 1604 14369 1657
rect 16426 1640 16457 1661
rect 16847 1640 16883 1661
rect 16090 1631 16127 1640
rect 16269 1639 16306 1640
rect 16090 1613 16099 1631
rect 16117 1613 16127 1631
rect 14388 1604 14425 1605
rect 14338 1595 14425 1604
rect 14338 1575 14396 1595
rect 14416 1575 14425 1595
rect 14338 1565 14425 1575
rect 14484 1595 14521 1605
rect 14484 1575 14492 1595
rect 14512 1575 14521 1595
rect 14338 1564 14369 1565
rect 14484 1504 14521 1575
rect 15739 1599 15776 1609
rect 16090 1603 16127 1613
rect 15739 1581 15748 1599
rect 15766 1581 15776 1599
rect 15739 1572 15776 1581
rect 15739 1548 15774 1572
rect 16091 1568 16127 1603
rect 16268 1630 16306 1639
rect 16268 1610 16277 1630
rect 16297 1610 16306 1630
rect 16268 1602 16306 1610
rect 16372 1634 16457 1640
rect 16482 1639 16519 1640
rect 16372 1614 16380 1634
rect 16400 1614 16457 1634
rect 16372 1606 16457 1614
rect 16481 1630 16519 1639
rect 16481 1610 16490 1630
rect 16510 1610 16519 1630
rect 16372 1605 16408 1606
rect 16481 1602 16519 1610
rect 16585 1634 16670 1640
rect 16690 1639 16727 1640
rect 16585 1614 16593 1634
rect 16613 1633 16670 1634
rect 16613 1614 16642 1633
rect 16585 1613 16642 1614
rect 16663 1613 16670 1633
rect 16585 1606 16670 1613
rect 16689 1630 16727 1639
rect 16689 1610 16698 1630
rect 16718 1610 16727 1630
rect 16585 1605 16621 1606
rect 16689 1602 16727 1610
rect 16793 1634 16937 1640
rect 16793 1614 16801 1634
rect 16821 1633 16909 1634
rect 16821 1614 16849 1633
rect 16793 1612 16849 1614
rect 16871 1614 16909 1633
rect 16929 1614 16937 1634
rect 16871 1612 16937 1614
rect 16793 1606 16937 1612
rect 16793 1605 16829 1606
rect 16901 1605 16937 1606
rect 17003 1639 17040 1640
rect 17003 1638 17041 1639
rect 17003 1630 17067 1638
rect 17003 1610 17012 1630
rect 17032 1616 17067 1630
rect 17087 1616 17090 1636
rect 17032 1611 17090 1616
rect 17032 1610 17067 1611
rect 16269 1573 16306 1602
rect 15737 1524 15774 1548
rect 15736 1518 15774 1524
rect 14271 1480 14521 1504
rect 15147 1500 15774 1518
rect 14729 1483 14897 1484
rect 15148 1483 15172 1500
rect 14729 1457 15173 1483
rect 14729 1455 14897 1457
rect 14729 1277 14756 1455
rect 14796 1417 14860 1429
rect 15136 1425 15173 1457
rect 15344 1456 15593 1478
rect 15344 1425 15381 1456
rect 15557 1454 15593 1456
rect 15736 1459 15774 1500
rect 16089 1527 16127 1568
rect 16270 1571 16306 1573
rect 16482 1571 16519 1602
rect 16270 1549 16519 1571
rect 16690 1570 16727 1602
rect 17003 1598 17067 1610
rect 17107 1572 17134 1750
rect 16966 1570 17134 1572
rect 16690 1544 17134 1570
rect 16691 1527 16715 1544
rect 16966 1543 17134 1544
rect 16089 1509 16716 1527
rect 17342 1523 17592 1547
rect 16089 1503 16127 1509
rect 16089 1479 16126 1503
rect 15557 1425 15594 1454
rect 14796 1416 14831 1417
rect 14773 1411 14831 1416
rect 14773 1391 14776 1411
rect 14796 1397 14831 1411
rect 14851 1397 14860 1417
rect 14796 1389 14860 1397
rect 14822 1388 14860 1389
rect 14823 1387 14860 1388
rect 14926 1421 14962 1422
rect 15034 1421 15070 1422
rect 14926 1415 15070 1421
rect 14926 1413 14992 1415
rect 14926 1393 14934 1413
rect 14954 1394 14992 1413
rect 15014 1413 15070 1415
rect 15014 1394 15042 1413
rect 14954 1393 15042 1394
rect 15062 1393 15070 1413
rect 14926 1387 15070 1393
rect 15136 1417 15174 1425
rect 15242 1421 15278 1422
rect 15136 1397 15145 1417
rect 15165 1397 15174 1417
rect 15136 1388 15174 1397
rect 15193 1414 15278 1421
rect 15193 1394 15200 1414
rect 15221 1413 15278 1414
rect 15221 1394 15250 1413
rect 15193 1393 15250 1394
rect 15270 1393 15278 1413
rect 15136 1387 15173 1388
rect 15193 1387 15278 1393
rect 15344 1417 15382 1425
rect 15455 1421 15491 1422
rect 15344 1397 15353 1417
rect 15373 1397 15382 1417
rect 15344 1388 15382 1397
rect 15406 1413 15491 1421
rect 15406 1393 15463 1413
rect 15483 1393 15491 1413
rect 15344 1387 15381 1388
rect 15406 1387 15491 1393
rect 15557 1417 15595 1425
rect 15557 1397 15566 1417
rect 15586 1397 15595 1417
rect 15557 1388 15595 1397
rect 15736 1424 15772 1459
rect 16089 1455 16124 1479
rect 16087 1446 16124 1455
rect 16087 1428 16097 1446
rect 16115 1428 16124 1446
rect 15736 1414 15773 1424
rect 16087 1418 16124 1428
rect 17342 1452 17379 1523
rect 17494 1462 17525 1463
rect 17342 1432 17351 1452
rect 17371 1432 17379 1452
rect 17342 1422 17379 1432
rect 17438 1452 17525 1462
rect 17438 1432 17447 1452
rect 17467 1432 17525 1452
rect 17438 1423 17525 1432
rect 17438 1422 17475 1423
rect 15736 1396 15746 1414
rect 15764 1396 15773 1414
rect 15557 1387 15594 1388
rect 15736 1387 15773 1396
rect 14980 1366 15016 1387
rect 15406 1366 15437 1387
rect 17494 1370 17525 1423
rect 17555 1452 17592 1523
rect 17763 1528 18156 1548
rect 18176 1528 18179 1548
rect 17763 1523 18179 1528
rect 17763 1522 18104 1523
rect 17707 1462 17738 1463
rect 17555 1432 17564 1452
rect 17584 1432 17592 1452
rect 17555 1422 17592 1432
rect 17651 1455 17738 1462
rect 17651 1452 17712 1455
rect 17651 1432 17660 1452
rect 17680 1435 17712 1452
rect 17733 1435 17738 1455
rect 17680 1432 17738 1435
rect 17651 1425 17738 1432
rect 17763 1452 17800 1522
rect 18066 1521 18103 1522
rect 17915 1462 17951 1463
rect 17763 1432 17772 1452
rect 17792 1432 17800 1452
rect 17651 1423 17707 1425
rect 17651 1422 17688 1423
rect 17763 1422 17800 1432
rect 17859 1452 18007 1462
rect 18107 1459 18203 1461
rect 17859 1432 17868 1452
rect 17888 1432 17978 1452
rect 17998 1432 18007 1452
rect 17859 1423 18007 1432
rect 18065 1452 18203 1459
rect 18065 1432 18074 1452
rect 18094 1432 18203 1452
rect 18065 1423 18203 1432
rect 17859 1422 17896 1423
rect 17915 1371 17951 1423
rect 17970 1422 18007 1423
rect 18066 1422 18103 1423
rect 17386 1369 17427 1370
rect 14813 1362 14913 1366
rect 14813 1358 14875 1362
rect 14813 1332 14820 1358
rect 14846 1336 14875 1358
rect 14901 1336 14913 1362
rect 14846 1332 14913 1336
rect 14813 1329 14913 1332
rect 14981 1329 15016 1366
rect 15078 1363 15437 1366
rect 15078 1358 15300 1363
rect 15078 1334 15091 1358
rect 15115 1339 15300 1358
rect 15324 1339 15437 1363
rect 15115 1334 15437 1339
rect 15078 1330 15437 1334
rect 15504 1358 15653 1366
rect 15504 1338 15515 1358
rect 15535 1338 15653 1358
rect 17278 1362 17427 1369
rect 16090 1354 16127 1356
rect 16090 1353 16738 1354
rect 15504 1331 15653 1338
rect 16089 1347 16738 1353
rect 15504 1330 15545 1331
rect 14828 1277 14865 1278
rect 14924 1277 14961 1278
rect 14980 1277 15016 1329
rect 15035 1277 15072 1278
rect 14728 1268 14866 1277
rect 12984 1259 13016 1264
rect 11764 1241 11860 1243
rect 11516 1214 11525 1234
rect 11545 1214 11635 1234
rect 11655 1214 11664 1234
rect 11516 1205 11664 1214
rect 11722 1234 11860 1241
rect 12477 1238 12923 1253
rect 12753 1237 12923 1238
rect 11722 1214 11731 1234
rect 11751 1214 11860 1234
rect 11722 1205 11860 1214
rect 11516 1204 11553 1205
rect 11572 1153 11608 1205
rect 11627 1204 11664 1205
rect 11723 1204 11760 1205
rect 11043 1151 11084 1152
rect 10366 1093 10403 1095
rect 10294 1085 10320 1086
rect 10363 1085 10403 1093
rect 9111 1068 9260 1075
rect 10363 1073 10375 1085
rect 10354 1068 10375 1073
rect 9111 1067 9152 1068
rect 9770 1067 10375 1068
rect 10393 1067 10403 1085
rect 8435 1014 8472 1015
rect 8531 1014 8568 1015
rect 8587 1014 8623 1066
rect 8642 1014 8679 1015
rect 8335 1005 8473 1014
rect 8335 985 8444 1005
rect 8464 985 8473 1005
rect 8335 978 8473 985
rect 8531 1005 8679 1014
rect 8531 985 8540 1005
rect 8560 985 8650 1005
rect 8670 985 8679 1005
rect 8335 976 8431 978
rect 8531 975 8679 985
rect 8738 1005 8775 1015
rect 8850 1014 8887 1015
rect 8831 1012 8887 1014
rect 8738 985 8746 1005
rect 8766 985 8775 1005
rect 8587 974 8623 975
rect 8435 915 8472 916
rect 8738 915 8775 985
rect 8800 1005 8887 1012
rect 8800 1002 8858 1005
rect 8800 982 8805 1002
rect 8826 985 8858 1002
rect 8878 985 8887 1005
rect 8826 982 8887 985
rect 8800 975 8887 982
rect 8946 1005 8983 1015
rect 8946 985 8954 1005
rect 8974 985 8983 1005
rect 8800 974 8831 975
rect 8434 914 8775 915
rect 8359 909 8775 914
rect 8359 889 8362 909
rect 8382 889 8775 909
rect 8946 914 8983 985
rect 9013 1014 9044 1067
rect 9770 1058 10403 1067
rect 9770 1051 10402 1058
rect 9770 1049 9832 1051
rect 9348 1039 9516 1040
rect 9770 1039 9792 1049
rect 9063 1014 9100 1015
rect 9013 1005 9100 1014
rect 9013 985 9071 1005
rect 9091 985 9100 1005
rect 9013 975 9100 985
rect 9159 1005 9196 1015
rect 9159 985 9167 1005
rect 9187 985 9196 1005
rect 9013 974 9044 975
rect 9159 914 9196 985
rect 8946 890 9196 914
rect 9348 1013 9792 1039
rect 9348 1011 9516 1013
rect 9348 833 9375 1011
rect 9415 973 9479 985
rect 9755 981 9792 1013
rect 9963 1012 10212 1034
rect 9963 981 10000 1012
rect 10176 1010 10212 1012
rect 10176 981 10213 1010
rect 9415 972 9450 973
rect 9392 967 9450 972
rect 9392 947 9395 967
rect 9415 953 9450 967
rect 9470 953 9479 973
rect 9415 945 9479 953
rect 9441 944 9479 945
rect 9442 943 9479 944
rect 9545 977 9581 978
rect 9653 977 9689 978
rect 9545 969 9689 977
rect 9545 949 9553 969
rect 9573 949 9602 969
rect 9545 948 9602 949
rect 9624 949 9661 969
rect 9681 949 9689 969
rect 9624 948 9689 949
rect 9545 943 9689 948
rect 9755 973 9793 981
rect 9861 977 9897 978
rect 9755 953 9764 973
rect 9784 953 9793 973
rect 9755 944 9793 953
rect 9812 970 9897 977
rect 9812 950 9819 970
rect 9840 969 9897 970
rect 9840 950 9869 969
rect 9812 949 9869 950
rect 9889 949 9897 969
rect 9755 943 9792 944
rect 9812 943 9897 949
rect 9963 973 10001 981
rect 10074 977 10110 978
rect 9963 953 9972 973
rect 9992 953 10001 973
rect 9963 944 10001 953
rect 10025 969 10110 977
rect 10025 949 10082 969
rect 10102 949 10110 969
rect 9963 943 10000 944
rect 10025 943 10110 949
rect 10176 973 10214 981
rect 10176 953 10185 973
rect 10205 953 10214 973
rect 10176 944 10214 953
rect 10176 943 10213 944
rect 9599 922 9635 943
rect 10025 922 10056 943
rect 9432 918 9532 922
rect 9432 914 9494 918
rect 9432 888 9439 914
rect 9465 892 9494 914
rect 9520 892 9532 918
rect 9465 888 9532 892
rect 9432 885 9532 888
rect 9600 885 9635 922
rect 9697 919 10056 922
rect 9697 914 9919 919
rect 9697 890 9710 914
rect 9734 895 9919 914
rect 9943 895 10056 919
rect 9734 890 10056 895
rect 9697 886 10056 890
rect 10123 914 10272 922
rect 10123 894 10134 914
rect 10154 894 10272 914
rect 10123 887 10272 894
rect 10363 902 10402 1051
rect 10805 987 10844 1136
rect 10935 1144 11084 1151
rect 10935 1124 11053 1144
rect 11073 1124 11084 1144
rect 10935 1116 11084 1124
rect 11151 1148 11510 1152
rect 11151 1143 11473 1148
rect 11151 1119 11264 1143
rect 11288 1124 11473 1143
rect 11497 1124 11510 1148
rect 11288 1119 11510 1124
rect 11151 1116 11510 1119
rect 11572 1116 11607 1153
rect 11675 1150 11775 1153
rect 11675 1146 11742 1150
rect 11675 1120 11687 1146
rect 11713 1124 11742 1146
rect 11768 1124 11775 1150
rect 11713 1120 11775 1124
rect 11675 1116 11775 1120
rect 11151 1095 11182 1116
rect 11572 1095 11608 1116
rect 10994 1094 11031 1095
rect 10993 1085 11031 1094
rect 10993 1065 11002 1085
rect 11022 1065 11031 1085
rect 10993 1057 11031 1065
rect 11097 1089 11182 1095
rect 11207 1094 11244 1095
rect 11097 1069 11105 1089
rect 11125 1069 11182 1089
rect 11097 1061 11182 1069
rect 11206 1085 11244 1094
rect 11206 1065 11215 1085
rect 11235 1065 11244 1085
rect 11097 1060 11133 1061
rect 11206 1057 11244 1065
rect 11310 1089 11395 1095
rect 11415 1094 11452 1095
rect 11310 1069 11318 1089
rect 11338 1088 11395 1089
rect 11338 1069 11367 1088
rect 11310 1068 11367 1069
rect 11388 1068 11395 1088
rect 11310 1061 11395 1068
rect 11414 1085 11452 1094
rect 11414 1065 11423 1085
rect 11443 1065 11452 1085
rect 11310 1060 11346 1061
rect 11414 1057 11452 1065
rect 11518 1090 11662 1095
rect 11518 1089 11583 1090
rect 11518 1069 11526 1089
rect 11546 1069 11583 1089
rect 11605 1089 11662 1090
rect 11605 1069 11634 1089
rect 11654 1069 11662 1089
rect 11518 1061 11662 1069
rect 11518 1060 11554 1061
rect 11626 1060 11662 1061
rect 11728 1094 11765 1095
rect 11728 1093 11766 1094
rect 11728 1085 11792 1093
rect 11728 1065 11737 1085
rect 11757 1071 11792 1085
rect 11812 1071 11815 1091
rect 11757 1066 11815 1071
rect 11757 1065 11792 1066
rect 10994 1028 11031 1057
rect 10995 1026 11031 1028
rect 11207 1026 11244 1057
rect 10995 1004 11244 1026
rect 11415 1025 11452 1057
rect 11728 1053 11792 1065
rect 11832 1027 11859 1205
rect 11691 1025 11859 1027
rect 11415 999 11859 1025
rect 12011 1124 12261 1148
rect 12011 1053 12048 1124
rect 12163 1063 12194 1064
rect 12011 1033 12020 1053
rect 12040 1033 12048 1053
rect 12011 1023 12048 1033
rect 12107 1053 12194 1063
rect 12107 1033 12116 1053
rect 12136 1033 12194 1053
rect 12107 1024 12194 1033
rect 12107 1023 12144 1024
rect 11415 989 11437 999
rect 11691 998 11859 999
rect 11375 987 11437 989
rect 10805 980 11437 987
rect 10804 971 11437 980
rect 12163 971 12194 1024
rect 12224 1053 12261 1124
rect 12432 1129 12825 1149
rect 12845 1129 12848 1149
rect 12432 1124 12848 1129
rect 12432 1123 12773 1124
rect 12376 1063 12407 1064
rect 12224 1033 12233 1053
rect 12253 1033 12261 1053
rect 12224 1023 12261 1033
rect 12320 1056 12407 1063
rect 12320 1053 12381 1056
rect 12320 1033 12329 1053
rect 12349 1036 12381 1053
rect 12402 1036 12407 1056
rect 12349 1033 12407 1036
rect 12320 1026 12407 1033
rect 12432 1053 12469 1123
rect 12735 1122 12772 1123
rect 12584 1063 12620 1064
rect 12432 1033 12441 1053
rect 12461 1033 12469 1053
rect 12320 1024 12376 1026
rect 12320 1023 12357 1024
rect 12432 1023 12469 1033
rect 12528 1053 12676 1063
rect 12776 1060 12872 1062
rect 12528 1033 12537 1053
rect 12557 1033 12647 1053
rect 12667 1033 12676 1053
rect 12528 1024 12676 1033
rect 12734 1053 12872 1060
rect 12734 1033 12743 1053
rect 12763 1033 12872 1053
rect 12734 1024 12872 1033
rect 12528 1023 12565 1024
rect 12584 972 12620 1024
rect 12639 1023 12676 1024
rect 12735 1023 12772 1024
rect 10804 953 10814 971
rect 10832 970 11437 971
rect 12055 970 12096 971
rect 10832 965 10853 970
rect 10832 953 10844 965
rect 11947 963 12096 970
rect 10804 945 10844 953
rect 10887 952 10913 953
rect 10804 943 10841 945
rect 10123 886 10164 887
rect 9447 833 9484 834
rect 9543 833 9580 834
rect 9599 833 9635 885
rect 9654 833 9691 834
rect 7512 788 7517 814
rect 7536 788 7543 814
rect 9347 824 9485 833
rect 9347 804 9456 824
rect 9476 804 9485 824
rect 9347 797 9485 804
rect 9543 824 9691 833
rect 9543 804 9552 824
rect 9572 804 9662 824
rect 9682 804 9691 824
rect 9347 795 9443 797
rect 9543 794 9691 804
rect 9750 824 9787 834
rect 9862 833 9899 834
rect 9843 831 9899 833
rect 9750 804 9758 824
rect 9778 804 9787 824
rect 9599 793 9635 794
rect 7512 785 7543 788
rect 6341 761 6479 770
rect 6135 760 6172 761
rect 6191 709 6227 761
rect 6246 760 6283 761
rect 6342 760 6379 761
rect 5662 707 5703 708
rect 4469 685 5118 691
rect 5554 700 5703 707
rect 4469 684 5117 685
rect 5080 682 5117 684
rect 5554 680 5672 700
rect 5692 680 5703 700
rect 5554 672 5703 680
rect 5770 704 6129 708
rect 5770 699 6092 704
rect 5770 675 5883 699
rect 5907 680 6092 699
rect 6116 680 6129 704
rect 5907 675 6129 680
rect 5770 672 6129 675
rect 6191 672 6226 709
rect 6294 706 6394 709
rect 6294 702 6361 706
rect 6294 676 6306 702
rect 6332 680 6361 702
rect 6387 680 6394 706
rect 6332 676 6394 680
rect 6294 672 6394 676
rect 5770 651 5801 672
rect 6191 651 6227 672
rect 5434 642 5471 651
rect 5613 650 5650 651
rect 5434 624 5443 642
rect 5461 624 5471 642
rect 5083 618 5120 620
rect 1029 602 1197 604
rect 753 576 1197 602
rect 754 550 778 576
rect 1029 575 1197 576
rect 5078 610 5120 618
rect 5434 614 5471 624
rect 5078 592 5092 610
rect 5110 592 5120 610
rect 5078 583 5120 592
rect 747 542 787 550
rect 747 535 756 542
rect 152 520 756 535
rect 779 520 787 542
rect 152 517 787 520
rect 152 511 190 517
rect 747 505 787 517
rect 5078 542 5119 583
rect 5435 579 5471 614
rect 5612 641 5650 650
rect 5612 621 5621 641
rect 5641 621 5650 641
rect 5612 613 5650 621
rect 5716 645 5801 651
rect 5826 650 5863 651
rect 5716 625 5724 645
rect 5744 625 5801 645
rect 5716 617 5801 625
rect 5825 641 5863 650
rect 5825 621 5834 641
rect 5854 621 5863 641
rect 5716 616 5752 617
rect 5825 613 5863 621
rect 5929 645 6014 651
rect 6034 650 6071 651
rect 5929 625 5937 645
rect 5957 644 6014 645
rect 5957 625 5986 644
rect 5929 624 5986 625
rect 6007 624 6014 644
rect 5929 617 6014 624
rect 6033 641 6071 650
rect 6033 621 6042 641
rect 6062 621 6071 641
rect 5929 616 5965 617
rect 6033 613 6071 621
rect 6137 645 6281 651
rect 6137 625 6145 645
rect 6165 644 6253 645
rect 6165 625 6193 644
rect 6137 623 6193 625
rect 6215 625 6253 644
rect 6273 625 6281 645
rect 6215 623 6281 625
rect 6137 617 6281 623
rect 6137 616 6173 617
rect 6245 616 6281 617
rect 6347 650 6384 651
rect 6347 649 6385 650
rect 6347 641 6411 649
rect 6347 621 6356 641
rect 6376 627 6411 641
rect 6431 627 6434 647
rect 6376 622 6434 627
rect 6376 621 6411 622
rect 5613 584 5650 613
rect 5078 520 5089 542
rect 5112 520 5119 542
rect 5078 515 5119 520
rect 5433 514 5471 579
rect 5614 582 5650 584
rect 5826 582 5863 613
rect 5614 560 5863 582
rect 6034 581 6071 613
rect 6347 609 6411 621
rect 6451 583 6478 761
rect 9447 734 9484 735
rect 9750 734 9787 804
rect 9812 824 9899 831
rect 9812 821 9870 824
rect 9812 801 9817 821
rect 9838 804 9870 821
rect 9890 804 9899 824
rect 9838 801 9899 804
rect 9812 794 9899 801
rect 9958 824 9995 834
rect 9958 804 9966 824
rect 9986 804 9995 824
rect 9812 793 9843 794
rect 9446 733 9787 734
rect 9371 728 9787 733
rect 9371 708 9374 728
rect 9394 708 9787 728
rect 9958 733 9995 804
rect 10025 833 10056 886
rect 10363 884 10373 902
rect 10391 884 10402 902
rect 10887 934 11441 952
rect 11947 943 12065 963
rect 12085 943 12096 963
rect 11947 935 12096 943
rect 12163 967 12522 971
rect 12163 962 12485 967
rect 12163 938 12276 962
rect 12300 943 12485 962
rect 12509 943 12522 967
rect 12300 938 12522 943
rect 12163 935 12522 938
rect 12584 935 12619 972
rect 12687 969 12787 972
rect 12687 965 12754 969
rect 12687 939 12699 965
rect 12725 943 12754 965
rect 12780 943 12787 969
rect 12725 939 12787 943
rect 12687 935 12787 939
rect 10363 875 10400 884
rect 10807 875 10844 881
rect 10887 875 10913 934
rect 11420 915 11441 934
rect 10807 872 10913 875
rect 10807 854 10816 872
rect 10834 858 10913 872
rect 10998 890 11248 914
rect 10834 856 10910 858
rect 10834 854 10844 856
rect 10807 844 10844 854
rect 10075 833 10112 834
rect 10025 824 10112 833
rect 10025 804 10083 824
rect 10103 804 10112 824
rect 10025 794 10112 804
rect 10171 824 10208 834
rect 10171 804 10179 824
rect 10199 804 10208 824
rect 10366 809 10403 813
rect 10025 793 10056 794
rect 10171 733 10208 804
rect 9958 709 10208 733
rect 10364 803 10403 809
rect 10364 785 10375 803
rect 10393 785 10403 803
rect 10364 776 10403 785
rect 10812 779 10843 844
rect 10998 819 11035 890
rect 11150 829 11181 830
rect 10998 799 11007 819
rect 11027 799 11035 819
rect 10998 789 11035 799
rect 11094 819 11181 829
rect 11094 799 11103 819
rect 11123 799 11181 819
rect 11094 790 11181 799
rect 11094 789 11131 790
rect 9750 685 9787 708
rect 10364 698 10399 776
rect 10811 770 10848 779
rect 10811 752 10821 770
rect 10839 752 10848 770
rect 10811 742 10848 752
rect 11150 737 11181 790
rect 11211 819 11248 890
rect 11419 895 11812 915
rect 11832 895 11835 915
rect 12163 914 12194 935
rect 12584 914 12620 935
rect 12006 913 12043 914
rect 11419 890 11835 895
rect 12005 904 12043 913
rect 11419 889 11760 890
rect 11363 829 11394 830
rect 11211 799 11220 819
rect 11240 799 11248 819
rect 11211 789 11248 799
rect 11307 822 11394 829
rect 11307 819 11368 822
rect 11307 799 11316 819
rect 11336 802 11368 819
rect 11389 802 11394 822
rect 11336 799 11394 802
rect 11307 792 11394 799
rect 11419 819 11456 889
rect 11722 888 11759 889
rect 12005 884 12014 904
rect 12034 884 12043 904
rect 12005 876 12043 884
rect 12109 908 12194 914
rect 12219 913 12256 914
rect 12109 888 12117 908
rect 12137 888 12194 908
rect 12109 880 12194 888
rect 12218 904 12256 913
rect 12218 884 12227 904
rect 12247 884 12256 904
rect 12109 879 12145 880
rect 12218 876 12256 884
rect 12322 908 12407 914
rect 12427 913 12464 914
rect 12322 888 12330 908
rect 12350 907 12407 908
rect 12350 888 12379 907
rect 12322 887 12379 888
rect 12400 887 12407 907
rect 12322 880 12407 887
rect 12426 904 12464 913
rect 12426 884 12435 904
rect 12455 884 12464 904
rect 12322 879 12358 880
rect 12426 876 12464 884
rect 12530 909 12674 914
rect 12530 908 12589 909
rect 12530 888 12538 908
rect 12558 889 12589 908
rect 12613 908 12674 909
rect 12613 889 12646 908
rect 12558 888 12646 889
rect 12666 888 12674 908
rect 12530 880 12674 888
rect 12530 879 12566 880
rect 12638 879 12674 880
rect 12740 913 12777 914
rect 12740 912 12778 913
rect 12740 904 12804 912
rect 12740 884 12749 904
rect 12769 890 12804 904
rect 12824 890 12827 910
rect 12769 885 12827 890
rect 12769 884 12804 885
rect 12006 847 12043 876
rect 12007 845 12043 847
rect 12219 845 12256 876
rect 11571 829 11607 830
rect 11419 799 11428 819
rect 11448 799 11456 819
rect 11307 790 11363 792
rect 11307 789 11344 790
rect 11419 789 11456 799
rect 11515 819 11663 829
rect 11763 826 11859 828
rect 11515 799 11524 819
rect 11544 799 11634 819
rect 11654 799 11663 819
rect 11515 790 11663 799
rect 11721 819 11859 826
rect 12007 823 12256 845
rect 12427 844 12464 876
rect 12740 872 12804 884
rect 12844 846 12871 1024
rect 12703 844 12871 846
rect 12427 840 12871 844
rect 11721 799 11730 819
rect 11750 799 11859 819
rect 12427 821 12476 840
rect 12496 821 12871 840
rect 12427 818 12871 821
rect 12703 817 12871 818
rect 12892 843 12923 1237
rect 12984 1241 12989 1259
rect 13009 1241 13016 1259
rect 12984 1236 13016 1241
rect 12987 1234 13016 1236
rect 13716 1249 13884 1250
rect 13716 1246 14160 1249
rect 13716 1227 14091 1246
rect 14111 1227 14160 1246
rect 14728 1248 14837 1268
rect 14857 1248 14866 1268
rect 13716 1223 14160 1227
rect 13716 1221 13884 1223
rect 13716 1043 13743 1221
rect 13783 1183 13847 1195
rect 14123 1191 14160 1223
rect 14331 1222 14580 1244
rect 14728 1241 14866 1248
rect 14924 1268 15072 1277
rect 14924 1248 14933 1268
rect 14953 1248 15043 1268
rect 15063 1248 15072 1268
rect 14728 1239 14824 1241
rect 14924 1238 15072 1248
rect 15131 1268 15168 1278
rect 15243 1277 15280 1278
rect 15224 1275 15280 1277
rect 15131 1248 15139 1268
rect 15159 1248 15168 1268
rect 14980 1237 15016 1238
rect 14331 1191 14368 1222
rect 14544 1220 14580 1222
rect 14544 1191 14581 1220
rect 13783 1182 13818 1183
rect 13760 1177 13818 1182
rect 13760 1157 13763 1177
rect 13783 1163 13818 1177
rect 13838 1163 13847 1183
rect 13783 1155 13847 1163
rect 13809 1154 13847 1155
rect 13810 1153 13847 1154
rect 13913 1187 13949 1188
rect 14021 1187 14057 1188
rect 13913 1179 14057 1187
rect 13913 1159 13921 1179
rect 13941 1159 13973 1179
rect 13997 1159 14029 1179
rect 14049 1159 14057 1179
rect 13913 1153 14057 1159
rect 14123 1183 14161 1191
rect 14229 1187 14265 1188
rect 14123 1163 14132 1183
rect 14152 1163 14161 1183
rect 14123 1154 14161 1163
rect 14180 1180 14265 1187
rect 14180 1160 14187 1180
rect 14208 1179 14265 1180
rect 14208 1160 14237 1179
rect 14180 1159 14237 1160
rect 14257 1159 14265 1179
rect 14123 1153 14160 1154
rect 14180 1153 14265 1159
rect 14331 1183 14369 1191
rect 14442 1187 14478 1188
rect 14331 1163 14340 1183
rect 14360 1163 14369 1183
rect 14331 1154 14369 1163
rect 14393 1179 14478 1187
rect 14393 1159 14450 1179
rect 14470 1159 14478 1179
rect 14331 1153 14368 1154
rect 14393 1153 14478 1159
rect 14544 1183 14582 1191
rect 14544 1163 14553 1183
rect 14573 1163 14582 1183
rect 14828 1178 14865 1179
rect 15131 1178 15168 1248
rect 15193 1268 15280 1275
rect 15193 1265 15251 1268
rect 15193 1245 15198 1265
rect 15219 1248 15251 1265
rect 15271 1248 15280 1268
rect 15219 1245 15280 1248
rect 15193 1238 15280 1245
rect 15339 1268 15376 1278
rect 15339 1248 15347 1268
rect 15367 1248 15376 1268
rect 15193 1237 15224 1238
rect 14827 1177 15168 1178
rect 14544 1154 14582 1163
rect 14752 1172 15168 1177
rect 14544 1153 14581 1154
rect 13967 1132 14003 1153
rect 14393 1132 14424 1153
rect 14752 1152 14755 1172
rect 14775 1152 15168 1172
rect 15339 1177 15376 1248
rect 15406 1277 15437 1330
rect 16089 1329 16099 1347
rect 16117 1333 16738 1347
rect 17278 1342 17396 1362
rect 17416 1342 17427 1362
rect 17278 1334 17427 1342
rect 17494 1366 17853 1370
rect 17494 1361 17816 1366
rect 17494 1337 17607 1361
rect 17631 1342 17816 1361
rect 17840 1342 17853 1366
rect 17631 1337 17853 1342
rect 17494 1334 17853 1337
rect 17915 1334 17950 1371
rect 18018 1368 18118 1371
rect 18018 1364 18085 1368
rect 18018 1338 18030 1364
rect 18056 1342 18085 1364
rect 18111 1342 18118 1368
rect 18056 1338 18118 1342
rect 18018 1334 18118 1338
rect 16117 1329 16127 1333
rect 16568 1332 16738 1333
rect 15739 1315 15776 1325
rect 15739 1297 15748 1315
rect 15766 1297 15776 1315
rect 15739 1288 15776 1297
rect 16089 1319 16127 1329
rect 15456 1277 15493 1278
rect 15406 1268 15493 1277
rect 15406 1248 15464 1268
rect 15484 1248 15493 1268
rect 15406 1238 15493 1248
rect 15552 1268 15589 1278
rect 15552 1248 15560 1268
rect 15580 1248 15589 1268
rect 15406 1237 15437 1238
rect 15552 1177 15589 1248
rect 15744 1223 15775 1288
rect 16089 1241 16124 1319
rect 16701 1309 16738 1332
rect 17494 1313 17525 1334
rect 17915 1313 17951 1334
rect 17337 1312 17374 1313
rect 16085 1232 16124 1241
rect 15743 1213 15780 1223
rect 15743 1211 15753 1213
rect 15677 1209 15753 1211
rect 15339 1153 15589 1177
rect 15674 1195 15753 1209
rect 15771 1195 15780 1213
rect 16085 1214 16095 1232
rect 16113 1214 16124 1232
rect 16085 1208 16124 1214
rect 16280 1284 16530 1308
rect 16280 1213 16317 1284
rect 16432 1223 16463 1224
rect 16085 1204 16122 1208
rect 15674 1192 15780 1195
rect 15146 1133 15167 1152
rect 15674 1133 15700 1192
rect 15743 1186 15780 1192
rect 16280 1193 16289 1213
rect 16309 1193 16317 1213
rect 16280 1183 16317 1193
rect 16376 1213 16463 1223
rect 16376 1193 16385 1213
rect 16405 1193 16463 1213
rect 16376 1184 16463 1193
rect 16376 1183 16413 1184
rect 16088 1133 16125 1142
rect 13800 1128 13900 1132
rect 13800 1124 13862 1128
rect 13800 1098 13807 1124
rect 13833 1102 13862 1124
rect 13888 1102 13900 1128
rect 13833 1098 13900 1102
rect 13800 1095 13900 1098
rect 13968 1095 14003 1132
rect 14065 1129 14424 1132
rect 14065 1124 14287 1129
rect 14065 1100 14078 1124
rect 14102 1105 14287 1124
rect 14311 1105 14424 1129
rect 14102 1100 14424 1105
rect 14065 1096 14424 1100
rect 14491 1124 14640 1132
rect 14491 1104 14502 1124
rect 14522 1104 14640 1124
rect 15146 1115 15700 1133
rect 15746 1122 15783 1124
rect 15674 1114 15700 1115
rect 15743 1114 15783 1122
rect 14491 1097 14640 1104
rect 15743 1102 15755 1114
rect 15734 1097 15755 1102
rect 14491 1096 14532 1097
rect 15150 1096 15755 1097
rect 15773 1096 15783 1114
rect 13815 1043 13852 1044
rect 13911 1043 13948 1044
rect 13967 1043 14003 1095
rect 14022 1043 14059 1044
rect 13715 1034 13853 1043
rect 13715 1014 13824 1034
rect 13844 1014 13853 1034
rect 13715 1007 13853 1014
rect 13911 1034 14059 1043
rect 13911 1014 13920 1034
rect 13940 1014 14030 1034
rect 14050 1014 14059 1034
rect 13715 1005 13811 1007
rect 13911 1004 14059 1014
rect 14118 1034 14155 1044
rect 14230 1043 14267 1044
rect 14211 1041 14267 1043
rect 14118 1014 14126 1034
rect 14146 1014 14155 1034
rect 13967 1003 14003 1004
rect 13815 944 13852 945
rect 14118 944 14155 1014
rect 14180 1034 14267 1041
rect 14180 1031 14238 1034
rect 14180 1011 14185 1031
rect 14206 1014 14238 1031
rect 14258 1014 14267 1034
rect 14206 1011 14267 1014
rect 14180 1004 14267 1011
rect 14326 1034 14363 1044
rect 14326 1014 14334 1034
rect 14354 1014 14363 1034
rect 14180 1003 14211 1004
rect 13814 943 14155 944
rect 13739 938 14155 943
rect 13739 918 13742 938
rect 13762 918 14155 938
rect 14326 943 14363 1014
rect 14393 1043 14424 1096
rect 15150 1087 15783 1096
rect 16086 1115 16097 1133
rect 16115 1115 16125 1133
rect 16432 1131 16463 1184
rect 16493 1213 16530 1284
rect 16701 1289 17094 1309
rect 17114 1289 17117 1309
rect 16701 1284 17117 1289
rect 17336 1303 17374 1312
rect 16701 1283 17042 1284
rect 17336 1283 17345 1303
rect 17365 1283 17374 1303
rect 16645 1223 16676 1224
rect 16493 1193 16502 1213
rect 16522 1193 16530 1213
rect 16493 1183 16530 1193
rect 16589 1216 16676 1223
rect 16589 1213 16650 1216
rect 16589 1193 16598 1213
rect 16618 1196 16650 1213
rect 16671 1196 16676 1216
rect 16618 1193 16676 1196
rect 16589 1186 16676 1193
rect 16701 1213 16738 1283
rect 17004 1282 17041 1283
rect 17336 1275 17374 1283
rect 17440 1307 17525 1313
rect 17550 1312 17587 1313
rect 17440 1287 17448 1307
rect 17468 1287 17525 1307
rect 17440 1279 17525 1287
rect 17549 1303 17587 1312
rect 17549 1283 17558 1303
rect 17578 1283 17587 1303
rect 17440 1278 17476 1279
rect 17549 1275 17587 1283
rect 17653 1307 17738 1313
rect 17758 1312 17795 1313
rect 17653 1287 17661 1307
rect 17681 1306 17738 1307
rect 17681 1287 17710 1306
rect 17653 1286 17710 1287
rect 17731 1286 17738 1306
rect 17653 1279 17738 1286
rect 17757 1303 17795 1312
rect 17757 1283 17766 1303
rect 17786 1283 17795 1303
rect 17653 1278 17689 1279
rect 17757 1275 17795 1283
rect 17861 1307 18005 1313
rect 17861 1287 17869 1307
rect 17889 1306 17977 1307
rect 17889 1287 17922 1306
rect 17945 1287 17977 1306
rect 17997 1287 18005 1307
rect 17861 1279 18005 1287
rect 17861 1278 17897 1279
rect 17969 1278 18005 1279
rect 18071 1312 18108 1313
rect 18071 1311 18109 1312
rect 18071 1303 18135 1311
rect 18071 1283 18080 1303
rect 18100 1289 18135 1303
rect 18155 1289 18158 1309
rect 18100 1284 18158 1289
rect 18100 1283 18135 1284
rect 17337 1246 17374 1275
rect 17338 1244 17374 1246
rect 17550 1244 17587 1275
rect 16853 1223 16889 1224
rect 16701 1193 16710 1213
rect 16730 1193 16738 1213
rect 16589 1184 16645 1186
rect 16589 1183 16626 1184
rect 16701 1183 16738 1193
rect 16797 1213 16945 1223
rect 17338 1222 17587 1244
rect 17758 1243 17795 1275
rect 18071 1271 18135 1283
rect 18175 1245 18202 1423
rect 18034 1243 18202 1245
rect 17758 1232 18202 1243
rect 18265 1243 18295 2244
rect 18384 2237 18421 2248
rect 20005 2237 20032 2415
rect 20072 2377 20136 2389
rect 20412 2385 20449 2417
rect 20620 2416 20869 2438
rect 20620 2385 20657 2416
rect 20833 2414 20869 2416
rect 21012 2419 21050 2460
rect 20833 2385 20870 2414
rect 20072 2376 20107 2377
rect 20049 2371 20107 2376
rect 20049 2351 20052 2371
rect 20072 2357 20107 2371
rect 20127 2357 20136 2377
rect 20072 2349 20136 2357
rect 20098 2348 20136 2349
rect 20099 2347 20136 2348
rect 20202 2381 20238 2382
rect 20310 2381 20346 2382
rect 20202 2375 20346 2381
rect 20202 2373 20268 2375
rect 20202 2353 20210 2373
rect 20230 2354 20268 2373
rect 20290 2373 20346 2375
rect 20290 2354 20318 2373
rect 20230 2353 20318 2354
rect 20338 2353 20346 2373
rect 20202 2347 20346 2353
rect 20412 2377 20450 2385
rect 20518 2381 20554 2382
rect 20412 2357 20421 2377
rect 20441 2357 20450 2377
rect 20412 2348 20450 2357
rect 20469 2374 20554 2381
rect 20469 2354 20476 2374
rect 20497 2373 20554 2374
rect 20497 2354 20526 2373
rect 20469 2353 20526 2354
rect 20546 2353 20554 2373
rect 20412 2347 20449 2348
rect 20469 2347 20554 2353
rect 20620 2377 20658 2385
rect 20731 2381 20767 2382
rect 20620 2357 20629 2377
rect 20649 2357 20658 2377
rect 20620 2348 20658 2357
rect 20682 2373 20767 2381
rect 20682 2353 20739 2373
rect 20759 2353 20767 2373
rect 20620 2347 20657 2348
rect 20682 2347 20767 2353
rect 20833 2377 20871 2385
rect 20833 2357 20842 2377
rect 20862 2357 20871 2377
rect 20833 2348 20871 2357
rect 21012 2384 21048 2419
rect 21012 2374 21049 2384
rect 21012 2356 21022 2374
rect 21040 2356 21049 2374
rect 20833 2347 20870 2348
rect 21012 2347 21049 2356
rect 20256 2326 20292 2347
rect 20682 2326 20713 2347
rect 20089 2322 20189 2326
rect 20089 2318 20151 2322
rect 20089 2292 20096 2318
rect 20122 2296 20151 2318
rect 20177 2296 20189 2322
rect 20122 2292 20189 2296
rect 20089 2289 20189 2292
rect 20257 2289 20292 2326
rect 20354 2323 20713 2326
rect 20354 2318 20576 2323
rect 20354 2294 20367 2318
rect 20391 2299 20576 2318
rect 20600 2299 20713 2323
rect 20391 2294 20713 2299
rect 20354 2290 20713 2294
rect 20780 2318 20929 2326
rect 20780 2298 20791 2318
rect 20811 2298 20929 2318
rect 20780 2291 20929 2298
rect 20780 2290 20821 2291
rect 20104 2237 20141 2238
rect 20200 2237 20237 2238
rect 20256 2237 20292 2289
rect 20311 2237 20348 2238
rect 20004 2228 20142 2237
rect 18940 2210 18971 2213
rect 18940 2184 18947 2210
rect 18966 2184 18971 2210
rect 18940 1790 18971 2184
rect 18992 2209 19160 2210
rect 18992 2206 19436 2209
rect 18992 2187 19367 2206
rect 19387 2187 19436 2206
rect 20004 2208 20113 2228
rect 20133 2208 20142 2228
rect 18992 2183 19436 2187
rect 18992 2181 19160 2183
rect 18992 2003 19019 2181
rect 19059 2143 19123 2155
rect 19399 2151 19436 2183
rect 19607 2182 19856 2204
rect 20004 2201 20142 2208
rect 20200 2228 20348 2237
rect 20200 2208 20209 2228
rect 20229 2208 20319 2228
rect 20339 2208 20348 2228
rect 20004 2199 20100 2201
rect 20200 2198 20348 2208
rect 20407 2228 20444 2238
rect 20519 2237 20556 2238
rect 20500 2235 20556 2237
rect 20407 2208 20415 2228
rect 20435 2208 20444 2228
rect 20256 2197 20292 2198
rect 19607 2151 19644 2182
rect 19820 2180 19856 2182
rect 19820 2151 19857 2180
rect 19059 2142 19094 2143
rect 19036 2137 19094 2142
rect 19036 2117 19039 2137
rect 19059 2123 19094 2137
rect 19114 2123 19123 2143
rect 19059 2115 19123 2123
rect 19085 2114 19123 2115
rect 19086 2113 19123 2114
rect 19189 2147 19225 2148
rect 19297 2147 19333 2148
rect 19189 2139 19333 2147
rect 19189 2119 19197 2139
rect 19217 2138 19305 2139
rect 19217 2119 19250 2138
rect 19189 2118 19250 2119
rect 19274 2119 19305 2138
rect 19325 2119 19333 2139
rect 19274 2118 19333 2119
rect 19189 2113 19333 2118
rect 19399 2143 19437 2151
rect 19505 2147 19541 2148
rect 19399 2123 19408 2143
rect 19428 2123 19437 2143
rect 19399 2114 19437 2123
rect 19456 2140 19541 2147
rect 19456 2120 19463 2140
rect 19484 2139 19541 2140
rect 19484 2120 19513 2139
rect 19456 2119 19513 2120
rect 19533 2119 19541 2139
rect 19399 2113 19436 2114
rect 19456 2113 19541 2119
rect 19607 2143 19645 2151
rect 19718 2147 19754 2148
rect 19607 2123 19616 2143
rect 19636 2123 19645 2143
rect 19607 2114 19645 2123
rect 19669 2139 19754 2147
rect 19669 2119 19726 2139
rect 19746 2119 19754 2139
rect 19607 2113 19644 2114
rect 19669 2113 19754 2119
rect 19820 2143 19858 2151
rect 19820 2123 19829 2143
rect 19849 2123 19858 2143
rect 20104 2138 20141 2139
rect 20407 2138 20444 2208
rect 20469 2228 20556 2235
rect 20469 2225 20527 2228
rect 20469 2205 20474 2225
rect 20495 2208 20527 2225
rect 20547 2208 20556 2228
rect 20495 2205 20556 2208
rect 20469 2198 20556 2205
rect 20615 2228 20652 2238
rect 20615 2208 20623 2228
rect 20643 2208 20652 2228
rect 20469 2197 20500 2198
rect 20103 2137 20444 2138
rect 19820 2114 19858 2123
rect 20028 2132 20444 2137
rect 19820 2113 19857 2114
rect 19243 2092 19279 2113
rect 19669 2092 19700 2113
rect 20028 2112 20031 2132
rect 20051 2112 20444 2132
rect 20615 2137 20652 2208
rect 20682 2237 20713 2290
rect 21015 2275 21052 2285
rect 21015 2257 21024 2275
rect 21042 2257 21052 2275
rect 21015 2248 21052 2257
rect 20732 2237 20769 2238
rect 20682 2228 20769 2237
rect 20682 2208 20740 2228
rect 20760 2208 20769 2228
rect 20682 2198 20769 2208
rect 20828 2228 20865 2238
rect 20828 2208 20836 2228
rect 20856 2208 20865 2228
rect 20682 2197 20713 2198
rect 20828 2137 20865 2208
rect 21020 2183 21051 2248
rect 21019 2173 21056 2183
rect 21019 2171 21029 2173
rect 20953 2169 21029 2171
rect 20615 2113 20865 2137
rect 20950 2155 21029 2169
rect 21047 2155 21056 2173
rect 20950 2152 21056 2155
rect 20422 2093 20443 2112
rect 20950 2093 20976 2152
rect 21019 2146 21056 2152
rect 19076 2088 19176 2092
rect 19076 2084 19138 2088
rect 19076 2058 19083 2084
rect 19109 2062 19138 2084
rect 19164 2062 19176 2088
rect 19109 2058 19176 2062
rect 19076 2055 19176 2058
rect 19244 2055 19279 2092
rect 19341 2089 19700 2092
rect 19341 2084 19563 2089
rect 19341 2060 19354 2084
rect 19378 2065 19563 2084
rect 19587 2065 19700 2089
rect 19378 2060 19700 2065
rect 19341 2056 19700 2060
rect 19767 2084 19916 2092
rect 19767 2064 19778 2084
rect 19798 2064 19916 2084
rect 20422 2075 20976 2093
rect 21022 2082 21059 2084
rect 20950 2074 20976 2075
rect 21019 2074 21059 2082
rect 19767 2057 19916 2064
rect 21019 2062 21031 2074
rect 21010 2057 21031 2062
rect 19767 2056 19808 2057
rect 20426 2056 21031 2057
rect 21049 2056 21059 2074
rect 19091 2003 19128 2004
rect 19187 2003 19224 2004
rect 19243 2003 19279 2055
rect 19298 2003 19335 2004
rect 18991 1994 19129 2003
rect 18991 1974 19100 1994
rect 19120 1974 19129 1994
rect 18991 1967 19129 1974
rect 19187 1994 19335 2003
rect 19187 1974 19196 1994
rect 19216 1974 19306 1994
rect 19326 1974 19335 1994
rect 18991 1965 19087 1967
rect 19187 1964 19335 1974
rect 19394 1994 19431 2004
rect 19506 2003 19543 2004
rect 19487 2001 19543 2003
rect 19394 1974 19402 1994
rect 19422 1974 19431 1994
rect 19243 1963 19279 1964
rect 19091 1904 19128 1905
rect 19394 1904 19431 1974
rect 19456 1994 19543 2001
rect 19456 1991 19514 1994
rect 19456 1971 19461 1991
rect 19482 1974 19514 1991
rect 19534 1974 19543 1994
rect 19482 1971 19543 1974
rect 19456 1964 19543 1971
rect 19602 1994 19639 2004
rect 19602 1974 19610 1994
rect 19630 1974 19639 1994
rect 19456 1963 19487 1964
rect 19090 1903 19431 1904
rect 19015 1898 19431 1903
rect 19015 1878 19018 1898
rect 19038 1878 19431 1898
rect 19602 1903 19639 1974
rect 19669 2003 19700 2056
rect 20426 2047 21059 2056
rect 20426 2040 21058 2047
rect 20426 2038 20488 2040
rect 20004 2028 20172 2029
rect 20426 2028 20448 2038
rect 19719 2003 19756 2004
rect 19669 1994 19756 2003
rect 19669 1974 19727 1994
rect 19747 1974 19756 1994
rect 19669 1964 19756 1974
rect 19815 1994 19852 2004
rect 19815 1974 19823 1994
rect 19843 1974 19852 1994
rect 19669 1963 19700 1964
rect 19815 1903 19852 1974
rect 19602 1879 19852 1903
rect 20004 2002 20448 2028
rect 20004 2000 20172 2002
rect 20004 1822 20031 2000
rect 20071 1962 20135 1974
rect 20411 1970 20448 2002
rect 20619 2001 20868 2023
rect 20619 1970 20656 2001
rect 20832 1999 20868 2001
rect 20832 1970 20869 1999
rect 20071 1961 20106 1962
rect 20048 1956 20106 1961
rect 20048 1936 20051 1956
rect 20071 1942 20106 1956
rect 20126 1942 20135 1962
rect 20071 1934 20135 1942
rect 20097 1933 20135 1934
rect 20098 1932 20135 1933
rect 20201 1966 20237 1967
rect 20309 1966 20345 1967
rect 20201 1958 20345 1966
rect 20201 1938 20209 1958
rect 20229 1938 20258 1958
rect 20201 1937 20258 1938
rect 20280 1938 20317 1958
rect 20337 1938 20345 1958
rect 20280 1937 20345 1938
rect 20201 1932 20345 1937
rect 20411 1962 20449 1970
rect 20517 1966 20553 1967
rect 20411 1942 20420 1962
rect 20440 1942 20449 1962
rect 20411 1933 20449 1942
rect 20468 1959 20553 1966
rect 20468 1939 20475 1959
rect 20496 1958 20553 1959
rect 20496 1939 20525 1958
rect 20468 1938 20525 1939
rect 20545 1938 20553 1958
rect 20411 1932 20448 1933
rect 20468 1932 20553 1938
rect 20619 1962 20657 1970
rect 20730 1966 20766 1967
rect 20619 1942 20628 1962
rect 20648 1942 20657 1962
rect 20619 1933 20657 1942
rect 20681 1958 20766 1966
rect 20681 1938 20738 1958
rect 20758 1938 20766 1958
rect 20619 1932 20656 1933
rect 20681 1932 20766 1938
rect 20832 1962 20870 1970
rect 20832 1942 20841 1962
rect 20861 1942 20870 1962
rect 20832 1933 20870 1942
rect 20832 1932 20869 1933
rect 20255 1911 20291 1932
rect 20681 1911 20712 1932
rect 20088 1907 20188 1911
rect 20088 1903 20150 1907
rect 20088 1877 20095 1903
rect 20121 1881 20150 1903
rect 20176 1881 20188 1907
rect 20121 1877 20188 1881
rect 20088 1874 20188 1877
rect 20256 1874 20291 1911
rect 20353 1908 20712 1911
rect 20353 1903 20575 1908
rect 20353 1879 20366 1903
rect 20390 1884 20575 1903
rect 20599 1884 20712 1908
rect 20390 1879 20712 1884
rect 20353 1875 20712 1879
rect 20779 1903 20928 1911
rect 20779 1883 20790 1903
rect 20810 1883 20928 1903
rect 20779 1876 20928 1883
rect 21019 1891 21058 2040
rect 20779 1875 20820 1876
rect 20103 1822 20140 1823
rect 20199 1822 20236 1823
rect 20255 1822 20291 1874
rect 20310 1822 20347 1823
rect 20003 1813 20141 1822
rect 20003 1793 20112 1813
rect 20132 1793 20141 1813
rect 18940 1789 19110 1790
rect 18940 1774 19386 1789
rect 20003 1786 20141 1793
rect 20199 1813 20347 1822
rect 20199 1793 20208 1813
rect 20228 1793 20318 1813
rect 20338 1793 20347 1813
rect 20003 1784 20099 1786
rect 18942 1763 19386 1774
rect 18942 1761 19110 1763
rect 18942 1583 18969 1761
rect 19009 1723 19073 1735
rect 19349 1731 19386 1763
rect 19557 1762 19806 1784
rect 20199 1783 20347 1793
rect 20406 1813 20443 1823
rect 20518 1822 20555 1823
rect 20499 1820 20555 1822
rect 20406 1793 20414 1813
rect 20434 1793 20443 1813
rect 20255 1782 20291 1783
rect 19557 1731 19594 1762
rect 19770 1760 19806 1762
rect 19770 1731 19807 1760
rect 19009 1722 19044 1723
rect 18986 1717 19044 1722
rect 18986 1697 18989 1717
rect 19009 1703 19044 1717
rect 19064 1703 19073 1723
rect 19009 1695 19073 1703
rect 19035 1694 19073 1695
rect 19036 1693 19073 1694
rect 19139 1727 19175 1728
rect 19247 1727 19283 1728
rect 19139 1719 19283 1727
rect 19139 1699 19147 1719
rect 19167 1718 19255 1719
rect 19167 1701 19195 1718
rect 19219 1701 19255 1718
rect 19167 1699 19255 1701
rect 19275 1699 19283 1719
rect 19139 1693 19283 1699
rect 19349 1723 19387 1731
rect 19455 1727 19491 1728
rect 19349 1703 19358 1723
rect 19378 1703 19387 1723
rect 19349 1694 19387 1703
rect 19406 1720 19491 1727
rect 19406 1700 19413 1720
rect 19434 1719 19491 1720
rect 19434 1700 19463 1719
rect 19406 1699 19463 1700
rect 19483 1699 19491 1719
rect 19349 1693 19386 1694
rect 19406 1693 19491 1699
rect 19557 1723 19595 1731
rect 19668 1727 19704 1728
rect 19557 1703 19566 1723
rect 19586 1703 19595 1723
rect 19557 1694 19595 1703
rect 19619 1719 19704 1727
rect 19619 1699 19676 1719
rect 19696 1699 19704 1719
rect 19557 1693 19594 1694
rect 19619 1693 19704 1699
rect 19770 1723 19808 1731
rect 20103 1723 20140 1724
rect 20406 1723 20443 1793
rect 20468 1813 20555 1820
rect 20468 1810 20526 1813
rect 20468 1790 20473 1810
rect 20494 1793 20526 1810
rect 20546 1793 20555 1813
rect 20494 1790 20555 1793
rect 20468 1783 20555 1790
rect 20614 1813 20651 1823
rect 20614 1793 20622 1813
rect 20642 1793 20651 1813
rect 20468 1782 20499 1783
rect 19770 1703 19779 1723
rect 19799 1703 19808 1723
rect 20102 1722 20443 1723
rect 19770 1694 19808 1703
rect 20027 1717 20443 1722
rect 20027 1697 20030 1717
rect 20050 1697 20443 1717
rect 20614 1722 20651 1793
rect 20681 1822 20712 1875
rect 21019 1873 21029 1891
rect 21047 1873 21058 1891
rect 21019 1864 21056 1873
rect 20731 1822 20768 1823
rect 20681 1813 20768 1822
rect 20681 1793 20739 1813
rect 20759 1793 20768 1813
rect 20681 1783 20768 1793
rect 20827 1813 20864 1823
rect 20827 1793 20835 1813
rect 20855 1793 20864 1813
rect 21022 1798 21059 1802
rect 20681 1782 20712 1783
rect 20827 1722 20864 1793
rect 20614 1698 20864 1722
rect 21020 1792 21059 1798
rect 21020 1774 21031 1792
rect 21049 1774 21059 1792
rect 21020 1765 21059 1774
rect 19770 1693 19807 1694
rect 19193 1672 19229 1693
rect 19619 1672 19650 1693
rect 20406 1674 20443 1697
rect 21020 1687 21055 1765
rect 21017 1677 21055 1687
rect 20406 1673 20576 1674
rect 21017 1673 21027 1677
rect 19026 1668 19126 1672
rect 19026 1664 19088 1668
rect 19026 1638 19033 1664
rect 19059 1642 19088 1664
rect 19114 1642 19126 1668
rect 19059 1638 19126 1642
rect 19026 1635 19126 1638
rect 19194 1635 19229 1672
rect 19291 1669 19650 1672
rect 19291 1664 19513 1669
rect 19291 1640 19304 1664
rect 19328 1645 19513 1664
rect 19537 1645 19650 1669
rect 19328 1640 19650 1645
rect 19291 1636 19650 1640
rect 19717 1664 19866 1672
rect 19717 1644 19728 1664
rect 19748 1644 19866 1664
rect 20406 1659 21027 1673
rect 21045 1659 21055 1677
rect 20406 1653 21055 1659
rect 20406 1652 21054 1653
rect 21017 1650 21054 1652
rect 19717 1637 19866 1644
rect 19717 1636 19758 1637
rect 19041 1583 19078 1584
rect 19137 1583 19174 1584
rect 19193 1583 19229 1635
rect 19248 1583 19285 1584
rect 18941 1574 19079 1583
rect 18941 1554 19050 1574
rect 19070 1554 19079 1574
rect 18941 1547 19079 1554
rect 19137 1574 19285 1583
rect 19137 1554 19146 1574
rect 19166 1554 19256 1574
rect 19276 1554 19285 1574
rect 18941 1545 19037 1547
rect 19137 1544 19285 1554
rect 19344 1574 19381 1584
rect 19456 1583 19493 1584
rect 19437 1581 19493 1583
rect 19344 1554 19352 1574
rect 19372 1554 19381 1574
rect 19193 1543 19229 1544
rect 19041 1484 19078 1485
rect 19344 1484 19381 1554
rect 19406 1574 19493 1581
rect 19406 1571 19464 1574
rect 19406 1551 19411 1571
rect 19432 1554 19464 1571
rect 19484 1554 19493 1574
rect 19432 1551 19493 1554
rect 19406 1544 19493 1551
rect 19552 1574 19589 1584
rect 19552 1554 19560 1574
rect 19580 1554 19589 1574
rect 19406 1543 19437 1544
rect 19040 1483 19381 1484
rect 18965 1478 19381 1483
rect 18965 1458 18968 1478
rect 18988 1458 19381 1478
rect 19552 1483 19589 1554
rect 19619 1583 19650 1636
rect 19669 1583 19706 1584
rect 19619 1574 19706 1583
rect 19619 1554 19677 1574
rect 19697 1554 19706 1574
rect 19619 1544 19706 1554
rect 19765 1574 19802 1584
rect 19765 1554 19773 1574
rect 19793 1554 19802 1574
rect 19619 1543 19650 1544
rect 19765 1483 19802 1554
rect 21020 1578 21057 1588
rect 21020 1560 21029 1578
rect 21047 1560 21057 1578
rect 21020 1551 21057 1560
rect 21020 1527 21055 1551
rect 21018 1503 21055 1527
rect 21017 1497 21055 1503
rect 19552 1459 19802 1483
rect 20428 1479 21055 1497
rect 20010 1462 20178 1463
rect 20429 1462 20453 1479
rect 20010 1436 20454 1462
rect 20010 1434 20178 1436
rect 20010 1256 20037 1434
rect 20077 1396 20141 1408
rect 20417 1404 20454 1436
rect 20625 1435 20874 1457
rect 20625 1404 20662 1435
rect 20838 1433 20874 1435
rect 21017 1438 21055 1479
rect 20838 1404 20875 1433
rect 20077 1395 20112 1396
rect 20054 1390 20112 1395
rect 20054 1370 20057 1390
rect 20077 1376 20112 1390
rect 20132 1376 20141 1396
rect 20077 1368 20141 1376
rect 20103 1367 20141 1368
rect 20104 1366 20141 1367
rect 20207 1400 20243 1401
rect 20315 1400 20351 1401
rect 20207 1394 20351 1400
rect 20207 1392 20273 1394
rect 20207 1372 20215 1392
rect 20235 1373 20273 1392
rect 20295 1392 20351 1394
rect 20295 1373 20323 1392
rect 20235 1372 20323 1373
rect 20343 1372 20351 1392
rect 20207 1366 20351 1372
rect 20417 1396 20455 1404
rect 20523 1400 20559 1401
rect 20417 1376 20426 1396
rect 20446 1376 20455 1396
rect 20417 1367 20455 1376
rect 20474 1393 20559 1400
rect 20474 1373 20481 1393
rect 20502 1392 20559 1393
rect 20502 1373 20531 1392
rect 20474 1372 20531 1373
rect 20551 1372 20559 1392
rect 20417 1366 20454 1367
rect 20474 1366 20559 1372
rect 20625 1396 20663 1404
rect 20736 1400 20772 1401
rect 20625 1376 20634 1396
rect 20654 1376 20663 1396
rect 20625 1367 20663 1376
rect 20687 1392 20772 1400
rect 20687 1372 20744 1392
rect 20764 1372 20772 1392
rect 20625 1366 20662 1367
rect 20687 1366 20772 1372
rect 20838 1396 20876 1404
rect 20838 1376 20847 1396
rect 20867 1376 20876 1396
rect 20838 1367 20876 1376
rect 21017 1403 21053 1438
rect 21017 1393 21054 1403
rect 21017 1375 21027 1393
rect 21045 1375 21054 1393
rect 20838 1366 20875 1367
rect 21017 1366 21054 1375
rect 20261 1345 20297 1366
rect 20687 1345 20718 1366
rect 20094 1341 20194 1345
rect 20094 1337 20156 1341
rect 20094 1311 20101 1337
rect 20127 1315 20156 1337
rect 20182 1315 20194 1341
rect 20127 1311 20194 1315
rect 20094 1308 20194 1311
rect 20262 1308 20297 1345
rect 20359 1342 20718 1345
rect 20359 1337 20581 1342
rect 20359 1313 20372 1337
rect 20396 1318 20581 1337
rect 20605 1318 20718 1342
rect 20396 1313 20718 1318
rect 20359 1309 20718 1313
rect 20785 1337 20934 1345
rect 20785 1317 20796 1337
rect 20816 1317 20934 1337
rect 20785 1310 20934 1317
rect 20785 1309 20826 1310
rect 20109 1256 20146 1257
rect 20205 1256 20242 1257
rect 20261 1256 20297 1308
rect 20316 1256 20353 1257
rect 20009 1247 20147 1256
rect 18265 1238 18297 1243
rect 17045 1220 17141 1222
rect 16797 1193 16806 1213
rect 16826 1193 16916 1213
rect 16936 1193 16945 1213
rect 16797 1184 16945 1193
rect 17003 1213 17141 1220
rect 17758 1217 18204 1232
rect 18034 1216 18204 1217
rect 17003 1193 17012 1213
rect 17032 1193 17141 1213
rect 17003 1184 17141 1193
rect 16797 1183 16834 1184
rect 16853 1132 16889 1184
rect 16908 1183 16945 1184
rect 17004 1183 17041 1184
rect 16324 1130 16365 1131
rect 15150 1080 15782 1087
rect 15150 1078 15212 1080
rect 14728 1068 14896 1069
rect 15150 1068 15172 1078
rect 14443 1043 14480 1044
rect 14393 1034 14480 1043
rect 14393 1014 14451 1034
rect 14471 1014 14480 1034
rect 14393 1004 14480 1014
rect 14539 1034 14576 1044
rect 14539 1014 14547 1034
rect 14567 1014 14576 1034
rect 14393 1003 14424 1004
rect 14539 943 14576 1014
rect 14326 919 14576 943
rect 14728 1042 15172 1068
rect 14728 1040 14896 1042
rect 14728 862 14755 1040
rect 14795 1002 14859 1014
rect 15135 1010 15172 1042
rect 15343 1041 15592 1063
rect 15343 1010 15380 1041
rect 15556 1039 15592 1041
rect 15556 1010 15593 1039
rect 14795 1001 14830 1002
rect 14772 996 14830 1001
rect 14772 976 14775 996
rect 14795 982 14830 996
rect 14850 982 14859 1002
rect 14795 974 14859 982
rect 14821 973 14859 974
rect 14822 972 14859 973
rect 14925 1006 14961 1007
rect 15033 1006 15069 1007
rect 14925 998 15069 1006
rect 14925 978 14933 998
rect 14953 978 14982 998
rect 14925 977 14982 978
rect 15004 978 15041 998
rect 15061 978 15069 998
rect 15004 977 15069 978
rect 14925 972 15069 977
rect 15135 1002 15173 1010
rect 15241 1006 15277 1007
rect 15135 982 15144 1002
rect 15164 982 15173 1002
rect 15135 973 15173 982
rect 15192 999 15277 1006
rect 15192 979 15199 999
rect 15220 998 15277 999
rect 15220 979 15249 998
rect 15192 978 15249 979
rect 15269 978 15277 998
rect 15135 972 15172 973
rect 15192 972 15277 978
rect 15343 1002 15381 1010
rect 15454 1006 15490 1007
rect 15343 982 15352 1002
rect 15372 982 15381 1002
rect 15343 973 15381 982
rect 15405 998 15490 1006
rect 15405 978 15462 998
rect 15482 978 15490 998
rect 15343 972 15380 973
rect 15405 972 15490 978
rect 15556 1002 15594 1010
rect 15556 982 15565 1002
rect 15585 982 15594 1002
rect 15556 973 15594 982
rect 15556 972 15593 973
rect 14979 951 15015 972
rect 15405 951 15436 972
rect 14812 947 14912 951
rect 14812 943 14874 947
rect 14812 917 14819 943
rect 14845 921 14874 943
rect 14900 921 14912 947
rect 14845 917 14912 921
rect 14812 914 14912 917
rect 14980 914 15015 951
rect 15077 948 15436 951
rect 15077 943 15299 948
rect 15077 919 15090 943
rect 15114 924 15299 943
rect 15323 924 15436 948
rect 15114 919 15436 924
rect 15077 915 15436 919
rect 15503 943 15652 951
rect 15503 923 15514 943
rect 15534 923 15652 943
rect 15503 916 15652 923
rect 15743 931 15782 1080
rect 16086 966 16125 1115
rect 16216 1123 16365 1130
rect 16216 1103 16334 1123
rect 16354 1103 16365 1123
rect 16216 1095 16365 1103
rect 16432 1127 16791 1131
rect 16432 1122 16754 1127
rect 16432 1098 16545 1122
rect 16569 1103 16754 1122
rect 16778 1103 16791 1127
rect 16569 1098 16791 1103
rect 16432 1095 16791 1098
rect 16853 1095 16888 1132
rect 16956 1129 17056 1132
rect 16956 1125 17023 1129
rect 16956 1099 16968 1125
rect 16994 1103 17023 1125
rect 17049 1103 17056 1129
rect 16994 1099 17056 1103
rect 16956 1095 17056 1099
rect 16432 1074 16463 1095
rect 16853 1074 16889 1095
rect 16275 1073 16312 1074
rect 16274 1064 16312 1073
rect 16274 1044 16283 1064
rect 16303 1044 16312 1064
rect 16274 1036 16312 1044
rect 16378 1068 16463 1074
rect 16488 1073 16525 1074
rect 16378 1048 16386 1068
rect 16406 1048 16463 1068
rect 16378 1040 16463 1048
rect 16487 1064 16525 1073
rect 16487 1044 16496 1064
rect 16516 1044 16525 1064
rect 16378 1039 16414 1040
rect 16487 1036 16525 1044
rect 16591 1068 16676 1074
rect 16696 1073 16733 1074
rect 16591 1048 16599 1068
rect 16619 1067 16676 1068
rect 16619 1048 16648 1067
rect 16591 1047 16648 1048
rect 16669 1047 16676 1067
rect 16591 1040 16676 1047
rect 16695 1064 16733 1073
rect 16695 1044 16704 1064
rect 16724 1044 16733 1064
rect 16591 1039 16627 1040
rect 16695 1036 16733 1044
rect 16799 1069 16943 1074
rect 16799 1068 16864 1069
rect 16799 1048 16807 1068
rect 16827 1048 16864 1068
rect 16886 1068 16943 1069
rect 16886 1048 16915 1068
rect 16935 1048 16943 1068
rect 16799 1040 16943 1048
rect 16799 1039 16835 1040
rect 16907 1039 16943 1040
rect 17009 1073 17046 1074
rect 17009 1072 17047 1073
rect 17009 1064 17073 1072
rect 17009 1044 17018 1064
rect 17038 1050 17073 1064
rect 17093 1050 17096 1070
rect 17038 1045 17096 1050
rect 17038 1044 17073 1045
rect 16275 1007 16312 1036
rect 16276 1005 16312 1007
rect 16488 1005 16525 1036
rect 16276 983 16525 1005
rect 16696 1004 16733 1036
rect 17009 1032 17073 1044
rect 17113 1006 17140 1184
rect 16972 1004 17140 1006
rect 16696 978 17140 1004
rect 17292 1103 17542 1127
rect 17292 1032 17329 1103
rect 17444 1042 17475 1043
rect 17292 1012 17301 1032
rect 17321 1012 17329 1032
rect 17292 1002 17329 1012
rect 17388 1032 17475 1042
rect 17388 1012 17397 1032
rect 17417 1012 17475 1032
rect 17388 1003 17475 1012
rect 17388 1002 17425 1003
rect 16696 968 16718 978
rect 16972 977 17140 978
rect 16656 966 16718 968
rect 16086 959 16718 966
rect 15503 915 15544 916
rect 14827 862 14864 863
rect 14923 862 14960 863
rect 14979 862 15015 914
rect 15034 862 15071 863
rect 12892 817 12897 843
rect 12916 817 12923 843
rect 14727 853 14865 862
rect 14727 833 14836 853
rect 14856 833 14865 853
rect 14727 826 14865 833
rect 14923 853 15071 862
rect 14923 833 14932 853
rect 14952 833 15042 853
rect 15062 833 15071 853
rect 14727 824 14823 826
rect 14923 823 15071 833
rect 15130 853 15167 863
rect 15242 862 15279 863
rect 15223 860 15279 862
rect 15130 833 15138 853
rect 15158 833 15167 853
rect 14979 822 15015 823
rect 12892 814 12923 817
rect 11721 790 11859 799
rect 11515 789 11552 790
rect 11571 738 11607 790
rect 11626 789 11663 790
rect 11722 789 11759 790
rect 11042 736 11083 737
rect 10934 729 11083 736
rect 10934 709 11052 729
rect 11072 709 11083 729
rect 10934 701 11083 709
rect 11150 733 11509 737
rect 11150 728 11472 733
rect 11150 704 11263 728
rect 11287 709 11472 728
rect 11496 709 11509 733
rect 11287 704 11509 709
rect 11150 701 11509 704
rect 11571 701 11606 738
rect 11674 735 11774 738
rect 11674 731 11741 735
rect 11674 705 11686 731
rect 11712 709 11741 731
rect 11767 709 11774 735
rect 11712 705 11774 709
rect 11674 701 11774 705
rect 10361 688 10399 698
rect 9750 684 9920 685
rect 10361 684 10371 688
rect 9750 670 10371 684
rect 10389 670 10399 688
rect 11150 680 11181 701
rect 11571 680 11607 701
rect 9750 664 10399 670
rect 10814 671 10851 680
rect 10993 679 11030 680
rect 9750 663 10398 664
rect 10361 661 10398 663
rect 10814 653 10823 671
rect 10841 653 10851 671
rect 10814 643 10851 653
rect 10815 608 10851 643
rect 10992 670 11030 679
rect 10992 650 11001 670
rect 11021 650 11030 670
rect 10992 642 11030 650
rect 11096 674 11181 680
rect 11206 679 11243 680
rect 11096 654 11104 674
rect 11124 654 11181 674
rect 11096 646 11181 654
rect 11205 670 11243 679
rect 11205 650 11214 670
rect 11234 650 11243 670
rect 11096 645 11132 646
rect 11205 642 11243 650
rect 11309 674 11394 680
rect 11414 679 11451 680
rect 11309 654 11317 674
rect 11337 673 11394 674
rect 11337 654 11366 673
rect 11309 653 11366 654
rect 11387 653 11394 673
rect 11309 646 11394 653
rect 11413 670 11451 679
rect 11413 650 11422 670
rect 11442 650 11451 670
rect 11309 645 11345 646
rect 11413 642 11451 650
rect 11517 674 11661 680
rect 11517 654 11525 674
rect 11545 673 11633 674
rect 11545 654 11573 673
rect 11517 652 11573 654
rect 11595 654 11633 673
rect 11653 654 11661 674
rect 11595 652 11661 654
rect 11517 646 11661 652
rect 11517 645 11553 646
rect 11625 645 11661 646
rect 11727 679 11764 680
rect 11727 678 11765 679
rect 11727 670 11791 678
rect 11727 650 11736 670
rect 11756 656 11791 670
rect 11811 656 11814 676
rect 11756 651 11814 656
rect 11756 650 11791 651
rect 10993 613 11030 642
rect 10364 597 10401 599
rect 6310 581 6478 583
rect 6034 555 6478 581
rect 6035 529 6059 555
rect 6310 554 6478 555
rect 10359 589 10401 597
rect 10359 571 10373 589
rect 10391 571 10401 589
rect 10359 562 10401 571
rect 6028 521 6068 529
rect 6028 514 6037 521
rect 5433 499 6037 514
rect 6060 499 6068 521
rect 5433 496 6068 499
rect 5433 490 5471 496
rect 6028 484 6068 496
rect 10359 521 10400 562
rect 10359 499 10370 521
rect 10393 499 10400 521
rect 10813 543 10851 608
rect 10994 611 11030 613
rect 11206 611 11243 642
rect 10994 589 11243 611
rect 11414 610 11451 642
rect 11727 638 11791 650
rect 11831 612 11858 790
rect 14827 763 14864 764
rect 15130 763 15167 833
rect 15192 853 15279 860
rect 15192 850 15250 853
rect 15192 830 15197 850
rect 15218 833 15250 850
rect 15270 833 15279 853
rect 15218 830 15279 833
rect 15192 823 15279 830
rect 15338 853 15375 863
rect 15338 833 15346 853
rect 15366 833 15375 853
rect 15192 822 15223 823
rect 14826 762 15167 763
rect 14751 757 15167 762
rect 14751 737 14754 757
rect 14774 737 15167 757
rect 15338 762 15375 833
rect 15405 862 15436 915
rect 15743 913 15753 931
rect 15771 913 15782 931
rect 16085 950 16718 959
rect 17444 950 17475 1003
rect 17505 1032 17542 1103
rect 17713 1108 18106 1128
rect 18126 1108 18129 1128
rect 17713 1103 18129 1108
rect 17713 1102 18054 1103
rect 17657 1042 17688 1043
rect 17505 1012 17514 1032
rect 17534 1012 17542 1032
rect 17505 1002 17542 1012
rect 17601 1035 17688 1042
rect 17601 1032 17662 1035
rect 17601 1012 17610 1032
rect 17630 1015 17662 1032
rect 17683 1015 17688 1035
rect 17630 1012 17688 1015
rect 17601 1005 17688 1012
rect 17713 1032 17750 1102
rect 18016 1101 18053 1102
rect 17865 1042 17901 1043
rect 17713 1012 17722 1032
rect 17742 1012 17750 1032
rect 17601 1003 17657 1005
rect 17601 1002 17638 1003
rect 17713 1002 17750 1012
rect 17809 1032 17957 1042
rect 18057 1039 18153 1041
rect 17809 1012 17818 1032
rect 17838 1012 17928 1032
rect 17948 1012 17957 1032
rect 17809 1003 17957 1012
rect 18015 1032 18153 1039
rect 18015 1012 18024 1032
rect 18044 1012 18153 1032
rect 18015 1003 18153 1012
rect 17809 1002 17846 1003
rect 17865 951 17901 1003
rect 17920 1002 17957 1003
rect 18016 1002 18053 1003
rect 16085 932 16095 950
rect 16113 949 16718 950
rect 17336 949 17377 950
rect 16113 944 16134 949
rect 16113 932 16125 944
rect 17228 942 17377 949
rect 16085 924 16125 932
rect 16168 931 16194 932
rect 16085 922 16122 924
rect 16168 913 16722 931
rect 17228 922 17346 942
rect 17366 922 17377 942
rect 17228 914 17377 922
rect 17444 946 17803 950
rect 17444 941 17766 946
rect 17444 917 17557 941
rect 17581 922 17766 941
rect 17790 922 17803 946
rect 17581 917 17803 922
rect 17444 914 17803 917
rect 17865 914 17900 951
rect 17968 948 18068 951
rect 17968 944 18035 948
rect 17968 918 17980 944
rect 18006 922 18035 944
rect 18061 922 18068 948
rect 18006 918 18068 922
rect 17968 914 18068 918
rect 15743 904 15780 913
rect 15455 862 15492 863
rect 15405 853 15492 862
rect 15405 833 15463 853
rect 15483 833 15492 853
rect 15405 823 15492 833
rect 15551 853 15588 863
rect 15551 833 15559 853
rect 15579 833 15588 853
rect 16088 854 16125 860
rect 16168 854 16194 913
rect 16701 894 16722 913
rect 16088 851 16194 854
rect 15746 838 15783 842
rect 15405 822 15436 823
rect 15551 762 15588 833
rect 15338 738 15588 762
rect 15744 832 15783 838
rect 15744 814 15755 832
rect 15773 814 15783 832
rect 16088 833 16097 851
rect 16115 837 16194 851
rect 16279 869 16529 893
rect 16115 835 16191 837
rect 16115 833 16125 835
rect 16088 823 16125 833
rect 15744 805 15783 814
rect 15130 714 15167 737
rect 15744 727 15779 805
rect 16093 758 16124 823
rect 16279 798 16316 869
rect 16431 808 16462 809
rect 16279 778 16288 798
rect 16308 778 16316 798
rect 16279 768 16316 778
rect 16375 798 16462 808
rect 16375 778 16384 798
rect 16404 778 16462 798
rect 16375 769 16462 778
rect 16375 768 16412 769
rect 15741 717 15779 727
rect 16092 749 16129 758
rect 16092 731 16102 749
rect 16120 731 16129 749
rect 16092 721 16129 731
rect 15130 713 15300 714
rect 15741 713 15751 717
rect 15130 699 15751 713
rect 15769 699 15779 717
rect 16431 716 16462 769
rect 16492 798 16529 869
rect 16700 874 17093 894
rect 17113 874 17116 894
rect 17444 893 17475 914
rect 17865 893 17901 914
rect 17287 892 17324 893
rect 16700 869 17116 874
rect 17286 883 17324 892
rect 16700 868 17041 869
rect 16644 808 16675 809
rect 16492 778 16501 798
rect 16521 778 16529 798
rect 16492 768 16529 778
rect 16588 801 16675 808
rect 16588 798 16649 801
rect 16588 778 16597 798
rect 16617 781 16649 798
rect 16670 781 16675 801
rect 16617 778 16675 781
rect 16588 771 16675 778
rect 16700 798 16737 868
rect 17003 867 17040 868
rect 17286 863 17295 883
rect 17315 863 17324 883
rect 17286 855 17324 863
rect 17390 887 17475 893
rect 17500 892 17537 893
rect 17390 867 17398 887
rect 17418 867 17475 887
rect 17390 859 17475 867
rect 17499 883 17537 892
rect 17499 863 17508 883
rect 17528 863 17537 883
rect 17390 858 17426 859
rect 17499 855 17537 863
rect 17603 887 17688 893
rect 17708 892 17745 893
rect 17603 867 17611 887
rect 17631 886 17688 887
rect 17631 867 17660 886
rect 17603 866 17660 867
rect 17681 866 17688 886
rect 17603 859 17688 866
rect 17707 883 17745 892
rect 17707 863 17716 883
rect 17736 863 17745 883
rect 17603 858 17639 859
rect 17707 855 17745 863
rect 17811 888 17955 893
rect 17811 887 17870 888
rect 17811 867 17819 887
rect 17839 868 17870 887
rect 17894 887 17955 888
rect 17894 868 17927 887
rect 17839 867 17927 868
rect 17947 867 17955 887
rect 17811 859 17955 867
rect 17811 858 17847 859
rect 17919 858 17955 859
rect 18021 892 18058 893
rect 18021 891 18059 892
rect 18021 883 18085 891
rect 18021 863 18030 883
rect 18050 869 18085 883
rect 18105 869 18108 889
rect 18050 864 18108 869
rect 18050 863 18085 864
rect 17287 826 17324 855
rect 17288 824 17324 826
rect 17500 824 17537 855
rect 16852 808 16888 809
rect 16700 778 16709 798
rect 16729 778 16737 798
rect 16588 769 16644 771
rect 16588 768 16625 769
rect 16700 768 16737 778
rect 16796 798 16944 808
rect 17044 805 17140 807
rect 16796 778 16805 798
rect 16825 778 16915 798
rect 16935 778 16944 798
rect 16796 769 16944 778
rect 17002 798 17140 805
rect 17288 802 17537 824
rect 17708 823 17745 855
rect 18021 851 18085 863
rect 18125 825 18152 1003
rect 17984 823 18152 825
rect 17708 819 18152 823
rect 17002 778 17011 798
rect 17031 778 17140 798
rect 17708 800 17757 819
rect 17777 800 18152 819
rect 17708 797 18152 800
rect 17984 796 18152 797
rect 18173 822 18204 1216
rect 18265 1220 18270 1238
rect 18290 1220 18297 1238
rect 18265 1215 18297 1220
rect 18268 1213 18297 1215
rect 18997 1228 19165 1229
rect 18997 1225 19441 1228
rect 18997 1206 19372 1225
rect 19392 1206 19441 1225
rect 20009 1227 20118 1247
rect 20138 1227 20147 1247
rect 18997 1202 19441 1206
rect 18997 1200 19165 1202
rect 18997 1022 19024 1200
rect 19064 1162 19128 1174
rect 19404 1170 19441 1202
rect 19612 1201 19861 1223
rect 20009 1220 20147 1227
rect 20205 1247 20353 1256
rect 20205 1227 20214 1247
rect 20234 1227 20324 1247
rect 20344 1227 20353 1247
rect 20009 1218 20105 1220
rect 20205 1217 20353 1227
rect 20412 1247 20449 1257
rect 20524 1256 20561 1257
rect 20505 1254 20561 1256
rect 20412 1227 20420 1247
rect 20440 1227 20449 1247
rect 20261 1216 20297 1217
rect 19612 1170 19649 1201
rect 19825 1199 19861 1201
rect 19825 1170 19862 1199
rect 19064 1161 19099 1162
rect 19041 1156 19099 1161
rect 19041 1136 19044 1156
rect 19064 1142 19099 1156
rect 19119 1142 19128 1162
rect 19064 1134 19128 1142
rect 19090 1133 19128 1134
rect 19091 1132 19128 1133
rect 19194 1166 19230 1167
rect 19302 1166 19338 1167
rect 19194 1158 19338 1166
rect 19194 1138 19202 1158
rect 19222 1138 19254 1158
rect 19278 1138 19310 1158
rect 19330 1138 19338 1158
rect 19194 1132 19338 1138
rect 19404 1162 19442 1170
rect 19510 1166 19546 1167
rect 19404 1142 19413 1162
rect 19433 1142 19442 1162
rect 19404 1133 19442 1142
rect 19461 1159 19546 1166
rect 19461 1139 19468 1159
rect 19489 1158 19546 1159
rect 19489 1139 19518 1158
rect 19461 1138 19518 1139
rect 19538 1138 19546 1158
rect 19404 1132 19441 1133
rect 19461 1132 19546 1138
rect 19612 1162 19650 1170
rect 19723 1166 19759 1167
rect 19612 1142 19621 1162
rect 19641 1142 19650 1162
rect 19612 1133 19650 1142
rect 19674 1158 19759 1166
rect 19674 1138 19731 1158
rect 19751 1138 19759 1158
rect 19612 1132 19649 1133
rect 19674 1132 19759 1138
rect 19825 1162 19863 1170
rect 19825 1142 19834 1162
rect 19854 1142 19863 1162
rect 20109 1157 20146 1158
rect 20412 1157 20449 1227
rect 20474 1247 20561 1254
rect 20474 1244 20532 1247
rect 20474 1224 20479 1244
rect 20500 1227 20532 1244
rect 20552 1227 20561 1247
rect 20500 1224 20561 1227
rect 20474 1217 20561 1224
rect 20620 1247 20657 1257
rect 20620 1227 20628 1247
rect 20648 1227 20657 1247
rect 20474 1216 20505 1217
rect 20108 1156 20449 1157
rect 19825 1133 19863 1142
rect 20033 1151 20449 1156
rect 19825 1132 19862 1133
rect 19248 1111 19284 1132
rect 19674 1111 19705 1132
rect 20033 1131 20036 1151
rect 20056 1131 20449 1151
rect 20620 1156 20657 1227
rect 20687 1256 20718 1309
rect 21020 1294 21057 1304
rect 21020 1276 21029 1294
rect 21047 1276 21057 1294
rect 21020 1267 21057 1276
rect 20737 1256 20774 1257
rect 20687 1247 20774 1256
rect 20687 1227 20745 1247
rect 20765 1227 20774 1247
rect 20687 1217 20774 1227
rect 20833 1247 20870 1257
rect 20833 1227 20841 1247
rect 20861 1227 20870 1247
rect 20687 1216 20718 1217
rect 20833 1156 20870 1227
rect 21025 1202 21056 1267
rect 21024 1192 21061 1202
rect 21024 1190 21034 1192
rect 20958 1188 21034 1190
rect 20620 1132 20870 1156
rect 20955 1174 21034 1188
rect 21052 1174 21061 1192
rect 20955 1171 21061 1174
rect 20427 1112 20448 1131
rect 20955 1112 20981 1171
rect 21024 1165 21061 1171
rect 19081 1107 19181 1111
rect 19081 1103 19143 1107
rect 19081 1077 19088 1103
rect 19114 1081 19143 1103
rect 19169 1081 19181 1107
rect 19114 1077 19181 1081
rect 19081 1074 19181 1077
rect 19249 1074 19284 1111
rect 19346 1108 19705 1111
rect 19346 1103 19568 1108
rect 19346 1079 19359 1103
rect 19383 1084 19568 1103
rect 19592 1084 19705 1108
rect 19383 1079 19705 1084
rect 19346 1075 19705 1079
rect 19772 1103 19921 1111
rect 19772 1083 19783 1103
rect 19803 1083 19921 1103
rect 20427 1094 20981 1112
rect 21027 1101 21064 1103
rect 20955 1093 20981 1094
rect 21024 1093 21064 1101
rect 19772 1076 19921 1083
rect 21024 1081 21036 1093
rect 21015 1076 21036 1081
rect 19772 1075 19813 1076
rect 20431 1075 21036 1076
rect 21054 1075 21064 1093
rect 19096 1022 19133 1023
rect 19192 1022 19229 1023
rect 19248 1022 19284 1074
rect 19303 1022 19340 1023
rect 18996 1013 19134 1022
rect 18996 993 19105 1013
rect 19125 993 19134 1013
rect 18996 986 19134 993
rect 19192 1013 19340 1022
rect 19192 993 19201 1013
rect 19221 993 19311 1013
rect 19331 993 19340 1013
rect 18996 984 19092 986
rect 19192 983 19340 993
rect 19399 1013 19436 1023
rect 19511 1022 19548 1023
rect 19492 1020 19548 1022
rect 19399 993 19407 1013
rect 19427 993 19436 1013
rect 19248 982 19284 983
rect 19096 923 19133 924
rect 19399 923 19436 993
rect 19461 1013 19548 1020
rect 19461 1010 19519 1013
rect 19461 990 19466 1010
rect 19487 993 19519 1010
rect 19539 993 19548 1013
rect 19487 990 19548 993
rect 19461 983 19548 990
rect 19607 1013 19644 1023
rect 19607 993 19615 1013
rect 19635 993 19644 1013
rect 19461 982 19492 983
rect 19095 922 19436 923
rect 19020 917 19436 922
rect 19020 897 19023 917
rect 19043 897 19436 917
rect 19607 922 19644 993
rect 19674 1022 19705 1075
rect 20431 1066 21064 1075
rect 20431 1059 21063 1066
rect 20431 1057 20493 1059
rect 20009 1047 20177 1048
rect 20431 1047 20453 1057
rect 19724 1022 19761 1023
rect 19674 1013 19761 1022
rect 19674 993 19732 1013
rect 19752 993 19761 1013
rect 19674 983 19761 993
rect 19820 1013 19857 1023
rect 19820 993 19828 1013
rect 19848 993 19857 1013
rect 19674 982 19705 983
rect 19820 922 19857 993
rect 19607 898 19857 922
rect 20009 1021 20453 1047
rect 20009 1019 20177 1021
rect 20009 841 20036 1019
rect 20076 981 20140 993
rect 20416 989 20453 1021
rect 20624 1020 20873 1042
rect 20624 989 20661 1020
rect 20837 1018 20873 1020
rect 20837 989 20874 1018
rect 20076 980 20111 981
rect 20053 975 20111 980
rect 20053 955 20056 975
rect 20076 961 20111 975
rect 20131 961 20140 981
rect 20076 953 20140 961
rect 20102 952 20140 953
rect 20103 951 20140 952
rect 20206 985 20242 986
rect 20314 985 20350 986
rect 20206 977 20350 985
rect 20206 957 20214 977
rect 20234 957 20263 977
rect 20206 956 20263 957
rect 20285 957 20322 977
rect 20342 957 20350 977
rect 20285 956 20350 957
rect 20206 951 20350 956
rect 20416 981 20454 989
rect 20522 985 20558 986
rect 20416 961 20425 981
rect 20445 961 20454 981
rect 20416 952 20454 961
rect 20473 978 20558 985
rect 20473 958 20480 978
rect 20501 977 20558 978
rect 20501 958 20530 977
rect 20473 957 20530 958
rect 20550 957 20558 977
rect 20416 951 20453 952
rect 20473 951 20558 957
rect 20624 981 20662 989
rect 20735 985 20771 986
rect 20624 961 20633 981
rect 20653 961 20662 981
rect 20624 952 20662 961
rect 20686 977 20771 985
rect 20686 957 20743 977
rect 20763 957 20771 977
rect 20624 951 20661 952
rect 20686 951 20771 957
rect 20837 981 20875 989
rect 20837 961 20846 981
rect 20866 961 20875 981
rect 20837 952 20875 961
rect 20837 951 20874 952
rect 20260 930 20296 951
rect 20686 930 20717 951
rect 20093 926 20193 930
rect 20093 922 20155 926
rect 20093 896 20100 922
rect 20126 900 20155 922
rect 20181 900 20193 926
rect 20126 896 20193 900
rect 20093 893 20193 896
rect 20261 893 20296 930
rect 20358 927 20717 930
rect 20358 922 20580 927
rect 20358 898 20371 922
rect 20395 903 20580 922
rect 20604 903 20717 927
rect 20395 898 20717 903
rect 20358 894 20717 898
rect 20784 922 20933 930
rect 20784 902 20795 922
rect 20815 902 20933 922
rect 20784 895 20933 902
rect 21024 910 21063 1059
rect 20784 894 20825 895
rect 20108 841 20145 842
rect 20204 841 20241 842
rect 20260 841 20296 893
rect 20315 841 20352 842
rect 18173 796 18178 822
rect 18197 796 18204 822
rect 20008 832 20146 841
rect 20008 812 20117 832
rect 20137 812 20146 832
rect 20008 805 20146 812
rect 20204 832 20352 841
rect 20204 812 20213 832
rect 20233 812 20323 832
rect 20343 812 20352 832
rect 20008 803 20104 805
rect 20204 802 20352 812
rect 20411 832 20448 842
rect 20523 841 20560 842
rect 20504 839 20560 841
rect 20411 812 20419 832
rect 20439 812 20448 832
rect 20260 801 20296 802
rect 18173 793 18204 796
rect 17002 769 17140 778
rect 16796 768 16833 769
rect 16852 717 16888 769
rect 16907 768 16944 769
rect 17003 768 17040 769
rect 16323 715 16364 716
rect 15130 693 15779 699
rect 16215 708 16364 715
rect 15130 692 15778 693
rect 15741 690 15778 692
rect 16215 688 16333 708
rect 16353 688 16364 708
rect 16215 680 16364 688
rect 16431 712 16790 716
rect 16431 707 16753 712
rect 16431 683 16544 707
rect 16568 688 16753 707
rect 16777 688 16790 712
rect 16568 683 16790 688
rect 16431 680 16790 683
rect 16852 680 16887 717
rect 16955 714 17055 717
rect 16955 710 17022 714
rect 16955 684 16967 710
rect 16993 688 17022 710
rect 17048 688 17055 714
rect 16993 684 17055 688
rect 16955 680 17055 684
rect 16431 659 16462 680
rect 16852 659 16888 680
rect 16095 650 16132 659
rect 16274 658 16311 659
rect 16095 632 16104 650
rect 16122 632 16132 650
rect 15744 626 15781 628
rect 11690 610 11858 612
rect 11414 584 11858 610
rect 11415 558 11439 584
rect 11690 583 11858 584
rect 15739 618 15781 626
rect 16095 622 16132 632
rect 15739 600 15753 618
rect 15771 600 15781 618
rect 15739 591 15781 600
rect 11408 550 11448 558
rect 11408 543 11417 550
rect 10813 528 11417 543
rect 11440 528 11448 550
rect 10813 525 11448 528
rect 10813 519 10851 525
rect 11408 513 11448 525
rect 15739 550 15780 591
rect 16096 587 16132 622
rect 16273 649 16311 658
rect 16273 629 16282 649
rect 16302 629 16311 649
rect 16273 621 16311 629
rect 16377 653 16462 659
rect 16487 658 16524 659
rect 16377 633 16385 653
rect 16405 633 16462 653
rect 16377 625 16462 633
rect 16486 649 16524 658
rect 16486 629 16495 649
rect 16515 629 16524 649
rect 16377 624 16413 625
rect 16486 621 16524 629
rect 16590 653 16675 659
rect 16695 658 16732 659
rect 16590 633 16598 653
rect 16618 652 16675 653
rect 16618 633 16647 652
rect 16590 632 16647 633
rect 16668 632 16675 652
rect 16590 625 16675 632
rect 16694 649 16732 658
rect 16694 629 16703 649
rect 16723 629 16732 649
rect 16590 624 16626 625
rect 16694 621 16732 629
rect 16798 653 16942 659
rect 16798 633 16806 653
rect 16826 652 16914 653
rect 16826 633 16854 652
rect 16798 631 16854 633
rect 16876 633 16914 652
rect 16934 633 16942 653
rect 16876 631 16942 633
rect 16798 625 16942 631
rect 16798 624 16834 625
rect 16906 624 16942 625
rect 17008 658 17045 659
rect 17008 657 17046 658
rect 17008 649 17072 657
rect 17008 629 17017 649
rect 17037 635 17072 649
rect 17092 635 17095 655
rect 17037 630 17095 635
rect 17037 629 17072 630
rect 16274 592 16311 621
rect 15739 528 15750 550
rect 15773 528 15780 550
rect 15739 523 15780 528
rect 16094 522 16132 587
rect 16275 590 16311 592
rect 16487 590 16524 621
rect 16275 568 16524 590
rect 16695 589 16732 621
rect 17008 617 17072 629
rect 17112 591 17139 769
rect 20108 742 20145 743
rect 20411 742 20448 812
rect 20473 832 20560 839
rect 20473 829 20531 832
rect 20473 809 20478 829
rect 20499 812 20531 829
rect 20551 812 20560 832
rect 20499 809 20560 812
rect 20473 802 20560 809
rect 20619 832 20656 842
rect 20619 812 20627 832
rect 20647 812 20656 832
rect 20473 801 20504 802
rect 20107 741 20448 742
rect 20032 736 20448 741
rect 20032 716 20035 736
rect 20055 716 20448 736
rect 20619 741 20656 812
rect 20686 841 20717 894
rect 21024 892 21034 910
rect 21052 892 21063 910
rect 21024 883 21061 892
rect 20736 841 20773 842
rect 20686 832 20773 841
rect 20686 812 20744 832
rect 20764 812 20773 832
rect 20686 802 20773 812
rect 20832 832 20869 842
rect 20832 812 20840 832
rect 20860 812 20869 832
rect 21027 817 21064 821
rect 20686 801 20717 802
rect 20832 741 20869 812
rect 20619 717 20869 741
rect 21025 811 21064 817
rect 21025 793 21036 811
rect 21054 793 21064 811
rect 21025 784 21064 793
rect 20411 693 20448 716
rect 21025 706 21060 784
rect 21022 696 21060 706
rect 20411 692 20581 693
rect 21022 692 21032 696
rect 20411 678 21032 692
rect 21050 678 21060 696
rect 20411 672 21060 678
rect 20411 671 21059 672
rect 21022 669 21059 671
rect 21025 605 21062 607
rect 16971 589 17139 591
rect 16695 563 17139 589
rect 16696 537 16720 563
rect 16971 562 17139 563
rect 21020 597 21062 605
rect 21020 579 21034 597
rect 21052 579 21062 597
rect 21020 570 21062 579
rect 16689 529 16729 537
rect 16689 522 16698 529
rect 10359 494 10400 499
rect 16094 507 16698 522
rect 16721 507 16729 529
rect 16094 504 16729 507
rect 16094 498 16132 504
rect 16689 492 16729 504
rect 21020 529 21061 570
rect 21020 507 21031 529
rect 21054 507 21061 529
rect 21020 502 21061 507
rect 1740 401 1990 425
rect 1740 330 1777 401
rect 1892 340 1923 341
rect 1740 310 1749 330
rect 1769 310 1777 330
rect 1740 300 1777 310
rect 1836 330 1923 340
rect 1836 310 1845 330
rect 1865 310 1923 330
rect 1836 301 1923 310
rect 1836 300 1873 301
rect 1892 248 1923 301
rect 1953 330 1990 401
rect 2161 406 2554 426
rect 2574 406 2577 426
rect 2161 401 2577 406
rect 12401 409 12651 433
rect 2161 400 2502 401
rect 2105 340 2136 341
rect 1953 310 1962 330
rect 1982 310 1990 330
rect 1953 300 1990 310
rect 2049 333 2136 340
rect 2049 330 2110 333
rect 2049 310 2058 330
rect 2078 313 2110 330
rect 2131 313 2136 333
rect 2078 310 2136 313
rect 2049 303 2136 310
rect 2161 330 2198 400
rect 2464 399 2501 400
rect 7021 380 7271 404
rect 2313 340 2349 341
rect 2161 310 2170 330
rect 2190 310 2198 330
rect 2049 301 2105 303
rect 2049 300 2086 301
rect 2161 300 2198 310
rect 2257 330 2405 340
rect 2505 337 2601 339
rect 2257 310 2266 330
rect 2286 310 2376 330
rect 2396 310 2405 330
rect 2257 301 2405 310
rect 2463 336 2601 337
rect 2463 331 2687 336
rect 2463 330 2651 331
rect 2463 310 2472 330
rect 2492 311 2651 330
rect 2679 311 2687 331
rect 2492 310 2687 311
rect 2463 303 2687 310
rect 4830 313 5080 337
rect 2463 301 2601 303
rect 2257 300 2294 301
rect 2313 249 2349 301
rect 2368 300 2405 301
rect 2464 300 2501 301
rect 1784 247 1825 248
rect 1676 240 1825 247
rect 1676 220 1794 240
rect 1814 220 1825 240
rect 1676 212 1825 220
rect 1892 244 2251 248
rect 1892 239 2214 244
rect 1892 215 2005 239
rect 2029 220 2214 239
rect 2238 220 2251 244
rect 2029 215 2251 220
rect 1892 212 2251 215
rect 2313 212 2348 249
rect 2416 246 2516 249
rect 2416 242 2483 246
rect 2416 216 2428 242
rect 2454 220 2483 242
rect 2509 220 2516 246
rect 2454 216 2516 220
rect 2416 212 2516 216
rect 1892 191 1923 212
rect 2313 191 2349 212
rect 1735 190 1772 191
rect 1734 181 1772 190
rect 1734 161 1743 181
rect 1763 161 1772 181
rect 1734 153 1772 161
rect 1838 185 1923 191
rect 1948 190 1985 191
rect 1838 165 1846 185
rect 1866 165 1923 185
rect 1838 157 1923 165
rect 1947 181 1985 190
rect 1947 161 1956 181
rect 1976 161 1985 181
rect 1838 156 1874 157
rect 1947 153 1985 161
rect 2051 185 2136 191
rect 2156 190 2193 191
rect 2051 165 2059 185
rect 2079 184 2136 185
rect 2079 165 2108 184
rect 2051 164 2108 165
rect 2129 164 2136 184
rect 2051 157 2136 164
rect 2155 181 2193 190
rect 2155 161 2164 181
rect 2184 161 2193 181
rect 2051 156 2087 157
rect 2155 153 2193 161
rect 2259 185 2403 191
rect 2259 165 2267 185
rect 2287 184 2375 185
rect 2287 165 2322 184
rect 2259 162 2322 165
rect 2347 165 2375 184
rect 2395 165 2403 185
rect 2347 162 2403 165
rect 2259 157 2403 162
rect 2259 156 2295 157
rect 2367 156 2403 157
rect 2469 190 2506 191
rect 2469 189 2507 190
rect 2469 181 2533 189
rect 2469 161 2478 181
rect 2498 167 2533 181
rect 2553 167 2556 187
rect 2498 162 2556 167
rect 2498 161 2533 162
rect 1735 124 1772 153
rect 1736 122 1772 124
rect 1948 122 1985 153
rect 1736 100 1985 122
rect 2156 121 2193 153
rect 2469 149 2533 161
rect 2573 123 2600 301
rect 4830 242 4867 313
rect 4982 252 5013 253
rect 4830 222 4839 242
rect 4859 222 4867 242
rect 4830 212 4867 222
rect 4926 242 5013 252
rect 4926 222 4935 242
rect 4955 222 5013 242
rect 4926 213 5013 222
rect 4926 212 4963 213
rect 4982 160 5013 213
rect 5043 242 5080 313
rect 5251 318 5644 338
rect 5664 318 5667 338
rect 5251 313 5667 318
rect 5251 312 5592 313
rect 5195 252 5226 253
rect 5043 222 5052 242
rect 5072 222 5080 242
rect 5043 212 5080 222
rect 5139 245 5226 252
rect 5139 242 5200 245
rect 5139 222 5148 242
rect 5168 225 5200 242
rect 5221 225 5226 245
rect 5168 222 5226 225
rect 5139 215 5226 222
rect 5251 242 5288 312
rect 5554 311 5591 312
rect 7021 309 7058 380
rect 7173 319 7204 320
rect 7021 289 7030 309
rect 7050 289 7058 309
rect 7021 279 7058 289
rect 7117 309 7204 319
rect 7117 289 7126 309
rect 7146 289 7204 309
rect 7117 280 7204 289
rect 7117 279 7154 280
rect 5403 252 5439 253
rect 5251 222 5260 242
rect 5280 222 5288 242
rect 5139 213 5195 215
rect 5139 212 5176 213
rect 5251 212 5288 222
rect 5347 242 5495 252
rect 5595 249 5691 251
rect 5347 222 5356 242
rect 5376 222 5466 242
rect 5486 222 5495 242
rect 5347 213 5495 222
rect 5553 242 5691 249
rect 5553 222 5562 242
rect 5582 222 5691 242
rect 7173 227 7204 280
rect 7234 309 7271 380
rect 7442 385 7835 405
rect 7855 385 7858 405
rect 7442 380 7858 385
rect 7442 379 7783 380
rect 7386 319 7417 320
rect 7234 289 7243 309
rect 7263 289 7271 309
rect 7234 279 7271 289
rect 7330 312 7417 319
rect 7330 309 7391 312
rect 7330 289 7339 309
rect 7359 292 7391 309
rect 7412 292 7417 312
rect 7359 289 7417 292
rect 7330 282 7417 289
rect 7442 309 7479 379
rect 7745 378 7782 379
rect 12401 338 12438 409
rect 12553 348 12584 349
rect 7594 319 7630 320
rect 7442 289 7451 309
rect 7471 289 7479 309
rect 7330 280 7386 282
rect 7330 279 7367 280
rect 7442 279 7479 289
rect 7538 309 7686 319
rect 7786 316 7882 318
rect 7538 289 7547 309
rect 7567 289 7657 309
rect 7677 289 7686 309
rect 7538 280 7686 289
rect 7744 315 7882 316
rect 7744 310 7968 315
rect 7744 309 7932 310
rect 7744 289 7753 309
rect 7773 290 7932 309
rect 7960 290 7968 310
rect 7773 289 7968 290
rect 7744 282 7968 289
rect 10091 306 10341 330
rect 7744 280 7882 282
rect 7538 279 7575 280
rect 7594 228 7630 280
rect 7649 279 7686 280
rect 7745 279 7782 280
rect 7065 226 7106 227
rect 5553 213 5691 222
rect 6957 219 7106 226
rect 5347 212 5384 213
rect 5403 161 5439 213
rect 5458 212 5495 213
rect 5554 212 5591 213
rect 4874 159 4915 160
rect 4766 152 4915 159
rect 4766 132 4884 152
rect 4904 132 4915 152
rect 4766 124 4915 132
rect 4982 156 5341 160
rect 4982 151 5304 156
rect 4982 127 5095 151
rect 5119 132 5304 151
rect 5328 132 5341 156
rect 5119 127 5341 132
rect 4982 124 5341 127
rect 5403 124 5438 161
rect 5506 158 5606 161
rect 5506 154 5573 158
rect 5506 128 5518 154
rect 5544 132 5573 154
rect 5599 132 5606 158
rect 5544 128 5606 132
rect 5506 124 5606 128
rect 2432 121 2600 123
rect 2156 95 2600 121
rect 4982 103 5013 124
rect 5403 103 5439 124
rect 4825 102 4862 103
rect 2432 94 2600 95
rect 4824 93 4862 102
rect 4824 73 4833 93
rect 4853 73 4862 93
rect 4824 65 4862 73
rect 4928 97 5013 103
rect 5038 102 5075 103
rect 4928 77 4936 97
rect 4956 77 5013 97
rect 4928 69 5013 77
rect 5037 93 5075 102
rect 5037 73 5046 93
rect 5066 73 5075 93
rect 4928 68 4964 69
rect 5037 65 5075 73
rect 5141 97 5226 103
rect 5246 102 5283 103
rect 5141 77 5149 97
rect 5169 96 5226 97
rect 5169 77 5198 96
rect 5141 76 5198 77
rect 5219 76 5226 96
rect 5141 69 5226 76
rect 5245 93 5283 102
rect 5245 73 5254 93
rect 5274 73 5283 93
rect 5141 68 5177 69
rect 5245 65 5283 73
rect 5349 97 5493 103
rect 5349 77 5357 97
rect 5377 93 5465 97
rect 5377 77 5409 93
rect 5349 76 5409 77
rect 5430 77 5465 93
rect 5485 77 5493 97
rect 5430 76 5493 77
rect 5349 69 5493 76
rect 5349 68 5385 69
rect 5457 68 5493 69
rect 5559 102 5596 103
rect 5559 101 5597 102
rect 5559 93 5623 101
rect 5559 73 5568 93
rect 5588 79 5623 93
rect 5643 79 5646 99
rect 5588 74 5646 79
rect 5588 73 5623 74
rect 4825 36 4862 65
rect 4826 34 4862 36
rect 5038 34 5075 65
rect 4826 12 5075 34
rect 5246 33 5283 65
rect 5559 61 5623 73
rect 5663 35 5690 213
rect 6957 199 7075 219
rect 7095 199 7106 219
rect 6957 191 7106 199
rect 7173 223 7532 227
rect 7173 218 7495 223
rect 7173 194 7286 218
rect 7310 199 7495 218
rect 7519 199 7532 223
rect 7310 194 7532 199
rect 7173 191 7532 194
rect 7594 191 7629 228
rect 7697 225 7797 228
rect 7697 221 7764 225
rect 7697 195 7709 221
rect 7735 199 7764 221
rect 7790 199 7797 225
rect 7735 195 7797 199
rect 7697 191 7797 195
rect 7173 170 7204 191
rect 7594 170 7630 191
rect 7016 169 7053 170
rect 7015 160 7053 169
rect 7015 140 7024 160
rect 7044 140 7053 160
rect 7015 132 7053 140
rect 7119 164 7204 170
rect 7229 169 7266 170
rect 7119 144 7127 164
rect 7147 144 7204 164
rect 7119 136 7204 144
rect 7228 160 7266 169
rect 7228 140 7237 160
rect 7257 140 7266 160
rect 7119 135 7155 136
rect 7228 132 7266 140
rect 7332 164 7417 170
rect 7437 169 7474 170
rect 7332 144 7340 164
rect 7360 163 7417 164
rect 7360 144 7389 163
rect 7332 143 7389 144
rect 7410 143 7417 163
rect 7332 136 7417 143
rect 7436 160 7474 169
rect 7436 140 7445 160
rect 7465 140 7474 160
rect 7332 135 7368 136
rect 7436 132 7474 140
rect 7540 164 7684 170
rect 7540 144 7548 164
rect 7568 163 7656 164
rect 7568 144 7603 163
rect 7540 141 7603 144
rect 7628 144 7656 163
rect 7676 144 7684 164
rect 7628 141 7684 144
rect 7540 136 7684 141
rect 7540 135 7576 136
rect 7648 135 7684 136
rect 7750 169 7787 170
rect 7750 168 7788 169
rect 7750 160 7814 168
rect 7750 140 7759 160
rect 7779 146 7814 160
rect 7834 146 7837 166
rect 7779 141 7837 146
rect 7779 140 7814 141
rect 7016 103 7053 132
rect 7017 101 7053 103
rect 7229 101 7266 132
rect 7017 79 7266 101
rect 7437 100 7474 132
rect 7750 128 7814 140
rect 7854 124 7881 280
rect 10091 235 10128 306
rect 10243 245 10274 246
rect 10091 215 10100 235
rect 10120 215 10128 235
rect 10091 205 10128 215
rect 10187 235 10274 245
rect 10187 215 10196 235
rect 10216 215 10274 235
rect 10187 206 10274 215
rect 10187 205 10224 206
rect 10243 153 10274 206
rect 10304 235 10341 306
rect 10512 311 10905 331
rect 10925 311 10928 331
rect 10512 306 10928 311
rect 12401 318 12410 338
rect 12430 318 12438 338
rect 12401 308 12438 318
rect 12497 338 12584 348
rect 12497 318 12506 338
rect 12526 318 12584 338
rect 12497 309 12584 318
rect 12497 308 12534 309
rect 10512 305 10853 306
rect 10456 245 10487 246
rect 10304 215 10313 235
rect 10333 215 10341 235
rect 10304 205 10341 215
rect 10400 238 10487 245
rect 10400 235 10461 238
rect 10400 215 10409 235
rect 10429 218 10461 235
rect 10482 218 10487 238
rect 10429 215 10487 218
rect 10400 208 10487 215
rect 10512 235 10549 305
rect 10815 304 10852 305
rect 12553 256 12584 309
rect 12614 338 12651 409
rect 12822 414 13215 434
rect 13235 414 13238 434
rect 12822 409 13238 414
rect 12822 408 13163 409
rect 12766 348 12797 349
rect 12614 318 12623 338
rect 12643 318 12651 338
rect 12614 308 12651 318
rect 12710 341 12797 348
rect 12710 338 12771 341
rect 12710 318 12719 338
rect 12739 321 12771 338
rect 12792 321 12797 341
rect 12739 318 12797 321
rect 12710 311 12797 318
rect 12822 338 12859 408
rect 13125 407 13162 408
rect 17682 388 17932 412
rect 12974 348 13010 349
rect 12822 318 12831 338
rect 12851 318 12859 338
rect 12710 309 12766 311
rect 12710 308 12747 309
rect 12822 308 12859 318
rect 12918 338 13066 348
rect 13166 345 13262 347
rect 12918 318 12927 338
rect 12947 318 13037 338
rect 13057 318 13066 338
rect 12918 309 13066 318
rect 13124 344 13262 345
rect 13124 339 13348 344
rect 13124 338 13312 339
rect 13124 318 13133 338
rect 13153 319 13312 338
rect 13340 319 13348 339
rect 13153 318 13348 319
rect 13124 311 13348 318
rect 15491 321 15741 345
rect 13124 309 13262 311
rect 12918 308 12955 309
rect 12974 257 13010 309
rect 13029 308 13066 309
rect 13125 308 13162 309
rect 12445 255 12486 256
rect 12337 248 12486 255
rect 10664 245 10700 246
rect 10512 215 10521 235
rect 10541 215 10549 235
rect 10400 206 10456 208
rect 10400 205 10437 206
rect 10512 205 10549 215
rect 10608 235 10756 245
rect 10856 242 10952 244
rect 10608 215 10617 235
rect 10637 215 10727 235
rect 10747 215 10756 235
rect 10608 206 10756 215
rect 10814 235 10952 242
rect 10814 215 10823 235
rect 10843 215 10952 235
rect 12337 228 12455 248
rect 12475 228 12486 248
rect 12337 220 12486 228
rect 12553 252 12912 256
rect 12553 247 12875 252
rect 12553 223 12666 247
rect 12690 228 12875 247
rect 12899 228 12912 252
rect 12690 223 12912 228
rect 12553 220 12912 223
rect 12974 220 13009 257
rect 13077 254 13177 257
rect 13077 250 13144 254
rect 13077 224 13089 250
rect 13115 228 13144 250
rect 13170 228 13177 254
rect 13115 224 13177 228
rect 13077 220 13177 224
rect 10814 206 10952 215
rect 10608 205 10645 206
rect 10664 154 10700 206
rect 10719 205 10756 206
rect 10815 205 10852 206
rect 10135 152 10176 153
rect 10027 145 10176 152
rect 10027 125 10145 145
rect 10165 125 10176 145
rect 7851 101 7882 124
rect 10027 117 10176 125
rect 10243 149 10602 153
rect 10243 144 10565 149
rect 10243 120 10356 144
rect 10380 125 10565 144
rect 10589 125 10602 149
rect 10380 120 10602 125
rect 10243 117 10602 120
rect 10664 117 10699 154
rect 10767 151 10867 154
rect 10767 147 10834 151
rect 10767 121 10779 147
rect 10805 125 10834 147
rect 10860 125 10867 151
rect 10805 121 10867 125
rect 10767 117 10867 121
rect 7579 100 7882 101
rect 7437 75 7882 100
rect 10243 96 10274 117
rect 10664 96 10700 117
rect 10086 95 10123 96
rect 10085 86 10123 95
rect 7437 74 7622 75
rect 10085 66 10094 86
rect 10114 66 10123 86
rect 10085 58 10123 66
rect 10189 90 10274 96
rect 10299 95 10336 96
rect 10189 70 10197 90
rect 10217 70 10274 90
rect 10189 62 10274 70
rect 10298 86 10336 95
rect 10298 66 10307 86
rect 10327 66 10336 86
rect 10189 61 10225 62
rect 10298 58 10336 66
rect 10402 90 10487 96
rect 10507 95 10544 96
rect 10402 70 10410 90
rect 10430 89 10487 90
rect 10430 70 10459 89
rect 10402 69 10459 70
rect 10480 69 10487 89
rect 10402 62 10487 69
rect 10506 86 10544 95
rect 10506 66 10515 86
rect 10535 66 10544 86
rect 10402 61 10438 62
rect 10506 58 10544 66
rect 10610 91 10754 96
rect 10610 90 10668 91
rect 10610 70 10618 90
rect 10638 70 10668 90
rect 10610 68 10668 70
rect 10696 90 10754 91
rect 10696 70 10726 90
rect 10746 70 10754 90
rect 10696 68 10754 70
rect 10610 62 10754 68
rect 10610 61 10646 62
rect 10718 61 10754 62
rect 10820 95 10857 96
rect 10820 94 10858 95
rect 10820 86 10884 94
rect 10820 66 10829 86
rect 10849 72 10884 86
rect 10904 72 10907 92
rect 10849 67 10907 72
rect 10849 66 10884 67
rect 5522 33 5690 35
rect 5246 26 5690 33
rect 10086 29 10123 58
rect 5246 9 5659 26
rect 5683 9 5690 26
rect 5246 7 5690 9
rect 5522 6 5690 7
rect 10087 27 10123 29
rect 10299 27 10336 58
rect 10087 5 10336 27
rect 10507 26 10544 58
rect 10820 54 10884 66
rect 10924 36 10951 206
rect 12553 199 12584 220
rect 12974 199 13010 220
rect 12396 198 12433 199
rect 12395 189 12433 198
rect 12395 169 12404 189
rect 12424 169 12433 189
rect 12395 161 12433 169
rect 12499 193 12584 199
rect 12609 198 12646 199
rect 12499 173 12507 193
rect 12527 173 12584 193
rect 12499 165 12584 173
rect 12608 189 12646 198
rect 12608 169 12617 189
rect 12637 169 12646 189
rect 12499 164 12535 165
rect 12608 161 12646 169
rect 12712 193 12797 199
rect 12817 198 12854 199
rect 12712 173 12720 193
rect 12740 192 12797 193
rect 12740 173 12769 192
rect 12712 172 12769 173
rect 12790 172 12797 192
rect 12712 165 12797 172
rect 12816 189 12854 198
rect 12816 169 12825 189
rect 12845 169 12854 189
rect 12712 164 12748 165
rect 12816 161 12854 169
rect 12920 193 13064 199
rect 12920 173 12928 193
rect 12948 192 13036 193
rect 12948 173 12983 192
rect 12920 170 12983 173
rect 13008 173 13036 192
rect 13056 173 13064 193
rect 13008 170 13064 173
rect 12920 165 13064 170
rect 12920 164 12956 165
rect 13028 164 13064 165
rect 13130 198 13167 199
rect 13130 197 13168 198
rect 13130 189 13194 197
rect 13130 169 13139 189
rect 13159 175 13194 189
rect 13214 175 13217 195
rect 13159 170 13217 175
rect 13159 169 13194 170
rect 12396 132 12433 161
rect 12397 130 12433 132
rect 12609 130 12646 161
rect 12397 108 12646 130
rect 12817 129 12854 161
rect 13130 157 13194 169
rect 13234 131 13261 309
rect 15491 250 15528 321
rect 15643 260 15674 261
rect 15491 230 15500 250
rect 15520 230 15528 250
rect 15491 220 15528 230
rect 15587 250 15674 260
rect 15587 230 15596 250
rect 15616 230 15674 250
rect 15587 221 15674 230
rect 15587 220 15624 221
rect 15643 168 15674 221
rect 15704 250 15741 321
rect 15912 326 16305 346
rect 16325 326 16328 346
rect 15912 321 16328 326
rect 15912 320 16253 321
rect 15856 260 15887 261
rect 15704 230 15713 250
rect 15733 230 15741 250
rect 15704 220 15741 230
rect 15800 253 15887 260
rect 15800 250 15861 253
rect 15800 230 15809 250
rect 15829 233 15861 250
rect 15882 233 15887 253
rect 15829 230 15887 233
rect 15800 223 15887 230
rect 15912 250 15949 320
rect 16215 319 16252 320
rect 17682 317 17719 388
rect 17834 327 17865 328
rect 17682 297 17691 317
rect 17711 297 17719 317
rect 17682 287 17719 297
rect 17778 317 17865 327
rect 17778 297 17787 317
rect 17807 297 17865 317
rect 17778 288 17865 297
rect 17778 287 17815 288
rect 16064 260 16100 261
rect 15912 230 15921 250
rect 15941 230 15949 250
rect 15800 221 15856 223
rect 15800 220 15837 221
rect 15912 220 15949 230
rect 16008 250 16156 260
rect 16256 257 16352 259
rect 16008 230 16017 250
rect 16037 230 16127 250
rect 16147 230 16156 250
rect 16008 221 16156 230
rect 16214 250 16352 257
rect 16214 230 16223 250
rect 16243 230 16352 250
rect 17834 235 17865 288
rect 17895 317 17932 388
rect 18103 393 18496 413
rect 18516 393 18519 413
rect 18103 388 18519 393
rect 18103 387 18444 388
rect 18047 327 18078 328
rect 17895 297 17904 317
rect 17924 297 17932 317
rect 17895 287 17932 297
rect 17991 320 18078 327
rect 17991 317 18052 320
rect 17991 297 18000 317
rect 18020 300 18052 317
rect 18073 300 18078 320
rect 18020 297 18078 300
rect 17991 290 18078 297
rect 18103 317 18140 387
rect 18406 386 18443 387
rect 18255 327 18291 328
rect 18103 297 18112 317
rect 18132 297 18140 317
rect 17991 288 18047 290
rect 17991 287 18028 288
rect 18103 287 18140 297
rect 18199 317 18347 327
rect 18447 324 18543 326
rect 18199 297 18208 317
rect 18228 297 18318 317
rect 18338 297 18347 317
rect 18199 288 18347 297
rect 18405 323 18543 324
rect 18405 318 18629 323
rect 18405 317 18593 318
rect 18405 297 18414 317
rect 18434 298 18593 317
rect 18621 298 18629 318
rect 18434 297 18629 298
rect 18405 290 18629 297
rect 18405 288 18543 290
rect 18199 287 18236 288
rect 18255 236 18291 288
rect 18310 287 18347 288
rect 18406 287 18443 288
rect 17726 234 17767 235
rect 16214 221 16352 230
rect 17618 227 17767 234
rect 16008 220 16045 221
rect 16064 169 16100 221
rect 16119 220 16156 221
rect 16215 220 16252 221
rect 15535 167 15576 168
rect 15427 160 15576 167
rect 15427 140 15545 160
rect 15565 140 15576 160
rect 15427 132 15576 140
rect 15643 164 16002 168
rect 15643 159 15965 164
rect 15643 135 15756 159
rect 15780 140 15965 159
rect 15989 140 16002 164
rect 15780 135 16002 140
rect 15643 132 16002 135
rect 16064 132 16099 169
rect 16167 166 16267 169
rect 16167 162 16234 166
rect 16167 136 16179 162
rect 16205 140 16234 162
rect 16260 140 16267 166
rect 16205 136 16267 140
rect 16167 132 16267 136
rect 13093 129 13261 131
rect 12817 103 13261 129
rect 15643 111 15674 132
rect 16064 111 16100 132
rect 15486 110 15523 111
rect 13093 102 13261 103
rect 15485 101 15523 110
rect 15485 81 15494 101
rect 15514 81 15523 101
rect 15485 73 15523 81
rect 15589 105 15674 111
rect 15699 110 15736 111
rect 15589 85 15597 105
rect 15617 85 15674 105
rect 15589 77 15674 85
rect 15698 101 15736 110
rect 15698 81 15707 101
rect 15727 81 15736 101
rect 15589 76 15625 77
rect 15698 73 15736 81
rect 15802 105 15887 111
rect 15907 110 15944 111
rect 15802 85 15810 105
rect 15830 104 15887 105
rect 15830 85 15859 104
rect 15802 84 15859 85
rect 15880 84 15887 104
rect 15802 77 15887 84
rect 15906 101 15944 110
rect 15906 81 15915 101
rect 15935 81 15944 101
rect 15802 76 15838 77
rect 15906 73 15944 81
rect 16010 105 16154 111
rect 16010 85 16018 105
rect 16038 101 16126 105
rect 16038 85 16070 101
rect 16010 84 16070 85
rect 16091 85 16126 101
rect 16146 85 16154 105
rect 16091 84 16154 85
rect 16010 77 16154 84
rect 16010 76 16046 77
rect 16118 76 16154 77
rect 16220 110 16257 111
rect 16220 109 16258 110
rect 16220 101 16284 109
rect 16220 81 16229 101
rect 16249 87 16284 101
rect 16304 87 16307 107
rect 16249 82 16307 87
rect 16249 81 16284 82
rect 15486 44 15523 73
rect 10921 28 10951 36
rect 10783 26 10951 28
rect 10507 0 10951 26
rect 15487 42 15523 44
rect 15699 42 15736 73
rect 15487 20 15736 42
rect 15907 41 15944 73
rect 16220 69 16284 81
rect 16324 43 16351 221
rect 17618 207 17736 227
rect 17756 207 17767 227
rect 17618 199 17767 207
rect 17834 231 18193 235
rect 17834 226 18156 231
rect 17834 202 17947 226
rect 17971 207 18156 226
rect 18180 207 18193 231
rect 17971 202 18193 207
rect 17834 199 18193 202
rect 18255 199 18290 236
rect 18358 233 18458 236
rect 18358 229 18425 233
rect 18358 203 18370 229
rect 18396 207 18425 229
rect 18451 207 18458 233
rect 18396 203 18458 207
rect 18358 199 18458 203
rect 17834 178 17865 199
rect 18255 178 18291 199
rect 17677 177 17714 178
rect 17676 168 17714 177
rect 17676 148 17685 168
rect 17705 148 17714 168
rect 17676 140 17714 148
rect 17780 172 17865 178
rect 17890 177 17927 178
rect 17780 152 17788 172
rect 17808 152 17865 172
rect 17780 144 17865 152
rect 17889 168 17927 177
rect 17889 148 17898 168
rect 17918 148 17927 168
rect 17780 143 17816 144
rect 17889 140 17927 148
rect 17993 172 18078 178
rect 18098 177 18135 178
rect 17993 152 18001 172
rect 18021 171 18078 172
rect 18021 152 18050 171
rect 17993 151 18050 152
rect 18071 151 18078 171
rect 17993 144 18078 151
rect 18097 168 18135 177
rect 18097 148 18106 168
rect 18126 148 18135 168
rect 17993 143 18029 144
rect 18097 140 18135 148
rect 18201 172 18345 178
rect 18201 152 18209 172
rect 18229 171 18317 172
rect 18229 152 18264 171
rect 18201 149 18264 152
rect 18289 152 18317 171
rect 18337 152 18345 172
rect 18289 149 18345 152
rect 18201 144 18345 149
rect 18201 143 18237 144
rect 18309 143 18345 144
rect 18411 177 18448 178
rect 18411 176 18449 177
rect 18411 168 18475 176
rect 18411 148 18420 168
rect 18440 154 18475 168
rect 18495 154 18498 174
rect 18440 149 18498 154
rect 18440 148 18475 149
rect 17677 111 17714 140
rect 17678 109 17714 111
rect 17890 109 17927 140
rect 17678 87 17927 109
rect 18098 108 18135 140
rect 18411 136 18475 148
rect 18515 132 18542 288
rect 18512 109 18543 132
rect 18240 108 18543 109
rect 18098 83 18543 108
rect 18098 82 18283 83
rect 16183 41 16351 43
rect 15907 34 16351 41
rect 15907 17 16320 34
rect 16344 17 16351 34
rect 15907 15 16351 17
rect 16183 14 16351 15
rect 10783 -1 10951 0
rect 10921 -24 10951 -1
rect 10921 -45 10925 -24
rect 10945 -45 10951 -24
rect 10921 -52 10951 -45
<< viali >>
rect 1115 8160 1135 8180
rect 671 8067 692 8087
rect 4078 8241 4098 8261
rect 4294 8244 4316 8265
rect 4502 8244 4523 8264
rect 4122 8182 4148 8208
rect 2973 8074 2992 8100
rect 1044 7974 1070 8000
rect 669 7918 690 7938
rect 885 7919 907 7940
rect 1094 7921 1114 7941
rect 2127 7979 2147 7999
rect 1683 7886 1704 7906
rect 2056 7793 2082 7819
rect 1114 7745 1134 7765
rect 670 7652 691 7672
rect 1681 7737 1702 7757
rect 1892 7738 1916 7758
rect 2106 7740 2126 7760
rect 1778 7671 1798 7690
rect 2880 7658 2900 7676
rect 3393 8077 3413 8096
rect 3065 8007 3085 8027
rect 3276 8008 3300 8028
rect 3489 8010 3510 8030
rect 4500 8095 4521 8115
rect 4057 8002 4077 8022
rect 3109 7948 3135 7974
rect 3487 7861 3508 7881
rect 3044 7768 3064 7788
rect 6396 8139 6416 8159
rect 5952 8046 5973 8066
rect 9359 8220 9379 8240
rect 9575 8223 9597 8244
rect 9783 8223 9804 8243
rect 9403 8161 9429 8187
rect 8254 8053 8273 8079
rect 4077 7826 4097 7846
rect 4284 7827 4306 7848
rect 4501 7829 4522 7849
rect 4121 7767 4147 7793
rect 6325 7953 6351 7979
rect 5950 7897 5971 7917
rect 6166 7898 6188 7919
rect 6375 7900 6395 7920
rect 1043 7559 1069 7585
rect 668 7503 689 7523
rect 875 7502 897 7523
rect 1093 7506 1113 7526
rect 2182 7418 2202 7438
rect 1738 7325 1759 7345
rect 2111 7232 2137 7258
rect 1120 7179 1140 7199
rect 676 7086 697 7106
rect 1736 7176 1757 7196
rect 1951 7178 1975 7195
rect 2161 7179 2181 7199
rect 1049 6993 1075 7019
rect 674 6937 695 6957
rect 890 6938 912 6959
rect 1099 6940 1119 6960
rect 2132 6998 2152 7018
rect 1688 6905 1709 6925
rect 2061 6812 2087 6838
rect 1119 6764 1139 6784
rect 675 6671 696 6691
rect 1686 6756 1707 6776
rect 1896 6758 1920 6778
rect 2111 6759 2131 6779
rect 1783 6690 1803 6709
rect 2204 6686 2223 6712
rect 1048 6578 1074 6604
rect 673 6522 694 6542
rect 880 6521 902 6542
rect 1098 6525 1118 6545
rect 3015 7587 3035 7607
rect 3225 7590 3248 7609
rect 3439 7590 3460 7610
rect 4499 7680 4520 7700
rect 4056 7587 4076 7607
rect 7408 7958 7428 7978
rect 6964 7865 6985 7885
rect 7337 7772 7363 7798
rect 3059 7528 3085 7554
rect 6395 7724 6415 7744
rect 5951 7631 5972 7651
rect 6962 7716 6983 7736
rect 7173 7717 7197 7737
rect 7387 7719 7407 7739
rect 7059 7650 7079 7669
rect 8161 7637 8181 7655
rect 8674 8056 8694 8075
rect 8346 7986 8366 8006
rect 8557 7987 8581 8007
rect 8770 7989 8791 8009
rect 9781 8074 9802 8094
rect 9338 7981 9358 8001
rect 8390 7927 8416 7953
rect 11776 8168 11796 8188
rect 11332 8075 11353 8095
rect 14739 8249 14759 8269
rect 14955 8252 14977 8273
rect 15163 8252 15184 8272
rect 14783 8190 14809 8216
rect 13634 8082 13653 8108
rect 8768 7840 8789 7860
rect 8325 7747 8345 7767
rect 9358 7805 9378 7825
rect 9565 7806 9587 7827
rect 9782 7808 9803 7828
rect 9402 7746 9428 7772
rect 11705 7982 11731 8008
rect 11330 7926 11351 7946
rect 11546 7927 11568 7948
rect 11755 7929 11775 7949
rect 12788 7987 12808 8007
rect 12344 7894 12365 7914
rect 6324 7538 6350 7564
rect 3437 7441 3458 7461
rect 2994 7348 3014 7368
rect 5949 7482 5970 7502
rect 6156 7481 6178 7502
rect 6374 7485 6394 7505
rect 4083 7260 4103 7280
rect 4299 7263 4321 7284
rect 4507 7263 4528 7283
rect 7463 7397 7483 7417
rect 7019 7304 7040 7324
rect 4127 7201 4153 7227
rect 3398 7096 3418 7115
rect 3070 7026 3090 7046
rect 3280 7028 3304 7048
rect 3494 7029 3515 7049
rect 4505 7114 4526 7134
rect 4062 7021 4082 7041
rect 7392 7211 7418 7237
rect 3114 6967 3140 6993
rect 3492 6880 3513 6900
rect 3049 6787 3069 6807
rect 6401 7158 6421 7178
rect 5957 7065 5978 7085
rect 7017 7155 7038 7175
rect 7232 7157 7256 7174
rect 7442 7158 7462 7178
rect 4082 6845 4102 6865
rect 4289 6846 4311 6867
rect 4506 6848 4527 6868
rect 4126 6786 4152 6812
rect 6330 6972 6356 6998
rect 5955 6916 5976 6936
rect 6171 6917 6193 6938
rect 6380 6919 6400 6939
rect 2757 6629 2780 6648
rect 2347 6486 2367 6506
rect 1903 6393 1924 6413
rect 2276 6300 2302 6326
rect 1901 6244 1922 6264
rect 2110 6243 2135 6269
rect 2326 6247 2346 6267
rect 1127 6200 1147 6220
rect 683 6107 704 6127
rect 1056 6014 1082 6040
rect 681 5958 702 5978
rect 897 5959 919 5980
rect 1106 5961 1126 5981
rect 2139 6019 2159 6039
rect 1695 5926 1716 5946
rect 2068 5833 2094 5859
rect 1126 5785 1146 5805
rect 682 5692 703 5712
rect 1693 5777 1714 5797
rect 1904 5778 1928 5798
rect 2118 5780 2138 5800
rect 1790 5711 1810 5730
rect 1055 5599 1081 5625
rect 680 5543 701 5563
rect 887 5542 909 5563
rect 1105 5546 1125 5566
rect 2194 5458 2214 5478
rect 1750 5365 1771 5385
rect 2123 5272 2149 5298
rect 1132 5219 1152 5239
rect 688 5126 709 5146
rect 1748 5216 1769 5236
rect 1960 5217 1983 5236
rect 2173 5219 2193 5239
rect 1061 5033 1087 5059
rect 686 4977 707 4997
rect 902 4978 924 4999
rect 1111 4980 1131 5000
rect 2144 5038 2164 5058
rect 1700 4945 1721 4965
rect 2073 4852 2099 4878
rect 1131 4804 1151 4824
rect 687 4711 708 4731
rect 1698 4796 1719 4816
rect 1908 4798 1932 4818
rect 2123 4799 2143 4819
rect 1795 4730 1815 4749
rect 2308 5150 2328 5168
rect 2216 4726 2235 4752
rect 4504 6699 4525 6719
rect 4061 6606 4081 6626
rect 7413 6977 7433 6997
rect 6969 6884 6990 6904
rect 7342 6791 7368 6817
rect 2862 6559 2882 6579
rect 3069 6561 3092 6580
rect 3286 6562 3307 6582
rect 6400 6743 6420 6763
rect 5956 6650 5977 6670
rect 6967 6735 6988 6755
rect 7177 6737 7201 6757
rect 7392 6738 7412 6758
rect 7064 6669 7084 6688
rect 7485 6665 7504 6691
rect 6329 6557 6355 6583
rect 2906 6500 2932 6526
rect 3284 6413 3305 6433
rect 2841 6320 2861 6340
rect 5954 6501 5975 6521
rect 6161 6500 6183 6521
rect 6379 6504 6399 6524
rect 8296 7566 8316 7586
rect 8506 7569 8529 7588
rect 8720 7569 8741 7589
rect 9780 7659 9801 7679
rect 9337 7566 9357 7586
rect 12717 7801 12743 7827
rect 11775 7753 11795 7773
rect 11331 7660 11352 7680
rect 12342 7745 12363 7765
rect 12553 7746 12577 7766
rect 12767 7748 12787 7768
rect 12439 7679 12459 7698
rect 13541 7666 13561 7684
rect 14054 8085 14074 8104
rect 13726 8015 13746 8035
rect 13937 8016 13961 8036
rect 14150 8018 14171 8038
rect 15161 8103 15182 8123
rect 14718 8010 14738 8030
rect 13770 7956 13796 7982
rect 14148 7869 14169 7889
rect 13705 7776 13725 7796
rect 17057 8147 17077 8167
rect 16613 8054 16634 8074
rect 20020 8228 20040 8248
rect 20236 8231 20258 8252
rect 20444 8231 20465 8251
rect 20064 8169 20090 8195
rect 18915 8061 18934 8087
rect 14738 7834 14758 7854
rect 14945 7835 14967 7856
rect 15162 7837 15183 7857
rect 14782 7775 14808 7801
rect 16986 7961 17012 7987
rect 16611 7905 16632 7925
rect 16827 7906 16849 7927
rect 17036 7908 17056 7928
rect 11704 7567 11730 7593
rect 8340 7507 8366 7533
rect 8718 7420 8739 7440
rect 8275 7327 8295 7347
rect 11329 7511 11350 7531
rect 11536 7510 11558 7531
rect 11754 7514 11774 7534
rect 9364 7239 9384 7259
rect 9580 7242 9602 7263
rect 9788 7242 9809 7262
rect 12843 7426 12863 7446
rect 12399 7333 12420 7353
rect 12772 7240 12798 7266
rect 9408 7180 9434 7206
rect 8679 7075 8699 7094
rect 8351 7005 8371 7025
rect 8561 7007 8585 7027
rect 8775 7008 8796 7028
rect 9786 7093 9807 7113
rect 9343 7000 9363 7020
rect 8395 6946 8421 6972
rect 11781 7187 11801 7207
rect 11337 7094 11358 7114
rect 12397 7184 12418 7204
rect 12612 7186 12636 7203
rect 12822 7187 12842 7207
rect 8773 6859 8794 6879
rect 8330 6766 8350 6786
rect 9363 6824 9383 6844
rect 9570 6825 9592 6846
rect 9787 6827 9808 6847
rect 9407 6765 9433 6791
rect 11710 7001 11736 7027
rect 11335 6945 11356 6965
rect 11551 6946 11573 6967
rect 11760 6948 11780 6968
rect 12793 7006 12813 7026
rect 12349 6913 12370 6933
rect 8038 6608 8061 6627
rect 4090 6281 4110 6301
rect 4306 6284 4328 6305
rect 4514 6284 4535 6304
rect 7628 6465 7648 6485
rect 7184 6372 7205 6392
rect 7557 6279 7583 6305
rect 4134 6222 4160 6248
rect 2985 6114 3004 6140
rect 3405 6117 3425 6136
rect 3077 6047 3097 6067
rect 3288 6048 3312 6068
rect 3501 6050 3522 6070
rect 4512 6135 4533 6155
rect 4069 6042 4089 6062
rect 7182 6223 7203 6243
rect 7391 6222 7416 6248
rect 7607 6226 7627 6246
rect 3121 5988 3147 6014
rect 3499 5901 3520 5921
rect 3056 5808 3076 5828
rect 6408 6179 6428 6199
rect 5964 6086 5985 6106
rect 4089 5866 4109 5886
rect 4296 5867 4318 5888
rect 4513 5869 4534 5889
rect 4133 5807 4159 5833
rect 6337 5993 6363 6019
rect 5962 5937 5983 5957
rect 6178 5938 6200 5959
rect 6387 5940 6407 5960
rect 3027 5627 3047 5647
rect 3233 5631 3257 5648
rect 3451 5630 3472 5650
rect 4511 5720 4532 5740
rect 4068 5627 4088 5647
rect 7420 5998 7440 6018
rect 6976 5905 6997 5925
rect 7349 5812 7375 5838
rect 3071 5568 3097 5594
rect 6407 5764 6427 5784
rect 5963 5671 5984 5691
rect 6974 5756 6995 5776
rect 7185 5757 7209 5777
rect 7399 5759 7419 5779
rect 7071 5690 7091 5709
rect 6336 5578 6362 5604
rect 3449 5481 3470 5501
rect 3006 5388 3026 5408
rect 5961 5522 5982 5542
rect 6168 5521 6190 5542
rect 6386 5525 6406 5545
rect 4095 5300 4115 5320
rect 4311 5303 4333 5324
rect 4519 5303 4540 5323
rect 7475 5437 7495 5457
rect 7031 5344 7052 5364
rect 4139 5241 4165 5267
rect 3410 5136 3430 5155
rect 3082 5066 3102 5086
rect 3292 5068 3316 5088
rect 3506 5069 3527 5089
rect 4517 5154 4538 5174
rect 4074 5061 4094 5081
rect 7404 5251 7430 5277
rect 3126 5007 3152 5033
rect 3504 4920 3525 4940
rect 3061 4827 3081 4847
rect 6413 5198 6433 5218
rect 5969 5105 5990 5125
rect 7029 5195 7050 5215
rect 7241 5196 7264 5215
rect 7454 5198 7474 5218
rect 4094 4885 4114 4905
rect 4301 4886 4323 4907
rect 4518 4888 4539 4908
rect 4138 4826 4164 4852
rect 6342 5012 6368 5038
rect 5967 4956 5988 4976
rect 6183 4957 6205 4978
rect 6392 4959 6412 4979
rect 1060 4618 1086 4644
rect 685 4562 706 4582
rect 892 4561 914 4582
rect 1110 4565 1130 4585
rect 4516 4739 4537 4759
rect 2787 4634 2807 4654
rect 2991 4635 3017 4654
rect 3211 4637 3232 4657
rect 4073 4646 4093 4666
rect 7425 5017 7445 5037
rect 6981 4924 7002 4944
rect 7354 4831 7380 4857
rect 2831 4575 2857 4601
rect 6412 4783 6432 4803
rect 5968 4690 5989 4710
rect 6979 4775 7000 4795
rect 7189 4777 7213 4797
rect 7404 4778 7424 4798
rect 7076 4709 7096 4728
rect 7589 5129 7609 5147
rect 7497 4705 7516 4731
rect 9785 6678 9806 6698
rect 9342 6585 9362 6605
rect 12722 6820 12748 6846
rect 8143 6538 8163 6558
rect 8350 6540 8373 6559
rect 8567 6541 8588 6561
rect 11780 6772 11800 6792
rect 11336 6679 11357 6699
rect 12347 6764 12368 6784
rect 12557 6766 12581 6786
rect 12772 6767 12792 6787
rect 12444 6698 12464 6717
rect 12865 6694 12884 6720
rect 11709 6586 11735 6612
rect 8187 6479 8213 6505
rect 11334 6530 11355 6550
rect 11541 6529 11563 6550
rect 11759 6533 11779 6553
rect 8565 6392 8586 6412
rect 8122 6299 8142 6319
rect 13676 7595 13696 7615
rect 13886 7598 13909 7617
rect 14100 7598 14121 7618
rect 15160 7688 15181 7708
rect 14717 7595 14737 7615
rect 18069 7966 18089 7986
rect 17625 7873 17646 7893
rect 17998 7780 18024 7806
rect 13720 7536 13746 7562
rect 17056 7732 17076 7752
rect 16612 7639 16633 7659
rect 17623 7724 17644 7744
rect 17834 7725 17858 7745
rect 18048 7727 18068 7747
rect 17720 7658 17740 7677
rect 18822 7645 18842 7663
rect 19335 8064 19355 8083
rect 19007 7994 19027 8014
rect 19218 7995 19242 8015
rect 19431 7997 19452 8017
rect 20442 8082 20463 8102
rect 19999 7989 20019 8009
rect 19051 7935 19077 7961
rect 19429 7848 19450 7868
rect 18986 7755 19006 7775
rect 20019 7813 20039 7833
rect 20226 7814 20248 7835
rect 20443 7816 20464 7836
rect 20063 7754 20089 7780
rect 16985 7546 17011 7572
rect 14098 7449 14119 7469
rect 13655 7356 13675 7376
rect 16610 7490 16631 7510
rect 16817 7489 16839 7510
rect 17035 7493 17055 7513
rect 14744 7268 14764 7288
rect 14960 7271 14982 7292
rect 15168 7271 15189 7291
rect 18124 7405 18144 7425
rect 17680 7312 17701 7332
rect 14788 7209 14814 7235
rect 14059 7104 14079 7123
rect 13731 7034 13751 7054
rect 13941 7036 13965 7056
rect 14155 7037 14176 7057
rect 15166 7122 15187 7142
rect 14723 7029 14743 7049
rect 18053 7219 18079 7245
rect 13775 6975 13801 7001
rect 14153 6888 14174 6908
rect 13710 6795 13730 6815
rect 17062 7166 17082 7186
rect 16618 7073 16639 7093
rect 17678 7163 17699 7183
rect 17893 7165 17917 7182
rect 18103 7166 18123 7186
rect 14743 6853 14763 6873
rect 14950 6854 14972 6875
rect 15167 6856 15188 6876
rect 14787 6794 14813 6820
rect 16991 6980 17017 7006
rect 16616 6924 16637 6944
rect 16832 6925 16854 6946
rect 17041 6927 17061 6947
rect 13418 6637 13441 6656
rect 13008 6494 13028 6514
rect 12564 6401 12585 6421
rect 9371 6260 9391 6280
rect 9587 6263 9609 6284
rect 9795 6263 9816 6283
rect 12937 6308 12963 6334
rect 9415 6201 9441 6227
rect 8266 6093 8285 6119
rect 8686 6096 8706 6115
rect 8358 6026 8378 6046
rect 8569 6027 8593 6047
rect 8782 6029 8803 6049
rect 9793 6114 9814 6134
rect 9350 6021 9370 6041
rect 12562 6252 12583 6272
rect 12771 6251 12796 6277
rect 12987 6255 13007 6275
rect 8402 5967 8428 5993
rect 11788 6208 11808 6228
rect 11344 6115 11365 6135
rect 8780 5880 8801 5900
rect 8337 5787 8357 5807
rect 9370 5845 9390 5865
rect 9577 5846 9599 5867
rect 9794 5848 9815 5868
rect 9414 5786 9440 5812
rect 11717 6022 11743 6048
rect 11342 5966 11363 5986
rect 11558 5967 11580 5988
rect 11767 5969 11787 5989
rect 12800 6027 12820 6047
rect 12356 5934 12377 5954
rect 8308 5606 8328 5626
rect 8514 5610 8538 5627
rect 8732 5609 8753 5629
rect 9792 5699 9813 5719
rect 9349 5606 9369 5626
rect 12729 5841 12755 5867
rect 11787 5793 11807 5813
rect 11343 5700 11364 5720
rect 12354 5785 12375 5805
rect 12565 5786 12589 5806
rect 12779 5788 12799 5808
rect 12451 5719 12471 5738
rect 11716 5607 11742 5633
rect 8352 5547 8378 5573
rect 8730 5460 8751 5480
rect 8287 5367 8307 5387
rect 11341 5551 11362 5571
rect 11548 5550 11570 5571
rect 11766 5554 11786 5574
rect 9376 5279 9396 5299
rect 9592 5282 9614 5303
rect 9800 5282 9821 5302
rect 12855 5466 12875 5486
rect 12411 5373 12432 5393
rect 12784 5280 12810 5306
rect 9420 5220 9446 5246
rect 8691 5115 8711 5134
rect 8363 5045 8383 5065
rect 8573 5047 8597 5067
rect 8787 5048 8808 5068
rect 9798 5133 9819 5153
rect 9355 5040 9375 5060
rect 8407 4986 8433 5012
rect 11793 5227 11813 5247
rect 11349 5134 11370 5154
rect 12409 5224 12430 5244
rect 12621 5225 12644 5244
rect 12834 5227 12854 5247
rect 8785 4899 8806 4919
rect 8342 4806 8362 4826
rect 9375 4864 9395 4884
rect 9582 4865 9604 4886
rect 9799 4867 9820 4887
rect 9419 4805 9445 4831
rect 11722 5041 11748 5067
rect 11347 4985 11368 5005
rect 11563 4986 11585 5007
rect 11772 4988 11792 5008
rect 12805 5046 12825 5066
rect 12361 4953 12382 4973
rect 6341 4597 6367 4623
rect 2442 4494 2462 4514
rect 1998 4401 2019 4421
rect 3209 4488 3230 4508
rect 2766 4395 2786 4415
rect 5966 4541 5987 4561
rect 6173 4540 6195 4561
rect 6391 4544 6411 4564
rect 9797 4718 9818 4738
rect 8068 4613 8088 4633
rect 8272 4614 8298 4633
rect 8492 4616 8513 4636
rect 9354 4625 9374 4645
rect 12734 4860 12760 4886
rect 11792 4812 11812 4832
rect 11348 4719 11369 4739
rect 12359 4804 12380 4824
rect 12569 4806 12593 4826
rect 12784 4807 12804 4827
rect 12456 4738 12476 4757
rect 12969 5158 12989 5176
rect 12877 4734 12896 4760
rect 15165 6707 15186 6727
rect 14722 6614 14742 6634
rect 18074 6985 18094 7005
rect 17630 6892 17651 6912
rect 18003 6799 18029 6825
rect 13523 6567 13543 6587
rect 13730 6569 13753 6588
rect 13947 6570 13968 6590
rect 17061 6751 17081 6771
rect 16617 6658 16638 6678
rect 17628 6743 17649 6763
rect 17838 6745 17862 6765
rect 18053 6746 18073 6766
rect 17725 6677 17745 6696
rect 18146 6673 18165 6699
rect 16990 6565 17016 6591
rect 13567 6508 13593 6534
rect 13945 6421 13966 6441
rect 13502 6328 13522 6348
rect 16615 6509 16636 6529
rect 16822 6508 16844 6529
rect 17040 6512 17060 6532
rect 18957 7574 18977 7594
rect 19167 7577 19190 7596
rect 19381 7577 19402 7597
rect 20441 7667 20462 7687
rect 19998 7574 20018 7594
rect 19001 7515 19027 7541
rect 19379 7428 19400 7448
rect 18936 7335 18956 7355
rect 20025 7247 20045 7267
rect 20241 7250 20263 7271
rect 20449 7250 20470 7270
rect 20069 7188 20095 7214
rect 19340 7083 19360 7102
rect 19012 7013 19032 7033
rect 19222 7015 19246 7035
rect 19436 7016 19457 7036
rect 20447 7101 20468 7121
rect 20004 7008 20024 7028
rect 19056 6954 19082 6980
rect 19434 6867 19455 6887
rect 18991 6774 19011 6794
rect 20024 6832 20044 6852
rect 20231 6833 20253 6854
rect 20448 6835 20469 6855
rect 20068 6773 20094 6799
rect 18699 6616 18722 6635
rect 14751 6289 14771 6309
rect 14967 6292 14989 6313
rect 15175 6292 15196 6312
rect 18289 6473 18309 6493
rect 17845 6380 17866 6400
rect 18218 6287 18244 6313
rect 14795 6230 14821 6256
rect 13646 6122 13665 6148
rect 14066 6125 14086 6144
rect 13738 6055 13758 6075
rect 13949 6056 13973 6076
rect 14162 6058 14183 6078
rect 15173 6143 15194 6163
rect 14730 6050 14750 6070
rect 17843 6231 17864 6251
rect 18052 6230 18077 6256
rect 18268 6234 18288 6254
rect 13782 5996 13808 6022
rect 14160 5909 14181 5929
rect 13717 5816 13737 5836
rect 17069 6187 17089 6207
rect 16625 6094 16646 6114
rect 14750 5874 14770 5894
rect 14957 5875 14979 5896
rect 15174 5877 15195 5897
rect 14794 5815 14820 5841
rect 16998 6001 17024 6027
rect 16623 5945 16644 5965
rect 16839 5946 16861 5967
rect 17048 5948 17068 5968
rect 13688 5635 13708 5655
rect 13894 5639 13918 5656
rect 14112 5638 14133 5658
rect 15172 5728 15193 5748
rect 14729 5635 14749 5655
rect 18081 6006 18101 6026
rect 17637 5913 17658 5933
rect 18010 5820 18036 5846
rect 13732 5576 13758 5602
rect 17068 5772 17088 5792
rect 16624 5679 16645 5699
rect 17635 5764 17656 5784
rect 17846 5765 17870 5785
rect 18060 5767 18080 5787
rect 17732 5698 17752 5717
rect 16997 5586 17023 5612
rect 14110 5489 14131 5509
rect 13667 5396 13687 5416
rect 16622 5530 16643 5550
rect 16829 5529 16851 5550
rect 17047 5533 17067 5553
rect 14756 5308 14776 5328
rect 14972 5311 14994 5332
rect 15180 5311 15201 5331
rect 18136 5445 18156 5465
rect 17692 5352 17713 5372
rect 14800 5249 14826 5275
rect 14071 5144 14091 5163
rect 13743 5074 13763 5094
rect 13953 5076 13977 5096
rect 14167 5077 14188 5097
rect 15178 5162 15199 5182
rect 14735 5069 14755 5089
rect 18065 5259 18091 5285
rect 13787 5015 13813 5041
rect 14165 4928 14186 4948
rect 13722 4835 13742 4855
rect 17074 5206 17094 5226
rect 16630 5113 16651 5133
rect 17690 5203 17711 5223
rect 17902 5204 17925 5223
rect 18115 5206 18135 5226
rect 14755 4893 14775 4913
rect 14962 4894 14984 4915
rect 15179 4896 15200 4916
rect 14799 4834 14825 4860
rect 17003 5020 17029 5046
rect 16628 4964 16649 4984
rect 16844 4965 16866 4986
rect 17053 4967 17073 4987
rect 11721 4626 11747 4652
rect 8112 4554 8138 4580
rect 2371 4308 2397 4334
rect 1135 4243 1155 4263
rect 1996 4252 2017 4272
rect 2211 4255 2237 4274
rect 2421 4255 2441 4275
rect 691 4150 712 4170
rect 4098 4324 4118 4344
rect 4314 4327 4336 4348
rect 4522 4327 4543 4347
rect 7723 4473 7743 4493
rect 7279 4380 7300 4400
rect 8490 4467 8511 4487
rect 8047 4374 8067 4394
rect 11346 4570 11367 4590
rect 11553 4569 11575 4590
rect 11771 4573 11791 4593
rect 15177 4747 15198 4767
rect 13448 4642 13468 4662
rect 13652 4643 13678 4662
rect 13872 4645 13893 4665
rect 14734 4654 14754 4674
rect 18086 5025 18106 5045
rect 17642 4932 17663 4952
rect 18015 4839 18041 4865
rect 13492 4583 13518 4609
rect 17073 4791 17093 4811
rect 16629 4698 16650 4718
rect 17640 4783 17661 4803
rect 17850 4785 17874 4805
rect 18065 4786 18085 4806
rect 17737 4717 17757 4736
rect 18250 5137 18270 5155
rect 18158 4713 18177 4739
rect 20446 6686 20467 6706
rect 20003 6593 20023 6613
rect 18804 6546 18824 6566
rect 19011 6548 19034 6567
rect 19228 6549 19249 6569
rect 18848 6487 18874 6513
rect 19226 6400 19247 6420
rect 18783 6307 18803 6327
rect 20032 6268 20052 6288
rect 20248 6271 20270 6292
rect 20456 6271 20477 6291
rect 20076 6209 20102 6235
rect 18927 6101 18946 6127
rect 19347 6104 19367 6123
rect 19019 6034 19039 6054
rect 19230 6035 19254 6055
rect 19443 6037 19464 6057
rect 20454 6122 20475 6142
rect 20011 6029 20031 6049
rect 19063 5975 19089 6001
rect 19441 5888 19462 5908
rect 18998 5795 19018 5815
rect 20031 5853 20051 5873
rect 20238 5854 20260 5875
rect 20455 5856 20476 5876
rect 20075 5794 20101 5820
rect 18969 5614 18989 5634
rect 19175 5618 19199 5635
rect 19393 5617 19414 5637
rect 20453 5707 20474 5727
rect 20010 5614 20030 5634
rect 19013 5555 19039 5581
rect 19391 5468 19412 5488
rect 18948 5375 18968 5395
rect 20037 5287 20057 5307
rect 20253 5290 20275 5311
rect 20461 5290 20482 5310
rect 20081 5228 20107 5254
rect 19352 5123 19372 5142
rect 19024 5053 19044 5073
rect 19234 5055 19258 5075
rect 19448 5056 19469 5076
rect 20459 5141 20480 5161
rect 20016 5048 20036 5068
rect 19068 4994 19094 5020
rect 19446 4907 19467 4927
rect 19003 4814 19023 4834
rect 20036 4872 20056 4892
rect 20243 4873 20265 4894
rect 20460 4875 20481 4895
rect 20080 4813 20106 4839
rect 17002 4605 17028 4631
rect 4142 4265 4168 4291
rect 1064 4057 1090 4083
rect 689 4001 710 4021
rect 905 4002 927 4023
rect 1114 4004 1134 4024
rect 2147 4062 2167 4082
rect 1703 3969 1724 3989
rect 2076 3876 2102 3902
rect 1134 3828 1154 3848
rect 690 3735 711 3755
rect 1701 3820 1722 3840
rect 1912 3821 1936 3841
rect 2126 3823 2146 3843
rect 1798 3754 1818 3773
rect 1063 3642 1089 3668
rect 688 3586 709 3606
rect 895 3585 917 3606
rect 1113 3589 1133 3609
rect 2202 3501 2222 3521
rect 1758 3408 1779 3428
rect 2131 3315 2157 3341
rect 1140 3262 1160 3282
rect 696 3169 717 3189
rect 1756 3259 1777 3279
rect 1971 3261 1995 3278
rect 2181 3262 2201 3282
rect 1069 3076 1095 3102
rect 694 3020 715 3040
rect 910 3021 932 3042
rect 1119 3023 1139 3043
rect 2152 3081 2172 3101
rect 1708 2988 1729 3008
rect 2081 2895 2107 2921
rect 1139 2847 1159 2867
rect 695 2754 716 2774
rect 1706 2839 1727 2859
rect 1916 2841 1940 2861
rect 2131 2842 2151 2862
rect 1803 2773 1823 2792
rect 2224 2769 2243 2795
rect 1068 2661 1094 2687
rect 693 2605 714 2625
rect 900 2604 922 2625
rect 1118 2608 1138 2628
rect 2367 2569 2387 2589
rect 1923 2476 1944 2496
rect 2296 2383 2322 2409
rect 1921 2327 1942 2347
rect 2136 2329 2159 2348
rect 2346 2330 2366 2350
rect 1147 2283 1167 2303
rect 703 2190 724 2210
rect 2993 4157 3012 4183
rect 2900 3741 2920 3759
rect 3413 4160 3433 4179
rect 3085 4090 3105 4110
rect 3296 4091 3320 4111
rect 3509 4093 3530 4113
rect 4520 4178 4541 4198
rect 4077 4085 4097 4105
rect 7652 4287 7678 4313
rect 3129 4031 3155 4057
rect 3507 3944 3528 3964
rect 3064 3851 3084 3871
rect 6416 4222 6436 4242
rect 7277 4231 7298 4251
rect 7492 4234 7518 4253
rect 7702 4234 7722 4254
rect 5972 4129 5993 4149
rect 9379 4303 9399 4323
rect 9595 4306 9617 4327
rect 9803 4306 9824 4326
rect 13103 4502 13123 4522
rect 12659 4409 12680 4429
rect 13870 4496 13891 4516
rect 13427 4403 13447 4423
rect 16627 4549 16648 4569
rect 16834 4548 16856 4569
rect 17052 4552 17072 4572
rect 20458 4726 20479 4746
rect 18729 4621 18749 4641
rect 18933 4622 18959 4641
rect 19153 4624 19174 4644
rect 20015 4633 20035 4653
rect 18773 4562 18799 4588
rect 13032 4316 13058 4342
rect 9423 4244 9449 4270
rect 4097 3909 4117 3929
rect 4304 3910 4326 3931
rect 4521 3912 4542 3932
rect 4141 3850 4167 3876
rect 6345 4036 6371 4062
rect 5970 3980 5991 4000
rect 6186 3981 6208 4002
rect 6395 3983 6415 4003
rect 3035 3670 3055 3690
rect 3245 3673 3268 3692
rect 3459 3673 3480 3693
rect 4519 3763 4540 3783
rect 4076 3670 4096 3690
rect 7428 4041 7448 4061
rect 6984 3948 7005 3968
rect 7357 3855 7383 3881
rect 3079 3611 3105 3637
rect 6415 3807 6435 3827
rect 5971 3714 5992 3734
rect 6982 3799 7003 3819
rect 7193 3800 7217 3820
rect 7407 3802 7427 3822
rect 7079 3733 7099 3752
rect 6344 3621 6370 3647
rect 3457 3524 3478 3544
rect 3014 3431 3034 3451
rect 5969 3565 5990 3585
rect 6176 3564 6198 3585
rect 6394 3568 6414 3588
rect 4103 3343 4123 3363
rect 4319 3346 4341 3367
rect 4527 3346 4548 3366
rect 7483 3480 7503 3500
rect 7039 3387 7060 3407
rect 4147 3284 4173 3310
rect 3418 3179 3438 3198
rect 3090 3109 3110 3129
rect 3300 3111 3324 3131
rect 3514 3112 3535 3132
rect 4525 3197 4546 3217
rect 4082 3104 4102 3124
rect 7412 3294 7438 3320
rect 3134 3050 3160 3076
rect 3512 2963 3533 2983
rect 3069 2870 3089 2890
rect 6421 3241 6441 3261
rect 5977 3148 5998 3168
rect 7037 3238 7058 3258
rect 7252 3240 7276 3257
rect 7462 3241 7482 3261
rect 4102 2928 4122 2948
rect 4309 2929 4331 2950
rect 4526 2931 4547 2951
rect 4146 2869 4172 2895
rect 6350 3055 6376 3081
rect 5975 2999 5996 3019
rect 6191 3000 6213 3021
rect 6400 3002 6420 3022
rect 4524 2782 4545 2802
rect 4081 2689 4101 2709
rect 7433 3060 7453 3080
rect 6989 2967 7010 2987
rect 7362 2874 7388 2900
rect 2882 2642 2902 2662
rect 3093 2640 3118 2666
rect 3306 2645 3327 2665
rect 6420 2826 6440 2846
rect 5976 2733 5997 2753
rect 6987 2818 7008 2838
rect 7197 2820 7221 2840
rect 7412 2821 7432 2841
rect 7084 2752 7104 2771
rect 7505 2748 7524 2774
rect 6349 2640 6375 2666
rect 2926 2583 2952 2609
rect 3304 2496 3325 2516
rect 2861 2403 2881 2423
rect 5974 2584 5995 2604
rect 6181 2583 6203 2604
rect 6399 2587 6419 2607
rect 2448 2261 2471 2280
rect 1076 2097 1102 2123
rect 701 2041 722 2061
rect 917 2042 939 2063
rect 1126 2044 1146 2064
rect 2159 2102 2179 2122
rect 1715 2009 1736 2029
rect 2088 1916 2114 1942
rect 1146 1868 1166 1888
rect 702 1775 723 1795
rect 1713 1860 1734 1880
rect 1924 1861 1948 1881
rect 2138 1863 2158 1883
rect 1810 1794 1830 1813
rect 1075 1682 1101 1708
rect 700 1626 721 1646
rect 907 1625 929 1646
rect 1125 1629 1145 1649
rect 2214 1541 2234 1561
rect 1770 1448 1791 1468
rect 2143 1355 2169 1381
rect 1152 1302 1172 1322
rect 708 1209 729 1229
rect 1768 1299 1789 1319
rect 1980 1300 2003 1319
rect 2193 1302 2213 1322
rect 4110 2364 4130 2384
rect 4326 2367 4348 2388
rect 4534 2367 4555 2387
rect 7648 2548 7668 2568
rect 7204 2455 7225 2475
rect 7577 2362 7603 2388
rect 4154 2305 4180 2331
rect 3005 2197 3024 2223
rect 3425 2200 3445 2219
rect 3097 2130 3117 2150
rect 3308 2131 3332 2151
rect 3521 2133 3542 2153
rect 4532 2218 4553 2238
rect 4089 2125 4109 2145
rect 7202 2306 7223 2326
rect 7417 2308 7440 2327
rect 7627 2309 7647 2329
rect 3141 2071 3167 2097
rect 3519 1984 3540 2004
rect 3076 1891 3096 1911
rect 6428 2262 6448 2282
rect 5984 2169 6005 2189
rect 8274 4136 8293 4162
rect 8181 3720 8201 3738
rect 8694 4139 8714 4158
rect 8366 4069 8386 4089
rect 8577 4070 8601 4090
rect 8790 4072 8811 4092
rect 9801 4157 9822 4177
rect 9358 4064 9378 4084
rect 8410 4010 8436 4036
rect 11796 4251 11816 4271
rect 12657 4260 12678 4280
rect 12872 4263 12898 4282
rect 13082 4263 13102 4283
rect 11352 4158 11373 4178
rect 14759 4332 14779 4352
rect 14975 4335 14997 4356
rect 15183 4335 15204 4355
rect 18384 4481 18404 4501
rect 17940 4388 17961 4408
rect 19151 4475 19172 4495
rect 18708 4382 18728 4402
rect 14803 4273 14829 4299
rect 8788 3923 8809 3943
rect 8345 3830 8365 3850
rect 9378 3888 9398 3908
rect 9585 3889 9607 3910
rect 9802 3891 9823 3911
rect 9422 3829 9448 3855
rect 11725 4065 11751 4091
rect 11350 4009 11371 4029
rect 11566 4010 11588 4031
rect 11775 4012 11795 4032
rect 12808 4070 12828 4090
rect 12364 3977 12385 3997
rect 8316 3649 8336 3669
rect 8526 3652 8549 3671
rect 8740 3652 8761 3672
rect 9800 3742 9821 3762
rect 9357 3649 9377 3669
rect 12737 3884 12763 3910
rect 11795 3836 11815 3856
rect 11351 3743 11372 3763
rect 12362 3828 12383 3848
rect 12573 3829 12597 3849
rect 12787 3831 12807 3851
rect 12459 3762 12479 3781
rect 11724 3650 11750 3676
rect 8360 3590 8386 3616
rect 8738 3503 8759 3523
rect 8295 3410 8315 3430
rect 11349 3594 11370 3614
rect 11556 3593 11578 3614
rect 11774 3597 11794 3617
rect 9384 3322 9404 3342
rect 9600 3325 9622 3346
rect 9808 3325 9829 3345
rect 12863 3509 12883 3529
rect 12419 3416 12440 3436
rect 12792 3323 12818 3349
rect 9428 3263 9454 3289
rect 8699 3158 8719 3177
rect 8371 3088 8391 3108
rect 8581 3090 8605 3110
rect 8795 3091 8816 3111
rect 9806 3176 9827 3196
rect 9363 3083 9383 3103
rect 8415 3029 8441 3055
rect 11801 3270 11821 3290
rect 11357 3177 11378 3197
rect 12417 3267 12438 3287
rect 12632 3269 12656 3286
rect 12842 3270 12862 3290
rect 8793 2942 8814 2962
rect 8350 2849 8370 2869
rect 9383 2907 9403 2927
rect 9590 2908 9612 2929
rect 9807 2910 9828 2930
rect 9427 2848 9453 2874
rect 11730 3084 11756 3110
rect 11355 3028 11376 3048
rect 11571 3029 11593 3050
rect 11780 3031 11800 3051
rect 12813 3089 12833 3109
rect 12369 2996 12390 3016
rect 9805 2761 9826 2781
rect 9362 2668 9382 2688
rect 12742 2903 12768 2929
rect 8163 2621 8183 2641
rect 8374 2619 8399 2645
rect 8587 2624 8608 2644
rect 11800 2855 11820 2875
rect 11356 2762 11377 2782
rect 12367 2847 12388 2867
rect 12577 2849 12601 2869
rect 12792 2850 12812 2870
rect 12464 2781 12484 2800
rect 12885 2777 12904 2803
rect 11729 2669 11755 2695
rect 8207 2562 8233 2588
rect 11354 2613 11375 2633
rect 11561 2612 11583 2633
rect 11779 2616 11799 2636
rect 8585 2475 8606 2495
rect 8142 2382 8162 2402
rect 7729 2240 7752 2259
rect 4109 1949 4129 1969
rect 4316 1950 4338 1971
rect 4533 1952 4554 1972
rect 4153 1890 4179 1916
rect 6357 2076 6383 2102
rect 5982 2020 6003 2040
rect 6198 2021 6220 2042
rect 6407 2023 6427 2043
rect 3047 1710 3067 1730
rect 3253 1714 3277 1731
rect 3471 1713 3492 1733
rect 4531 1803 4552 1823
rect 4088 1710 4108 1730
rect 7440 2081 7460 2101
rect 6996 1988 7017 2008
rect 7369 1895 7395 1921
rect 3091 1651 3117 1677
rect 6427 1847 6447 1867
rect 5983 1754 6004 1774
rect 6994 1839 7015 1859
rect 7205 1840 7229 1860
rect 7419 1842 7439 1862
rect 7091 1773 7111 1792
rect 6356 1661 6382 1687
rect 3469 1564 3490 1584
rect 3026 1471 3046 1491
rect 5981 1605 6002 1625
rect 6188 1604 6210 1625
rect 6406 1608 6426 1628
rect 4115 1383 4135 1403
rect 4331 1386 4353 1407
rect 4539 1386 4560 1406
rect 7495 1520 7515 1540
rect 7051 1427 7072 1447
rect 4159 1324 4185 1350
rect 1081 1116 1107 1142
rect 706 1060 727 1080
rect 922 1061 944 1082
rect 1131 1063 1151 1083
rect 2164 1121 2184 1141
rect 1720 1028 1741 1048
rect 2093 935 2119 961
rect 1151 887 1171 907
rect 707 794 728 814
rect 1718 879 1739 899
rect 1928 881 1952 901
rect 2143 882 2163 902
rect 1815 813 1835 832
rect 2328 1233 2348 1251
rect 3430 1219 3450 1238
rect 3102 1149 3122 1169
rect 3312 1151 3336 1171
rect 3526 1152 3547 1172
rect 4537 1237 4558 1257
rect 4094 1144 4114 1164
rect 7424 1334 7450 1360
rect 3146 1090 3172 1116
rect 3524 1003 3545 1023
rect 3081 910 3101 930
rect 6433 1281 6453 1301
rect 5989 1188 6010 1208
rect 7049 1278 7070 1298
rect 7261 1279 7284 1298
rect 7474 1281 7494 1301
rect 13028 2577 13048 2597
rect 12584 2484 12605 2504
rect 9391 2343 9411 2363
rect 9607 2346 9629 2367
rect 9815 2346 9836 2366
rect 12957 2391 12983 2417
rect 9435 2284 9461 2310
rect 8286 2176 8305 2202
rect 8706 2179 8726 2198
rect 8378 2109 8398 2129
rect 8589 2110 8613 2130
rect 8802 2112 8823 2132
rect 9813 2197 9834 2217
rect 9370 2104 9390 2124
rect 12582 2335 12603 2355
rect 12797 2337 12820 2356
rect 13007 2338 13027 2358
rect 8422 2050 8448 2076
rect 11808 2291 11828 2311
rect 11364 2198 11385 2218
rect 13654 4165 13673 4191
rect 13561 3749 13581 3767
rect 14074 4168 14094 4187
rect 13746 4098 13766 4118
rect 13957 4099 13981 4119
rect 14170 4101 14191 4121
rect 15181 4186 15202 4206
rect 14738 4093 14758 4113
rect 18313 4295 18339 4321
rect 13790 4039 13816 4065
rect 14168 3952 14189 3972
rect 13725 3859 13745 3879
rect 17077 4230 17097 4250
rect 17938 4239 17959 4259
rect 18153 4242 18179 4261
rect 18363 4242 18383 4262
rect 16633 4137 16654 4157
rect 20040 4311 20060 4331
rect 20256 4314 20278 4335
rect 20464 4314 20485 4334
rect 20084 4252 20110 4278
rect 14758 3917 14778 3937
rect 14965 3918 14987 3939
rect 15182 3920 15203 3940
rect 14802 3858 14828 3884
rect 17006 4044 17032 4070
rect 16631 3988 16652 4008
rect 16847 3989 16869 4010
rect 17056 3991 17076 4011
rect 13696 3678 13716 3698
rect 13906 3681 13929 3700
rect 14120 3681 14141 3701
rect 15180 3771 15201 3791
rect 14737 3678 14757 3698
rect 18089 4049 18109 4069
rect 17645 3956 17666 3976
rect 18018 3863 18044 3889
rect 13740 3619 13766 3645
rect 17076 3815 17096 3835
rect 16632 3722 16653 3742
rect 17643 3807 17664 3827
rect 17854 3808 17878 3828
rect 18068 3810 18088 3830
rect 17740 3741 17760 3760
rect 17005 3629 17031 3655
rect 14118 3532 14139 3552
rect 13675 3439 13695 3459
rect 16630 3573 16651 3593
rect 16837 3572 16859 3593
rect 17055 3576 17075 3596
rect 14764 3351 14784 3371
rect 14980 3354 15002 3375
rect 15188 3354 15209 3374
rect 18144 3488 18164 3508
rect 17700 3395 17721 3415
rect 14808 3292 14834 3318
rect 14079 3187 14099 3206
rect 13751 3117 13771 3137
rect 13961 3119 13985 3139
rect 14175 3120 14196 3140
rect 15186 3205 15207 3225
rect 14743 3112 14763 3132
rect 18073 3302 18099 3328
rect 13795 3058 13821 3084
rect 14173 2971 14194 2991
rect 13730 2878 13750 2898
rect 17082 3249 17102 3269
rect 16638 3156 16659 3176
rect 17698 3246 17719 3266
rect 17913 3248 17937 3265
rect 18123 3249 18143 3269
rect 14763 2936 14783 2956
rect 14970 2937 14992 2958
rect 15187 2939 15208 2959
rect 14807 2877 14833 2903
rect 17011 3063 17037 3089
rect 16636 3007 16657 3027
rect 16852 3008 16874 3029
rect 17061 3010 17081 3030
rect 15185 2790 15206 2810
rect 14742 2697 14762 2717
rect 18094 3068 18114 3088
rect 17650 2975 17671 2995
rect 18023 2882 18049 2908
rect 13543 2650 13563 2670
rect 13754 2648 13779 2674
rect 13967 2653 13988 2673
rect 17081 2834 17101 2854
rect 16637 2741 16658 2761
rect 17648 2826 17669 2846
rect 17858 2828 17882 2848
rect 18073 2829 18093 2849
rect 17745 2760 17765 2779
rect 18166 2756 18185 2782
rect 17010 2648 17036 2674
rect 13587 2591 13613 2617
rect 13965 2504 13986 2524
rect 13522 2411 13542 2431
rect 16635 2592 16656 2612
rect 16842 2591 16864 2612
rect 17060 2595 17080 2615
rect 13109 2269 13132 2288
rect 8800 1963 8821 1983
rect 8357 1870 8377 1890
rect 9390 1928 9410 1948
rect 9597 1929 9619 1950
rect 9814 1931 9835 1951
rect 9434 1869 9460 1895
rect 11737 2105 11763 2131
rect 11362 2049 11383 2069
rect 11578 2050 11600 2071
rect 11787 2052 11807 2072
rect 12820 2110 12840 2130
rect 12376 2017 12397 2037
rect 8328 1689 8348 1709
rect 8534 1693 8558 1710
rect 8752 1692 8773 1712
rect 9812 1782 9833 1802
rect 9369 1689 9389 1709
rect 12749 1924 12775 1950
rect 11807 1876 11827 1896
rect 11363 1783 11384 1803
rect 12374 1868 12395 1888
rect 12585 1869 12609 1889
rect 12799 1871 12819 1891
rect 12471 1802 12491 1821
rect 11736 1690 11762 1716
rect 8372 1630 8398 1656
rect 8750 1543 8771 1563
rect 8307 1450 8327 1470
rect 11361 1634 11382 1654
rect 11568 1633 11590 1654
rect 11786 1637 11806 1657
rect 9396 1362 9416 1382
rect 9612 1365 9634 1386
rect 9820 1365 9841 1385
rect 12875 1549 12895 1569
rect 12431 1456 12452 1476
rect 12804 1363 12830 1389
rect 9440 1303 9466 1329
rect 4114 968 4134 988
rect 4321 969 4343 990
rect 4538 971 4559 991
rect 4158 909 4184 935
rect 6362 1095 6388 1121
rect 5987 1039 6008 1059
rect 6203 1040 6225 1061
rect 6412 1042 6432 1062
rect 2236 809 2255 835
rect 1080 701 1106 727
rect 705 645 726 665
rect 912 644 934 665
rect 1130 648 1150 668
rect 4536 822 4557 842
rect 4093 729 4113 749
rect 7445 1100 7465 1120
rect 7001 1007 7022 1027
rect 7374 914 7400 940
rect 6432 866 6452 886
rect 5988 773 6009 793
rect 6999 858 7020 878
rect 7209 860 7233 880
rect 7424 861 7444 881
rect 7096 792 7116 811
rect 7609 1212 7629 1230
rect 8711 1198 8731 1217
rect 8383 1128 8403 1148
rect 8593 1130 8617 1150
rect 8807 1131 8828 1151
rect 9818 1216 9839 1236
rect 9375 1123 9395 1143
rect 8427 1069 8453 1095
rect 11813 1310 11833 1330
rect 11369 1217 11390 1237
rect 12429 1307 12450 1327
rect 12641 1308 12664 1327
rect 12854 1310 12874 1330
rect 14771 2372 14791 2392
rect 14987 2375 15009 2396
rect 15195 2375 15216 2395
rect 18309 2556 18329 2576
rect 17865 2463 17886 2483
rect 18238 2370 18264 2396
rect 14815 2313 14841 2339
rect 13666 2205 13685 2231
rect 14086 2208 14106 2227
rect 13758 2138 13778 2158
rect 13969 2139 13993 2159
rect 14182 2141 14203 2161
rect 15193 2226 15214 2246
rect 14750 2133 14770 2153
rect 17863 2314 17884 2334
rect 18078 2316 18101 2335
rect 18288 2317 18308 2337
rect 13802 2079 13828 2105
rect 14180 1992 14201 2012
rect 13737 1899 13757 1919
rect 17089 2270 17109 2290
rect 16645 2177 16666 2197
rect 18935 4144 18954 4170
rect 18842 3728 18862 3746
rect 19355 4147 19375 4166
rect 19027 4077 19047 4097
rect 19238 4078 19262 4098
rect 19451 4080 19472 4100
rect 20462 4165 20483 4185
rect 20019 4072 20039 4092
rect 19071 4018 19097 4044
rect 19449 3931 19470 3951
rect 19006 3838 19026 3858
rect 20039 3896 20059 3916
rect 20246 3897 20268 3918
rect 20463 3899 20484 3919
rect 20083 3837 20109 3863
rect 18977 3657 18997 3677
rect 19187 3660 19210 3679
rect 19401 3660 19422 3680
rect 20461 3750 20482 3770
rect 20018 3657 20038 3677
rect 19021 3598 19047 3624
rect 19399 3511 19420 3531
rect 18956 3418 18976 3438
rect 20045 3330 20065 3350
rect 20261 3333 20283 3354
rect 20469 3333 20490 3353
rect 20089 3271 20115 3297
rect 19360 3166 19380 3185
rect 19032 3096 19052 3116
rect 19242 3098 19266 3118
rect 19456 3099 19477 3119
rect 20467 3184 20488 3204
rect 20024 3091 20044 3111
rect 19076 3037 19102 3063
rect 19454 2950 19475 2970
rect 19011 2857 19031 2877
rect 20044 2915 20064 2935
rect 20251 2916 20273 2937
rect 20468 2918 20489 2938
rect 20088 2856 20114 2882
rect 20466 2769 20487 2789
rect 20023 2676 20043 2696
rect 18824 2629 18844 2649
rect 19035 2627 19060 2653
rect 19248 2632 19269 2652
rect 18868 2570 18894 2596
rect 19246 2483 19267 2503
rect 18803 2390 18823 2410
rect 18390 2248 18413 2267
rect 14770 1957 14790 1977
rect 14977 1958 14999 1979
rect 15194 1960 15215 1980
rect 14814 1898 14840 1924
rect 17018 2084 17044 2110
rect 16643 2028 16664 2048
rect 16859 2029 16881 2050
rect 17068 2031 17088 2051
rect 13708 1718 13728 1738
rect 13914 1722 13938 1739
rect 14132 1721 14153 1741
rect 15192 1811 15213 1831
rect 14749 1718 14769 1738
rect 18101 2089 18121 2109
rect 17657 1996 17678 2016
rect 18030 1903 18056 1929
rect 13752 1659 13778 1685
rect 17088 1855 17108 1875
rect 16644 1762 16665 1782
rect 17655 1847 17676 1867
rect 17866 1848 17890 1868
rect 18080 1850 18100 1870
rect 17752 1781 17772 1800
rect 17017 1669 17043 1695
rect 14130 1572 14151 1592
rect 13687 1479 13707 1499
rect 16642 1613 16663 1633
rect 16849 1612 16871 1633
rect 17067 1616 17087 1636
rect 14776 1391 14796 1411
rect 14992 1394 15014 1415
rect 15200 1394 15221 1414
rect 18156 1528 18176 1548
rect 17712 1435 17733 1455
rect 14820 1332 14846 1358
rect 8805 982 8826 1002
rect 8362 889 8382 909
rect 9395 947 9415 967
rect 9602 948 9624 969
rect 9819 950 9840 970
rect 9439 888 9465 914
rect 11742 1124 11768 1150
rect 11367 1068 11388 1088
rect 11583 1069 11605 1090
rect 11792 1071 11812 1091
rect 12825 1129 12845 1149
rect 12381 1036 12402 1056
rect 7517 788 7536 814
rect 6361 680 6387 706
rect 756 520 779 542
rect 5986 624 6007 644
rect 6193 623 6215 644
rect 6411 627 6431 647
rect 5089 520 5112 542
rect 9817 801 9838 821
rect 9374 708 9394 728
rect 12754 943 12780 969
rect 11812 895 11832 915
rect 11368 802 11389 822
rect 12379 887 12400 907
rect 12589 889 12613 909
rect 12804 890 12824 910
rect 12476 821 12496 840
rect 12989 1241 13009 1259
rect 14091 1227 14111 1246
rect 13763 1157 13783 1177
rect 13973 1159 13997 1179
rect 14187 1160 14208 1180
rect 15198 1245 15219 1265
rect 14755 1152 14775 1172
rect 18085 1342 18111 1368
rect 13807 1098 13833 1124
rect 14185 1011 14206 1031
rect 13742 918 13762 938
rect 17094 1289 17114 1309
rect 16650 1196 16671 1216
rect 17710 1286 17731 1306
rect 17922 1287 17945 1306
rect 18135 1289 18155 1309
rect 20052 2351 20072 2371
rect 20268 2354 20290 2375
rect 20476 2354 20497 2374
rect 20096 2292 20122 2318
rect 18947 2184 18966 2210
rect 19367 2187 19387 2206
rect 19039 2117 19059 2137
rect 19250 2118 19274 2138
rect 19463 2120 19484 2140
rect 20474 2205 20495 2225
rect 20031 2112 20051 2132
rect 19083 2058 19109 2084
rect 19461 1971 19482 1991
rect 19018 1878 19038 1898
rect 20051 1936 20071 1956
rect 20258 1937 20280 1958
rect 20475 1939 20496 1959
rect 20095 1877 20121 1903
rect 18989 1697 19009 1717
rect 19195 1701 19219 1718
rect 19413 1700 19434 1720
rect 20473 1790 20494 1810
rect 20030 1697 20050 1717
rect 19033 1638 19059 1664
rect 19411 1551 19432 1571
rect 18968 1458 18988 1478
rect 20057 1370 20077 1390
rect 20273 1373 20295 1394
rect 20481 1373 20502 1393
rect 20101 1311 20127 1337
rect 14775 976 14795 996
rect 14982 977 15004 998
rect 15199 979 15220 999
rect 14819 917 14845 943
rect 17023 1103 17049 1129
rect 16648 1047 16669 1067
rect 16864 1048 16886 1069
rect 17073 1050 17093 1070
rect 12897 817 12916 843
rect 11741 709 11767 735
rect 11366 653 11387 673
rect 11573 652 11595 673
rect 11791 656 11811 676
rect 6037 499 6060 521
rect 10370 499 10393 521
rect 15197 830 15218 850
rect 14754 737 14774 757
rect 18106 1108 18126 1128
rect 17662 1015 17683 1035
rect 18035 922 18061 948
rect 17093 874 17113 894
rect 16649 781 16670 801
rect 17660 866 17681 886
rect 17870 868 17894 888
rect 18085 869 18105 889
rect 17757 800 17777 819
rect 18270 1220 18290 1238
rect 19372 1206 19392 1225
rect 19044 1136 19064 1156
rect 19254 1138 19278 1158
rect 19468 1139 19489 1159
rect 20479 1224 20500 1244
rect 20036 1131 20056 1151
rect 19088 1077 19114 1103
rect 19466 990 19487 1010
rect 19023 897 19043 917
rect 20056 955 20076 975
rect 20263 956 20285 977
rect 20480 958 20501 978
rect 20100 896 20126 922
rect 18178 796 18197 822
rect 17022 688 17048 714
rect 11417 528 11440 550
rect 16647 632 16668 652
rect 16854 631 16876 652
rect 17072 635 17092 655
rect 15750 528 15773 550
rect 20478 809 20499 829
rect 20035 716 20055 736
rect 16698 507 16721 529
rect 21031 507 21054 529
rect 2554 406 2574 426
rect 2110 313 2131 333
rect 2651 311 2679 331
rect 2483 220 2509 246
rect 2108 164 2129 184
rect 2322 162 2347 184
rect 2533 167 2553 187
rect 5644 318 5664 338
rect 5200 225 5221 245
rect 7835 385 7855 405
rect 7391 292 7412 312
rect 7932 290 7960 310
rect 5573 132 5599 158
rect 5198 76 5219 96
rect 5409 76 5430 93
rect 5623 79 5643 99
rect 7764 199 7790 225
rect 7389 143 7410 163
rect 7603 141 7628 163
rect 7814 146 7834 166
rect 10905 311 10925 331
rect 10461 218 10482 238
rect 13215 414 13235 434
rect 12771 321 12792 341
rect 13312 319 13340 339
rect 13144 228 13170 254
rect 10834 125 10860 151
rect 10459 69 10480 89
rect 10668 68 10696 91
rect 10884 72 10904 92
rect 5659 9 5683 26
rect 12769 172 12790 192
rect 12983 170 13008 192
rect 13194 175 13214 195
rect 16305 326 16325 346
rect 15861 233 15882 253
rect 18496 393 18516 413
rect 18052 300 18073 320
rect 18593 298 18621 318
rect 16234 140 16260 166
rect 15859 84 15880 104
rect 16070 84 16091 101
rect 16284 87 16304 107
rect 18425 207 18451 233
rect 18050 151 18071 171
rect 18264 149 18289 171
rect 18475 154 18495 174
rect 16320 17 16344 34
rect 10925 -45 10945 -24
<< metal1 >>
rect 14575 8343 14984 8344
rect 3914 8335 4323 8336
rect 3908 8306 4323 8335
rect 9195 8314 9604 8315
rect 1111 8185 1143 8186
rect 1108 8180 1143 8185
rect 1108 8160 1115 8180
rect 1135 8160 1143 8180
rect 1108 8152 1143 8160
rect 3908 8155 3948 8306
rect 4282 8273 4323 8306
rect 9189 8285 9604 8314
rect 4070 8268 4105 8269
rect 664 8087 696 8094
rect 664 8067 671 8087
rect 692 8067 696 8087
rect 664 8002 696 8067
rect 1034 8002 1074 8003
rect 664 8000 1076 8002
rect 664 7974 1044 8000
rect 1070 7974 1076 8000
rect 664 7966 1076 7974
rect 664 7938 696 7966
rect 1109 7946 1143 8152
rect 3385 8127 3948 8155
rect 4049 8261 4105 8268
rect 4049 8241 4078 8261
rect 4098 8241 4105 8261
rect 4049 8236 4105 8241
rect 4278 8265 4328 8273
rect 4278 8244 4294 8265
rect 4316 8244 4328 8265
rect 2964 8100 3311 8104
rect 2964 8074 2973 8100
rect 2992 8074 3311 8100
rect 3386 8099 3420 8127
rect 2964 8069 3311 8074
rect 3385 8096 3421 8099
rect 3385 8077 3393 8096
rect 3413 8077 3421 8096
rect 3385 8073 3421 8077
rect 3271 8039 3311 8069
rect 3057 8034 3092 8035
rect 664 7918 669 7938
rect 690 7918 696 7938
rect 664 7911 696 7918
rect 873 7940 913 7945
rect 873 7919 885 7940
rect 907 7919 913 7940
rect 873 7907 913 7919
rect 1087 7941 1143 7946
rect 1087 7921 1094 7941
rect 1114 7921 1143 7941
rect 1087 7914 1143 7921
rect 1200 8015 2157 8034
rect 3036 8027 3092 8034
rect 1087 7913 1122 7914
rect 879 7875 907 7907
rect 1200 7875 1231 8015
rect 2120 7999 2155 8015
rect 2120 7979 2127 7999
rect 2147 7979 2155 7999
rect 2120 7971 2155 7979
rect 879 7844 1231 7875
rect 1676 7906 1708 7913
rect 1676 7886 1683 7906
rect 1704 7886 1708 7906
rect 1676 7821 1708 7886
rect 2046 7821 2086 7822
rect 1676 7819 2088 7821
rect 1676 7793 2056 7819
rect 2082 7793 2088 7819
rect 1676 7785 2088 7793
rect 1110 7770 1142 7771
rect 1107 7765 1142 7770
rect 1107 7745 1114 7765
rect 1134 7745 1142 7765
rect 1107 7737 1142 7745
rect 663 7672 695 7679
rect 663 7652 670 7672
rect 691 7652 695 7672
rect 663 7587 695 7652
rect 1033 7587 1073 7588
rect 663 7585 1075 7587
rect 663 7559 1043 7585
rect 1069 7559 1075 7585
rect 663 7551 1075 7559
rect 663 7523 695 7551
rect 663 7503 668 7523
rect 689 7503 695 7523
rect 663 7496 695 7503
rect 863 7523 913 7532
rect 1108 7531 1142 7737
rect 1676 7757 1708 7785
rect 1676 7737 1681 7757
rect 1702 7737 1708 7757
rect 1676 7730 1708 7737
rect 1883 7758 1925 7766
rect 2121 7765 2155 7971
rect 1883 7738 1892 7758
rect 1916 7738 1925 7758
rect 1883 7726 1925 7738
rect 2099 7760 2155 7765
rect 2099 7740 2106 7760
rect 2126 7740 2155 7760
rect 3036 8007 3065 8027
rect 3085 8007 3092 8027
rect 3036 8002 3092 8007
rect 3268 8028 3311 8039
rect 3268 8008 3276 8028
rect 3300 8022 3311 8028
rect 3483 8030 3515 8037
rect 3300 8008 3310 8022
rect 3036 7796 3070 8002
rect 3268 7999 3310 8008
rect 3483 8010 3489 8030
rect 3510 8010 3515 8030
rect 3483 7982 3515 8010
rect 4049 8030 4083 8236
rect 4278 8235 4328 8244
rect 4496 8264 4528 8271
rect 4496 8244 4502 8264
rect 4523 8244 4528 8264
rect 4496 8216 4528 8244
rect 4116 8208 4528 8216
rect 4116 8182 4122 8208
rect 4148 8182 4528 8208
rect 4116 8180 4528 8182
rect 4118 8179 4158 8180
rect 4496 8115 4528 8180
rect 6392 8164 6424 8165
rect 6389 8159 6424 8164
rect 6389 8139 6396 8159
rect 6416 8139 6424 8159
rect 6389 8131 6424 8139
rect 9189 8134 9229 8285
rect 9563 8252 9604 8285
rect 14569 8314 14984 8343
rect 19856 8322 20265 8323
rect 9351 8247 9386 8248
rect 4496 8095 4500 8115
rect 4521 8095 4528 8115
rect 4496 8088 4528 8095
rect 5945 8066 5977 8073
rect 5945 8046 5952 8066
rect 5973 8046 5977 8066
rect 4049 8022 4084 8030
rect 4049 8002 4057 8022
rect 4077 8002 4084 8022
rect 4049 7997 4084 8002
rect 4049 7996 4081 7997
rect 3103 7974 3515 7982
rect 3103 7948 3109 7974
rect 3135 7948 3515 7974
rect 3103 7946 3515 7948
rect 3105 7945 3145 7946
rect 3483 7881 3515 7946
rect 5945 7981 5977 8046
rect 6315 7981 6355 7982
rect 5945 7979 6357 7981
rect 5945 7953 6325 7979
rect 6351 7953 6357 7979
rect 5945 7945 6357 7953
rect 3483 7861 3487 7881
rect 3508 7861 3515 7881
rect 3483 7854 3515 7861
rect 3960 7892 4312 7923
rect 3036 7788 3071 7796
rect 3036 7768 3044 7788
rect 3064 7768 3071 7788
rect 3036 7752 3071 7768
rect 3960 7752 3991 7892
rect 4284 7860 4312 7892
rect 5945 7917 5977 7945
rect 6390 7925 6424 8131
rect 8666 8106 9229 8134
rect 9330 8240 9386 8247
rect 9330 8220 9359 8240
rect 9379 8220 9386 8240
rect 9330 8215 9386 8220
rect 9559 8244 9609 8252
rect 9559 8223 9575 8244
rect 9597 8223 9609 8244
rect 8245 8079 8592 8083
rect 8245 8053 8254 8079
rect 8273 8053 8592 8079
rect 8667 8078 8701 8106
rect 8245 8048 8592 8053
rect 8666 8075 8702 8078
rect 8666 8056 8674 8075
rect 8694 8056 8702 8075
rect 8666 8052 8702 8056
rect 8552 8018 8592 8048
rect 8338 8013 8373 8014
rect 5945 7897 5950 7917
rect 5971 7897 5977 7917
rect 5945 7890 5977 7897
rect 6154 7919 6194 7924
rect 6154 7898 6166 7919
rect 6188 7898 6194 7919
rect 6154 7886 6194 7898
rect 6368 7920 6424 7925
rect 6368 7900 6375 7920
rect 6395 7900 6424 7920
rect 6368 7893 6424 7900
rect 6481 7994 7438 8013
rect 8317 8006 8373 8013
rect 6368 7892 6403 7893
rect 4069 7853 4104 7854
rect 2099 7733 2155 7740
rect 3034 7733 3991 7752
rect 4048 7846 4104 7853
rect 4048 7826 4077 7846
rect 4097 7826 4104 7846
rect 4048 7821 4104 7826
rect 4278 7848 4318 7860
rect 4278 7827 4284 7848
rect 4306 7827 4318 7848
rect 4278 7822 4318 7827
rect 4495 7849 4527 7856
rect 4495 7829 4501 7849
rect 4522 7829 4527 7849
rect 2099 7732 2134 7733
rect 1885 7697 1920 7726
rect 1885 7696 2195 7697
rect 1770 7690 1806 7694
rect 1770 7671 1778 7690
rect 1798 7671 1806 7690
rect 1770 7668 1806 7671
rect 1771 7640 1805 7668
rect 1885 7662 2212 7696
rect 863 7502 875 7523
rect 897 7502 913 7523
rect 863 7494 913 7502
rect 1086 7526 1142 7531
rect 1086 7506 1093 7526
rect 1113 7506 1142 7526
rect 1086 7499 1142 7506
rect 1243 7612 1806 7640
rect 1086 7498 1121 7499
rect 868 7461 909 7494
rect 1243 7461 1283 7612
rect 868 7432 1283 7461
rect 2172 7438 2212 7662
rect 2873 7681 2902 7683
rect 2873 7676 3246 7681
rect 2873 7658 2880 7676
rect 2900 7658 3246 7676
rect 2873 7653 3246 7658
rect 2878 7651 3246 7653
rect 3007 7614 3042 7615
rect 3222 7614 3246 7651
rect 868 7431 1277 7432
rect 2172 7418 2182 7438
rect 2202 7418 2212 7438
rect 2172 7408 2212 7418
rect 2986 7607 3042 7614
rect 2986 7587 3015 7607
rect 3035 7587 3042 7607
rect 2986 7582 3042 7587
rect 3217 7609 3254 7614
rect 3217 7590 3225 7609
rect 3248 7590 3254 7609
rect 3217 7584 3254 7590
rect 3433 7610 3465 7617
rect 3433 7590 3439 7610
rect 3460 7590 3465 7610
rect 1731 7345 1763 7352
rect 1731 7325 1738 7345
rect 1759 7325 1763 7345
rect 1731 7260 1763 7325
rect 2101 7260 2141 7261
rect 1731 7258 2143 7260
rect 1731 7232 2111 7258
rect 2137 7232 2143 7258
rect 1731 7224 2143 7232
rect 1116 7204 1148 7205
rect 1113 7199 1148 7204
rect 1113 7179 1120 7199
rect 1140 7179 1148 7199
rect 1113 7171 1148 7179
rect 669 7106 701 7113
rect 669 7086 676 7106
rect 697 7086 701 7106
rect 669 7021 701 7086
rect 1039 7021 1079 7022
rect 669 7019 1081 7021
rect 669 6993 1049 7019
rect 1075 6993 1081 7019
rect 669 6985 1081 6993
rect 669 6957 701 6985
rect 1114 6965 1148 7171
rect 1731 7196 1763 7224
rect 1731 7176 1736 7196
rect 1757 7176 1763 7196
rect 1731 7169 1763 7176
rect 1942 7195 1980 7207
rect 2176 7204 2210 7408
rect 2986 7378 3020 7582
rect 3433 7562 3465 7590
rect 4048 7615 4082 7821
rect 4495 7801 4527 7829
rect 6160 7854 6188 7886
rect 6481 7854 6512 7994
rect 7401 7978 7436 7994
rect 7401 7958 7408 7978
rect 7428 7958 7436 7978
rect 7401 7950 7436 7958
rect 6160 7823 6512 7854
rect 6957 7885 6989 7892
rect 6957 7865 6964 7885
rect 6985 7865 6989 7885
rect 4115 7793 4527 7801
rect 4115 7767 4121 7793
rect 4147 7767 4527 7793
rect 4115 7765 4527 7767
rect 4117 7764 4157 7765
rect 4495 7700 4527 7765
rect 6957 7800 6989 7865
rect 7327 7800 7367 7801
rect 6957 7798 7369 7800
rect 6957 7772 7337 7798
rect 7363 7772 7369 7798
rect 6957 7764 7369 7772
rect 6391 7749 6423 7750
rect 6388 7744 6423 7749
rect 6388 7724 6395 7744
rect 6415 7724 6423 7744
rect 6388 7716 6423 7724
rect 4495 7680 4499 7700
rect 4520 7680 4527 7700
rect 4495 7673 4527 7680
rect 5944 7651 5976 7658
rect 5944 7631 5951 7651
rect 5972 7631 5976 7651
rect 4048 7607 4083 7615
rect 4048 7587 4056 7607
rect 4076 7587 4083 7607
rect 4048 7582 4083 7587
rect 4048 7581 4080 7582
rect 3053 7554 3465 7562
rect 3053 7528 3059 7554
rect 3085 7528 3465 7554
rect 3053 7526 3465 7528
rect 3055 7525 3095 7526
rect 3433 7461 3465 7526
rect 5944 7566 5976 7631
rect 6314 7566 6354 7567
rect 5944 7564 6356 7566
rect 5944 7538 6324 7564
rect 6350 7538 6356 7564
rect 5944 7530 6356 7538
rect 5944 7502 5976 7530
rect 5944 7482 5949 7502
rect 5970 7482 5976 7502
rect 5944 7475 5976 7482
rect 6144 7502 6194 7511
rect 6389 7510 6423 7716
rect 6957 7736 6989 7764
rect 6957 7716 6962 7736
rect 6983 7716 6989 7736
rect 6957 7709 6989 7716
rect 7164 7737 7206 7745
rect 7402 7744 7436 7950
rect 7164 7717 7173 7737
rect 7197 7717 7206 7737
rect 7164 7705 7206 7717
rect 7380 7739 7436 7744
rect 7380 7719 7387 7739
rect 7407 7719 7436 7739
rect 8317 7986 8346 8006
rect 8366 7986 8373 8006
rect 8317 7981 8373 7986
rect 8549 8007 8592 8018
rect 8549 7987 8557 8007
rect 8581 8001 8592 8007
rect 8764 8009 8796 8016
rect 8581 7987 8591 8001
rect 8317 7775 8351 7981
rect 8549 7978 8591 7987
rect 8764 7989 8770 8009
rect 8791 7989 8796 8009
rect 8764 7961 8796 7989
rect 9330 8009 9364 8215
rect 9559 8214 9609 8223
rect 9777 8243 9809 8250
rect 9777 8223 9783 8243
rect 9804 8223 9809 8243
rect 9777 8195 9809 8223
rect 9397 8187 9809 8195
rect 11772 8193 11804 8194
rect 9397 8161 9403 8187
rect 9429 8161 9809 8187
rect 9397 8159 9809 8161
rect 11769 8188 11804 8193
rect 11769 8168 11776 8188
rect 11796 8168 11804 8188
rect 11769 8160 11804 8168
rect 14569 8163 14609 8314
rect 14943 8281 14984 8314
rect 19850 8293 20265 8322
rect 14731 8276 14766 8277
rect 9399 8158 9439 8159
rect 9777 8094 9809 8159
rect 9777 8074 9781 8094
rect 9802 8074 9809 8094
rect 9777 8067 9809 8074
rect 11325 8095 11357 8102
rect 11325 8075 11332 8095
rect 11353 8075 11357 8095
rect 11325 8010 11357 8075
rect 11695 8010 11735 8011
rect 9330 8001 9365 8009
rect 9330 7981 9338 8001
rect 9358 7981 9365 8001
rect 9330 7976 9365 7981
rect 11325 8008 11737 8010
rect 11325 7982 11705 8008
rect 11731 7982 11737 8008
rect 9330 7975 9362 7976
rect 8384 7953 8796 7961
rect 8384 7927 8390 7953
rect 8416 7927 8796 7953
rect 8384 7925 8796 7927
rect 8386 7924 8426 7925
rect 8764 7860 8796 7925
rect 11325 7974 11737 7982
rect 11325 7946 11357 7974
rect 11770 7954 11804 8160
rect 14046 8135 14609 8163
rect 14710 8269 14766 8276
rect 14710 8249 14739 8269
rect 14759 8249 14766 8269
rect 14710 8244 14766 8249
rect 14939 8273 14989 8281
rect 14939 8252 14955 8273
rect 14977 8252 14989 8273
rect 13625 8108 13972 8112
rect 13625 8082 13634 8108
rect 13653 8082 13972 8108
rect 14047 8107 14081 8135
rect 13625 8077 13972 8082
rect 14046 8104 14082 8107
rect 14046 8085 14054 8104
rect 14074 8085 14082 8104
rect 14046 8081 14082 8085
rect 13932 8047 13972 8077
rect 13718 8042 13753 8043
rect 11325 7926 11330 7946
rect 11351 7926 11357 7946
rect 11325 7919 11357 7926
rect 11534 7948 11574 7953
rect 11534 7927 11546 7948
rect 11568 7927 11574 7948
rect 11534 7915 11574 7927
rect 11748 7949 11804 7954
rect 11748 7929 11755 7949
rect 11775 7929 11804 7949
rect 11748 7922 11804 7929
rect 11861 8023 12818 8042
rect 13697 8035 13753 8042
rect 11748 7921 11783 7922
rect 8764 7840 8768 7860
rect 8789 7840 8796 7860
rect 8764 7833 8796 7840
rect 9241 7871 9593 7902
rect 8317 7767 8352 7775
rect 8317 7747 8325 7767
rect 8345 7747 8352 7767
rect 8317 7731 8352 7747
rect 9241 7731 9272 7871
rect 9565 7839 9593 7871
rect 11540 7883 11568 7915
rect 11861 7883 11892 8023
rect 12781 8007 12816 8023
rect 12781 7987 12788 8007
rect 12808 7987 12816 8007
rect 12781 7979 12816 7987
rect 11540 7852 11892 7883
rect 12337 7914 12369 7921
rect 12337 7894 12344 7914
rect 12365 7894 12369 7914
rect 9350 7832 9385 7833
rect 7380 7712 7436 7719
rect 8315 7712 9272 7731
rect 9329 7825 9385 7832
rect 9329 7805 9358 7825
rect 9378 7805 9385 7825
rect 9329 7800 9385 7805
rect 9559 7827 9599 7839
rect 9559 7806 9565 7827
rect 9587 7806 9599 7827
rect 9559 7801 9599 7806
rect 9776 7828 9808 7835
rect 9776 7808 9782 7828
rect 9803 7808 9808 7828
rect 7380 7711 7415 7712
rect 7166 7676 7201 7705
rect 7166 7675 7476 7676
rect 7051 7669 7087 7673
rect 7051 7650 7059 7669
rect 7079 7650 7087 7669
rect 7051 7647 7087 7650
rect 7052 7619 7086 7647
rect 7166 7641 7493 7675
rect 6144 7481 6156 7502
rect 6178 7481 6194 7502
rect 6144 7473 6194 7481
rect 6367 7505 6423 7510
rect 6367 7485 6374 7505
rect 6394 7485 6423 7505
rect 6367 7478 6423 7485
rect 6524 7591 7087 7619
rect 6367 7477 6402 7478
rect 3433 7441 3437 7461
rect 3458 7441 3465 7461
rect 3433 7434 3465 7441
rect 6149 7440 6190 7473
rect 6524 7440 6564 7591
rect 6149 7411 6564 7440
rect 7453 7417 7493 7641
rect 8154 7660 8183 7662
rect 8154 7655 8527 7660
rect 8154 7637 8161 7655
rect 8181 7637 8527 7655
rect 8154 7632 8527 7637
rect 8159 7630 8527 7632
rect 8288 7593 8323 7594
rect 8503 7593 8527 7630
rect 6149 7410 6558 7411
rect 7453 7397 7463 7417
rect 7483 7397 7493 7417
rect 7453 7387 7493 7397
rect 8267 7586 8323 7593
rect 8267 7566 8296 7586
rect 8316 7566 8323 7586
rect 8267 7561 8323 7566
rect 8498 7588 8535 7593
rect 8498 7569 8506 7588
rect 8529 7569 8535 7588
rect 8498 7563 8535 7569
rect 8714 7589 8746 7596
rect 8714 7569 8720 7589
rect 8741 7569 8746 7589
rect 1942 7178 1951 7195
rect 1975 7178 1980 7195
rect 1942 7135 1980 7178
rect 2154 7199 2210 7204
rect 2154 7179 2161 7199
rect 2181 7179 2210 7199
rect 2154 7172 2210 7179
rect 2984 7368 3024 7378
rect 2984 7348 2994 7368
rect 3014 7348 3024 7368
rect 3919 7354 4328 7355
rect 2154 7171 2189 7172
rect 2288 7135 2372 7140
rect 1942 7106 2372 7135
rect 669 6937 674 6957
rect 695 6937 701 6957
rect 669 6930 701 6937
rect 878 6959 918 6964
rect 878 6938 890 6959
rect 912 6938 918 6959
rect 878 6926 918 6938
rect 1092 6960 1148 6965
rect 1092 6940 1099 6960
rect 1119 6940 1148 6960
rect 1092 6933 1148 6940
rect 1205 7034 2162 7053
rect 1092 6932 1127 6933
rect 884 6894 912 6926
rect 1205 6894 1236 7034
rect 2125 7018 2160 7034
rect 2125 6998 2132 7018
rect 2152 6998 2160 7018
rect 2125 6990 2160 6998
rect 884 6863 1236 6894
rect 1681 6925 1713 6932
rect 1681 6905 1688 6925
rect 1709 6905 1713 6925
rect 1681 6840 1713 6905
rect 2051 6840 2091 6841
rect 1681 6838 2093 6840
rect 1681 6812 2061 6838
rect 2087 6812 2093 6838
rect 1681 6804 2093 6812
rect 1115 6789 1147 6790
rect 1112 6784 1147 6789
rect 1112 6764 1119 6784
rect 1139 6764 1147 6784
rect 1112 6756 1147 6764
rect 668 6691 700 6698
rect 668 6671 675 6691
rect 696 6671 700 6691
rect 668 6606 700 6671
rect 1038 6606 1078 6607
rect 668 6604 1080 6606
rect 668 6578 1048 6604
rect 1074 6578 1080 6604
rect 668 6570 1080 6578
rect 668 6542 700 6570
rect 668 6522 673 6542
rect 694 6522 700 6542
rect 668 6515 700 6522
rect 868 6542 918 6551
rect 1113 6550 1147 6756
rect 1681 6776 1713 6804
rect 1681 6756 1686 6776
rect 1707 6756 1713 6776
rect 1886 6778 1928 6787
rect 2126 6784 2160 6990
rect 1886 6764 1896 6778
rect 1681 6749 1713 6756
rect 1885 6758 1896 6764
rect 1920 6758 1928 6778
rect 1885 6747 1928 6758
rect 2104 6779 2160 6784
rect 2104 6759 2111 6779
rect 2131 6759 2160 6779
rect 2104 6752 2160 6759
rect 2104 6751 2139 6752
rect 1885 6717 1925 6747
rect 1775 6709 1811 6713
rect 1775 6690 1783 6709
rect 1803 6690 1811 6709
rect 1775 6687 1811 6690
rect 1885 6712 2232 6717
rect 1776 6659 1810 6687
rect 1885 6686 2204 6712
rect 2223 6686 2232 6712
rect 1885 6682 2232 6686
rect 868 6521 880 6542
rect 902 6521 918 6542
rect 868 6513 918 6521
rect 1091 6545 1147 6550
rect 1091 6525 1098 6545
rect 1118 6525 1147 6545
rect 1091 6518 1147 6525
rect 1248 6631 1811 6659
rect 1091 6517 1126 6518
rect 873 6480 914 6513
rect 1248 6480 1288 6631
rect 2337 6512 2372 7106
rect 2984 7124 3024 7348
rect 3913 7325 4328 7354
rect 3913 7174 3953 7325
rect 4287 7292 4328 7325
rect 7012 7324 7044 7331
rect 7012 7304 7019 7324
rect 7040 7304 7044 7324
rect 4075 7287 4110 7288
rect 3390 7146 3953 7174
rect 4054 7280 4110 7287
rect 4054 7260 4083 7280
rect 4103 7260 4110 7280
rect 4054 7255 4110 7260
rect 4283 7284 4333 7292
rect 4283 7263 4299 7284
rect 4321 7263 4333 7284
rect 2984 7090 3311 7124
rect 3391 7118 3425 7146
rect 3390 7115 3426 7118
rect 3390 7096 3398 7115
rect 3418 7096 3426 7115
rect 3390 7092 3426 7096
rect 3001 7089 3311 7090
rect 3276 7060 3311 7089
rect 3062 7053 3097 7054
rect 3041 7046 3097 7053
rect 3041 7026 3070 7046
rect 3090 7026 3097 7046
rect 3041 7021 3097 7026
rect 3271 7048 3313 7060
rect 3271 7028 3280 7048
rect 3304 7028 3313 7048
rect 3041 6815 3075 7021
rect 3271 7020 3313 7028
rect 3488 7049 3520 7056
rect 3488 7029 3494 7049
rect 3515 7029 3520 7049
rect 3488 7001 3520 7029
rect 4054 7049 4088 7255
rect 4283 7254 4333 7263
rect 4501 7283 4533 7290
rect 4501 7263 4507 7283
rect 4528 7263 4533 7283
rect 4501 7235 4533 7263
rect 4121 7227 4533 7235
rect 4121 7201 4127 7227
rect 4153 7201 4533 7227
rect 4121 7199 4533 7201
rect 4123 7198 4163 7199
rect 4501 7134 4533 7199
rect 7012 7239 7044 7304
rect 7382 7239 7422 7240
rect 7012 7237 7424 7239
rect 7012 7211 7392 7237
rect 7418 7211 7424 7237
rect 7012 7203 7424 7211
rect 6397 7183 6429 7184
rect 6394 7178 6429 7183
rect 6394 7158 6401 7178
rect 6421 7158 6429 7178
rect 6394 7150 6429 7158
rect 4501 7114 4505 7134
rect 4526 7114 4533 7134
rect 4501 7107 4533 7114
rect 5950 7085 5982 7092
rect 5950 7065 5957 7085
rect 5978 7065 5982 7085
rect 4054 7041 4089 7049
rect 4054 7021 4062 7041
rect 4082 7021 4089 7041
rect 4054 7016 4089 7021
rect 4054 7015 4086 7016
rect 3108 6993 3520 7001
rect 3108 6967 3114 6993
rect 3140 6967 3520 6993
rect 3108 6965 3520 6967
rect 3110 6964 3150 6965
rect 3488 6900 3520 6965
rect 5950 7000 5982 7065
rect 6320 7000 6360 7001
rect 5950 6998 6362 7000
rect 5950 6972 6330 6998
rect 6356 6972 6362 6998
rect 5950 6964 6362 6972
rect 3488 6880 3492 6900
rect 3513 6880 3520 6900
rect 3488 6873 3520 6880
rect 3965 6911 4317 6942
rect 3041 6807 3076 6815
rect 3041 6787 3049 6807
rect 3069 6787 3076 6807
rect 3041 6771 3076 6787
rect 3965 6771 3996 6911
rect 4289 6879 4317 6911
rect 5950 6936 5982 6964
rect 6395 6944 6429 7150
rect 7012 7175 7044 7203
rect 7012 7155 7017 7175
rect 7038 7155 7044 7175
rect 7012 7148 7044 7155
rect 7223 7174 7261 7186
rect 7457 7183 7491 7387
rect 8267 7357 8301 7561
rect 8714 7541 8746 7569
rect 9329 7594 9363 7800
rect 9776 7780 9808 7808
rect 9396 7772 9808 7780
rect 12337 7829 12369 7894
rect 12707 7829 12747 7830
rect 12337 7827 12749 7829
rect 12337 7801 12717 7827
rect 12743 7801 12749 7827
rect 12337 7793 12749 7801
rect 11771 7778 11803 7779
rect 9396 7746 9402 7772
rect 9428 7746 9808 7772
rect 9396 7744 9808 7746
rect 11768 7773 11803 7778
rect 11768 7753 11775 7773
rect 11795 7753 11803 7773
rect 11768 7745 11803 7753
rect 9398 7743 9438 7744
rect 9776 7679 9808 7744
rect 9776 7659 9780 7679
rect 9801 7659 9808 7679
rect 9776 7652 9808 7659
rect 11324 7680 11356 7687
rect 11324 7660 11331 7680
rect 11352 7660 11356 7680
rect 11324 7595 11356 7660
rect 11694 7595 11734 7596
rect 9329 7586 9364 7594
rect 9329 7566 9337 7586
rect 9357 7566 9364 7586
rect 9329 7561 9364 7566
rect 11324 7593 11736 7595
rect 11324 7567 11704 7593
rect 11730 7567 11736 7593
rect 9329 7560 9361 7561
rect 8334 7533 8746 7541
rect 8334 7507 8340 7533
rect 8366 7507 8746 7533
rect 8334 7505 8746 7507
rect 8336 7504 8376 7505
rect 8714 7440 8746 7505
rect 11324 7559 11736 7567
rect 11324 7531 11356 7559
rect 11324 7511 11329 7531
rect 11350 7511 11356 7531
rect 11324 7504 11356 7511
rect 11524 7531 11574 7540
rect 11769 7539 11803 7745
rect 12337 7765 12369 7793
rect 12337 7745 12342 7765
rect 12363 7745 12369 7765
rect 12337 7738 12369 7745
rect 12544 7766 12586 7774
rect 12782 7773 12816 7979
rect 12544 7746 12553 7766
rect 12577 7746 12586 7766
rect 12544 7734 12586 7746
rect 12760 7768 12816 7773
rect 12760 7748 12767 7768
rect 12787 7748 12816 7768
rect 13697 8015 13726 8035
rect 13746 8015 13753 8035
rect 13697 8010 13753 8015
rect 13929 8036 13972 8047
rect 13929 8016 13937 8036
rect 13961 8030 13972 8036
rect 14144 8038 14176 8045
rect 13961 8016 13971 8030
rect 13697 7804 13731 8010
rect 13929 8007 13971 8016
rect 14144 8018 14150 8038
rect 14171 8018 14176 8038
rect 14144 7990 14176 8018
rect 14710 8038 14744 8244
rect 14939 8243 14989 8252
rect 15157 8272 15189 8279
rect 15157 8252 15163 8272
rect 15184 8252 15189 8272
rect 15157 8224 15189 8252
rect 14777 8216 15189 8224
rect 14777 8190 14783 8216
rect 14809 8190 15189 8216
rect 14777 8188 15189 8190
rect 14779 8187 14819 8188
rect 15157 8123 15189 8188
rect 17053 8172 17085 8173
rect 17050 8167 17085 8172
rect 17050 8147 17057 8167
rect 17077 8147 17085 8167
rect 17050 8139 17085 8147
rect 19850 8142 19890 8293
rect 20224 8260 20265 8293
rect 20012 8255 20047 8256
rect 15157 8103 15161 8123
rect 15182 8103 15189 8123
rect 15157 8096 15189 8103
rect 16606 8074 16638 8081
rect 16606 8054 16613 8074
rect 16634 8054 16638 8074
rect 14710 8030 14745 8038
rect 14710 8010 14718 8030
rect 14738 8010 14745 8030
rect 14710 8005 14745 8010
rect 14710 8004 14742 8005
rect 13764 7982 14176 7990
rect 13764 7956 13770 7982
rect 13796 7956 14176 7982
rect 13764 7954 14176 7956
rect 13766 7953 13806 7954
rect 14144 7889 14176 7954
rect 16606 7989 16638 8054
rect 16976 7989 17016 7990
rect 16606 7987 17018 7989
rect 16606 7961 16986 7987
rect 17012 7961 17018 7987
rect 16606 7953 17018 7961
rect 14144 7869 14148 7889
rect 14169 7869 14176 7889
rect 14144 7862 14176 7869
rect 14621 7900 14973 7931
rect 13697 7796 13732 7804
rect 13697 7776 13705 7796
rect 13725 7776 13732 7796
rect 13697 7760 13732 7776
rect 14621 7760 14652 7900
rect 14945 7868 14973 7900
rect 16606 7925 16638 7953
rect 17051 7933 17085 8139
rect 19327 8114 19890 8142
rect 19991 8248 20047 8255
rect 19991 8228 20020 8248
rect 20040 8228 20047 8248
rect 19991 8223 20047 8228
rect 20220 8252 20270 8260
rect 20220 8231 20236 8252
rect 20258 8231 20270 8252
rect 18906 8087 19253 8091
rect 18906 8061 18915 8087
rect 18934 8061 19253 8087
rect 19328 8086 19362 8114
rect 18906 8056 19253 8061
rect 19327 8083 19363 8086
rect 19327 8064 19335 8083
rect 19355 8064 19363 8083
rect 19327 8060 19363 8064
rect 19213 8026 19253 8056
rect 18999 8021 19034 8022
rect 16606 7905 16611 7925
rect 16632 7905 16638 7925
rect 16606 7898 16638 7905
rect 16815 7927 16855 7932
rect 16815 7906 16827 7927
rect 16849 7906 16855 7927
rect 16815 7894 16855 7906
rect 17029 7928 17085 7933
rect 17029 7908 17036 7928
rect 17056 7908 17085 7928
rect 17029 7901 17085 7908
rect 17142 8002 18099 8021
rect 18978 8014 19034 8021
rect 17029 7900 17064 7901
rect 14730 7861 14765 7862
rect 12760 7741 12816 7748
rect 13695 7741 14652 7760
rect 14709 7854 14765 7861
rect 14709 7834 14738 7854
rect 14758 7834 14765 7854
rect 14709 7829 14765 7834
rect 14939 7856 14979 7868
rect 14939 7835 14945 7856
rect 14967 7835 14979 7856
rect 14939 7830 14979 7835
rect 15156 7857 15188 7864
rect 15156 7837 15162 7857
rect 15183 7837 15188 7857
rect 12760 7740 12795 7741
rect 12546 7705 12581 7734
rect 12546 7704 12856 7705
rect 12431 7698 12467 7702
rect 12431 7679 12439 7698
rect 12459 7679 12467 7698
rect 12431 7676 12467 7679
rect 12432 7648 12466 7676
rect 12546 7670 12873 7704
rect 11524 7510 11536 7531
rect 11558 7510 11574 7531
rect 11524 7502 11574 7510
rect 11747 7534 11803 7539
rect 11747 7514 11754 7534
rect 11774 7514 11803 7534
rect 11747 7507 11803 7514
rect 11904 7620 12467 7648
rect 11747 7506 11782 7507
rect 8714 7420 8718 7440
rect 8739 7420 8746 7440
rect 11529 7469 11570 7502
rect 11904 7469 11944 7620
rect 11529 7440 11944 7469
rect 12833 7446 12873 7670
rect 13534 7689 13563 7691
rect 13534 7684 13907 7689
rect 13534 7666 13541 7684
rect 13561 7666 13907 7684
rect 13534 7661 13907 7666
rect 13539 7659 13907 7661
rect 13668 7622 13703 7623
rect 13883 7622 13907 7659
rect 11529 7439 11938 7440
rect 8714 7413 8746 7420
rect 12833 7426 12843 7446
rect 12863 7426 12873 7446
rect 12833 7416 12873 7426
rect 13647 7615 13703 7622
rect 13647 7595 13676 7615
rect 13696 7595 13703 7615
rect 13647 7590 13703 7595
rect 13878 7617 13915 7622
rect 13878 7598 13886 7617
rect 13909 7598 13915 7617
rect 13878 7592 13915 7598
rect 14094 7618 14126 7625
rect 14094 7598 14100 7618
rect 14121 7598 14126 7618
rect 7223 7157 7232 7174
rect 7256 7157 7261 7174
rect 7223 7114 7261 7157
rect 7435 7178 7491 7183
rect 7435 7158 7442 7178
rect 7462 7158 7491 7178
rect 7435 7151 7491 7158
rect 8265 7347 8305 7357
rect 8265 7327 8275 7347
rect 8295 7327 8305 7347
rect 12392 7353 12424 7360
rect 9200 7333 9609 7334
rect 7435 7150 7470 7151
rect 7569 7114 7653 7119
rect 7223 7085 7653 7114
rect 5950 6916 5955 6936
rect 5976 6916 5982 6936
rect 5950 6909 5982 6916
rect 6159 6938 6199 6943
rect 6159 6917 6171 6938
rect 6193 6917 6199 6938
rect 6159 6905 6199 6917
rect 6373 6939 6429 6944
rect 6373 6919 6380 6939
rect 6400 6919 6429 6939
rect 6373 6912 6429 6919
rect 6486 7013 7443 7032
rect 6373 6911 6408 6912
rect 4074 6872 4109 6873
rect 3039 6752 3996 6771
rect 4053 6865 4109 6872
rect 4053 6845 4082 6865
rect 4102 6845 4109 6865
rect 4053 6840 4109 6845
rect 4283 6867 4323 6879
rect 4283 6846 4289 6867
rect 4311 6846 4323 6867
rect 4283 6841 4323 6846
rect 4500 6868 4532 6875
rect 4500 6848 4506 6868
rect 4527 6848 4532 6868
rect 2749 6654 2786 6659
rect 2749 6648 3096 6654
rect 2749 6629 2757 6648
rect 2780 6629 3096 6648
rect 2749 6624 3096 6629
rect 2749 6618 2786 6624
rect 3066 6593 3096 6624
rect 4053 6634 4087 6840
rect 4500 6820 4532 6848
rect 6165 6873 6193 6905
rect 6486 6873 6517 7013
rect 7406 6997 7441 7013
rect 7406 6977 7413 6997
rect 7433 6977 7441 6997
rect 7406 6969 7441 6977
rect 6165 6842 6517 6873
rect 6962 6904 6994 6911
rect 6962 6884 6969 6904
rect 6990 6884 6994 6904
rect 4120 6812 4532 6820
rect 4120 6786 4126 6812
rect 4152 6786 4532 6812
rect 4120 6784 4532 6786
rect 4122 6783 4162 6784
rect 4500 6719 4532 6784
rect 6962 6819 6994 6884
rect 7332 6819 7372 6820
rect 6962 6817 7374 6819
rect 6962 6791 7342 6817
rect 7368 6791 7374 6817
rect 6962 6783 7374 6791
rect 6396 6768 6428 6769
rect 6393 6763 6428 6768
rect 6393 6743 6400 6763
rect 6420 6743 6428 6763
rect 6393 6735 6428 6743
rect 4500 6699 4504 6719
rect 4525 6699 4532 6719
rect 4500 6692 4532 6699
rect 5949 6670 5981 6677
rect 5949 6650 5956 6670
rect 5977 6650 5981 6670
rect 4053 6626 4088 6634
rect 4053 6606 4061 6626
rect 4081 6606 4088 6626
rect 4053 6601 4088 6606
rect 4053 6600 4085 6601
rect 2854 6586 2889 6587
rect 2833 6579 2889 6586
rect 2833 6559 2862 6579
rect 2882 6559 2889 6579
rect 2833 6554 2889 6559
rect 3064 6580 3103 6593
rect 3064 6561 3069 6580
rect 3092 6561 3103 6580
rect 3064 6555 3103 6561
rect 3280 6582 3312 6589
rect 3280 6562 3286 6582
rect 3307 6562 3312 6582
rect 2337 6506 2375 6512
rect 2337 6486 2347 6506
rect 2367 6486 2375 6506
rect 2337 6484 2375 6486
rect 873 6451 1288 6480
rect 2340 6478 2375 6484
rect 873 6450 1282 6451
rect 1896 6413 1928 6420
rect 1896 6393 1903 6413
rect 1924 6393 1928 6413
rect 1896 6328 1928 6393
rect 2266 6328 2306 6329
rect 1896 6326 2308 6328
rect 1896 6300 2276 6326
rect 2302 6300 2308 6326
rect 1896 6292 2308 6300
rect 1896 6264 1928 6292
rect 1896 6244 1901 6264
rect 1922 6244 1928 6264
rect 1896 6237 1928 6244
rect 2100 6269 2147 6275
rect 2341 6272 2375 6478
rect 2833 6348 2867 6554
rect 3280 6534 3312 6562
rect 2900 6526 3312 6534
rect 2900 6500 2906 6526
rect 2932 6500 3312 6526
rect 2900 6498 3312 6500
rect 2902 6497 2942 6498
rect 3280 6433 3312 6498
rect 5949 6585 5981 6650
rect 6319 6585 6359 6586
rect 5949 6583 6361 6585
rect 5949 6557 6329 6583
rect 6355 6557 6361 6583
rect 5949 6549 6361 6557
rect 5949 6521 5981 6549
rect 5949 6501 5954 6521
rect 5975 6501 5981 6521
rect 5949 6494 5981 6501
rect 6149 6521 6199 6530
rect 6394 6529 6428 6735
rect 6962 6755 6994 6783
rect 6962 6735 6967 6755
rect 6988 6735 6994 6755
rect 7167 6757 7209 6766
rect 7407 6763 7441 6969
rect 7167 6743 7177 6757
rect 6962 6728 6994 6735
rect 7166 6737 7177 6743
rect 7201 6737 7209 6757
rect 7166 6726 7209 6737
rect 7385 6758 7441 6763
rect 7385 6738 7392 6758
rect 7412 6738 7441 6758
rect 7385 6731 7441 6738
rect 7385 6730 7420 6731
rect 7166 6696 7206 6726
rect 7056 6688 7092 6692
rect 7056 6669 7064 6688
rect 7084 6669 7092 6688
rect 7056 6666 7092 6669
rect 7166 6691 7513 6696
rect 7057 6638 7091 6666
rect 7166 6665 7485 6691
rect 7504 6665 7513 6691
rect 7166 6661 7513 6665
rect 6149 6500 6161 6521
rect 6183 6500 6199 6521
rect 6149 6492 6199 6500
rect 6372 6524 6428 6529
rect 6372 6504 6379 6524
rect 6399 6504 6428 6524
rect 6372 6497 6428 6504
rect 6529 6610 7092 6638
rect 6372 6496 6407 6497
rect 3280 6413 3284 6433
rect 3305 6413 3312 6433
rect 6154 6459 6195 6492
rect 6529 6459 6569 6610
rect 7618 6491 7653 7085
rect 8265 7103 8305 7327
rect 9194 7304 9609 7333
rect 9194 7153 9234 7304
rect 9568 7271 9609 7304
rect 12392 7333 12399 7353
rect 12420 7333 12424 7353
rect 9356 7266 9391 7267
rect 8671 7125 9234 7153
rect 9335 7259 9391 7266
rect 9335 7239 9364 7259
rect 9384 7239 9391 7259
rect 9335 7234 9391 7239
rect 9564 7263 9614 7271
rect 9564 7242 9580 7263
rect 9602 7242 9614 7263
rect 8265 7069 8592 7103
rect 8672 7097 8706 7125
rect 8671 7094 8707 7097
rect 8671 7075 8679 7094
rect 8699 7075 8707 7094
rect 8671 7071 8707 7075
rect 8282 7068 8592 7069
rect 8557 7039 8592 7068
rect 8343 7032 8378 7033
rect 8322 7025 8378 7032
rect 8322 7005 8351 7025
rect 8371 7005 8378 7025
rect 8322 7000 8378 7005
rect 8552 7027 8594 7039
rect 8552 7007 8561 7027
rect 8585 7007 8594 7027
rect 8322 6794 8356 7000
rect 8552 6999 8594 7007
rect 8769 7028 8801 7035
rect 8769 7008 8775 7028
rect 8796 7008 8801 7028
rect 8769 6980 8801 7008
rect 9335 7028 9369 7234
rect 9564 7233 9614 7242
rect 9782 7262 9814 7269
rect 9782 7242 9788 7262
rect 9809 7242 9814 7262
rect 9782 7214 9814 7242
rect 9402 7206 9814 7214
rect 12392 7268 12424 7333
rect 12762 7268 12802 7269
rect 12392 7266 12804 7268
rect 12392 7240 12772 7266
rect 12798 7240 12804 7266
rect 12392 7232 12804 7240
rect 11777 7212 11809 7213
rect 9402 7180 9408 7206
rect 9434 7180 9814 7206
rect 9402 7178 9814 7180
rect 11774 7207 11809 7212
rect 11774 7187 11781 7207
rect 11801 7187 11809 7207
rect 11774 7179 11809 7187
rect 9404 7177 9444 7178
rect 9782 7113 9814 7178
rect 9782 7093 9786 7113
rect 9807 7093 9814 7113
rect 9782 7086 9814 7093
rect 11330 7114 11362 7121
rect 11330 7094 11337 7114
rect 11358 7094 11362 7114
rect 11330 7029 11362 7094
rect 11700 7029 11740 7030
rect 9335 7020 9370 7028
rect 9335 7000 9343 7020
rect 9363 7000 9370 7020
rect 9335 6995 9370 7000
rect 11330 7027 11742 7029
rect 11330 7001 11710 7027
rect 11736 7001 11742 7027
rect 9335 6994 9367 6995
rect 8389 6972 8801 6980
rect 8389 6946 8395 6972
rect 8421 6946 8801 6972
rect 8389 6944 8801 6946
rect 8391 6943 8431 6944
rect 8769 6879 8801 6944
rect 11330 6993 11742 7001
rect 11330 6965 11362 6993
rect 11775 6973 11809 7179
rect 12392 7204 12424 7232
rect 12392 7184 12397 7204
rect 12418 7184 12424 7204
rect 12392 7177 12424 7184
rect 12603 7203 12641 7215
rect 12837 7212 12871 7416
rect 13647 7386 13681 7590
rect 14094 7570 14126 7598
rect 14709 7623 14743 7829
rect 15156 7809 15188 7837
rect 16821 7862 16849 7894
rect 17142 7862 17173 8002
rect 18062 7986 18097 8002
rect 18062 7966 18069 7986
rect 18089 7966 18097 7986
rect 18062 7958 18097 7966
rect 16821 7831 17173 7862
rect 17618 7893 17650 7900
rect 17618 7873 17625 7893
rect 17646 7873 17650 7893
rect 14776 7801 15188 7809
rect 14776 7775 14782 7801
rect 14808 7775 15188 7801
rect 14776 7773 15188 7775
rect 14778 7772 14818 7773
rect 15156 7708 15188 7773
rect 17618 7808 17650 7873
rect 17988 7808 18028 7809
rect 17618 7806 18030 7808
rect 17618 7780 17998 7806
rect 18024 7780 18030 7806
rect 17618 7772 18030 7780
rect 17052 7757 17084 7758
rect 17049 7752 17084 7757
rect 17049 7732 17056 7752
rect 17076 7732 17084 7752
rect 17049 7724 17084 7732
rect 15156 7688 15160 7708
rect 15181 7688 15188 7708
rect 15156 7681 15188 7688
rect 16605 7659 16637 7666
rect 16605 7639 16612 7659
rect 16633 7639 16637 7659
rect 14709 7615 14744 7623
rect 14709 7595 14717 7615
rect 14737 7595 14744 7615
rect 14709 7590 14744 7595
rect 14709 7589 14741 7590
rect 13714 7562 14126 7570
rect 13714 7536 13720 7562
rect 13746 7536 14126 7562
rect 13714 7534 14126 7536
rect 13716 7533 13756 7534
rect 14094 7469 14126 7534
rect 16605 7574 16637 7639
rect 16975 7574 17015 7575
rect 16605 7572 17017 7574
rect 16605 7546 16985 7572
rect 17011 7546 17017 7572
rect 16605 7538 17017 7546
rect 16605 7510 16637 7538
rect 16605 7490 16610 7510
rect 16631 7490 16637 7510
rect 16605 7483 16637 7490
rect 16805 7510 16855 7519
rect 17050 7518 17084 7724
rect 17618 7744 17650 7772
rect 17618 7724 17623 7744
rect 17644 7724 17650 7744
rect 17618 7717 17650 7724
rect 17825 7745 17867 7753
rect 18063 7752 18097 7958
rect 17825 7725 17834 7745
rect 17858 7725 17867 7745
rect 17825 7713 17867 7725
rect 18041 7747 18097 7752
rect 18041 7727 18048 7747
rect 18068 7727 18097 7747
rect 18978 7994 19007 8014
rect 19027 7994 19034 8014
rect 18978 7989 19034 7994
rect 19210 8015 19253 8026
rect 19210 7995 19218 8015
rect 19242 8009 19253 8015
rect 19425 8017 19457 8024
rect 19242 7995 19252 8009
rect 18978 7783 19012 7989
rect 19210 7986 19252 7995
rect 19425 7997 19431 8017
rect 19452 7997 19457 8017
rect 19425 7969 19457 7997
rect 19991 8017 20025 8223
rect 20220 8222 20270 8231
rect 20438 8251 20470 8258
rect 20438 8231 20444 8251
rect 20465 8231 20470 8251
rect 20438 8203 20470 8231
rect 20058 8195 20470 8203
rect 20058 8169 20064 8195
rect 20090 8169 20470 8195
rect 20058 8167 20470 8169
rect 20060 8166 20100 8167
rect 20438 8102 20470 8167
rect 20438 8082 20442 8102
rect 20463 8082 20470 8102
rect 20438 8075 20470 8082
rect 19991 8009 20026 8017
rect 19991 7989 19999 8009
rect 20019 7989 20026 8009
rect 19991 7984 20026 7989
rect 19991 7983 20023 7984
rect 19045 7961 19457 7969
rect 19045 7935 19051 7961
rect 19077 7935 19457 7961
rect 19045 7933 19457 7935
rect 19047 7932 19087 7933
rect 19425 7868 19457 7933
rect 19425 7848 19429 7868
rect 19450 7848 19457 7868
rect 19425 7841 19457 7848
rect 19902 7879 20254 7910
rect 18978 7775 19013 7783
rect 18978 7755 18986 7775
rect 19006 7755 19013 7775
rect 18978 7739 19013 7755
rect 19902 7739 19933 7879
rect 20226 7847 20254 7879
rect 20011 7840 20046 7841
rect 18041 7720 18097 7727
rect 18976 7720 19933 7739
rect 19990 7833 20046 7840
rect 19990 7813 20019 7833
rect 20039 7813 20046 7833
rect 19990 7808 20046 7813
rect 20220 7835 20260 7847
rect 20220 7814 20226 7835
rect 20248 7814 20260 7835
rect 20220 7809 20260 7814
rect 20437 7836 20469 7843
rect 20437 7816 20443 7836
rect 20464 7816 20469 7836
rect 18041 7719 18076 7720
rect 17827 7684 17862 7713
rect 17827 7683 18137 7684
rect 17712 7677 17748 7681
rect 17712 7658 17720 7677
rect 17740 7658 17748 7677
rect 17712 7655 17748 7658
rect 17713 7627 17747 7655
rect 17827 7649 18154 7683
rect 16805 7489 16817 7510
rect 16839 7489 16855 7510
rect 16805 7481 16855 7489
rect 17028 7513 17084 7518
rect 17028 7493 17035 7513
rect 17055 7493 17084 7513
rect 17028 7486 17084 7493
rect 17185 7599 17748 7627
rect 17028 7485 17063 7486
rect 14094 7449 14098 7469
rect 14119 7449 14126 7469
rect 14094 7442 14126 7449
rect 16810 7448 16851 7481
rect 17185 7448 17225 7599
rect 16810 7419 17225 7448
rect 18114 7425 18154 7649
rect 18815 7668 18844 7670
rect 18815 7663 19188 7668
rect 18815 7645 18822 7663
rect 18842 7645 19188 7663
rect 18815 7640 19188 7645
rect 18820 7638 19188 7640
rect 18949 7601 18984 7602
rect 19164 7601 19188 7638
rect 16810 7418 17219 7419
rect 18114 7405 18124 7425
rect 18144 7405 18154 7425
rect 18114 7395 18154 7405
rect 18928 7594 18984 7601
rect 18928 7574 18957 7594
rect 18977 7574 18984 7594
rect 18928 7569 18984 7574
rect 19159 7596 19196 7601
rect 19159 7577 19167 7596
rect 19190 7577 19196 7596
rect 19159 7571 19196 7577
rect 19375 7597 19407 7604
rect 19375 7577 19381 7597
rect 19402 7577 19407 7597
rect 12603 7186 12612 7203
rect 12636 7186 12641 7203
rect 12603 7143 12641 7186
rect 12815 7207 12871 7212
rect 12815 7187 12822 7207
rect 12842 7187 12871 7207
rect 12815 7180 12871 7187
rect 13645 7376 13685 7386
rect 13645 7356 13655 7376
rect 13675 7356 13685 7376
rect 14580 7362 14989 7363
rect 12815 7179 12850 7180
rect 12949 7143 13033 7148
rect 12603 7114 13033 7143
rect 11330 6945 11335 6965
rect 11356 6945 11362 6965
rect 11330 6938 11362 6945
rect 11539 6967 11579 6972
rect 11539 6946 11551 6967
rect 11573 6946 11579 6967
rect 11539 6934 11579 6946
rect 11753 6968 11809 6973
rect 11753 6948 11760 6968
rect 11780 6948 11809 6968
rect 11753 6941 11809 6948
rect 11866 7042 12823 7061
rect 11753 6940 11788 6941
rect 8769 6859 8773 6879
rect 8794 6859 8801 6879
rect 8769 6852 8801 6859
rect 9246 6890 9598 6921
rect 8322 6786 8357 6794
rect 8322 6766 8330 6786
rect 8350 6766 8357 6786
rect 8322 6750 8357 6766
rect 9246 6750 9277 6890
rect 9570 6858 9598 6890
rect 11545 6902 11573 6934
rect 11866 6902 11897 7042
rect 12786 7026 12821 7042
rect 12786 7006 12793 7026
rect 12813 7006 12821 7026
rect 12786 6998 12821 7006
rect 11545 6871 11897 6902
rect 12342 6933 12374 6940
rect 12342 6913 12349 6933
rect 12370 6913 12374 6933
rect 9355 6851 9390 6852
rect 8320 6731 9277 6750
rect 9334 6844 9390 6851
rect 9334 6824 9363 6844
rect 9383 6824 9390 6844
rect 9334 6819 9390 6824
rect 9564 6846 9604 6858
rect 9564 6825 9570 6846
rect 9592 6825 9604 6846
rect 9564 6820 9604 6825
rect 9781 6847 9813 6854
rect 9781 6827 9787 6847
rect 9808 6827 9813 6847
rect 8030 6633 8067 6638
rect 8030 6627 8377 6633
rect 8030 6608 8038 6627
rect 8061 6608 8377 6627
rect 8030 6603 8377 6608
rect 8030 6597 8067 6603
rect 8347 6572 8377 6603
rect 9334 6613 9368 6819
rect 9781 6799 9813 6827
rect 9401 6791 9813 6799
rect 12342 6848 12374 6913
rect 12712 6848 12752 6849
rect 12342 6846 12754 6848
rect 12342 6820 12722 6846
rect 12748 6820 12754 6846
rect 12342 6812 12754 6820
rect 11776 6797 11808 6798
rect 9401 6765 9407 6791
rect 9433 6765 9813 6791
rect 9401 6763 9813 6765
rect 11773 6792 11808 6797
rect 11773 6772 11780 6792
rect 11800 6772 11808 6792
rect 11773 6764 11808 6772
rect 9403 6762 9443 6763
rect 9781 6698 9813 6763
rect 9781 6678 9785 6698
rect 9806 6678 9813 6698
rect 9781 6671 9813 6678
rect 11329 6699 11361 6706
rect 11329 6679 11336 6699
rect 11357 6679 11361 6699
rect 11329 6614 11361 6679
rect 11699 6614 11739 6615
rect 9334 6605 9369 6613
rect 9334 6585 9342 6605
rect 9362 6585 9369 6605
rect 9334 6580 9369 6585
rect 11329 6612 11741 6614
rect 11329 6586 11709 6612
rect 11735 6586 11741 6612
rect 9334 6579 9366 6580
rect 11329 6578 11741 6586
rect 8135 6565 8170 6566
rect 8114 6558 8170 6565
rect 8114 6538 8143 6558
rect 8163 6538 8170 6558
rect 8114 6533 8170 6538
rect 8345 6559 8384 6572
rect 8345 6540 8350 6559
rect 8373 6540 8384 6559
rect 8345 6534 8384 6540
rect 8561 6561 8593 6568
rect 8561 6541 8567 6561
rect 8588 6541 8593 6561
rect 7618 6485 7656 6491
rect 7618 6465 7628 6485
rect 7648 6465 7656 6485
rect 7618 6463 7656 6465
rect 6154 6430 6569 6459
rect 7621 6457 7656 6463
rect 6154 6429 6563 6430
rect 3280 6406 3312 6413
rect 7177 6392 7209 6399
rect 3926 6375 4335 6376
rect 2833 6342 2868 6348
rect 3920 6346 4335 6375
rect 2833 6340 2871 6342
rect 2833 6320 2841 6340
rect 2861 6320 2871 6340
rect 2833 6314 2871 6320
rect 2100 6243 2110 6269
rect 2135 6243 2147 6269
rect 2100 6241 2147 6243
rect 2319 6267 2375 6272
rect 2319 6247 2326 6267
rect 2346 6247 2375 6267
rect 1123 6225 1155 6226
rect 1120 6220 1155 6225
rect 1120 6200 1127 6220
rect 1147 6200 1155 6220
rect 1120 6192 1155 6200
rect 676 6127 708 6134
rect 676 6107 683 6127
rect 704 6107 708 6127
rect 676 6042 708 6107
rect 1046 6042 1086 6043
rect 676 6040 1088 6042
rect 676 6014 1056 6040
rect 1082 6014 1088 6040
rect 676 6006 1088 6014
rect 676 5978 708 6006
rect 1121 5986 1155 6192
rect 2105 6206 2142 6241
rect 2319 6240 2375 6247
rect 2319 6239 2354 6240
rect 2439 6206 2471 6208
rect 2105 6173 2475 6206
rect 676 5958 681 5978
rect 702 5958 708 5978
rect 676 5951 708 5958
rect 885 5980 925 5985
rect 885 5959 897 5980
rect 919 5959 925 5980
rect 885 5947 925 5959
rect 1099 5981 1155 5986
rect 1099 5961 1106 5981
rect 1126 5961 1155 5981
rect 1099 5954 1155 5961
rect 1212 6055 2169 6074
rect 1099 5953 1134 5954
rect 891 5915 919 5947
rect 1212 5915 1243 6055
rect 2132 6039 2167 6055
rect 2132 6019 2139 6039
rect 2159 6019 2167 6039
rect 2132 6011 2167 6019
rect 891 5884 1243 5915
rect 1688 5946 1720 5953
rect 1688 5926 1695 5946
rect 1716 5926 1720 5946
rect 1688 5861 1720 5926
rect 2058 5861 2098 5862
rect 1688 5859 2100 5861
rect 1688 5833 2068 5859
rect 2094 5833 2100 5859
rect 1688 5825 2100 5833
rect 1122 5810 1154 5811
rect 1119 5805 1154 5810
rect 1119 5785 1126 5805
rect 1146 5785 1154 5805
rect 1119 5777 1154 5785
rect 675 5712 707 5719
rect 675 5692 682 5712
rect 703 5692 707 5712
rect 675 5627 707 5692
rect 1045 5627 1085 5628
rect 675 5625 1087 5627
rect 675 5599 1055 5625
rect 1081 5599 1087 5625
rect 675 5591 1087 5599
rect 675 5563 707 5591
rect 675 5543 680 5563
rect 701 5543 707 5563
rect 675 5536 707 5543
rect 875 5563 925 5572
rect 1120 5571 1154 5777
rect 1688 5797 1720 5825
rect 1688 5777 1693 5797
rect 1714 5777 1720 5797
rect 1688 5770 1720 5777
rect 1895 5798 1937 5806
rect 2133 5805 2167 6011
rect 1895 5778 1904 5798
rect 1928 5778 1937 5798
rect 1895 5766 1937 5778
rect 2111 5800 2167 5805
rect 2111 5780 2118 5800
rect 2138 5780 2167 5800
rect 2111 5773 2167 5780
rect 2111 5772 2146 5773
rect 1897 5737 1932 5766
rect 1897 5736 2207 5737
rect 1782 5730 1818 5734
rect 1782 5711 1790 5730
rect 1810 5711 1818 5730
rect 1782 5708 1818 5711
rect 1783 5680 1817 5708
rect 1897 5702 2224 5736
rect 875 5542 887 5563
rect 909 5542 925 5563
rect 875 5534 925 5542
rect 1098 5566 1154 5571
rect 1098 5546 1105 5566
rect 1125 5546 1154 5566
rect 1098 5539 1154 5546
rect 1255 5652 1818 5680
rect 1098 5538 1133 5539
rect 880 5501 921 5534
rect 1255 5501 1295 5652
rect 880 5472 1295 5501
rect 2184 5478 2224 5702
rect 880 5471 1289 5472
rect 2184 5458 2194 5478
rect 2214 5458 2224 5478
rect 2184 5448 2224 5458
rect 1743 5385 1775 5392
rect 1743 5365 1750 5385
rect 1771 5365 1775 5385
rect 1743 5300 1775 5365
rect 2113 5300 2153 5301
rect 1743 5298 2155 5300
rect 1743 5272 2123 5298
rect 2149 5272 2155 5298
rect 1743 5264 2155 5272
rect 1128 5244 1160 5245
rect 1125 5239 1160 5244
rect 1125 5219 1132 5239
rect 1152 5219 1160 5239
rect 1125 5211 1160 5219
rect 681 5146 713 5153
rect 681 5126 688 5146
rect 709 5126 713 5146
rect 681 5061 713 5126
rect 1051 5061 1091 5062
rect 681 5059 1093 5061
rect 681 5033 1061 5059
rect 1087 5033 1093 5059
rect 681 5025 1093 5033
rect 681 4997 713 5025
rect 1126 5005 1160 5211
rect 1743 5236 1775 5264
rect 2188 5244 2222 5448
rect 1743 5216 1748 5236
rect 1769 5216 1775 5236
rect 1743 5209 1775 5216
rect 1954 5236 1991 5242
rect 1954 5217 1960 5236
rect 1983 5217 1991 5236
rect 1954 5212 1991 5217
rect 2166 5239 2222 5244
rect 2166 5219 2173 5239
rect 2193 5219 2222 5239
rect 2166 5212 2222 5219
rect 1962 5175 1986 5212
rect 2166 5211 2201 5212
rect 1962 5173 2330 5175
rect 1962 5168 2335 5173
rect 1962 5150 2308 5168
rect 2328 5150 2335 5168
rect 1962 5145 2335 5150
rect 2306 5143 2335 5145
rect 681 4977 686 4997
rect 707 4977 713 4997
rect 681 4970 713 4977
rect 890 4999 930 5004
rect 890 4978 902 4999
rect 924 4978 930 4999
rect 890 4966 930 4978
rect 1104 5000 1160 5005
rect 1104 4980 1111 5000
rect 1131 4980 1160 5000
rect 1104 4973 1160 4980
rect 1217 5074 2174 5093
rect 1104 4972 1139 4973
rect 896 4934 924 4966
rect 1217 4934 1248 5074
rect 2137 5058 2172 5074
rect 2137 5038 2144 5058
rect 2164 5038 2172 5058
rect 2137 5030 2172 5038
rect 896 4903 1248 4934
rect 1693 4965 1725 4972
rect 1693 4945 1700 4965
rect 1721 4945 1725 4965
rect 1693 4880 1725 4945
rect 2063 4880 2103 4881
rect 1693 4878 2105 4880
rect 1693 4852 2073 4878
rect 2099 4852 2105 4878
rect 1693 4844 2105 4852
rect 1127 4829 1159 4830
rect 1124 4824 1159 4829
rect 1124 4804 1131 4824
rect 1151 4804 1159 4824
rect 1124 4796 1159 4804
rect 680 4731 712 4738
rect 680 4711 687 4731
rect 708 4711 712 4731
rect 680 4646 712 4711
rect 1050 4646 1090 4647
rect 680 4644 1092 4646
rect 680 4618 1060 4644
rect 1086 4618 1092 4644
rect 680 4610 1092 4618
rect 680 4582 712 4610
rect 680 4562 685 4582
rect 706 4562 712 4582
rect 680 4555 712 4562
rect 880 4582 930 4591
rect 1125 4590 1159 4796
rect 1693 4816 1725 4844
rect 1693 4796 1698 4816
rect 1719 4796 1725 4816
rect 1898 4818 1940 4827
rect 2138 4824 2172 5030
rect 1898 4804 1908 4818
rect 1693 4789 1725 4796
rect 1897 4798 1908 4804
rect 1932 4798 1940 4818
rect 1897 4787 1940 4798
rect 2116 4819 2172 4824
rect 2116 4799 2123 4819
rect 2143 4799 2172 4819
rect 2116 4792 2172 4799
rect 2116 4791 2151 4792
rect 1897 4757 1937 4787
rect 1787 4749 1823 4753
rect 1787 4730 1795 4749
rect 1815 4730 1823 4749
rect 1787 4727 1823 4730
rect 1897 4752 2244 4757
rect 1788 4699 1822 4727
rect 1897 4726 2216 4752
rect 2235 4726 2244 4752
rect 1897 4722 2244 4726
rect 880 4561 892 4582
rect 914 4561 930 4582
rect 880 4553 930 4561
rect 1103 4585 1159 4590
rect 1103 4565 1110 4585
rect 1130 4565 1159 4585
rect 1103 4558 1159 4565
rect 1260 4671 1823 4699
rect 1103 4557 1138 4558
rect 885 4520 926 4553
rect 1260 4520 1300 4671
rect 2439 4520 2471 6173
rect 2836 5720 2871 6314
rect 3920 6195 3960 6346
rect 4294 6313 4335 6346
rect 7177 6372 7184 6392
rect 7205 6372 7209 6392
rect 4082 6308 4117 6309
rect 3397 6167 3960 6195
rect 4061 6301 4117 6308
rect 4061 6281 4090 6301
rect 4110 6281 4117 6301
rect 4061 6276 4117 6281
rect 4290 6305 4340 6313
rect 4290 6284 4306 6305
rect 4328 6284 4340 6305
rect 2976 6140 3323 6144
rect 2976 6114 2985 6140
rect 3004 6114 3323 6140
rect 3398 6139 3432 6167
rect 2976 6109 3323 6114
rect 3397 6136 3433 6139
rect 3397 6117 3405 6136
rect 3425 6117 3433 6136
rect 3397 6113 3433 6117
rect 3283 6079 3323 6109
rect 3069 6074 3104 6075
rect 3048 6067 3104 6074
rect 3048 6047 3077 6067
rect 3097 6047 3104 6067
rect 3048 6042 3104 6047
rect 3280 6068 3323 6079
rect 3280 6048 3288 6068
rect 3312 6062 3323 6068
rect 3495 6070 3527 6077
rect 3312 6048 3322 6062
rect 3048 5836 3082 6042
rect 3280 6039 3322 6048
rect 3495 6050 3501 6070
rect 3522 6050 3527 6070
rect 3495 6022 3527 6050
rect 4061 6070 4095 6276
rect 4290 6275 4340 6284
rect 4508 6304 4540 6311
rect 4508 6284 4514 6304
rect 4535 6284 4540 6304
rect 4508 6256 4540 6284
rect 4128 6248 4540 6256
rect 4128 6222 4134 6248
rect 4160 6222 4540 6248
rect 4128 6220 4540 6222
rect 4130 6219 4170 6220
rect 4508 6155 4540 6220
rect 7177 6307 7209 6372
rect 7547 6307 7587 6308
rect 7177 6305 7589 6307
rect 7177 6279 7557 6305
rect 7583 6279 7589 6305
rect 7177 6271 7589 6279
rect 7177 6243 7209 6271
rect 7177 6223 7182 6243
rect 7203 6223 7209 6243
rect 7177 6216 7209 6223
rect 7381 6248 7428 6254
rect 7622 6251 7656 6457
rect 8114 6327 8148 6533
rect 8561 6513 8593 6541
rect 11329 6550 11361 6578
rect 11329 6530 11334 6550
rect 11355 6530 11361 6550
rect 11329 6523 11361 6530
rect 11529 6550 11579 6559
rect 11774 6558 11808 6764
rect 12342 6784 12374 6812
rect 12342 6764 12347 6784
rect 12368 6764 12374 6784
rect 12547 6786 12589 6795
rect 12787 6792 12821 6998
rect 12547 6772 12557 6786
rect 12342 6757 12374 6764
rect 12546 6766 12557 6772
rect 12581 6766 12589 6786
rect 12546 6755 12589 6766
rect 12765 6787 12821 6792
rect 12765 6767 12772 6787
rect 12792 6767 12821 6787
rect 12765 6760 12821 6767
rect 12765 6759 12800 6760
rect 12546 6725 12586 6755
rect 12436 6717 12472 6721
rect 12436 6698 12444 6717
rect 12464 6698 12472 6717
rect 12436 6695 12472 6698
rect 12546 6720 12893 6725
rect 12437 6667 12471 6695
rect 12546 6694 12865 6720
rect 12884 6694 12893 6720
rect 12546 6690 12893 6694
rect 11529 6529 11541 6550
rect 11563 6529 11579 6550
rect 11529 6521 11579 6529
rect 11752 6553 11808 6558
rect 11752 6533 11759 6553
rect 11779 6533 11808 6553
rect 11752 6526 11808 6533
rect 11909 6639 12472 6667
rect 11752 6525 11787 6526
rect 8181 6505 8593 6513
rect 8181 6479 8187 6505
rect 8213 6479 8593 6505
rect 8181 6477 8593 6479
rect 8183 6476 8223 6477
rect 8561 6412 8593 6477
rect 11534 6488 11575 6521
rect 11909 6488 11949 6639
rect 12998 6520 13033 7114
rect 13645 7132 13685 7356
rect 14574 7333 14989 7362
rect 14574 7182 14614 7333
rect 14948 7300 14989 7333
rect 17673 7332 17705 7339
rect 17673 7312 17680 7332
rect 17701 7312 17705 7332
rect 14736 7295 14771 7296
rect 14051 7154 14614 7182
rect 14715 7288 14771 7295
rect 14715 7268 14744 7288
rect 14764 7268 14771 7288
rect 14715 7263 14771 7268
rect 14944 7292 14994 7300
rect 14944 7271 14960 7292
rect 14982 7271 14994 7292
rect 13645 7098 13972 7132
rect 14052 7126 14086 7154
rect 14051 7123 14087 7126
rect 14051 7104 14059 7123
rect 14079 7104 14087 7123
rect 14051 7100 14087 7104
rect 13662 7097 13972 7098
rect 13937 7068 13972 7097
rect 13723 7061 13758 7062
rect 13702 7054 13758 7061
rect 13702 7034 13731 7054
rect 13751 7034 13758 7054
rect 13702 7029 13758 7034
rect 13932 7056 13974 7068
rect 13932 7036 13941 7056
rect 13965 7036 13974 7056
rect 13702 6823 13736 7029
rect 13932 7028 13974 7036
rect 14149 7057 14181 7064
rect 14149 7037 14155 7057
rect 14176 7037 14181 7057
rect 14149 7009 14181 7037
rect 14715 7057 14749 7263
rect 14944 7262 14994 7271
rect 15162 7291 15194 7298
rect 15162 7271 15168 7291
rect 15189 7271 15194 7291
rect 15162 7243 15194 7271
rect 14782 7235 15194 7243
rect 14782 7209 14788 7235
rect 14814 7209 15194 7235
rect 14782 7207 15194 7209
rect 14784 7206 14824 7207
rect 15162 7142 15194 7207
rect 17673 7247 17705 7312
rect 18043 7247 18083 7248
rect 17673 7245 18085 7247
rect 17673 7219 18053 7245
rect 18079 7219 18085 7245
rect 17673 7211 18085 7219
rect 17058 7191 17090 7192
rect 17055 7186 17090 7191
rect 17055 7166 17062 7186
rect 17082 7166 17090 7186
rect 17055 7158 17090 7166
rect 15162 7122 15166 7142
rect 15187 7122 15194 7142
rect 15162 7115 15194 7122
rect 16611 7093 16643 7100
rect 16611 7073 16618 7093
rect 16639 7073 16643 7093
rect 14715 7049 14750 7057
rect 14715 7029 14723 7049
rect 14743 7029 14750 7049
rect 14715 7024 14750 7029
rect 14715 7023 14747 7024
rect 13769 7001 14181 7009
rect 13769 6975 13775 7001
rect 13801 6975 14181 7001
rect 13769 6973 14181 6975
rect 13771 6972 13811 6973
rect 14149 6908 14181 6973
rect 16611 7008 16643 7073
rect 16981 7008 17021 7009
rect 16611 7006 17023 7008
rect 16611 6980 16991 7006
rect 17017 6980 17023 7006
rect 16611 6972 17023 6980
rect 14149 6888 14153 6908
rect 14174 6888 14181 6908
rect 14149 6881 14181 6888
rect 14626 6919 14978 6950
rect 13702 6815 13737 6823
rect 13702 6795 13710 6815
rect 13730 6795 13737 6815
rect 13702 6779 13737 6795
rect 14626 6779 14657 6919
rect 14950 6887 14978 6919
rect 16611 6944 16643 6972
rect 17056 6952 17090 7158
rect 17673 7183 17705 7211
rect 17673 7163 17678 7183
rect 17699 7163 17705 7183
rect 17673 7156 17705 7163
rect 17884 7182 17922 7194
rect 18118 7191 18152 7395
rect 18928 7365 18962 7569
rect 19375 7549 19407 7577
rect 19990 7602 20024 7808
rect 20437 7788 20469 7816
rect 20057 7780 20469 7788
rect 20057 7754 20063 7780
rect 20089 7754 20469 7780
rect 20057 7752 20469 7754
rect 20059 7751 20099 7752
rect 20437 7687 20469 7752
rect 20437 7667 20441 7687
rect 20462 7667 20469 7687
rect 20437 7660 20469 7667
rect 19990 7594 20025 7602
rect 19990 7574 19998 7594
rect 20018 7574 20025 7594
rect 19990 7569 20025 7574
rect 19990 7568 20022 7569
rect 18995 7541 19407 7549
rect 18995 7515 19001 7541
rect 19027 7515 19407 7541
rect 18995 7513 19407 7515
rect 18997 7512 19037 7513
rect 19375 7448 19407 7513
rect 19375 7428 19379 7448
rect 19400 7428 19407 7448
rect 19375 7421 19407 7428
rect 17884 7165 17893 7182
rect 17917 7165 17922 7182
rect 17884 7122 17922 7165
rect 18096 7186 18152 7191
rect 18096 7166 18103 7186
rect 18123 7166 18152 7186
rect 18096 7159 18152 7166
rect 18926 7355 18966 7365
rect 18926 7335 18936 7355
rect 18956 7335 18966 7355
rect 19861 7341 20270 7342
rect 18096 7158 18131 7159
rect 18230 7122 18314 7127
rect 17884 7093 18314 7122
rect 16611 6924 16616 6944
rect 16637 6924 16643 6944
rect 16611 6917 16643 6924
rect 16820 6946 16860 6951
rect 16820 6925 16832 6946
rect 16854 6925 16860 6946
rect 16820 6913 16860 6925
rect 17034 6947 17090 6952
rect 17034 6927 17041 6947
rect 17061 6927 17090 6947
rect 17034 6920 17090 6927
rect 17147 7021 18104 7040
rect 17034 6919 17069 6920
rect 14735 6880 14770 6881
rect 13700 6760 14657 6779
rect 14714 6873 14770 6880
rect 14714 6853 14743 6873
rect 14763 6853 14770 6873
rect 14714 6848 14770 6853
rect 14944 6875 14984 6887
rect 14944 6854 14950 6875
rect 14972 6854 14984 6875
rect 14944 6849 14984 6854
rect 15161 6876 15193 6883
rect 15161 6856 15167 6876
rect 15188 6856 15193 6876
rect 13410 6662 13447 6667
rect 13410 6656 13757 6662
rect 13410 6637 13418 6656
rect 13441 6637 13757 6656
rect 13410 6632 13757 6637
rect 13410 6626 13447 6632
rect 13727 6601 13757 6632
rect 14714 6642 14748 6848
rect 15161 6828 15193 6856
rect 16826 6881 16854 6913
rect 17147 6881 17178 7021
rect 18067 7005 18102 7021
rect 18067 6985 18074 7005
rect 18094 6985 18102 7005
rect 18067 6977 18102 6985
rect 16826 6850 17178 6881
rect 17623 6912 17655 6919
rect 17623 6892 17630 6912
rect 17651 6892 17655 6912
rect 14781 6820 15193 6828
rect 14781 6794 14787 6820
rect 14813 6794 15193 6820
rect 14781 6792 15193 6794
rect 14783 6791 14823 6792
rect 15161 6727 15193 6792
rect 17623 6827 17655 6892
rect 17993 6827 18033 6828
rect 17623 6825 18035 6827
rect 17623 6799 18003 6825
rect 18029 6799 18035 6825
rect 17623 6791 18035 6799
rect 17057 6776 17089 6777
rect 17054 6771 17089 6776
rect 17054 6751 17061 6771
rect 17081 6751 17089 6771
rect 17054 6743 17089 6751
rect 15161 6707 15165 6727
rect 15186 6707 15193 6727
rect 15161 6700 15193 6707
rect 16610 6678 16642 6685
rect 16610 6658 16617 6678
rect 16638 6658 16642 6678
rect 14714 6634 14749 6642
rect 14714 6614 14722 6634
rect 14742 6614 14749 6634
rect 14714 6609 14749 6614
rect 14714 6608 14746 6609
rect 13515 6594 13550 6595
rect 13494 6587 13550 6594
rect 13494 6567 13523 6587
rect 13543 6567 13550 6587
rect 13494 6562 13550 6567
rect 13725 6588 13764 6601
rect 13725 6569 13730 6588
rect 13753 6569 13764 6588
rect 13725 6563 13764 6569
rect 13941 6590 13973 6597
rect 13941 6570 13947 6590
rect 13968 6570 13973 6590
rect 12998 6514 13036 6520
rect 12998 6494 13008 6514
rect 13028 6494 13036 6514
rect 12998 6492 13036 6494
rect 11534 6459 11949 6488
rect 13001 6486 13036 6492
rect 11534 6458 11943 6459
rect 8561 6392 8565 6412
rect 8586 6392 8593 6412
rect 8561 6385 8593 6392
rect 12557 6421 12589 6428
rect 12557 6401 12564 6421
rect 12585 6401 12589 6421
rect 9207 6354 9616 6355
rect 8114 6321 8149 6327
rect 9201 6325 9616 6354
rect 8114 6319 8152 6321
rect 8114 6299 8122 6319
rect 8142 6299 8152 6319
rect 8114 6293 8152 6299
rect 7381 6222 7391 6248
rect 7416 6222 7428 6248
rect 7381 6220 7428 6222
rect 7600 6246 7656 6251
rect 7600 6226 7607 6246
rect 7627 6226 7656 6246
rect 6404 6204 6436 6205
rect 6401 6199 6436 6204
rect 6401 6179 6408 6199
rect 6428 6179 6436 6199
rect 6401 6171 6436 6179
rect 4508 6135 4512 6155
rect 4533 6135 4540 6155
rect 4508 6128 4540 6135
rect 5957 6106 5989 6113
rect 5957 6086 5964 6106
rect 5985 6086 5989 6106
rect 4061 6062 4096 6070
rect 4061 6042 4069 6062
rect 4089 6042 4096 6062
rect 4061 6037 4096 6042
rect 4061 6036 4093 6037
rect 3115 6014 3527 6022
rect 3115 5988 3121 6014
rect 3147 5988 3527 6014
rect 3115 5986 3527 5988
rect 3117 5985 3157 5986
rect 3495 5921 3527 5986
rect 5957 6021 5989 6086
rect 6327 6021 6367 6022
rect 5957 6019 6369 6021
rect 5957 5993 6337 6019
rect 6363 5993 6369 6019
rect 5957 5985 6369 5993
rect 3495 5901 3499 5921
rect 3520 5901 3527 5921
rect 3495 5894 3527 5901
rect 3972 5932 4324 5963
rect 3048 5828 3083 5836
rect 3048 5808 3056 5828
rect 3076 5808 3083 5828
rect 3048 5792 3083 5808
rect 3972 5792 4003 5932
rect 4296 5900 4324 5932
rect 5957 5957 5989 5985
rect 6402 5965 6436 6171
rect 7386 6185 7423 6220
rect 7600 6219 7656 6226
rect 7600 6218 7635 6219
rect 7720 6185 7752 6187
rect 7386 6152 7756 6185
rect 5957 5937 5962 5957
rect 5983 5937 5989 5957
rect 5957 5930 5989 5937
rect 6166 5959 6206 5964
rect 6166 5938 6178 5959
rect 6200 5938 6206 5959
rect 6166 5926 6206 5938
rect 6380 5960 6436 5965
rect 6380 5940 6387 5960
rect 6407 5940 6436 5960
rect 6380 5933 6436 5940
rect 6493 6034 7450 6053
rect 6380 5932 6415 5933
rect 4081 5893 4116 5894
rect 3046 5773 4003 5792
rect 4060 5886 4116 5893
rect 4060 5866 4089 5886
rect 4109 5866 4116 5886
rect 4060 5861 4116 5866
rect 4290 5888 4330 5900
rect 4290 5867 4296 5888
rect 4318 5867 4330 5888
rect 4290 5862 4330 5867
rect 4507 5889 4539 5896
rect 4507 5869 4513 5889
rect 4534 5869 4539 5889
rect 2836 5691 3266 5720
rect 2836 5686 2920 5691
rect 3019 5654 3054 5655
rect 2998 5647 3054 5654
rect 2998 5627 3027 5647
rect 3047 5627 3054 5647
rect 2998 5622 3054 5627
rect 3228 5648 3266 5691
rect 3228 5631 3233 5648
rect 3257 5631 3266 5648
rect 2998 5418 3032 5622
rect 3228 5619 3266 5631
rect 3445 5650 3477 5657
rect 3445 5630 3451 5650
rect 3472 5630 3477 5650
rect 3445 5602 3477 5630
rect 4060 5655 4094 5861
rect 4507 5841 4539 5869
rect 6172 5894 6200 5926
rect 6493 5894 6524 6034
rect 7413 6018 7448 6034
rect 7413 5998 7420 6018
rect 7440 5998 7448 6018
rect 7413 5990 7448 5998
rect 6172 5863 6524 5894
rect 6969 5925 7001 5932
rect 6969 5905 6976 5925
rect 6997 5905 7001 5925
rect 4127 5833 4539 5841
rect 4127 5807 4133 5833
rect 4159 5807 4539 5833
rect 4127 5805 4539 5807
rect 4129 5804 4169 5805
rect 4507 5740 4539 5805
rect 6969 5840 7001 5905
rect 7339 5840 7379 5841
rect 6969 5838 7381 5840
rect 6969 5812 7349 5838
rect 7375 5812 7381 5838
rect 6969 5804 7381 5812
rect 6403 5789 6435 5790
rect 6400 5784 6435 5789
rect 6400 5764 6407 5784
rect 6427 5764 6435 5784
rect 6400 5756 6435 5764
rect 4507 5720 4511 5740
rect 4532 5720 4539 5740
rect 4507 5713 4539 5720
rect 5956 5691 5988 5698
rect 5956 5671 5963 5691
rect 5984 5671 5988 5691
rect 4060 5647 4095 5655
rect 4060 5627 4068 5647
rect 4088 5627 4095 5647
rect 4060 5622 4095 5627
rect 4060 5621 4092 5622
rect 3065 5594 3477 5602
rect 3065 5568 3071 5594
rect 3097 5568 3477 5594
rect 3065 5566 3477 5568
rect 3067 5565 3107 5566
rect 3445 5501 3477 5566
rect 5956 5606 5988 5671
rect 6326 5606 6366 5607
rect 5956 5604 6368 5606
rect 5956 5578 6336 5604
rect 6362 5578 6368 5604
rect 5956 5570 6368 5578
rect 5956 5542 5988 5570
rect 5956 5522 5961 5542
rect 5982 5522 5988 5542
rect 5956 5515 5988 5522
rect 6156 5542 6206 5551
rect 6401 5550 6435 5756
rect 6969 5776 7001 5804
rect 6969 5756 6974 5776
rect 6995 5756 7001 5776
rect 6969 5749 7001 5756
rect 7176 5777 7218 5785
rect 7414 5784 7448 5990
rect 7176 5757 7185 5777
rect 7209 5757 7218 5777
rect 7176 5745 7218 5757
rect 7392 5779 7448 5784
rect 7392 5759 7399 5779
rect 7419 5759 7448 5779
rect 7392 5752 7448 5759
rect 7392 5751 7427 5752
rect 7178 5716 7213 5745
rect 7178 5715 7488 5716
rect 7063 5709 7099 5713
rect 7063 5690 7071 5709
rect 7091 5690 7099 5709
rect 7063 5687 7099 5690
rect 7064 5659 7098 5687
rect 7178 5681 7505 5715
rect 6156 5521 6168 5542
rect 6190 5521 6206 5542
rect 6156 5513 6206 5521
rect 6379 5545 6435 5550
rect 6379 5525 6386 5545
rect 6406 5525 6435 5545
rect 6379 5518 6435 5525
rect 6536 5631 7099 5659
rect 6379 5517 6414 5518
rect 3445 5481 3449 5501
rect 3470 5481 3477 5501
rect 3445 5474 3477 5481
rect 6161 5480 6202 5513
rect 6536 5480 6576 5631
rect 6161 5451 6576 5480
rect 7465 5457 7505 5681
rect 6161 5450 6570 5451
rect 7465 5437 7475 5457
rect 7495 5437 7505 5457
rect 7465 5427 7505 5437
rect 2996 5408 3036 5418
rect 2996 5388 3006 5408
rect 3026 5388 3036 5408
rect 3931 5394 4340 5395
rect 2996 5164 3036 5388
rect 3925 5365 4340 5394
rect 3925 5214 3965 5365
rect 4299 5332 4340 5365
rect 7024 5364 7056 5371
rect 7024 5344 7031 5364
rect 7052 5344 7056 5364
rect 4087 5327 4122 5328
rect 3402 5186 3965 5214
rect 4066 5320 4122 5327
rect 4066 5300 4095 5320
rect 4115 5300 4122 5320
rect 4066 5295 4122 5300
rect 4295 5324 4345 5332
rect 4295 5303 4311 5324
rect 4333 5303 4345 5324
rect 2996 5130 3323 5164
rect 3403 5158 3437 5186
rect 3402 5155 3438 5158
rect 3402 5136 3410 5155
rect 3430 5136 3438 5155
rect 3402 5132 3438 5136
rect 3013 5129 3323 5130
rect 3288 5100 3323 5129
rect 3074 5093 3109 5094
rect 3053 5086 3109 5093
rect 3053 5066 3082 5086
rect 3102 5066 3109 5086
rect 3053 5061 3109 5066
rect 3283 5088 3325 5100
rect 3283 5068 3292 5088
rect 3316 5068 3325 5088
rect 3053 4855 3087 5061
rect 3283 5060 3325 5068
rect 3500 5089 3532 5096
rect 3500 5069 3506 5089
rect 3527 5069 3532 5089
rect 3500 5041 3532 5069
rect 4066 5089 4100 5295
rect 4295 5294 4345 5303
rect 4513 5323 4545 5330
rect 4513 5303 4519 5323
rect 4540 5303 4545 5323
rect 4513 5275 4545 5303
rect 4133 5267 4545 5275
rect 4133 5241 4139 5267
rect 4165 5241 4545 5267
rect 4133 5239 4545 5241
rect 4135 5238 4175 5239
rect 4513 5174 4545 5239
rect 7024 5279 7056 5344
rect 7394 5279 7434 5280
rect 7024 5277 7436 5279
rect 7024 5251 7404 5277
rect 7430 5251 7436 5277
rect 7024 5243 7436 5251
rect 6409 5223 6441 5224
rect 6406 5218 6441 5223
rect 6406 5198 6413 5218
rect 6433 5198 6441 5218
rect 6406 5190 6441 5198
rect 4513 5154 4517 5174
rect 4538 5154 4545 5174
rect 4513 5147 4545 5154
rect 5962 5125 5994 5132
rect 5962 5105 5969 5125
rect 5990 5105 5994 5125
rect 4066 5081 4101 5089
rect 4066 5061 4074 5081
rect 4094 5061 4101 5081
rect 4066 5056 4101 5061
rect 4066 5055 4098 5056
rect 3120 5033 3532 5041
rect 3120 5007 3126 5033
rect 3152 5007 3532 5033
rect 3120 5005 3532 5007
rect 3122 5004 3162 5005
rect 3500 4940 3532 5005
rect 5962 5040 5994 5105
rect 6332 5040 6372 5041
rect 5962 5038 6374 5040
rect 5962 5012 6342 5038
rect 6368 5012 6374 5038
rect 5962 5004 6374 5012
rect 3500 4920 3504 4940
rect 3525 4920 3532 4940
rect 3500 4913 3532 4920
rect 3977 4951 4329 4982
rect 3053 4847 3088 4855
rect 3053 4827 3061 4847
rect 3081 4827 3088 4847
rect 3053 4811 3088 4827
rect 3977 4811 4008 4951
rect 4301 4919 4329 4951
rect 5962 4976 5994 5004
rect 6407 4984 6441 5190
rect 7024 5215 7056 5243
rect 7469 5223 7503 5427
rect 7024 5195 7029 5215
rect 7050 5195 7056 5215
rect 7024 5188 7056 5195
rect 7235 5215 7272 5221
rect 7235 5196 7241 5215
rect 7264 5196 7272 5215
rect 7235 5191 7272 5196
rect 7447 5218 7503 5223
rect 7447 5198 7454 5218
rect 7474 5198 7503 5218
rect 7447 5191 7503 5198
rect 7243 5154 7267 5191
rect 7447 5190 7482 5191
rect 7243 5152 7611 5154
rect 7243 5147 7616 5152
rect 7243 5129 7589 5147
rect 7609 5129 7616 5147
rect 7243 5124 7616 5129
rect 7587 5122 7616 5124
rect 5962 4956 5967 4976
rect 5988 4956 5994 4976
rect 5962 4949 5994 4956
rect 6171 4978 6211 4983
rect 6171 4957 6183 4978
rect 6205 4957 6211 4978
rect 6171 4945 6211 4957
rect 6385 4979 6441 4984
rect 6385 4959 6392 4979
rect 6412 4959 6441 4979
rect 6385 4952 6441 4959
rect 6498 5053 7455 5072
rect 6385 4951 6420 4952
rect 4086 4912 4121 4913
rect 3051 4792 4008 4811
rect 4065 4905 4121 4912
rect 4065 4885 4094 4905
rect 4114 4885 4121 4905
rect 4065 4880 4121 4885
rect 4295 4907 4335 4919
rect 4295 4886 4301 4907
rect 4323 4886 4335 4907
rect 4295 4881 4335 4886
rect 4512 4908 4544 4915
rect 4512 4888 4518 4908
rect 4539 4888 4544 4908
rect 2649 4735 2734 4738
rect 2642 4731 2734 4735
rect 2642 4730 3023 4731
rect 2642 4700 2649 4730
rect 2686 4701 3023 4730
rect 2686 4700 2734 4701
rect 2642 4698 2734 4700
rect 2642 4695 2727 4698
rect 2988 4663 3023 4701
rect 4065 4674 4099 4880
rect 4512 4860 4544 4888
rect 6177 4913 6205 4945
rect 6498 4913 6529 5053
rect 7418 5037 7453 5053
rect 7418 5017 7425 5037
rect 7445 5017 7453 5037
rect 7418 5009 7453 5017
rect 6177 4882 6529 4913
rect 6974 4944 7006 4951
rect 6974 4924 6981 4944
rect 7002 4924 7006 4944
rect 4132 4852 4544 4860
rect 4132 4826 4138 4852
rect 4164 4826 4544 4852
rect 4132 4824 4544 4826
rect 4134 4823 4174 4824
rect 4512 4759 4544 4824
rect 6974 4859 7006 4924
rect 7344 4859 7384 4860
rect 6974 4857 7386 4859
rect 6974 4831 7354 4857
rect 7380 4831 7386 4857
rect 6974 4823 7386 4831
rect 6408 4808 6440 4809
rect 6405 4803 6440 4808
rect 6405 4783 6412 4803
rect 6432 4783 6440 4803
rect 6405 4775 6440 4783
rect 4512 4739 4516 4759
rect 4537 4739 4544 4759
rect 4512 4732 4544 4739
rect 5961 4710 5993 4717
rect 5961 4690 5968 4710
rect 5989 4690 5993 4710
rect 4065 4666 4100 4674
rect 2779 4661 2814 4662
rect 885 4491 1300 4520
rect 2438 4519 2471 4520
rect 2435 4514 2471 4519
rect 2435 4494 2442 4514
rect 2462 4494 2471 4514
rect 885 4490 1294 4491
rect 2435 4489 2471 4494
rect 2758 4654 2814 4661
rect 2758 4634 2787 4654
rect 2807 4634 2814 4654
rect 2758 4629 2814 4634
rect 2983 4654 3032 4663
rect 2983 4635 2991 4654
rect 3017 4635 3032 4654
rect 2435 4486 2470 4489
rect 1991 4421 2023 4428
rect 1991 4401 1998 4421
rect 2019 4401 2023 4421
rect 1991 4336 2023 4401
rect 2361 4336 2401 4337
rect 1991 4334 2403 4336
rect 1991 4308 2371 4334
rect 2397 4308 2403 4334
rect 1991 4300 2403 4308
rect 1991 4272 2023 4300
rect 1131 4268 1163 4269
rect 1128 4263 1163 4268
rect 1128 4243 1135 4263
rect 1155 4243 1163 4263
rect 1991 4252 1996 4272
rect 2017 4252 2023 4272
rect 1991 4245 2023 4252
rect 2196 4274 2245 4284
rect 2436 4280 2470 4486
rect 2758 4423 2792 4629
rect 2983 4625 3032 4635
rect 3205 4657 3237 4664
rect 3205 4637 3211 4657
rect 3232 4637 3237 4657
rect 4065 4646 4073 4666
rect 4093 4646 4100 4666
rect 4065 4641 4100 4646
rect 4065 4640 4097 4641
rect 3205 4609 3237 4637
rect 2825 4601 3237 4609
rect 2825 4575 2831 4601
rect 2857 4575 3237 4601
rect 2825 4573 3237 4575
rect 2827 4572 2867 4573
rect 3205 4508 3237 4573
rect 5961 4625 5993 4690
rect 6331 4625 6371 4626
rect 5961 4623 6373 4625
rect 5961 4597 6341 4623
rect 6367 4597 6373 4623
rect 5961 4589 6373 4597
rect 5961 4561 5993 4589
rect 5961 4541 5966 4561
rect 5987 4541 5993 4561
rect 5961 4534 5993 4541
rect 6161 4561 6211 4570
rect 6406 4569 6440 4775
rect 6974 4795 7006 4823
rect 6974 4775 6979 4795
rect 7000 4775 7006 4795
rect 7179 4797 7221 4806
rect 7419 4803 7453 5009
rect 7179 4783 7189 4797
rect 6974 4768 7006 4775
rect 7178 4777 7189 4783
rect 7213 4777 7221 4797
rect 7178 4766 7221 4777
rect 7397 4798 7453 4803
rect 7397 4778 7404 4798
rect 7424 4778 7453 4798
rect 7397 4771 7453 4778
rect 7397 4770 7432 4771
rect 7178 4736 7218 4766
rect 7068 4728 7104 4732
rect 7068 4709 7076 4728
rect 7096 4709 7104 4728
rect 7068 4706 7104 4709
rect 7178 4731 7525 4736
rect 7069 4678 7103 4706
rect 7178 4705 7497 4731
rect 7516 4705 7525 4731
rect 7178 4701 7525 4705
rect 6161 4540 6173 4561
rect 6195 4540 6211 4561
rect 6161 4532 6211 4540
rect 6384 4564 6440 4569
rect 6384 4544 6391 4564
rect 6411 4544 6440 4564
rect 6384 4537 6440 4544
rect 6541 4650 7104 4678
rect 6384 4536 6419 4537
rect 3205 4488 3209 4508
rect 3230 4488 3237 4508
rect 3205 4481 3237 4488
rect 6166 4499 6207 4532
rect 6541 4499 6581 4650
rect 7720 4499 7752 6152
rect 8117 5699 8152 6293
rect 9201 6174 9241 6325
rect 9575 6292 9616 6325
rect 12557 6336 12589 6401
rect 12927 6336 12967 6337
rect 12557 6334 12969 6336
rect 12557 6308 12937 6334
rect 12963 6308 12969 6334
rect 12557 6300 12969 6308
rect 9363 6287 9398 6288
rect 8678 6146 9241 6174
rect 9342 6280 9398 6287
rect 9342 6260 9371 6280
rect 9391 6260 9398 6280
rect 9342 6255 9398 6260
rect 9571 6284 9621 6292
rect 9571 6263 9587 6284
rect 9609 6263 9621 6284
rect 8257 6119 8604 6123
rect 8257 6093 8266 6119
rect 8285 6093 8604 6119
rect 8679 6118 8713 6146
rect 8257 6088 8604 6093
rect 8678 6115 8714 6118
rect 8678 6096 8686 6115
rect 8706 6096 8714 6115
rect 8678 6092 8714 6096
rect 8564 6058 8604 6088
rect 8350 6053 8385 6054
rect 8329 6046 8385 6053
rect 8329 6026 8358 6046
rect 8378 6026 8385 6046
rect 8329 6021 8385 6026
rect 8561 6047 8604 6058
rect 8561 6027 8569 6047
rect 8593 6041 8604 6047
rect 8776 6049 8808 6056
rect 8593 6027 8603 6041
rect 8329 5815 8363 6021
rect 8561 6018 8603 6027
rect 8776 6029 8782 6049
rect 8803 6029 8808 6049
rect 8776 6001 8808 6029
rect 9342 6049 9376 6255
rect 9571 6254 9621 6263
rect 9789 6283 9821 6290
rect 9789 6263 9795 6283
rect 9816 6263 9821 6283
rect 9789 6235 9821 6263
rect 12557 6272 12589 6300
rect 12557 6252 12562 6272
rect 12583 6252 12589 6272
rect 12557 6245 12589 6252
rect 12761 6277 12808 6283
rect 13002 6280 13036 6486
rect 13494 6356 13528 6562
rect 13941 6542 13973 6570
rect 13561 6534 13973 6542
rect 13561 6508 13567 6534
rect 13593 6508 13973 6534
rect 13561 6506 13973 6508
rect 13563 6505 13603 6506
rect 13941 6441 13973 6506
rect 16610 6593 16642 6658
rect 16980 6593 17020 6594
rect 16610 6591 17022 6593
rect 16610 6565 16990 6591
rect 17016 6565 17022 6591
rect 16610 6557 17022 6565
rect 16610 6529 16642 6557
rect 16610 6509 16615 6529
rect 16636 6509 16642 6529
rect 16610 6502 16642 6509
rect 16810 6529 16860 6538
rect 17055 6537 17089 6743
rect 17623 6763 17655 6791
rect 17623 6743 17628 6763
rect 17649 6743 17655 6763
rect 17828 6765 17870 6774
rect 18068 6771 18102 6977
rect 17828 6751 17838 6765
rect 17623 6736 17655 6743
rect 17827 6745 17838 6751
rect 17862 6745 17870 6765
rect 17827 6734 17870 6745
rect 18046 6766 18102 6771
rect 18046 6746 18053 6766
rect 18073 6746 18102 6766
rect 18046 6739 18102 6746
rect 18046 6738 18081 6739
rect 17827 6704 17867 6734
rect 17717 6696 17753 6700
rect 17717 6677 17725 6696
rect 17745 6677 17753 6696
rect 17717 6674 17753 6677
rect 17827 6699 18174 6704
rect 17718 6646 17752 6674
rect 17827 6673 18146 6699
rect 18165 6673 18174 6699
rect 17827 6669 18174 6673
rect 16810 6508 16822 6529
rect 16844 6508 16860 6529
rect 16810 6500 16860 6508
rect 17033 6532 17089 6537
rect 17033 6512 17040 6532
rect 17060 6512 17089 6532
rect 17033 6505 17089 6512
rect 17190 6618 17753 6646
rect 17033 6504 17068 6505
rect 13941 6421 13945 6441
rect 13966 6421 13973 6441
rect 16815 6467 16856 6500
rect 17190 6467 17230 6618
rect 18279 6499 18314 7093
rect 18926 7111 18966 7335
rect 19855 7312 20270 7341
rect 19855 7161 19895 7312
rect 20229 7279 20270 7312
rect 20017 7274 20052 7275
rect 19332 7133 19895 7161
rect 19996 7267 20052 7274
rect 19996 7247 20025 7267
rect 20045 7247 20052 7267
rect 19996 7242 20052 7247
rect 20225 7271 20275 7279
rect 20225 7250 20241 7271
rect 20263 7250 20275 7271
rect 18926 7077 19253 7111
rect 19333 7105 19367 7133
rect 19332 7102 19368 7105
rect 19332 7083 19340 7102
rect 19360 7083 19368 7102
rect 19332 7079 19368 7083
rect 18943 7076 19253 7077
rect 19218 7047 19253 7076
rect 19004 7040 19039 7041
rect 18983 7033 19039 7040
rect 18983 7013 19012 7033
rect 19032 7013 19039 7033
rect 18983 7008 19039 7013
rect 19213 7035 19255 7047
rect 19213 7015 19222 7035
rect 19246 7015 19255 7035
rect 18983 6802 19017 7008
rect 19213 7007 19255 7015
rect 19430 7036 19462 7043
rect 19430 7016 19436 7036
rect 19457 7016 19462 7036
rect 19430 6988 19462 7016
rect 19996 7036 20030 7242
rect 20225 7241 20275 7250
rect 20443 7270 20475 7277
rect 20443 7250 20449 7270
rect 20470 7250 20475 7270
rect 20443 7222 20475 7250
rect 20063 7214 20475 7222
rect 20063 7188 20069 7214
rect 20095 7188 20475 7214
rect 20063 7186 20475 7188
rect 20065 7185 20105 7186
rect 20443 7121 20475 7186
rect 20443 7101 20447 7121
rect 20468 7101 20475 7121
rect 20443 7094 20475 7101
rect 19996 7028 20031 7036
rect 19996 7008 20004 7028
rect 20024 7008 20031 7028
rect 19996 7003 20031 7008
rect 19996 7002 20028 7003
rect 19050 6980 19462 6988
rect 19050 6954 19056 6980
rect 19082 6954 19462 6980
rect 19050 6952 19462 6954
rect 19052 6951 19092 6952
rect 19430 6887 19462 6952
rect 19430 6867 19434 6887
rect 19455 6867 19462 6887
rect 19430 6860 19462 6867
rect 19907 6898 20259 6929
rect 18983 6794 19018 6802
rect 18983 6774 18991 6794
rect 19011 6774 19018 6794
rect 18983 6758 19018 6774
rect 19907 6758 19938 6898
rect 20231 6866 20259 6898
rect 20016 6859 20051 6860
rect 18981 6739 19938 6758
rect 19995 6852 20051 6859
rect 19995 6832 20024 6852
rect 20044 6832 20051 6852
rect 19995 6827 20051 6832
rect 20225 6854 20265 6866
rect 20225 6833 20231 6854
rect 20253 6833 20265 6854
rect 20225 6828 20265 6833
rect 20442 6855 20474 6862
rect 20442 6835 20448 6855
rect 20469 6835 20474 6855
rect 18691 6641 18728 6646
rect 18691 6635 19038 6641
rect 18691 6616 18699 6635
rect 18722 6616 19038 6635
rect 18691 6611 19038 6616
rect 18691 6605 18728 6611
rect 19008 6580 19038 6611
rect 19995 6621 20029 6827
rect 20442 6807 20474 6835
rect 20062 6799 20474 6807
rect 20062 6773 20068 6799
rect 20094 6773 20474 6799
rect 20062 6771 20474 6773
rect 20064 6770 20104 6771
rect 20442 6706 20474 6771
rect 20442 6686 20446 6706
rect 20467 6686 20474 6706
rect 20442 6679 20474 6686
rect 19995 6613 20030 6621
rect 19995 6593 20003 6613
rect 20023 6593 20030 6613
rect 19995 6588 20030 6593
rect 19995 6587 20027 6588
rect 18796 6573 18831 6574
rect 18775 6566 18831 6573
rect 18775 6546 18804 6566
rect 18824 6546 18831 6566
rect 18775 6541 18831 6546
rect 19006 6567 19045 6580
rect 19006 6548 19011 6567
rect 19034 6548 19045 6567
rect 19006 6542 19045 6548
rect 19222 6569 19254 6576
rect 19222 6549 19228 6569
rect 19249 6549 19254 6569
rect 18279 6493 18317 6499
rect 18279 6473 18289 6493
rect 18309 6473 18317 6493
rect 18279 6471 18317 6473
rect 16815 6438 17230 6467
rect 18282 6465 18317 6471
rect 16815 6437 17224 6438
rect 13941 6414 13973 6421
rect 17838 6400 17870 6407
rect 14587 6383 14996 6384
rect 13494 6350 13529 6356
rect 14581 6354 14996 6383
rect 13494 6348 13532 6350
rect 13494 6328 13502 6348
rect 13522 6328 13532 6348
rect 13494 6322 13532 6328
rect 12761 6251 12771 6277
rect 12796 6251 12808 6277
rect 12761 6249 12808 6251
rect 12980 6275 13036 6280
rect 12980 6255 12987 6275
rect 13007 6255 13036 6275
rect 9409 6227 9821 6235
rect 11784 6233 11816 6234
rect 9409 6201 9415 6227
rect 9441 6201 9821 6227
rect 9409 6199 9821 6201
rect 11781 6228 11816 6233
rect 11781 6208 11788 6228
rect 11808 6208 11816 6228
rect 11781 6200 11816 6208
rect 9411 6198 9451 6199
rect 9789 6134 9821 6199
rect 9789 6114 9793 6134
rect 9814 6114 9821 6134
rect 9789 6107 9821 6114
rect 11337 6135 11369 6142
rect 11337 6115 11344 6135
rect 11365 6115 11369 6135
rect 11337 6050 11369 6115
rect 11707 6050 11747 6051
rect 9342 6041 9377 6049
rect 9342 6021 9350 6041
rect 9370 6021 9377 6041
rect 9342 6016 9377 6021
rect 11337 6048 11749 6050
rect 11337 6022 11717 6048
rect 11743 6022 11749 6048
rect 9342 6015 9374 6016
rect 8396 5993 8808 6001
rect 8396 5967 8402 5993
rect 8428 5967 8808 5993
rect 8396 5965 8808 5967
rect 8398 5964 8438 5965
rect 8776 5900 8808 5965
rect 11337 6014 11749 6022
rect 11337 5986 11369 6014
rect 11782 5994 11816 6200
rect 12766 6214 12803 6249
rect 12980 6248 13036 6255
rect 12980 6247 13015 6248
rect 13100 6214 13132 6216
rect 12766 6181 13136 6214
rect 11337 5966 11342 5986
rect 11363 5966 11369 5986
rect 11337 5959 11369 5966
rect 11546 5988 11586 5993
rect 11546 5967 11558 5988
rect 11580 5967 11586 5988
rect 11546 5955 11586 5967
rect 11760 5989 11816 5994
rect 11760 5969 11767 5989
rect 11787 5969 11816 5989
rect 11760 5962 11816 5969
rect 11873 6063 12830 6082
rect 11760 5961 11795 5962
rect 8776 5880 8780 5900
rect 8801 5880 8808 5900
rect 8776 5873 8808 5880
rect 9253 5911 9605 5942
rect 8329 5807 8364 5815
rect 8329 5787 8337 5807
rect 8357 5787 8364 5807
rect 8329 5771 8364 5787
rect 9253 5771 9284 5911
rect 9577 5879 9605 5911
rect 11552 5923 11580 5955
rect 11873 5923 11904 6063
rect 12793 6047 12828 6063
rect 12793 6027 12800 6047
rect 12820 6027 12828 6047
rect 12793 6019 12828 6027
rect 11552 5892 11904 5923
rect 12349 5954 12381 5961
rect 12349 5934 12356 5954
rect 12377 5934 12381 5954
rect 9362 5872 9397 5873
rect 8327 5752 9284 5771
rect 9341 5865 9397 5872
rect 9341 5845 9370 5865
rect 9390 5845 9397 5865
rect 9341 5840 9397 5845
rect 9571 5867 9611 5879
rect 9571 5846 9577 5867
rect 9599 5846 9611 5867
rect 9571 5841 9611 5846
rect 9788 5868 9820 5875
rect 9788 5848 9794 5868
rect 9815 5848 9820 5868
rect 8117 5670 8547 5699
rect 8117 5665 8201 5670
rect 8300 5633 8335 5634
rect 8279 5626 8335 5633
rect 8279 5606 8308 5626
rect 8328 5606 8335 5626
rect 8279 5601 8335 5606
rect 8509 5627 8547 5670
rect 8509 5610 8514 5627
rect 8538 5610 8547 5627
rect 8279 5397 8313 5601
rect 8509 5598 8547 5610
rect 8726 5629 8758 5636
rect 8726 5609 8732 5629
rect 8753 5609 8758 5629
rect 8726 5581 8758 5609
rect 9341 5634 9375 5840
rect 9788 5820 9820 5848
rect 9408 5812 9820 5820
rect 12349 5869 12381 5934
rect 12719 5869 12759 5870
rect 12349 5867 12761 5869
rect 12349 5841 12729 5867
rect 12755 5841 12761 5867
rect 12349 5833 12761 5841
rect 11783 5818 11815 5819
rect 9408 5786 9414 5812
rect 9440 5786 9820 5812
rect 9408 5784 9820 5786
rect 11780 5813 11815 5818
rect 11780 5793 11787 5813
rect 11807 5793 11815 5813
rect 11780 5785 11815 5793
rect 9410 5783 9450 5784
rect 9788 5719 9820 5784
rect 9788 5699 9792 5719
rect 9813 5699 9820 5719
rect 9788 5692 9820 5699
rect 11336 5720 11368 5727
rect 11336 5700 11343 5720
rect 11364 5700 11368 5720
rect 11336 5635 11368 5700
rect 11706 5635 11746 5636
rect 9341 5626 9376 5634
rect 9341 5606 9349 5626
rect 9369 5606 9376 5626
rect 9341 5601 9376 5606
rect 11336 5633 11748 5635
rect 11336 5607 11716 5633
rect 11742 5607 11748 5633
rect 9341 5600 9373 5601
rect 8346 5573 8758 5581
rect 8346 5547 8352 5573
rect 8378 5547 8758 5573
rect 8346 5545 8758 5547
rect 8348 5544 8388 5545
rect 8726 5480 8758 5545
rect 11336 5599 11748 5607
rect 11336 5571 11368 5599
rect 11336 5551 11341 5571
rect 11362 5551 11368 5571
rect 11336 5544 11368 5551
rect 11536 5571 11586 5580
rect 11781 5579 11815 5785
rect 12349 5805 12381 5833
rect 12349 5785 12354 5805
rect 12375 5785 12381 5805
rect 12349 5778 12381 5785
rect 12556 5806 12598 5814
rect 12794 5813 12828 6019
rect 12556 5786 12565 5806
rect 12589 5786 12598 5806
rect 12556 5774 12598 5786
rect 12772 5808 12828 5813
rect 12772 5788 12779 5808
rect 12799 5788 12828 5808
rect 12772 5781 12828 5788
rect 12772 5780 12807 5781
rect 12558 5745 12593 5774
rect 12558 5744 12868 5745
rect 12443 5738 12479 5742
rect 12443 5719 12451 5738
rect 12471 5719 12479 5738
rect 12443 5716 12479 5719
rect 12444 5688 12478 5716
rect 12558 5710 12885 5744
rect 11536 5550 11548 5571
rect 11570 5550 11586 5571
rect 11536 5542 11586 5550
rect 11759 5574 11815 5579
rect 11759 5554 11766 5574
rect 11786 5554 11815 5574
rect 11759 5547 11815 5554
rect 11916 5660 12479 5688
rect 11759 5546 11794 5547
rect 8726 5460 8730 5480
rect 8751 5460 8758 5480
rect 11541 5509 11582 5542
rect 11916 5509 11956 5660
rect 11541 5480 11956 5509
rect 12845 5486 12885 5710
rect 11541 5479 11950 5480
rect 8726 5453 8758 5460
rect 12845 5466 12855 5486
rect 12875 5466 12885 5486
rect 12845 5456 12885 5466
rect 8277 5387 8317 5397
rect 8277 5367 8287 5387
rect 8307 5367 8317 5387
rect 12404 5393 12436 5400
rect 9212 5373 9621 5374
rect 8277 5143 8317 5367
rect 9206 5344 9621 5373
rect 9206 5193 9246 5344
rect 9580 5311 9621 5344
rect 12404 5373 12411 5393
rect 12432 5373 12436 5393
rect 9368 5306 9403 5307
rect 8683 5165 9246 5193
rect 9347 5299 9403 5306
rect 9347 5279 9376 5299
rect 9396 5279 9403 5299
rect 9347 5274 9403 5279
rect 9576 5303 9626 5311
rect 9576 5282 9592 5303
rect 9614 5282 9626 5303
rect 8277 5109 8604 5143
rect 8684 5137 8718 5165
rect 8683 5134 8719 5137
rect 8683 5115 8691 5134
rect 8711 5115 8719 5134
rect 8683 5111 8719 5115
rect 8294 5108 8604 5109
rect 8569 5079 8604 5108
rect 8355 5072 8390 5073
rect 8334 5065 8390 5072
rect 8334 5045 8363 5065
rect 8383 5045 8390 5065
rect 8334 5040 8390 5045
rect 8564 5067 8606 5079
rect 8564 5047 8573 5067
rect 8597 5047 8606 5067
rect 8334 4834 8368 5040
rect 8564 5039 8606 5047
rect 8781 5068 8813 5075
rect 8781 5048 8787 5068
rect 8808 5048 8813 5068
rect 8781 5020 8813 5048
rect 9347 5068 9381 5274
rect 9576 5273 9626 5282
rect 9794 5302 9826 5309
rect 9794 5282 9800 5302
rect 9821 5282 9826 5302
rect 9794 5254 9826 5282
rect 9414 5246 9826 5254
rect 12404 5308 12436 5373
rect 12774 5308 12814 5309
rect 12404 5306 12816 5308
rect 12404 5280 12784 5306
rect 12810 5280 12816 5306
rect 12404 5272 12816 5280
rect 11789 5252 11821 5253
rect 9414 5220 9420 5246
rect 9446 5220 9826 5246
rect 9414 5218 9826 5220
rect 11786 5247 11821 5252
rect 11786 5227 11793 5247
rect 11813 5227 11821 5247
rect 11786 5219 11821 5227
rect 9416 5217 9456 5218
rect 9794 5153 9826 5218
rect 9794 5133 9798 5153
rect 9819 5133 9826 5153
rect 9794 5126 9826 5133
rect 11342 5154 11374 5161
rect 11342 5134 11349 5154
rect 11370 5134 11374 5154
rect 11342 5069 11374 5134
rect 11712 5069 11752 5070
rect 9347 5060 9382 5068
rect 9347 5040 9355 5060
rect 9375 5040 9382 5060
rect 9347 5035 9382 5040
rect 11342 5067 11754 5069
rect 11342 5041 11722 5067
rect 11748 5041 11754 5067
rect 9347 5034 9379 5035
rect 8401 5012 8813 5020
rect 8401 4986 8407 5012
rect 8433 4986 8813 5012
rect 8401 4984 8813 4986
rect 8403 4983 8443 4984
rect 8781 4919 8813 4984
rect 11342 5033 11754 5041
rect 11342 5005 11374 5033
rect 11787 5013 11821 5219
rect 12404 5244 12436 5272
rect 12849 5252 12883 5456
rect 12404 5224 12409 5244
rect 12430 5224 12436 5244
rect 12404 5217 12436 5224
rect 12615 5244 12652 5250
rect 12615 5225 12621 5244
rect 12644 5225 12652 5244
rect 12615 5220 12652 5225
rect 12827 5247 12883 5252
rect 12827 5227 12834 5247
rect 12854 5227 12883 5247
rect 12827 5220 12883 5227
rect 12623 5183 12647 5220
rect 12827 5219 12862 5220
rect 12623 5181 12991 5183
rect 12623 5176 12996 5181
rect 12623 5158 12969 5176
rect 12989 5158 12996 5176
rect 12623 5153 12996 5158
rect 12967 5151 12996 5153
rect 11342 4985 11347 5005
rect 11368 4985 11374 5005
rect 11342 4978 11374 4985
rect 11551 5007 11591 5012
rect 11551 4986 11563 5007
rect 11585 4986 11591 5007
rect 11551 4974 11591 4986
rect 11765 5008 11821 5013
rect 11765 4988 11772 5008
rect 11792 4988 11821 5008
rect 11765 4981 11821 4988
rect 11878 5082 12835 5101
rect 11765 4980 11800 4981
rect 8781 4899 8785 4919
rect 8806 4899 8813 4919
rect 8781 4892 8813 4899
rect 9258 4930 9610 4961
rect 8334 4826 8369 4834
rect 8334 4806 8342 4826
rect 8362 4806 8369 4826
rect 8334 4790 8369 4806
rect 9258 4790 9289 4930
rect 9582 4898 9610 4930
rect 11557 4942 11585 4974
rect 11878 4942 11909 5082
rect 12798 5066 12833 5082
rect 12798 5046 12805 5066
rect 12825 5046 12833 5066
rect 12798 5038 12833 5046
rect 11557 4911 11909 4942
rect 12354 4973 12386 4980
rect 12354 4953 12361 4973
rect 12382 4953 12386 4973
rect 9367 4891 9402 4892
rect 8332 4771 9289 4790
rect 9346 4884 9402 4891
rect 9346 4864 9375 4884
rect 9395 4864 9402 4884
rect 9346 4859 9402 4864
rect 9576 4886 9616 4898
rect 9576 4865 9582 4886
rect 9604 4865 9616 4886
rect 9576 4860 9616 4865
rect 9793 4887 9825 4894
rect 9793 4867 9799 4887
rect 9820 4867 9825 4887
rect 7930 4714 8015 4717
rect 7923 4710 8015 4714
rect 7923 4709 8304 4710
rect 7923 4679 7930 4709
rect 7967 4680 8304 4709
rect 7967 4679 8015 4680
rect 7923 4677 8015 4679
rect 7923 4674 8008 4677
rect 8269 4642 8304 4680
rect 9346 4653 9380 4859
rect 9793 4839 9825 4867
rect 9413 4831 9825 4839
rect 12354 4888 12386 4953
rect 12724 4888 12764 4889
rect 12354 4886 12766 4888
rect 12354 4860 12734 4886
rect 12760 4860 12766 4886
rect 12354 4852 12766 4860
rect 11788 4837 11820 4838
rect 9413 4805 9419 4831
rect 9445 4805 9825 4831
rect 9413 4803 9825 4805
rect 11785 4832 11820 4837
rect 11785 4812 11792 4832
rect 11812 4812 11820 4832
rect 11785 4804 11820 4812
rect 9415 4802 9455 4803
rect 9793 4738 9825 4803
rect 9793 4718 9797 4738
rect 9818 4718 9825 4738
rect 9793 4711 9825 4718
rect 11341 4739 11373 4746
rect 11341 4719 11348 4739
rect 11369 4719 11373 4739
rect 11341 4654 11373 4719
rect 11711 4654 11751 4655
rect 9346 4645 9381 4653
rect 8060 4640 8095 4641
rect 6166 4470 6581 4499
rect 7719 4498 7752 4499
rect 7716 4493 7752 4498
rect 7716 4473 7723 4493
rect 7743 4473 7752 4493
rect 6166 4469 6575 4470
rect 7716 4468 7752 4473
rect 8039 4633 8095 4640
rect 8039 4613 8068 4633
rect 8088 4613 8095 4633
rect 8039 4608 8095 4613
rect 8264 4633 8313 4642
rect 8264 4614 8272 4633
rect 8298 4614 8313 4633
rect 7716 4465 7751 4468
rect 2758 4420 2793 4423
rect 2196 4255 2211 4274
rect 2237 4255 2245 4274
rect 2196 4246 2245 4255
rect 2414 4275 2470 4280
rect 2414 4255 2421 4275
rect 2441 4255 2470 4275
rect 2414 4248 2470 4255
rect 2757 4415 2793 4420
rect 3934 4418 4343 4419
rect 2757 4395 2766 4415
rect 2786 4395 2793 4415
rect 2757 4390 2793 4395
rect 2757 4389 2790 4390
rect 3928 4389 4343 4418
rect 2414 4247 2449 4248
rect 1128 4235 1163 4243
rect 684 4170 716 4177
rect 684 4150 691 4170
rect 712 4150 716 4170
rect 684 4085 716 4150
rect 1054 4085 1094 4086
rect 684 4083 1096 4085
rect 684 4057 1064 4083
rect 1090 4057 1096 4083
rect 684 4049 1096 4057
rect 684 4021 716 4049
rect 1129 4029 1163 4235
rect 2205 4208 2240 4246
rect 2463 4208 2586 4213
rect 2205 4207 2586 4208
rect 2205 4179 2548 4207
rect 2582 4206 2586 4207
rect 2582 4179 2587 4206
rect 2205 4178 2587 4179
rect 2463 4173 2587 4178
rect 684 4001 689 4021
rect 710 4001 716 4021
rect 684 3994 716 4001
rect 893 4023 933 4028
rect 893 4002 905 4023
rect 927 4002 933 4023
rect 893 3990 933 4002
rect 1107 4024 1163 4029
rect 1107 4004 1114 4024
rect 1134 4004 1163 4024
rect 1107 3997 1163 4004
rect 1220 4098 2177 4117
rect 1107 3996 1142 3997
rect 899 3958 927 3990
rect 1220 3958 1251 4098
rect 2140 4082 2175 4098
rect 2140 4062 2147 4082
rect 2167 4062 2175 4082
rect 2140 4054 2175 4062
rect 899 3927 1251 3958
rect 1696 3989 1728 3996
rect 1696 3969 1703 3989
rect 1724 3969 1728 3989
rect 1696 3904 1728 3969
rect 2066 3904 2106 3905
rect 1696 3902 2108 3904
rect 1696 3876 2076 3902
rect 2102 3876 2108 3902
rect 1696 3868 2108 3876
rect 1130 3853 1162 3854
rect 1127 3848 1162 3853
rect 1127 3828 1134 3848
rect 1154 3828 1162 3848
rect 1127 3820 1162 3828
rect 683 3755 715 3762
rect 683 3735 690 3755
rect 711 3735 715 3755
rect 683 3670 715 3735
rect 1053 3670 1093 3671
rect 683 3668 1095 3670
rect 683 3642 1063 3668
rect 1089 3642 1095 3668
rect 683 3634 1095 3642
rect 683 3606 715 3634
rect 683 3586 688 3606
rect 709 3586 715 3606
rect 683 3579 715 3586
rect 883 3606 933 3615
rect 1128 3614 1162 3820
rect 1696 3840 1728 3868
rect 1696 3820 1701 3840
rect 1722 3820 1728 3840
rect 1696 3813 1728 3820
rect 1903 3841 1945 3849
rect 2141 3848 2175 4054
rect 1903 3821 1912 3841
rect 1936 3821 1945 3841
rect 1903 3809 1945 3821
rect 2119 3843 2175 3848
rect 2119 3823 2126 3843
rect 2146 3823 2175 3843
rect 2119 3816 2175 3823
rect 2119 3815 2154 3816
rect 1905 3780 1940 3809
rect 1905 3779 2215 3780
rect 1790 3773 1826 3777
rect 1790 3754 1798 3773
rect 1818 3754 1826 3773
rect 1790 3751 1826 3754
rect 1791 3723 1825 3751
rect 1905 3745 2232 3779
rect 883 3585 895 3606
rect 917 3585 933 3606
rect 883 3577 933 3585
rect 1106 3609 1162 3614
rect 1106 3589 1113 3609
rect 1133 3589 1162 3609
rect 1106 3582 1162 3589
rect 1263 3695 1826 3723
rect 1106 3581 1141 3582
rect 888 3544 929 3577
rect 1263 3544 1303 3695
rect 888 3515 1303 3544
rect 2192 3521 2232 3745
rect 888 3514 1297 3515
rect 2192 3501 2202 3521
rect 2222 3501 2232 3521
rect 2192 3491 2232 3501
rect 1751 3428 1783 3435
rect 1751 3408 1758 3428
rect 1779 3408 1783 3428
rect 1751 3343 1783 3408
rect 2121 3343 2161 3344
rect 1751 3341 2163 3343
rect 1751 3315 2131 3341
rect 2157 3315 2163 3341
rect 1751 3307 2163 3315
rect 1136 3287 1168 3288
rect 1133 3282 1168 3287
rect 1133 3262 1140 3282
rect 1160 3262 1168 3282
rect 1133 3254 1168 3262
rect 689 3189 721 3196
rect 689 3169 696 3189
rect 717 3169 721 3189
rect 689 3104 721 3169
rect 1059 3104 1099 3105
rect 689 3102 1101 3104
rect 689 3076 1069 3102
rect 1095 3076 1101 3102
rect 689 3068 1101 3076
rect 689 3040 721 3068
rect 1134 3048 1168 3254
rect 1751 3279 1783 3307
rect 1751 3259 1756 3279
rect 1777 3259 1783 3279
rect 1751 3252 1783 3259
rect 1962 3278 2000 3290
rect 2196 3287 2230 3491
rect 1962 3261 1971 3278
rect 1995 3261 2000 3278
rect 1962 3218 2000 3261
rect 2174 3282 2230 3287
rect 2174 3262 2181 3282
rect 2201 3262 2230 3282
rect 2174 3255 2230 3262
rect 2174 3254 2209 3255
rect 2308 3218 2392 3223
rect 1962 3189 2392 3218
rect 689 3020 694 3040
rect 715 3020 721 3040
rect 689 3013 721 3020
rect 898 3042 938 3047
rect 898 3021 910 3042
rect 932 3021 938 3042
rect 898 3009 938 3021
rect 1112 3043 1168 3048
rect 1112 3023 1119 3043
rect 1139 3023 1168 3043
rect 1112 3016 1168 3023
rect 1225 3117 2182 3136
rect 1112 3015 1147 3016
rect 904 2977 932 3009
rect 1225 2977 1256 3117
rect 2145 3101 2180 3117
rect 2145 3081 2152 3101
rect 2172 3081 2180 3101
rect 2145 3073 2180 3081
rect 904 2946 1256 2977
rect 1701 3008 1733 3015
rect 1701 2988 1708 3008
rect 1729 2988 1733 3008
rect 1701 2923 1733 2988
rect 2071 2923 2111 2924
rect 1701 2921 2113 2923
rect 1701 2895 2081 2921
rect 2107 2895 2113 2921
rect 1701 2887 2113 2895
rect 1135 2872 1167 2873
rect 1132 2867 1167 2872
rect 1132 2847 1139 2867
rect 1159 2847 1167 2867
rect 1132 2839 1167 2847
rect 688 2774 720 2781
rect 688 2754 695 2774
rect 716 2754 720 2774
rect 688 2689 720 2754
rect 1058 2689 1098 2690
rect 688 2687 1100 2689
rect 688 2661 1068 2687
rect 1094 2661 1100 2687
rect 688 2653 1100 2661
rect 688 2625 720 2653
rect 688 2605 693 2625
rect 714 2605 720 2625
rect 688 2598 720 2605
rect 888 2625 938 2634
rect 1133 2633 1167 2839
rect 1701 2859 1733 2887
rect 1701 2839 1706 2859
rect 1727 2839 1733 2859
rect 1906 2861 1948 2870
rect 2146 2867 2180 3073
rect 1906 2847 1916 2861
rect 1701 2832 1733 2839
rect 1905 2841 1916 2847
rect 1940 2841 1948 2861
rect 1905 2830 1948 2841
rect 2124 2862 2180 2867
rect 2124 2842 2131 2862
rect 2151 2842 2180 2862
rect 2124 2835 2180 2842
rect 2124 2834 2159 2835
rect 1905 2800 1945 2830
rect 1795 2792 1831 2796
rect 1795 2773 1803 2792
rect 1823 2773 1831 2792
rect 1795 2770 1831 2773
rect 1905 2795 2252 2800
rect 1796 2742 1830 2770
rect 1905 2769 2224 2795
rect 2243 2769 2252 2795
rect 1905 2765 2252 2769
rect 888 2604 900 2625
rect 922 2604 938 2625
rect 888 2596 938 2604
rect 1111 2628 1167 2633
rect 1111 2608 1118 2628
rect 1138 2608 1167 2628
rect 1111 2601 1167 2608
rect 1268 2714 1831 2742
rect 1111 2600 1146 2601
rect 893 2563 934 2596
rect 1268 2563 1308 2714
rect 2357 2595 2392 3189
rect 2757 2736 2789 4389
rect 3928 4238 3968 4389
rect 4302 4356 4343 4389
rect 7272 4400 7304 4407
rect 7272 4380 7279 4400
rect 7300 4380 7304 4400
rect 4090 4351 4125 4352
rect 3405 4210 3968 4238
rect 4069 4344 4125 4351
rect 4069 4324 4098 4344
rect 4118 4324 4125 4344
rect 4069 4319 4125 4324
rect 4298 4348 4348 4356
rect 4298 4327 4314 4348
rect 4336 4327 4348 4348
rect 2984 4183 3331 4187
rect 2984 4157 2993 4183
rect 3012 4157 3331 4183
rect 3406 4182 3440 4210
rect 2984 4152 3331 4157
rect 3405 4179 3441 4182
rect 3405 4160 3413 4179
rect 3433 4160 3441 4179
rect 3405 4156 3441 4160
rect 3291 4122 3331 4152
rect 3077 4117 3112 4118
rect 3056 4110 3112 4117
rect 3056 4090 3085 4110
rect 3105 4090 3112 4110
rect 3056 4085 3112 4090
rect 3288 4111 3331 4122
rect 3288 4091 3296 4111
rect 3320 4105 3331 4111
rect 3503 4113 3535 4120
rect 3320 4091 3330 4105
rect 3056 3879 3090 4085
rect 3288 4082 3330 4091
rect 3503 4093 3509 4113
rect 3530 4093 3535 4113
rect 3503 4065 3535 4093
rect 4069 4113 4103 4319
rect 4298 4318 4348 4327
rect 4516 4347 4548 4354
rect 4516 4327 4522 4347
rect 4543 4327 4548 4347
rect 4516 4299 4548 4327
rect 4136 4291 4548 4299
rect 4136 4265 4142 4291
rect 4168 4265 4548 4291
rect 4136 4263 4548 4265
rect 4138 4262 4178 4263
rect 4516 4198 4548 4263
rect 7272 4315 7304 4380
rect 7642 4315 7682 4316
rect 7272 4313 7684 4315
rect 7272 4287 7652 4313
rect 7678 4287 7684 4313
rect 7272 4279 7684 4287
rect 7272 4251 7304 4279
rect 6412 4247 6444 4248
rect 6409 4242 6444 4247
rect 6409 4222 6416 4242
rect 6436 4222 6444 4242
rect 7272 4231 7277 4251
rect 7298 4231 7304 4251
rect 7272 4224 7304 4231
rect 7477 4253 7526 4263
rect 7717 4259 7751 4465
rect 8039 4402 8073 4608
rect 8264 4604 8313 4614
rect 8486 4636 8518 4643
rect 8486 4616 8492 4636
rect 8513 4616 8518 4636
rect 9346 4625 9354 4645
rect 9374 4625 9381 4645
rect 9346 4620 9381 4625
rect 11341 4652 11753 4654
rect 11341 4626 11721 4652
rect 11747 4626 11753 4652
rect 9346 4619 9378 4620
rect 8486 4588 8518 4616
rect 8106 4580 8518 4588
rect 8106 4554 8112 4580
rect 8138 4554 8518 4580
rect 11341 4618 11753 4626
rect 11341 4590 11373 4618
rect 11341 4570 11346 4590
rect 11367 4570 11373 4590
rect 11341 4563 11373 4570
rect 11541 4590 11591 4599
rect 11786 4598 11820 4804
rect 12354 4824 12386 4852
rect 12354 4804 12359 4824
rect 12380 4804 12386 4824
rect 12559 4826 12601 4835
rect 12799 4832 12833 5038
rect 12559 4812 12569 4826
rect 12354 4797 12386 4804
rect 12558 4806 12569 4812
rect 12593 4806 12601 4826
rect 12558 4795 12601 4806
rect 12777 4827 12833 4832
rect 12777 4807 12784 4827
rect 12804 4807 12833 4827
rect 12777 4800 12833 4807
rect 12777 4799 12812 4800
rect 12558 4765 12598 4795
rect 12448 4757 12484 4761
rect 12448 4738 12456 4757
rect 12476 4738 12484 4757
rect 12448 4735 12484 4738
rect 12558 4760 12905 4765
rect 12449 4707 12483 4735
rect 12558 4734 12877 4760
rect 12896 4734 12905 4760
rect 12558 4730 12905 4734
rect 11541 4569 11553 4590
rect 11575 4569 11591 4590
rect 11541 4561 11591 4569
rect 11764 4593 11820 4598
rect 11764 4573 11771 4593
rect 11791 4573 11820 4593
rect 11764 4566 11820 4573
rect 11921 4679 12484 4707
rect 11764 4565 11799 4566
rect 8106 4552 8518 4554
rect 8108 4551 8148 4552
rect 8486 4487 8518 4552
rect 11546 4528 11587 4561
rect 11921 4528 11961 4679
rect 13100 4528 13132 6181
rect 13497 5728 13532 6322
rect 14581 6203 14621 6354
rect 14955 6321 14996 6354
rect 17838 6380 17845 6400
rect 17866 6380 17870 6400
rect 14743 6316 14778 6317
rect 14058 6175 14621 6203
rect 14722 6309 14778 6316
rect 14722 6289 14751 6309
rect 14771 6289 14778 6309
rect 14722 6284 14778 6289
rect 14951 6313 15001 6321
rect 14951 6292 14967 6313
rect 14989 6292 15001 6313
rect 13637 6148 13984 6152
rect 13637 6122 13646 6148
rect 13665 6122 13984 6148
rect 14059 6147 14093 6175
rect 13637 6117 13984 6122
rect 14058 6144 14094 6147
rect 14058 6125 14066 6144
rect 14086 6125 14094 6144
rect 14058 6121 14094 6125
rect 13944 6087 13984 6117
rect 13730 6082 13765 6083
rect 13709 6075 13765 6082
rect 13709 6055 13738 6075
rect 13758 6055 13765 6075
rect 13709 6050 13765 6055
rect 13941 6076 13984 6087
rect 13941 6056 13949 6076
rect 13973 6070 13984 6076
rect 14156 6078 14188 6085
rect 13973 6056 13983 6070
rect 13709 5844 13743 6050
rect 13941 6047 13983 6056
rect 14156 6058 14162 6078
rect 14183 6058 14188 6078
rect 14156 6030 14188 6058
rect 14722 6078 14756 6284
rect 14951 6283 15001 6292
rect 15169 6312 15201 6319
rect 15169 6292 15175 6312
rect 15196 6292 15201 6312
rect 15169 6264 15201 6292
rect 14789 6256 15201 6264
rect 14789 6230 14795 6256
rect 14821 6230 15201 6256
rect 14789 6228 15201 6230
rect 14791 6227 14831 6228
rect 15169 6163 15201 6228
rect 17838 6315 17870 6380
rect 18208 6315 18248 6316
rect 17838 6313 18250 6315
rect 17838 6287 18218 6313
rect 18244 6287 18250 6313
rect 17838 6279 18250 6287
rect 17838 6251 17870 6279
rect 17838 6231 17843 6251
rect 17864 6231 17870 6251
rect 17838 6224 17870 6231
rect 18042 6256 18089 6262
rect 18283 6259 18317 6465
rect 18775 6335 18809 6541
rect 19222 6521 19254 6549
rect 18842 6513 19254 6521
rect 18842 6487 18848 6513
rect 18874 6487 19254 6513
rect 18842 6485 19254 6487
rect 18844 6484 18884 6485
rect 19222 6420 19254 6485
rect 19222 6400 19226 6420
rect 19247 6400 19254 6420
rect 19222 6393 19254 6400
rect 19868 6362 20277 6363
rect 18775 6329 18810 6335
rect 19862 6333 20277 6362
rect 18775 6327 18813 6329
rect 18775 6307 18783 6327
rect 18803 6307 18813 6327
rect 18775 6301 18813 6307
rect 18042 6230 18052 6256
rect 18077 6230 18089 6256
rect 18042 6228 18089 6230
rect 18261 6254 18317 6259
rect 18261 6234 18268 6254
rect 18288 6234 18317 6254
rect 17065 6212 17097 6213
rect 17062 6207 17097 6212
rect 17062 6187 17069 6207
rect 17089 6187 17097 6207
rect 17062 6179 17097 6187
rect 15169 6143 15173 6163
rect 15194 6143 15201 6163
rect 15169 6136 15201 6143
rect 16618 6114 16650 6121
rect 16618 6094 16625 6114
rect 16646 6094 16650 6114
rect 14722 6070 14757 6078
rect 14722 6050 14730 6070
rect 14750 6050 14757 6070
rect 14722 6045 14757 6050
rect 14722 6044 14754 6045
rect 13776 6022 14188 6030
rect 13776 5996 13782 6022
rect 13808 5996 14188 6022
rect 13776 5994 14188 5996
rect 13778 5993 13818 5994
rect 14156 5929 14188 5994
rect 16618 6029 16650 6094
rect 16988 6029 17028 6030
rect 16618 6027 17030 6029
rect 16618 6001 16998 6027
rect 17024 6001 17030 6027
rect 16618 5993 17030 6001
rect 14156 5909 14160 5929
rect 14181 5909 14188 5929
rect 14156 5902 14188 5909
rect 14633 5940 14985 5971
rect 13709 5836 13744 5844
rect 13709 5816 13717 5836
rect 13737 5816 13744 5836
rect 13709 5800 13744 5816
rect 14633 5800 14664 5940
rect 14957 5908 14985 5940
rect 16618 5965 16650 5993
rect 17063 5973 17097 6179
rect 18047 6193 18084 6228
rect 18261 6227 18317 6234
rect 18261 6226 18296 6227
rect 18381 6193 18413 6195
rect 18047 6160 18417 6193
rect 16618 5945 16623 5965
rect 16644 5945 16650 5965
rect 16618 5938 16650 5945
rect 16827 5967 16867 5972
rect 16827 5946 16839 5967
rect 16861 5946 16867 5967
rect 16827 5934 16867 5946
rect 17041 5968 17097 5973
rect 17041 5948 17048 5968
rect 17068 5948 17097 5968
rect 17041 5941 17097 5948
rect 17154 6042 18111 6061
rect 17041 5940 17076 5941
rect 14742 5901 14777 5902
rect 13707 5781 14664 5800
rect 14721 5894 14777 5901
rect 14721 5874 14750 5894
rect 14770 5874 14777 5894
rect 14721 5869 14777 5874
rect 14951 5896 14991 5908
rect 14951 5875 14957 5896
rect 14979 5875 14991 5896
rect 14951 5870 14991 5875
rect 15168 5897 15200 5904
rect 15168 5877 15174 5897
rect 15195 5877 15200 5897
rect 13497 5699 13927 5728
rect 13497 5694 13581 5699
rect 13680 5662 13715 5663
rect 13659 5655 13715 5662
rect 13659 5635 13688 5655
rect 13708 5635 13715 5655
rect 13659 5630 13715 5635
rect 13889 5656 13927 5699
rect 13889 5639 13894 5656
rect 13918 5639 13927 5656
rect 13659 5426 13693 5630
rect 13889 5627 13927 5639
rect 14106 5658 14138 5665
rect 14106 5638 14112 5658
rect 14133 5638 14138 5658
rect 14106 5610 14138 5638
rect 14721 5663 14755 5869
rect 15168 5849 15200 5877
rect 16833 5902 16861 5934
rect 17154 5902 17185 6042
rect 18074 6026 18109 6042
rect 18074 6006 18081 6026
rect 18101 6006 18109 6026
rect 18074 5998 18109 6006
rect 16833 5871 17185 5902
rect 17630 5933 17662 5940
rect 17630 5913 17637 5933
rect 17658 5913 17662 5933
rect 14788 5841 15200 5849
rect 14788 5815 14794 5841
rect 14820 5815 15200 5841
rect 14788 5813 15200 5815
rect 14790 5812 14830 5813
rect 15168 5748 15200 5813
rect 17630 5848 17662 5913
rect 18000 5848 18040 5849
rect 17630 5846 18042 5848
rect 17630 5820 18010 5846
rect 18036 5820 18042 5846
rect 17630 5812 18042 5820
rect 17064 5797 17096 5798
rect 17061 5792 17096 5797
rect 17061 5772 17068 5792
rect 17088 5772 17096 5792
rect 17061 5764 17096 5772
rect 15168 5728 15172 5748
rect 15193 5728 15200 5748
rect 15168 5721 15200 5728
rect 16617 5699 16649 5706
rect 16617 5679 16624 5699
rect 16645 5679 16649 5699
rect 14721 5655 14756 5663
rect 14721 5635 14729 5655
rect 14749 5635 14756 5655
rect 14721 5630 14756 5635
rect 14721 5629 14753 5630
rect 13726 5602 14138 5610
rect 13726 5576 13732 5602
rect 13758 5576 14138 5602
rect 13726 5574 14138 5576
rect 13728 5573 13768 5574
rect 14106 5509 14138 5574
rect 16617 5614 16649 5679
rect 16987 5614 17027 5615
rect 16617 5612 17029 5614
rect 16617 5586 16997 5612
rect 17023 5586 17029 5612
rect 16617 5578 17029 5586
rect 16617 5550 16649 5578
rect 16617 5530 16622 5550
rect 16643 5530 16649 5550
rect 16617 5523 16649 5530
rect 16817 5550 16867 5559
rect 17062 5558 17096 5764
rect 17630 5784 17662 5812
rect 17630 5764 17635 5784
rect 17656 5764 17662 5784
rect 17630 5757 17662 5764
rect 17837 5785 17879 5793
rect 18075 5792 18109 5998
rect 17837 5765 17846 5785
rect 17870 5765 17879 5785
rect 17837 5753 17879 5765
rect 18053 5787 18109 5792
rect 18053 5767 18060 5787
rect 18080 5767 18109 5787
rect 18053 5760 18109 5767
rect 18053 5759 18088 5760
rect 17839 5724 17874 5753
rect 17839 5723 18149 5724
rect 17724 5717 17760 5721
rect 17724 5698 17732 5717
rect 17752 5698 17760 5717
rect 17724 5695 17760 5698
rect 17725 5667 17759 5695
rect 17839 5689 18166 5723
rect 16817 5529 16829 5550
rect 16851 5529 16867 5550
rect 16817 5521 16867 5529
rect 17040 5553 17096 5558
rect 17040 5533 17047 5553
rect 17067 5533 17096 5553
rect 17040 5526 17096 5533
rect 17197 5639 17760 5667
rect 17040 5525 17075 5526
rect 14106 5489 14110 5509
rect 14131 5489 14138 5509
rect 14106 5482 14138 5489
rect 16822 5488 16863 5521
rect 17197 5488 17237 5639
rect 16822 5459 17237 5488
rect 18126 5465 18166 5689
rect 16822 5458 17231 5459
rect 18126 5445 18136 5465
rect 18156 5445 18166 5465
rect 18126 5435 18166 5445
rect 13657 5416 13697 5426
rect 13657 5396 13667 5416
rect 13687 5396 13697 5416
rect 14592 5402 15001 5403
rect 13657 5172 13697 5396
rect 14586 5373 15001 5402
rect 14586 5222 14626 5373
rect 14960 5340 15001 5373
rect 17685 5372 17717 5379
rect 17685 5352 17692 5372
rect 17713 5352 17717 5372
rect 14748 5335 14783 5336
rect 14063 5194 14626 5222
rect 14727 5328 14783 5335
rect 14727 5308 14756 5328
rect 14776 5308 14783 5328
rect 14727 5303 14783 5308
rect 14956 5332 15006 5340
rect 14956 5311 14972 5332
rect 14994 5311 15006 5332
rect 13657 5138 13984 5172
rect 14064 5166 14098 5194
rect 14063 5163 14099 5166
rect 14063 5144 14071 5163
rect 14091 5144 14099 5163
rect 14063 5140 14099 5144
rect 13674 5137 13984 5138
rect 13949 5108 13984 5137
rect 13735 5101 13770 5102
rect 13714 5094 13770 5101
rect 13714 5074 13743 5094
rect 13763 5074 13770 5094
rect 13714 5069 13770 5074
rect 13944 5096 13986 5108
rect 13944 5076 13953 5096
rect 13977 5076 13986 5096
rect 13714 4863 13748 5069
rect 13944 5068 13986 5076
rect 14161 5097 14193 5104
rect 14161 5077 14167 5097
rect 14188 5077 14193 5097
rect 14161 5049 14193 5077
rect 14727 5097 14761 5303
rect 14956 5302 15006 5311
rect 15174 5331 15206 5338
rect 15174 5311 15180 5331
rect 15201 5311 15206 5331
rect 15174 5283 15206 5311
rect 14794 5275 15206 5283
rect 14794 5249 14800 5275
rect 14826 5249 15206 5275
rect 14794 5247 15206 5249
rect 14796 5246 14836 5247
rect 15174 5182 15206 5247
rect 17685 5287 17717 5352
rect 18055 5287 18095 5288
rect 17685 5285 18097 5287
rect 17685 5259 18065 5285
rect 18091 5259 18097 5285
rect 17685 5251 18097 5259
rect 17070 5231 17102 5232
rect 17067 5226 17102 5231
rect 17067 5206 17074 5226
rect 17094 5206 17102 5226
rect 17067 5198 17102 5206
rect 15174 5162 15178 5182
rect 15199 5162 15206 5182
rect 15174 5155 15206 5162
rect 16623 5133 16655 5140
rect 16623 5113 16630 5133
rect 16651 5113 16655 5133
rect 14727 5089 14762 5097
rect 14727 5069 14735 5089
rect 14755 5069 14762 5089
rect 14727 5064 14762 5069
rect 14727 5063 14759 5064
rect 13781 5041 14193 5049
rect 13781 5015 13787 5041
rect 13813 5015 14193 5041
rect 13781 5013 14193 5015
rect 13783 5012 13823 5013
rect 14161 4948 14193 5013
rect 16623 5048 16655 5113
rect 16993 5048 17033 5049
rect 16623 5046 17035 5048
rect 16623 5020 17003 5046
rect 17029 5020 17035 5046
rect 16623 5012 17035 5020
rect 14161 4928 14165 4948
rect 14186 4928 14193 4948
rect 14161 4921 14193 4928
rect 14638 4959 14990 4990
rect 13714 4855 13749 4863
rect 13714 4835 13722 4855
rect 13742 4835 13749 4855
rect 13714 4819 13749 4835
rect 14638 4819 14669 4959
rect 14962 4927 14990 4959
rect 16623 4984 16655 5012
rect 17068 4992 17102 5198
rect 17685 5223 17717 5251
rect 18130 5231 18164 5435
rect 17685 5203 17690 5223
rect 17711 5203 17717 5223
rect 17685 5196 17717 5203
rect 17896 5223 17933 5229
rect 17896 5204 17902 5223
rect 17925 5204 17933 5223
rect 17896 5199 17933 5204
rect 18108 5226 18164 5231
rect 18108 5206 18115 5226
rect 18135 5206 18164 5226
rect 18108 5199 18164 5206
rect 17904 5162 17928 5199
rect 18108 5198 18143 5199
rect 17904 5160 18272 5162
rect 17904 5155 18277 5160
rect 17904 5137 18250 5155
rect 18270 5137 18277 5155
rect 17904 5132 18277 5137
rect 18248 5130 18277 5132
rect 16623 4964 16628 4984
rect 16649 4964 16655 4984
rect 16623 4957 16655 4964
rect 16832 4986 16872 4991
rect 16832 4965 16844 4986
rect 16866 4965 16872 4986
rect 16832 4953 16872 4965
rect 17046 4987 17102 4992
rect 17046 4967 17053 4987
rect 17073 4967 17102 4987
rect 17046 4960 17102 4967
rect 17159 5061 18116 5080
rect 17046 4959 17081 4960
rect 14747 4920 14782 4921
rect 13712 4800 14669 4819
rect 14726 4913 14782 4920
rect 14726 4893 14755 4913
rect 14775 4893 14782 4913
rect 14726 4888 14782 4893
rect 14956 4915 14996 4927
rect 14956 4894 14962 4915
rect 14984 4894 14996 4915
rect 14956 4889 14996 4894
rect 15173 4916 15205 4923
rect 15173 4896 15179 4916
rect 15200 4896 15205 4916
rect 13310 4743 13395 4746
rect 13303 4739 13395 4743
rect 13303 4738 13684 4739
rect 13303 4708 13310 4738
rect 13347 4709 13684 4738
rect 13347 4708 13395 4709
rect 13303 4706 13395 4708
rect 13303 4703 13388 4706
rect 13649 4671 13684 4709
rect 14726 4682 14760 4888
rect 15173 4868 15205 4896
rect 16838 4921 16866 4953
rect 17159 4921 17190 5061
rect 18079 5045 18114 5061
rect 18079 5025 18086 5045
rect 18106 5025 18114 5045
rect 18079 5017 18114 5025
rect 16838 4890 17190 4921
rect 17635 4952 17667 4959
rect 17635 4932 17642 4952
rect 17663 4932 17667 4952
rect 14793 4860 15205 4868
rect 14793 4834 14799 4860
rect 14825 4834 15205 4860
rect 14793 4832 15205 4834
rect 14795 4831 14835 4832
rect 15173 4767 15205 4832
rect 17635 4867 17667 4932
rect 18005 4867 18045 4868
rect 17635 4865 18047 4867
rect 17635 4839 18015 4865
rect 18041 4839 18047 4865
rect 17635 4831 18047 4839
rect 17069 4816 17101 4817
rect 17066 4811 17101 4816
rect 17066 4791 17073 4811
rect 17093 4791 17101 4811
rect 17066 4783 17101 4791
rect 15173 4747 15177 4767
rect 15198 4747 15205 4767
rect 15173 4740 15205 4747
rect 16622 4718 16654 4725
rect 16622 4698 16629 4718
rect 16650 4698 16654 4718
rect 14726 4674 14761 4682
rect 13440 4669 13475 4670
rect 11546 4499 11961 4528
rect 13099 4527 13132 4528
rect 13096 4522 13132 4527
rect 13096 4502 13103 4522
rect 13123 4502 13132 4522
rect 11546 4498 11955 4499
rect 13096 4497 13132 4502
rect 13419 4662 13475 4669
rect 13419 4642 13448 4662
rect 13468 4642 13475 4662
rect 13419 4637 13475 4642
rect 13644 4662 13693 4671
rect 13644 4643 13652 4662
rect 13678 4643 13693 4662
rect 13096 4494 13131 4497
rect 8486 4467 8490 4487
rect 8511 4467 8518 4487
rect 8486 4460 8518 4467
rect 12652 4429 12684 4436
rect 12652 4409 12659 4429
rect 12680 4409 12684 4429
rect 8039 4399 8074 4402
rect 7477 4234 7492 4253
rect 7518 4234 7526 4253
rect 7477 4225 7526 4234
rect 7695 4254 7751 4259
rect 7695 4234 7702 4254
rect 7722 4234 7751 4254
rect 7695 4227 7751 4234
rect 8038 4394 8074 4399
rect 9215 4397 9624 4398
rect 8038 4374 8047 4394
rect 8067 4374 8074 4394
rect 8038 4369 8074 4374
rect 8038 4368 8071 4369
rect 9209 4368 9624 4397
rect 7695 4226 7730 4227
rect 6409 4214 6444 4222
rect 4516 4178 4520 4198
rect 4541 4178 4548 4198
rect 4516 4171 4548 4178
rect 5965 4149 5997 4156
rect 5965 4129 5972 4149
rect 5993 4129 5997 4149
rect 4069 4105 4104 4113
rect 4069 4085 4077 4105
rect 4097 4085 4104 4105
rect 4069 4080 4104 4085
rect 4069 4079 4101 4080
rect 3123 4057 3535 4065
rect 3123 4031 3129 4057
rect 3155 4031 3535 4057
rect 3123 4029 3535 4031
rect 3125 4028 3165 4029
rect 3503 3964 3535 4029
rect 5965 4064 5997 4129
rect 6335 4064 6375 4065
rect 5965 4062 6377 4064
rect 5965 4036 6345 4062
rect 6371 4036 6377 4062
rect 5965 4028 6377 4036
rect 3503 3944 3507 3964
rect 3528 3944 3535 3964
rect 3503 3937 3535 3944
rect 3980 3975 4332 4006
rect 3056 3871 3091 3879
rect 3056 3851 3064 3871
rect 3084 3851 3091 3871
rect 3056 3835 3091 3851
rect 3980 3835 4011 3975
rect 4304 3943 4332 3975
rect 5965 4000 5997 4028
rect 6410 4008 6444 4214
rect 7486 4187 7521 4225
rect 7744 4187 7867 4192
rect 7486 4186 7867 4187
rect 7486 4158 7829 4186
rect 7863 4185 7867 4186
rect 7863 4158 7868 4185
rect 7486 4157 7868 4158
rect 7744 4152 7868 4157
rect 5965 3980 5970 4000
rect 5991 3980 5997 4000
rect 5965 3973 5997 3980
rect 6174 4002 6214 4007
rect 6174 3981 6186 4002
rect 6208 3981 6214 4002
rect 6174 3969 6214 3981
rect 6388 4003 6444 4008
rect 6388 3983 6395 4003
rect 6415 3983 6444 4003
rect 6388 3976 6444 3983
rect 6501 4077 7458 4096
rect 6388 3975 6423 3976
rect 4089 3936 4124 3937
rect 3054 3816 4011 3835
rect 4068 3929 4124 3936
rect 4068 3909 4097 3929
rect 4117 3909 4124 3929
rect 4068 3904 4124 3909
rect 4298 3931 4338 3943
rect 4298 3910 4304 3931
rect 4326 3910 4338 3931
rect 4298 3905 4338 3910
rect 4515 3932 4547 3939
rect 4515 3912 4521 3932
rect 4542 3912 4547 3932
rect 2893 3764 2922 3766
rect 2893 3759 3266 3764
rect 2893 3741 2900 3759
rect 2920 3741 3266 3759
rect 2893 3736 3266 3741
rect 2898 3734 3266 3736
rect 3027 3697 3062 3698
rect 3242 3697 3266 3734
rect 3006 3690 3062 3697
rect 3006 3670 3035 3690
rect 3055 3670 3062 3690
rect 3006 3665 3062 3670
rect 3237 3692 3274 3697
rect 3237 3673 3245 3692
rect 3268 3673 3274 3692
rect 3237 3667 3274 3673
rect 3453 3693 3485 3700
rect 3453 3673 3459 3693
rect 3480 3673 3485 3693
rect 3006 3461 3040 3665
rect 3453 3645 3485 3673
rect 4068 3698 4102 3904
rect 4515 3884 4547 3912
rect 6180 3937 6208 3969
rect 6501 3937 6532 4077
rect 7421 4061 7456 4077
rect 7421 4041 7428 4061
rect 7448 4041 7456 4061
rect 7421 4033 7456 4041
rect 6180 3906 6532 3937
rect 6977 3968 7009 3975
rect 6977 3948 6984 3968
rect 7005 3948 7009 3968
rect 4135 3876 4547 3884
rect 4135 3850 4141 3876
rect 4167 3850 4547 3876
rect 4135 3848 4547 3850
rect 4137 3847 4177 3848
rect 4515 3783 4547 3848
rect 6977 3883 7009 3948
rect 7347 3883 7387 3884
rect 6977 3881 7389 3883
rect 6977 3855 7357 3881
rect 7383 3855 7389 3881
rect 6977 3847 7389 3855
rect 6411 3832 6443 3833
rect 6408 3827 6443 3832
rect 6408 3807 6415 3827
rect 6435 3807 6443 3827
rect 6408 3799 6443 3807
rect 4515 3763 4519 3783
rect 4540 3763 4547 3783
rect 4515 3756 4547 3763
rect 5964 3734 5996 3741
rect 5964 3714 5971 3734
rect 5992 3714 5996 3734
rect 4068 3690 4103 3698
rect 4068 3670 4076 3690
rect 4096 3670 4103 3690
rect 4068 3665 4103 3670
rect 4068 3664 4100 3665
rect 3073 3637 3485 3645
rect 3073 3611 3079 3637
rect 3105 3611 3485 3637
rect 3073 3609 3485 3611
rect 3075 3608 3115 3609
rect 3453 3544 3485 3609
rect 5964 3649 5996 3714
rect 6334 3649 6374 3650
rect 5964 3647 6376 3649
rect 5964 3621 6344 3647
rect 6370 3621 6376 3647
rect 5964 3613 6376 3621
rect 5964 3585 5996 3613
rect 5964 3565 5969 3585
rect 5990 3565 5996 3585
rect 5964 3558 5996 3565
rect 6164 3585 6214 3594
rect 6409 3593 6443 3799
rect 6977 3819 7009 3847
rect 6977 3799 6982 3819
rect 7003 3799 7009 3819
rect 6977 3792 7009 3799
rect 7184 3820 7226 3828
rect 7422 3827 7456 4033
rect 7184 3800 7193 3820
rect 7217 3800 7226 3820
rect 7184 3788 7226 3800
rect 7400 3822 7456 3827
rect 7400 3802 7407 3822
rect 7427 3802 7456 3822
rect 7400 3795 7456 3802
rect 7400 3794 7435 3795
rect 7186 3759 7221 3788
rect 7186 3758 7496 3759
rect 7071 3752 7107 3756
rect 7071 3733 7079 3752
rect 7099 3733 7107 3752
rect 7071 3730 7107 3733
rect 7072 3702 7106 3730
rect 7186 3724 7513 3758
rect 6164 3564 6176 3585
rect 6198 3564 6214 3585
rect 6164 3556 6214 3564
rect 6387 3588 6443 3593
rect 6387 3568 6394 3588
rect 6414 3568 6443 3588
rect 6387 3561 6443 3568
rect 6544 3674 7107 3702
rect 6387 3560 6422 3561
rect 3453 3524 3457 3544
rect 3478 3524 3485 3544
rect 3453 3517 3485 3524
rect 6169 3523 6210 3556
rect 6544 3523 6584 3674
rect 6169 3494 6584 3523
rect 7473 3500 7513 3724
rect 6169 3493 6578 3494
rect 7473 3480 7483 3500
rect 7503 3480 7513 3500
rect 7473 3470 7513 3480
rect 3004 3451 3044 3461
rect 3004 3431 3014 3451
rect 3034 3431 3044 3451
rect 3939 3437 4348 3438
rect 3004 3207 3044 3431
rect 3933 3408 4348 3437
rect 3933 3257 3973 3408
rect 4307 3375 4348 3408
rect 7032 3407 7064 3414
rect 7032 3387 7039 3407
rect 7060 3387 7064 3407
rect 4095 3370 4130 3371
rect 3410 3229 3973 3257
rect 4074 3363 4130 3370
rect 4074 3343 4103 3363
rect 4123 3343 4130 3363
rect 4074 3338 4130 3343
rect 4303 3367 4353 3375
rect 4303 3346 4319 3367
rect 4341 3346 4353 3367
rect 3004 3173 3331 3207
rect 3411 3201 3445 3229
rect 3410 3198 3446 3201
rect 3410 3179 3418 3198
rect 3438 3179 3446 3198
rect 3410 3175 3446 3179
rect 3021 3172 3331 3173
rect 3296 3143 3331 3172
rect 3082 3136 3117 3137
rect 3061 3129 3117 3136
rect 3061 3109 3090 3129
rect 3110 3109 3117 3129
rect 3061 3104 3117 3109
rect 3291 3131 3333 3143
rect 3291 3111 3300 3131
rect 3324 3111 3333 3131
rect 3061 2898 3095 3104
rect 3291 3103 3333 3111
rect 3508 3132 3540 3139
rect 3508 3112 3514 3132
rect 3535 3112 3540 3132
rect 3508 3084 3540 3112
rect 4074 3132 4108 3338
rect 4303 3337 4353 3346
rect 4521 3366 4553 3373
rect 4521 3346 4527 3366
rect 4548 3346 4553 3366
rect 4521 3318 4553 3346
rect 4141 3310 4553 3318
rect 4141 3284 4147 3310
rect 4173 3284 4553 3310
rect 4141 3282 4553 3284
rect 4143 3281 4183 3282
rect 4521 3217 4553 3282
rect 7032 3322 7064 3387
rect 7402 3322 7442 3323
rect 7032 3320 7444 3322
rect 7032 3294 7412 3320
rect 7438 3294 7444 3320
rect 7032 3286 7444 3294
rect 6417 3266 6449 3267
rect 6414 3261 6449 3266
rect 6414 3241 6421 3261
rect 6441 3241 6449 3261
rect 6414 3233 6449 3241
rect 4521 3197 4525 3217
rect 4546 3197 4553 3217
rect 4521 3190 4553 3197
rect 5970 3168 6002 3175
rect 5970 3148 5977 3168
rect 5998 3148 6002 3168
rect 4074 3124 4109 3132
rect 4074 3104 4082 3124
rect 4102 3104 4109 3124
rect 4074 3099 4109 3104
rect 4074 3098 4106 3099
rect 3128 3076 3540 3084
rect 3128 3050 3134 3076
rect 3160 3050 3540 3076
rect 3128 3048 3540 3050
rect 3130 3047 3170 3048
rect 3508 2983 3540 3048
rect 5970 3083 6002 3148
rect 6340 3083 6380 3084
rect 5970 3081 6382 3083
rect 5970 3055 6350 3081
rect 6376 3055 6382 3081
rect 5970 3047 6382 3055
rect 3508 2963 3512 2983
rect 3533 2963 3540 2983
rect 3508 2956 3540 2963
rect 3985 2994 4337 3025
rect 3061 2890 3096 2898
rect 3061 2870 3069 2890
rect 3089 2870 3096 2890
rect 3061 2854 3096 2870
rect 3985 2854 4016 2994
rect 4309 2962 4337 2994
rect 5970 3019 6002 3047
rect 6415 3027 6449 3233
rect 7032 3258 7064 3286
rect 7032 3238 7037 3258
rect 7058 3238 7064 3258
rect 7032 3231 7064 3238
rect 7243 3257 7281 3269
rect 7477 3266 7511 3470
rect 7243 3240 7252 3257
rect 7276 3240 7281 3257
rect 7243 3197 7281 3240
rect 7455 3261 7511 3266
rect 7455 3241 7462 3261
rect 7482 3241 7511 3261
rect 7455 3234 7511 3241
rect 7455 3233 7490 3234
rect 7589 3197 7673 3202
rect 7243 3168 7673 3197
rect 5970 2999 5975 3019
rect 5996 2999 6002 3019
rect 5970 2992 6002 2999
rect 6179 3021 6219 3026
rect 6179 3000 6191 3021
rect 6213 3000 6219 3021
rect 6179 2988 6219 3000
rect 6393 3022 6449 3027
rect 6393 3002 6400 3022
rect 6420 3002 6449 3022
rect 6393 2995 6449 3002
rect 6506 3096 7463 3115
rect 6393 2994 6428 2995
rect 4094 2955 4129 2956
rect 3059 2835 4016 2854
rect 4073 2948 4129 2955
rect 4073 2928 4102 2948
rect 4122 2928 4129 2948
rect 4073 2923 4129 2928
rect 4303 2950 4343 2962
rect 4303 2929 4309 2950
rect 4331 2929 4343 2950
rect 4303 2924 4343 2929
rect 4520 2951 4552 2958
rect 4520 2931 4526 2951
rect 4547 2931 4552 2951
rect 2753 2703 3123 2736
rect 2757 2701 2789 2703
rect 2874 2669 2909 2670
rect 2853 2662 2909 2669
rect 3086 2668 3123 2703
rect 4073 2717 4107 2923
rect 4520 2903 4552 2931
rect 6185 2956 6213 2988
rect 6506 2956 6537 3096
rect 7426 3080 7461 3096
rect 7426 3060 7433 3080
rect 7453 3060 7461 3080
rect 7426 3052 7461 3060
rect 6185 2925 6537 2956
rect 6982 2987 7014 2994
rect 6982 2967 6989 2987
rect 7010 2967 7014 2987
rect 4140 2895 4552 2903
rect 4140 2869 4146 2895
rect 4172 2869 4552 2895
rect 4140 2867 4552 2869
rect 4142 2866 4182 2867
rect 4520 2802 4552 2867
rect 6982 2902 7014 2967
rect 7352 2902 7392 2903
rect 6982 2900 7394 2902
rect 6982 2874 7362 2900
rect 7388 2874 7394 2900
rect 6982 2866 7394 2874
rect 6416 2851 6448 2852
rect 6413 2846 6448 2851
rect 6413 2826 6420 2846
rect 6440 2826 6448 2846
rect 6413 2818 6448 2826
rect 4520 2782 4524 2802
rect 4545 2782 4552 2802
rect 4520 2775 4552 2782
rect 5969 2753 6001 2760
rect 5969 2733 5976 2753
rect 5997 2733 6001 2753
rect 4073 2709 4108 2717
rect 4073 2689 4081 2709
rect 4101 2689 4108 2709
rect 4073 2684 4108 2689
rect 4073 2683 4105 2684
rect 2853 2642 2882 2662
rect 2902 2642 2909 2662
rect 2853 2637 2909 2642
rect 3081 2666 3128 2668
rect 3081 2640 3093 2666
rect 3118 2640 3128 2666
rect 2357 2589 2395 2595
rect 2357 2569 2367 2589
rect 2387 2569 2395 2589
rect 2357 2567 2395 2569
rect 893 2534 1308 2563
rect 2360 2561 2395 2567
rect 893 2533 1302 2534
rect 1916 2496 1948 2503
rect 1916 2476 1923 2496
rect 1944 2476 1948 2496
rect 1916 2411 1948 2476
rect 2286 2411 2326 2412
rect 1916 2409 2328 2411
rect 1916 2383 2296 2409
rect 2322 2383 2328 2409
rect 1916 2375 2328 2383
rect 1916 2347 1948 2375
rect 2361 2355 2395 2561
rect 2853 2431 2887 2637
rect 3081 2634 3128 2640
rect 3300 2665 3332 2672
rect 3300 2645 3306 2665
rect 3327 2645 3332 2665
rect 3300 2617 3332 2645
rect 2920 2609 3332 2617
rect 2920 2583 2926 2609
rect 2952 2583 3332 2609
rect 2920 2581 3332 2583
rect 2922 2580 2962 2581
rect 3300 2516 3332 2581
rect 5969 2668 6001 2733
rect 6339 2668 6379 2669
rect 5969 2666 6381 2668
rect 5969 2640 6349 2666
rect 6375 2640 6381 2666
rect 5969 2632 6381 2640
rect 5969 2604 6001 2632
rect 5969 2584 5974 2604
rect 5995 2584 6001 2604
rect 5969 2577 6001 2584
rect 6169 2604 6219 2613
rect 6414 2612 6448 2818
rect 6982 2838 7014 2866
rect 6982 2818 6987 2838
rect 7008 2818 7014 2838
rect 7187 2840 7229 2849
rect 7427 2846 7461 3052
rect 7187 2826 7197 2840
rect 6982 2811 7014 2818
rect 7186 2820 7197 2826
rect 7221 2820 7229 2840
rect 7186 2809 7229 2820
rect 7405 2841 7461 2846
rect 7405 2821 7412 2841
rect 7432 2821 7461 2841
rect 7405 2814 7461 2821
rect 7405 2813 7440 2814
rect 7186 2779 7226 2809
rect 7076 2771 7112 2775
rect 7076 2752 7084 2771
rect 7104 2752 7112 2771
rect 7076 2749 7112 2752
rect 7186 2774 7533 2779
rect 7077 2721 7111 2749
rect 7186 2748 7505 2774
rect 7524 2748 7533 2774
rect 7186 2744 7533 2748
rect 6169 2583 6181 2604
rect 6203 2583 6219 2604
rect 6169 2575 6219 2583
rect 6392 2607 6448 2612
rect 6392 2587 6399 2607
rect 6419 2587 6448 2607
rect 6392 2580 6448 2587
rect 6549 2693 7112 2721
rect 6392 2579 6427 2580
rect 3300 2496 3304 2516
rect 3325 2496 3332 2516
rect 6174 2542 6215 2575
rect 6549 2542 6589 2693
rect 7638 2574 7673 3168
rect 8038 2715 8070 4368
rect 9209 4217 9249 4368
rect 9583 4335 9624 4368
rect 12652 4344 12684 4409
rect 13022 4344 13062 4345
rect 12652 4342 13064 4344
rect 9371 4330 9406 4331
rect 8686 4189 9249 4217
rect 9350 4323 9406 4330
rect 9350 4303 9379 4323
rect 9399 4303 9406 4323
rect 9350 4298 9406 4303
rect 9579 4327 9629 4335
rect 9579 4306 9595 4327
rect 9617 4306 9629 4327
rect 8265 4162 8612 4166
rect 8265 4136 8274 4162
rect 8293 4136 8612 4162
rect 8687 4161 8721 4189
rect 8265 4131 8612 4136
rect 8686 4158 8722 4161
rect 8686 4139 8694 4158
rect 8714 4139 8722 4158
rect 8686 4135 8722 4139
rect 8572 4101 8612 4131
rect 8358 4096 8393 4097
rect 8337 4089 8393 4096
rect 8337 4069 8366 4089
rect 8386 4069 8393 4089
rect 8337 4064 8393 4069
rect 8569 4090 8612 4101
rect 8569 4070 8577 4090
rect 8601 4084 8612 4090
rect 8784 4092 8816 4099
rect 8601 4070 8611 4084
rect 8337 3858 8371 4064
rect 8569 4061 8611 4070
rect 8784 4072 8790 4092
rect 8811 4072 8816 4092
rect 8784 4044 8816 4072
rect 9350 4092 9384 4298
rect 9579 4297 9629 4306
rect 9797 4326 9829 4333
rect 9797 4306 9803 4326
rect 9824 4306 9829 4326
rect 9797 4278 9829 4306
rect 9417 4270 9829 4278
rect 12652 4316 13032 4342
rect 13058 4316 13064 4342
rect 12652 4308 13064 4316
rect 12652 4280 12684 4308
rect 11792 4276 11824 4277
rect 9417 4244 9423 4270
rect 9449 4244 9829 4270
rect 9417 4242 9829 4244
rect 11789 4271 11824 4276
rect 11789 4251 11796 4271
rect 11816 4251 11824 4271
rect 12652 4260 12657 4280
rect 12678 4260 12684 4280
rect 12652 4253 12684 4260
rect 12857 4282 12906 4292
rect 13097 4288 13131 4494
rect 13419 4431 13453 4637
rect 13644 4633 13693 4643
rect 13866 4665 13898 4672
rect 13866 4645 13872 4665
rect 13893 4645 13898 4665
rect 14726 4654 14734 4674
rect 14754 4654 14761 4674
rect 14726 4649 14761 4654
rect 14726 4648 14758 4649
rect 13866 4617 13898 4645
rect 13486 4609 13898 4617
rect 13486 4583 13492 4609
rect 13518 4583 13898 4609
rect 13486 4581 13898 4583
rect 13488 4580 13528 4581
rect 13866 4516 13898 4581
rect 16622 4633 16654 4698
rect 16992 4633 17032 4634
rect 16622 4631 17034 4633
rect 16622 4605 17002 4631
rect 17028 4605 17034 4631
rect 16622 4597 17034 4605
rect 16622 4569 16654 4597
rect 16622 4549 16627 4569
rect 16648 4549 16654 4569
rect 16622 4542 16654 4549
rect 16822 4569 16872 4578
rect 17067 4577 17101 4783
rect 17635 4803 17667 4831
rect 17635 4783 17640 4803
rect 17661 4783 17667 4803
rect 17840 4805 17882 4814
rect 18080 4811 18114 5017
rect 17840 4791 17850 4805
rect 17635 4776 17667 4783
rect 17839 4785 17850 4791
rect 17874 4785 17882 4805
rect 17839 4774 17882 4785
rect 18058 4806 18114 4811
rect 18058 4786 18065 4806
rect 18085 4786 18114 4806
rect 18058 4779 18114 4786
rect 18058 4778 18093 4779
rect 17839 4744 17879 4774
rect 17729 4736 17765 4740
rect 17729 4717 17737 4736
rect 17757 4717 17765 4736
rect 17729 4714 17765 4717
rect 17839 4739 18186 4744
rect 17730 4686 17764 4714
rect 17839 4713 18158 4739
rect 18177 4713 18186 4739
rect 17839 4709 18186 4713
rect 16822 4548 16834 4569
rect 16856 4548 16872 4569
rect 16822 4540 16872 4548
rect 17045 4572 17101 4577
rect 17045 4552 17052 4572
rect 17072 4552 17101 4572
rect 17045 4545 17101 4552
rect 17202 4658 17765 4686
rect 17045 4544 17080 4545
rect 13866 4496 13870 4516
rect 13891 4496 13898 4516
rect 13866 4489 13898 4496
rect 16827 4507 16868 4540
rect 17202 4507 17242 4658
rect 18381 4507 18413 6160
rect 18778 5707 18813 6301
rect 19862 6182 19902 6333
rect 20236 6300 20277 6333
rect 20024 6295 20059 6296
rect 19339 6154 19902 6182
rect 20003 6288 20059 6295
rect 20003 6268 20032 6288
rect 20052 6268 20059 6288
rect 20003 6263 20059 6268
rect 20232 6292 20282 6300
rect 20232 6271 20248 6292
rect 20270 6271 20282 6292
rect 18918 6127 19265 6131
rect 18918 6101 18927 6127
rect 18946 6101 19265 6127
rect 19340 6126 19374 6154
rect 18918 6096 19265 6101
rect 19339 6123 19375 6126
rect 19339 6104 19347 6123
rect 19367 6104 19375 6123
rect 19339 6100 19375 6104
rect 19225 6066 19265 6096
rect 19011 6061 19046 6062
rect 18990 6054 19046 6061
rect 18990 6034 19019 6054
rect 19039 6034 19046 6054
rect 18990 6029 19046 6034
rect 19222 6055 19265 6066
rect 19222 6035 19230 6055
rect 19254 6049 19265 6055
rect 19437 6057 19469 6064
rect 19254 6035 19264 6049
rect 18990 5823 19024 6029
rect 19222 6026 19264 6035
rect 19437 6037 19443 6057
rect 19464 6037 19469 6057
rect 19437 6009 19469 6037
rect 20003 6057 20037 6263
rect 20232 6262 20282 6271
rect 20450 6291 20482 6298
rect 20450 6271 20456 6291
rect 20477 6271 20482 6291
rect 20450 6243 20482 6271
rect 20070 6235 20482 6243
rect 20070 6209 20076 6235
rect 20102 6209 20482 6235
rect 20070 6207 20482 6209
rect 20072 6206 20112 6207
rect 20450 6142 20482 6207
rect 20450 6122 20454 6142
rect 20475 6122 20482 6142
rect 20450 6115 20482 6122
rect 20003 6049 20038 6057
rect 20003 6029 20011 6049
rect 20031 6029 20038 6049
rect 20003 6024 20038 6029
rect 20003 6023 20035 6024
rect 19057 6001 19469 6009
rect 19057 5975 19063 6001
rect 19089 5975 19469 6001
rect 19057 5973 19469 5975
rect 19059 5972 19099 5973
rect 19437 5908 19469 5973
rect 19437 5888 19441 5908
rect 19462 5888 19469 5908
rect 19437 5881 19469 5888
rect 19914 5919 20266 5950
rect 18990 5815 19025 5823
rect 18990 5795 18998 5815
rect 19018 5795 19025 5815
rect 18990 5779 19025 5795
rect 19914 5779 19945 5919
rect 20238 5887 20266 5919
rect 20023 5880 20058 5881
rect 18988 5760 19945 5779
rect 20002 5873 20058 5880
rect 20002 5853 20031 5873
rect 20051 5853 20058 5873
rect 20002 5848 20058 5853
rect 20232 5875 20272 5887
rect 20232 5854 20238 5875
rect 20260 5854 20272 5875
rect 20232 5849 20272 5854
rect 20449 5876 20481 5883
rect 20449 5856 20455 5876
rect 20476 5856 20481 5876
rect 18778 5678 19208 5707
rect 18778 5673 18862 5678
rect 18961 5641 18996 5642
rect 18940 5634 18996 5641
rect 18940 5614 18969 5634
rect 18989 5614 18996 5634
rect 18940 5609 18996 5614
rect 19170 5635 19208 5678
rect 19170 5618 19175 5635
rect 19199 5618 19208 5635
rect 18940 5405 18974 5609
rect 19170 5606 19208 5618
rect 19387 5637 19419 5644
rect 19387 5617 19393 5637
rect 19414 5617 19419 5637
rect 19387 5589 19419 5617
rect 20002 5642 20036 5848
rect 20449 5828 20481 5856
rect 20069 5820 20481 5828
rect 20069 5794 20075 5820
rect 20101 5794 20481 5820
rect 20069 5792 20481 5794
rect 20071 5791 20111 5792
rect 20449 5727 20481 5792
rect 20449 5707 20453 5727
rect 20474 5707 20481 5727
rect 20449 5700 20481 5707
rect 20002 5634 20037 5642
rect 20002 5614 20010 5634
rect 20030 5614 20037 5634
rect 20002 5609 20037 5614
rect 20002 5608 20034 5609
rect 19007 5581 19419 5589
rect 19007 5555 19013 5581
rect 19039 5555 19419 5581
rect 19007 5553 19419 5555
rect 19009 5552 19049 5553
rect 19387 5488 19419 5553
rect 19387 5468 19391 5488
rect 19412 5468 19419 5488
rect 19387 5461 19419 5468
rect 18938 5395 18978 5405
rect 18938 5375 18948 5395
rect 18968 5375 18978 5395
rect 19873 5381 20282 5382
rect 18938 5151 18978 5375
rect 19867 5352 20282 5381
rect 19867 5201 19907 5352
rect 20241 5319 20282 5352
rect 20029 5314 20064 5315
rect 19344 5173 19907 5201
rect 20008 5307 20064 5314
rect 20008 5287 20037 5307
rect 20057 5287 20064 5307
rect 20008 5282 20064 5287
rect 20237 5311 20287 5319
rect 20237 5290 20253 5311
rect 20275 5290 20287 5311
rect 18938 5117 19265 5151
rect 19345 5145 19379 5173
rect 19344 5142 19380 5145
rect 19344 5123 19352 5142
rect 19372 5123 19380 5142
rect 19344 5119 19380 5123
rect 18955 5116 19265 5117
rect 19230 5087 19265 5116
rect 19016 5080 19051 5081
rect 18995 5073 19051 5080
rect 18995 5053 19024 5073
rect 19044 5053 19051 5073
rect 18995 5048 19051 5053
rect 19225 5075 19267 5087
rect 19225 5055 19234 5075
rect 19258 5055 19267 5075
rect 18995 4842 19029 5048
rect 19225 5047 19267 5055
rect 19442 5076 19474 5083
rect 19442 5056 19448 5076
rect 19469 5056 19474 5076
rect 19442 5028 19474 5056
rect 20008 5076 20042 5282
rect 20237 5281 20287 5290
rect 20455 5310 20487 5317
rect 20455 5290 20461 5310
rect 20482 5290 20487 5310
rect 20455 5262 20487 5290
rect 20075 5254 20487 5262
rect 20075 5228 20081 5254
rect 20107 5228 20487 5254
rect 20075 5226 20487 5228
rect 20077 5225 20117 5226
rect 20455 5161 20487 5226
rect 20455 5141 20459 5161
rect 20480 5141 20487 5161
rect 20455 5134 20487 5141
rect 20008 5068 20043 5076
rect 20008 5048 20016 5068
rect 20036 5048 20043 5068
rect 20008 5043 20043 5048
rect 20008 5042 20040 5043
rect 19062 5020 19474 5028
rect 19062 4994 19068 5020
rect 19094 4994 19474 5020
rect 19062 4992 19474 4994
rect 19064 4991 19104 4992
rect 19442 4927 19474 4992
rect 19442 4907 19446 4927
rect 19467 4907 19474 4927
rect 19442 4900 19474 4907
rect 19919 4938 20271 4969
rect 18995 4834 19030 4842
rect 18995 4814 19003 4834
rect 19023 4814 19030 4834
rect 18995 4798 19030 4814
rect 19919 4798 19950 4938
rect 20243 4906 20271 4938
rect 20028 4899 20063 4900
rect 18993 4779 19950 4798
rect 20007 4892 20063 4899
rect 20007 4872 20036 4892
rect 20056 4872 20063 4892
rect 20007 4867 20063 4872
rect 20237 4894 20277 4906
rect 20237 4873 20243 4894
rect 20265 4873 20277 4894
rect 20237 4868 20277 4873
rect 20454 4895 20486 4902
rect 20454 4875 20460 4895
rect 20481 4875 20486 4895
rect 18591 4722 18676 4725
rect 18584 4718 18676 4722
rect 18584 4717 18965 4718
rect 18584 4687 18591 4717
rect 18628 4688 18965 4717
rect 18628 4687 18676 4688
rect 18584 4685 18676 4687
rect 18584 4682 18669 4685
rect 18930 4650 18965 4688
rect 20007 4661 20041 4867
rect 20454 4847 20486 4875
rect 20074 4839 20486 4847
rect 20074 4813 20080 4839
rect 20106 4813 20486 4839
rect 20074 4811 20486 4813
rect 20076 4810 20116 4811
rect 20454 4746 20486 4811
rect 20454 4726 20458 4746
rect 20479 4726 20486 4746
rect 20454 4719 20486 4726
rect 20007 4653 20042 4661
rect 18721 4648 18756 4649
rect 16827 4478 17242 4507
rect 18380 4506 18413 4507
rect 18377 4501 18413 4506
rect 18377 4481 18384 4501
rect 18404 4481 18413 4501
rect 16827 4477 17236 4478
rect 18377 4476 18413 4481
rect 18700 4641 18756 4648
rect 18700 4621 18729 4641
rect 18749 4621 18756 4641
rect 18700 4616 18756 4621
rect 18925 4641 18974 4650
rect 18925 4622 18933 4641
rect 18959 4622 18974 4641
rect 18377 4473 18412 4476
rect 13419 4428 13454 4431
rect 12857 4263 12872 4282
rect 12898 4263 12906 4282
rect 12857 4254 12906 4263
rect 13075 4283 13131 4288
rect 13075 4263 13082 4283
rect 13102 4263 13131 4283
rect 13075 4256 13131 4263
rect 13418 4423 13454 4428
rect 14595 4426 15004 4427
rect 13418 4403 13427 4423
rect 13447 4403 13454 4423
rect 13418 4398 13454 4403
rect 13418 4397 13451 4398
rect 14589 4397 15004 4426
rect 13075 4255 13110 4256
rect 11789 4243 11824 4251
rect 9419 4241 9459 4242
rect 9797 4177 9829 4242
rect 9797 4157 9801 4177
rect 9822 4157 9829 4177
rect 9797 4150 9829 4157
rect 11345 4178 11377 4185
rect 11345 4158 11352 4178
rect 11373 4158 11377 4178
rect 11345 4093 11377 4158
rect 11715 4093 11755 4094
rect 9350 4084 9385 4092
rect 9350 4064 9358 4084
rect 9378 4064 9385 4084
rect 9350 4059 9385 4064
rect 11345 4091 11757 4093
rect 11345 4065 11725 4091
rect 11751 4065 11757 4091
rect 9350 4058 9382 4059
rect 8404 4036 8816 4044
rect 8404 4010 8410 4036
rect 8436 4010 8816 4036
rect 8404 4008 8816 4010
rect 8406 4007 8446 4008
rect 8784 3943 8816 4008
rect 11345 4057 11757 4065
rect 11345 4029 11377 4057
rect 11790 4037 11824 4243
rect 12866 4216 12901 4254
rect 13124 4216 13247 4221
rect 12866 4215 13247 4216
rect 12866 4187 13209 4215
rect 13243 4214 13247 4215
rect 13243 4187 13248 4214
rect 12866 4186 13248 4187
rect 13124 4181 13248 4186
rect 11345 4009 11350 4029
rect 11371 4009 11377 4029
rect 11345 4002 11377 4009
rect 11554 4031 11594 4036
rect 11554 4010 11566 4031
rect 11588 4010 11594 4031
rect 11554 3998 11594 4010
rect 11768 4032 11824 4037
rect 11768 4012 11775 4032
rect 11795 4012 11824 4032
rect 11768 4005 11824 4012
rect 11881 4106 12838 4125
rect 11768 4004 11803 4005
rect 8784 3923 8788 3943
rect 8809 3923 8816 3943
rect 8784 3916 8816 3923
rect 9261 3954 9613 3985
rect 8337 3850 8372 3858
rect 8337 3830 8345 3850
rect 8365 3830 8372 3850
rect 8337 3814 8372 3830
rect 9261 3814 9292 3954
rect 9585 3922 9613 3954
rect 11560 3966 11588 3998
rect 11881 3966 11912 4106
rect 12801 4090 12836 4106
rect 12801 4070 12808 4090
rect 12828 4070 12836 4090
rect 12801 4062 12836 4070
rect 11560 3935 11912 3966
rect 12357 3997 12389 4004
rect 12357 3977 12364 3997
rect 12385 3977 12389 3997
rect 9370 3915 9405 3916
rect 8335 3795 9292 3814
rect 9349 3908 9405 3915
rect 9349 3888 9378 3908
rect 9398 3888 9405 3908
rect 9349 3883 9405 3888
rect 9579 3910 9619 3922
rect 9579 3889 9585 3910
rect 9607 3889 9619 3910
rect 9579 3884 9619 3889
rect 9796 3911 9828 3918
rect 9796 3891 9802 3911
rect 9823 3891 9828 3911
rect 8174 3743 8203 3745
rect 8174 3738 8547 3743
rect 8174 3720 8181 3738
rect 8201 3720 8547 3738
rect 8174 3715 8547 3720
rect 8179 3713 8547 3715
rect 8308 3676 8343 3677
rect 8523 3676 8547 3713
rect 8287 3669 8343 3676
rect 8287 3649 8316 3669
rect 8336 3649 8343 3669
rect 8287 3644 8343 3649
rect 8518 3671 8555 3676
rect 8518 3652 8526 3671
rect 8549 3652 8555 3671
rect 8518 3646 8555 3652
rect 8734 3672 8766 3679
rect 8734 3652 8740 3672
rect 8761 3652 8766 3672
rect 8287 3440 8321 3644
rect 8734 3624 8766 3652
rect 9349 3677 9383 3883
rect 9796 3863 9828 3891
rect 9416 3855 9828 3863
rect 12357 3912 12389 3977
rect 12727 3912 12767 3913
rect 12357 3910 12769 3912
rect 12357 3884 12737 3910
rect 12763 3884 12769 3910
rect 12357 3876 12769 3884
rect 11791 3861 11823 3862
rect 9416 3829 9422 3855
rect 9448 3829 9828 3855
rect 9416 3827 9828 3829
rect 11788 3856 11823 3861
rect 11788 3836 11795 3856
rect 11815 3836 11823 3856
rect 11788 3828 11823 3836
rect 9418 3826 9458 3827
rect 9796 3762 9828 3827
rect 9796 3742 9800 3762
rect 9821 3742 9828 3762
rect 9796 3735 9828 3742
rect 11344 3763 11376 3770
rect 11344 3743 11351 3763
rect 11372 3743 11376 3763
rect 11344 3678 11376 3743
rect 11714 3678 11754 3679
rect 9349 3669 9384 3677
rect 9349 3649 9357 3669
rect 9377 3649 9384 3669
rect 9349 3644 9384 3649
rect 11344 3676 11756 3678
rect 11344 3650 11724 3676
rect 11750 3650 11756 3676
rect 9349 3643 9381 3644
rect 8354 3616 8766 3624
rect 8354 3590 8360 3616
rect 8386 3590 8766 3616
rect 8354 3588 8766 3590
rect 8356 3587 8396 3588
rect 8734 3523 8766 3588
rect 11344 3642 11756 3650
rect 11344 3614 11376 3642
rect 11344 3594 11349 3614
rect 11370 3594 11376 3614
rect 11344 3587 11376 3594
rect 11544 3614 11594 3623
rect 11789 3622 11823 3828
rect 12357 3848 12389 3876
rect 12357 3828 12362 3848
rect 12383 3828 12389 3848
rect 12357 3821 12389 3828
rect 12564 3849 12606 3857
rect 12802 3856 12836 4062
rect 12564 3829 12573 3849
rect 12597 3829 12606 3849
rect 12564 3817 12606 3829
rect 12780 3851 12836 3856
rect 12780 3831 12787 3851
rect 12807 3831 12836 3851
rect 12780 3824 12836 3831
rect 12780 3823 12815 3824
rect 12566 3788 12601 3817
rect 12566 3787 12876 3788
rect 12451 3781 12487 3785
rect 12451 3762 12459 3781
rect 12479 3762 12487 3781
rect 12451 3759 12487 3762
rect 12452 3731 12486 3759
rect 12566 3753 12893 3787
rect 11544 3593 11556 3614
rect 11578 3593 11594 3614
rect 11544 3585 11594 3593
rect 11767 3617 11823 3622
rect 11767 3597 11774 3617
rect 11794 3597 11823 3617
rect 11767 3590 11823 3597
rect 11924 3703 12487 3731
rect 11767 3589 11802 3590
rect 8734 3503 8738 3523
rect 8759 3503 8766 3523
rect 11549 3552 11590 3585
rect 11924 3552 11964 3703
rect 11549 3523 11964 3552
rect 12853 3529 12893 3753
rect 11549 3522 11958 3523
rect 8734 3496 8766 3503
rect 12853 3509 12863 3529
rect 12883 3509 12893 3529
rect 12853 3499 12893 3509
rect 8285 3430 8325 3440
rect 8285 3410 8295 3430
rect 8315 3410 8325 3430
rect 12412 3436 12444 3443
rect 9220 3416 9629 3417
rect 8285 3186 8325 3410
rect 9214 3387 9629 3416
rect 9214 3236 9254 3387
rect 9588 3354 9629 3387
rect 12412 3416 12419 3436
rect 12440 3416 12444 3436
rect 9376 3349 9411 3350
rect 8691 3208 9254 3236
rect 9355 3342 9411 3349
rect 9355 3322 9384 3342
rect 9404 3322 9411 3342
rect 9355 3317 9411 3322
rect 9584 3346 9634 3354
rect 9584 3325 9600 3346
rect 9622 3325 9634 3346
rect 8285 3152 8612 3186
rect 8692 3180 8726 3208
rect 8691 3177 8727 3180
rect 8691 3158 8699 3177
rect 8719 3158 8727 3177
rect 8691 3154 8727 3158
rect 8302 3151 8612 3152
rect 8577 3122 8612 3151
rect 8363 3115 8398 3116
rect 8342 3108 8398 3115
rect 8342 3088 8371 3108
rect 8391 3088 8398 3108
rect 8342 3083 8398 3088
rect 8572 3110 8614 3122
rect 8572 3090 8581 3110
rect 8605 3090 8614 3110
rect 8342 2877 8376 3083
rect 8572 3082 8614 3090
rect 8789 3111 8821 3118
rect 8789 3091 8795 3111
rect 8816 3091 8821 3111
rect 8789 3063 8821 3091
rect 9355 3111 9389 3317
rect 9584 3316 9634 3325
rect 9802 3345 9834 3352
rect 9802 3325 9808 3345
rect 9829 3325 9834 3345
rect 9802 3297 9834 3325
rect 9422 3289 9834 3297
rect 12412 3351 12444 3416
rect 12782 3351 12822 3352
rect 12412 3349 12824 3351
rect 12412 3323 12792 3349
rect 12818 3323 12824 3349
rect 12412 3315 12824 3323
rect 11797 3295 11829 3296
rect 9422 3263 9428 3289
rect 9454 3263 9834 3289
rect 9422 3261 9834 3263
rect 11794 3290 11829 3295
rect 11794 3270 11801 3290
rect 11821 3270 11829 3290
rect 11794 3262 11829 3270
rect 9424 3260 9464 3261
rect 9802 3196 9834 3261
rect 9802 3176 9806 3196
rect 9827 3176 9834 3196
rect 9802 3169 9834 3176
rect 11350 3197 11382 3204
rect 11350 3177 11357 3197
rect 11378 3177 11382 3197
rect 11350 3112 11382 3177
rect 11720 3112 11760 3113
rect 9355 3103 9390 3111
rect 9355 3083 9363 3103
rect 9383 3083 9390 3103
rect 9355 3078 9390 3083
rect 11350 3110 11762 3112
rect 11350 3084 11730 3110
rect 11756 3084 11762 3110
rect 9355 3077 9387 3078
rect 8409 3055 8821 3063
rect 8409 3029 8415 3055
rect 8441 3029 8821 3055
rect 8409 3027 8821 3029
rect 8411 3026 8451 3027
rect 8789 2962 8821 3027
rect 11350 3076 11762 3084
rect 11350 3048 11382 3076
rect 11795 3056 11829 3262
rect 12412 3287 12444 3315
rect 12412 3267 12417 3287
rect 12438 3267 12444 3287
rect 12412 3260 12444 3267
rect 12623 3286 12661 3298
rect 12857 3295 12891 3499
rect 12623 3269 12632 3286
rect 12656 3269 12661 3286
rect 12623 3226 12661 3269
rect 12835 3290 12891 3295
rect 12835 3270 12842 3290
rect 12862 3270 12891 3290
rect 12835 3263 12891 3270
rect 12835 3262 12870 3263
rect 12969 3226 13053 3231
rect 12623 3197 13053 3226
rect 11350 3028 11355 3048
rect 11376 3028 11382 3048
rect 11350 3021 11382 3028
rect 11559 3050 11599 3055
rect 11559 3029 11571 3050
rect 11593 3029 11599 3050
rect 11559 3017 11599 3029
rect 11773 3051 11829 3056
rect 11773 3031 11780 3051
rect 11800 3031 11829 3051
rect 11773 3024 11829 3031
rect 11886 3125 12843 3144
rect 11773 3023 11808 3024
rect 8789 2942 8793 2962
rect 8814 2942 8821 2962
rect 8789 2935 8821 2942
rect 9266 2973 9618 3004
rect 8342 2869 8377 2877
rect 8342 2849 8350 2869
rect 8370 2849 8377 2869
rect 8342 2833 8377 2849
rect 9266 2833 9297 2973
rect 9590 2941 9618 2973
rect 11565 2985 11593 3017
rect 11886 2985 11917 3125
rect 12806 3109 12841 3125
rect 12806 3089 12813 3109
rect 12833 3089 12841 3109
rect 12806 3081 12841 3089
rect 11565 2954 11917 2985
rect 12362 3016 12394 3023
rect 12362 2996 12369 3016
rect 12390 2996 12394 3016
rect 9375 2934 9410 2935
rect 8340 2814 9297 2833
rect 9354 2927 9410 2934
rect 9354 2907 9383 2927
rect 9403 2907 9410 2927
rect 9354 2902 9410 2907
rect 9584 2929 9624 2941
rect 9584 2908 9590 2929
rect 9612 2908 9624 2929
rect 9584 2903 9624 2908
rect 9801 2930 9833 2937
rect 9801 2910 9807 2930
rect 9828 2910 9833 2930
rect 8034 2682 8404 2715
rect 8038 2680 8070 2682
rect 8155 2648 8190 2649
rect 8134 2641 8190 2648
rect 8367 2647 8404 2682
rect 9354 2696 9388 2902
rect 9801 2882 9833 2910
rect 9421 2874 9833 2882
rect 12362 2931 12394 2996
rect 12732 2931 12772 2932
rect 12362 2929 12774 2931
rect 12362 2903 12742 2929
rect 12768 2903 12774 2929
rect 12362 2895 12774 2903
rect 11796 2880 11828 2881
rect 9421 2848 9427 2874
rect 9453 2848 9833 2874
rect 9421 2846 9833 2848
rect 11793 2875 11828 2880
rect 11793 2855 11800 2875
rect 11820 2855 11828 2875
rect 11793 2847 11828 2855
rect 9423 2845 9463 2846
rect 9801 2781 9833 2846
rect 9801 2761 9805 2781
rect 9826 2761 9833 2781
rect 9801 2754 9833 2761
rect 11349 2782 11381 2789
rect 11349 2762 11356 2782
rect 11377 2762 11381 2782
rect 11349 2697 11381 2762
rect 11719 2697 11759 2698
rect 9354 2688 9389 2696
rect 9354 2668 9362 2688
rect 9382 2668 9389 2688
rect 9354 2663 9389 2668
rect 11349 2695 11761 2697
rect 11349 2669 11729 2695
rect 11755 2669 11761 2695
rect 9354 2662 9386 2663
rect 11349 2661 11761 2669
rect 8134 2621 8163 2641
rect 8183 2621 8190 2641
rect 8134 2616 8190 2621
rect 8362 2645 8409 2647
rect 8362 2619 8374 2645
rect 8399 2619 8409 2645
rect 7638 2568 7676 2574
rect 7638 2548 7648 2568
rect 7668 2548 7676 2568
rect 7638 2546 7676 2548
rect 6174 2513 6589 2542
rect 7641 2540 7676 2546
rect 6174 2512 6583 2513
rect 3300 2489 3332 2496
rect 7197 2475 7229 2482
rect 3946 2458 4355 2459
rect 2853 2425 2888 2431
rect 3940 2429 4355 2458
rect 2853 2423 2891 2425
rect 2853 2403 2861 2423
rect 2881 2403 2891 2423
rect 2853 2397 2891 2403
rect 1916 2327 1921 2347
rect 1942 2327 1948 2347
rect 1916 2320 1948 2327
rect 2125 2348 2164 2354
rect 2125 2329 2136 2348
rect 2159 2329 2164 2348
rect 2125 2316 2164 2329
rect 2339 2350 2395 2355
rect 2339 2330 2346 2350
rect 2366 2330 2395 2350
rect 2339 2323 2395 2330
rect 2339 2322 2374 2323
rect 1143 2308 1175 2309
rect 1140 2303 1175 2308
rect 1140 2283 1147 2303
rect 1167 2283 1175 2303
rect 1140 2275 1175 2283
rect 696 2210 728 2217
rect 696 2190 703 2210
rect 724 2190 728 2210
rect 696 2125 728 2190
rect 1066 2125 1106 2126
rect 696 2123 1108 2125
rect 696 2097 1076 2123
rect 1102 2097 1108 2123
rect 696 2089 1108 2097
rect 696 2061 728 2089
rect 1141 2069 1175 2275
rect 2132 2285 2162 2316
rect 2442 2285 2479 2291
rect 2132 2280 2479 2285
rect 2132 2261 2448 2280
rect 2471 2261 2479 2280
rect 2132 2255 2479 2261
rect 2442 2250 2479 2255
rect 696 2041 701 2061
rect 722 2041 728 2061
rect 696 2034 728 2041
rect 905 2063 945 2068
rect 905 2042 917 2063
rect 939 2042 945 2063
rect 905 2030 945 2042
rect 1119 2064 1175 2069
rect 1119 2044 1126 2064
rect 1146 2044 1175 2064
rect 1119 2037 1175 2044
rect 1232 2138 2189 2157
rect 1119 2036 1154 2037
rect 911 1998 939 2030
rect 1232 1998 1263 2138
rect 2152 2122 2187 2138
rect 2152 2102 2159 2122
rect 2179 2102 2187 2122
rect 2152 2094 2187 2102
rect 911 1967 1263 1998
rect 1708 2029 1740 2036
rect 1708 2009 1715 2029
rect 1736 2009 1740 2029
rect 1708 1944 1740 2009
rect 2078 1944 2118 1945
rect 1708 1942 2120 1944
rect 1708 1916 2088 1942
rect 2114 1916 2120 1942
rect 1708 1908 2120 1916
rect 1142 1893 1174 1894
rect 1139 1888 1174 1893
rect 1139 1868 1146 1888
rect 1166 1868 1174 1888
rect 1139 1860 1174 1868
rect 695 1795 727 1802
rect 695 1775 702 1795
rect 723 1775 727 1795
rect 695 1710 727 1775
rect 1065 1710 1105 1711
rect 695 1708 1107 1710
rect 695 1682 1075 1708
rect 1101 1682 1107 1708
rect 695 1674 1107 1682
rect 695 1646 727 1674
rect 695 1626 700 1646
rect 721 1626 727 1646
rect 695 1619 727 1626
rect 895 1646 945 1655
rect 1140 1654 1174 1860
rect 1708 1880 1740 1908
rect 1708 1860 1713 1880
rect 1734 1860 1740 1880
rect 1708 1853 1740 1860
rect 1915 1881 1957 1889
rect 2153 1888 2187 2094
rect 1915 1861 1924 1881
rect 1948 1861 1957 1881
rect 1915 1849 1957 1861
rect 2131 1883 2187 1888
rect 2131 1863 2138 1883
rect 2158 1863 2187 1883
rect 2131 1856 2187 1863
rect 2131 1855 2166 1856
rect 1917 1820 1952 1849
rect 1917 1819 2227 1820
rect 1802 1813 1838 1817
rect 1802 1794 1810 1813
rect 1830 1794 1838 1813
rect 1802 1791 1838 1794
rect 1803 1763 1837 1791
rect 1917 1785 2244 1819
rect 895 1625 907 1646
rect 929 1625 945 1646
rect 895 1617 945 1625
rect 1118 1649 1174 1654
rect 1118 1629 1125 1649
rect 1145 1629 1174 1649
rect 1118 1622 1174 1629
rect 1275 1735 1838 1763
rect 1118 1621 1153 1622
rect 900 1584 941 1617
rect 1275 1584 1315 1735
rect 900 1555 1315 1584
rect 2204 1561 2244 1785
rect 2856 1803 2891 2397
rect 3940 2278 3980 2429
rect 4314 2396 4355 2429
rect 7197 2455 7204 2475
rect 7225 2455 7229 2475
rect 4102 2391 4137 2392
rect 3417 2250 3980 2278
rect 4081 2384 4137 2391
rect 4081 2364 4110 2384
rect 4130 2364 4137 2384
rect 4081 2359 4137 2364
rect 4310 2388 4360 2396
rect 4310 2367 4326 2388
rect 4348 2367 4360 2388
rect 2996 2223 3343 2227
rect 2996 2197 3005 2223
rect 3024 2197 3343 2223
rect 3418 2222 3452 2250
rect 2996 2192 3343 2197
rect 3417 2219 3453 2222
rect 3417 2200 3425 2219
rect 3445 2200 3453 2219
rect 3417 2196 3453 2200
rect 3303 2162 3343 2192
rect 3089 2157 3124 2158
rect 3068 2150 3124 2157
rect 3068 2130 3097 2150
rect 3117 2130 3124 2150
rect 3068 2125 3124 2130
rect 3300 2151 3343 2162
rect 3300 2131 3308 2151
rect 3332 2145 3343 2151
rect 3515 2153 3547 2160
rect 3332 2131 3342 2145
rect 3068 1919 3102 2125
rect 3300 2122 3342 2131
rect 3515 2133 3521 2153
rect 3542 2133 3547 2153
rect 3515 2105 3547 2133
rect 4081 2153 4115 2359
rect 4310 2358 4360 2367
rect 4528 2387 4560 2394
rect 4528 2367 4534 2387
rect 4555 2367 4560 2387
rect 4528 2339 4560 2367
rect 4148 2331 4560 2339
rect 4148 2305 4154 2331
rect 4180 2305 4560 2331
rect 4148 2303 4560 2305
rect 4150 2302 4190 2303
rect 4528 2238 4560 2303
rect 7197 2390 7229 2455
rect 7567 2390 7607 2391
rect 7197 2388 7609 2390
rect 7197 2362 7577 2388
rect 7603 2362 7609 2388
rect 7197 2354 7609 2362
rect 7197 2326 7229 2354
rect 7642 2334 7676 2540
rect 8134 2410 8168 2616
rect 8362 2613 8409 2619
rect 8581 2644 8613 2651
rect 8581 2624 8587 2644
rect 8608 2624 8613 2644
rect 8581 2596 8613 2624
rect 11349 2633 11381 2661
rect 11349 2613 11354 2633
rect 11375 2613 11381 2633
rect 11349 2606 11381 2613
rect 11549 2633 11599 2642
rect 11794 2641 11828 2847
rect 12362 2867 12394 2895
rect 12362 2847 12367 2867
rect 12388 2847 12394 2867
rect 12567 2869 12609 2878
rect 12807 2875 12841 3081
rect 12567 2855 12577 2869
rect 12362 2840 12394 2847
rect 12566 2849 12577 2855
rect 12601 2849 12609 2869
rect 12566 2838 12609 2849
rect 12785 2870 12841 2875
rect 12785 2850 12792 2870
rect 12812 2850 12841 2870
rect 12785 2843 12841 2850
rect 12785 2842 12820 2843
rect 12566 2808 12606 2838
rect 12456 2800 12492 2804
rect 12456 2781 12464 2800
rect 12484 2781 12492 2800
rect 12456 2778 12492 2781
rect 12566 2803 12913 2808
rect 12457 2750 12491 2778
rect 12566 2777 12885 2803
rect 12904 2777 12913 2803
rect 12566 2773 12913 2777
rect 11549 2612 11561 2633
rect 11583 2612 11599 2633
rect 11549 2604 11599 2612
rect 11772 2636 11828 2641
rect 11772 2616 11779 2636
rect 11799 2616 11828 2636
rect 11772 2609 11828 2616
rect 11929 2722 12492 2750
rect 11772 2608 11807 2609
rect 8201 2588 8613 2596
rect 8201 2562 8207 2588
rect 8233 2562 8613 2588
rect 8201 2560 8613 2562
rect 8203 2559 8243 2560
rect 8581 2495 8613 2560
rect 11554 2571 11595 2604
rect 11929 2571 11969 2722
rect 13018 2603 13053 3197
rect 13418 2744 13450 4397
rect 14589 4246 14629 4397
rect 14963 4364 15004 4397
rect 17933 4408 17965 4415
rect 17933 4388 17940 4408
rect 17961 4388 17965 4408
rect 14751 4359 14786 4360
rect 14066 4218 14629 4246
rect 14730 4352 14786 4359
rect 14730 4332 14759 4352
rect 14779 4332 14786 4352
rect 14730 4327 14786 4332
rect 14959 4356 15009 4364
rect 14959 4335 14975 4356
rect 14997 4335 15009 4356
rect 13645 4191 13992 4195
rect 13645 4165 13654 4191
rect 13673 4165 13992 4191
rect 14067 4190 14101 4218
rect 13645 4160 13992 4165
rect 14066 4187 14102 4190
rect 14066 4168 14074 4187
rect 14094 4168 14102 4187
rect 14066 4164 14102 4168
rect 13952 4130 13992 4160
rect 13738 4125 13773 4126
rect 13717 4118 13773 4125
rect 13717 4098 13746 4118
rect 13766 4098 13773 4118
rect 13717 4093 13773 4098
rect 13949 4119 13992 4130
rect 13949 4099 13957 4119
rect 13981 4113 13992 4119
rect 14164 4121 14196 4128
rect 13981 4099 13991 4113
rect 13717 3887 13751 4093
rect 13949 4090 13991 4099
rect 14164 4101 14170 4121
rect 14191 4101 14196 4121
rect 14164 4073 14196 4101
rect 14730 4121 14764 4327
rect 14959 4326 15009 4335
rect 15177 4355 15209 4362
rect 15177 4335 15183 4355
rect 15204 4335 15209 4355
rect 15177 4307 15209 4335
rect 14797 4299 15209 4307
rect 14797 4273 14803 4299
rect 14829 4273 15209 4299
rect 14797 4271 15209 4273
rect 14799 4270 14839 4271
rect 15177 4206 15209 4271
rect 17933 4323 17965 4388
rect 18303 4323 18343 4324
rect 17933 4321 18345 4323
rect 17933 4295 18313 4321
rect 18339 4295 18345 4321
rect 17933 4287 18345 4295
rect 17933 4259 17965 4287
rect 17073 4255 17105 4256
rect 17070 4250 17105 4255
rect 17070 4230 17077 4250
rect 17097 4230 17105 4250
rect 17933 4239 17938 4259
rect 17959 4239 17965 4259
rect 17933 4232 17965 4239
rect 18138 4261 18187 4271
rect 18378 4267 18412 4473
rect 18700 4410 18734 4616
rect 18925 4612 18974 4622
rect 19147 4644 19179 4651
rect 19147 4624 19153 4644
rect 19174 4624 19179 4644
rect 20007 4633 20015 4653
rect 20035 4633 20042 4653
rect 20007 4628 20042 4633
rect 20007 4627 20039 4628
rect 19147 4596 19179 4624
rect 18767 4588 19179 4596
rect 18767 4562 18773 4588
rect 18799 4562 19179 4588
rect 18767 4560 19179 4562
rect 18769 4559 18809 4560
rect 19147 4495 19179 4560
rect 19147 4475 19151 4495
rect 19172 4475 19179 4495
rect 19147 4468 19179 4475
rect 18700 4407 18735 4410
rect 18138 4242 18153 4261
rect 18179 4242 18187 4261
rect 18138 4233 18187 4242
rect 18356 4262 18412 4267
rect 18356 4242 18363 4262
rect 18383 4242 18412 4262
rect 18356 4235 18412 4242
rect 18699 4402 18735 4407
rect 19876 4405 20285 4406
rect 18699 4382 18708 4402
rect 18728 4382 18735 4402
rect 18699 4377 18735 4382
rect 18699 4376 18732 4377
rect 19870 4376 20285 4405
rect 18356 4234 18391 4235
rect 17070 4222 17105 4230
rect 15177 4186 15181 4206
rect 15202 4186 15209 4206
rect 15177 4179 15209 4186
rect 16626 4157 16658 4164
rect 16626 4137 16633 4157
rect 16654 4137 16658 4157
rect 14730 4113 14765 4121
rect 14730 4093 14738 4113
rect 14758 4093 14765 4113
rect 14730 4088 14765 4093
rect 14730 4087 14762 4088
rect 13784 4065 14196 4073
rect 13784 4039 13790 4065
rect 13816 4039 14196 4065
rect 13784 4037 14196 4039
rect 13786 4036 13826 4037
rect 14164 3972 14196 4037
rect 16626 4072 16658 4137
rect 16996 4072 17036 4073
rect 16626 4070 17038 4072
rect 16626 4044 17006 4070
rect 17032 4044 17038 4070
rect 16626 4036 17038 4044
rect 14164 3952 14168 3972
rect 14189 3952 14196 3972
rect 14164 3945 14196 3952
rect 14641 3983 14993 4014
rect 13717 3879 13752 3887
rect 13717 3859 13725 3879
rect 13745 3859 13752 3879
rect 13717 3843 13752 3859
rect 14641 3843 14672 3983
rect 14965 3951 14993 3983
rect 16626 4008 16658 4036
rect 17071 4016 17105 4222
rect 18147 4195 18182 4233
rect 18405 4195 18528 4200
rect 18147 4194 18528 4195
rect 18147 4166 18490 4194
rect 18524 4193 18528 4194
rect 18524 4166 18529 4193
rect 18147 4165 18529 4166
rect 18405 4160 18529 4165
rect 16626 3988 16631 4008
rect 16652 3988 16658 4008
rect 16626 3981 16658 3988
rect 16835 4010 16875 4015
rect 16835 3989 16847 4010
rect 16869 3989 16875 4010
rect 16835 3977 16875 3989
rect 17049 4011 17105 4016
rect 17049 3991 17056 4011
rect 17076 3991 17105 4011
rect 17049 3984 17105 3991
rect 17162 4085 18119 4104
rect 17049 3983 17084 3984
rect 14750 3944 14785 3945
rect 13715 3824 14672 3843
rect 14729 3937 14785 3944
rect 14729 3917 14758 3937
rect 14778 3917 14785 3937
rect 14729 3912 14785 3917
rect 14959 3939 14999 3951
rect 14959 3918 14965 3939
rect 14987 3918 14999 3939
rect 14959 3913 14999 3918
rect 15176 3940 15208 3947
rect 15176 3920 15182 3940
rect 15203 3920 15208 3940
rect 13554 3772 13583 3774
rect 13554 3767 13927 3772
rect 13554 3749 13561 3767
rect 13581 3749 13927 3767
rect 13554 3744 13927 3749
rect 13559 3742 13927 3744
rect 13688 3705 13723 3706
rect 13903 3705 13927 3742
rect 13667 3698 13723 3705
rect 13667 3678 13696 3698
rect 13716 3678 13723 3698
rect 13667 3673 13723 3678
rect 13898 3700 13935 3705
rect 13898 3681 13906 3700
rect 13929 3681 13935 3700
rect 13898 3675 13935 3681
rect 14114 3701 14146 3708
rect 14114 3681 14120 3701
rect 14141 3681 14146 3701
rect 13667 3469 13701 3673
rect 14114 3653 14146 3681
rect 14729 3706 14763 3912
rect 15176 3892 15208 3920
rect 16841 3945 16869 3977
rect 17162 3945 17193 4085
rect 18082 4069 18117 4085
rect 18082 4049 18089 4069
rect 18109 4049 18117 4069
rect 18082 4041 18117 4049
rect 16841 3914 17193 3945
rect 17638 3976 17670 3983
rect 17638 3956 17645 3976
rect 17666 3956 17670 3976
rect 14796 3884 15208 3892
rect 14796 3858 14802 3884
rect 14828 3858 15208 3884
rect 14796 3856 15208 3858
rect 14798 3855 14838 3856
rect 15176 3791 15208 3856
rect 17638 3891 17670 3956
rect 18008 3891 18048 3892
rect 17638 3889 18050 3891
rect 17638 3863 18018 3889
rect 18044 3863 18050 3889
rect 17638 3855 18050 3863
rect 17072 3840 17104 3841
rect 17069 3835 17104 3840
rect 17069 3815 17076 3835
rect 17096 3815 17104 3835
rect 17069 3807 17104 3815
rect 15176 3771 15180 3791
rect 15201 3771 15208 3791
rect 15176 3764 15208 3771
rect 16625 3742 16657 3749
rect 16625 3722 16632 3742
rect 16653 3722 16657 3742
rect 14729 3698 14764 3706
rect 14729 3678 14737 3698
rect 14757 3678 14764 3698
rect 14729 3673 14764 3678
rect 14729 3672 14761 3673
rect 13734 3645 14146 3653
rect 13734 3619 13740 3645
rect 13766 3619 14146 3645
rect 13734 3617 14146 3619
rect 13736 3616 13776 3617
rect 14114 3552 14146 3617
rect 16625 3657 16657 3722
rect 16995 3657 17035 3658
rect 16625 3655 17037 3657
rect 16625 3629 17005 3655
rect 17031 3629 17037 3655
rect 16625 3621 17037 3629
rect 16625 3593 16657 3621
rect 16625 3573 16630 3593
rect 16651 3573 16657 3593
rect 16625 3566 16657 3573
rect 16825 3593 16875 3602
rect 17070 3601 17104 3807
rect 17638 3827 17670 3855
rect 17638 3807 17643 3827
rect 17664 3807 17670 3827
rect 17638 3800 17670 3807
rect 17845 3828 17887 3836
rect 18083 3835 18117 4041
rect 17845 3808 17854 3828
rect 17878 3808 17887 3828
rect 17845 3796 17887 3808
rect 18061 3830 18117 3835
rect 18061 3810 18068 3830
rect 18088 3810 18117 3830
rect 18061 3803 18117 3810
rect 18061 3802 18096 3803
rect 17847 3767 17882 3796
rect 17847 3766 18157 3767
rect 17732 3760 17768 3764
rect 17732 3741 17740 3760
rect 17760 3741 17768 3760
rect 17732 3738 17768 3741
rect 17733 3710 17767 3738
rect 17847 3732 18174 3766
rect 16825 3572 16837 3593
rect 16859 3572 16875 3593
rect 16825 3564 16875 3572
rect 17048 3596 17104 3601
rect 17048 3576 17055 3596
rect 17075 3576 17104 3596
rect 17048 3569 17104 3576
rect 17205 3682 17768 3710
rect 17048 3568 17083 3569
rect 14114 3532 14118 3552
rect 14139 3532 14146 3552
rect 14114 3525 14146 3532
rect 16830 3531 16871 3564
rect 17205 3531 17245 3682
rect 16830 3502 17245 3531
rect 18134 3508 18174 3732
rect 16830 3501 17239 3502
rect 18134 3488 18144 3508
rect 18164 3488 18174 3508
rect 18134 3478 18174 3488
rect 13665 3459 13705 3469
rect 13665 3439 13675 3459
rect 13695 3439 13705 3459
rect 14600 3445 15009 3446
rect 13665 3215 13705 3439
rect 14594 3416 15009 3445
rect 14594 3265 14634 3416
rect 14968 3383 15009 3416
rect 17693 3415 17725 3422
rect 17693 3395 17700 3415
rect 17721 3395 17725 3415
rect 14756 3378 14791 3379
rect 14071 3237 14634 3265
rect 14735 3371 14791 3378
rect 14735 3351 14764 3371
rect 14784 3351 14791 3371
rect 14735 3346 14791 3351
rect 14964 3375 15014 3383
rect 14964 3354 14980 3375
rect 15002 3354 15014 3375
rect 13665 3181 13992 3215
rect 14072 3209 14106 3237
rect 14071 3206 14107 3209
rect 14071 3187 14079 3206
rect 14099 3187 14107 3206
rect 14071 3183 14107 3187
rect 13682 3180 13992 3181
rect 13957 3151 13992 3180
rect 13743 3144 13778 3145
rect 13722 3137 13778 3144
rect 13722 3117 13751 3137
rect 13771 3117 13778 3137
rect 13722 3112 13778 3117
rect 13952 3139 13994 3151
rect 13952 3119 13961 3139
rect 13985 3119 13994 3139
rect 13722 2906 13756 3112
rect 13952 3111 13994 3119
rect 14169 3140 14201 3147
rect 14169 3120 14175 3140
rect 14196 3120 14201 3140
rect 14169 3092 14201 3120
rect 14735 3140 14769 3346
rect 14964 3345 15014 3354
rect 15182 3374 15214 3381
rect 15182 3354 15188 3374
rect 15209 3354 15214 3374
rect 15182 3326 15214 3354
rect 14802 3318 15214 3326
rect 14802 3292 14808 3318
rect 14834 3292 15214 3318
rect 14802 3290 15214 3292
rect 14804 3289 14844 3290
rect 15182 3225 15214 3290
rect 17693 3330 17725 3395
rect 18063 3330 18103 3331
rect 17693 3328 18105 3330
rect 17693 3302 18073 3328
rect 18099 3302 18105 3328
rect 17693 3294 18105 3302
rect 17078 3274 17110 3275
rect 17075 3269 17110 3274
rect 17075 3249 17082 3269
rect 17102 3249 17110 3269
rect 17075 3241 17110 3249
rect 15182 3205 15186 3225
rect 15207 3205 15214 3225
rect 15182 3198 15214 3205
rect 16631 3176 16663 3183
rect 16631 3156 16638 3176
rect 16659 3156 16663 3176
rect 14735 3132 14770 3140
rect 14735 3112 14743 3132
rect 14763 3112 14770 3132
rect 14735 3107 14770 3112
rect 14735 3106 14767 3107
rect 13789 3084 14201 3092
rect 13789 3058 13795 3084
rect 13821 3058 14201 3084
rect 13789 3056 14201 3058
rect 13791 3055 13831 3056
rect 14169 2991 14201 3056
rect 16631 3091 16663 3156
rect 17001 3091 17041 3092
rect 16631 3089 17043 3091
rect 16631 3063 17011 3089
rect 17037 3063 17043 3089
rect 16631 3055 17043 3063
rect 14169 2971 14173 2991
rect 14194 2971 14201 2991
rect 14169 2964 14201 2971
rect 14646 3002 14998 3033
rect 13722 2898 13757 2906
rect 13722 2878 13730 2898
rect 13750 2878 13757 2898
rect 13722 2862 13757 2878
rect 14646 2862 14677 3002
rect 14970 2970 14998 3002
rect 16631 3027 16663 3055
rect 17076 3035 17110 3241
rect 17693 3266 17725 3294
rect 17693 3246 17698 3266
rect 17719 3246 17725 3266
rect 17693 3239 17725 3246
rect 17904 3265 17942 3277
rect 18138 3274 18172 3478
rect 17904 3248 17913 3265
rect 17937 3248 17942 3265
rect 17904 3205 17942 3248
rect 18116 3269 18172 3274
rect 18116 3249 18123 3269
rect 18143 3249 18172 3269
rect 18116 3242 18172 3249
rect 18116 3241 18151 3242
rect 18250 3205 18334 3210
rect 17904 3176 18334 3205
rect 16631 3007 16636 3027
rect 16657 3007 16663 3027
rect 16631 3000 16663 3007
rect 16840 3029 16880 3034
rect 16840 3008 16852 3029
rect 16874 3008 16880 3029
rect 16840 2996 16880 3008
rect 17054 3030 17110 3035
rect 17054 3010 17061 3030
rect 17081 3010 17110 3030
rect 17054 3003 17110 3010
rect 17167 3104 18124 3123
rect 17054 3002 17089 3003
rect 14755 2963 14790 2964
rect 13720 2843 14677 2862
rect 14734 2956 14790 2963
rect 14734 2936 14763 2956
rect 14783 2936 14790 2956
rect 14734 2931 14790 2936
rect 14964 2958 15004 2970
rect 14964 2937 14970 2958
rect 14992 2937 15004 2958
rect 14964 2932 15004 2937
rect 15181 2959 15213 2966
rect 15181 2939 15187 2959
rect 15208 2939 15213 2959
rect 13414 2711 13784 2744
rect 13418 2709 13450 2711
rect 13535 2677 13570 2678
rect 13514 2670 13570 2677
rect 13747 2676 13784 2711
rect 14734 2725 14768 2931
rect 15181 2911 15213 2939
rect 16846 2964 16874 2996
rect 17167 2964 17198 3104
rect 18087 3088 18122 3104
rect 18087 3068 18094 3088
rect 18114 3068 18122 3088
rect 18087 3060 18122 3068
rect 16846 2933 17198 2964
rect 17643 2995 17675 3002
rect 17643 2975 17650 2995
rect 17671 2975 17675 2995
rect 14801 2903 15213 2911
rect 14801 2877 14807 2903
rect 14833 2877 15213 2903
rect 14801 2875 15213 2877
rect 14803 2874 14843 2875
rect 15181 2810 15213 2875
rect 17643 2910 17675 2975
rect 18013 2910 18053 2911
rect 17643 2908 18055 2910
rect 17643 2882 18023 2908
rect 18049 2882 18055 2908
rect 17643 2874 18055 2882
rect 17077 2859 17109 2860
rect 17074 2854 17109 2859
rect 17074 2834 17081 2854
rect 17101 2834 17109 2854
rect 17074 2826 17109 2834
rect 15181 2790 15185 2810
rect 15206 2790 15213 2810
rect 15181 2783 15213 2790
rect 16630 2761 16662 2768
rect 16630 2741 16637 2761
rect 16658 2741 16662 2761
rect 14734 2717 14769 2725
rect 14734 2697 14742 2717
rect 14762 2697 14769 2717
rect 14734 2692 14769 2697
rect 14734 2691 14766 2692
rect 13514 2650 13543 2670
rect 13563 2650 13570 2670
rect 13514 2645 13570 2650
rect 13742 2674 13789 2676
rect 13742 2648 13754 2674
rect 13779 2648 13789 2674
rect 13018 2597 13056 2603
rect 13018 2577 13028 2597
rect 13048 2577 13056 2597
rect 13018 2575 13056 2577
rect 11554 2542 11969 2571
rect 13021 2569 13056 2575
rect 11554 2541 11963 2542
rect 8581 2475 8585 2495
rect 8606 2475 8613 2495
rect 8581 2468 8613 2475
rect 12577 2504 12609 2511
rect 12577 2484 12584 2504
rect 12605 2484 12609 2504
rect 9227 2437 9636 2438
rect 8134 2404 8169 2410
rect 9221 2408 9636 2437
rect 8134 2402 8172 2404
rect 8134 2382 8142 2402
rect 8162 2382 8172 2402
rect 8134 2376 8172 2382
rect 7197 2306 7202 2326
rect 7223 2306 7229 2326
rect 7197 2299 7229 2306
rect 7406 2327 7445 2333
rect 7406 2308 7417 2327
rect 7440 2308 7445 2327
rect 7406 2295 7445 2308
rect 7620 2329 7676 2334
rect 7620 2309 7627 2329
rect 7647 2309 7676 2329
rect 7620 2302 7676 2309
rect 7620 2301 7655 2302
rect 6424 2287 6456 2288
rect 6421 2282 6456 2287
rect 6421 2262 6428 2282
rect 6448 2262 6456 2282
rect 6421 2254 6456 2262
rect 4528 2218 4532 2238
rect 4553 2218 4560 2238
rect 4528 2211 4560 2218
rect 5977 2189 6009 2196
rect 5977 2169 5984 2189
rect 6005 2169 6009 2189
rect 4081 2145 4116 2153
rect 4081 2125 4089 2145
rect 4109 2125 4116 2145
rect 4081 2120 4116 2125
rect 4081 2119 4113 2120
rect 3135 2097 3547 2105
rect 3135 2071 3141 2097
rect 3167 2071 3547 2097
rect 3135 2069 3547 2071
rect 3137 2068 3177 2069
rect 3515 2004 3547 2069
rect 5977 2104 6009 2169
rect 6347 2104 6387 2105
rect 5977 2102 6389 2104
rect 5977 2076 6357 2102
rect 6383 2076 6389 2102
rect 5977 2068 6389 2076
rect 3515 1984 3519 2004
rect 3540 1984 3547 2004
rect 3515 1977 3547 1984
rect 3992 2015 4344 2046
rect 3068 1911 3103 1919
rect 3068 1891 3076 1911
rect 3096 1891 3103 1911
rect 3068 1875 3103 1891
rect 3992 1875 4023 2015
rect 4316 1983 4344 2015
rect 5977 2040 6009 2068
rect 6422 2048 6456 2254
rect 7413 2264 7443 2295
rect 7723 2264 7760 2270
rect 7413 2259 7760 2264
rect 7413 2240 7729 2259
rect 7752 2240 7760 2259
rect 7413 2234 7760 2240
rect 7723 2229 7760 2234
rect 5977 2020 5982 2040
rect 6003 2020 6009 2040
rect 5977 2013 6009 2020
rect 6186 2042 6226 2047
rect 6186 2021 6198 2042
rect 6220 2021 6226 2042
rect 6186 2009 6226 2021
rect 6400 2043 6456 2048
rect 6400 2023 6407 2043
rect 6427 2023 6456 2043
rect 6400 2016 6456 2023
rect 6513 2117 7470 2136
rect 6400 2015 6435 2016
rect 4101 1976 4136 1977
rect 3066 1856 4023 1875
rect 4080 1969 4136 1976
rect 4080 1949 4109 1969
rect 4129 1949 4136 1969
rect 4080 1944 4136 1949
rect 4310 1971 4350 1983
rect 4310 1950 4316 1971
rect 4338 1950 4350 1971
rect 4310 1945 4350 1950
rect 4527 1972 4559 1979
rect 4527 1952 4533 1972
rect 4554 1952 4559 1972
rect 2856 1774 3286 1803
rect 2856 1769 2940 1774
rect 3039 1737 3074 1738
rect 900 1554 1309 1555
rect 2204 1541 2214 1561
rect 2234 1541 2244 1561
rect 2204 1531 2244 1541
rect 3018 1730 3074 1737
rect 3018 1710 3047 1730
rect 3067 1710 3074 1730
rect 3018 1705 3074 1710
rect 3248 1731 3286 1774
rect 3248 1714 3253 1731
rect 3277 1714 3286 1731
rect 1763 1468 1795 1475
rect 1763 1448 1770 1468
rect 1791 1448 1795 1468
rect 1763 1383 1795 1448
rect 2133 1383 2173 1384
rect 1763 1381 2175 1383
rect 1763 1355 2143 1381
rect 2169 1355 2175 1381
rect 1763 1347 2175 1355
rect 1148 1327 1180 1328
rect 1145 1322 1180 1327
rect 1145 1302 1152 1322
rect 1172 1302 1180 1322
rect 1145 1294 1180 1302
rect 701 1229 733 1236
rect 701 1209 708 1229
rect 729 1209 733 1229
rect 701 1144 733 1209
rect 1071 1144 1111 1145
rect 701 1142 1113 1144
rect 701 1116 1081 1142
rect 1107 1116 1113 1142
rect 701 1108 1113 1116
rect 701 1080 733 1108
rect 1146 1088 1180 1294
rect 1763 1319 1795 1347
rect 2208 1327 2242 1531
rect 3018 1501 3052 1705
rect 3248 1702 3286 1714
rect 3465 1733 3497 1740
rect 3465 1713 3471 1733
rect 3492 1713 3497 1733
rect 3465 1685 3497 1713
rect 4080 1738 4114 1944
rect 4527 1924 4559 1952
rect 6192 1977 6220 2009
rect 6513 1977 6544 2117
rect 7433 2101 7468 2117
rect 7433 2081 7440 2101
rect 7460 2081 7468 2101
rect 7433 2073 7468 2081
rect 6192 1946 6544 1977
rect 6989 2008 7021 2015
rect 6989 1988 6996 2008
rect 7017 1988 7021 2008
rect 4147 1916 4559 1924
rect 4147 1890 4153 1916
rect 4179 1890 4559 1916
rect 4147 1888 4559 1890
rect 4149 1887 4189 1888
rect 4527 1823 4559 1888
rect 6989 1923 7021 1988
rect 7359 1923 7399 1924
rect 6989 1921 7401 1923
rect 6989 1895 7369 1921
rect 7395 1895 7401 1921
rect 6989 1887 7401 1895
rect 6423 1872 6455 1873
rect 6420 1867 6455 1872
rect 6420 1847 6427 1867
rect 6447 1847 6455 1867
rect 6420 1839 6455 1847
rect 4527 1803 4531 1823
rect 4552 1803 4559 1823
rect 4527 1796 4559 1803
rect 5976 1774 6008 1781
rect 5976 1754 5983 1774
rect 6004 1754 6008 1774
rect 4080 1730 4115 1738
rect 4080 1710 4088 1730
rect 4108 1710 4115 1730
rect 4080 1705 4115 1710
rect 4080 1704 4112 1705
rect 3085 1677 3497 1685
rect 3085 1651 3091 1677
rect 3117 1651 3497 1677
rect 3085 1649 3497 1651
rect 3087 1648 3127 1649
rect 3465 1584 3497 1649
rect 5976 1689 6008 1754
rect 6346 1689 6386 1690
rect 5976 1687 6388 1689
rect 5976 1661 6356 1687
rect 6382 1661 6388 1687
rect 5976 1653 6388 1661
rect 5976 1625 6008 1653
rect 5976 1605 5981 1625
rect 6002 1605 6008 1625
rect 5976 1598 6008 1605
rect 6176 1625 6226 1634
rect 6421 1633 6455 1839
rect 6989 1859 7021 1887
rect 6989 1839 6994 1859
rect 7015 1839 7021 1859
rect 6989 1832 7021 1839
rect 7196 1860 7238 1868
rect 7434 1867 7468 2073
rect 7196 1840 7205 1860
rect 7229 1840 7238 1860
rect 7196 1828 7238 1840
rect 7412 1862 7468 1867
rect 7412 1842 7419 1862
rect 7439 1842 7468 1862
rect 7412 1835 7468 1842
rect 7412 1834 7447 1835
rect 7198 1799 7233 1828
rect 7198 1798 7508 1799
rect 7083 1792 7119 1796
rect 7083 1773 7091 1792
rect 7111 1773 7119 1792
rect 7083 1770 7119 1773
rect 7084 1742 7118 1770
rect 7198 1764 7525 1798
rect 6176 1604 6188 1625
rect 6210 1604 6226 1625
rect 6176 1596 6226 1604
rect 6399 1628 6455 1633
rect 6399 1608 6406 1628
rect 6426 1608 6455 1628
rect 6399 1601 6455 1608
rect 6556 1714 7119 1742
rect 6399 1600 6434 1601
rect 3465 1564 3469 1584
rect 3490 1564 3497 1584
rect 3465 1557 3497 1564
rect 6181 1563 6222 1596
rect 6556 1563 6596 1714
rect 6181 1534 6596 1563
rect 7485 1540 7525 1764
rect 8137 1782 8172 2376
rect 9221 2257 9261 2408
rect 9595 2375 9636 2408
rect 12577 2419 12609 2484
rect 12947 2419 12987 2420
rect 12577 2417 12989 2419
rect 12577 2391 12957 2417
rect 12983 2391 12989 2417
rect 12577 2383 12989 2391
rect 9383 2370 9418 2371
rect 8698 2229 9261 2257
rect 9362 2363 9418 2370
rect 9362 2343 9391 2363
rect 9411 2343 9418 2363
rect 9362 2338 9418 2343
rect 9591 2367 9641 2375
rect 9591 2346 9607 2367
rect 9629 2346 9641 2367
rect 8277 2202 8624 2206
rect 8277 2176 8286 2202
rect 8305 2176 8624 2202
rect 8699 2201 8733 2229
rect 8277 2171 8624 2176
rect 8698 2198 8734 2201
rect 8698 2179 8706 2198
rect 8726 2179 8734 2198
rect 8698 2175 8734 2179
rect 8584 2141 8624 2171
rect 8370 2136 8405 2137
rect 8349 2129 8405 2136
rect 8349 2109 8378 2129
rect 8398 2109 8405 2129
rect 8349 2104 8405 2109
rect 8581 2130 8624 2141
rect 8581 2110 8589 2130
rect 8613 2124 8624 2130
rect 8796 2132 8828 2139
rect 8613 2110 8623 2124
rect 8349 1898 8383 2104
rect 8581 2101 8623 2110
rect 8796 2112 8802 2132
rect 8823 2112 8828 2132
rect 8796 2084 8828 2112
rect 9362 2132 9396 2338
rect 9591 2337 9641 2346
rect 9809 2366 9841 2373
rect 9809 2346 9815 2366
rect 9836 2346 9841 2366
rect 9809 2318 9841 2346
rect 12577 2355 12609 2383
rect 13022 2363 13056 2569
rect 13514 2439 13548 2645
rect 13742 2642 13789 2648
rect 13961 2673 13993 2680
rect 13961 2653 13967 2673
rect 13988 2653 13993 2673
rect 13961 2625 13993 2653
rect 13581 2617 13993 2625
rect 13581 2591 13587 2617
rect 13613 2591 13993 2617
rect 13581 2589 13993 2591
rect 13583 2588 13623 2589
rect 13961 2524 13993 2589
rect 16630 2676 16662 2741
rect 17000 2676 17040 2677
rect 16630 2674 17042 2676
rect 16630 2648 17010 2674
rect 17036 2648 17042 2674
rect 16630 2640 17042 2648
rect 16630 2612 16662 2640
rect 16630 2592 16635 2612
rect 16656 2592 16662 2612
rect 16630 2585 16662 2592
rect 16830 2612 16880 2621
rect 17075 2620 17109 2826
rect 17643 2846 17675 2874
rect 17643 2826 17648 2846
rect 17669 2826 17675 2846
rect 17848 2848 17890 2857
rect 18088 2854 18122 3060
rect 17848 2834 17858 2848
rect 17643 2819 17675 2826
rect 17847 2828 17858 2834
rect 17882 2828 17890 2848
rect 17847 2817 17890 2828
rect 18066 2849 18122 2854
rect 18066 2829 18073 2849
rect 18093 2829 18122 2849
rect 18066 2822 18122 2829
rect 18066 2821 18101 2822
rect 17847 2787 17887 2817
rect 17737 2779 17773 2783
rect 17737 2760 17745 2779
rect 17765 2760 17773 2779
rect 17737 2757 17773 2760
rect 17847 2782 18194 2787
rect 17738 2729 17772 2757
rect 17847 2756 18166 2782
rect 18185 2756 18194 2782
rect 17847 2752 18194 2756
rect 16830 2591 16842 2612
rect 16864 2591 16880 2612
rect 16830 2583 16880 2591
rect 17053 2615 17109 2620
rect 17053 2595 17060 2615
rect 17080 2595 17109 2615
rect 17053 2588 17109 2595
rect 17210 2701 17773 2729
rect 17053 2587 17088 2588
rect 13961 2504 13965 2524
rect 13986 2504 13993 2524
rect 16835 2550 16876 2583
rect 17210 2550 17250 2701
rect 18299 2582 18334 3176
rect 18699 2723 18731 4376
rect 19870 4225 19910 4376
rect 20244 4343 20285 4376
rect 20032 4338 20067 4339
rect 19347 4197 19910 4225
rect 20011 4331 20067 4338
rect 20011 4311 20040 4331
rect 20060 4311 20067 4331
rect 20011 4306 20067 4311
rect 20240 4335 20290 4343
rect 20240 4314 20256 4335
rect 20278 4314 20290 4335
rect 18926 4170 19273 4174
rect 18926 4144 18935 4170
rect 18954 4144 19273 4170
rect 19348 4169 19382 4197
rect 18926 4139 19273 4144
rect 19347 4166 19383 4169
rect 19347 4147 19355 4166
rect 19375 4147 19383 4166
rect 19347 4143 19383 4147
rect 19233 4109 19273 4139
rect 19019 4104 19054 4105
rect 18998 4097 19054 4104
rect 18998 4077 19027 4097
rect 19047 4077 19054 4097
rect 18998 4072 19054 4077
rect 19230 4098 19273 4109
rect 19230 4078 19238 4098
rect 19262 4092 19273 4098
rect 19445 4100 19477 4107
rect 19262 4078 19272 4092
rect 18998 3866 19032 4072
rect 19230 4069 19272 4078
rect 19445 4080 19451 4100
rect 19472 4080 19477 4100
rect 19445 4052 19477 4080
rect 20011 4100 20045 4306
rect 20240 4305 20290 4314
rect 20458 4334 20490 4341
rect 20458 4314 20464 4334
rect 20485 4314 20490 4334
rect 20458 4286 20490 4314
rect 20078 4278 20490 4286
rect 20078 4252 20084 4278
rect 20110 4252 20490 4278
rect 20078 4250 20490 4252
rect 20080 4249 20120 4250
rect 20458 4185 20490 4250
rect 20458 4165 20462 4185
rect 20483 4165 20490 4185
rect 20458 4158 20490 4165
rect 20011 4092 20046 4100
rect 20011 4072 20019 4092
rect 20039 4072 20046 4092
rect 20011 4067 20046 4072
rect 20011 4066 20043 4067
rect 19065 4044 19477 4052
rect 19065 4018 19071 4044
rect 19097 4018 19477 4044
rect 19065 4016 19477 4018
rect 19067 4015 19107 4016
rect 19445 3951 19477 4016
rect 19445 3931 19449 3951
rect 19470 3931 19477 3951
rect 19445 3924 19477 3931
rect 19922 3962 20274 3993
rect 18998 3858 19033 3866
rect 18998 3838 19006 3858
rect 19026 3838 19033 3858
rect 18998 3822 19033 3838
rect 19922 3822 19953 3962
rect 20246 3930 20274 3962
rect 20031 3923 20066 3924
rect 18996 3803 19953 3822
rect 20010 3916 20066 3923
rect 20010 3896 20039 3916
rect 20059 3896 20066 3916
rect 20010 3891 20066 3896
rect 20240 3918 20280 3930
rect 20240 3897 20246 3918
rect 20268 3897 20280 3918
rect 20240 3892 20280 3897
rect 20457 3919 20489 3926
rect 20457 3899 20463 3919
rect 20484 3899 20489 3919
rect 18835 3751 18864 3753
rect 18835 3746 19208 3751
rect 18835 3728 18842 3746
rect 18862 3728 19208 3746
rect 18835 3723 19208 3728
rect 18840 3721 19208 3723
rect 18969 3684 19004 3685
rect 19184 3684 19208 3721
rect 18948 3677 19004 3684
rect 18948 3657 18977 3677
rect 18997 3657 19004 3677
rect 18948 3652 19004 3657
rect 19179 3679 19216 3684
rect 19179 3660 19187 3679
rect 19210 3660 19216 3679
rect 19179 3654 19216 3660
rect 19395 3680 19427 3687
rect 19395 3660 19401 3680
rect 19422 3660 19427 3680
rect 18948 3448 18982 3652
rect 19395 3632 19427 3660
rect 20010 3685 20044 3891
rect 20457 3871 20489 3899
rect 20077 3863 20489 3871
rect 20077 3837 20083 3863
rect 20109 3837 20489 3863
rect 20077 3835 20489 3837
rect 20079 3834 20119 3835
rect 20457 3770 20489 3835
rect 20457 3750 20461 3770
rect 20482 3750 20489 3770
rect 20457 3743 20489 3750
rect 20010 3677 20045 3685
rect 20010 3657 20018 3677
rect 20038 3657 20045 3677
rect 20010 3652 20045 3657
rect 20010 3651 20042 3652
rect 19015 3624 19427 3632
rect 19015 3598 19021 3624
rect 19047 3598 19427 3624
rect 19015 3596 19427 3598
rect 19017 3595 19057 3596
rect 19395 3531 19427 3596
rect 19395 3511 19399 3531
rect 19420 3511 19427 3531
rect 19395 3504 19427 3511
rect 18946 3438 18986 3448
rect 18946 3418 18956 3438
rect 18976 3418 18986 3438
rect 19881 3424 20290 3425
rect 18946 3194 18986 3418
rect 19875 3395 20290 3424
rect 19875 3244 19915 3395
rect 20249 3362 20290 3395
rect 20037 3357 20072 3358
rect 19352 3216 19915 3244
rect 20016 3350 20072 3357
rect 20016 3330 20045 3350
rect 20065 3330 20072 3350
rect 20016 3325 20072 3330
rect 20245 3354 20295 3362
rect 20245 3333 20261 3354
rect 20283 3333 20295 3354
rect 18946 3160 19273 3194
rect 19353 3188 19387 3216
rect 19352 3185 19388 3188
rect 19352 3166 19360 3185
rect 19380 3166 19388 3185
rect 19352 3162 19388 3166
rect 18963 3159 19273 3160
rect 19238 3130 19273 3159
rect 19024 3123 19059 3124
rect 19003 3116 19059 3123
rect 19003 3096 19032 3116
rect 19052 3096 19059 3116
rect 19003 3091 19059 3096
rect 19233 3118 19275 3130
rect 19233 3098 19242 3118
rect 19266 3098 19275 3118
rect 19003 2885 19037 3091
rect 19233 3090 19275 3098
rect 19450 3119 19482 3126
rect 19450 3099 19456 3119
rect 19477 3099 19482 3119
rect 19450 3071 19482 3099
rect 20016 3119 20050 3325
rect 20245 3324 20295 3333
rect 20463 3353 20495 3360
rect 20463 3333 20469 3353
rect 20490 3333 20495 3353
rect 20463 3305 20495 3333
rect 20083 3297 20495 3305
rect 20083 3271 20089 3297
rect 20115 3271 20495 3297
rect 20083 3269 20495 3271
rect 20085 3268 20125 3269
rect 20463 3204 20495 3269
rect 20463 3184 20467 3204
rect 20488 3184 20495 3204
rect 20463 3177 20495 3184
rect 20016 3111 20051 3119
rect 20016 3091 20024 3111
rect 20044 3091 20051 3111
rect 20016 3086 20051 3091
rect 20016 3085 20048 3086
rect 19070 3063 19482 3071
rect 19070 3037 19076 3063
rect 19102 3037 19482 3063
rect 19070 3035 19482 3037
rect 19072 3034 19112 3035
rect 19450 2970 19482 3035
rect 19450 2950 19454 2970
rect 19475 2950 19482 2970
rect 19450 2943 19482 2950
rect 19927 2981 20279 3012
rect 19003 2877 19038 2885
rect 19003 2857 19011 2877
rect 19031 2857 19038 2877
rect 19003 2841 19038 2857
rect 19927 2841 19958 2981
rect 20251 2949 20279 2981
rect 20036 2942 20071 2943
rect 19001 2822 19958 2841
rect 20015 2935 20071 2942
rect 20015 2915 20044 2935
rect 20064 2915 20071 2935
rect 20015 2910 20071 2915
rect 20245 2937 20285 2949
rect 20245 2916 20251 2937
rect 20273 2916 20285 2937
rect 20245 2911 20285 2916
rect 20462 2938 20494 2945
rect 20462 2918 20468 2938
rect 20489 2918 20494 2938
rect 18695 2690 19065 2723
rect 18699 2688 18731 2690
rect 18816 2656 18851 2657
rect 18795 2649 18851 2656
rect 19028 2655 19065 2690
rect 20015 2704 20049 2910
rect 20462 2890 20494 2918
rect 20082 2882 20494 2890
rect 20082 2856 20088 2882
rect 20114 2856 20494 2882
rect 20082 2854 20494 2856
rect 20084 2853 20124 2854
rect 20462 2789 20494 2854
rect 20462 2769 20466 2789
rect 20487 2769 20494 2789
rect 20462 2762 20494 2769
rect 20015 2696 20050 2704
rect 20015 2676 20023 2696
rect 20043 2676 20050 2696
rect 20015 2671 20050 2676
rect 20015 2670 20047 2671
rect 18795 2629 18824 2649
rect 18844 2629 18851 2649
rect 18795 2624 18851 2629
rect 19023 2653 19070 2655
rect 19023 2627 19035 2653
rect 19060 2627 19070 2653
rect 18299 2576 18337 2582
rect 18299 2556 18309 2576
rect 18329 2556 18337 2576
rect 18299 2554 18337 2556
rect 16835 2521 17250 2550
rect 18302 2548 18337 2554
rect 16835 2520 17244 2521
rect 13961 2497 13993 2504
rect 17858 2483 17890 2490
rect 14607 2466 15016 2467
rect 13514 2433 13549 2439
rect 14601 2437 15016 2466
rect 13514 2431 13552 2433
rect 13514 2411 13522 2431
rect 13542 2411 13552 2431
rect 13514 2405 13552 2411
rect 12577 2335 12582 2355
rect 12603 2335 12609 2355
rect 12577 2328 12609 2335
rect 12786 2356 12825 2362
rect 12786 2337 12797 2356
rect 12820 2337 12825 2356
rect 12786 2324 12825 2337
rect 13000 2358 13056 2363
rect 13000 2338 13007 2358
rect 13027 2338 13056 2358
rect 13000 2331 13056 2338
rect 13000 2330 13035 2331
rect 9429 2310 9841 2318
rect 11804 2316 11836 2317
rect 9429 2284 9435 2310
rect 9461 2284 9841 2310
rect 9429 2282 9841 2284
rect 11801 2311 11836 2316
rect 11801 2291 11808 2311
rect 11828 2291 11836 2311
rect 11801 2283 11836 2291
rect 9431 2281 9471 2282
rect 9809 2217 9841 2282
rect 9809 2197 9813 2217
rect 9834 2197 9841 2217
rect 9809 2190 9841 2197
rect 11357 2218 11389 2225
rect 11357 2198 11364 2218
rect 11385 2198 11389 2218
rect 11357 2133 11389 2198
rect 11727 2133 11767 2134
rect 9362 2124 9397 2132
rect 9362 2104 9370 2124
rect 9390 2104 9397 2124
rect 9362 2099 9397 2104
rect 11357 2131 11769 2133
rect 11357 2105 11737 2131
rect 11763 2105 11769 2131
rect 9362 2098 9394 2099
rect 8416 2076 8828 2084
rect 8416 2050 8422 2076
rect 8448 2050 8828 2076
rect 8416 2048 8828 2050
rect 8418 2047 8458 2048
rect 8796 1983 8828 2048
rect 11357 2097 11769 2105
rect 11357 2069 11389 2097
rect 11802 2077 11836 2283
rect 12793 2293 12823 2324
rect 13103 2293 13140 2299
rect 12793 2288 13140 2293
rect 12793 2269 13109 2288
rect 13132 2269 13140 2288
rect 12793 2263 13140 2269
rect 13103 2258 13140 2263
rect 11357 2049 11362 2069
rect 11383 2049 11389 2069
rect 11357 2042 11389 2049
rect 11566 2071 11606 2076
rect 11566 2050 11578 2071
rect 11600 2050 11606 2071
rect 11566 2038 11606 2050
rect 11780 2072 11836 2077
rect 11780 2052 11787 2072
rect 11807 2052 11836 2072
rect 11780 2045 11836 2052
rect 11893 2146 12850 2165
rect 11780 2044 11815 2045
rect 8796 1963 8800 1983
rect 8821 1963 8828 1983
rect 8796 1956 8828 1963
rect 9273 1994 9625 2025
rect 8349 1890 8384 1898
rect 8349 1870 8357 1890
rect 8377 1870 8384 1890
rect 8349 1854 8384 1870
rect 9273 1854 9304 1994
rect 9597 1962 9625 1994
rect 11572 2006 11600 2038
rect 11893 2006 11924 2146
rect 12813 2130 12848 2146
rect 12813 2110 12820 2130
rect 12840 2110 12848 2130
rect 12813 2102 12848 2110
rect 11572 1975 11924 2006
rect 12369 2037 12401 2044
rect 12369 2017 12376 2037
rect 12397 2017 12401 2037
rect 9382 1955 9417 1956
rect 8347 1835 9304 1854
rect 9361 1948 9417 1955
rect 9361 1928 9390 1948
rect 9410 1928 9417 1948
rect 9361 1923 9417 1928
rect 9591 1950 9631 1962
rect 9591 1929 9597 1950
rect 9619 1929 9631 1950
rect 9591 1924 9631 1929
rect 9808 1951 9840 1958
rect 9808 1931 9814 1951
rect 9835 1931 9840 1951
rect 8137 1753 8567 1782
rect 8137 1748 8221 1753
rect 8320 1716 8355 1717
rect 6181 1533 6590 1534
rect 7485 1520 7495 1540
rect 7515 1520 7525 1540
rect 7485 1510 7525 1520
rect 8299 1709 8355 1716
rect 8299 1689 8328 1709
rect 8348 1689 8355 1709
rect 8299 1684 8355 1689
rect 8529 1710 8567 1753
rect 8529 1693 8534 1710
rect 8558 1693 8567 1710
rect 1763 1299 1768 1319
rect 1789 1299 1795 1319
rect 1763 1292 1795 1299
rect 1974 1319 2011 1325
rect 1974 1300 1980 1319
rect 2003 1300 2011 1319
rect 1974 1295 2011 1300
rect 2186 1322 2242 1327
rect 2186 1302 2193 1322
rect 2213 1302 2242 1322
rect 2186 1295 2242 1302
rect 3016 1491 3056 1501
rect 3016 1471 3026 1491
rect 3046 1471 3056 1491
rect 3951 1477 4360 1478
rect 1982 1258 2006 1295
rect 2186 1294 2221 1295
rect 1982 1256 2350 1258
rect 1982 1251 2355 1256
rect 1982 1233 2328 1251
rect 2348 1233 2355 1251
rect 1982 1228 2355 1233
rect 2326 1226 2355 1228
rect 3016 1247 3056 1471
rect 3945 1448 4360 1477
rect 3945 1297 3985 1448
rect 4319 1415 4360 1448
rect 7044 1447 7076 1454
rect 7044 1427 7051 1447
rect 7072 1427 7076 1447
rect 4107 1410 4142 1411
rect 3422 1269 3985 1297
rect 4086 1403 4142 1410
rect 4086 1383 4115 1403
rect 4135 1383 4142 1403
rect 4086 1378 4142 1383
rect 4315 1407 4365 1415
rect 4315 1386 4331 1407
rect 4353 1386 4365 1407
rect 3016 1213 3343 1247
rect 3423 1241 3457 1269
rect 3422 1238 3458 1241
rect 3422 1219 3430 1238
rect 3450 1219 3458 1238
rect 3422 1215 3458 1219
rect 3033 1212 3343 1213
rect 3308 1183 3343 1212
rect 3094 1176 3129 1177
rect 701 1060 706 1080
rect 727 1060 733 1080
rect 701 1053 733 1060
rect 910 1082 950 1087
rect 910 1061 922 1082
rect 944 1061 950 1082
rect 910 1049 950 1061
rect 1124 1083 1180 1088
rect 1124 1063 1131 1083
rect 1151 1063 1180 1083
rect 1124 1056 1180 1063
rect 1237 1157 2194 1176
rect 3073 1169 3129 1176
rect 1124 1055 1159 1056
rect 916 1017 944 1049
rect 1237 1017 1268 1157
rect 2157 1141 2192 1157
rect 2157 1121 2164 1141
rect 2184 1121 2192 1141
rect 2157 1113 2192 1121
rect 916 986 1268 1017
rect 1713 1048 1745 1055
rect 1713 1028 1720 1048
rect 1741 1028 1745 1048
rect 1713 963 1745 1028
rect 2083 963 2123 964
rect 1713 961 2125 963
rect 1713 935 2093 961
rect 2119 935 2125 961
rect 1713 927 2125 935
rect 1147 912 1179 913
rect 1144 907 1179 912
rect 1144 887 1151 907
rect 1171 887 1179 907
rect 1144 879 1179 887
rect 700 814 732 821
rect 700 794 707 814
rect 728 794 732 814
rect 700 729 732 794
rect 1070 729 1110 730
rect 700 727 1112 729
rect 700 701 1080 727
rect 1106 701 1112 727
rect 700 693 1112 701
rect 700 665 732 693
rect 700 645 705 665
rect 726 645 732 665
rect 700 638 732 645
rect 900 665 950 674
rect 1145 673 1179 879
rect 1713 899 1745 927
rect 1713 879 1718 899
rect 1739 879 1745 899
rect 1918 901 1960 910
rect 2158 907 2192 1113
rect 1918 887 1928 901
rect 1713 872 1745 879
rect 1917 881 1928 887
rect 1952 881 1960 901
rect 1917 870 1960 881
rect 2136 902 2192 907
rect 2136 882 2143 902
rect 2163 882 2192 902
rect 3073 1149 3102 1169
rect 3122 1149 3129 1169
rect 3073 1144 3129 1149
rect 3303 1171 3345 1183
rect 3303 1151 3312 1171
rect 3336 1151 3345 1171
rect 3073 938 3107 1144
rect 3303 1143 3345 1151
rect 3520 1172 3552 1179
rect 3520 1152 3526 1172
rect 3547 1152 3552 1172
rect 3520 1124 3552 1152
rect 4086 1172 4120 1378
rect 4315 1377 4365 1386
rect 4533 1406 4565 1413
rect 4533 1386 4539 1406
rect 4560 1386 4565 1406
rect 4533 1358 4565 1386
rect 4153 1350 4565 1358
rect 4153 1324 4159 1350
rect 4185 1324 4565 1350
rect 4153 1322 4565 1324
rect 4155 1321 4195 1322
rect 4533 1257 4565 1322
rect 7044 1362 7076 1427
rect 7414 1362 7454 1363
rect 7044 1360 7456 1362
rect 7044 1334 7424 1360
rect 7450 1334 7456 1360
rect 7044 1326 7456 1334
rect 6429 1306 6461 1307
rect 6426 1301 6461 1306
rect 6426 1281 6433 1301
rect 6453 1281 6461 1301
rect 6426 1273 6461 1281
rect 4533 1237 4537 1257
rect 4558 1237 4565 1257
rect 4533 1230 4565 1237
rect 5982 1208 6014 1215
rect 5982 1188 5989 1208
rect 6010 1188 6014 1208
rect 4086 1164 4121 1172
rect 4086 1144 4094 1164
rect 4114 1144 4121 1164
rect 4086 1139 4121 1144
rect 4086 1138 4118 1139
rect 3140 1116 3552 1124
rect 3140 1090 3146 1116
rect 3172 1090 3552 1116
rect 3140 1088 3552 1090
rect 3142 1087 3182 1088
rect 3520 1023 3552 1088
rect 5982 1123 6014 1188
rect 6352 1123 6392 1124
rect 5982 1121 6394 1123
rect 5982 1095 6362 1121
rect 6388 1095 6394 1121
rect 5982 1087 6394 1095
rect 3520 1003 3524 1023
rect 3545 1003 3552 1023
rect 3520 996 3552 1003
rect 3997 1034 4349 1065
rect 3073 930 3108 938
rect 3073 910 3081 930
rect 3101 910 3108 930
rect 3073 894 3108 910
rect 3997 894 4028 1034
rect 4321 1002 4349 1034
rect 5982 1059 6014 1087
rect 6427 1067 6461 1273
rect 7044 1298 7076 1326
rect 7489 1306 7523 1510
rect 8299 1480 8333 1684
rect 8529 1681 8567 1693
rect 8746 1712 8778 1719
rect 8746 1692 8752 1712
rect 8773 1692 8778 1712
rect 8746 1664 8778 1692
rect 9361 1717 9395 1923
rect 9808 1903 9840 1931
rect 9428 1895 9840 1903
rect 12369 1952 12401 2017
rect 12739 1952 12779 1953
rect 12369 1950 12781 1952
rect 12369 1924 12749 1950
rect 12775 1924 12781 1950
rect 12369 1916 12781 1924
rect 11803 1901 11835 1902
rect 9428 1869 9434 1895
rect 9460 1869 9840 1895
rect 9428 1867 9840 1869
rect 11800 1896 11835 1901
rect 11800 1876 11807 1896
rect 11827 1876 11835 1896
rect 11800 1868 11835 1876
rect 9430 1866 9470 1867
rect 9808 1802 9840 1867
rect 9808 1782 9812 1802
rect 9833 1782 9840 1802
rect 9808 1775 9840 1782
rect 11356 1803 11388 1810
rect 11356 1783 11363 1803
rect 11384 1783 11388 1803
rect 11356 1718 11388 1783
rect 11726 1718 11766 1719
rect 9361 1709 9396 1717
rect 9361 1689 9369 1709
rect 9389 1689 9396 1709
rect 9361 1684 9396 1689
rect 11356 1716 11768 1718
rect 11356 1690 11736 1716
rect 11762 1690 11768 1716
rect 9361 1683 9393 1684
rect 8366 1656 8778 1664
rect 8366 1630 8372 1656
rect 8398 1630 8778 1656
rect 8366 1628 8778 1630
rect 8368 1627 8408 1628
rect 8746 1563 8778 1628
rect 11356 1682 11768 1690
rect 11356 1654 11388 1682
rect 11356 1634 11361 1654
rect 11382 1634 11388 1654
rect 11356 1627 11388 1634
rect 11556 1654 11606 1663
rect 11801 1662 11835 1868
rect 12369 1888 12401 1916
rect 12369 1868 12374 1888
rect 12395 1868 12401 1888
rect 12369 1861 12401 1868
rect 12576 1889 12618 1897
rect 12814 1896 12848 2102
rect 12576 1869 12585 1889
rect 12609 1869 12618 1889
rect 12576 1857 12618 1869
rect 12792 1891 12848 1896
rect 12792 1871 12799 1891
rect 12819 1871 12848 1891
rect 12792 1864 12848 1871
rect 12792 1863 12827 1864
rect 12578 1828 12613 1857
rect 12578 1827 12888 1828
rect 12463 1821 12499 1825
rect 12463 1802 12471 1821
rect 12491 1802 12499 1821
rect 12463 1799 12499 1802
rect 12464 1771 12498 1799
rect 12578 1793 12905 1827
rect 11556 1633 11568 1654
rect 11590 1633 11606 1654
rect 11556 1625 11606 1633
rect 11779 1657 11835 1662
rect 11779 1637 11786 1657
rect 11806 1637 11835 1657
rect 11779 1630 11835 1637
rect 11936 1743 12499 1771
rect 11779 1629 11814 1630
rect 8746 1543 8750 1563
rect 8771 1543 8778 1563
rect 11561 1592 11602 1625
rect 11936 1592 11976 1743
rect 11561 1563 11976 1592
rect 12865 1569 12905 1793
rect 13517 1811 13552 2405
rect 14601 2286 14641 2437
rect 14975 2404 15016 2437
rect 17858 2463 17865 2483
rect 17886 2463 17890 2483
rect 14763 2399 14798 2400
rect 14078 2258 14641 2286
rect 14742 2392 14798 2399
rect 14742 2372 14771 2392
rect 14791 2372 14798 2392
rect 14742 2367 14798 2372
rect 14971 2396 15021 2404
rect 14971 2375 14987 2396
rect 15009 2375 15021 2396
rect 13657 2231 14004 2235
rect 13657 2205 13666 2231
rect 13685 2205 14004 2231
rect 14079 2230 14113 2258
rect 13657 2200 14004 2205
rect 14078 2227 14114 2230
rect 14078 2208 14086 2227
rect 14106 2208 14114 2227
rect 14078 2204 14114 2208
rect 13964 2170 14004 2200
rect 13750 2165 13785 2166
rect 13729 2158 13785 2165
rect 13729 2138 13758 2158
rect 13778 2138 13785 2158
rect 13729 2133 13785 2138
rect 13961 2159 14004 2170
rect 13961 2139 13969 2159
rect 13993 2153 14004 2159
rect 14176 2161 14208 2168
rect 13993 2139 14003 2153
rect 13729 1927 13763 2133
rect 13961 2130 14003 2139
rect 14176 2141 14182 2161
rect 14203 2141 14208 2161
rect 14176 2113 14208 2141
rect 14742 2161 14776 2367
rect 14971 2366 15021 2375
rect 15189 2395 15221 2402
rect 15189 2375 15195 2395
rect 15216 2375 15221 2395
rect 15189 2347 15221 2375
rect 14809 2339 15221 2347
rect 14809 2313 14815 2339
rect 14841 2313 15221 2339
rect 14809 2311 15221 2313
rect 14811 2310 14851 2311
rect 15189 2246 15221 2311
rect 17858 2398 17890 2463
rect 18228 2398 18268 2399
rect 17858 2396 18270 2398
rect 17858 2370 18238 2396
rect 18264 2370 18270 2396
rect 17858 2362 18270 2370
rect 17858 2334 17890 2362
rect 18303 2342 18337 2548
rect 18795 2418 18829 2624
rect 19023 2621 19070 2627
rect 19242 2652 19274 2659
rect 19242 2632 19248 2652
rect 19269 2632 19274 2652
rect 19242 2604 19274 2632
rect 18862 2596 19274 2604
rect 18862 2570 18868 2596
rect 18894 2570 19274 2596
rect 18862 2568 19274 2570
rect 18864 2567 18904 2568
rect 19242 2503 19274 2568
rect 19242 2483 19246 2503
rect 19267 2483 19274 2503
rect 19242 2476 19274 2483
rect 19888 2445 20297 2446
rect 18795 2412 18830 2418
rect 19882 2416 20297 2445
rect 18795 2410 18833 2412
rect 18795 2390 18803 2410
rect 18823 2390 18833 2410
rect 18795 2384 18833 2390
rect 17858 2314 17863 2334
rect 17884 2314 17890 2334
rect 17858 2307 17890 2314
rect 18067 2335 18106 2341
rect 18067 2316 18078 2335
rect 18101 2316 18106 2335
rect 18067 2303 18106 2316
rect 18281 2337 18337 2342
rect 18281 2317 18288 2337
rect 18308 2317 18337 2337
rect 18281 2310 18337 2317
rect 18281 2309 18316 2310
rect 17085 2295 17117 2296
rect 17082 2290 17117 2295
rect 17082 2270 17089 2290
rect 17109 2270 17117 2290
rect 17082 2262 17117 2270
rect 15189 2226 15193 2246
rect 15214 2226 15221 2246
rect 15189 2219 15221 2226
rect 16638 2197 16670 2204
rect 16638 2177 16645 2197
rect 16666 2177 16670 2197
rect 14742 2153 14777 2161
rect 14742 2133 14750 2153
rect 14770 2133 14777 2153
rect 14742 2128 14777 2133
rect 14742 2127 14774 2128
rect 13796 2105 14208 2113
rect 13796 2079 13802 2105
rect 13828 2079 14208 2105
rect 13796 2077 14208 2079
rect 13798 2076 13838 2077
rect 14176 2012 14208 2077
rect 16638 2112 16670 2177
rect 17008 2112 17048 2113
rect 16638 2110 17050 2112
rect 16638 2084 17018 2110
rect 17044 2084 17050 2110
rect 16638 2076 17050 2084
rect 14176 1992 14180 2012
rect 14201 1992 14208 2012
rect 14176 1985 14208 1992
rect 14653 2023 15005 2054
rect 13729 1919 13764 1927
rect 13729 1899 13737 1919
rect 13757 1899 13764 1919
rect 13729 1883 13764 1899
rect 14653 1883 14684 2023
rect 14977 1991 15005 2023
rect 16638 2048 16670 2076
rect 17083 2056 17117 2262
rect 18074 2272 18104 2303
rect 18384 2272 18421 2278
rect 18074 2267 18421 2272
rect 18074 2248 18390 2267
rect 18413 2248 18421 2267
rect 18074 2242 18421 2248
rect 18384 2237 18421 2242
rect 16638 2028 16643 2048
rect 16664 2028 16670 2048
rect 16638 2021 16670 2028
rect 16847 2050 16887 2055
rect 16847 2029 16859 2050
rect 16881 2029 16887 2050
rect 16847 2017 16887 2029
rect 17061 2051 17117 2056
rect 17061 2031 17068 2051
rect 17088 2031 17117 2051
rect 17061 2024 17117 2031
rect 17174 2125 18131 2144
rect 17061 2023 17096 2024
rect 14762 1984 14797 1985
rect 13727 1864 14684 1883
rect 14741 1977 14797 1984
rect 14741 1957 14770 1977
rect 14790 1957 14797 1977
rect 14741 1952 14797 1957
rect 14971 1979 15011 1991
rect 14971 1958 14977 1979
rect 14999 1958 15011 1979
rect 14971 1953 15011 1958
rect 15188 1980 15220 1987
rect 15188 1960 15194 1980
rect 15215 1960 15220 1980
rect 13517 1782 13947 1811
rect 13517 1777 13601 1782
rect 13700 1745 13735 1746
rect 11561 1562 11970 1563
rect 8746 1536 8778 1543
rect 12865 1549 12875 1569
rect 12895 1549 12905 1569
rect 12865 1539 12905 1549
rect 13679 1738 13735 1745
rect 13679 1718 13708 1738
rect 13728 1718 13735 1738
rect 13679 1713 13735 1718
rect 13909 1739 13947 1782
rect 13909 1722 13914 1739
rect 13938 1722 13947 1739
rect 7044 1278 7049 1298
rect 7070 1278 7076 1298
rect 7044 1271 7076 1278
rect 7255 1298 7292 1304
rect 7255 1279 7261 1298
rect 7284 1279 7292 1298
rect 7255 1274 7292 1279
rect 7467 1301 7523 1306
rect 7467 1281 7474 1301
rect 7494 1281 7523 1301
rect 7467 1274 7523 1281
rect 8297 1470 8337 1480
rect 8297 1450 8307 1470
rect 8327 1450 8337 1470
rect 12424 1476 12456 1483
rect 9232 1456 9641 1457
rect 7263 1237 7287 1274
rect 7467 1273 7502 1274
rect 7263 1235 7631 1237
rect 7263 1230 7636 1235
rect 7263 1212 7609 1230
rect 7629 1212 7636 1230
rect 7263 1207 7636 1212
rect 7607 1205 7636 1207
rect 8297 1226 8337 1450
rect 9226 1427 9641 1456
rect 9226 1276 9266 1427
rect 9600 1394 9641 1427
rect 12424 1456 12431 1476
rect 12452 1456 12456 1476
rect 9388 1389 9423 1390
rect 8703 1248 9266 1276
rect 9367 1382 9423 1389
rect 9367 1362 9396 1382
rect 9416 1362 9423 1382
rect 9367 1357 9423 1362
rect 9596 1386 9646 1394
rect 9596 1365 9612 1386
rect 9634 1365 9646 1386
rect 8297 1192 8624 1226
rect 8704 1220 8738 1248
rect 8703 1217 8739 1220
rect 8703 1198 8711 1217
rect 8731 1198 8739 1217
rect 8703 1194 8739 1198
rect 8314 1191 8624 1192
rect 8589 1162 8624 1191
rect 8375 1155 8410 1156
rect 5982 1039 5987 1059
rect 6008 1039 6014 1059
rect 5982 1032 6014 1039
rect 6191 1061 6231 1066
rect 6191 1040 6203 1061
rect 6225 1040 6231 1061
rect 6191 1028 6231 1040
rect 6405 1062 6461 1067
rect 6405 1042 6412 1062
rect 6432 1042 6461 1062
rect 6405 1035 6461 1042
rect 6518 1136 7475 1155
rect 8354 1148 8410 1155
rect 6405 1034 6440 1035
rect 4106 995 4141 996
rect 2136 875 2192 882
rect 3071 875 4028 894
rect 4085 988 4141 995
rect 4085 968 4114 988
rect 4134 968 4141 988
rect 4085 963 4141 968
rect 4315 990 4355 1002
rect 4315 969 4321 990
rect 4343 969 4355 990
rect 4315 964 4355 969
rect 4532 991 4564 998
rect 4532 971 4538 991
rect 4559 971 4564 991
rect 2136 874 2171 875
rect 1917 840 1957 870
rect 1807 832 1843 836
rect 1807 813 1815 832
rect 1835 813 1843 832
rect 1807 810 1843 813
rect 1917 835 2264 840
rect 1808 782 1842 810
rect 1917 809 2236 835
rect 2255 809 2264 835
rect 1917 805 2264 809
rect 900 644 912 665
rect 934 644 950 665
rect 900 636 950 644
rect 1123 668 1179 673
rect 1123 648 1130 668
rect 1150 648 1179 668
rect 1123 641 1179 648
rect 1280 754 1843 782
rect 4085 757 4119 963
rect 4532 943 4564 971
rect 6197 996 6225 1028
rect 6518 996 6549 1136
rect 7438 1120 7473 1136
rect 7438 1100 7445 1120
rect 7465 1100 7473 1120
rect 7438 1092 7473 1100
rect 6197 965 6549 996
rect 6994 1027 7026 1034
rect 6994 1007 7001 1027
rect 7022 1007 7026 1027
rect 4152 935 4564 943
rect 4152 909 4158 935
rect 4184 909 4564 935
rect 4152 907 4564 909
rect 4154 906 4194 907
rect 4532 842 4564 907
rect 6994 942 7026 1007
rect 7364 942 7404 943
rect 6994 940 7406 942
rect 6994 914 7374 940
rect 7400 914 7406 940
rect 6994 906 7406 914
rect 6428 891 6460 892
rect 6425 886 6460 891
rect 6425 866 6432 886
rect 6452 866 6460 886
rect 6425 858 6460 866
rect 4532 822 4536 842
rect 4557 822 4564 842
rect 4532 815 4564 822
rect 5981 793 6013 800
rect 5981 773 5988 793
rect 6009 773 6013 793
rect 1123 640 1158 641
rect 905 603 946 636
rect 1280 603 1320 754
rect 4085 749 4120 757
rect 4085 729 4093 749
rect 4113 729 4120 749
rect 4085 724 4120 729
rect 4085 723 4117 724
rect 5981 708 6013 773
rect 6351 708 6391 709
rect 5981 706 6393 708
rect 5981 680 6361 706
rect 6387 680 6393 706
rect 5981 672 6393 680
rect 5981 644 6013 672
rect 5981 624 5986 644
rect 6007 624 6013 644
rect 5981 617 6013 624
rect 6181 644 6231 653
rect 6426 652 6460 858
rect 6994 878 7026 906
rect 6994 858 6999 878
rect 7020 858 7026 878
rect 7199 880 7241 889
rect 7439 886 7473 1092
rect 7199 866 7209 880
rect 6994 851 7026 858
rect 7198 860 7209 866
rect 7233 860 7241 880
rect 7198 849 7241 860
rect 7417 881 7473 886
rect 7417 861 7424 881
rect 7444 861 7473 881
rect 8354 1128 8383 1148
rect 8403 1128 8410 1148
rect 8354 1123 8410 1128
rect 8584 1150 8626 1162
rect 8584 1130 8593 1150
rect 8617 1130 8626 1150
rect 8354 917 8388 1123
rect 8584 1122 8626 1130
rect 8801 1151 8833 1158
rect 8801 1131 8807 1151
rect 8828 1131 8833 1151
rect 8801 1103 8833 1131
rect 9367 1151 9401 1357
rect 9596 1356 9646 1365
rect 9814 1385 9846 1392
rect 9814 1365 9820 1385
rect 9841 1365 9846 1385
rect 9814 1337 9846 1365
rect 9434 1329 9846 1337
rect 12424 1391 12456 1456
rect 12794 1391 12834 1392
rect 12424 1389 12836 1391
rect 12424 1363 12804 1389
rect 12830 1363 12836 1389
rect 12424 1355 12836 1363
rect 11809 1335 11841 1336
rect 9434 1303 9440 1329
rect 9466 1303 9846 1329
rect 9434 1301 9846 1303
rect 11806 1330 11841 1335
rect 11806 1310 11813 1330
rect 11833 1310 11841 1330
rect 11806 1302 11841 1310
rect 9436 1300 9476 1301
rect 9814 1236 9846 1301
rect 9814 1216 9818 1236
rect 9839 1216 9846 1236
rect 9814 1209 9846 1216
rect 11362 1237 11394 1244
rect 11362 1217 11369 1237
rect 11390 1217 11394 1237
rect 11362 1152 11394 1217
rect 11732 1152 11772 1153
rect 9367 1143 9402 1151
rect 9367 1123 9375 1143
rect 9395 1123 9402 1143
rect 9367 1118 9402 1123
rect 11362 1150 11774 1152
rect 11362 1124 11742 1150
rect 11768 1124 11774 1150
rect 9367 1117 9399 1118
rect 8421 1095 8833 1103
rect 8421 1069 8427 1095
rect 8453 1069 8833 1095
rect 8421 1067 8833 1069
rect 8423 1066 8463 1067
rect 8801 1002 8833 1067
rect 11362 1116 11774 1124
rect 11362 1088 11394 1116
rect 11807 1096 11841 1302
rect 12424 1327 12456 1355
rect 12869 1335 12903 1539
rect 13679 1509 13713 1713
rect 13909 1710 13947 1722
rect 14126 1741 14158 1748
rect 14126 1721 14132 1741
rect 14153 1721 14158 1741
rect 14126 1693 14158 1721
rect 14741 1746 14775 1952
rect 15188 1932 15220 1960
rect 16853 1985 16881 2017
rect 17174 1985 17205 2125
rect 18094 2109 18129 2125
rect 18094 2089 18101 2109
rect 18121 2089 18129 2109
rect 18094 2081 18129 2089
rect 16853 1954 17205 1985
rect 17650 2016 17682 2023
rect 17650 1996 17657 2016
rect 17678 1996 17682 2016
rect 14808 1924 15220 1932
rect 14808 1898 14814 1924
rect 14840 1898 15220 1924
rect 14808 1896 15220 1898
rect 14810 1895 14850 1896
rect 15188 1831 15220 1896
rect 17650 1931 17682 1996
rect 18020 1931 18060 1932
rect 17650 1929 18062 1931
rect 17650 1903 18030 1929
rect 18056 1903 18062 1929
rect 17650 1895 18062 1903
rect 17084 1880 17116 1881
rect 17081 1875 17116 1880
rect 17081 1855 17088 1875
rect 17108 1855 17116 1875
rect 17081 1847 17116 1855
rect 15188 1811 15192 1831
rect 15213 1811 15220 1831
rect 15188 1804 15220 1811
rect 16637 1782 16669 1789
rect 16637 1762 16644 1782
rect 16665 1762 16669 1782
rect 14741 1738 14776 1746
rect 14741 1718 14749 1738
rect 14769 1718 14776 1738
rect 14741 1713 14776 1718
rect 14741 1712 14773 1713
rect 13746 1685 14158 1693
rect 13746 1659 13752 1685
rect 13778 1659 14158 1685
rect 13746 1657 14158 1659
rect 13748 1656 13788 1657
rect 14126 1592 14158 1657
rect 16637 1697 16669 1762
rect 17007 1697 17047 1698
rect 16637 1695 17049 1697
rect 16637 1669 17017 1695
rect 17043 1669 17049 1695
rect 16637 1661 17049 1669
rect 16637 1633 16669 1661
rect 16637 1613 16642 1633
rect 16663 1613 16669 1633
rect 16637 1606 16669 1613
rect 16837 1633 16887 1642
rect 17082 1641 17116 1847
rect 17650 1867 17682 1895
rect 17650 1847 17655 1867
rect 17676 1847 17682 1867
rect 17650 1840 17682 1847
rect 17857 1868 17899 1876
rect 18095 1875 18129 2081
rect 17857 1848 17866 1868
rect 17890 1848 17899 1868
rect 17857 1836 17899 1848
rect 18073 1870 18129 1875
rect 18073 1850 18080 1870
rect 18100 1850 18129 1870
rect 18073 1843 18129 1850
rect 18073 1842 18108 1843
rect 17859 1807 17894 1836
rect 17859 1806 18169 1807
rect 17744 1800 17780 1804
rect 17744 1781 17752 1800
rect 17772 1781 17780 1800
rect 17744 1778 17780 1781
rect 17745 1750 17779 1778
rect 17859 1772 18186 1806
rect 16837 1612 16849 1633
rect 16871 1612 16887 1633
rect 16837 1604 16887 1612
rect 17060 1636 17116 1641
rect 17060 1616 17067 1636
rect 17087 1616 17116 1636
rect 17060 1609 17116 1616
rect 17217 1722 17780 1750
rect 17060 1608 17095 1609
rect 14126 1572 14130 1592
rect 14151 1572 14158 1592
rect 14126 1565 14158 1572
rect 16842 1571 16883 1604
rect 17217 1571 17257 1722
rect 16842 1542 17257 1571
rect 18146 1548 18186 1772
rect 18798 1790 18833 2384
rect 19882 2265 19922 2416
rect 20256 2383 20297 2416
rect 20044 2378 20079 2379
rect 19359 2237 19922 2265
rect 20023 2371 20079 2378
rect 20023 2351 20052 2371
rect 20072 2351 20079 2371
rect 20023 2346 20079 2351
rect 20252 2375 20302 2383
rect 20252 2354 20268 2375
rect 20290 2354 20302 2375
rect 18938 2210 19285 2214
rect 18938 2184 18947 2210
rect 18966 2184 19285 2210
rect 19360 2209 19394 2237
rect 18938 2179 19285 2184
rect 19359 2206 19395 2209
rect 19359 2187 19367 2206
rect 19387 2187 19395 2206
rect 19359 2183 19395 2187
rect 19245 2149 19285 2179
rect 19031 2144 19066 2145
rect 19010 2137 19066 2144
rect 19010 2117 19039 2137
rect 19059 2117 19066 2137
rect 19010 2112 19066 2117
rect 19242 2138 19285 2149
rect 19242 2118 19250 2138
rect 19274 2132 19285 2138
rect 19457 2140 19489 2147
rect 19274 2118 19284 2132
rect 19010 1906 19044 2112
rect 19242 2109 19284 2118
rect 19457 2120 19463 2140
rect 19484 2120 19489 2140
rect 19457 2092 19489 2120
rect 20023 2140 20057 2346
rect 20252 2345 20302 2354
rect 20470 2374 20502 2381
rect 20470 2354 20476 2374
rect 20497 2354 20502 2374
rect 20470 2326 20502 2354
rect 20090 2318 20502 2326
rect 20090 2292 20096 2318
rect 20122 2292 20502 2318
rect 20090 2290 20502 2292
rect 20092 2289 20132 2290
rect 20470 2225 20502 2290
rect 20470 2205 20474 2225
rect 20495 2205 20502 2225
rect 20470 2198 20502 2205
rect 20023 2132 20058 2140
rect 20023 2112 20031 2132
rect 20051 2112 20058 2132
rect 20023 2107 20058 2112
rect 20023 2106 20055 2107
rect 19077 2084 19489 2092
rect 19077 2058 19083 2084
rect 19109 2058 19489 2084
rect 19077 2056 19489 2058
rect 19079 2055 19119 2056
rect 19457 1991 19489 2056
rect 19457 1971 19461 1991
rect 19482 1971 19489 1991
rect 19457 1964 19489 1971
rect 19934 2002 20286 2033
rect 19010 1898 19045 1906
rect 19010 1878 19018 1898
rect 19038 1878 19045 1898
rect 19010 1862 19045 1878
rect 19934 1862 19965 2002
rect 20258 1970 20286 2002
rect 20043 1963 20078 1964
rect 19008 1843 19965 1862
rect 20022 1956 20078 1963
rect 20022 1936 20051 1956
rect 20071 1936 20078 1956
rect 20022 1931 20078 1936
rect 20252 1958 20292 1970
rect 20252 1937 20258 1958
rect 20280 1937 20292 1958
rect 20252 1932 20292 1937
rect 20469 1959 20501 1966
rect 20469 1939 20475 1959
rect 20496 1939 20501 1959
rect 18798 1761 19228 1790
rect 18798 1756 18882 1761
rect 18981 1724 19016 1725
rect 16842 1541 17251 1542
rect 18146 1528 18156 1548
rect 18176 1528 18186 1548
rect 18146 1518 18186 1528
rect 18960 1717 19016 1724
rect 18960 1697 18989 1717
rect 19009 1697 19016 1717
rect 18960 1692 19016 1697
rect 19190 1718 19228 1761
rect 19190 1701 19195 1718
rect 19219 1701 19228 1718
rect 12424 1307 12429 1327
rect 12450 1307 12456 1327
rect 12424 1300 12456 1307
rect 12635 1327 12672 1333
rect 12635 1308 12641 1327
rect 12664 1308 12672 1327
rect 12635 1303 12672 1308
rect 12847 1330 12903 1335
rect 12847 1310 12854 1330
rect 12874 1310 12903 1330
rect 12847 1303 12903 1310
rect 13677 1499 13717 1509
rect 13677 1479 13687 1499
rect 13707 1479 13717 1499
rect 14612 1485 15021 1486
rect 12643 1266 12667 1303
rect 12847 1302 12882 1303
rect 12643 1264 13011 1266
rect 12643 1259 13016 1264
rect 12643 1241 12989 1259
rect 13009 1241 13016 1259
rect 12643 1236 13016 1241
rect 12987 1234 13016 1236
rect 13677 1255 13717 1479
rect 14606 1456 15021 1485
rect 14606 1305 14646 1456
rect 14980 1423 15021 1456
rect 17705 1455 17737 1462
rect 17705 1435 17712 1455
rect 17733 1435 17737 1455
rect 14768 1418 14803 1419
rect 14083 1277 14646 1305
rect 14747 1411 14803 1418
rect 14747 1391 14776 1411
rect 14796 1391 14803 1411
rect 14747 1386 14803 1391
rect 14976 1415 15026 1423
rect 14976 1394 14992 1415
rect 15014 1394 15026 1415
rect 13677 1221 14004 1255
rect 14084 1249 14118 1277
rect 14083 1246 14119 1249
rect 14083 1227 14091 1246
rect 14111 1227 14119 1246
rect 14083 1223 14119 1227
rect 13694 1220 14004 1221
rect 13969 1191 14004 1220
rect 13755 1184 13790 1185
rect 11362 1068 11367 1088
rect 11388 1068 11394 1088
rect 11362 1061 11394 1068
rect 11571 1090 11611 1095
rect 11571 1069 11583 1090
rect 11605 1069 11611 1090
rect 11571 1057 11611 1069
rect 11785 1091 11841 1096
rect 11785 1071 11792 1091
rect 11812 1071 11841 1091
rect 11785 1064 11841 1071
rect 11898 1165 12855 1184
rect 13734 1177 13790 1184
rect 11785 1063 11820 1064
rect 8801 982 8805 1002
rect 8826 982 8833 1002
rect 8801 975 8833 982
rect 9278 1013 9630 1044
rect 8354 909 8389 917
rect 8354 889 8362 909
rect 8382 889 8389 909
rect 8354 873 8389 889
rect 9278 873 9309 1013
rect 9602 981 9630 1013
rect 11577 1025 11605 1057
rect 11898 1025 11929 1165
rect 12818 1149 12853 1165
rect 12818 1129 12825 1149
rect 12845 1129 12853 1149
rect 12818 1121 12853 1129
rect 11577 994 11929 1025
rect 12374 1056 12406 1063
rect 12374 1036 12381 1056
rect 12402 1036 12406 1056
rect 9387 974 9422 975
rect 7417 854 7473 861
rect 8352 854 9309 873
rect 9366 967 9422 974
rect 9366 947 9395 967
rect 9415 947 9422 967
rect 9366 942 9422 947
rect 9596 969 9636 981
rect 9596 948 9602 969
rect 9624 948 9636 969
rect 9596 943 9636 948
rect 9813 970 9845 977
rect 9813 950 9819 970
rect 9840 950 9845 970
rect 7417 853 7452 854
rect 7198 819 7238 849
rect 7088 811 7124 815
rect 7088 792 7096 811
rect 7116 792 7124 811
rect 7088 789 7124 792
rect 7198 814 7545 819
rect 7089 761 7123 789
rect 7198 788 7517 814
rect 7536 788 7545 814
rect 7198 784 7545 788
rect 6181 623 6193 644
rect 6215 623 6231 644
rect 6181 615 6231 623
rect 6404 647 6460 652
rect 6404 627 6411 647
rect 6431 627 6460 647
rect 6404 620 6460 627
rect 6561 733 7124 761
rect 9366 736 9400 942
rect 9813 922 9845 950
rect 9433 914 9845 922
rect 12374 971 12406 1036
rect 12744 971 12784 972
rect 12374 969 12786 971
rect 12374 943 12754 969
rect 12780 943 12786 969
rect 12374 935 12786 943
rect 11808 920 11840 921
rect 9433 888 9439 914
rect 9465 888 9845 914
rect 9433 886 9845 888
rect 11805 915 11840 920
rect 11805 895 11812 915
rect 11832 895 11840 915
rect 11805 887 11840 895
rect 9435 885 9475 886
rect 9813 821 9845 886
rect 9813 801 9817 821
rect 9838 801 9845 821
rect 9813 794 9845 801
rect 11361 822 11393 829
rect 11361 802 11368 822
rect 11389 802 11393 822
rect 11361 737 11393 802
rect 11731 737 11771 738
rect 6404 619 6439 620
rect 905 574 1320 603
rect 6186 582 6227 615
rect 6561 582 6601 733
rect 9366 728 9401 736
rect 9366 708 9374 728
rect 9394 708 9401 728
rect 9366 703 9401 708
rect 11361 735 11773 737
rect 11361 709 11741 735
rect 11767 709 11773 735
rect 9366 702 9398 703
rect 11361 701 11773 709
rect 11361 673 11393 701
rect 11361 653 11366 673
rect 11387 653 11393 673
rect 11361 646 11393 653
rect 11561 673 11611 682
rect 11806 681 11840 887
rect 12374 907 12406 935
rect 12374 887 12379 907
rect 12400 887 12406 907
rect 12579 909 12621 918
rect 12819 915 12853 1121
rect 12579 895 12589 909
rect 12374 880 12406 887
rect 12578 889 12589 895
rect 12613 889 12621 909
rect 12578 878 12621 889
rect 12797 910 12853 915
rect 12797 890 12804 910
rect 12824 890 12853 910
rect 13734 1157 13763 1177
rect 13783 1157 13790 1177
rect 13734 1152 13790 1157
rect 13964 1179 14006 1191
rect 13964 1159 13973 1179
rect 13997 1159 14006 1179
rect 13734 946 13768 1152
rect 13964 1151 14006 1159
rect 14181 1180 14213 1187
rect 14181 1160 14187 1180
rect 14208 1160 14213 1180
rect 14181 1132 14213 1160
rect 14747 1180 14781 1386
rect 14976 1385 15026 1394
rect 15194 1414 15226 1421
rect 15194 1394 15200 1414
rect 15221 1394 15226 1414
rect 15194 1366 15226 1394
rect 14814 1358 15226 1366
rect 14814 1332 14820 1358
rect 14846 1332 15226 1358
rect 14814 1330 15226 1332
rect 14816 1329 14856 1330
rect 15194 1265 15226 1330
rect 17705 1370 17737 1435
rect 18075 1370 18115 1371
rect 17705 1368 18117 1370
rect 17705 1342 18085 1368
rect 18111 1342 18117 1368
rect 17705 1334 18117 1342
rect 17090 1314 17122 1315
rect 17087 1309 17122 1314
rect 17087 1289 17094 1309
rect 17114 1289 17122 1309
rect 17087 1281 17122 1289
rect 15194 1245 15198 1265
rect 15219 1245 15226 1265
rect 15194 1238 15226 1245
rect 16643 1216 16675 1223
rect 16643 1196 16650 1216
rect 16671 1196 16675 1216
rect 14747 1172 14782 1180
rect 14747 1152 14755 1172
rect 14775 1152 14782 1172
rect 14747 1147 14782 1152
rect 14747 1146 14779 1147
rect 13801 1124 14213 1132
rect 13801 1098 13807 1124
rect 13833 1098 14213 1124
rect 13801 1096 14213 1098
rect 13803 1095 13843 1096
rect 14181 1031 14213 1096
rect 16643 1131 16675 1196
rect 17013 1131 17053 1132
rect 16643 1129 17055 1131
rect 16643 1103 17023 1129
rect 17049 1103 17055 1129
rect 16643 1095 17055 1103
rect 14181 1011 14185 1031
rect 14206 1011 14213 1031
rect 14181 1004 14213 1011
rect 14658 1042 15010 1073
rect 13734 938 13769 946
rect 13734 918 13742 938
rect 13762 918 13769 938
rect 13734 902 13769 918
rect 14658 902 14689 1042
rect 14982 1010 15010 1042
rect 16643 1067 16675 1095
rect 17088 1075 17122 1281
rect 17705 1306 17737 1334
rect 18150 1314 18184 1518
rect 18960 1488 18994 1692
rect 19190 1689 19228 1701
rect 19407 1720 19439 1727
rect 19407 1700 19413 1720
rect 19434 1700 19439 1720
rect 19407 1672 19439 1700
rect 20022 1725 20056 1931
rect 20469 1911 20501 1939
rect 20089 1903 20501 1911
rect 20089 1877 20095 1903
rect 20121 1877 20501 1903
rect 20089 1875 20501 1877
rect 20091 1874 20131 1875
rect 20469 1810 20501 1875
rect 20469 1790 20473 1810
rect 20494 1790 20501 1810
rect 20469 1783 20501 1790
rect 20022 1717 20057 1725
rect 20022 1697 20030 1717
rect 20050 1697 20057 1717
rect 20022 1692 20057 1697
rect 20022 1691 20054 1692
rect 19027 1664 19439 1672
rect 19027 1638 19033 1664
rect 19059 1638 19439 1664
rect 19027 1636 19439 1638
rect 19029 1635 19069 1636
rect 19407 1571 19439 1636
rect 19407 1551 19411 1571
rect 19432 1551 19439 1571
rect 19407 1544 19439 1551
rect 17705 1286 17710 1306
rect 17731 1286 17737 1306
rect 17705 1279 17737 1286
rect 17916 1306 17953 1312
rect 17916 1287 17922 1306
rect 17945 1287 17953 1306
rect 17916 1282 17953 1287
rect 18128 1309 18184 1314
rect 18128 1289 18135 1309
rect 18155 1289 18184 1309
rect 18128 1282 18184 1289
rect 18958 1478 18998 1488
rect 18958 1458 18968 1478
rect 18988 1458 18998 1478
rect 19893 1464 20302 1465
rect 17924 1245 17948 1282
rect 18128 1281 18163 1282
rect 17924 1243 18292 1245
rect 17924 1238 18297 1243
rect 17924 1220 18270 1238
rect 18290 1220 18297 1238
rect 17924 1215 18297 1220
rect 18268 1213 18297 1215
rect 18958 1234 18998 1458
rect 19887 1435 20302 1464
rect 19887 1284 19927 1435
rect 20261 1402 20302 1435
rect 20049 1397 20084 1398
rect 19364 1256 19927 1284
rect 20028 1390 20084 1397
rect 20028 1370 20057 1390
rect 20077 1370 20084 1390
rect 20028 1365 20084 1370
rect 20257 1394 20307 1402
rect 20257 1373 20273 1394
rect 20295 1373 20307 1394
rect 18958 1200 19285 1234
rect 19365 1228 19399 1256
rect 19364 1225 19400 1228
rect 19364 1206 19372 1225
rect 19392 1206 19400 1225
rect 19364 1202 19400 1206
rect 18975 1199 19285 1200
rect 19250 1170 19285 1199
rect 19036 1163 19071 1164
rect 16643 1047 16648 1067
rect 16669 1047 16675 1067
rect 16643 1040 16675 1047
rect 16852 1069 16892 1074
rect 16852 1048 16864 1069
rect 16886 1048 16892 1069
rect 16852 1036 16892 1048
rect 17066 1070 17122 1075
rect 17066 1050 17073 1070
rect 17093 1050 17122 1070
rect 17066 1043 17122 1050
rect 17179 1144 18136 1163
rect 19015 1156 19071 1163
rect 17066 1042 17101 1043
rect 14767 1003 14802 1004
rect 12797 883 12853 890
rect 13732 883 14689 902
rect 14746 996 14802 1003
rect 14746 976 14775 996
rect 14795 976 14802 996
rect 14746 971 14802 976
rect 14976 998 15016 1010
rect 14976 977 14982 998
rect 15004 977 15016 998
rect 14976 972 15016 977
rect 15193 999 15225 1006
rect 15193 979 15199 999
rect 15220 979 15225 999
rect 12797 882 12832 883
rect 12578 848 12618 878
rect 12468 840 12504 844
rect 12468 821 12476 840
rect 12496 821 12504 840
rect 12468 818 12504 821
rect 12578 843 12925 848
rect 12469 790 12503 818
rect 12578 817 12897 843
rect 12916 817 12925 843
rect 12578 813 12925 817
rect 11561 652 11573 673
rect 11595 652 11611 673
rect 11561 644 11611 652
rect 11784 676 11840 681
rect 11784 656 11791 676
rect 11811 656 11840 676
rect 11784 649 11840 656
rect 11941 762 12504 790
rect 14746 765 14780 971
rect 15193 951 15225 979
rect 16858 1004 16886 1036
rect 17179 1004 17210 1144
rect 18099 1128 18134 1144
rect 18099 1108 18106 1128
rect 18126 1108 18134 1128
rect 18099 1100 18134 1108
rect 16858 973 17210 1004
rect 17655 1035 17687 1042
rect 17655 1015 17662 1035
rect 17683 1015 17687 1035
rect 14813 943 15225 951
rect 14813 917 14819 943
rect 14845 917 15225 943
rect 14813 915 15225 917
rect 14815 914 14855 915
rect 15193 850 15225 915
rect 17655 950 17687 1015
rect 18025 950 18065 951
rect 17655 948 18067 950
rect 17655 922 18035 948
rect 18061 922 18067 948
rect 17655 914 18067 922
rect 17089 899 17121 900
rect 17086 894 17121 899
rect 17086 874 17093 894
rect 17113 874 17121 894
rect 17086 866 17121 874
rect 15193 830 15197 850
rect 15218 830 15225 850
rect 15193 823 15225 830
rect 16642 801 16674 808
rect 16642 781 16649 801
rect 16670 781 16674 801
rect 11784 648 11819 649
rect 905 573 1314 574
rect 6186 553 6601 582
rect 11566 611 11607 644
rect 11941 611 11981 762
rect 14746 757 14781 765
rect 14746 737 14754 757
rect 14774 737 14781 757
rect 14746 732 14781 737
rect 14746 731 14778 732
rect 16642 716 16674 781
rect 17012 716 17052 717
rect 16642 714 17054 716
rect 16642 688 17022 714
rect 17048 688 17054 714
rect 16642 680 17054 688
rect 16642 652 16674 680
rect 16642 632 16647 652
rect 16668 632 16674 652
rect 16642 625 16674 632
rect 16842 652 16892 661
rect 17087 660 17121 866
rect 17655 886 17687 914
rect 17655 866 17660 886
rect 17681 866 17687 886
rect 17860 888 17902 897
rect 18100 894 18134 1100
rect 17860 874 17870 888
rect 17655 859 17687 866
rect 17859 868 17870 874
rect 17894 868 17902 888
rect 17859 857 17902 868
rect 18078 889 18134 894
rect 18078 869 18085 889
rect 18105 869 18134 889
rect 19015 1136 19044 1156
rect 19064 1136 19071 1156
rect 19015 1131 19071 1136
rect 19245 1158 19287 1170
rect 19245 1138 19254 1158
rect 19278 1138 19287 1158
rect 19015 925 19049 1131
rect 19245 1130 19287 1138
rect 19462 1159 19494 1166
rect 19462 1139 19468 1159
rect 19489 1139 19494 1159
rect 19462 1111 19494 1139
rect 20028 1159 20062 1365
rect 20257 1364 20307 1373
rect 20475 1393 20507 1400
rect 20475 1373 20481 1393
rect 20502 1373 20507 1393
rect 20475 1345 20507 1373
rect 20095 1337 20507 1345
rect 20095 1311 20101 1337
rect 20127 1311 20507 1337
rect 20095 1309 20507 1311
rect 20097 1308 20137 1309
rect 20475 1244 20507 1309
rect 20475 1224 20479 1244
rect 20500 1224 20507 1244
rect 20475 1217 20507 1224
rect 20028 1151 20063 1159
rect 20028 1131 20036 1151
rect 20056 1131 20063 1151
rect 20028 1126 20063 1131
rect 20028 1125 20060 1126
rect 19082 1103 19494 1111
rect 19082 1077 19088 1103
rect 19114 1077 19494 1103
rect 19082 1075 19494 1077
rect 19084 1074 19124 1075
rect 19462 1010 19494 1075
rect 19462 990 19466 1010
rect 19487 990 19494 1010
rect 19462 983 19494 990
rect 19939 1021 20291 1052
rect 19015 917 19050 925
rect 19015 897 19023 917
rect 19043 897 19050 917
rect 19015 881 19050 897
rect 19939 881 19970 1021
rect 20263 989 20291 1021
rect 20048 982 20083 983
rect 18078 862 18134 869
rect 19013 862 19970 881
rect 20027 975 20083 982
rect 20027 955 20056 975
rect 20076 955 20083 975
rect 20027 950 20083 955
rect 20257 977 20297 989
rect 20257 956 20263 977
rect 20285 956 20297 977
rect 20257 951 20297 956
rect 20474 978 20506 985
rect 20474 958 20480 978
rect 20501 958 20506 978
rect 18078 861 18113 862
rect 17859 827 17899 857
rect 17749 819 17785 823
rect 17749 800 17757 819
rect 17777 800 17785 819
rect 17749 797 17785 800
rect 17859 822 18206 827
rect 17750 769 17784 797
rect 17859 796 18178 822
rect 18197 796 18206 822
rect 17859 792 18206 796
rect 16842 631 16854 652
rect 16876 631 16892 652
rect 16842 623 16892 631
rect 17065 655 17121 660
rect 17065 635 17072 655
rect 17092 635 17121 655
rect 17065 628 17121 635
rect 17222 741 17785 769
rect 20027 744 20061 950
rect 20474 930 20506 958
rect 20094 922 20506 930
rect 20094 896 20100 922
rect 20126 896 20506 922
rect 20094 894 20506 896
rect 20096 893 20136 894
rect 20474 829 20506 894
rect 20474 809 20478 829
rect 20499 809 20506 829
rect 20474 802 20506 809
rect 17065 627 17100 628
rect 11566 582 11981 611
rect 16847 590 16888 623
rect 17222 590 17262 741
rect 20027 736 20062 744
rect 20027 716 20035 736
rect 20055 716 20062 736
rect 20027 711 20062 716
rect 20027 710 20059 711
rect 11566 581 11975 582
rect 16847 561 17262 590
rect 16847 560 17256 561
rect 11408 553 11448 558
rect 6186 552 6595 553
rect 11355 550 15780 553
rect 747 545 787 550
rect 694 542 5119 545
rect 694 520 756 542
rect 779 520 5089 542
rect 5112 520 5119 542
rect 6028 524 6068 529
rect 11355 528 11417 550
rect 11440 528 15750 550
rect 15773 528 15780 550
rect 16689 532 16729 537
rect 694 515 5119 520
rect 5975 521 10400 524
rect 11355 523 15780 528
rect 16636 529 21061 532
rect 747 505 787 515
rect 5975 499 6037 521
rect 6060 499 10370 521
rect 10393 499 10400 521
rect 11408 513 11448 523
rect 16636 507 16698 529
rect 16721 507 21031 529
rect 21054 507 21061 529
rect 16636 502 21061 507
rect 5975 494 10400 499
rect 6028 484 6068 494
rect 16689 492 16729 502
rect 13204 481 13253 485
rect 13204 480 13214 481
rect 2543 473 2592 477
rect 2543 472 2553 473
rect 2543 443 2552 472
rect 2584 443 2592 473
rect 2543 442 2592 443
rect 2542 434 2592 442
rect 2542 426 2591 434
rect 2542 406 2554 426
rect 2574 406 2591 426
rect 2542 399 2591 406
rect 2646 425 2694 428
rect 2547 398 2582 399
rect 2103 333 2135 340
rect 2103 313 2110 333
rect 2131 313 2135 333
rect 2103 248 2135 313
rect 2473 248 2513 249
rect 2103 246 2515 248
rect 2103 220 2483 246
rect 2509 220 2515 246
rect 2103 212 2515 220
rect 2103 184 2135 212
rect 2548 192 2582 398
rect 2646 398 2649 425
rect 2684 398 2694 425
rect 2646 331 2694 398
rect 2646 311 2651 331
rect 2679 311 2694 331
rect 2646 301 2694 311
rect 2775 418 2811 463
rect 7824 452 7873 456
rect 7824 451 7834 452
rect 5636 418 5672 424
rect 7824 422 7833 451
rect 7865 422 7873 452
rect 13204 451 13213 480
rect 13245 451 13253 481
rect 13204 450 13253 451
rect 7824 421 7873 422
rect 2775 390 5672 418
rect 2103 164 2108 184
rect 2129 164 2135 184
rect 2103 157 2135 164
rect 2311 184 2355 191
rect 2311 162 2322 184
rect 2347 162 2355 184
rect 2311 154 2355 162
rect 2526 187 2582 192
rect 2526 167 2533 187
rect 2553 167 2582 187
rect 2526 160 2582 167
rect 2526 159 2561 160
rect 2317 124 2342 154
rect 2775 126 2813 390
rect 5636 338 5672 390
rect 7823 413 7873 421
rect 13203 442 13253 450
rect 13203 434 13252 442
rect 13203 414 13215 434
rect 13235 414 13252 434
rect 7823 405 7872 413
rect 13203 407 13252 414
rect 13307 433 13355 436
rect 7823 385 7835 405
rect 7855 385 7872 405
rect 7823 378 7872 385
rect 7927 404 7975 407
rect 13208 406 13243 407
rect 7828 377 7863 378
rect 5636 318 5644 338
rect 5664 318 5672 338
rect 5636 315 5672 318
rect 5637 310 5672 315
rect 5193 245 5225 252
rect 5193 225 5200 245
rect 5221 225 5225 245
rect 5193 160 5225 225
rect 5563 160 5603 161
rect 5193 158 5605 160
rect 5193 132 5573 158
rect 5599 132 5605 158
rect 2725 124 2814 126
rect 2317 91 2814 124
rect 2725 87 2814 91
rect 5193 124 5605 132
rect 5193 96 5225 124
rect 5638 104 5672 310
rect 7384 312 7416 319
rect 7384 292 7391 312
rect 7412 292 7416 312
rect 7384 227 7416 292
rect 7754 227 7794 228
rect 7384 225 7796 227
rect 7384 199 7764 225
rect 7790 199 7796 225
rect 7384 191 7796 199
rect 7384 163 7416 191
rect 7829 171 7863 377
rect 7927 377 7930 404
rect 7965 377 7975 404
rect 7927 310 7975 377
rect 9892 345 10934 374
rect 7927 290 7932 310
rect 7960 290 7975 310
rect 7927 280 7975 290
rect 7384 143 7389 163
rect 7410 143 7416 163
rect 7384 136 7416 143
rect 7592 163 7636 170
rect 7592 141 7603 163
rect 7628 141 7636 163
rect 7592 133 7636 141
rect 7807 166 7863 171
rect 7807 146 7814 166
rect 7834 146 7863 166
rect 7807 139 7863 146
rect 7807 138 7842 139
rect 5193 76 5198 96
rect 5219 76 5225 96
rect 5193 69 5225 76
rect 5399 93 5444 102
rect 5399 76 5409 93
rect 5430 76 5444 93
rect 5399 49 5444 76
rect 5616 99 5672 104
rect 5616 79 5623 99
rect 5643 79 5672 99
rect 5616 72 5672 79
rect 7598 104 7623 133
rect 7598 73 7622 104
rect 6914 72 7622 73
rect 5616 71 5651 72
rect 5796 71 7622 72
rect 5397 9 5444 49
rect 5787 70 7622 71
rect 5787 51 7621 70
rect 5787 40 6959 51
rect 5787 34 5834 40
rect 5395 5 5444 9
rect 5650 26 5834 34
rect 5650 9 5659 26
rect 5683 9 5834 26
rect 5395 -25 5443 5
rect 5650 1 5834 9
rect 5650 0 5833 1
rect 5395 -42 5441 -25
rect 9894 -42 9922 345
rect 10897 331 10934 345
rect 10897 311 10905 331
rect 10925 311 10934 331
rect 10897 281 10934 311
rect 12764 341 12796 348
rect 12764 321 12771 341
rect 12792 321 12796 341
rect 10454 238 10486 245
rect 10454 218 10461 238
rect 10482 218 10486 238
rect 10454 153 10486 218
rect 10824 153 10864 154
rect 10454 151 10866 153
rect 10454 125 10834 151
rect 10860 125 10866 151
rect 10454 117 10866 125
rect 10454 89 10486 117
rect 10454 69 10459 89
rect 10480 69 10486 89
rect 10454 62 10486 69
rect 10659 91 10709 99
rect 10899 97 10933 281
rect 12764 256 12796 321
rect 13134 256 13174 257
rect 12764 254 13176 256
rect 12764 228 13144 254
rect 13170 228 13176 254
rect 12764 220 13176 228
rect 12764 192 12796 220
rect 13209 200 13243 406
rect 13307 406 13310 433
rect 13345 406 13355 433
rect 13307 339 13355 406
rect 13307 319 13312 339
rect 13340 319 13355 339
rect 13307 309 13355 319
rect 13436 426 13472 471
rect 18485 460 18534 464
rect 18485 459 18495 460
rect 16297 426 16333 432
rect 18485 430 18494 459
rect 18526 430 18534 460
rect 18485 429 18534 430
rect 13436 398 16333 426
rect 12764 172 12769 192
rect 12790 172 12796 192
rect 12764 165 12796 172
rect 12972 192 13016 199
rect 12972 170 12983 192
rect 13008 170 13016 192
rect 12972 162 13016 170
rect 13187 195 13243 200
rect 13187 175 13194 195
rect 13214 175 13243 195
rect 13187 168 13243 175
rect 13187 167 13222 168
rect 12978 132 13003 162
rect 13436 134 13474 398
rect 16297 346 16333 398
rect 18484 421 18534 429
rect 18484 413 18533 421
rect 18484 393 18496 413
rect 18516 393 18533 413
rect 18484 386 18533 393
rect 18588 412 18636 415
rect 18489 385 18524 386
rect 16297 326 16305 346
rect 16325 326 16333 346
rect 16297 323 16333 326
rect 16298 318 16333 323
rect 15854 253 15886 260
rect 15854 233 15861 253
rect 15882 233 15886 253
rect 15854 168 15886 233
rect 16224 168 16264 169
rect 15854 166 16266 168
rect 15854 140 16234 166
rect 16260 140 16266 166
rect 13386 132 13475 134
rect 12978 99 13475 132
rect 10659 68 10668 91
rect 10696 68 10709 91
rect 10659 58 10709 68
rect 10877 92 10933 97
rect 13386 95 13475 99
rect 15854 132 16266 140
rect 15854 104 15886 132
rect 16299 112 16333 318
rect 18045 320 18077 327
rect 18045 300 18052 320
rect 18073 300 18077 320
rect 18045 235 18077 300
rect 18415 235 18455 236
rect 18045 233 18457 235
rect 18045 207 18425 233
rect 18451 207 18457 233
rect 18045 199 18457 207
rect 18045 171 18077 199
rect 18490 179 18524 385
rect 18588 385 18591 412
rect 18626 385 18636 412
rect 18588 318 18636 385
rect 18588 298 18593 318
rect 18621 298 18636 318
rect 18588 288 18636 298
rect 18045 151 18050 171
rect 18071 151 18077 171
rect 18045 144 18077 151
rect 18253 171 18297 178
rect 18253 149 18264 171
rect 18289 149 18297 171
rect 18253 141 18297 149
rect 18468 174 18524 179
rect 18468 154 18475 174
rect 18495 154 18524 174
rect 18468 147 18524 154
rect 18468 146 18503 147
rect 10877 72 10884 92
rect 10904 72 10933 92
rect 15854 84 15859 104
rect 15880 84 15886 104
rect 15854 77 15886 84
rect 16060 101 16105 110
rect 16060 84 16070 101
rect 16091 84 16105 101
rect 10877 65 10933 72
rect 10877 64 10912 65
rect 5395 -65 9929 -42
rect 10660 -58 10692 58
rect 16060 47 16105 84
rect 16277 107 16333 112
rect 16277 87 16284 107
rect 16304 87 16333 107
rect 16277 80 16333 87
rect 18259 112 18284 141
rect 18259 81 18283 112
rect 17575 80 18283 81
rect 16277 79 16312 80
rect 16457 79 18283 80
rect 16057 13 16105 47
rect 16448 78 18283 79
rect 16448 59 18282 78
rect 16448 48 17620 59
rect 16448 42 16495 48
rect 16311 34 16495 42
rect 16311 17 16320 34
rect 16344 17 16495 34
rect 10920 -14 10951 -6
rect 10912 -20 10951 -14
rect 16057 -20 16103 13
rect 16311 9 16495 17
rect 16311 8 16494 9
rect 10912 -24 16104 -20
rect 10912 -45 10925 -24
rect 10945 -45 16104 -24
rect 10912 -49 16104 -45
rect 10912 -50 10951 -49
rect 10912 -57 10947 -50
rect 9894 -71 9922 -65
<< via1 >>
rect 2649 4700 2686 4730
rect 7930 4679 7967 4709
rect 2548 4179 2582 4207
rect 13310 4708 13347 4738
rect 7829 4158 7863 4186
rect 18591 4687 18628 4717
rect 13209 4187 13243 4215
rect 18490 4166 18524 4194
rect 13214 480 13245 481
rect 2553 472 2584 473
rect 2552 443 2584 472
rect 2649 398 2684 425
rect 7834 451 7865 452
rect 7833 422 7865 451
rect 13213 451 13245 480
rect 7930 377 7965 404
rect 13310 406 13345 433
rect 18495 459 18526 460
rect 18494 430 18526 459
rect 18591 385 18626 412
<< metal2 >>
rect 13305 4738 13354 4744
rect 2644 4730 2693 4736
rect 2644 4700 2649 4730
rect 2686 4700 2693 4730
rect 2542 4207 2587 4213
rect 2542 4179 2548 4207
rect 2582 4179 2587 4207
rect 2542 569 2587 4179
rect 2644 600 2693 4700
rect 7925 4709 7974 4715
rect 7925 4679 7930 4709
rect 7967 4679 7974 4709
rect 7823 4186 7868 4192
rect 7823 4158 7829 4186
rect 7863 4158 7868 4186
rect 2548 477 2586 569
rect 2543 473 2592 477
rect 2543 472 2553 473
rect 2543 443 2552 472
rect 2584 443 2592 473
rect 2543 434 2592 443
rect 2646 425 2692 600
rect 7823 548 7868 4158
rect 7925 579 7974 4679
rect 13305 4708 13310 4738
rect 13347 4708 13354 4738
rect 13203 4215 13248 4221
rect 13203 4187 13209 4215
rect 13243 4187 13248 4215
rect 7829 456 7867 548
rect 2646 398 2649 425
rect 2684 398 2692 425
rect 7824 452 7873 456
rect 7824 451 7834 452
rect 7824 422 7833 451
rect 7865 422 7873 452
rect 7824 413 7873 422
rect 2646 383 2692 398
rect 7927 404 7973 579
rect 13203 577 13248 4187
rect 13305 608 13354 4708
rect 18586 4717 18635 4723
rect 18586 4687 18591 4717
rect 18628 4687 18635 4717
rect 18484 4194 18529 4200
rect 18484 4166 18490 4194
rect 18524 4166 18529 4194
rect 13209 485 13247 577
rect 13204 481 13253 485
rect 13204 480 13214 481
rect 13204 451 13213 480
rect 13245 451 13253 481
rect 13204 442 13253 451
rect 7927 377 7930 404
rect 7965 377 7973 404
rect 13307 433 13353 608
rect 18484 556 18529 4166
rect 18586 587 18635 4687
rect 18490 464 18528 556
rect 13307 406 13310 433
rect 13345 406 13353 433
rect 18485 460 18534 464
rect 18485 459 18495 460
rect 18485 430 18494 459
rect 18526 430 18534 460
rect 18485 421 18534 430
rect 13307 391 13353 406
rect 18588 412 18634 587
rect 7927 362 7973 377
rect 18588 385 18591 412
rect 18626 385 18634 412
rect 18588 370 18634 385
<< labels >>
rlabel locali 304 8164 333 8170 1 vdd
rlabel locali 517 8161 546 8167 1 vdd
rlabel locali 250 7976 272 7991 1 d0
rlabel nwell 671 8131 694 8134 1 vdd
rlabel locali 301 7865 330 7871 1 gnd
rlabel locali 514 7865 543 7871 1 gnd
rlabel space 611 7860 640 7869 1 gnd
rlabel locali 303 7749 332 7755 1 vdd
rlabel locali 516 7746 545 7752 1 vdd
rlabel locali 249 7561 271 7576 1 d0
rlabel nwell 670 7716 693 7719 1 vdd
rlabel locali 300 7450 329 7456 1 gnd
rlabel locali 513 7450 542 7456 1 gnd
rlabel space 610 7445 639 7454 1 gnd
rlabel locali 1316 7983 1345 7989 1 vdd
rlabel locali 1529 7980 1558 7986 1 vdd
rlabel nwell 1683 7950 1706 7953 1 vdd
rlabel locali 1313 7684 1342 7690 1 gnd
rlabel locali 1526 7684 1555 7690 1 gnd
rlabel space 1623 7679 1652 7688 1 gnd
rlabel locali 1254 7794 1301 7815 1 d1
rlabel locali 116 8356 141 8365 1 vref
rlabel locali 309 7183 338 7189 1 vdd
rlabel locali 522 7180 551 7186 1 vdd
rlabel locali 255 6995 277 7010 1 d0
rlabel nwell 676 7150 699 7153 1 vdd
rlabel locali 306 6884 335 6890 1 gnd
rlabel locali 519 6884 548 6890 1 gnd
rlabel space 616 6879 645 6888 1 gnd
rlabel locali 308 6768 337 6774 1 vdd
rlabel locali 521 6765 550 6771 1 vdd
rlabel locali 254 6580 276 6595 1 d0
rlabel nwell 675 6735 698 6738 1 vdd
rlabel locali 305 6469 334 6475 1 gnd
rlabel locali 518 6469 547 6475 1 gnd
rlabel locali 1321 7002 1350 7008 1 vdd
rlabel locali 1534 6999 1563 7005 1 vdd
rlabel nwell 1688 6969 1711 6972 1 vdd
rlabel locali 1318 6703 1347 6709 1 gnd
rlabel locali 1531 6703 1560 6709 1 gnd
rlabel space 1628 6698 1657 6707 1 gnd
rlabel locali 1259 6813 1306 6834 1 d1
rlabel locali 1371 7422 1400 7428 1 vdd
rlabel locali 1584 7419 1613 7425 1 vdd
rlabel nwell 1738 7389 1761 7392 1 vdd
rlabel locali 1368 7123 1397 7129 1 gnd
rlabel locali 1581 7123 1610 7129 1 gnd
rlabel space 1678 7118 1707 7127 1 gnd
rlabel locali 1314 7234 1337 7249 1 d2
rlabel space 615 6464 644 6473 1 gnd
rlabel locali 1326 5274 1349 5289 1 d2
rlabel space 1690 5158 1719 5167 1 gnd
rlabel locali 1593 5163 1622 5169 1 gnd
rlabel locali 1380 5163 1409 5169 1 gnd
rlabel nwell 1750 5429 1773 5432 1 vdd
rlabel locali 1596 5459 1625 5465 1 vdd
rlabel locali 1383 5462 1412 5468 1 vdd
rlabel locali 1271 4853 1318 4874 1 d1
rlabel space 1640 4738 1669 4747 1 gnd
rlabel locali 1543 4743 1572 4749 1 gnd
rlabel locali 1330 4743 1359 4749 1 gnd
rlabel nwell 1700 5009 1723 5012 1 vdd
rlabel locali 1546 5039 1575 5045 1 vdd
rlabel locali 1333 5042 1362 5048 1 vdd
rlabel space 627 4504 656 4513 1 gnd
rlabel locali 530 4509 559 4515 1 gnd
rlabel locali 317 4509 346 4515 1 gnd
rlabel nwell 687 4775 710 4778 1 vdd
rlabel locali 266 4620 288 4635 1 d0
rlabel locali 533 4805 562 4811 1 vdd
rlabel locali 320 4808 349 4814 1 vdd
rlabel space 628 4919 657 4928 1 gnd
rlabel locali 531 4924 560 4930 1 gnd
rlabel locali 318 4924 347 4930 1 gnd
rlabel nwell 688 5190 711 5193 1 vdd
rlabel locali 267 5035 289 5050 1 d0
rlabel locali 534 5220 563 5226 1 vdd
rlabel locali 321 5223 350 5229 1 vdd
rlabel locali 1266 5834 1313 5855 1 d1
rlabel space 1635 5719 1664 5728 1 gnd
rlabel locali 1538 5724 1567 5730 1 gnd
rlabel locali 1325 5724 1354 5730 1 gnd
rlabel nwell 1695 5990 1718 5993 1 vdd
rlabel locali 1541 6020 1570 6026 1 vdd
rlabel locali 1328 6023 1357 6029 1 vdd
rlabel space 622 5485 651 5494 1 gnd
rlabel locali 525 5490 554 5496 1 gnd
rlabel locali 312 5490 341 5496 1 gnd
rlabel nwell 682 5756 705 5759 1 vdd
rlabel locali 261 5601 283 5616 1 d0
rlabel locali 528 5786 557 5792 1 vdd
rlabel locali 315 5789 344 5795 1 vdd
rlabel space 623 5900 652 5909 1 gnd
rlabel locali 526 5905 555 5911 1 gnd
rlabel locali 313 5905 342 5911 1 gnd
rlabel nwell 683 6171 706 6174 1 vdd
rlabel locali 262 6016 284 6031 1 d0
rlabel locali 529 6201 558 6207 1 vdd
rlabel locali 316 6204 345 6210 1 vdd
rlabel locali 1536 6490 1565 6496 1 vdd
rlabel locali 1749 6487 1778 6493 1 vdd
rlabel nwell 1903 6457 1926 6460 1 vdd
rlabel locali 1533 6191 1562 6197 1 gnd
rlabel locali 1746 6191 1775 6197 1 gnd
rlabel space 1843 6186 1872 6195 1 gnd
rlabel locali 1474 6300 1506 6319 1 d3
rlabel locali 1494 2383 1526 2402 1 d3
rlabel space 1863 2269 1892 2278 1 gnd
rlabel locali 1766 2274 1795 2280 1 gnd
rlabel locali 1553 2274 1582 2280 1 gnd
rlabel nwell 1923 2540 1946 2543 1 vdd
rlabel locali 1769 2570 1798 2576 1 vdd
rlabel locali 1556 2573 1585 2579 1 vdd
rlabel locali 336 2287 365 2293 1 vdd
rlabel locali 549 2284 578 2290 1 vdd
rlabel locali 282 2099 304 2114 1 d0
rlabel nwell 703 2254 726 2257 1 vdd
rlabel locali 333 1988 362 1994 1 gnd
rlabel locali 546 1988 575 1994 1 gnd
rlabel space 643 1983 672 1992 1 gnd
rlabel locali 335 1872 364 1878 1 vdd
rlabel locali 548 1869 577 1875 1 vdd
rlabel locali 281 1684 303 1699 1 d0
rlabel nwell 702 1839 725 1842 1 vdd
rlabel locali 332 1573 361 1579 1 gnd
rlabel locali 545 1573 574 1579 1 gnd
rlabel space 642 1568 671 1577 1 gnd
rlabel locali 1348 2106 1377 2112 1 vdd
rlabel locali 1561 2103 1590 2109 1 vdd
rlabel nwell 1715 2073 1738 2076 1 vdd
rlabel locali 1345 1807 1374 1813 1 gnd
rlabel locali 1558 1807 1587 1813 1 gnd
rlabel space 1655 1802 1684 1811 1 gnd
rlabel locali 1286 1917 1333 1938 1 d1
rlabel locali 341 1306 370 1312 1 vdd
rlabel locali 554 1303 583 1309 1 vdd
rlabel locali 287 1118 309 1133 1 d0
rlabel nwell 708 1273 731 1276 1 vdd
rlabel locali 338 1007 367 1013 1 gnd
rlabel locali 551 1007 580 1013 1 gnd
rlabel space 648 1002 677 1011 1 gnd
rlabel locali 340 891 369 897 1 vdd
rlabel locali 553 888 582 894 1 vdd
rlabel locali 286 703 308 718 1 d0
rlabel nwell 707 858 730 861 1 vdd
rlabel locali 337 592 366 598 1 gnd
rlabel locali 550 592 579 598 1 gnd
rlabel space 647 587 676 596 1 gnd
rlabel locali 1353 1125 1382 1131 1 vdd
rlabel locali 1566 1122 1595 1128 1 vdd
rlabel nwell 1720 1092 1743 1095 1 vdd
rlabel locali 1350 826 1379 832 1 gnd
rlabel locali 1563 826 1592 832 1 gnd
rlabel space 1660 821 1689 830 1 gnd
rlabel locali 1291 936 1338 957 1 d1
rlabel locali 1403 1545 1432 1551 1 vdd
rlabel locali 1616 1542 1645 1548 1 vdd
rlabel nwell 1770 1512 1793 1515 1 vdd
rlabel locali 1400 1246 1429 1252 1 gnd
rlabel locali 1613 1246 1642 1252 1 gnd
rlabel space 1710 1241 1739 1250 1 gnd
rlabel locali 1346 1357 1369 1372 1 d2
rlabel space 635 2547 664 2556 1 gnd
rlabel locali 1334 3317 1357 3332 1 d2
rlabel space 1698 3201 1727 3210 1 gnd
rlabel locali 1601 3206 1630 3212 1 gnd
rlabel locali 1388 3206 1417 3212 1 gnd
rlabel nwell 1758 3472 1781 3475 1 vdd
rlabel locali 1604 3502 1633 3508 1 vdd
rlabel locali 1391 3505 1420 3511 1 vdd
rlabel locali 1279 2896 1326 2917 1 d1
rlabel space 1648 2781 1677 2790 1 gnd
rlabel locali 1551 2786 1580 2792 1 gnd
rlabel locali 1338 2786 1367 2792 1 gnd
rlabel nwell 1708 3052 1731 3055 1 vdd
rlabel locali 1554 3082 1583 3088 1 vdd
rlabel locali 1341 3085 1370 3091 1 vdd
rlabel locali 538 2552 567 2558 1 gnd
rlabel locali 325 2552 354 2558 1 gnd
rlabel nwell 695 2818 718 2821 1 vdd
rlabel locali 274 2663 296 2678 1 d0
rlabel locali 541 2848 570 2854 1 vdd
rlabel locali 328 2851 357 2857 1 vdd
rlabel space 636 2962 665 2971 1 gnd
rlabel locali 539 2967 568 2973 1 gnd
rlabel locali 326 2967 355 2973 1 gnd
rlabel nwell 696 3233 719 3236 1 vdd
rlabel locali 275 3078 297 3093 1 d0
rlabel locali 542 3263 571 3269 1 vdd
rlabel locali 329 3266 358 3272 1 vdd
rlabel locali 1274 3877 1321 3898 1 d1
rlabel space 1643 3762 1672 3771 1 gnd
rlabel locali 1546 3767 1575 3773 1 gnd
rlabel locali 1333 3767 1362 3773 1 gnd
rlabel nwell 1703 4033 1726 4036 1 vdd
rlabel locali 1549 4063 1578 4069 1 vdd
rlabel locali 1336 4066 1365 4072 1 vdd
rlabel space 630 3528 659 3537 1 gnd
rlabel locali 533 3533 562 3539 1 gnd
rlabel locali 320 3533 349 3539 1 gnd
rlabel nwell 690 3799 713 3802 1 vdd
rlabel locali 269 3644 291 3659 1 d0
rlabel locali 536 3829 565 3835 1 vdd
rlabel locali 323 3832 352 3838 1 vdd
rlabel space 631 3943 660 3952 1 gnd
rlabel locali 534 3948 563 3954 1 gnd
rlabel locali 321 3948 350 3954 1 gnd
rlabel nwell 691 4214 714 4217 1 vdd
rlabel locali 270 4059 292 4074 1 d0
rlabel locali 537 4244 566 4250 1 vdd
rlabel locali 324 4247 353 4253 1 vdd
rlabel locali 1631 4498 1660 4504 1 vdd
rlabel locali 1844 4495 1873 4501 1 vdd
rlabel nwell 1998 4465 2021 4468 1 vdd
rlabel locali 1628 4199 1657 4205 1 gnd
rlabel locali 1841 4199 1870 4205 1 gnd
rlabel space 1938 4194 1967 4203 1 gnd
rlabel locali 1573 4304 1595 4328 1 d4
rlabel locali 4895 739 4924 745 5 vdd
rlabel locali 4682 742 4711 748 5 vdd
rlabel locali 4956 918 4978 933 5 d0
rlabel nwell 4534 775 4557 778 5 vdd
rlabel locali 4898 1038 4927 1044 5 gnd
rlabel locali 4685 1038 4714 1044 5 gnd
rlabel space 4588 1040 4617 1049 5 gnd
rlabel locali 4896 1154 4925 1160 5 vdd
rlabel locali 4683 1157 4712 1163 5 vdd
rlabel locali 4957 1333 4979 1348 5 d0
rlabel nwell 4535 1190 4558 1193 5 vdd
rlabel locali 4899 1453 4928 1459 5 gnd
rlabel locali 4686 1453 4715 1459 5 gnd
rlabel space 4589 1455 4618 1464 5 gnd
rlabel locali 3883 920 3912 926 5 vdd
rlabel locali 3670 923 3699 929 5 vdd
rlabel nwell 3522 956 3545 959 5 vdd
rlabel locali 3886 1219 3915 1225 5 gnd
rlabel locali 3673 1219 3702 1225 5 gnd
rlabel space 3576 1221 3605 1230 5 gnd
rlabel locali 3927 1094 3974 1115 5 d1
rlabel locali 4890 1720 4919 1726 5 vdd
rlabel locali 4677 1723 4706 1729 5 vdd
rlabel locali 4951 1899 4973 1914 5 d0
rlabel nwell 4529 1756 4552 1759 5 vdd
rlabel locali 4893 2019 4922 2025 5 gnd
rlabel locali 4680 2019 4709 2025 5 gnd
rlabel space 4583 2021 4612 2030 5 gnd
rlabel locali 4891 2135 4920 2141 5 vdd
rlabel locali 4678 2138 4707 2144 5 vdd
rlabel locali 4952 2314 4974 2329 5 d0
rlabel nwell 4530 2171 4553 2174 5 vdd
rlabel locali 4894 2434 4923 2440 5 gnd
rlabel locali 4681 2434 4710 2440 5 gnd
rlabel locali 3878 1901 3907 1907 5 vdd
rlabel locali 3665 1904 3694 1910 5 vdd
rlabel nwell 3517 1937 3540 1940 5 vdd
rlabel locali 3881 2200 3910 2206 5 gnd
rlabel locali 3668 2200 3697 2206 5 gnd
rlabel space 3571 2202 3600 2211 5 gnd
rlabel locali 3922 2075 3969 2096 5 d1
rlabel locali 3828 1481 3857 1487 5 vdd
rlabel locali 3615 1484 3644 1490 5 vdd
rlabel nwell 3467 1517 3490 1520 5 vdd
rlabel locali 3831 1780 3860 1786 5 gnd
rlabel locali 3618 1780 3647 1786 5 gnd
rlabel space 3521 1782 3550 1791 5 gnd
rlabel locali 3891 1660 3914 1675 5 d2
rlabel space 4584 2436 4613 2445 5 gnd
rlabel locali 3879 3620 3902 3635 5 d2
rlabel space 3509 3742 3538 3751 5 gnd
rlabel locali 3606 3740 3635 3746 5 gnd
rlabel locali 3819 3740 3848 3746 5 gnd
rlabel nwell 3455 3477 3478 3480 5 vdd
rlabel locali 3603 3444 3632 3450 5 vdd
rlabel locali 3816 3441 3845 3447 5 vdd
rlabel locali 3910 4035 3957 4056 5 d1
rlabel space 3559 4162 3588 4171 5 gnd
rlabel locali 3656 4160 3685 4166 5 gnd
rlabel locali 3869 4160 3898 4166 5 gnd
rlabel nwell 3505 3897 3528 3900 5 vdd
rlabel locali 3653 3864 3682 3870 5 vdd
rlabel locali 3866 3861 3895 3867 5 vdd
rlabel space 4572 4396 4601 4405 5 gnd
rlabel locali 4669 4394 4698 4400 5 gnd
rlabel locali 4882 4394 4911 4400 5 gnd
rlabel nwell 4518 4131 4541 4134 5 vdd
rlabel locali 4940 4274 4962 4289 5 d0
rlabel locali 4666 4098 4695 4104 5 vdd
rlabel locali 4879 4095 4908 4101 5 vdd
rlabel space 4571 3981 4600 3990 5 gnd
rlabel locali 4668 3979 4697 3985 5 gnd
rlabel locali 4881 3979 4910 3985 5 gnd
rlabel nwell 4517 3716 4540 3719 5 vdd
rlabel locali 4939 3859 4961 3874 5 d0
rlabel locali 4665 3683 4694 3689 5 vdd
rlabel locali 4878 3680 4907 3686 5 vdd
rlabel locali 3915 3054 3962 3075 5 d1
rlabel space 3564 3181 3593 3190 5 gnd
rlabel locali 3661 3179 3690 3185 5 gnd
rlabel locali 3874 3179 3903 3185 5 gnd
rlabel nwell 3510 2916 3533 2919 5 vdd
rlabel locali 3658 2883 3687 2889 5 vdd
rlabel locali 3871 2880 3900 2886 5 vdd
rlabel space 4577 3415 4606 3424 5 gnd
rlabel locali 4674 3413 4703 3419 5 gnd
rlabel locali 4887 3413 4916 3419 5 gnd
rlabel nwell 4523 3150 4546 3153 5 vdd
rlabel locali 4945 3293 4967 3308 5 d0
rlabel locali 4671 3117 4700 3123 5 vdd
rlabel locali 4884 3114 4913 3120 5 vdd
rlabel space 4576 3000 4605 3009 5 gnd
rlabel locali 4673 2998 4702 3004 5 gnd
rlabel locali 4886 2998 4915 3004 5 gnd
rlabel nwell 4522 2735 4545 2738 5 vdd
rlabel locali 4944 2878 4966 2893 5 d0
rlabel locali 4670 2702 4699 2708 5 vdd
rlabel locali 4883 2699 4912 2705 5 vdd
rlabel locali 3663 2413 3692 2419 5 vdd
rlabel locali 3450 2416 3479 2422 5 vdd
rlabel nwell 3302 2449 3325 2452 5 vdd
rlabel locali 3666 2712 3695 2718 5 gnd
rlabel locali 3453 2712 3482 2718 5 gnd
rlabel space 3356 2714 3385 2723 5 gnd
rlabel locali 3722 2590 3754 2609 5 d3
rlabel locali 3702 6507 3734 6526 5 d3
rlabel space 3336 6631 3365 6640 5 gnd
rlabel locali 3433 6629 3462 6635 5 gnd
rlabel locali 3646 6629 3675 6635 5 gnd
rlabel nwell 3282 6366 3305 6369 5 vdd
rlabel locali 3430 6333 3459 6339 5 vdd
rlabel locali 3643 6330 3672 6336 5 vdd
rlabel locali 4863 6616 4892 6622 5 vdd
rlabel locali 4650 6619 4679 6625 5 vdd
rlabel locali 4924 6795 4946 6810 5 d0
rlabel nwell 4502 6652 4525 6655 5 vdd
rlabel locali 4866 6915 4895 6921 5 gnd
rlabel locali 4653 6915 4682 6921 5 gnd
rlabel space 4556 6917 4585 6926 5 gnd
rlabel locali 4864 7031 4893 7037 5 vdd
rlabel locali 4651 7034 4680 7040 5 vdd
rlabel locali 4925 7210 4947 7225 5 d0
rlabel nwell 4503 7067 4526 7070 5 vdd
rlabel locali 4867 7330 4896 7336 5 gnd
rlabel locali 4654 7330 4683 7336 5 gnd
rlabel space 4557 7332 4586 7341 5 gnd
rlabel locali 3851 6797 3880 6803 5 vdd
rlabel locali 3638 6800 3667 6806 5 vdd
rlabel nwell 3490 6833 3513 6836 5 vdd
rlabel locali 3854 7096 3883 7102 5 gnd
rlabel locali 3641 7096 3670 7102 5 gnd
rlabel space 3544 7098 3573 7107 5 gnd
rlabel locali 3895 6971 3942 6992 5 d1
rlabel locali 4858 7597 4887 7603 5 vdd
rlabel locali 4645 7600 4674 7606 5 vdd
rlabel locali 4919 7776 4941 7791 5 d0
rlabel nwell 4497 7633 4520 7636 5 vdd
rlabel locali 4861 7896 4890 7902 5 gnd
rlabel locali 4648 7896 4677 7902 5 gnd
rlabel space 4551 7898 4580 7907 5 gnd
rlabel locali 4859 8012 4888 8018 5 vdd
rlabel locali 4646 8015 4675 8021 5 vdd
rlabel locali 4920 8191 4942 8206 5 d0
rlabel nwell 4498 8048 4521 8051 5 vdd
rlabel locali 4862 8311 4891 8317 5 gnd
rlabel locali 4649 8311 4678 8317 5 gnd
rlabel space 4552 8313 4581 8322 5 gnd
rlabel locali 3846 7778 3875 7784 5 vdd
rlabel locali 3633 7781 3662 7787 5 vdd
rlabel nwell 3485 7814 3508 7817 5 vdd
rlabel locali 3849 8077 3878 8083 5 gnd
rlabel locali 3636 8077 3665 8083 5 gnd
rlabel space 3539 8079 3568 8088 5 gnd
rlabel locali 3890 7952 3937 7973 5 d1
rlabel locali 3796 7358 3825 7364 5 vdd
rlabel locali 3583 7361 3612 7367 5 vdd
rlabel nwell 3435 7394 3458 7397 5 vdd
rlabel locali 3799 7657 3828 7663 5 gnd
rlabel locali 3586 7657 3615 7663 5 gnd
rlabel space 3489 7659 3518 7668 5 gnd
rlabel locali 3859 7537 3882 7552 5 d2
rlabel space 4564 6353 4593 6362 5 gnd
rlabel locali 3871 5577 3894 5592 5 d2
rlabel space 3501 5699 3530 5708 5 gnd
rlabel locali 3598 5697 3627 5703 5 gnd
rlabel locali 3811 5697 3840 5703 5 gnd
rlabel nwell 3447 5434 3470 5437 5 vdd
rlabel locali 3595 5401 3624 5407 5 vdd
rlabel locali 3808 5398 3837 5404 5 vdd
rlabel locali 3902 5992 3949 6013 5 d1
rlabel space 3551 6119 3580 6128 5 gnd
rlabel locali 3648 6117 3677 6123 5 gnd
rlabel locali 3861 6117 3890 6123 5 gnd
rlabel nwell 3497 5854 3520 5857 5 vdd
rlabel locali 3645 5821 3674 5827 5 vdd
rlabel locali 3858 5818 3887 5824 5 vdd
rlabel locali 4661 6351 4690 6357 5 gnd
rlabel locali 4874 6351 4903 6357 5 gnd
rlabel nwell 4510 6088 4533 6091 5 vdd
rlabel locali 4932 6231 4954 6246 5 d0
rlabel locali 4658 6055 4687 6061 5 vdd
rlabel locali 4871 6052 4900 6058 5 vdd
rlabel space 4563 5938 4592 5947 5 gnd
rlabel locali 4660 5936 4689 5942 5 gnd
rlabel locali 4873 5936 4902 5942 5 gnd
rlabel nwell 4509 5673 4532 5676 5 vdd
rlabel locali 4931 5816 4953 5831 5 d0
rlabel locali 4657 5640 4686 5646 5 vdd
rlabel locali 4870 5637 4899 5643 5 vdd
rlabel locali 3907 5011 3954 5032 5 d1
rlabel space 3556 5138 3585 5147 5 gnd
rlabel locali 3653 5136 3682 5142 5 gnd
rlabel locali 3866 5136 3895 5142 5 gnd
rlabel nwell 3502 4873 3525 4876 5 vdd
rlabel locali 3650 4840 3679 4846 5 vdd
rlabel locali 3863 4837 3892 4843 5 vdd
rlabel space 4569 5372 4598 5381 5 gnd
rlabel locali 4666 5370 4695 5376 5 gnd
rlabel locali 4879 5370 4908 5376 5 gnd
rlabel nwell 4515 5107 4538 5110 5 vdd
rlabel locali 4937 5250 4959 5265 5 d0
rlabel locali 4663 5074 4692 5080 5 vdd
rlabel locali 4876 5071 4905 5077 5 vdd
rlabel space 4568 4957 4597 4966 5 gnd
rlabel locali 4665 4955 4694 4961 5 gnd
rlabel locali 4878 4955 4907 4961 5 gnd
rlabel nwell 4514 4692 4537 4695 5 vdd
rlabel locali 4936 4835 4958 4850 5 d0
rlabel locali 4662 4659 4691 4665 5 vdd
rlabel locali 4875 4656 4904 4662 5 vdd
rlabel locali 3568 4405 3597 4411 5 vdd
rlabel locali 3355 4408 3384 4414 5 vdd
rlabel nwell 3207 4441 3230 4444 5 vdd
rlabel locali 3571 4704 3600 4710 5 gnd
rlabel locali 3358 4704 3387 4710 5 gnd
rlabel space 3261 4706 3290 4715 5 gnd
rlabel locali 3633 4581 3655 4605 5 d4
rlabel locali 1743 410 1772 416 1 vdd
rlabel locali 1956 407 1985 413 1 vdd
rlabel nwell 2110 377 2133 380 1 vdd
rlabel locali 1740 111 1769 117 1 gnd
rlabel locali 1953 111 1982 117 1 gnd
rlabel space 2050 106 2079 115 1 gnd
rlabel locali 1685 219 1709 236 1 d5
rlabel locali 5585 8143 5614 8149 1 vdd
rlabel locali 5798 8140 5827 8146 1 vdd
rlabel locali 5531 7955 5553 7970 1 d0
rlabel nwell 5952 8110 5975 8113 1 vdd
rlabel locali 5582 7844 5611 7850 1 gnd
rlabel locali 5795 7844 5824 7850 1 gnd
rlabel space 5892 7839 5921 7848 1 gnd
rlabel locali 5584 7728 5613 7734 1 vdd
rlabel locali 5797 7725 5826 7731 1 vdd
rlabel locali 5530 7540 5552 7555 1 d0
rlabel nwell 5951 7695 5974 7698 1 vdd
rlabel locali 5581 7429 5610 7435 1 gnd
rlabel locali 5794 7429 5823 7435 1 gnd
rlabel space 5891 7424 5920 7433 1 gnd
rlabel locali 6597 7962 6626 7968 1 vdd
rlabel locali 6810 7959 6839 7965 1 vdd
rlabel nwell 6964 7929 6987 7932 1 vdd
rlabel locali 6594 7663 6623 7669 1 gnd
rlabel locali 6807 7663 6836 7669 1 gnd
rlabel space 6904 7658 6933 7667 1 gnd
rlabel locali 6535 7773 6582 7794 1 d1
rlabel locali 5590 7162 5619 7168 1 vdd
rlabel locali 5803 7159 5832 7165 1 vdd
rlabel locali 5536 6974 5558 6989 1 d0
rlabel nwell 5957 7129 5980 7132 1 vdd
rlabel locali 5587 6863 5616 6869 1 gnd
rlabel locali 5800 6863 5829 6869 1 gnd
rlabel space 5897 6858 5926 6867 1 gnd
rlabel locali 5589 6747 5618 6753 1 vdd
rlabel locali 5802 6744 5831 6750 1 vdd
rlabel locali 5535 6559 5557 6574 1 d0
rlabel nwell 5956 6714 5979 6717 1 vdd
rlabel locali 5586 6448 5615 6454 1 gnd
rlabel locali 5799 6448 5828 6454 1 gnd
rlabel locali 6602 6981 6631 6987 1 vdd
rlabel locali 6815 6978 6844 6984 1 vdd
rlabel nwell 6969 6948 6992 6951 1 vdd
rlabel locali 6599 6682 6628 6688 1 gnd
rlabel locali 6812 6682 6841 6688 1 gnd
rlabel space 6909 6677 6938 6686 1 gnd
rlabel locali 6540 6792 6587 6813 1 d1
rlabel locali 6652 7401 6681 7407 1 vdd
rlabel locali 6865 7398 6894 7404 1 vdd
rlabel nwell 7019 7368 7042 7371 1 vdd
rlabel locali 6649 7102 6678 7108 1 gnd
rlabel locali 6862 7102 6891 7108 1 gnd
rlabel space 6959 7097 6988 7106 1 gnd
rlabel locali 6595 7213 6618 7228 1 d2
rlabel space 5896 6443 5925 6452 1 gnd
rlabel locali 6607 5253 6630 5268 1 d2
rlabel space 6971 5137 7000 5146 1 gnd
rlabel locali 6874 5142 6903 5148 1 gnd
rlabel locali 6661 5142 6690 5148 1 gnd
rlabel nwell 7031 5408 7054 5411 1 vdd
rlabel locali 6877 5438 6906 5444 1 vdd
rlabel locali 6664 5441 6693 5447 1 vdd
rlabel locali 6552 4832 6599 4853 1 d1
rlabel space 6921 4717 6950 4726 1 gnd
rlabel locali 6824 4722 6853 4728 1 gnd
rlabel locali 6611 4722 6640 4728 1 gnd
rlabel nwell 6981 4988 7004 4991 1 vdd
rlabel locali 6827 5018 6856 5024 1 vdd
rlabel locali 6614 5021 6643 5027 1 vdd
rlabel space 5908 4483 5937 4492 1 gnd
rlabel locali 5811 4488 5840 4494 1 gnd
rlabel locali 5598 4488 5627 4494 1 gnd
rlabel nwell 5968 4754 5991 4757 1 vdd
rlabel locali 5547 4599 5569 4614 1 d0
rlabel locali 5814 4784 5843 4790 1 vdd
rlabel locali 5601 4787 5630 4793 1 vdd
rlabel space 5909 4898 5938 4907 1 gnd
rlabel locali 5812 4903 5841 4909 1 gnd
rlabel locali 5599 4903 5628 4909 1 gnd
rlabel nwell 5969 5169 5992 5172 1 vdd
rlabel locali 5548 5014 5570 5029 1 d0
rlabel locali 5815 5199 5844 5205 1 vdd
rlabel locali 5602 5202 5631 5208 1 vdd
rlabel locali 6547 5813 6594 5834 1 d1
rlabel space 6916 5698 6945 5707 1 gnd
rlabel locali 6819 5703 6848 5709 1 gnd
rlabel locali 6606 5703 6635 5709 1 gnd
rlabel nwell 6976 5969 6999 5972 1 vdd
rlabel locali 6822 5999 6851 6005 1 vdd
rlabel locali 6609 6002 6638 6008 1 vdd
rlabel space 5903 5464 5932 5473 1 gnd
rlabel locali 5806 5469 5835 5475 1 gnd
rlabel locali 5593 5469 5622 5475 1 gnd
rlabel nwell 5963 5735 5986 5738 1 vdd
rlabel locali 5542 5580 5564 5595 1 d0
rlabel locali 5809 5765 5838 5771 1 vdd
rlabel locali 5596 5768 5625 5774 1 vdd
rlabel space 5904 5879 5933 5888 1 gnd
rlabel locali 5807 5884 5836 5890 1 gnd
rlabel locali 5594 5884 5623 5890 1 gnd
rlabel nwell 5964 6150 5987 6153 1 vdd
rlabel locali 5543 5995 5565 6010 1 d0
rlabel locali 5810 6180 5839 6186 1 vdd
rlabel locali 5597 6183 5626 6189 1 vdd
rlabel locali 6817 6469 6846 6475 1 vdd
rlabel locali 7030 6466 7059 6472 1 vdd
rlabel nwell 7184 6436 7207 6439 1 vdd
rlabel locali 6814 6170 6843 6176 1 gnd
rlabel locali 7027 6170 7056 6176 1 gnd
rlabel space 7124 6165 7153 6174 1 gnd
rlabel locali 6755 6279 6787 6298 1 d3
rlabel locali 6775 2362 6807 2381 1 d3
rlabel space 7144 2248 7173 2257 1 gnd
rlabel locali 7047 2253 7076 2259 1 gnd
rlabel locali 6834 2253 6863 2259 1 gnd
rlabel nwell 7204 2519 7227 2522 1 vdd
rlabel locali 7050 2549 7079 2555 1 vdd
rlabel locali 6837 2552 6866 2558 1 vdd
rlabel locali 5617 2266 5646 2272 1 vdd
rlabel locali 5830 2263 5859 2269 1 vdd
rlabel locali 5563 2078 5585 2093 1 d0
rlabel nwell 5984 2233 6007 2236 1 vdd
rlabel locali 5614 1967 5643 1973 1 gnd
rlabel locali 5827 1967 5856 1973 1 gnd
rlabel space 5924 1962 5953 1971 1 gnd
rlabel locali 5616 1851 5645 1857 1 vdd
rlabel locali 5829 1848 5858 1854 1 vdd
rlabel locali 5562 1663 5584 1678 1 d0
rlabel nwell 5983 1818 6006 1821 1 vdd
rlabel locali 5613 1552 5642 1558 1 gnd
rlabel locali 5826 1552 5855 1558 1 gnd
rlabel space 5923 1547 5952 1556 1 gnd
rlabel locali 6629 2085 6658 2091 1 vdd
rlabel locali 6842 2082 6871 2088 1 vdd
rlabel nwell 6996 2052 7019 2055 1 vdd
rlabel locali 6626 1786 6655 1792 1 gnd
rlabel locali 6839 1786 6868 1792 1 gnd
rlabel space 6936 1781 6965 1790 1 gnd
rlabel locali 6567 1896 6614 1917 1 d1
rlabel locali 5622 1285 5651 1291 1 vdd
rlabel locali 5835 1282 5864 1288 1 vdd
rlabel locali 5568 1097 5590 1112 1 d0
rlabel nwell 5989 1252 6012 1255 1 vdd
rlabel locali 5619 986 5648 992 1 gnd
rlabel locali 5832 986 5861 992 1 gnd
rlabel space 5929 981 5958 990 1 gnd
rlabel locali 5621 870 5650 876 1 vdd
rlabel locali 5834 867 5863 873 1 vdd
rlabel locali 5567 682 5589 697 1 d0
rlabel nwell 5988 837 6011 840 1 vdd
rlabel locali 5618 571 5647 577 1 gnd
rlabel locali 5831 571 5860 577 1 gnd
rlabel space 5928 566 5957 575 1 gnd
rlabel locali 6634 1104 6663 1110 1 vdd
rlabel locali 6847 1101 6876 1107 1 vdd
rlabel nwell 7001 1071 7024 1074 1 vdd
rlabel locali 6631 805 6660 811 1 gnd
rlabel locali 6844 805 6873 811 1 gnd
rlabel space 6941 800 6970 809 1 gnd
rlabel locali 6572 915 6619 936 1 d1
rlabel locali 6684 1524 6713 1530 1 vdd
rlabel locali 6897 1521 6926 1527 1 vdd
rlabel nwell 7051 1491 7074 1494 1 vdd
rlabel locali 6681 1225 6710 1231 1 gnd
rlabel locali 6894 1225 6923 1231 1 gnd
rlabel space 6991 1220 7020 1229 1 gnd
rlabel locali 6627 1336 6650 1351 1 d2
rlabel space 5916 2526 5945 2535 1 gnd
rlabel locali 6615 3296 6638 3311 1 d2
rlabel space 6979 3180 7008 3189 1 gnd
rlabel locali 6882 3185 6911 3191 1 gnd
rlabel locali 6669 3185 6698 3191 1 gnd
rlabel nwell 7039 3451 7062 3454 1 vdd
rlabel locali 6885 3481 6914 3487 1 vdd
rlabel locali 6672 3484 6701 3490 1 vdd
rlabel locali 6560 2875 6607 2896 1 d1
rlabel space 6929 2760 6958 2769 1 gnd
rlabel locali 6832 2765 6861 2771 1 gnd
rlabel locali 6619 2765 6648 2771 1 gnd
rlabel nwell 6989 3031 7012 3034 1 vdd
rlabel locali 6835 3061 6864 3067 1 vdd
rlabel locali 6622 3064 6651 3070 1 vdd
rlabel locali 5819 2531 5848 2537 1 gnd
rlabel locali 5606 2531 5635 2537 1 gnd
rlabel nwell 5976 2797 5999 2800 1 vdd
rlabel locali 5555 2642 5577 2657 1 d0
rlabel locali 5822 2827 5851 2833 1 vdd
rlabel locali 5609 2830 5638 2836 1 vdd
rlabel space 5917 2941 5946 2950 1 gnd
rlabel locali 5820 2946 5849 2952 1 gnd
rlabel locali 5607 2946 5636 2952 1 gnd
rlabel nwell 5977 3212 6000 3215 1 vdd
rlabel locali 5556 3057 5578 3072 1 d0
rlabel locali 5823 3242 5852 3248 1 vdd
rlabel locali 5610 3245 5639 3251 1 vdd
rlabel locali 6555 3856 6602 3877 1 d1
rlabel space 6924 3741 6953 3750 1 gnd
rlabel locali 6827 3746 6856 3752 1 gnd
rlabel locali 6614 3746 6643 3752 1 gnd
rlabel nwell 6984 4012 7007 4015 1 vdd
rlabel locali 6830 4042 6859 4048 1 vdd
rlabel locali 6617 4045 6646 4051 1 vdd
rlabel space 5911 3507 5940 3516 1 gnd
rlabel locali 5814 3512 5843 3518 1 gnd
rlabel locali 5601 3512 5630 3518 1 gnd
rlabel nwell 5971 3778 5994 3781 1 vdd
rlabel locali 5550 3623 5572 3638 1 d0
rlabel locali 5817 3808 5846 3814 1 vdd
rlabel locali 5604 3811 5633 3817 1 vdd
rlabel space 5912 3922 5941 3931 1 gnd
rlabel locali 5815 3927 5844 3933 1 gnd
rlabel locali 5602 3927 5631 3933 1 gnd
rlabel nwell 5972 4193 5995 4196 1 vdd
rlabel locali 5551 4038 5573 4053 1 d0
rlabel locali 5818 4223 5847 4229 1 vdd
rlabel locali 5605 4226 5634 4232 1 vdd
rlabel locali 6912 4477 6941 4483 1 vdd
rlabel locali 7125 4474 7154 4480 1 vdd
rlabel nwell 7279 4444 7302 4447 1 vdd
rlabel locali 6909 4178 6938 4184 1 gnd
rlabel locali 7122 4178 7151 4184 1 gnd
rlabel space 7219 4173 7248 4182 1 gnd
rlabel locali 6854 4283 6876 4307 1 d4
rlabel locali 10176 718 10205 724 5 vdd
rlabel locali 9963 721 9992 727 5 vdd
rlabel locali 10237 897 10259 912 5 d0
rlabel nwell 9815 754 9838 757 5 vdd
rlabel locali 10179 1017 10208 1023 5 gnd
rlabel locali 9966 1017 9995 1023 5 gnd
rlabel space 9869 1019 9898 1028 5 gnd
rlabel locali 10177 1133 10206 1139 5 vdd
rlabel locali 9964 1136 9993 1142 5 vdd
rlabel locali 10238 1312 10260 1327 5 d0
rlabel nwell 9816 1169 9839 1172 5 vdd
rlabel locali 10180 1432 10209 1438 5 gnd
rlabel locali 9967 1432 9996 1438 5 gnd
rlabel space 9870 1434 9899 1443 5 gnd
rlabel locali 9164 899 9193 905 5 vdd
rlabel locali 8951 902 8980 908 5 vdd
rlabel nwell 8803 935 8826 938 5 vdd
rlabel locali 9167 1198 9196 1204 5 gnd
rlabel locali 8954 1198 8983 1204 5 gnd
rlabel space 8857 1200 8886 1209 5 gnd
rlabel locali 9208 1073 9255 1094 5 d1
rlabel locali 10171 1699 10200 1705 5 vdd
rlabel locali 9958 1702 9987 1708 5 vdd
rlabel locali 10232 1878 10254 1893 5 d0
rlabel nwell 9810 1735 9833 1738 5 vdd
rlabel locali 10174 1998 10203 2004 5 gnd
rlabel locali 9961 1998 9990 2004 5 gnd
rlabel space 9864 2000 9893 2009 5 gnd
rlabel locali 10172 2114 10201 2120 5 vdd
rlabel locali 9959 2117 9988 2123 5 vdd
rlabel locali 10233 2293 10255 2308 5 d0
rlabel nwell 9811 2150 9834 2153 5 vdd
rlabel locali 10175 2413 10204 2419 5 gnd
rlabel locali 9962 2413 9991 2419 5 gnd
rlabel locali 9159 1880 9188 1886 5 vdd
rlabel locali 8946 1883 8975 1889 5 vdd
rlabel nwell 8798 1916 8821 1919 5 vdd
rlabel locali 9162 2179 9191 2185 5 gnd
rlabel locali 8949 2179 8978 2185 5 gnd
rlabel space 8852 2181 8881 2190 5 gnd
rlabel locali 9203 2054 9250 2075 5 d1
rlabel locali 9109 1460 9138 1466 5 vdd
rlabel locali 8896 1463 8925 1469 5 vdd
rlabel nwell 8748 1496 8771 1499 5 vdd
rlabel locali 9112 1759 9141 1765 5 gnd
rlabel locali 8899 1759 8928 1765 5 gnd
rlabel space 8802 1761 8831 1770 5 gnd
rlabel locali 9172 1639 9195 1654 5 d2
rlabel space 9865 2415 9894 2424 5 gnd
rlabel locali 9160 3599 9183 3614 5 d2
rlabel space 8790 3721 8819 3730 5 gnd
rlabel locali 8887 3719 8916 3725 5 gnd
rlabel locali 9100 3719 9129 3725 5 gnd
rlabel nwell 8736 3456 8759 3459 5 vdd
rlabel locali 8884 3423 8913 3429 5 vdd
rlabel locali 9097 3420 9126 3426 5 vdd
rlabel locali 9191 4014 9238 4035 5 d1
rlabel space 8840 4141 8869 4150 5 gnd
rlabel locali 8937 4139 8966 4145 5 gnd
rlabel locali 9150 4139 9179 4145 5 gnd
rlabel nwell 8786 3876 8809 3879 5 vdd
rlabel locali 8934 3843 8963 3849 5 vdd
rlabel locali 9147 3840 9176 3846 5 vdd
rlabel space 9853 4375 9882 4384 5 gnd
rlabel locali 9950 4373 9979 4379 5 gnd
rlabel locali 10163 4373 10192 4379 5 gnd
rlabel nwell 9799 4110 9822 4113 5 vdd
rlabel locali 10221 4253 10243 4268 5 d0
rlabel locali 9947 4077 9976 4083 5 vdd
rlabel locali 10160 4074 10189 4080 5 vdd
rlabel space 9852 3960 9881 3969 5 gnd
rlabel locali 9949 3958 9978 3964 5 gnd
rlabel locali 10162 3958 10191 3964 5 gnd
rlabel nwell 9798 3695 9821 3698 5 vdd
rlabel locali 10220 3838 10242 3853 5 d0
rlabel locali 9946 3662 9975 3668 5 vdd
rlabel locali 10159 3659 10188 3665 5 vdd
rlabel locali 9196 3033 9243 3054 5 d1
rlabel space 8845 3160 8874 3169 5 gnd
rlabel locali 8942 3158 8971 3164 5 gnd
rlabel locali 9155 3158 9184 3164 5 gnd
rlabel nwell 8791 2895 8814 2898 5 vdd
rlabel locali 8939 2862 8968 2868 5 vdd
rlabel locali 9152 2859 9181 2865 5 vdd
rlabel space 9858 3394 9887 3403 5 gnd
rlabel locali 9955 3392 9984 3398 5 gnd
rlabel locali 10168 3392 10197 3398 5 gnd
rlabel nwell 9804 3129 9827 3132 5 vdd
rlabel locali 10226 3272 10248 3287 5 d0
rlabel locali 9952 3096 9981 3102 5 vdd
rlabel locali 10165 3093 10194 3099 5 vdd
rlabel space 9857 2979 9886 2988 5 gnd
rlabel locali 9954 2977 9983 2983 5 gnd
rlabel locali 10167 2977 10196 2983 5 gnd
rlabel nwell 9803 2714 9826 2717 5 vdd
rlabel locali 10225 2857 10247 2872 5 d0
rlabel locali 9951 2681 9980 2687 5 vdd
rlabel locali 10164 2678 10193 2684 5 vdd
rlabel locali 8944 2392 8973 2398 5 vdd
rlabel locali 8731 2395 8760 2401 5 vdd
rlabel nwell 8583 2428 8606 2431 5 vdd
rlabel locali 8947 2691 8976 2697 5 gnd
rlabel locali 8734 2691 8763 2697 5 gnd
rlabel space 8637 2693 8666 2702 5 gnd
rlabel locali 9003 2569 9035 2588 5 d3
rlabel locali 8983 6486 9015 6505 5 d3
rlabel space 8617 6610 8646 6619 5 gnd
rlabel locali 8714 6608 8743 6614 5 gnd
rlabel locali 8927 6608 8956 6614 5 gnd
rlabel nwell 8563 6345 8586 6348 5 vdd
rlabel locali 8711 6312 8740 6318 5 vdd
rlabel locali 8924 6309 8953 6315 5 vdd
rlabel locali 10144 6595 10173 6601 5 vdd
rlabel locali 9931 6598 9960 6604 5 vdd
rlabel locali 10205 6774 10227 6789 5 d0
rlabel nwell 9783 6631 9806 6634 5 vdd
rlabel locali 10147 6894 10176 6900 5 gnd
rlabel locali 9934 6894 9963 6900 5 gnd
rlabel space 9837 6896 9866 6905 5 gnd
rlabel locali 10145 7010 10174 7016 5 vdd
rlabel locali 9932 7013 9961 7019 5 vdd
rlabel locali 10206 7189 10228 7204 5 d0
rlabel nwell 9784 7046 9807 7049 5 vdd
rlabel locali 10148 7309 10177 7315 5 gnd
rlabel locali 9935 7309 9964 7315 5 gnd
rlabel space 9838 7311 9867 7320 5 gnd
rlabel locali 9132 6776 9161 6782 5 vdd
rlabel locali 8919 6779 8948 6785 5 vdd
rlabel nwell 8771 6812 8794 6815 5 vdd
rlabel locali 9135 7075 9164 7081 5 gnd
rlabel locali 8922 7075 8951 7081 5 gnd
rlabel space 8825 7077 8854 7086 5 gnd
rlabel locali 9176 6950 9223 6971 5 d1
rlabel locali 10139 7576 10168 7582 5 vdd
rlabel locali 9926 7579 9955 7585 5 vdd
rlabel locali 10200 7755 10222 7770 5 d0
rlabel nwell 9778 7612 9801 7615 5 vdd
rlabel locali 10142 7875 10171 7881 5 gnd
rlabel locali 9929 7875 9958 7881 5 gnd
rlabel space 9832 7877 9861 7886 5 gnd
rlabel locali 10140 7991 10169 7997 5 vdd
rlabel locali 9927 7994 9956 8000 5 vdd
rlabel locali 10201 8170 10223 8185 5 d0
rlabel nwell 9779 8027 9802 8030 5 vdd
rlabel locali 10143 8290 10172 8296 5 gnd
rlabel locali 9930 8290 9959 8296 5 gnd
rlabel space 9833 8292 9862 8301 5 gnd
rlabel locali 9127 7757 9156 7763 5 vdd
rlabel locali 8914 7760 8943 7766 5 vdd
rlabel nwell 8766 7793 8789 7796 5 vdd
rlabel locali 9130 8056 9159 8062 5 gnd
rlabel locali 8917 8056 8946 8062 5 gnd
rlabel space 8820 8058 8849 8067 5 gnd
rlabel locali 9171 7931 9218 7952 5 d1
rlabel locali 9077 7337 9106 7343 5 vdd
rlabel locali 8864 7340 8893 7346 5 vdd
rlabel nwell 8716 7373 8739 7376 5 vdd
rlabel locali 9080 7636 9109 7642 5 gnd
rlabel locali 8867 7636 8896 7642 5 gnd
rlabel space 8770 7638 8799 7647 5 gnd
rlabel locali 9140 7516 9163 7531 5 d2
rlabel space 9845 6332 9874 6341 5 gnd
rlabel locali 9152 5556 9175 5571 5 d2
rlabel space 8782 5678 8811 5687 5 gnd
rlabel locali 8879 5676 8908 5682 5 gnd
rlabel locali 9092 5676 9121 5682 5 gnd
rlabel nwell 8728 5413 8751 5416 5 vdd
rlabel locali 8876 5380 8905 5386 5 vdd
rlabel locali 9089 5377 9118 5383 5 vdd
rlabel locali 9183 5971 9230 5992 5 d1
rlabel space 8832 6098 8861 6107 5 gnd
rlabel locali 8929 6096 8958 6102 5 gnd
rlabel locali 9142 6096 9171 6102 5 gnd
rlabel nwell 8778 5833 8801 5836 5 vdd
rlabel locali 8926 5800 8955 5806 5 vdd
rlabel locali 9139 5797 9168 5803 5 vdd
rlabel locali 9942 6330 9971 6336 5 gnd
rlabel locali 10155 6330 10184 6336 5 gnd
rlabel nwell 9791 6067 9814 6070 5 vdd
rlabel locali 10213 6210 10235 6225 5 d0
rlabel locali 9939 6034 9968 6040 5 vdd
rlabel locali 10152 6031 10181 6037 5 vdd
rlabel space 9844 5917 9873 5926 5 gnd
rlabel locali 9941 5915 9970 5921 5 gnd
rlabel locali 10154 5915 10183 5921 5 gnd
rlabel nwell 9790 5652 9813 5655 5 vdd
rlabel locali 10212 5795 10234 5810 5 d0
rlabel locali 9938 5619 9967 5625 5 vdd
rlabel locali 10151 5616 10180 5622 5 vdd
rlabel locali 9188 4990 9235 5011 5 d1
rlabel space 8837 5117 8866 5126 5 gnd
rlabel locali 8934 5115 8963 5121 5 gnd
rlabel locali 9147 5115 9176 5121 5 gnd
rlabel nwell 8783 4852 8806 4855 5 vdd
rlabel locali 8931 4819 8960 4825 5 vdd
rlabel locali 9144 4816 9173 4822 5 vdd
rlabel space 9850 5351 9879 5360 5 gnd
rlabel locali 9947 5349 9976 5355 5 gnd
rlabel locali 10160 5349 10189 5355 5 gnd
rlabel nwell 9796 5086 9819 5089 5 vdd
rlabel locali 10218 5229 10240 5244 5 d0
rlabel locali 9944 5053 9973 5059 5 vdd
rlabel locali 10157 5050 10186 5056 5 vdd
rlabel space 9849 4936 9878 4945 5 gnd
rlabel locali 9946 4934 9975 4940 5 gnd
rlabel locali 10159 4934 10188 4940 5 gnd
rlabel nwell 9795 4671 9818 4674 5 vdd
rlabel locali 10217 4814 10239 4829 5 d0
rlabel locali 9943 4638 9972 4644 5 vdd
rlabel locali 10156 4635 10185 4641 5 vdd
rlabel locali 8849 4384 8878 4390 5 vdd
rlabel locali 8636 4387 8665 4393 5 vdd
rlabel nwell 8488 4420 8511 4423 5 vdd
rlabel locali 8852 4683 8881 4689 5 gnd
rlabel locali 8639 4683 8668 4689 5 gnd
rlabel space 8542 4685 8571 4694 5 gnd
rlabel locali 8914 4560 8936 4584 5 d4
rlabel locali 7024 389 7053 395 1 vdd
rlabel locali 7237 386 7266 392 1 vdd
rlabel nwell 7391 356 7414 359 1 vdd
rlabel locali 7021 90 7050 96 1 gnd
rlabel locali 7234 90 7263 96 1 gnd
rlabel space 7331 85 7360 94 1 gnd
rlabel locali 6966 198 6990 215 1 d5
rlabel locali 4833 322 4862 328 1 vdd
rlabel locali 5046 319 5075 325 1 vdd
rlabel nwell 5200 289 5223 292 1 vdd
rlabel locali 4830 23 4859 29 1 gnd
rlabel locali 5043 23 5072 29 1 gnd
rlabel space 5140 18 5169 27 1 gnd
rlabel locali 4777 129 4796 149 1 d6
rlabel locali 10965 8172 10994 8178 1 vdd
rlabel locali 11178 8169 11207 8175 1 vdd
rlabel locali 10911 7984 10933 7999 1 d0
rlabel nwell 11332 8139 11355 8142 1 vdd
rlabel locali 10962 7873 10991 7879 1 gnd
rlabel locali 11175 7873 11204 7879 1 gnd
rlabel space 11272 7868 11301 7877 1 gnd
rlabel locali 10964 7757 10993 7763 1 vdd
rlabel locali 11177 7754 11206 7760 1 vdd
rlabel locali 10910 7569 10932 7584 1 d0
rlabel nwell 11331 7724 11354 7727 1 vdd
rlabel locali 10961 7458 10990 7464 1 gnd
rlabel locali 11174 7458 11203 7464 1 gnd
rlabel space 11271 7453 11300 7462 1 gnd
rlabel locali 11977 7991 12006 7997 1 vdd
rlabel locali 12190 7988 12219 7994 1 vdd
rlabel nwell 12344 7958 12367 7961 1 vdd
rlabel locali 11974 7692 12003 7698 1 gnd
rlabel locali 12187 7692 12216 7698 1 gnd
rlabel space 12284 7687 12313 7696 1 gnd
rlabel locali 11915 7802 11962 7823 1 d1
rlabel locali 10970 7191 10999 7197 1 vdd
rlabel locali 11183 7188 11212 7194 1 vdd
rlabel locali 10916 7003 10938 7018 1 d0
rlabel nwell 11337 7158 11360 7161 1 vdd
rlabel locali 10967 6892 10996 6898 1 gnd
rlabel locali 11180 6892 11209 6898 1 gnd
rlabel space 11277 6887 11306 6896 1 gnd
rlabel locali 10969 6776 10998 6782 1 vdd
rlabel locali 11182 6773 11211 6779 1 vdd
rlabel locali 10915 6588 10937 6603 1 d0
rlabel nwell 11336 6743 11359 6746 1 vdd
rlabel locali 10966 6477 10995 6483 1 gnd
rlabel locali 11179 6477 11208 6483 1 gnd
rlabel locali 11982 7010 12011 7016 1 vdd
rlabel locali 12195 7007 12224 7013 1 vdd
rlabel nwell 12349 6977 12372 6980 1 vdd
rlabel locali 11979 6711 12008 6717 1 gnd
rlabel locali 12192 6711 12221 6717 1 gnd
rlabel space 12289 6706 12318 6715 1 gnd
rlabel locali 11920 6821 11967 6842 1 d1
rlabel locali 12032 7430 12061 7436 1 vdd
rlabel locali 12245 7427 12274 7433 1 vdd
rlabel nwell 12399 7397 12422 7400 1 vdd
rlabel locali 12029 7131 12058 7137 1 gnd
rlabel locali 12242 7131 12271 7137 1 gnd
rlabel space 12339 7126 12368 7135 1 gnd
rlabel locali 11975 7242 11998 7257 1 d2
rlabel space 11276 6472 11305 6481 1 gnd
rlabel locali 11987 5282 12010 5297 1 d2
rlabel space 12351 5166 12380 5175 1 gnd
rlabel locali 12254 5171 12283 5177 1 gnd
rlabel locali 12041 5171 12070 5177 1 gnd
rlabel nwell 12411 5437 12434 5440 1 vdd
rlabel locali 12257 5467 12286 5473 1 vdd
rlabel locali 12044 5470 12073 5476 1 vdd
rlabel locali 11932 4861 11979 4882 1 d1
rlabel space 12301 4746 12330 4755 1 gnd
rlabel locali 12204 4751 12233 4757 1 gnd
rlabel locali 11991 4751 12020 4757 1 gnd
rlabel nwell 12361 5017 12384 5020 1 vdd
rlabel locali 12207 5047 12236 5053 1 vdd
rlabel locali 11994 5050 12023 5056 1 vdd
rlabel space 11288 4512 11317 4521 1 gnd
rlabel locali 11191 4517 11220 4523 1 gnd
rlabel locali 10978 4517 11007 4523 1 gnd
rlabel nwell 11348 4783 11371 4786 1 vdd
rlabel locali 10927 4628 10949 4643 1 d0
rlabel locali 11194 4813 11223 4819 1 vdd
rlabel locali 10981 4816 11010 4822 1 vdd
rlabel space 11289 4927 11318 4936 1 gnd
rlabel locali 11192 4932 11221 4938 1 gnd
rlabel locali 10979 4932 11008 4938 1 gnd
rlabel nwell 11349 5198 11372 5201 1 vdd
rlabel locali 10928 5043 10950 5058 1 d0
rlabel locali 11195 5228 11224 5234 1 vdd
rlabel locali 10982 5231 11011 5237 1 vdd
rlabel locali 11927 5842 11974 5863 1 d1
rlabel space 12296 5727 12325 5736 1 gnd
rlabel locali 12199 5732 12228 5738 1 gnd
rlabel locali 11986 5732 12015 5738 1 gnd
rlabel nwell 12356 5998 12379 6001 1 vdd
rlabel locali 12202 6028 12231 6034 1 vdd
rlabel locali 11989 6031 12018 6037 1 vdd
rlabel space 11283 5493 11312 5502 1 gnd
rlabel locali 11186 5498 11215 5504 1 gnd
rlabel locali 10973 5498 11002 5504 1 gnd
rlabel nwell 11343 5764 11366 5767 1 vdd
rlabel locali 10922 5609 10944 5624 1 d0
rlabel locali 11189 5794 11218 5800 1 vdd
rlabel locali 10976 5797 11005 5803 1 vdd
rlabel space 11284 5908 11313 5917 1 gnd
rlabel locali 11187 5913 11216 5919 1 gnd
rlabel locali 10974 5913 11003 5919 1 gnd
rlabel nwell 11344 6179 11367 6182 1 vdd
rlabel locali 10923 6024 10945 6039 1 d0
rlabel locali 11190 6209 11219 6215 1 vdd
rlabel locali 10977 6212 11006 6218 1 vdd
rlabel locali 12197 6498 12226 6504 1 vdd
rlabel locali 12410 6495 12439 6501 1 vdd
rlabel nwell 12564 6465 12587 6468 1 vdd
rlabel locali 12194 6199 12223 6205 1 gnd
rlabel locali 12407 6199 12436 6205 1 gnd
rlabel space 12504 6194 12533 6203 1 gnd
rlabel locali 12135 6308 12167 6327 1 d3
rlabel locali 12155 2391 12187 2410 1 d3
rlabel space 12524 2277 12553 2286 1 gnd
rlabel locali 12427 2282 12456 2288 1 gnd
rlabel locali 12214 2282 12243 2288 1 gnd
rlabel nwell 12584 2548 12607 2551 1 vdd
rlabel locali 12430 2578 12459 2584 1 vdd
rlabel locali 12217 2581 12246 2587 1 vdd
rlabel locali 10997 2295 11026 2301 1 vdd
rlabel locali 11210 2292 11239 2298 1 vdd
rlabel locali 10943 2107 10965 2122 1 d0
rlabel nwell 11364 2262 11387 2265 1 vdd
rlabel locali 10994 1996 11023 2002 1 gnd
rlabel locali 11207 1996 11236 2002 1 gnd
rlabel space 11304 1991 11333 2000 1 gnd
rlabel locali 10996 1880 11025 1886 1 vdd
rlabel locali 11209 1877 11238 1883 1 vdd
rlabel locali 10942 1692 10964 1707 1 d0
rlabel nwell 11363 1847 11386 1850 1 vdd
rlabel locali 10993 1581 11022 1587 1 gnd
rlabel locali 11206 1581 11235 1587 1 gnd
rlabel space 11303 1576 11332 1585 1 gnd
rlabel locali 12009 2114 12038 2120 1 vdd
rlabel locali 12222 2111 12251 2117 1 vdd
rlabel nwell 12376 2081 12399 2084 1 vdd
rlabel locali 12006 1815 12035 1821 1 gnd
rlabel locali 12219 1815 12248 1821 1 gnd
rlabel space 12316 1810 12345 1819 1 gnd
rlabel locali 11947 1925 11994 1946 1 d1
rlabel locali 11002 1314 11031 1320 1 vdd
rlabel locali 11215 1311 11244 1317 1 vdd
rlabel locali 10948 1126 10970 1141 1 d0
rlabel nwell 11369 1281 11392 1284 1 vdd
rlabel locali 10999 1015 11028 1021 1 gnd
rlabel locali 11212 1015 11241 1021 1 gnd
rlabel space 11309 1010 11338 1019 1 gnd
rlabel locali 11001 899 11030 905 1 vdd
rlabel locali 11214 896 11243 902 1 vdd
rlabel locali 10947 711 10969 726 1 d0
rlabel nwell 11368 866 11391 869 1 vdd
rlabel locali 10998 600 11027 606 1 gnd
rlabel locali 11211 600 11240 606 1 gnd
rlabel space 11308 595 11337 604 1 gnd
rlabel locali 12014 1133 12043 1139 1 vdd
rlabel locali 12227 1130 12256 1136 1 vdd
rlabel nwell 12381 1100 12404 1103 1 vdd
rlabel locali 12011 834 12040 840 1 gnd
rlabel locali 12224 834 12253 840 1 gnd
rlabel space 12321 829 12350 838 1 gnd
rlabel locali 11952 944 11999 965 1 d1
rlabel locali 12064 1553 12093 1559 1 vdd
rlabel locali 12277 1550 12306 1556 1 vdd
rlabel nwell 12431 1520 12454 1523 1 vdd
rlabel locali 12061 1254 12090 1260 1 gnd
rlabel locali 12274 1254 12303 1260 1 gnd
rlabel space 12371 1249 12400 1258 1 gnd
rlabel locali 12007 1365 12030 1380 1 d2
rlabel space 11296 2555 11325 2564 1 gnd
rlabel locali 11995 3325 12018 3340 1 d2
rlabel space 12359 3209 12388 3218 1 gnd
rlabel locali 12262 3214 12291 3220 1 gnd
rlabel locali 12049 3214 12078 3220 1 gnd
rlabel nwell 12419 3480 12442 3483 1 vdd
rlabel locali 12265 3510 12294 3516 1 vdd
rlabel locali 12052 3513 12081 3519 1 vdd
rlabel locali 11940 2904 11987 2925 1 d1
rlabel space 12309 2789 12338 2798 1 gnd
rlabel locali 12212 2794 12241 2800 1 gnd
rlabel locali 11999 2794 12028 2800 1 gnd
rlabel nwell 12369 3060 12392 3063 1 vdd
rlabel locali 12215 3090 12244 3096 1 vdd
rlabel locali 12002 3093 12031 3099 1 vdd
rlabel locali 11199 2560 11228 2566 1 gnd
rlabel locali 10986 2560 11015 2566 1 gnd
rlabel nwell 11356 2826 11379 2829 1 vdd
rlabel locali 10935 2671 10957 2686 1 d0
rlabel locali 11202 2856 11231 2862 1 vdd
rlabel locali 10989 2859 11018 2865 1 vdd
rlabel space 11297 2970 11326 2979 1 gnd
rlabel locali 11200 2975 11229 2981 1 gnd
rlabel locali 10987 2975 11016 2981 1 gnd
rlabel nwell 11357 3241 11380 3244 1 vdd
rlabel locali 10936 3086 10958 3101 1 d0
rlabel locali 11203 3271 11232 3277 1 vdd
rlabel locali 10990 3274 11019 3280 1 vdd
rlabel locali 11935 3885 11982 3906 1 d1
rlabel space 12304 3770 12333 3779 1 gnd
rlabel locali 12207 3775 12236 3781 1 gnd
rlabel locali 11994 3775 12023 3781 1 gnd
rlabel nwell 12364 4041 12387 4044 1 vdd
rlabel locali 12210 4071 12239 4077 1 vdd
rlabel locali 11997 4074 12026 4080 1 vdd
rlabel space 11291 3536 11320 3545 1 gnd
rlabel locali 11194 3541 11223 3547 1 gnd
rlabel locali 10981 3541 11010 3547 1 gnd
rlabel nwell 11351 3807 11374 3810 1 vdd
rlabel locali 10930 3652 10952 3667 1 d0
rlabel locali 11197 3837 11226 3843 1 vdd
rlabel locali 10984 3840 11013 3846 1 vdd
rlabel space 11292 3951 11321 3960 1 gnd
rlabel locali 11195 3956 11224 3962 1 gnd
rlabel locali 10982 3956 11011 3962 1 gnd
rlabel nwell 11352 4222 11375 4225 1 vdd
rlabel locali 10931 4067 10953 4082 1 d0
rlabel locali 11198 4252 11227 4258 1 vdd
rlabel locali 10985 4255 11014 4261 1 vdd
rlabel locali 12292 4506 12321 4512 1 vdd
rlabel locali 12505 4503 12534 4509 1 vdd
rlabel nwell 12659 4473 12682 4476 1 vdd
rlabel locali 12289 4207 12318 4213 1 gnd
rlabel locali 12502 4207 12531 4213 1 gnd
rlabel space 12599 4202 12628 4211 1 gnd
rlabel locali 12234 4312 12256 4336 1 d4
rlabel locali 15556 747 15585 753 5 vdd
rlabel locali 15343 750 15372 756 5 vdd
rlabel locali 15617 926 15639 941 5 d0
rlabel nwell 15195 783 15218 786 5 vdd
rlabel locali 15559 1046 15588 1052 5 gnd
rlabel locali 15346 1046 15375 1052 5 gnd
rlabel space 15249 1048 15278 1057 5 gnd
rlabel locali 15557 1162 15586 1168 5 vdd
rlabel locali 15344 1165 15373 1171 5 vdd
rlabel locali 15618 1341 15640 1356 5 d0
rlabel nwell 15196 1198 15219 1201 5 vdd
rlabel locali 15560 1461 15589 1467 5 gnd
rlabel locali 15347 1461 15376 1467 5 gnd
rlabel space 15250 1463 15279 1472 5 gnd
rlabel locali 14544 928 14573 934 5 vdd
rlabel locali 14331 931 14360 937 5 vdd
rlabel nwell 14183 964 14206 967 5 vdd
rlabel locali 14547 1227 14576 1233 5 gnd
rlabel locali 14334 1227 14363 1233 5 gnd
rlabel space 14237 1229 14266 1238 5 gnd
rlabel locali 14588 1102 14635 1123 5 d1
rlabel locali 15551 1728 15580 1734 5 vdd
rlabel locali 15338 1731 15367 1737 5 vdd
rlabel locali 15612 1907 15634 1922 5 d0
rlabel nwell 15190 1764 15213 1767 5 vdd
rlabel locali 15554 2027 15583 2033 5 gnd
rlabel locali 15341 2027 15370 2033 5 gnd
rlabel space 15244 2029 15273 2038 5 gnd
rlabel locali 15552 2143 15581 2149 5 vdd
rlabel locali 15339 2146 15368 2152 5 vdd
rlabel locali 15613 2322 15635 2337 5 d0
rlabel nwell 15191 2179 15214 2182 5 vdd
rlabel locali 15555 2442 15584 2448 5 gnd
rlabel locali 15342 2442 15371 2448 5 gnd
rlabel locali 14539 1909 14568 1915 5 vdd
rlabel locali 14326 1912 14355 1918 5 vdd
rlabel nwell 14178 1945 14201 1948 5 vdd
rlabel locali 14542 2208 14571 2214 5 gnd
rlabel locali 14329 2208 14358 2214 5 gnd
rlabel space 14232 2210 14261 2219 5 gnd
rlabel locali 14583 2083 14630 2104 5 d1
rlabel locali 14489 1489 14518 1495 5 vdd
rlabel locali 14276 1492 14305 1498 5 vdd
rlabel nwell 14128 1525 14151 1528 5 vdd
rlabel locali 14492 1788 14521 1794 5 gnd
rlabel locali 14279 1788 14308 1794 5 gnd
rlabel space 14182 1790 14211 1799 5 gnd
rlabel locali 14552 1668 14575 1683 5 d2
rlabel space 15245 2444 15274 2453 5 gnd
rlabel locali 14540 3628 14563 3643 5 d2
rlabel space 14170 3750 14199 3759 5 gnd
rlabel locali 14267 3748 14296 3754 5 gnd
rlabel locali 14480 3748 14509 3754 5 gnd
rlabel nwell 14116 3485 14139 3488 5 vdd
rlabel locali 14264 3452 14293 3458 5 vdd
rlabel locali 14477 3449 14506 3455 5 vdd
rlabel locali 14571 4043 14618 4064 5 d1
rlabel space 14220 4170 14249 4179 5 gnd
rlabel locali 14317 4168 14346 4174 5 gnd
rlabel locali 14530 4168 14559 4174 5 gnd
rlabel nwell 14166 3905 14189 3908 5 vdd
rlabel locali 14314 3872 14343 3878 5 vdd
rlabel locali 14527 3869 14556 3875 5 vdd
rlabel space 15233 4404 15262 4413 5 gnd
rlabel locali 15330 4402 15359 4408 5 gnd
rlabel locali 15543 4402 15572 4408 5 gnd
rlabel nwell 15179 4139 15202 4142 5 vdd
rlabel locali 15601 4282 15623 4297 5 d0
rlabel locali 15327 4106 15356 4112 5 vdd
rlabel locali 15540 4103 15569 4109 5 vdd
rlabel space 15232 3989 15261 3998 5 gnd
rlabel locali 15329 3987 15358 3993 5 gnd
rlabel locali 15542 3987 15571 3993 5 gnd
rlabel nwell 15178 3724 15201 3727 5 vdd
rlabel locali 15600 3867 15622 3882 5 d0
rlabel locali 15326 3691 15355 3697 5 vdd
rlabel locali 15539 3688 15568 3694 5 vdd
rlabel locali 14576 3062 14623 3083 5 d1
rlabel space 14225 3189 14254 3198 5 gnd
rlabel locali 14322 3187 14351 3193 5 gnd
rlabel locali 14535 3187 14564 3193 5 gnd
rlabel nwell 14171 2924 14194 2927 5 vdd
rlabel locali 14319 2891 14348 2897 5 vdd
rlabel locali 14532 2888 14561 2894 5 vdd
rlabel space 15238 3423 15267 3432 5 gnd
rlabel locali 15335 3421 15364 3427 5 gnd
rlabel locali 15548 3421 15577 3427 5 gnd
rlabel nwell 15184 3158 15207 3161 5 vdd
rlabel locali 15606 3301 15628 3316 5 d0
rlabel locali 15332 3125 15361 3131 5 vdd
rlabel locali 15545 3122 15574 3128 5 vdd
rlabel space 15237 3008 15266 3017 5 gnd
rlabel locali 15334 3006 15363 3012 5 gnd
rlabel locali 15547 3006 15576 3012 5 gnd
rlabel nwell 15183 2743 15206 2746 5 vdd
rlabel locali 15605 2886 15627 2901 5 d0
rlabel locali 15331 2710 15360 2716 5 vdd
rlabel locali 15544 2707 15573 2713 5 vdd
rlabel locali 14324 2421 14353 2427 5 vdd
rlabel locali 14111 2424 14140 2430 5 vdd
rlabel nwell 13963 2457 13986 2460 5 vdd
rlabel locali 14327 2720 14356 2726 5 gnd
rlabel locali 14114 2720 14143 2726 5 gnd
rlabel space 14017 2722 14046 2731 5 gnd
rlabel locali 14383 2598 14415 2617 5 d3
rlabel locali 14363 6515 14395 6534 5 d3
rlabel space 13997 6639 14026 6648 5 gnd
rlabel locali 14094 6637 14123 6643 5 gnd
rlabel locali 14307 6637 14336 6643 5 gnd
rlabel nwell 13943 6374 13966 6377 5 vdd
rlabel locali 14091 6341 14120 6347 5 vdd
rlabel locali 14304 6338 14333 6344 5 vdd
rlabel locali 15524 6624 15553 6630 5 vdd
rlabel locali 15311 6627 15340 6633 5 vdd
rlabel locali 15585 6803 15607 6818 5 d0
rlabel nwell 15163 6660 15186 6663 5 vdd
rlabel locali 15527 6923 15556 6929 5 gnd
rlabel locali 15314 6923 15343 6929 5 gnd
rlabel space 15217 6925 15246 6934 5 gnd
rlabel locali 15525 7039 15554 7045 5 vdd
rlabel locali 15312 7042 15341 7048 5 vdd
rlabel locali 15586 7218 15608 7233 5 d0
rlabel nwell 15164 7075 15187 7078 5 vdd
rlabel locali 15528 7338 15557 7344 5 gnd
rlabel locali 15315 7338 15344 7344 5 gnd
rlabel space 15218 7340 15247 7349 5 gnd
rlabel locali 14512 6805 14541 6811 5 vdd
rlabel locali 14299 6808 14328 6814 5 vdd
rlabel nwell 14151 6841 14174 6844 5 vdd
rlabel locali 14515 7104 14544 7110 5 gnd
rlabel locali 14302 7104 14331 7110 5 gnd
rlabel space 14205 7106 14234 7115 5 gnd
rlabel locali 14556 6979 14603 7000 5 d1
rlabel locali 15519 7605 15548 7611 5 vdd
rlabel locali 15306 7608 15335 7614 5 vdd
rlabel locali 15580 7784 15602 7799 5 d0
rlabel nwell 15158 7641 15181 7644 5 vdd
rlabel locali 15522 7904 15551 7910 5 gnd
rlabel locali 15309 7904 15338 7910 5 gnd
rlabel space 15212 7906 15241 7915 5 gnd
rlabel locali 15520 8020 15549 8026 5 vdd
rlabel locali 15307 8023 15336 8029 5 vdd
rlabel locali 15581 8199 15603 8214 5 d0
rlabel nwell 15159 8056 15182 8059 5 vdd
rlabel locali 15523 8319 15552 8325 5 gnd
rlabel locali 15310 8319 15339 8325 5 gnd
rlabel space 15213 8321 15242 8330 5 gnd
rlabel locali 14507 7786 14536 7792 5 vdd
rlabel locali 14294 7789 14323 7795 5 vdd
rlabel nwell 14146 7822 14169 7825 5 vdd
rlabel locali 14510 8085 14539 8091 5 gnd
rlabel locali 14297 8085 14326 8091 5 gnd
rlabel space 14200 8087 14229 8096 5 gnd
rlabel locali 14551 7960 14598 7981 5 d1
rlabel locali 14457 7366 14486 7372 5 vdd
rlabel locali 14244 7369 14273 7375 5 vdd
rlabel nwell 14096 7402 14119 7405 5 vdd
rlabel locali 14460 7665 14489 7671 5 gnd
rlabel locali 14247 7665 14276 7671 5 gnd
rlabel space 14150 7667 14179 7676 5 gnd
rlabel locali 14520 7545 14543 7560 5 d2
rlabel space 15225 6361 15254 6370 5 gnd
rlabel locali 14532 5585 14555 5600 5 d2
rlabel space 14162 5707 14191 5716 5 gnd
rlabel locali 14259 5705 14288 5711 5 gnd
rlabel locali 14472 5705 14501 5711 5 gnd
rlabel nwell 14108 5442 14131 5445 5 vdd
rlabel locali 14256 5409 14285 5415 5 vdd
rlabel locali 14469 5406 14498 5412 5 vdd
rlabel locali 14563 6000 14610 6021 5 d1
rlabel space 14212 6127 14241 6136 5 gnd
rlabel locali 14309 6125 14338 6131 5 gnd
rlabel locali 14522 6125 14551 6131 5 gnd
rlabel nwell 14158 5862 14181 5865 5 vdd
rlabel locali 14306 5829 14335 5835 5 vdd
rlabel locali 14519 5826 14548 5832 5 vdd
rlabel locali 15322 6359 15351 6365 5 gnd
rlabel locali 15535 6359 15564 6365 5 gnd
rlabel nwell 15171 6096 15194 6099 5 vdd
rlabel locali 15593 6239 15615 6254 5 d0
rlabel locali 15319 6063 15348 6069 5 vdd
rlabel locali 15532 6060 15561 6066 5 vdd
rlabel space 15224 5946 15253 5955 5 gnd
rlabel locali 15321 5944 15350 5950 5 gnd
rlabel locali 15534 5944 15563 5950 5 gnd
rlabel nwell 15170 5681 15193 5684 5 vdd
rlabel locali 15592 5824 15614 5839 5 d0
rlabel locali 15318 5648 15347 5654 5 vdd
rlabel locali 15531 5645 15560 5651 5 vdd
rlabel locali 14568 5019 14615 5040 5 d1
rlabel space 14217 5146 14246 5155 5 gnd
rlabel locali 14314 5144 14343 5150 5 gnd
rlabel locali 14527 5144 14556 5150 5 gnd
rlabel nwell 14163 4881 14186 4884 5 vdd
rlabel locali 14311 4848 14340 4854 5 vdd
rlabel locali 14524 4845 14553 4851 5 vdd
rlabel space 15230 5380 15259 5389 5 gnd
rlabel locali 15327 5378 15356 5384 5 gnd
rlabel locali 15540 5378 15569 5384 5 gnd
rlabel nwell 15176 5115 15199 5118 5 vdd
rlabel locali 15598 5258 15620 5273 5 d0
rlabel locali 15324 5082 15353 5088 5 vdd
rlabel locali 15537 5079 15566 5085 5 vdd
rlabel space 15229 4965 15258 4974 5 gnd
rlabel locali 15326 4963 15355 4969 5 gnd
rlabel locali 15539 4963 15568 4969 5 gnd
rlabel nwell 15175 4700 15198 4703 5 vdd
rlabel locali 15597 4843 15619 4858 5 d0
rlabel locali 15323 4667 15352 4673 5 vdd
rlabel locali 15536 4664 15565 4670 5 vdd
rlabel locali 14229 4413 14258 4419 5 vdd
rlabel locali 14016 4416 14045 4422 5 vdd
rlabel nwell 13868 4449 13891 4452 5 vdd
rlabel locali 14232 4712 14261 4718 5 gnd
rlabel locali 14019 4712 14048 4718 5 gnd
rlabel space 13922 4714 13951 4723 5 gnd
rlabel locali 14294 4589 14316 4613 5 d4
rlabel locali 12404 418 12433 424 1 vdd
rlabel locali 12617 415 12646 421 1 vdd
rlabel nwell 12771 385 12794 388 1 vdd
rlabel locali 12401 119 12430 125 1 gnd
rlabel locali 12614 119 12643 125 1 gnd
rlabel space 12711 114 12740 123 1 gnd
rlabel locali 12346 227 12370 244 1 d5
rlabel locali 16246 8151 16275 8157 1 vdd
rlabel locali 16459 8148 16488 8154 1 vdd
rlabel locali 16192 7963 16214 7978 1 d0
rlabel nwell 16613 8118 16636 8121 1 vdd
rlabel locali 16243 7852 16272 7858 1 gnd
rlabel locali 16456 7852 16485 7858 1 gnd
rlabel space 16553 7847 16582 7856 1 gnd
rlabel locali 16245 7736 16274 7742 1 vdd
rlabel locali 16458 7733 16487 7739 1 vdd
rlabel locali 16191 7548 16213 7563 1 d0
rlabel nwell 16612 7703 16635 7706 1 vdd
rlabel locali 16242 7437 16271 7443 1 gnd
rlabel locali 16455 7437 16484 7443 1 gnd
rlabel space 16552 7432 16581 7441 1 gnd
rlabel locali 17258 7970 17287 7976 1 vdd
rlabel locali 17471 7967 17500 7973 1 vdd
rlabel nwell 17625 7937 17648 7940 1 vdd
rlabel locali 17255 7671 17284 7677 1 gnd
rlabel locali 17468 7671 17497 7677 1 gnd
rlabel space 17565 7666 17594 7675 1 gnd
rlabel locali 17196 7781 17243 7802 1 d1
rlabel locali 16251 7170 16280 7176 1 vdd
rlabel locali 16464 7167 16493 7173 1 vdd
rlabel locali 16197 6982 16219 6997 1 d0
rlabel nwell 16618 7137 16641 7140 1 vdd
rlabel locali 16248 6871 16277 6877 1 gnd
rlabel locali 16461 6871 16490 6877 1 gnd
rlabel space 16558 6866 16587 6875 1 gnd
rlabel locali 16250 6755 16279 6761 1 vdd
rlabel locali 16463 6752 16492 6758 1 vdd
rlabel locali 16196 6567 16218 6582 1 d0
rlabel nwell 16617 6722 16640 6725 1 vdd
rlabel locali 16247 6456 16276 6462 1 gnd
rlabel locali 16460 6456 16489 6462 1 gnd
rlabel locali 17263 6989 17292 6995 1 vdd
rlabel locali 17476 6986 17505 6992 1 vdd
rlabel nwell 17630 6956 17653 6959 1 vdd
rlabel locali 17260 6690 17289 6696 1 gnd
rlabel locali 17473 6690 17502 6696 1 gnd
rlabel space 17570 6685 17599 6694 1 gnd
rlabel locali 17201 6800 17248 6821 1 d1
rlabel locali 17313 7409 17342 7415 1 vdd
rlabel locali 17526 7406 17555 7412 1 vdd
rlabel nwell 17680 7376 17703 7379 1 vdd
rlabel locali 17310 7110 17339 7116 1 gnd
rlabel locali 17523 7110 17552 7116 1 gnd
rlabel space 17620 7105 17649 7114 1 gnd
rlabel locali 17256 7221 17279 7236 1 d2
rlabel space 16557 6451 16586 6460 1 gnd
rlabel locali 17268 5261 17291 5276 1 d2
rlabel space 17632 5145 17661 5154 1 gnd
rlabel locali 17535 5150 17564 5156 1 gnd
rlabel locali 17322 5150 17351 5156 1 gnd
rlabel nwell 17692 5416 17715 5419 1 vdd
rlabel locali 17538 5446 17567 5452 1 vdd
rlabel locali 17325 5449 17354 5455 1 vdd
rlabel locali 17213 4840 17260 4861 1 d1
rlabel space 17582 4725 17611 4734 1 gnd
rlabel locali 17485 4730 17514 4736 1 gnd
rlabel locali 17272 4730 17301 4736 1 gnd
rlabel nwell 17642 4996 17665 4999 1 vdd
rlabel locali 17488 5026 17517 5032 1 vdd
rlabel locali 17275 5029 17304 5035 1 vdd
rlabel space 16569 4491 16598 4500 1 gnd
rlabel locali 16472 4496 16501 4502 1 gnd
rlabel locali 16259 4496 16288 4502 1 gnd
rlabel nwell 16629 4762 16652 4765 1 vdd
rlabel locali 16208 4607 16230 4622 1 d0
rlabel locali 16475 4792 16504 4798 1 vdd
rlabel locali 16262 4795 16291 4801 1 vdd
rlabel space 16570 4906 16599 4915 1 gnd
rlabel locali 16473 4911 16502 4917 1 gnd
rlabel locali 16260 4911 16289 4917 1 gnd
rlabel nwell 16630 5177 16653 5180 1 vdd
rlabel locali 16209 5022 16231 5037 1 d0
rlabel locali 16476 5207 16505 5213 1 vdd
rlabel locali 16263 5210 16292 5216 1 vdd
rlabel locali 17208 5821 17255 5842 1 d1
rlabel space 17577 5706 17606 5715 1 gnd
rlabel locali 17480 5711 17509 5717 1 gnd
rlabel locali 17267 5711 17296 5717 1 gnd
rlabel nwell 17637 5977 17660 5980 1 vdd
rlabel locali 17483 6007 17512 6013 1 vdd
rlabel locali 17270 6010 17299 6016 1 vdd
rlabel space 16564 5472 16593 5481 1 gnd
rlabel locali 16467 5477 16496 5483 1 gnd
rlabel locali 16254 5477 16283 5483 1 gnd
rlabel nwell 16624 5743 16647 5746 1 vdd
rlabel locali 16203 5588 16225 5603 1 d0
rlabel locali 16470 5773 16499 5779 1 vdd
rlabel locali 16257 5776 16286 5782 1 vdd
rlabel space 16565 5887 16594 5896 1 gnd
rlabel locali 16468 5892 16497 5898 1 gnd
rlabel locali 16255 5892 16284 5898 1 gnd
rlabel nwell 16625 6158 16648 6161 1 vdd
rlabel locali 16204 6003 16226 6018 1 d0
rlabel locali 16471 6188 16500 6194 1 vdd
rlabel locali 16258 6191 16287 6197 1 vdd
rlabel locali 17478 6477 17507 6483 1 vdd
rlabel locali 17691 6474 17720 6480 1 vdd
rlabel nwell 17845 6444 17868 6447 1 vdd
rlabel locali 17475 6178 17504 6184 1 gnd
rlabel locali 17688 6178 17717 6184 1 gnd
rlabel space 17785 6173 17814 6182 1 gnd
rlabel locali 17416 6287 17448 6306 1 d3
rlabel locali 17436 2370 17468 2389 1 d3
rlabel space 17805 2256 17834 2265 1 gnd
rlabel locali 17708 2261 17737 2267 1 gnd
rlabel locali 17495 2261 17524 2267 1 gnd
rlabel nwell 17865 2527 17888 2530 1 vdd
rlabel locali 17711 2557 17740 2563 1 vdd
rlabel locali 17498 2560 17527 2566 1 vdd
rlabel locali 16278 2274 16307 2280 1 vdd
rlabel locali 16491 2271 16520 2277 1 vdd
rlabel locali 16224 2086 16246 2101 1 d0
rlabel nwell 16645 2241 16668 2244 1 vdd
rlabel locali 16275 1975 16304 1981 1 gnd
rlabel locali 16488 1975 16517 1981 1 gnd
rlabel space 16585 1970 16614 1979 1 gnd
rlabel locali 16277 1859 16306 1865 1 vdd
rlabel locali 16490 1856 16519 1862 1 vdd
rlabel locali 16223 1671 16245 1686 1 d0
rlabel nwell 16644 1826 16667 1829 1 vdd
rlabel locali 16274 1560 16303 1566 1 gnd
rlabel locali 16487 1560 16516 1566 1 gnd
rlabel space 16584 1555 16613 1564 1 gnd
rlabel locali 17290 2093 17319 2099 1 vdd
rlabel locali 17503 2090 17532 2096 1 vdd
rlabel nwell 17657 2060 17680 2063 1 vdd
rlabel locali 17287 1794 17316 1800 1 gnd
rlabel locali 17500 1794 17529 1800 1 gnd
rlabel space 17597 1789 17626 1798 1 gnd
rlabel locali 17228 1904 17275 1925 1 d1
rlabel locali 16283 1293 16312 1299 1 vdd
rlabel locali 16496 1290 16525 1296 1 vdd
rlabel locali 16229 1105 16251 1120 1 d0
rlabel nwell 16650 1260 16673 1263 1 vdd
rlabel locali 16280 994 16309 1000 1 gnd
rlabel locali 16493 994 16522 1000 1 gnd
rlabel space 16590 989 16619 998 1 gnd
rlabel locali 16282 878 16311 884 1 vdd
rlabel locali 16495 875 16524 881 1 vdd
rlabel locali 16228 690 16250 705 1 d0
rlabel nwell 16649 845 16672 848 1 vdd
rlabel locali 16279 579 16308 585 1 gnd
rlabel locali 16492 579 16521 585 1 gnd
rlabel space 16589 574 16618 583 1 gnd
rlabel locali 17295 1112 17324 1118 1 vdd
rlabel locali 17508 1109 17537 1115 1 vdd
rlabel nwell 17662 1079 17685 1082 1 vdd
rlabel locali 17292 813 17321 819 1 gnd
rlabel locali 17505 813 17534 819 1 gnd
rlabel space 17602 808 17631 817 1 gnd
rlabel locali 17233 923 17280 944 1 d1
rlabel locali 17345 1532 17374 1538 1 vdd
rlabel locali 17558 1529 17587 1535 1 vdd
rlabel nwell 17712 1499 17735 1502 1 vdd
rlabel locali 17342 1233 17371 1239 1 gnd
rlabel locali 17555 1233 17584 1239 1 gnd
rlabel space 17652 1228 17681 1237 1 gnd
rlabel locali 17288 1344 17311 1359 1 d2
rlabel space 16577 2534 16606 2543 1 gnd
rlabel locali 17276 3304 17299 3319 1 d2
rlabel space 17640 3188 17669 3197 1 gnd
rlabel locali 17543 3193 17572 3199 1 gnd
rlabel locali 17330 3193 17359 3199 1 gnd
rlabel nwell 17700 3459 17723 3462 1 vdd
rlabel locali 17546 3489 17575 3495 1 vdd
rlabel locali 17333 3492 17362 3498 1 vdd
rlabel locali 17221 2883 17268 2904 1 d1
rlabel space 17590 2768 17619 2777 1 gnd
rlabel locali 17493 2773 17522 2779 1 gnd
rlabel locali 17280 2773 17309 2779 1 gnd
rlabel nwell 17650 3039 17673 3042 1 vdd
rlabel locali 17496 3069 17525 3075 1 vdd
rlabel locali 17283 3072 17312 3078 1 vdd
rlabel locali 16480 2539 16509 2545 1 gnd
rlabel locali 16267 2539 16296 2545 1 gnd
rlabel nwell 16637 2805 16660 2808 1 vdd
rlabel locali 16216 2650 16238 2665 1 d0
rlabel locali 16483 2835 16512 2841 1 vdd
rlabel locali 16270 2838 16299 2844 1 vdd
rlabel space 16578 2949 16607 2958 1 gnd
rlabel locali 16481 2954 16510 2960 1 gnd
rlabel locali 16268 2954 16297 2960 1 gnd
rlabel nwell 16638 3220 16661 3223 1 vdd
rlabel locali 16217 3065 16239 3080 1 d0
rlabel locali 16484 3250 16513 3256 1 vdd
rlabel locali 16271 3253 16300 3259 1 vdd
rlabel locali 17216 3864 17263 3885 1 d1
rlabel space 17585 3749 17614 3758 1 gnd
rlabel locali 17488 3754 17517 3760 1 gnd
rlabel locali 17275 3754 17304 3760 1 gnd
rlabel nwell 17645 4020 17668 4023 1 vdd
rlabel locali 17491 4050 17520 4056 1 vdd
rlabel locali 17278 4053 17307 4059 1 vdd
rlabel space 16572 3515 16601 3524 1 gnd
rlabel locali 16475 3520 16504 3526 1 gnd
rlabel locali 16262 3520 16291 3526 1 gnd
rlabel nwell 16632 3786 16655 3789 1 vdd
rlabel locali 16211 3631 16233 3646 1 d0
rlabel locali 16478 3816 16507 3822 1 vdd
rlabel locali 16265 3819 16294 3825 1 vdd
rlabel space 16573 3930 16602 3939 1 gnd
rlabel locali 16476 3935 16505 3941 1 gnd
rlabel locali 16263 3935 16292 3941 1 gnd
rlabel nwell 16633 4201 16656 4204 1 vdd
rlabel locali 16212 4046 16234 4061 1 d0
rlabel locali 16479 4231 16508 4237 1 vdd
rlabel locali 16266 4234 16295 4240 1 vdd
rlabel locali 17573 4485 17602 4491 1 vdd
rlabel locali 17786 4482 17815 4488 1 vdd
rlabel nwell 17940 4452 17963 4455 1 vdd
rlabel locali 17570 4186 17599 4192 1 gnd
rlabel locali 17783 4186 17812 4192 1 gnd
rlabel space 17880 4181 17909 4190 1 gnd
rlabel locali 17515 4291 17537 4315 1 d4
rlabel locali 20837 726 20866 732 5 vdd
rlabel locali 20624 729 20653 735 5 vdd
rlabel locali 20898 905 20920 920 5 d0
rlabel nwell 20476 762 20499 765 5 vdd
rlabel locali 20840 1025 20869 1031 5 gnd
rlabel locali 20627 1025 20656 1031 5 gnd
rlabel space 20530 1027 20559 1036 5 gnd
rlabel locali 20838 1141 20867 1147 5 vdd
rlabel locali 20625 1144 20654 1150 5 vdd
rlabel locali 20899 1320 20921 1335 5 d0
rlabel nwell 20477 1177 20500 1180 5 vdd
rlabel locali 20841 1440 20870 1446 5 gnd
rlabel locali 20628 1440 20657 1446 5 gnd
rlabel space 20531 1442 20560 1451 5 gnd
rlabel locali 19825 907 19854 913 5 vdd
rlabel locali 19612 910 19641 916 5 vdd
rlabel nwell 19464 943 19487 946 5 vdd
rlabel locali 19828 1206 19857 1212 5 gnd
rlabel locali 19615 1206 19644 1212 5 gnd
rlabel space 19518 1208 19547 1217 5 gnd
rlabel locali 19869 1081 19916 1102 5 d1
rlabel locali 20832 1707 20861 1713 5 vdd
rlabel locali 20619 1710 20648 1716 5 vdd
rlabel locali 20893 1886 20915 1901 5 d0
rlabel nwell 20471 1743 20494 1746 5 vdd
rlabel locali 20835 2006 20864 2012 5 gnd
rlabel locali 20622 2006 20651 2012 5 gnd
rlabel space 20525 2008 20554 2017 5 gnd
rlabel locali 20833 2122 20862 2128 5 vdd
rlabel locali 20620 2125 20649 2131 5 vdd
rlabel locali 20894 2301 20916 2316 5 d0
rlabel nwell 20472 2158 20495 2161 5 vdd
rlabel locali 20836 2421 20865 2427 5 gnd
rlabel locali 20623 2421 20652 2427 5 gnd
rlabel locali 19820 1888 19849 1894 5 vdd
rlabel locali 19607 1891 19636 1897 5 vdd
rlabel nwell 19459 1924 19482 1927 5 vdd
rlabel locali 19823 2187 19852 2193 5 gnd
rlabel locali 19610 2187 19639 2193 5 gnd
rlabel space 19513 2189 19542 2198 5 gnd
rlabel locali 19864 2062 19911 2083 5 d1
rlabel locali 19770 1468 19799 1474 5 vdd
rlabel locali 19557 1471 19586 1477 5 vdd
rlabel nwell 19409 1504 19432 1507 5 vdd
rlabel locali 19773 1767 19802 1773 5 gnd
rlabel locali 19560 1767 19589 1773 5 gnd
rlabel space 19463 1769 19492 1778 5 gnd
rlabel locali 19833 1647 19856 1662 5 d2
rlabel space 20526 2423 20555 2432 5 gnd
rlabel locali 19821 3607 19844 3622 5 d2
rlabel space 19451 3729 19480 3738 5 gnd
rlabel locali 19548 3727 19577 3733 5 gnd
rlabel locali 19761 3727 19790 3733 5 gnd
rlabel nwell 19397 3464 19420 3467 5 vdd
rlabel locali 19545 3431 19574 3437 5 vdd
rlabel locali 19758 3428 19787 3434 5 vdd
rlabel locali 19852 4022 19899 4043 5 d1
rlabel space 19501 4149 19530 4158 5 gnd
rlabel locali 19598 4147 19627 4153 5 gnd
rlabel locali 19811 4147 19840 4153 5 gnd
rlabel nwell 19447 3884 19470 3887 5 vdd
rlabel locali 19595 3851 19624 3857 5 vdd
rlabel locali 19808 3848 19837 3854 5 vdd
rlabel space 20514 4383 20543 4392 5 gnd
rlabel locali 20611 4381 20640 4387 5 gnd
rlabel locali 20824 4381 20853 4387 5 gnd
rlabel nwell 20460 4118 20483 4121 5 vdd
rlabel locali 20882 4261 20904 4276 5 d0
rlabel locali 20608 4085 20637 4091 5 vdd
rlabel locali 20821 4082 20850 4088 5 vdd
rlabel space 20513 3968 20542 3977 5 gnd
rlabel locali 20610 3966 20639 3972 5 gnd
rlabel locali 20823 3966 20852 3972 5 gnd
rlabel nwell 20459 3703 20482 3706 5 vdd
rlabel locali 20881 3846 20903 3861 5 d0
rlabel locali 20607 3670 20636 3676 5 vdd
rlabel locali 20820 3667 20849 3673 5 vdd
rlabel locali 19857 3041 19904 3062 5 d1
rlabel space 19506 3168 19535 3177 5 gnd
rlabel locali 19603 3166 19632 3172 5 gnd
rlabel locali 19816 3166 19845 3172 5 gnd
rlabel nwell 19452 2903 19475 2906 5 vdd
rlabel locali 19600 2870 19629 2876 5 vdd
rlabel locali 19813 2867 19842 2873 5 vdd
rlabel space 20519 3402 20548 3411 5 gnd
rlabel locali 20616 3400 20645 3406 5 gnd
rlabel locali 20829 3400 20858 3406 5 gnd
rlabel nwell 20465 3137 20488 3140 5 vdd
rlabel locali 20887 3280 20909 3295 5 d0
rlabel locali 20613 3104 20642 3110 5 vdd
rlabel locali 20826 3101 20855 3107 5 vdd
rlabel space 20518 2987 20547 2996 5 gnd
rlabel locali 20615 2985 20644 2991 5 gnd
rlabel locali 20828 2985 20857 2991 5 gnd
rlabel nwell 20464 2722 20487 2725 5 vdd
rlabel locali 20886 2865 20908 2880 5 d0
rlabel locali 20612 2689 20641 2695 5 vdd
rlabel locali 20825 2686 20854 2692 5 vdd
rlabel locali 19605 2400 19634 2406 5 vdd
rlabel locali 19392 2403 19421 2409 5 vdd
rlabel nwell 19244 2436 19267 2439 5 vdd
rlabel locali 19608 2699 19637 2705 5 gnd
rlabel locali 19395 2699 19424 2705 5 gnd
rlabel space 19298 2701 19327 2710 5 gnd
rlabel locali 19664 2577 19696 2596 5 d3
rlabel locali 19644 6494 19676 6513 5 d3
rlabel space 19278 6618 19307 6627 5 gnd
rlabel locali 19375 6616 19404 6622 5 gnd
rlabel locali 19588 6616 19617 6622 5 gnd
rlabel nwell 19224 6353 19247 6356 5 vdd
rlabel locali 19372 6320 19401 6326 5 vdd
rlabel locali 19585 6317 19614 6323 5 vdd
rlabel locali 20805 6603 20834 6609 5 vdd
rlabel locali 20592 6606 20621 6612 5 vdd
rlabel locali 20866 6782 20888 6797 5 d0
rlabel nwell 20444 6639 20467 6642 5 vdd
rlabel locali 20808 6902 20837 6908 5 gnd
rlabel locali 20595 6902 20624 6908 5 gnd
rlabel space 20498 6904 20527 6913 5 gnd
rlabel locali 20806 7018 20835 7024 5 vdd
rlabel locali 20593 7021 20622 7027 5 vdd
rlabel locali 20867 7197 20889 7212 5 d0
rlabel nwell 20445 7054 20468 7057 5 vdd
rlabel locali 20809 7317 20838 7323 5 gnd
rlabel locali 20596 7317 20625 7323 5 gnd
rlabel space 20499 7319 20528 7328 5 gnd
rlabel locali 19793 6784 19822 6790 5 vdd
rlabel locali 19580 6787 19609 6793 5 vdd
rlabel nwell 19432 6820 19455 6823 5 vdd
rlabel locali 19796 7083 19825 7089 5 gnd
rlabel locali 19583 7083 19612 7089 5 gnd
rlabel space 19486 7085 19515 7094 5 gnd
rlabel locali 19837 6958 19884 6979 5 d1
rlabel locali 20800 7584 20829 7590 5 vdd
rlabel locali 20587 7587 20616 7593 5 vdd
rlabel locali 20861 7763 20883 7778 5 d0
rlabel nwell 20439 7620 20462 7623 5 vdd
rlabel locali 20803 7883 20832 7889 5 gnd
rlabel locali 20590 7883 20619 7889 5 gnd
rlabel space 20493 7885 20522 7894 5 gnd
rlabel locali 20801 7999 20830 8005 5 vdd
rlabel locali 20588 8002 20617 8008 5 vdd
rlabel locali 20862 8178 20884 8193 5 d0
rlabel nwell 20440 8035 20463 8038 5 vdd
rlabel locali 20804 8298 20833 8304 5 gnd
rlabel locali 20591 8298 20620 8304 5 gnd
rlabel space 20494 8300 20523 8309 5 gnd
rlabel locali 19788 7765 19817 7771 5 vdd
rlabel locali 19575 7768 19604 7774 5 vdd
rlabel nwell 19427 7801 19450 7804 5 vdd
rlabel locali 19791 8064 19820 8070 5 gnd
rlabel locali 19578 8064 19607 8070 5 gnd
rlabel space 19481 8066 19510 8075 5 gnd
rlabel locali 19832 7939 19879 7960 5 d1
rlabel locali 20985 8340 21012 8353 5 gnd
rlabel locali 19738 7345 19767 7351 5 vdd
rlabel locali 19525 7348 19554 7354 5 vdd
rlabel nwell 19377 7381 19400 7384 5 vdd
rlabel locali 19741 7644 19770 7650 5 gnd
rlabel locali 19528 7644 19557 7650 5 gnd
rlabel space 19431 7646 19460 7655 5 gnd
rlabel locali 19801 7524 19824 7539 5 d2
rlabel space 20506 6340 20535 6349 5 gnd
rlabel locali 19813 5564 19836 5579 5 d2
rlabel space 19443 5686 19472 5695 5 gnd
rlabel locali 19540 5684 19569 5690 5 gnd
rlabel locali 19753 5684 19782 5690 5 gnd
rlabel nwell 19389 5421 19412 5424 5 vdd
rlabel locali 19537 5388 19566 5394 5 vdd
rlabel locali 19750 5385 19779 5391 5 vdd
rlabel locali 19844 5979 19891 6000 5 d1
rlabel space 19493 6106 19522 6115 5 gnd
rlabel locali 19590 6104 19619 6110 5 gnd
rlabel locali 19803 6104 19832 6110 5 gnd
rlabel nwell 19439 5841 19462 5844 5 vdd
rlabel locali 19587 5808 19616 5814 5 vdd
rlabel locali 19800 5805 19829 5811 5 vdd
rlabel locali 20603 6338 20632 6344 5 gnd
rlabel locali 20816 6338 20845 6344 5 gnd
rlabel nwell 20452 6075 20475 6078 5 vdd
rlabel locali 20874 6218 20896 6233 5 d0
rlabel locali 20600 6042 20629 6048 5 vdd
rlabel locali 20813 6039 20842 6045 5 vdd
rlabel space 20505 5925 20534 5934 5 gnd
rlabel locali 20602 5923 20631 5929 5 gnd
rlabel locali 20815 5923 20844 5929 5 gnd
rlabel nwell 20451 5660 20474 5663 5 vdd
rlabel locali 20873 5803 20895 5818 5 d0
rlabel locali 20599 5627 20628 5633 5 vdd
rlabel locali 20812 5624 20841 5630 5 vdd
rlabel locali 19849 4998 19896 5019 5 d1
rlabel space 19498 5125 19527 5134 5 gnd
rlabel locali 19595 5123 19624 5129 5 gnd
rlabel locali 19808 5123 19837 5129 5 gnd
rlabel nwell 19444 4860 19467 4863 5 vdd
rlabel locali 19592 4827 19621 4833 5 vdd
rlabel locali 19805 4824 19834 4830 5 vdd
rlabel space 20511 5359 20540 5368 5 gnd
rlabel locali 20608 5357 20637 5363 5 gnd
rlabel locali 20821 5357 20850 5363 5 gnd
rlabel nwell 20457 5094 20480 5097 5 vdd
rlabel locali 20879 5237 20901 5252 5 d0
rlabel locali 20605 5061 20634 5067 5 vdd
rlabel locali 20818 5058 20847 5064 5 vdd
rlabel space 20510 4944 20539 4953 5 gnd
rlabel locali 20607 4942 20636 4948 5 gnd
rlabel locali 20820 4942 20849 4948 5 gnd
rlabel nwell 20456 4679 20479 4682 5 vdd
rlabel locali 20878 4822 20900 4837 5 d0
rlabel locali 20604 4646 20633 4652 5 vdd
rlabel locali 20817 4643 20846 4649 5 vdd
rlabel locali 19510 4392 19539 4398 5 vdd
rlabel locali 19297 4395 19326 4401 5 vdd
rlabel nwell 19149 4428 19172 4431 5 vdd
rlabel locali 19513 4691 19542 4697 5 gnd
rlabel locali 19300 4691 19329 4697 5 gnd
rlabel space 19203 4693 19232 4702 5 gnd
rlabel locali 19575 4568 19597 4592 5 d4
rlabel locali 17685 397 17714 403 1 vdd
rlabel locali 17898 394 17927 400 1 vdd
rlabel nwell 18052 364 18075 367 1 vdd
rlabel locali 17682 98 17711 104 1 gnd
rlabel locali 17895 98 17924 104 1 gnd
rlabel space 17992 93 18021 102 1 gnd
rlabel locali 17627 206 17651 223 1 d5
rlabel locali 15494 330 15523 336 1 vdd
rlabel locali 15707 327 15736 333 1 vdd
rlabel nwell 15861 297 15884 300 1 vdd
rlabel locali 15491 31 15520 37 1 gnd
rlabel locali 15704 31 15733 37 1 gnd
rlabel space 15801 26 15830 35 1 gnd
rlabel locali 15438 137 15457 157 1 d6
rlabel locali 10094 315 10123 321 1 vdd
rlabel locali 10307 312 10336 318 1 vdd
rlabel locali 10670 162 10692 177 1 vout
rlabel nwell 10461 282 10484 285 1 vdd
rlabel locali 10091 16 10120 22 1 gnd
rlabel locali 10304 16 10333 22 1 gnd
rlabel space 10401 11 10430 20 1 gnd
rlabel locali 10038 128 10051 143 1 d7
<< end >>
