* SPICE3 file created from 9bit_DAC.ext - technology: sky130A

*.option scale=10000u

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_8352_5673# a_8456_4922# a_8411_4935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1 a_22931_906# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2 a_153_1298# a_153_1016# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3 a_12310_1924# a_12097_1924# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4 a_16058_7861# a_16547_7961# a_16755_7961# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5 a_24608_6887# a_25666_7108# a_25617_7298# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6 a_27168_6943# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7 a_11283_5041# a_11070_5041# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8 a_40557_5895# a_41615_6116# a_41570_6129# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9 a_1798_5391# a_1684_5272# a_1892_5272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X10 a_39066_4810# a_38853_4810# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X11 a_14815_2439# a_14818_1847# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X12 gnd d2 a_40748_7422# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X13 a_39056_6258# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X14 gnd a_9692_2220# a_9484_2220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X15 a_6093_7538# a_6898_7772# a_7067_7330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X16 a_16559_6001# a_16346_6001# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X17 a_22111_4589# a_21898_4589# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X18 a_10814_1306# a_11303_1124# a_11511_1124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X19 a_38068_1640# a_37855_1640# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X20 a_28180_6762# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X21 a_38265_4015# a_37844_4015# a_37568_4197# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X22 a_4133_5933# a_4390_5743# a_3121_6114# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X23 a_32580_1095# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X24 a_29697_2659# a_29911_1537# a_29862_1727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X25 vdd d3 a_40615_2477# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X26 gnd a_30137_7834# a_29929_7834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X27 a_27387_5549# a_27174_5549# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X28 vdd d3 a_29934_6386# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X29 a_17571_5820# a_17358_5820# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X30 a_622_5033# a_409_5033# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X31 a_3146_1216# a_4207_845# a_4162_858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X32 a_37856_2055# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X33 a_13492_4709# a_13636_2527# a_13591_2540# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X34 a_33555_7772# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X35 a_38250_6951# a_37829_6951# a_37553_6851# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X36 a_5906_4036# a_5693_4036# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X37 gnd d2 a_19290_1574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X38 a_16787_2084# a_17591_1903# a_17760_1461# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X39 a_17728_7338# a_17346_7780# a_16755_7961# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X40 gnd a_20320_7690# a_20112_7690# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X41 a_37580_1955# a_37582_1856# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X42 a_19067_5924# a_20125_6145# a_20080_6158# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X43 vdd d0 a_4395_4762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X44 a_7322_4287# a_7213_4287# a_7421_4287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X45 a_6094_7953# a_5673_7953# a_5397_7853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X46 gnd a_15044_6730# a_14836_6730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X47 gnd a_19345_1013# a_19137_1013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X48 a_23347_2354# a_23134_2354# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X49 a_9408_7306# a_9665_7116# a_8399_6895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X50 a_25633_5161# a_25886_5148# a_24620_4927# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X51 a_15904_140# a_17773_207# a_18095_207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X52 a_5422_3237# a_5422_2955# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X53 a_16572_3063# a_16359_3063# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X54 a_8427_1195# a_9488_824# a_9443_837# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X55 a_24635_1991# a_24888_1978# a_24585_1571# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X56 a_14791_6743# a_14787_6920# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X57 a_16366_2084# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X58 a_30929_2204# a_31182_2191# a_29916_1970# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X59 a_40550_6874# a_40803_6861# a_40491_7612# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X60 a_16791_688# a_17596_922# a_17755_1342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X61 a_26832_103# a_26411_103# a_26733_103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X62 a_7082_3294# a_6973_3294# a_7181_3294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X63 a_32983_3621# a_32562_3621# a_32294_3451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X64 a_26411_103# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X65 a_8211_2511# a_8464_2498# a_8112_4680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X66 a_11490_4626# a_12295_4860# a_12454_5280# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X67 a_37582_1856# a_37587_1470# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X68 a_16766_5586# a_17571_5820# a_17740_5378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X69 a_12467_3442# a_12085_3884# a_11494_4065# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X70 a_29921_989# a_30979_1210# a_30930_1400# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X71 a_9415_6327# a_9418_5735# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X72 a_40511_3695# a_40615_2944# a_40570_2957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X73 vdd d2 a_40748_7422# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X74 a_11479_7001# a_11058_7001# a_10782_6901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X75 vdd a_36534_6701# a_36326_6701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X76 vdd a_9692_2220# a_9484_2220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X77 a_40515_3518# a_40610_3925# a_40561_4115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X78 gnd d0 a_15072_2249# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X79 a_38037_7932# a_37824_7932# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X80 a_22307_6549# a_21886_6549# a_21620_6381# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X81 a_16792_1103# a_16371_1103# a_16095_1003# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X82 a_12442_7240# a_12070_6820# a_11478_6586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X83 vdd a_4378_7703# a_4170_7703# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X84 a_16552_6980# a_16339_6980# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X85 a_11493_3650# a_11072_3650# a_10804_3480# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X86 gnd d1 a_35517_7863# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X87 a_818_6993# a_397_6993# a_121_7175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X88 a_41573_3934# a_41583_3191# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X89 vdd d2 a_19290_1574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X90 a_22334_1653# a_23139_1887# a_23308_1445# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X91 gnd a_29934_6386# a_29726_6386# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X92 a_6702_4831# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X93 a_36310_1429# a_36567_1239# a_35301_1018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X94 a_32963_7538# a_32542_7538# a_32269_7754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X95 gnd d0 a_36529_7682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X96 vdd a_15044_6730# a_14836_6730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X97 a_22315_5985# a_21894_5985# a_21618_5885# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X98 gnd d0 a_9679_3765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X99 vdd a_19345_1013# a_19137_1013# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X100 a_5704_1661# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X101 a_24553_7448# a_24648_7855# a_24599_8045# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X102 a_39116_5230# a_38903_5230# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X103 a_832_3642# a_411_3642# a_138_3858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X104 a_16547_7961# a_16334_7961# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X105 gnd a_4395_4762# a_4187_4762# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X106 a_19056_7080# a_20117_6709# a_20068_6899# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X107 vdd d1 a_24861_6874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X108 a_32560_5012# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X109 a_14814_2024# a_14824_1281# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X110 a_8426_1999# a_9484_2220# a_9435_2410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X111 a_24599_8045# a_25660_7674# a_25611_7864# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X112 a_23174_5243# a_22961_5243# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X113 a_29866_1550# a_29961_1957# a_29912_2147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X114 gnd d1 a_14027_7892# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X115 a_16772_5020# a_16351_5020# a_16075_5202# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X116 a_32559_4597# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X117 gnd a_31170_4151# a_30962_4151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X118 a_32788_2076# a_32575_2076# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X119 a_14820_1458# a_15077_1268# a_13811_1047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X120 a_11473_7567# a_11052_7567# a_10779_7783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X121 gnd d1 a_19340_1994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X122 a_28703_4258# a_28490_4258# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X123 a_27596_5964# a_27175_5964# a_26899_6146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X124 a_29921_989# a_30979_1210# a_30934_1223# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X125 a_33642_1334# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X126 a_1818_1474# a_1436_1916# a_845_2097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X127 a_37562_5773# a_38048_5557# a_38256_5557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X128 a_11070_5041# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X129 gnd d0 a_36566_824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X130 a_5342_132# a_10395_125# a_10603_125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X131 a_20084_4762# a_20337_4749# a_19068_5120# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X132 a_32289_4432# a_32772_4597# a_32980_4597# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X133 vdd d0 a_20358_1247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X134 a_29912_2147# a_30169_1957# a_29866_1550# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X135 a_27380_6528# a_27167_6528# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X136 a_25627_5727# a_25880_5714# a_24611_6085# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X137 a_34031_7211# a_33610_7211# a_33932_7211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X138 a_8191_6428# a_8444_6415# a_8116_4503# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X139 a_27174_5549# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X140 vdd d0 a_25888_3757# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X141 a_28463_3265# a_28250_3265# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X142 a_24636_1187# a_25697_816# a_25648_1006# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X143 a_2252_220# a_5134_132# a_5342_132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X144 vdd a_29934_6386# a_29726_6386# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X145 a_34051_3294# a_34008_2362# a_34192_4287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X146 gnd d0 a_25881_6129# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X147 a_10796_5437# a_11277_5607# a_11485_5607# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X148 vdd d0 a_36529_7682# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X149 a_5693_4036# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X150 vdd d0 a_9679_3765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X151 a_32306_896# a_32792_680# a_33000_680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X152 a_17634_3302# a_17421_3302# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X153 gnd d0 a_15076_853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X154 vdd a_4395_4762# a_4187_4762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X155 a_35246_1579# a_35499_1566# a_35077_2688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X156 a_2926_2709# a_3140_1587# a_3095_1600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X157 a_20887_n19# a_20674_n19# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X158 a_23134_2354# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X159 a_24628_2970# a_24881_2957# a_24569_3708# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X160 a_35246_1579# a_35341_1986# a_35296_1999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X161 a_8426_1999# a_9484_2220# a_9439_2233# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X162 a_24599_8045# a_25660_7674# a_25615_7687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X163 a_37555_7347# a_37553_7133# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X164 a_14807_4222# a_15060_4209# a_13794_3988# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X165 a_12541_7240# a_12120_7240# a_12442_7240# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X166 a_24325_4495# a_24445_6407# a_24396_6597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X167 a_32543_7953# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X168 a_16063_6880# a_16065_6781# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X169 vdd a_31170_4151# a_30962_4151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X170 gnd d0 a_31166_4712# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X171 a_37582_2451# a_38061_2619# a_38269_2619# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X172 gnd d0 a_41836_3178# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X173 a_28683_1305# a_28262_1305# a_28589_1424# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X174 a_21611_6864# a_22100_6964# a_22308_6964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X175 a_13799_3007# a_14857_3228# a_14808_3418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X176 a_10816_925# a_11302_709# a_11510_709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X177 a_4153_2016# a_4410_1826# a_3141_2197# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X178 a_20076_6335# a_20079_5743# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X179 gnd d1 a_40815_4901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X180 a_30929_985# a_26933_666# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X181 a_23139_1887# a_22926_1887# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X182 a_16759_6565# a_17564_6799# a_17723_7219# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X183 a_34043_5251# a_33988_6279# a_34196_6279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X184 a_33957_3413# a_33575_3855# a_32984_4036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X185 a_32969_6972# a_32548_6972# a_32272_6872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X186 a_29842_5644# a_29946_4893# a_29901_4906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X187 gnd d0 a_20341_4188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X188 a_21652_687# a_22131_672# a_22339_672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X189 a_13732_5702# a_13836_4951# a_13787_5141# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X190 a_16085_3459# a_16566_3629# a_16774_3629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X191 a_23288_5362# a_23174_5243# a_23382_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X192 a_25636_2966# a_25648_2225# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X193 a_9407_8110# a_9660_8097# a_8394_7876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X194 a_604_7559# a_391_7559# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X195 a_39476_178# a_39263_178# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X196 a_27583_7509# a_28388_7743# a_28557_7301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X197 a_3126_5133# a_4187_4762# a_4138_4952# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X198 a_23124_4823# a_22911_4823# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X199 a_30905_6298# a_31162_6108# a_29896_5887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X200 a_21623_5186# a_21623_4904# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X201 a_16078_4226# a_16078_3944# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X202 a_25623_5904# a_25880_5714# a_24611_6085# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X203 gnd d0 a_9676_4741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X204 a_22126_1653# a_21913_1653# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X205 gnd a_15072_2249# a_14864_2249# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X206 a_37824_7932# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X207 a_32768_5993# a_32555_5993# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X208 vdd d1 a_19325_4930# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X209 a_22323_4028# a_21902_4028# a_21626_4210# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X210 a_16065_6781# a_16072_6397# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X211 a_8187_6605# a_8444_6415# a_8116_4503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X212 a_41579_3368# a_41836_3178# a_40570_2957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X213 gnd d1 a_19320_5911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X214 a_11511_1124# a_12315_943# a_12474_1363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X215 a_33780_5812# a_33567_5812# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X216 a_32304_1277# a_32793_1095# a_33001_1095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X217 a_30934_1223# a_30930_1400# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X218 a_21914_2068# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X219 gnd a_35517_7863# a_35309_7863# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X220 a_37560_5872# a_37562_5773# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X221 a_35061_6428# a_35259_7443# a_35210_7633# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X222 vdd d3 a_24673_2490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X223 a_23742_191# a_23321_191# a_23630_4279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X224 a_27584_7924# a_27163_7924# a_26887_7824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X225 a_39061_5791# a_38848_5791# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X226 a_33944_5251# a_33835_5251# a_34043_5251# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X227 a_10799_3866# a_10804_3480# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X228 a_35242_1756# a_35499_1566# a_35077_2688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X229 a_6985_1334# a_6772_1334# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X230 a_17987_6287# a_17566_6287# a_17834_5259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X231 a_23321_191# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X232 a_20072_6722# a_20068_6899# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X233 vdd a_8679_1986# a_8471_1986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X234 gnd a_9672_6137# a_9464_6137# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X235 a_35280_4136# a_35537_3946# a_35234_3539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X236 vdd d1 a_24893_997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X237 a_16334_7961# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X238 a_11278_6022# a_11065_6022# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X239 a_38277_2055# a_39081_1874# a_39250_1432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X240 a_26733_103# a_28602_170# a_28924_170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X241 a_28602_170# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X242 a_1892_5272# a_1471_5272# a_1793_5272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X243 vdd d0 a_31166_4712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X244 a_39473_4266# a_39364_4266# a_39572_4266# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X245 a_8415_3155# a_9476_2784# a_9427_2974# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X246 a_28413_2845# a_28200_2845# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X247 a_32781_3055# a_32568_3055# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X248 a_22106_5570# a_21893_5570# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X249 a_8116_4503# a_8369_4490# a_7434_199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X250 gnd d1 a_8672_2965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X251 gnd a_14027_7892# a_13819_7892# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X252 a_12290_5841# a_12077_5841# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X253 a_28207_1866# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X254 a_32575_2076# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X255 a_29701_2482# a_29954_2469# a_29602_4651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X256 a_30930_1400# a_30933_808# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X257 a_37562_5773# a_37567_5387# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X258 a_28490_4258# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X259 a_10809_2287# a_10809_2005# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X260 a_1801_3315# a_1429_2895# a_838_3076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X261 a_18868_2696# a_19082_1574# a_19033_1764# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X262 a_3095_1600# a_3190_2007# a_3145_2020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X263 a_35226_5496# a_35321_5903# a_35276_5916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X264 a_13790_4165# a_14047_3975# a_13744_3568# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X265 a_27199_651# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X266 a_14787_8139# a_15040_8126# a_13774_7905# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X267 a_3126_5133# a_4187_4762# a_4142_4775# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X268 gnd a_36566_824# a_36358_824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X269 vdd d0 a_9676_4741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X270 a_5886_7953# a_5673_7953# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X271 a_12913_228# a_15795_140# a_10504_125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X272 a_39074_2853# a_38861_2853# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X273 a_5399_7754# a_5885_7538# a_6093_7538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X274 vdd a_20358_1247# a_20150_1247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X275 a_16567_4044# a_16354_4044# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X276 a_33001_1095# a_32580_1095# a_32304_1277# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X277 a_41553_7851# a_41563_7108# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X278 a_30901_6685# a_31154_6672# a_29885_7043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X279 gnd d4 a_19030_4498# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X280 gnd d1 a_40818_3925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X281 a_31672_96# d7 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X282 a_4142_4775# a_4138_4952# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X283 a_28250_3265# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X284 a_17755_1342# a_17383_922# a_16791_688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X285 a_17383_922# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X286 a_35061_6428# a_35259_7443# a_35214_7456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X287 a_40515_3518# a_40768_3505# a_40362_2490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X288 a_38282_1074# a_37861_1074# a_37585_974# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X289 a_17723_7219# a_17614_7219# a_17822_7219# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X290 gnd d0 a_41830_3744# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X291 a_29916_1970# a_30974_2191# a_30925_2381# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X292 a_8390_8053# a_8647_7863# a_8344_7456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X293 a_16552_6980# a_16339_6980# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X294 a_17421_3302# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X295 a_39218_7309# a_38836_7751# a_38244_7517# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X296 a_5891_6972# a_5678_6972# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X297 a_26909_4403# a_27392_4568# a_27600_4568# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X298 gnd a_15076_853# a_14868_853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X299 a_6126_2076# a_5705_2076# a_5429_1976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X300 a_14794_5941# a_14804_5198# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X301 vdd d1 a_24876_3938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X302 a_8415_3155# a_9476_2784# a_9431_2797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X303 a_11511_1124# a_11090_1124# a_10814_1306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X304 a_813_7974# a_392_7974# a_116_8156# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X305 a_9406_7695# a_9402_7872# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X306 a_32995_1661# a_33800_1895# a_33969_1453# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X307 a_12447_7359# a_12065_7801# a_11474_7982# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X308 a_40338_6584# a_40552_5462# a_40503_5652# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X309 a_32284_5194# a_32773_5012# a_32981_5012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X310 a_37840_4576# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X311 a_16787_2084# a_16366_2084# a_16090_2266# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X312 gnd a_41836_3178# a_41628_3178# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X313 gnd d0 a_25868_7674# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X314 gnd a_31166_4712# a_30958_4712# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X315 vdd a_3383_4943# a_3175_4943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X316 gnd a_36550_4180# a_36342_4180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X317 a_32981_5012# a_33785_4831# a_33944_5251# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X318 gnd a_40780_1545# a_40572_1545# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X319 a_18868_2696# a_19082_1574# a_19037_1587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X320 gnd a_40815_4901# a_40607_4901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X321 a_12801_4316# a_12380_4316# a_12702_4316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X322 a_10789_6204# a_11278_6022# a_11486_6022# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X323 vdd a_8659_5903# a_8451_5903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X324 a_19025_3547# a_19278_3534# a_18872_2519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X325 a_32301_1877# a_32787_1661# a_32995_1661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X326 a_40573_2155# a_40830_1965# a_40527_1558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X327 a_14783_8316# a_15040_8126# a_13774_7905# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X328 a_26904_4883# a_26906_4784# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X329 a_33982_199# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X330 a_19025_3547# a_19120_3954# a_19075_3967# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X331 a_391_7559# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X332 a_1441_935# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X333 vdd d0 a_41816_7095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X334 a_30897_6862# a_31154_6672# a_29885_7043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X335 a_32555_5993# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X336 vdd a_19325_4930# a_19117_4930# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X337 a_128_5914# a_617_6014# a_825_6014# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X338 a_34982_4680# a_35239_4490# a_34304_199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X339 a_12561_3323# a_12140_3323# a_12462_3323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X340 vdd d0 a_20321_8105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X341 vdd d0 a_41830_3744# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X342 a_32579_680# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X343 a_36309_1014# a_32313_695# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X344 a_1459_7232# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X345 a_1429_2895# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X346 a_629_2661# a_416_2661# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X347 gnd d3 a_40615_2477# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X348 a_37573_3216# a_38062_3034# a_38270_3034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X349 a_19075_3967# a_20133_4188# a_20088_4201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X350 a_14807_3003# a_14819_2262# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X351 a_13770_8082# a_14027_7892# a_13724_7485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X352 a_13790_4165# a_14851_3794# a_14806_3807# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X353 a_13811_1047# a_14869_1268# a_14824_1281# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X354 vdd a_8672_2965# a_8464_2965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X355 a_13492_4709# a_13636_2527# a_13587_2717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X356 a_6772_1334# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X357 a_38270_3034# a_39074_2853# a_39233_3273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X358 a_11271_7001# a_11058_7001# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X359 a_32286_5408# a_32767_5578# a_32975_5578# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X360 a_16078_4226# a_16567_4044# a_16775_4044# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X361 a_27188_3026# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X362 vdd d0 a_25869_8089# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X363 a_32980_4597# a_32559_4597# a_32289_4432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X364 vdd a_24893_997# a_24685_997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X365 a_39124_3273# a_38911_3273# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X366 a_11065_6022# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X367 a_30917_4164# a_30913_4341# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X368 a_10802_2984# a_11291_3084# a_11499_3084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X369 a_6114_4036# a_6918_3855# a_7087_3413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X370 a_1654_935# a_1441_935# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X371 a_40338_6584# a_40552_5462# a_40507_5475# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X372 a_28200_2845# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X373 vdd d0 a_25868_7674# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X374 vdd a_31166_4712# a_30958_4712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X375 a_27375_7509# a_27162_7509# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X376 a_40495_7435# a_40748_7422# a_40342_6407# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X377 vdd a_36550_4180# a_36342_4180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X378 gnd d0 a_36546_4741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X379 a_642_1116# a_429_1116# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X380 vdd a_40780_1545# a_40572_1545# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X381 a_40358_2667# a_40615_2477# a_40263_4659# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X382 a_7181_3294# a_7138_2362# a_7322_4287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X383 a_5342_132# a_4921_132# a_5243_132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X384 a_19021_3724# a_19278_3534# a_18872_2519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X385 a_25616_6883# a_25628_6142# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X386 vdd d1 a_30169_1957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X387 a_6935_914# a_6722_914# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X388 a_8376_1579# a_8629_1566# a_8207_2688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X389 a_35289_2978# a_36347_3199# a_36298_3389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X390 a_8395_7072# a_9456_6701# a_9411_6714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X391 a_24616_5104# a_25677_4733# a_25628_4923# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X392 a_9432_3212# a_9428_3389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X393 a_38249_6536# a_39054_6770# a_39213_7190# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X394 gnd d1 a_24873_4914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X395 a_39585_178# a_40312_4469# a_40267_4482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X396 a_37843_3600# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X397 a_2926_2709# a_3183_2519# a_2831_4701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X398 a_28651_7182# a_28608_6250# a_28816_6250# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X399 a_16766_5586# a_16345_5586# a_16077_5416# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X400 gnd d0 a_31161_5693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X401 a_30913_4341# a_30916_3749# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X402 a_39344_1313# a_38923_1313# a_39250_1432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X403 a_5673_7953# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X404 a_36297_4193# a_36293_4370# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X405 a_36285_6327# a_36542_6137# a_35276_5916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X406 gnd d0 a_15056_4770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X407 a_13794_3988# a_14852_4209# a_14803_4399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X408 a_16354_4044# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X409 gnd a_40818_3925# a_40610_3925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X410 a_10395_125# a_10182_125# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X411 a_18848_6613# a_19062_5491# a_19017_5504# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X412 a_10779_7783# a_10784_7397# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X413 a_29846_5467# a_29941_5874# a_29896_5887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X414 a_12702_4316# a_12305_2391# a_12573_1363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X415 a_25637_3381# a_25894_3191# a_24628_2970# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X416 gnd a_30099_5454# a_29891_5454# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X417 a_9428_3389# a_9431_2797# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X418 a_36314_1252# a_36567_1239# a_35301_1018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X419 a_11297_1690# a_11084_1690# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X420 a_4125_7716# a_4121_7893# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X421 a_23119_5804# a_22906_5804# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X422 vdd a_24876_3938# a_24668_3938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X423 a_29606_4474# a_29859_4461# a_28924_170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X424 a_32567_2640# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X425 a_40491_7612# a_40748_7422# a_40342_6407# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X426 a_143_2877# a_629_2661# a_837_2661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X427 a_29896_5887# a_30954_6108# a_30909_6121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X428 a_1409_6812# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X429 vdd d0 a_36546_4741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X430 a_3141_2197# a_4202_1826# a_4153_2016# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X431 gnd a_25868_7674# a_25660_7674# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X432 a_38245_7932# a_37824_7932# a_37548_7832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X433 a_21886_6549# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X434 a_23534_191# a_23321_191# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X435 a_16779_2648# a_16358_2648# a_16085_2864# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X436 a_26919_1947# a_26921_1848# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X437 a_21645_1483# a_21643_1269# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X438 a_8372_1756# a_8629_1566# a_8207_2688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X439 a_39238_3392# a_39124_3273# a_39332_3273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X440 a_24616_5104# a_25677_4733# a_25632_4746# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X441 a_37570_3816# a_38056_3600# a_38264_3600# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X442 a_10504_125# a_15582_140# a_12913_228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X443 a_14824_1281# a_15077_1268# a_13811_1047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X444 a_10784_6802# a_11270_6586# a_11478_6586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X445 a_28812_4258# a_28703_4258# a_28911_4258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X446 a_15582_140# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X447 a_4138_6171# a_4134_6348# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X448 a_21894_5985# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X449 a_26889_7725# a_27375_7509# a_27583_7509# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X450 vdd a_41816_7095# a_41608_7095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X451 a_23132_2866# a_22919_2866# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X452 vdd d0 a_15056_4770# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X453 a_23194_1326# a_22981_1326# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X454 vdd a_36530_8097# a_36322_8097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X455 a_40545_7855# a_40798_7842# a_40495_7435# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X456 a_16563_4605# a_16350_4605# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X457 a_24604_7064# a_24861_6874# a_24549_7625# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X458 a_28408_3826# a_28195_3826# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X459 vdd d0 a_36566_824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X460 a_130_6410# a_609_6578# a_817_6578# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X461 a_36281_6714# a_36534_6701# a_35265_7072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X462 a_3129_4157# a_3386_3967# a_3083_3560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X463 a_36309_1014# a_36566_824# a_35297_1195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X464 gnd d0 a_20358_1247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X465 a_16075_4920# a_16077_4821# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X466 a_5424_3451# a_5422_3237# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X467 a_22340_1087# a_21919_1087# a_21643_987# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X468 a_26921_1848# a_26926_1462# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X469 a_7138_2362# a_6925_2362# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X470 a_9424_5169# a_9677_5156# a_8411_4935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X471 a_416_2661# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X472 a_35269_6895# a_36327_7116# a_36278_7306# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X473 gnd d0 a_25888_3757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X474 a_5910_2640# a_5697_2640# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X475 a_12315_943# a_12102_943# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X476 a_27616_2047# a_27195_2047# a_26919_1947# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X477 a_8426_1999# a_8679_1986# a_8376_1579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X478 a_4125_7716# a_4378_7703# a_3109_8074# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X479 a_23276_7322# a_22894_7764# a_22302_7530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X480 vdd a_30099_5454# a_29891_5454# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X481 a_35234_3539# a_35329_3946# a_35280_4136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X482 a_37548_8114# a_37548_7832# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X483 a_16097_1499# a_16095_1285# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X484 gnd d0 a_41811_8076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X485 a_37555_7347# a_38036_7517# a_38244_7517# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X486 gnd d4 a_8369_4490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X487 gnd a_9696_824# a_9488_824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X488 a_29602_4651# a_29859_4461# a_28924_170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X489 a_13744_3568# a_13839_3975# a_13794_3988# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X490 a_9438_1818# a_9691_1805# a_8422_2176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X491 a_13774_7905# a_14832_8126# a_14783_8316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X492 a_10796_5437# a_10794_5223# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X493 a_35280_4136# a_36341_3765# a_36292_3955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X494 a_10782_7183# a_10782_6901# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X495 a_845_2097# a_1649_1916# a_1818_1474# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X496 vdd d3 a_40595_6394# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X497 a_30912_3926# a_30922_3183# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X498 vdd a_25868_7674# a_25660_7674# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X499 a_27162_7509# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X500 a_26889_7725# a_26894_7339# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X501 a_29885_7043# a_30946_6672# a_30897_6862# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X502 a_16077_4821# a_16080_4440# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X503 gnd a_36546_4741# a_36338_4741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X504 gnd d1 a_30142_6853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X505 a_20093_3220# a_20089_3397# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X506 a_38277_2055# a_37856_2055# a_37580_2237# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X507 a_7118_6279# a_6905_6279# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X508 a_37860_659# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X509 a_13752_1785# a_14009_1595# a_13587_2717# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X510 a_6098_6557# a_5677_6557# a_5411_6389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X511 a_33773_6791# a_33560_6791# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X512 gnd a_4390_5743# a_4182_5743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X513 gnd a_30149_5874# a_29941_5874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X514 a_22315_5985# a_23119_5804# a_23288_5362# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X515 a_20088_2982# a_20345_2792# a_19076_3163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X516 a_41577_3757# a_41573_3934# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X517 a_849_701# a_1654_935# a_1813_1355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X518 gnd a_24873_4914# a_24665_4914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X519 a_38262_4991# a_37841_4991# a_37565_4891# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X520 a_34291_4287# a_33870_4287# a_34192_4287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X521 a_153_1016# a_155_917# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X522 a_1617_7793# a_1404_7793# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X523 a_5918_2076# a_5705_2076# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X524 vdd a_40835_984# a_40627_984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X525 a_38061_2619# a_37848_2619# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X526 a_3059_7654# a_3163_6903# a_3114_7093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X527 a_6106_5993# a_5685_5993# a_5409_5893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X528 gnd a_15056_4770# a_14848_4770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X529 a_6930_1895# a_6717_1895# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X530 a_26899_6146# a_26899_5864# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X531 a_22919_2866# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X532 a_8344_7456# a_8439_7863# a_8390_8053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X533 a_32279_6175# a_32279_5893# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X534 a_9420_5346# a_9677_5156# a_8411_4935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X535 a_33969_1453# a_33587_1895# a_32996_2076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X536 a_35269_6895# a_36327_7116# a_36282_7129# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X537 a_40342_6407# a_40595_6394# a_40267_4482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X538 gnd a_3391_2986# a_3183_2986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X539 a_14818_1847# a_14814_2024# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X540 a_41583_3191# a_41836_3178# a_40570_2957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X541 a_21631_3229# a_22120_3047# a_22328_3047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X542 vdd d1 a_8652_6882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X543 vdd d0 a_41811_8076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X544 a_32975_5578# a_33780_5812# a_33949_5370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X545 a_13806_2028# a_14059_2015# a_13756_1608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X546 a_34051_3294# a_33630_3294# a_33952_3294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X547 a_8390_8053# a_9451_7682# a_9402_7872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X548 a_17559_7780# a_17346_7780# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X549 a_40562_4914# a_40815_4901# a_40503_5652# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X550 a_33944_5251# a_33572_4831# a_32980_4597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X551 a_11084_1690# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X552 a_41590_2212# a_41586_2389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X553 vdd d0 a_4384_7137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X554 a_23112_6783# a_22899_6783# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X555 a_20996_n19# a_31672_96# a_26832_103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X556 a_32995_1661# a_32574_1661# a_32306_1491# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X557 a_13774_7905# a_14832_8126# a_14787_8139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X558 a_19001_7641# a_19105_6890# a_19056_7080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X559 gnd a_9679_3765# a_9471_3765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X560 a_27604_4007# a_28408_3826# a_28577_3384# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X561 a_35280_4136# a_36341_3765# a_36296_3778# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X562 a_22114_3613# a_21901_3613# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X563 a_11510_709# a_11089_709# a_10823_724# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X564 a_34982_4680# a_35126_2498# a_35077_2688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X565 a_1798_5391# a_1416_5833# a_824_5599# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X566 a_37844_4015# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X567 a_12479_1482# a_12097_1924# a_11506_2105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X568 a_3130_4956# a_3383_4943# a_3071_5694# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X569 a_22320_5004# a_21899_5004# a_21623_4904# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X570 a_40562_4914# a_41620_5135# a_41571_5325# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X571 vdd a_36546_4741# a_36338_4741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X572 gnd d0 a_31181_1776# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X573 a_29885_7043# a_30946_6672# a_30901_6685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X574 a_21902_4028# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X575 a_20093_3220# a_20346_3207# a_19080_2986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X576 a_32292_2955# a_32781_3055# a_32989_3055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X577 a_21645_888# a_21652_687# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X578 a_40527_1558# a_40622_1965# a_40573_2155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X579 a_38049_5972# a_37836_5972# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X580 vdd d1 a_40798_7842# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X581 a_22319_4589# a_21898_4589# a_21628_4424# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X582 vdd a_4390_5743# a_4182_5743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X583 a_12454_5280# a_12082_4860# a_11490_4626# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X584 a_5422_2955# a_5424_2856# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X585 a_33969_1453# a_33855_1334# a_34063_1334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X586 a_11505_1690# a_11084_1690# a_10816_1520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X587 a_13724_7485# a_13819_7892# a_13774_7905# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X588 a_9418_5735# a_9671_5722# a_8402_6093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X589 a_17740_5378# a_17358_5820# a_16766_5586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X590 a_10797_3965# a_11286_4065# a_11494_4065# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X591 vdd d4 a_35239_4490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X592 a_24416_2680# a_24673_2490# a_24321_4672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X593 a_5399_7754# a_5404_7368# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X594 a_38264_3600# a_39069_3834# a_39238_3392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X595 a_8427_1195# a_9488_824# a_9439_1014# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X596 a_37553_7133# a_38042_6951# a_38250_6951# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X597 a_36304_1995# a_36561_1805# a_35292_2176# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X598 a_11298_2105# a_11085_2105# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X599 a_32975_5578# a_32554_5578# a_32281_5794# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X600 a_19072_4943# a_19325_4930# a_19013_5681# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X601 a_26912_3208# a_26912_2926# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X602 a_1880_7232# a_1459_7232# a_1786_7351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X603 gnd d0 a_9691_1805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X604 a_32292_3237# a_32292_2955# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X605 a_19072_4943# a_20130_5164# a_20081_5354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X606 vdd a_15056_4770# a_14848_4770# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X607 a_16350_4605# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X608 a_24585_1571# a_24680_1978# a_24635_1991# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X609 a_1644_2383# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X610 a_7161_7211# a_7118_6279# a_7326_6279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X611 a_28195_3826# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X612 a_12310_1924# a_12097_1924# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X613 a_16058_8143# a_16547_7961# a_16755_7961# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X614 a_27168_6943# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X615 a_9418_5735# a_9414_5912# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X616 gnd a_20358_1247# a_20150_1247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X617 a_8419_2978# a_8672_2965# a_8360_3716# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X618 a_13802_2205# a_14059_2015# a_13756_1608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X619 a_408_4618# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X620 gnd d0 a_31175_3170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X621 a_637_2097# a_424_2097# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X622 a_26921_2443# a_27400_2611# a_27608_2611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X623 a_8390_8053# a_9451_7682# a_9406_7695# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X624 vdd d4 a_13749_4519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X625 a_5424_2856# a_5431_2472# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X626 a_36302_3212# a_36298_3389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X627 a_26924_966# a_26926_867# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X628 vdd a_9679_3765# a_9471_3765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X629 a_39086_893# a_38873_893# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X630 a_14814_2024# a_15071_1834# a_13802_2205# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X631 a_17743_3302# a_17371_2882# a_16779_2648# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X632 a_23382_5243# a_23327_6271# a_23535_6271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X633 a_5402_6872# a_5891_6972# a_6099_6972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X634 gnd d2 a_3316_7464# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X635 a_6910_5812# a_6697_5812# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X636 a_40562_4914# a_41620_5135# a_41575_5148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X637 vdd d0 a_31181_1776# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X638 a_2831_4701# a_2975_2519# a_2930_2532# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X639 a_27412_651# a_27199_651# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X640 a_17591_1903# a_17378_1903# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X641 a_16564_5020# a_16351_5020# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X642 a_7079_5370# a_6965_5251# a_7173_5251# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X643 a_38270_3034# a_37849_3034# a_37573_3216# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X644 a_21625_5400# a_21623_5186# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X645 a_16080_4440# a_16078_4226# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X646 a_40565_3938# a_40818_3925# a_40515_3518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X647 vdd d0 a_20352_1813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X648 gnd a_4383_6722# a_4175_6722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X649 a_11479_7001# a_12283_6820# a_12442_7240# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X650 gnd a_30142_6853# a_29934_6853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X651 a_27392_4568# a_27179_4568# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X652 a_9414_5912# a_9671_5722# a_8402_6093# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X653 a_34043_5251# a_33622_5251# a_33944_5251# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X654 a_39245_1313# a_38873_893# a_38281_659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X655 a_33560_6791# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X656 a_6114_4036# a_5693_4036# a_5417_4218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X657 a_21628_3829# a_22114_3613# a_22322_3613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X658 a_37861_1074# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X659 a_36298_3389# a_36301_2797# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X660 a_41577_3757# a_41830_3744# a_40561_4115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X661 a_34986_4503# a_35106_6415# a_35057_6605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X662 a_5911_3055# a_5698_3055# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X663 a_32547_6557# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X664 a_1404_7793# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X665 a_19072_4943# a_20130_5164# a_20085_5177# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X666 a_40503_5652# a_40607_4901# a_40562_4914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X667 a_17646_1342# a_17433_1342# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X668 a_5705_2076# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X669 a_29905_3126# a_30162_2936# a_29850_3687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X670 a_20073_7137# a_20326_7124# a_19060_6903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X671 a_833_4057# a_412_4057# a_136_3957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X672 a_24619_4128# a_24876_3938# a_24573_3531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X673 a_24640_1010# a_24893_997# a_24581_1748# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X674 a_28628_2333# a_28415_2333# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X675 vdd d0 a_31175_3170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X676 a_38053_4576# a_37840_4576# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X677 vdd d2 a_30107_3497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X678 a_5402_7154# a_5402_6872# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X679 a_19037_1587# a_19132_1994# a_19087_2007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X680 a_10777_7882# a_11266_7982# a_11474_7982# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X681 a_25615_7687# a_25868_7674# a_24599_8045# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X682 a_38037_7932# a_37824_7932# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X683 a_20087_3786# a_20340_3773# a_19071_4144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X684 a_32294_3451# a_32775_3621# a_32983_3621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X685 a_1719_4308# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X686 a_21613_7360# a_22094_7530# a_22302_7530# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X687 vdd a_15059_3794# a_14851_3794# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X688 a_13811_1047# a_14869_1268# a_14820_1458# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X689 a_1781_7232# a_1409_6812# a_817_6578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X690 vdd d2 a_3316_7464# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X691 a_30892_7843# a_30902_7100# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X692 a_16771_4605# a_17576_4839# a_17735_5259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X693 a_9444_1252# a_9440_1429# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X694 a_12462_3323# a_12090_2903# a_11499_3084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X695 a_10811_2501# a_10809_2287# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X696 a_2930_2532# a_3128_3547# a_3083_3560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X697 a_16097_1499# a_16578_1669# a_16786_1669# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X698 a_41559_7285# a_41816_7095# a_40550_6874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X699 a_39289_2341# a_39076_2341# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X700 a_616_5599# a_403_5599# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X701 a_38042_6951# a_37829_6951# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X702 a_16547_7961# a_16334_7961# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X703 a_35264_7876# a_36322_8097# a_36273_8287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X704 vdd a_8684_1005# a_8476_1005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X705 vdd a_4383_6722# a_4175_6722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X706 a_28608_6250# a_28395_6250# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X707 a_1479_3315# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X708 a_37836_5972# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X709 a_22335_2068# a_21914_2068# a_21638_2250# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X710 vdd a_40798_7842# a_40590_7842# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X711 a_27588_6528# a_27167_6528# a_26901_6360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X712 a_41573_3934# a_41830_3744# a_40561_4115# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X713 a_40578_1174# a_41639_803# a_41590_993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X714 gnd d1 a_35522_6882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X715 a_34986_4503# a_35106_6415# a_35061_6428# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X716 a_22339_672# a_23144_906# a_23303_1326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X717 a_40362_2490# a_40615_2477# a_40263_4659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X718 a_2153_220# a_2044_220# a_2252_220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X719 gnd a_35529_5903# a_35321_5903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X720 a_32792_680# a_32579_680# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X721 gnd d1 a_3366_7884# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X722 a_20069_7314# a_20326_7124# a_19060_6903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X723 a_138_3858# a_143_3472# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X724 a_11085_2105# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X725 a_36272_7872# a_36282_7129# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X726 a_22949_7203# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X727 a_24549_7625# a_24653_6874# a_24604_7064# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X728 a_9440_1429# a_9443_837# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X729 a_20079_5743# a_20075_5920# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X730 a_27596_5964# a_27175_5964# a_26899_5864# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X731 a_39585_178# a_40312_4469# a_40263_4659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X732 a_2930_2532# a_3183_2519# a_2831_4701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X733 a_3091_1777# a_3348_1587# a_2926_2709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X734 a_29834_7427# a_29929_7834# a_29880_8024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X735 a_13795_3184# a_14052_2994# a_13740_3745# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X736 a_35292_2176# a_35549_1986# a_35246_1579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X737 a_1818_1474# a_1436_1916# a_844_1682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X738 a_25611_7864# a_25868_7674# a_24599_8045# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X739 a_36289_6150# a_36542_6137# a_35276_5916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X740 gnd a_15060_4209# a_14852_4209# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X741 a_20083_3963# a_20340_3773# a_19071_4144# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X742 a_7434_199# a_7325_199# a_5243_132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X743 a_12447_7359# a_12333_7240# a_12541_7240# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X744 a_28455_5222# a_28242_5222# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X745 a_16078_3944# a_16080_3845# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X746 gnd a_31175_3170# a_30967_3170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X747 a_1831_220# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X748 a_3150_1039# a_3403_1026# a_3091_1777# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X749 a_424_2097# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X750 a_17748_3421# a_17634_3302# a_17842_3302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X751 vdd d0 a_4403_2805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X752 gnd d1 a_19308_7871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X753 a_33768_7772# a_33555_7772# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X754 vdd a_4410_1826# a_4202_1826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X755 a_16754_7546# a_16333_7546# a_16060_7762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X756 a_148_2279# a_148_1997# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X757 vdd d0 a_25905_816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X758 a_1813_1355# a_1441_935# a_850_1116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X759 gnd a_3316_7464# a_3108_7464# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X760 a_24620_4927# a_24873_4914# a_24561_5665# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X761 a_38056_3600# a_37843_3600# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X762 vdd d0 a_31155_7087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X763 vdd a_41847_803# a_41639_803# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X764 vdd d2 a_14009_1595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X765 gnd a_9660_8097# a_9452_8097# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X766 a_22095_7945# a_21882_7945# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X767 a_14799_6179# a_15052_6166# a_13786_5945# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X768 a_38923_1313# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X769 a_829_4618# a_1634_4852# a_1793_5272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X770 a_16351_5020# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X771 a_5898_5993# a_5685_5993# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X772 a_5411_5794# a_5897_5578# a_6105_5578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X773 gnd d0 a_41828_5135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X774 a_5709_680# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X775 vdd a_20352_1813# a_20144_1813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X776 a_37567_5387# a_37565_5173# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X777 a_36281_6714# a_36277_6891# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X778 a_22322_3613# a_23127_3847# a_23296_3405# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X779 a_3118_6916# a_4176_7137# a_4131_7150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X780 a_33949_5370# a_33567_5812# a_32976_5993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X781 a_39332_3273# a_39289_2341# a_39473_4266# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X782 a_21611_7146# a_22100_6964# a_22308_6964# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X783 gnd d0 a_20333_6145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X784 a_16077_5416# a_16558_5586# a_16766_5586# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X785 a_17735_5259# a_17626_5259# a_17834_5259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X786 gnd d0 a_41842_1784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X787 a_35214_7456# a_35309_7863# a_35264_7876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X788 a_39230_5349# a_38848_5791# a_38256_5557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X789 a_16095_1285# a_16095_1003# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X790 a_17433_1342# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X791 a_23402_1326# a_23347_2354# a_23531_4279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X792 a_28651_7182# a_28230_7182# a_28552_7182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X793 a_5417_4218# a_5417_3936# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X794 gnd d1 a_14059_2015# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X795 a_41563_7108# a_41559_7285# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X796 a_28415_2333# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X797 a_22315_5985# a_21894_5985# a_21618_6167# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X798 a_10794_5223# a_10794_4941# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X799 a_3146_1216# a_3403_1026# a_3091_1777# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X800 vdd a_31175_3170# a_30967_3170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X801 vdd a_30107_3497# a_29899_3497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X802 a_4162_858# a_4158_1035# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X803 a_12573_1363# a_12518_2391# a_12702_4316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X804 a_29606_4474# a_29726_6386# a_29677_6576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X805 a_32989_3055# a_32568_3055# a_32292_3237# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X806 a_37824_7932# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X807 a_12459_5399# a_12077_5841# a_11486_6022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X808 a_23144_906# a_22931_906# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X809 a_17842_3302# a_17799_2370# a_17983_4295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X810 a_5431_2472# a_5910_2640# a_6118_2640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X811 a_18868_2696# a_19125_2506# a_18773_4688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X812 a_33952_3294# a_33580_2874# a_32989_3055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X813 a_26892_6843# a_27381_6943# a_27589_6943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X814 a_18777_4511# a_18897_6423# a_18848_6613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X815 vdd a_3316_7464# a_3108_7464# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X816 a_14804_5198# a_14800_5375# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X817 a_23182_3286# a_22969_3286# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X818 a_33964_1334# a_33592_914# a_33000_680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X819 a_14795_6356# a_15052_6166# a_13786_5945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X820 a_39324_5230# a_39269_6258# a_39477_6258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X821 a_24628_2970# a_25686_3191# a_25637_3381# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X822 a_33592_914# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X823 a_3141_2197# a_3398_2007# a_3095_1600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X824 a_35272_6093# a_35529_5903# a_35226_5496# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X825 a_1806_3434# a_1424_3876# a_833_4057# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X826 a_40577_1978# a_41635_2199# a_41590_2212# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X827 gnd a_15040_8126# a_14832_8126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X828 a_28569_5341# a_28455_5222# a_28663_5222# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X829 a_39076_2341# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X830 a_20063_7880# a_20320_7690# a_19051_8061# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X831 a_41559_7285# a_41562_6693# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X832 a_403_5599# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X833 a_8407_5112# a_9468_4741# a_9419_4931# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X834 a_32773_5012# a_32560_5012# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X835 vdd d0 a_41828_5135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X836 a_28405_4802# a_28192_4802# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X837 a_12814_228# a_12705_228# a_12913_228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X838 a_16334_7961# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X839 a_28395_6250# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X840 gnd d1 a_8664_4922# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X841 a_27407_1632# a_27194_1632# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X842 a_27604_4007# a_27183_4007# a_26907_4189# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X843 vdd d3 a_29954_2469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X844 gnd a_35522_6882# a_35314_6882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X845 a_6110_4597# a_5689_4597# a_5416_4813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X846 vdd d0 a_20333_6145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X847 vdd d0 a_41842_1784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X848 a_12573_1363# a_12152_1363# a_12474_1363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X849 a_25632_4362# a_25635_3770# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X850 a_22894_7764# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X851 a_39104_7190# a_38891_7190# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X852 a_32969_6972# a_33773_6791# a_33932_7211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X853 a_17748_3421# a_17366_3863# a_16775_4044# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X854 a_13782_6122# a_14039_5932# a_13736_5525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X855 a_14800_5375# a_14803_4783# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X856 a_19087_2007# a_20145_2228# a_20100_2241# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X857 gnd a_3366_7884# a_3158_7884# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X858 gnd a_41811_8076# a_40545_7855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X859 a_849_701# a_428_701# a_162_716# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X860 a_21919_1087# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X861 a_13802_2205# a_14863_1834# a_14818_1847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X862 vdd d1 a_14059_2015# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X863 a_11077_2669# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X864 a_9428_3389# a_9685_3199# a_8419_2978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X865 a_428_701# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X866 a_35285_3155# a_35542_2965# a_35230_3716# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X867 a_11283_5041# a_11070_5041# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X868 a_1793_5272# a_1684_5272# a_1892_5272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X869 a_30916_3749# a_31169_3736# a_29900_4107# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X870 a_16090_2266# a_16579_2084# a_16787_2084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X871 a_29606_4474# a_29726_6386# a_29681_6399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X872 a_16559_6001# a_16346_6001# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X873 a_10814_1024# a_11303_1124# a_11511_1124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X874 a_6126_2076# a_6930_1895# a_7099_1453# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X875 a_27387_5549# a_27174_5549# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X876 gnd a_19308_7871# a_19100_7871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X877 vdd a_4403_2805# a_4195_2805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X878 a_31994_96# a_37072_111# a_37394_111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X879 a_18777_4511# a_18897_6423# a_18852_6436# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X880 a_40507_5475# a_40602_5882# a_40557_5895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X881 a_37072_111# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X882 a_37856_2055# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X883 a_33555_7772# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X884 a_20068_8118# a_20321_8105# a_19055_7884# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X885 a_32267_7853# a_32756_7953# a_32964_7953# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X886 a_5677_6557# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X887 a_12553_5280# a_12132_5280# a_12459_5399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X888 a_5906_4036# a_5693_4036# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X889 a_24420_2503# a_24618_3518# a_24573_3531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X890 a_12706_6308# a_12593_4316# a_12801_4316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X891 vdd a_15040_8126# a_14832_8126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X892 gnd d0 a_4384_7137# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X893 a_33870_4287# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X894 a_19071_4144# a_19328_3954# a_19025_3547# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X895 a_23347_2354# a_23134_2354# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X896 vdd a_31155_7087# a_30947_7087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X897 a_8407_5112# a_9468_4741# a_9423_4754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X898 gnd d1 a_3386_3967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X899 a_5891_6972# a_5678_6972# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X900 a_3075_5517# a_3170_5924# a_3125_5937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X901 a_22327_2632# a_21906_2632# a_21640_2464# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X902 a_40566_3134# a_41627_2763# a_41578_2953# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X903 a_4126_8131# a_4122_8308# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X904 a_16572_3063# a_16359_3063# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X905 a_15904_140# a_17773_207# a_18082_4295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X906 a_12706_6308# a_12285_6308# a_12553_5280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X907 gnd d1 a_40823_2944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X908 a_5685_5993# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X909 gnd a_41828_5135# a_41620_5135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X910 a_813_7974# a_392_7974# a_116_7874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X911 a_33932_7211# a_33560_6791# a_32969_6972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X912 gnd a_40830_1965# a_40622_1965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X913 a_12467_3442# a_12353_3323# a_12561_3323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X914 a_32983_3621# a_32562_3621# a_32289_3837# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X915 a_26832_103# a_26411_103# a_23742_191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X916 a_20674_n19# d8 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X917 a_5436_896# a_5443_695# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X918 a_8395_7072# a_8652_6882# a_8340_7633# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X919 a_26411_103# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X920 a_41554_8266# a_41811_8076# a_40545_7855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X921 a_39213_7190# a_38841_6770# a_38249_6536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X922 gnd a_20333_6145# a_20125_6145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X923 a_2835_4524# a_3088_4511# a_2153_220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X924 a_36314_1252# a_36310_1429# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X925 gnd a_41842_1784# a_41634_1784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X926 a_1786_7351# a_1404_7793# a_813_7974# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X927 gnd d0 a_20325_6709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X928 a_6131_1095# a_5710_1095# a_5434_995# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X929 a_19017_5504# a_19112_5911# a_19067_5924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X930 a_36277_8110# a_37548_8114# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X931 a_11479_7001# a_11058_7001# a_10782_7183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X932 a_38249_6536# a_37828_6536# a_37562_6368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X933 a_30912_3926# a_31169_3736# a_29900_4107# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X934 a_19076_3163# a_20137_2792# a_20088_2982# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X935 a_7067_7330# a_6685_7772# a_6093_7538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X936 a_38057_4015# a_37844_4015# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X937 a_16097_904# a_16104_703# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X938 a_4122_8308# a_4125_7716# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X939 a_16058_7861# a_16060_7762# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X940 a_33000_680# a_33805_914# a_33964_1334# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X941 vdd a_24888_1978# a_24680_1978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X942 a_22307_6549# a_21886_6549# a_21613_6765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X943 a_16792_1103# a_16371_1103# a_16095_1285# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X944 a_41578_2953# a_41590_2212# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X945 a_10784_7397# a_10782_7183# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X946 gnd d0 a_25873_6693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X947 vdd d0 a_41822_5701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X948 a_30916_3749# a_30912_3926# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X949 a_21898_4589# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X950 vdd a_8664_4922# a_8456_4922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X951 gnd d4 a_13749_4519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X952 a_36310_1429# a_36313_837# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X953 a_38262_4991# a_39066_4810# a_39225_5230# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X954 a_25631_3947# a_25641_3204# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X955 a_1900_3315# a_1479_3315# a_1801_3315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X956 a_21618_6167# a_21618_5885# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X957 a_16070_6183# a_16559_6001# a_16767_6001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X958 a_30933_808# a_31186_795# a_29917_1166# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X959 a_37582_1856# a_38068_1640# a_38276_1640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X960 a_5243_132# a_7112_199# a_7434_199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X961 a_40566_3134# a_41627_2763# a_41582_2776# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X962 a_7112_199# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X963 a_6106_5993# a_6910_5812# a_7079_5370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X964 gnd d2 a_8609_5483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X965 a_26901_5765# a_27387_5549# a_27595_5549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X966 vdd d0 a_9685_3199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X967 a_27400_2611# a_27187_2611# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X968 a_32560_5012# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X969 vdd a_41828_5135# a_41620_5135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X970 a_28192_4802# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X971 a_9431_2797# a_9427_2974# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X972 a_2831_4701# a_2975_2519# a_2926_2709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X973 gnd a_30087_7414# a_29879_7414# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X974 a_21628_4424# a_22111_4589# a_22319_4589# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X975 a_13740_3745# a_13844_2994# a_13799_3007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X976 a_27194_1632# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X977 a_30929_2204# a_30925_2381# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X978 vdd a_29954_2469# a_29746_2469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X979 a_24608_6887# a_25666_7108# a_25621_7121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X980 a_26901_6360# a_26899_6146# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X981 a_3134_3176# a_4195_2805# a_4150_2818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X982 a_41590_993# a_37594_674# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X983 gnd d0 a_25901_2212# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X984 a_13775_7101# a_14032_6911# a_13720_7662# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X985 a_32281_6389# a_32279_6175# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X986 vdd a_20333_6145# a_20125_6145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X987 a_2831_4701# a_3088_4511# a_2153_220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X988 vdd a_41842_1784# a_41634_1784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X989 a_16075_5202# a_16075_4920# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X990 vdd d1 a_35549_1986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X991 vdd d0 a_31150_8068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X992 a_14787_6920# a_14799_6179# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X993 a_35281_4935# a_36339_5156# a_36290_5346# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X994 a_5422_3237# a_5911_3055# a_6119_3055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X995 a_11070_5041# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X996 a_24619_4128# a_25680_3757# a_25635_3770# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X997 a_37567_5387# a_38048_5557# a_38256_5557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X998 a_38073_659# a_37860_659# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X999 a_10504_125# a_10395_125# a_10603_125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1000 a_24321_4672# a_24465_2490# a_24416_2680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1001 a_30897_8081# a_30893_8258# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1002 a_27380_6528# a_27167_6528# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1003 a_13786_5945# a_14844_6166# a_14795_6356# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1004 a_35292_2176# a_36353_1805# a_36304_1995# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1005 a_34031_7211# a_33610_7211# a_33937_7330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1006 a_27174_5549# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1007 a_5243_132# a_5134_132# a_5342_132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1008 a_32755_7538# a_32542_7538# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1009 a_39312_7190# a_38891_7190# a_39213_7190# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1010 a_6111_5012# a_5690_5012# a_5414_4912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1011 a_21631_3229# a_21631_2947# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1012 a_7325_199# a_7112_199# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1013 a_34063_1334# a_34008_2362# a_34192_4287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1014 gnd d1 a_30154_4893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1015 a_5693_4036# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1016 a_16345_5586# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1017 a_9419_4931# a_9427_4193# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1018 a_9427_4193# a_9680_4180# a_8414_3959# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1019 a_624_3642# a_411_3642# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1020 vdd d2 a_8609_5483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1021 a_23134_2354# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1022 a_36284_5912# a_36294_5169# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1023 vdd a_30087_7414# a_29879_7414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1024 a_2930_2532# a_3128_3547# a_3079_3737# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1025 a_20099_1826# a_20352_1813# a_19083_2184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1026 a_8207_2688# a_8464_2498# a_8112_4680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1027 a_26914_3422# a_26912_3208# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1028 a_32294_3451# a_32292_3237# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1029 gnd a_40823_2944# a_40615_2944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1030 gnd d2 a_35467_7443# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1031 vdd d0 a_25901_2212# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1032 a_11265_7567# a_11052_7567# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1033 a_4134_6348# a_4391_6158# a_3125_5937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1034 a_10823_724# a_11302_709# a_11510_709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1035 a_7434_199# a_8161_4490# a_8116_4503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1036 a_417_3076# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1037 a_21643_1269# a_22132_1087# a_22340_1087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1038 a_35281_4935# a_36339_5156# a_36294_5169# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1039 a_39230_5349# a_39116_5230# a_39324_5230# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1040 a_17983_4295# a_17586_2370# a_17854_1342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1041 a_24400_6420# a_24598_7435# a_24549_7625# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1042 gnd a_20325_6709# a_20117_6709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1043 a_18773_4688# a_18917_2506# a_18872_2519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1044 a_28400_5783# a_28187_5783# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1045 a_16097_904# a_16583_688# a_16791_688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1046 a_604_7559# a_391_7559# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1047 a_23283_5243# a_23174_5243# a_23382_5243# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1048 a_1429_2895# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1049 gnd d1 a_8659_5903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1050 vdd d0 a_4396_5177# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1051 a_23124_4823# a_22911_4823# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1052 gnd a_24861_6874# a_24653_6874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1053 a_13786_5945# a_14844_6166# a_14799_6179# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1054 a_28242_5222# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1055 a_27616_2047# a_28420_1866# a_28589_1424# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1056 a_22126_1653# a_21913_1653# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1057 gnd a_9691_1805# a_9483_1805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1058 gnd d2 a_13977_7472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1059 a_36296_3778# a_36549_3765# a_35280_4136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1060 gnd a_25873_6693# a_25665_6693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1061 vdd d1 a_8684_1005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1062 vdd a_41822_5701# a_41614_5701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1063 a_11485_5607# a_11064_5607# a_10796_5437# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1064 vdd d1 a_35529_5903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1065 a_21914_2068# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1066 a_19056_7080# a_20117_6709# a_20072_6722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1067 a_26899_5864# a_26901_5765# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1068 a_5902_4597# a_5689_4597# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1069 a_37565_5173# a_37565_4891# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1070 a_9423_4370# a_9680_4180# a_8414_3959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1071 a_32279_5893# a_32281_5794# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1072 a_40362_2490# a_40560_3505# a_40515_3518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1073 a_5436_1491# a_5434_1277# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1074 a_4150_2818# a_4146_2995# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1075 a_24565_5488# a_24660_5895# a_24615_5908# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1076 a_17773_207# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1077 a_1892_5272# a_1837_6300# a_2045_6300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1078 a_16065_6781# a_16551_6565# a_16759_6565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1079 a_824_5599# a_403_5599# a_130_5815# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1080 a_35272_6093# a_36333_5722# a_36284_5912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1081 a_5419_3837# a_5905_3621# a_6113_3621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1082 a_38276_1640# a_39081_1874# a_39250_1432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1083 a_14806_3807# a_15059_3794# a_13790_4165# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1084 a_34196_6279# a_34083_4287# a_34291_4287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1085 vdd d2 a_35467_7443# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1086 a_1892_5272# a_1471_5272# a_1798_5391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1087 a_38269_2619# a_37848_2619# a_37582_2451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1088 a_28413_2845# a_28200_2845# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1089 a_41575_5148# a_41571_5325# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1090 a_28475_1305# a_28262_1305# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1091 vdd d1 a_14039_5932# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1092 a_40550_6874# a_41608_7095# a_41559_7285# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1093 a_5416_4813# a_5419_4432# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1094 gnd d1 a_30157_3917# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1095 a_28207_1866# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1096 vdd a_4379_8118# a_4171_8118# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1097 a_23209_4279# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1098 a_34196_6279# a_33775_6279# a_34043_5251# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1099 a_33788_3855# a_33575_3855# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1100 a_23303_1326# a_22931_906# a_22339_672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1101 gnd d0 a_25893_2776# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1102 a_24400_6420# a_24598_7435# a_24553_7448# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1103 a_27621_1066# a_27200_1066# a_26924_966# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1104 a_8431_1018# a_8684_1005# a_8372_1756# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1105 a_5404_7368# a_5402_7154# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1106 a_23271_7203# a_22899_6783# a_22307_6549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1107 a_26901_5765# a_26906_5379# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1108 a_16774_3629# a_16353_3629# a_16085_3459# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1109 gnd d0 a_31169_3736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1110 gnd a_25900_1797# a_25692_1797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1111 a_35230_3716# a_35334_2965# a_35285_3155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1112 a_2045_6300# a_1624_6300# a_1892_5272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1113 a_153_1298# a_642_1116# a_850_1116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1114 a_33957_3413# a_33843_3294# a_34051_3294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1115 a_9406_7695# a_9659_7682# a_8390_8053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1116 a_32964_7953# a_32543_7953# a_32267_8135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1117 a_28557_7301# a_28175_7743# a_27583_7509# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1118 gnd a_24653_6407# a_24445_6407# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1119 a_3118_6916# a_4176_7137# a_4127_7327# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1120 gnd d0 a_9680_4180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1121 a_22115_4028# a_21902_4028# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1122 vdd d2 a_13977_7472# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1123 gnd d0 a_9665_7116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1124 a_3083_3560# a_3178_3967# a_3129_4157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1125 a_36292_3955# a_36549_3765# a_35280_4136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1126 a_5404_7368# a_5885_7538# a_6093_7538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1127 gnd d2 a_3328_5504# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1128 a_41571_5325# a_41574_4733# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1129 a_26912_2926# a_26914_2827# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1130 a_3129_4157# a_4190_3786# a_4141_3976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1131 a_12298_3884# a_12085_3884# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1132 a_21623_5186# a_22112_5004# a_22320_5004# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1133 vdd d1 a_8667_3946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1134 a_32292_2955# a_32294_2856# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1135 a_41575_5148# a_41828_5135# a_40562_4914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1136 a_20080_4939# a_20088_4201# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1137 a_38282_1074# a_37861_1074# a_37585_1256# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1138 a_14803_4399# a_15060_4209# a_13794_3988# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1139 a_118_7775# a_604_7559# a_812_7559# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1140 a_24325_4495# a_24445_6407# a_24400_6420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1141 gnd a_30154_4893# a_29946_4893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1142 a_22320_5004# a_23124_4823# a_23283_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1143 a_5922_680# a_5709_680# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1144 a_39218_7309# a_38836_7751# a_38245_7932# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1145 a_411_3642# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1146 a_4158_2254# a_4411_2241# a_3145_2020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1147 a_35272_6093# a_36333_5722# a_36288_5735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1148 a_41589_1797# a_41842_1784# a_40573_2155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1149 a_21640_1869# a_22126_1653# a_22334_1653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1150 a_6126_2076# a_5705_2076# a_5429_2258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1151 gnd a_9671_5722# a_9463_5722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1152 a_5923_1095# a_5710_1095# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1153 a_39572_4266# a_39151_4266# a_39473_4266# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1154 a_6130_680# a_6935_914# a_7094_1334# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1155 vdd a_36561_1805# a_36353_1805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1156 a_6898_7772# a_6685_7772# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1157 a_20085_5177# a_20338_5164# a_19072_4943# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1158 vdd d0 a_20341_4188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1159 gnd a_35467_7443# a_35259_7443# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1160 a_21894_5985# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1161 a_32284_4912# a_32773_5012# a_32981_5012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1162 a_33964_1334# a_33592_914# a_33001_1095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1163 a_24631_2168# a_24888_1978# a_24585_1571# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1164 a_845_2097# a_424_2097# a_148_1997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1165 a_11052_7567# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1166 a_8340_7633# a_8444_6882# a_8395_7072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1167 a_12479_1482# a_12097_1924# a_11505_1690# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1168 a_32294_2856# a_32301_2472# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1169 vdd d0 a_25893_2776# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1170 a_9403_8287# a_9660_8097# a_8394_7876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1171 vdd d0 a_31169_3736# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1172 a_32980_4597# a_33785_4831# a_33944_5251# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1173 a_13811_1047# a_14064_1034# a_13752_1785# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1174 gnd d3 a_29954_2469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1175 a_26912_3208# a_27401_3026# a_27609_3026# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1176 a_12801_4316# a_12380_4316# a_12706_6308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1177 a_9402_7872# a_9659_7682# a_8390_8053# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1178 a_10789_5922# a_11278_6022# a_11486_6022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1179 a_38049_5972# a_37836_5972# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1180 a_32306_1491# a_32787_1661# a_32995_1661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1181 vdd d0 a_15064_2813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1182 a_38256_5557# a_39061_5791# a_39230_5349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1183 vdd d0 a_9680_4180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1184 a_13807_1224# a_14868_853# a_14823_866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1185 a_14786_7724# a_15039_7711# a_13770_8082# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1186 a_391_7559# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1187 vdd d0 a_9665_7116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1188 a_16346_6001# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1189 a_18082_4295# a_17661_4295# a_17983_4295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1190 gnd a_9684_2784# a_9476_2784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1191 vdd a_15071_1834# a_14863_1834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1192 a_19087_2007# a_20145_2228# a_20096_2418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1193 a_21625_5400# a_22106_5570# a_22314_5570# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1194 vdd a_4396_5177# a_4188_5177# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1195 a_1793_5272# a_1421_4852# a_829_4618# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1196 a_20104_845# a_20100_1022# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1197 a_36313_837# a_36309_1014# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1198 a_36301_2797# a_36297_2974# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1199 a_25620_6706# a_25616_6883# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1200 a_27395_3592# a_27182_3592# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1201 a_12474_1363# a_12102_943# a_11511_1124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1202 gnd a_13977_7472# a_13769_7472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1203 a_28187_5783# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1204 a_3129_4157# a_4190_3786# a_4145_3799# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1205 a_41571_5325# a_41828_5135# a_40562_4914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1206 a_17760_1461# a_17378_1903# a_16787_2084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1207 a_17822_7219# a_17401_7219# a_17723_7219# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1208 a_8411_4935# a_8664_4922# a_8352_5673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1209 a_12561_3323# a_12140_3323# a_12467_3442# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1210 a_21640_2464# a_21638_2250# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1211 a_37573_2934# a_38062_3034# a_38270_3034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1212 vdd d1 a_40803_6861# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1213 gnd d2 a_35487_3526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1214 gnd d0 a_36555_3199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1215 a_22302_7530# a_21881_7530# a_21613_7360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1216 vdd d4 a_40520_4469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1217 a_35297_1195# a_35554_1005# a_35242_1756# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1218 a_40541_8032# a_41602_7661# a_41553_7851# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1219 a_4154_2431# a_4411_2241# a_3145_2020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1220 a_13720_7662# a_13824_6911# a_13779_6924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1221 a_30902_7100# a_30898_7277# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1222 vdd a_40810_5882# a_40602_5882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1223 a_41585_1974# a_41842_1784# a_40573_2155# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1224 a_20092_2805# a_20088_2982# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1225 vdd a_9671_5722# a_9463_5722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1226 a_38269_2619# a_39074_2853# a_39233_3273# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1227 a_39250_1432# a_39136_1313# a_39344_1313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1228 a_16078_3944# a_16567_4044# a_16775_4044# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1229 a_24420_2503# a_24618_3518# a_24569_3708# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1230 a_11303_1124# a_11090_1124# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1231 a_27188_3026# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1232 a_1818_1474# a_1704_1355# a_1912_1355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1233 a_12278_7801# a_12065_7801# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1234 vdd d2 a_19270_5491# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1235 a_20081_5354# a_20338_5164# a_19072_4943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1236 a_6113_3621# a_6918_3855# a_7087_3413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1237 vdd a_35467_7443# a_35259_7443# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1238 a_5402_7154# a_5891_6972# a_6099_6972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1239 a_6131_1095# a_6935_914# a_7094_1334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1240 gnd d1 a_8679_1986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1241 a_28200_2845# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1242 a_25624_6319# a_25881_6129# a_24615_5908# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1243 a_28262_1305# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1244 a_4134_6348# a_4137_5756# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1245 a_5419_4432# a_5417_4218# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1246 a_38262_4991# a_37841_4991# a_37565_5173# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1247 gnd a_30157_3917# a_29949_3917# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1248 a_641_701# a_428_701# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1249 vout a_20674_n19# a_20996_n19# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1250 a_29866_1550# a_29961_1957# a_29916_1970# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1251 gnd d2 a_13997_3555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1252 a_17591_1903# a_17378_1903# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1253 a_7193_1334# a_7138_2362# a_7322_4287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1254 a_19051_8061# a_20112_7690# a_20063_7880# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1255 a_13807_1224# a_14064_1034# a_13752_1785# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1256 a_642_1116# a_429_1116# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1257 a_7213_4287# a_7000_4287# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1258 a_33575_3855# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1259 a_5342_132# a_4921_132# a_2252_220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1260 gnd a_25893_2776# a_25685_2776# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1261 a_36289_4931# a_36297_4193# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1262 a_32287_4218# a_32776_4036# a_32984_4036# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1263 a_14782_7901# a_15039_7711# a_13770_8082# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1264 a_6106_5993# a_5685_5993# a_5409_6175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1265 gnd a_20340_3773# a_20132_3773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1266 a_17760_1461# a_17646_1342# a_17854_1342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1267 a_6930_1895# a_6717_1895# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1268 a_30898_7277# a_30901_6685# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1269 a_5903_5012# a_5690_5012# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1270 vdd a_9684_2784# a_9476_2784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1271 vdd d4 a_19030_4498# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1272 a_36282_7129# a_36278_7306# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1273 a_29897_5083# a_30154_4893# a_29842_5644# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1274 a_10777_8164# a_10777_7882# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1275 vdd a_13977_7472# a_13769_7472# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1276 a_818_6993# a_1622_6812# a_1781_7232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1277 gnd d0 a_4410_1826# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1278 a_29917_1166# a_30978_795# a_30933_808# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1279 a_825_6014# a_404_6014# a_128_5914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1280 a_39066_4810# a_38853_4810# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1281 a_11498_2669# a_12303_2903# a_12462_3323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1282 gnd a_3328_5504# a_3120_5504# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1283 a_21906_2632# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1284 a_38068_1640# a_37855_1640# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1285 vdd d0 a_31167_5127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1286 a_12085_3884# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1287 a_10395_125# a_10182_125# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1288 a_40570_2957# a_40823_2944# a_40511_3695# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1289 a_20088_4201# a_20084_4378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1290 vdd d2 a_35487_3526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1291 a_9427_2974# a_9439_2233# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1292 a_40541_8032# a_41602_7661# a_41557_7674# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1293 a_17571_5820# a_17358_5820# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1294 a_20079_5743# a_20332_5730# a_19063_6101# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1295 a_19088_1203# a_20149_832# a_20100_1022# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1296 vdd a_4399_4201# a_4191_4201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1297 a_28443_7182# a_28230_7182# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1298 a_36278_7306# a_36281_6714# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1299 a_4150_2818# a_4403_2805# a_3134_3176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1300 vdd d2 a_40768_3505# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1301 a_5710_1095# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1302 a_3109_8074# a_4170_7703# a_4125_7716# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1303 a_397_6993# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1304 a_3130_4956# a_4188_5177# a_4143_5190# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1305 vdd d1 a_24868_5895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1306 a_37828_6536# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1307 a_12705_228# a_12492_228# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1308 a_24624_3147# a_24881_2957# a_24569_3708# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1309 a_6685_7772# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1310 a_150_2493# a_629_2661# a_837_2661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1311 a_12462_3323# a_12090_2903# a_11498_2669# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1312 gnd d0 a_36535_7116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1313 vdd d2 a_13997_3555# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1314 a_148_1997# a_150_1898# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1315 a_1409_6812# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1316 a_21886_6549# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1317 a_133_5215# a_133_4933# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1318 vdd a_25893_2776# a_25685_2776# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1319 a_25620_6706# a_25873_6693# a_24604_7064# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1320 a_38042_6951# a_37829_6951# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1321 gnd d1 a_35537_3946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1322 a_28911_4258# a_28815_170# a_26733_103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1323 a_41565_5891# a_41822_5701# a_40553_6072# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1324 vdd a_20340_3773# a_20132_3773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1325 vdd a_30119_1537# a_29911_1537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1326 gnd a_29954_2469# a_29746_2469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1327 a_37836_5972# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1328 a_39233_3273# a_39124_3273# a_39332_3273# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1329 gnd d0 a_36549_3765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1330 vdd a_15064_2813# a_14856_2813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1331 a_24573_3531# a_24668_3938# a_24619_4128# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1332 a_39136_1313# a_38923_1313# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1333 gnd d0 a_31150_8068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1334 a_26894_7339# a_27375_7509# a_27583_7509# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1335 a_16338_6565# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1336 vdd a_25888_3757# a_25680_3757# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1337 a_23194_1326# a_22981_1326# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1338 gnd d0 a_15045_7145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1339 a_32272_6872# a_32274_6773# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1340 a_24619_4128# a_25680_3757# a_25631_3947# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1341 a_27182_3592# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1342 a_17743_3302# a_17371_2882# a_16780_3063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1343 gnd d1 a_14047_3975# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1344 a_41586_2389# a_41589_1797# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1345 a_12442_7240# a_12070_6820# a_11479_7001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1346 a_20075_5920# a_20332_5730# a_19063_6101# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1347 a_7138_2362# a_6925_2362# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1348 vdd a_40803_6861# a_40595_6861# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1349 a_5417_3936# a_5419_3837# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1350 a_11493_3650# a_11072_3650# a_10799_3866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1351 a_148_2279# a_637_2097# a_845_2097# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1352 gnd a_36555_3199# a_36347_3199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1353 vdd a_9664_6701# a_9456_6701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1354 gnd d0 a_15059_3794# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1355 a_23144_906# a_22931_906# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1356 a_6118_2640# a_5697_2640# a_5431_2472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1357 a_25648_2225# a_25901_2212# a_24635_1991# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1358 a_23276_7322# a_22894_7764# a_22303_7945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1359 a_33988_6279# a_33775_6279# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1360 a_27616_2047# a_27195_2047# a_26919_2229# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1361 gnd d0 a_9660_8097# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1362 gnd d1 a_3371_6903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1363 a_11090_1124# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1364 a_32287_4218# a_32287_3936# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1365 a_39116_5230# a_38903_5230# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1366 a_27601_4983# a_27180_4983# a_26904_4883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1367 a_23630_4279# a_23209_4279# a_23531_4279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1368 a_26894_6744# a_26901_6360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1369 a_12065_7801# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1370 vdd d0 a_36535_7116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1371 a_32274_6773# a_32281_6389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1372 a_29830_7604# a_29934_6853# a_29885_7043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1373 a_9440_1429# a_9697_1239# a_8431_1018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1374 a_28557_7301# a_28443_7182# a_28651_7182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1375 a_35289_2978# a_36347_3199# a_36302_3212# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1376 gnd a_13997_3555# a_13789_3555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1377 a_22095_7945# a_21882_7945# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1378 a_41562_6693# a_41558_6870# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1379 vdd d0 a_41831_4159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1380 a_10816_1520# a_11297_1690# a_11505_1690# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1381 gnd d1 a_19313_6890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1382 a_4138_6171# a_4391_6158# a_3125_5937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1383 vdd d0 a_36549_3765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1384 a_6098_6557# a_5677_6557# a_5404_6773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1385 gnd d0 a_31187_1210# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1386 gnd d3 a_35334_2498# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1387 a_38891_7190# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1388 a_22314_5570# a_23119_5804# a_23288_5362# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1389 a_5690_5012# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1390 a_13794_3988# a_14852_4209# a_14807_4222# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1391 a_23390_3286# a_22969_3286# a_23291_3286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1392 vdd d0 a_15045_7145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1393 a_5689_4597# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1394 a_5434_1277# a_5434_995# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1395 a_5918_2076# a_5705_2076# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1396 a_38061_2619# a_37848_2619# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1397 a_25635_3770# a_25631_3947# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1398 a_4146_2995# a_4158_2254# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1399 a_34291_4287# a_34195_199# a_34403_199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1400 a_817_6578# a_396_6578# a_130_6410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1401 gnd d0 a_4396_5177# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1402 gnd a_8597_7443# a_8389_7443# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1403 a_22100_6964# a_21887_6964# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1404 a_21620_6381# a_21618_6167# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1405 a_14803_4783# a_14799_4960# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1406 a_26832_103# a_31885_96# a_20996_n19# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1407 vdd a_20320_7690# a_20112_7690# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1408 vdd a_31167_5127# a_30959_5127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1409 a_3150_1039# a_4208_1260# a_4159_1450# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1410 gnd d1 a_3398_2007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1411 a_22919_2866# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1412 a_27376_7924# a_27163_7924# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1413 a_21631_2947# a_22120_3047# a_22328_3047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1414 gnd d1 a_40835_984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1415 a_25644_2402# a_25901_2212# a_24635_1991# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1416 vdd d1 a_30137_7834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1417 a_5419_4432# a_5902_4597# a_6110_4597# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1418 a_33944_5251# a_33572_4831# a_32981_5012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1419 a_32313_695# a_32792_680# a_33000_680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1420 a_13752_1785# a_13856_1034# a_13807_1224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1421 a_23308_1445# a_23194_1326# a_23402_1326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1422 a_28230_7182# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1423 a_32995_1661# a_32574_1661# a_32301_1877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1424 a_27603_3592# a_28408_3826# a_28577_3384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1425 a_26892_7125# a_27381_6943# a_27589_6943# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1426 a_35210_7633# a_35314_6882# a_35269_6895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1427 vdd a_24868_5895# a_24660_5895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1428 a_11510_709# a_11089_709# a_10816_925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1429 a_30925_2381# a_31182_2191# a_29916_1970# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1430 a_1798_5391# a_1416_5833# a_825_6014# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1431 a_17874_4295# a_17661_4295# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1432 a_37844_4015# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1433 a_40495_7435# a_40590_7842# a_40545_7855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1434 a_12541_7240# a_12120_7240# a_12447_7359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1435 a_22320_5004# a_21899_5004# a_21623_5186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1436 a_135_4834# a_621_4618# a_829_4618# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1437 vdd a_13997_3555# a_13789_3555# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1438 a_3063_7477# a_3158_7884# a_3113_7897# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1439 gnd a_36535_7116# a_36327_7116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1440 a_4921_132# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1441 a_5397_8135# a_5397_7853# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1442 gnd d0 a_15039_7711# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1443 a_13724_7485# a_13977_7472# a_13571_6457# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1444 a_16791_688# a_16370_688# a_16104_703# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1445 a_41585_1974# a_41595_1231# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1446 a_38069_2055# a_37856_2055# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1447 gnd a_35537_3946# a_35329_3946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1448 a_16370_688# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1449 a_35081_2511# a_35279_3526# a_35230_3716# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1450 vdd d0 a_31187_1210# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1451 a_8376_1579# a_8471_1986# a_8426_1999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1452 gnd a_4379_8118# a_4171_8118# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1453 a_34403_199# a_33982_199# a_34291_4287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1454 a_33964_1334# a_33855_1334# a_34063_1334# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1455 a_39081_1874# a_38868_1874# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1456 a_28425_885# a_28212_885# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1457 gnd a_20321_8105# a_20113_8105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1458 a_11069_4626# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1459 a_11298_2105# a_11085_2105# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1460 a_35277_5112# a_35534_4922# a_35222_5673# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1461 a_40582_997# a_41640_1218# a_41595_1231# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1462 a_37394_111# a_39263_178# a_39585_178# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1463 vdd a_8597_7443# a_8389_7443# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1464 gnd a_15045_7145# a_14837_7145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1465 a_9407_6891# a_9419_6150# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1466 a_39263_178# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1467 a_1912_1355# a_1491_1355# a_1813_1355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1468 gnd d0 a_25905_816# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1469 a_7094_1334# a_6722_914# a_6130_680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1470 a_3150_1039# a_4208_1260# a_4163_1273# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1471 a_7173_5251# a_7118_6279# a_7326_6279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1472 gnd a_14047_3975# a_13839_3975# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1473 a_20095_2003# a_20105_1260# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1474 a_3121_6114# a_3378_5924# a_3075_5517# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1475 vdd d0 a_9697_1239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1476 gnd d3 a_35314_6415# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1477 a_23370_7203# a_22949_7203# a_23271_7203# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1478 a_408_4618# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1479 vdd d0 a_20357_832# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1480 a_20100_1022# a_20357_832# a_19088_1203# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1481 a_13752_1785# a_13856_1034# a_13811_1047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1482 a_813_7974# a_1617_7793# a_1786_7351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1483 a_33775_6279# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1484 a_5898_5993# a_5685_5993# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1485 a_32984_4036# a_32563_4036# a_32287_3936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1486 a_24620_4927# a_25678_5148# a_25633_5161# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1487 a_19092_1026# a_20150_1247# a_20105_1260# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1488 a_17854_1342# a_17433_1342# a_17755_1342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1489 a_13787_5141# a_14044_4951# a_13732_5702# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1490 a_16583_688# a_16370_688# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1491 a_32267_8135# a_32756_7953# a_32964_7953# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1492 gnd a_8647_7863# a_8439_7863# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1493 a_6910_5812# a_6697_5812# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1494 a_26733_103# a_28602_170# a_28911_4258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1495 a_5434_1277# a_5923_1095# a_6131_1095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1496 a_13720_7662# a_13977_7472# a_13571_6457# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1497 a_22899_6783# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1498 vdd a_36535_7116# a_36327_7116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1499 a_16358_2648# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1500 vdd d0 a_15039_7711# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1501 a_8191_6428# a_8389_7443# a_8340_7633# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1502 a_40558_5091# a_41619_4720# a_41570_4910# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1503 a_28602_170# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1504 vdd d1 a_19340_1994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1505 a_36297_2974# a_36309_2233# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1506 a_30921_2768# a_31174_2755# a_29905_3126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1507 gnd d3 a_13824_6444# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1508 gnd a_29859_4461# a_29651_4461# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1509 a_10811_1906# a_10816_1520# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1510 a_21618_5885# a_21620_5786# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1511 a_7074_5251# a_6965_5251# a_7173_5251# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1512 a_3134_3176# a_3391_2986# a_3079_3737# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1513 a_16755_7961# a_17559_7780# a_17728_7338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1514 gnd d0 a_4390_5743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1515 a_35081_2511# a_35279_3526# a_35234_3539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1516 a_27392_4568# a_27179_4568# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1517 a_11494_4065# a_11073_4065# a_10797_3965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1518 a_8410_4136# a_8667_3946# a_8364_3539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1519 a_31885_96# a_31672_96# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1520 gnd a_19313_6890# a_19105_6890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1521 a_34043_5251# a_33622_5251# a_33949_5370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1522 a_37861_1074# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1523 a_21633_3443# a_22114_3613# a_22322_3613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1524 a_39238_3392# a_38856_3834# a_38264_3600# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1525 gnd a_35334_2498# a_35126_2498# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1526 vdd d2 a_3336_3547# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1527 a_5911_3055# a_5698_3055# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1528 a_32767_5578# a_32554_5578# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1529 a_26926_867# a_27412_651# a_27620_651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1530 a_1672_7232# a_1459_7232# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1531 a_30914_5140# a_30910_5317# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1532 vdd a_15045_7145# a_14837_7145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1533 a_32547_6557# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1534 a_16080_3845# a_16085_3459# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1535 a_5705_2076# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1536 gnd d0 a_36530_8097# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1537 a_37548_7832# a_38037_7932# a_38245_7932# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1538 gnd d1 a_3391_2986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1539 a_636_1682# a_423_1682# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1540 a_2041_4308# a_1644_2383# a_1912_1355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1541 a_19076_3163# a_19333_2973# a_19021_3724# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1542 gnd a_4396_5177# a_4188_5177# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1543 a_833_4057# a_412_4057# a_136_4239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1544 a_35284_3959# a_36342_4180# a_36293_4370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1545 a_15904_140# a_15795_140# a_10504_125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1546 a_40358_2667# a_40572_1545# a_40523_1735# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1547 a_28628_2333# a_28415_2333# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1548 gnd a_3398_2007# a_3190_2007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1549 vdd d3 a_35314_6415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1550 a_8356_5496# a_8451_5903# a_8406_5916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1551 a_27608_2611# a_27187_2611# a_26921_2443# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1552 a_24603_7868# a_25661_8089# a_25612_8279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1553 a_27163_7924# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1554 gnd a_40835_984# a_40627_984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1555 a_34982_4680# a_35126_2498# a_35081_2511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1556 a_13587_2717# a_13801_1595# a_13752_1785# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1557 vdd a_30137_7834# a_29929_7834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1558 a_10809_2287# a_11298_2105# a_11506_2105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1559 a_23535_6271# a_23114_6271# a_23382_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1560 a_1719_4308# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1561 gnd a_41810_7661# a_41602_7661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1562 gnd d4 a_40520_4469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1563 a_41591_1408# a_41594_816# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1564 a_20089_3397# a_20346_3207# a_19080_2986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1565 a_1781_7232# a_1409_6812# a_818_6993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1566 a_30910_5317# a_30913_4725# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1567 a_16090_2266# a_16090_1984# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1568 a_36294_5169# a_36290_5346# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1569 vdd a_13749_4519# a_13541_4519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1570 a_17661_4295# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1571 a_21631_2947# a_21633_2848# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1572 gnd a_41554_8266# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1573 a_8191_6428# a_8389_7443# a_8344_7456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1574 a_7062_7211# a_6690_6791# a_6098_6557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1575 a_40558_5091# a_41619_4720# a_41574_4733# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1576 a_30917_2945# a_31174_2755# a_29905_3126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1577 vdd d3 a_13824_6444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1578 a_10789_6204# a_10789_5922# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1579 vdd a_29859_4461# a_29651_4461# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1580 a_38062_3034# a_37849_3034# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1581 a_25631_3947# a_25888_3757# a_24619_4128# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1582 a_4151_3233# a_4147_3410# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1583 a_36309_2233# a_36562_2220# a_35296_1999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1584 vdd d0 a_4390_5743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1585 a_25628_6142# a_25881_6129# a_24615_5908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1586 a_1479_3315# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1587 a_38281_659# a_39086_893# a_39245_1313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1588 a_27588_6528# a_27167_6528# a_26894_6744# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1589 a_14811_2826# a_15064_2813# a_13795_3184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1590 a_121_7175# a_121_6893# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1591 a_39049_7751# a_38836_7751# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1592 a_40546_7051# a_40803_6861# a_40491_7612# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1593 a_21881_7530# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1594 a_17564_6799# a_17351_6799# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1595 a_14799_6179# a_14795_6356# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1596 a_20084_4762# a_20080_4939# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1597 a_11291_3084# a_11078_3084# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1598 a_6125_1661# a_6930_1895# a_7099_1453# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1599 a_4126_6912# a_4138_6171# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1600 a_17983_4295# a_17874_4295# a_18082_4295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1601 a_28212_885# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1602 a_33000_680# a_32579_680# a_32313_695# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1603 a_5414_5194# a_5903_5012# a_6111_5012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1604 a_19068_5120# a_20129_4749# a_20084_4762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1605 a_16075_5202# a_16564_5020# a_16772_5020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1606 a_11085_2105# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1607 a_22949_7203# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1608 a_35284_3959# a_36342_4180# a_36297_4193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1609 a_15795_140# a_15582_140# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1610 a_21633_2848# a_21640_2464# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1611 gnd a_9680_4180# a_9472_4180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1612 a_40358_2667# a_40572_1545# a_40527_1558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1613 a_3114_7093# a_3371_6903# a_3059_7654# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1614 a_6111_5012# a_6915_4831# a_7074_5251# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1615 gnd a_25905_816# a_25697_816# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1616 a_29701_2482# a_29899_3497# a_29850_3687# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1617 a_4147_3410# a_4150_2818# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1618 a_40515_3518# a_40610_3925# a_40565_3938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1619 a_5431_1877# a_5917_1661# a_6125_1661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1620 gnd d0 a_31182_2191# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1621 gnd a_35314_6415# a_35106_6415# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1622 gnd d0 a_31167_5127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1623 a_17743_3302# a_17634_3302# a_17842_3302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1624 vdd a_41810_7661# a_41602_7661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1625 a_31672_96# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1626 vdd d1 a_35517_7863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1627 vdd a_4391_6158# a_4183_6158# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1628 a_29854_3510# a_30107_3497# a_29701_2482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1629 a_5685_5993# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1630 a_17735_5259# a_17363_4839# a_16771_4605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1631 a_8112_4680# a_8369_4490# a_7434_199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1632 a_19056_7080# a_19313_6890# a_19001_7641# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1633 a_16786_1669# a_16365_1669# a_16097_1499# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1634 a_35242_1756# a_35346_1005# a_35297_1195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1635 a_28671_3265# a_28628_2333# a_28812_4258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1636 a_24553_7448# a_24648_7855# a_24603_7868# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1637 a_41565_5891# a_41575_5148# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1638 a_36305_2410# a_36562_2220# a_35296_1999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1639 a_28569_5341# a_28187_5783# a_27595_5549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1640 a_3130_4956# a_4188_5177# a_4139_5367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1641 a_32284_4912# a_32286_4813# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1642 gnd a_13824_6444# a_13616_6444# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1643 a_22127_2068# a_21914_2068# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1644 gnd d0 a_9677_5156# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1645 a_14812_3241# a_14808_3418# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1646 a_5416_5408# a_5897_5578# a_6105_5578# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1647 a_4162_858# a_4415_845# a_3146_1216# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1648 a_32760_6557# a_32547_6557# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1649 a_409_5033# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1650 a_32306_1491# a_32304_1277# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1651 vdd a_3336_3547# a_3128_3547# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1652 a_24636_1187# a_24893_997# a_24581_1748# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1653 gnd a_30119_1537# a_29911_1537# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1654 a_32554_5578# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1655 a_39344_1313# a_39289_2341# a_39473_4266# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1656 a_21611_7146# a_21611_6864# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1657 a_130_5815# a_616_5599# a_824_5599# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1658 vdd a_9680_4180# a_9472_4180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1659 a_14815_2439# a_15072_2249# a_13806_2028# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1660 a_28663_5222# a_28608_6250# a_28816_6250# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1661 a_40511_3695# a_40768_3505# a_40362_2490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1662 a_423_1682# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1663 a_24611_6085# a_24868_5895# a_24565_5488# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1664 vdd d0 a_41848_1218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1665 a_29916_1970# a_30974_2191# a_30929_2204# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1666 a_28415_2333# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1667 a_32286_4813# a_32289_4432# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1668 gnd a_25888_3757# a_25680_3757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1669 a_838_3076# a_1642_2895# a_1801_3315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1670 vdd a_35314_6415# a_35106_6415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1671 a_8419_2978# a_9477_3199# a_9428_3389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1672 a_14808_3418# a_14811_2826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1673 a_34195_199# a_33982_199# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1674 a_11270_6586# a_11057_6586# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1675 a_8211_2511# a_8409_3526# a_8360_3716# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1676 a_25621_7121# a_25617_7298# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1677 vdd d0 a_20353_2228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1678 gnd a_35479_5483# a_35271_5483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1679 a_41574_4733# a_41570_4910# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1680 a_10804_2885# a_11290_2669# a_11498_2669# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1681 a_9415_6327# a_9672_6137# a_8406_5916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1682 a_35264_7876# a_36322_8097# a_36277_8110# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1683 a_22308_6964# a_23112_6783# a_23271_7203# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1684 a_26924_1248# a_27413_1066# a_27621_1066# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1685 a_29681_6399# a_29879_7414# a_29830_7604# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1686 vdd a_13824_6444# a_13616_6444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1687 vdd d0 a_9677_5156# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1688 a_28564_5222# a_28455_5222# a_28663_5222# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1689 a_29602_4651# a_29746_2469# a_29701_2482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1690 a_32567_2640# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1691 a_25647_1810# a_25643_1987# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1692 gnd d0 a_15071_1834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1693 a_9407_8110# a_10777_8164# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1694 a_28405_4802# a_28192_4802# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1695 a_36301_2797# a_36554_2784# a_35285_3155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1696 gnd a_35239_4490# a_35031_4490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1697 a_38873_893# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1698 gnd d2 a_19258_7451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1699 a_30902_7100# a_31155_7087# a_29889_6866# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1700 a_9444_1252# a_9697_1239# a_8431_1018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1701 a_27407_1632# a_27194_1632# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1702 a_25617_7298# a_25620_6706# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1703 a_11490_4626# a_11069_4626# a_10799_4461# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1704 a_38836_7751# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1705 a_4145_3799# a_4398_3786# a_3129_4157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1706 a_23296_3405# a_22914_3847# a_22322_3613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1707 a_17834_5259# a_17413_5259# a_17735_5259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1708 gnd d0 a_25885_4733# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1709 a_12573_1363# a_12152_1363# a_12479_1482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1710 a_16060_7762# a_16065_7376# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1711 a_17351_6799# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1712 gnd d0 a_41831_4159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1713 a_5697_2640# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1714 a_35222_5673# a_35326_4922# a_35277_5112# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1715 a_37575_3430# a_38056_3600# a_38264_3600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1716 a_22894_7764# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1717 a_22314_5570# a_21893_5570# a_21625_5400# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1718 gnd d0 a_4404_3220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1719 a_21606_7845# a_22095_7945# a_22303_7945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1720 a_40553_6072# a_41614_5701# a_41565_5891# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1721 vdd a_15060_4209# a_14852_4209# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1722 a_23531_4279# a_23134_2354# a_23402_1326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1723 a_849_701# a_428_701# a_155_917# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1724 a_11077_2669# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1725 gnd d1 a_40810_5882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1726 a_13732_5702# a_13836_4951# a_13791_4964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1727 a_428_701# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1728 a_20089_3397# a_20092_2805# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1729 a_22339_672# a_21918_672# a_21652_687# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1730 gnd a_4411_2241# a_4203_2241# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1731 a_32964_7953# a_32543_7953# a_32267_7853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1732 a_13736_5525# a_13831_5932# a_13782_6122# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1733 a_8211_2511# a_8409_3526# a_8364_3539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1734 a_29905_3126# a_30966_2755# a_30917_2945# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1735 a_17346_7780# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1736 a_3121_6114# a_4182_5743# a_4133_5933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1737 gnd d1 a_30162_2936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1738 vdd a_4384_7137# a_4176_7137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1739 vdd a_35479_5483# a_35271_5483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1740 gnd a_31167_5127# a_30959_5127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1741 gnd d0 a_9671_5722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1742 a_31994_96# a_37072_111# a_34403_199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1743 a_33793_2874# a_33580_2874# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1744 vdd d1 a_19320_5911# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1745 a_135_5429# a_133_5215# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1746 gnd a_30169_1957# a_29961_1957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1747 vdd a_9660_8097# a_9452_8097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1748 a_14782_7901# a_14792_7158# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1749 vdd a_35517_7863# a_35309_7863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1750 a_41574_4349# a_41831_4159# a_40565_3938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1751 a_37072_111# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1752 a_39477_6258# a_39056_6258# a_39324_5230# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1753 a_33587_1895# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1754 gnd d0 a_20345_2792# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1755 a_5677_6557# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1756 a_29681_6399# a_29879_7414# a_29834_7427# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1757 a_9411_6714# a_9664_6701# a_8395_7072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1758 a_28552_7182# a_28180_6762# a_27588_6528# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1759 a_12702_4316# a_12593_4316# a_12801_4316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1760 a_1637_3876# a_1424_3876# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1761 a_32299_2258# a_32788_2076# a_32996_2076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1762 a_30925_2381# a_30928_1789# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1763 a_11474_7982# a_11053_7982# a_10777_7882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1764 a_27603_3592# a_27182_3592# a_26914_3422# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1765 a_3079_3737# a_3183_2986# a_3134_3176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1766 a_36297_2974# a_36554_2784# a_35285_3155# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1767 a_22120_3047# a_21907_3047# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1768 a_8399_6895# a_9457_7116# a_9408_7306# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1769 a_22327_2632# a_21906_2632# a_21633_2848# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1770 a_22969_3286# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1771 vdd d0 a_9696_824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1772 a_1857_2383# a_1644_2383# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1773 vdd d2 a_19258_7451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1774 a_8364_3539# a_8459_3946# a_8410_4136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1775 a_27396_4007# a_27183_4007# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1776 a_12706_6308# a_12285_6308# a_12541_7240# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1777 a_19017_5504# a_19270_5491# a_18848_6613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1778 a_4141_3976# a_4398_3786# a_3129_4157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1779 vdd d0 a_25885_4733# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1780 vdd d1 a_8672_2965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1781 a_21626_4210# a_21626_3928# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1782 vdd d0 a_31161_5693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1783 a_8410_4136# a_9471_3765# a_9422_3955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1784 a_17579_3863# a_17366_3863# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1785 a_12462_3323# a_12353_3323# a_12561_3323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1786 a_40582_997# a_40835_984# a_40523_1735# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1787 vdd d0 a_4404_3220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1788 a_4137_5756# a_4133_5933# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1789 a_19021_3724# a_19125_2973# a_19076_3163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1790 gnd d0 a_41847_803# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1791 vdd a_4411_2241# a_4203_2241# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1792 a_16755_7961# a_16334_7961# a_16058_8143# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1793 gnd a_9676_4741# a_9468_4741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1794 a_27601_4983# a_28405_4802# a_28564_5222# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1795 a_38249_6536# a_37828_6536# a_37555_6752# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1796 vdd a_41848_1218# a_41640_1218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1797 a_26921_1848# a_27407_1632# a_27615_1632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1798 a_7067_7330# a_6685_7772# a_6094_7953# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1799 a_30901_6685# a_30897_6862# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1800 a_38057_4015# a_37844_4015# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1801 a_40582_997# a_41640_1218# a_41591_1408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1802 a_29905_3126# a_30966_2755# a_30921_2768# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1803 a_6903_6791# a_6690_6791# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1804 a_3121_6114# a_4182_5743# a_4137_5756# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1805 a_16077_5416# a_16075_5202# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1806 a_32289_4432# a_32287_4218# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1807 a_29884_7847# a_30137_7834# a_29834_7427# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1808 vdd d0 a_9671_5722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1809 vdd d1 a_40818_3925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1810 a_39213_7190# a_39104_7190# a_39312_7190# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1811 a_7421_4287# a_7000_4287# a_7322_4287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1812 gnd d0 a_36547_5156# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1813 gnd d0 a_9697_1239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1814 vdd a_20353_2228# a_20145_2228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1815 a_13795_3184# a_14856_2813# a_14807_3003# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1816 a_17760_1461# a_17378_1903# a_16786_1669# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1817 a_17559_7780# a_17346_7780# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1818 a_11057_6586# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1819 a_25648_1006# a_25905_816# a_24636_1187# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1820 a_19092_1026# a_19345_1013# a_19033_1764# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1821 a_20073_7137# a_20069_7314# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1822 a_14791_6743# a_15044_6730# a_13775_7101# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1823 a_24620_4927# a_25678_5148# a_25629_5338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1824 a_1900_3315# a_1479_3315# a_1806_3434# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1825 a_8399_6895# a_9457_7116# a_9412_7129# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1826 a_16070_5901# a_16559_6001# a_16767_6001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1827 a_19092_1026# a_20150_1247# a_20101_1437# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1828 gnd d0 a_36561_1805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1829 a_6105_5578# a_6910_5812# a_7079_5370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1830 gnd d0 a_31162_6108# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1831 a_7181_3294# a_6760_3294# a_7082_3294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1832 a_26906_5379# a_27387_5549# a_27595_5549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1833 a_27400_2611# a_27187_2611# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1834 a_28192_4802# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1835 a_25652_829# a_25905_816# a_24636_1187# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1836 gnd a_19258_7451# a_19050_7451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1837 gnd d0 a_15057_5185# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1838 a_8410_4136# a_9471_3765# a_9426_3778# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1839 a_17755_1342# a_17383_922# a_16792_1103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1840 a_27194_1632# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1841 a_24631_2168# a_25692_1797# a_25643_1987# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1842 a_33843_3294# a_33630_3294# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1843 a_32775_3621# a_32562_3621# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1844 a_33567_5812# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1845 a_12454_5280# a_12082_4860# a_11491_5041# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1846 a_8112_4680# a_8256_2498# a_8207_2688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1847 a_37560_6154# a_37560_5872# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1848 a_133_4933# a_135_4834# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1849 a_5436_896# a_5922_680# a_6130_680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1850 a_17740_5378# a_17358_5820# a_16767_6001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1851 vdd a_9676_4741# a_9468_4741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1852 a_12298_3884# a_12085_3884# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1853 gnd a_4404_3220# a_4196_3220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1854 gnd a_35499_1566# a_35291_1566# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1855 a_20069_7314# a_20072_6722# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1856 a_36277_6891# a_36534_6701# a_35265_7072# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1857 a_5422_2955# a_5911_3055# a_6119_3055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1858 a_1786_7351# a_1672_7232# a_1880_7232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1859 gnd d2 a_3336_3547# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1860 a_40523_1735# a_40627_984# a_40582_997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1861 a_30924_1966# a_30934_1223# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1862 a_2252_220# a_1831_220# a_2153_220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1863 a_22099_6549# a_21886_6549# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1864 a_38073_659# a_37860_659# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1865 a_16584_1103# a_16371_1103# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1866 a_4121_7893# a_4378_7703# a_3109_8074# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1867 a_12283_6820# a_12070_6820# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1868 a_7099_1453# a_6985_1334# a_7193_1334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1869 a_32568_3055# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1870 vdd d4 a_8369_4490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1871 a_11285_3650# a_11072_3650# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1872 a_141_3258# a_630_3076# a_838_3076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1873 a_4163_1273# a_4159_1450# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1874 a_13571_6457# a_13824_6444# a_13496_4532# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1875 a_12077_5841# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1876 a_29842_5644# a_29946_4893# a_29897_5083# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1877 vdd d0 a_36547_5156# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1878 a_11499_3084# a_12303_2903# a_12462_3323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1879 gnd a_30162_2936# a_29954_2936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1880 gnd a_25869_8089# a_25661_8089# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1881 a_9434_1995# a_9691_1805# a_8422_2176# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1882 a_35301_1018# a_36359_1239# a_36314_1252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1883 a_33580_2874# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1884 a_4126_8131# a_5397_8135# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1885 a_32755_7538# a_32542_7538# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1886 a_41589_1797# a_41585_1974# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1887 gnd a_14009_1595# a_13801_1595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1888 a_22107_5985# a_21894_5985# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1889 a_6111_5012# a_5690_5012# a_5414_5194# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1890 a_19088_1203# a_19345_1013# a_19033_1764# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1891 a_14787_6920# a_15044_6730# a_13775_7101# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1892 a_38856_3834# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1893 gnd a_20345_2792# a_20137_2792# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1894 a_1424_3876# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1895 a_624_3642# a_411_3642# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1896 a_37568_4197# a_38057_4015# a_38265_4015# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1897 a_13806_2028# a_14864_2249# a_14819_2262# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1898 gnd a_13749_4519# a_13541_4519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1899 a_11078_3084# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1900 a_830_5033# a_409_5033# a_133_4933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1901 a_9427_4193# a_9423_4370# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1902 vdd d0 a_15057_5185# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1903 a_26907_3907# a_26909_3808# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1904 a_37573_3216# a_37573_2934# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1905 vdd a_19258_7451# a_19050_7451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1906 a_16564_5020# a_16351_5020# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1907 a_27183_4007# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1908 a_32287_3936# a_32289_3837# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1909 a_33001_1095# a_33805_914# a_33964_1334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1910 a_27620_651# a_27199_651# a_26933_666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1911 a_25635_3770# a_25888_3757# a_24619_4128# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1912 a_4159_1450# a_4162_858# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1913 vdd d0 a_20325_6709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1914 a_11265_7567# a_11052_7567# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1915 gnd a_8609_5483# a_8401_5483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1916 a_11478_6586# a_12283_6820# a_12442_7240# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1917 a_9439_1014# a_5443_695# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1918 a_27388_5964# a_27175_5964# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1919 a_17366_3863# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1920 a_417_3076# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1921 a_25648_1006# a_21652_687# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1922 vdd a_4404_3220# a_4196_3220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1923 vdd a_35499_1566# a_35291_1566# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1924 gnd d0 a_36541_5722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1925 a_7161_7211# a_6740_7211# a_7062_7211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1926 a_40338_6584# a_40595_6394# a_40267_4482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1927 a_38256_5557# a_37835_5557# a_37567_5387# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1928 a_844_1682# a_423_1682# a_150_1898# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1929 a_1912_1355# a_1857_2383# a_2041_4308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1930 a_19068_5120# a_20129_4749# a_20080_4939# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1931 vdd d1 a_24873_4914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1932 a_28242_5222# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1933 a_27615_1632# a_28420_1866# a_28589_1424# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1934 a_6690_6791# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1935 a_33823_7211# a_33610_7211# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1936 a_24611_6085# a_25672_5714# a_25623_5904# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1937 a_9423_4370# a_9426_3778# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1938 a_23535_6271# a_23422_4279# a_23630_4279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1939 a_8116_4503# a_8236_6415# a_8187_6605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1940 a_13567_6634# a_13824_6444# a_13496_4532# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1941 a_26904_5165# a_27393_4983# a_27601_4983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1942 a_35226_5496# a_35321_5903# a_35272_6093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1943 vdd a_40818_3925# a_40610_3925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1944 vdd a_9696_824# a_9488_824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1945 a_11485_5607# a_11064_5607# a_10791_5823# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1946 a_34192_4287# a_33795_2362# a_34063_1334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1947 gnd d1 a_35542_2965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1948 a_29889_6866# a_30947_7087# a_30898_7277# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1949 gnd a_36547_5156# a_36339_5156# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1950 gnd d0 a_4399_4201# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1951 gnd d0 a_15051_5751# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1952 a_27621_1066# a_28425_885# a_28584_1305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1953 gnd a_35549_1986# a_35341_1986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1954 a_37841_4991# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1955 a_3138_2999# a_4196_3220# a_4147_3410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1956 a_32304_1277# a_32304_995# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1957 gnd a_24673_2490# a_24465_2490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1958 gnd a_4391_6158# a_4183_6158# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1959 vdd d3 a_3183_2519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1960 a_24569_3708# a_24673_2957# a_24624_3147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1961 a_23296_3405# a_23182_3286# a_23390_3286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1962 a_16072_6397# a_16551_6565# a_16759_6565# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1963 a_17773_207# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1964 a_12333_7240# a_12120_7240# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1965 a_5424_3451# a_5905_3621# a_6113_3621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1966 a_29854_3510# a_29949_3917# a_29900_4107# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1967 gnd a_31162_6108# a_30954_6108# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1968 gnd d1 a_14052_2994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1969 a_38269_2619# a_37848_2619# a_37575_2835# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1970 vdd a_8609_5483# a_8401_5483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1971 gnd a_15057_5185# a_14849_5185# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1972 a_28475_1305# a_28262_1305# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1973 a_22308_6964# a_21887_6964# a_21611_7146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1974 a_3141_2197# a_4202_1826# a_4157_1839# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1975 a_33630_3294# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1976 gnd d1 a_19328_3954# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1977 a_32562_3621# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1978 a_17723_7219# a_17351_6799# a_16760_6980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1979 a_25633_5161# a_25629_5338# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1980 a_23209_4279# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1981 a_138_3858# a_624_3642# a_832_3642# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1982 a_34196_6279# a_33775_6279# a_34031_7211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1983 vdd d0 a_36541_5722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1984 a_33788_3855# a_33575_3855# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1985 vdd d0 a_9691_1805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1986 a_32274_6773# a_32760_6557# a_32968_6557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1987 a_16774_3629# a_16353_3629# a_16080_3845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1988 a_27621_1066# a_27200_1066# a_26924_1248# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1989 a_5397_7853# a_5399_7754# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1990 a_23382_5243# a_22961_5243# a_23283_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1991 a_8394_7876# a_9452_8097# a_9403_8287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1992 a_12085_3884# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1993 a_11058_7001# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1994 gnd a_3336_3547# a_3128_3547# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1995 a_153_1016# a_642_1116# a_850_1116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1996 a_28557_7301# a_28175_7743# a_27584_7924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1997 a_20996_n19# a_20887_n19# vout vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1998 a_24611_6085# a_25672_5714# a_25627_5727# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1999 a_32996_2076# a_32575_2076# a_32299_1976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2000 a_14819_2262# a_15072_2249# a_13806_2028# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2001 a_22115_4028# a_21902_4028# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2002 a_10779_7783# a_11265_7567# a_11473_7567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2003 a_12070_6820# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2004 a_8116_4503# a_8236_6415# a_8191_6428# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2005 a_16371_1103# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2006 a_16092_2480# a_16090_2266# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2007 a_40570_2957# a_41628_3178# a_41583_3191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2008 a_20105_1260# a_20101_1437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2009 a_32279_6175# a_32768_5993# a_32976_5993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2010 a_28911_4258# a_28490_4258# a_28812_4258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2011 a_11072_3650# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2012 gnd d0 a_41848_1218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2013 a_40541_8032# a_40798_7842# a_40495_7435# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2014 gnd a_8659_5903# a_8451_5903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2015 a_35264_7876# a_35517_7863# a_35214_7456# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2016 a_397_6993# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2017 a_12442_7240# a_12333_7240# a_12541_7240# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2018 a_10791_6418# a_10789_6204# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2019 vdd a_36547_5156# a_36339_5156# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2020 a_22100_6964# a_21887_6964# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2021 vdd d0 a_15051_5751# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2022 a_21623_4904# a_22112_5004# a_22320_5004# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2023 a_1831_220# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2024 a_25629_5338# a_25632_4746# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2025 a_123_7389# a_604_7559# a_812_7559# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2026 a_27376_7924# a_27163_7924# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2027 a_138_4453# a_136_4239# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2028 a_3138_2999# a_4196_3220# a_4151_3233# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2029 gnd d0 a_20353_2228# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2030 a_17779_6287# a_17566_6287# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2031 a_22319_4589# a_23124_4823# a_23283_5243# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2032 a_123_7389# a_121_7175# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2033 a_8422_2176# a_8679_1986# a_8376_1579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2034 a_9419_6150# a_9672_6137# a_8406_5916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2035 a_411_3642# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2036 a_35234_3539# a_35329_3946# a_35284_3959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2037 a_39250_1432# a_38868_1874# a_38276_1640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2038 a_21645_1483# a_22126_1653# a_22334_1653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2039 a_27595_5549# a_28400_5783# a_28569_5341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2040 a_28671_3265# a_28250_3265# a_28572_3265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2041 a_1684_5272# a_1471_5272# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2042 a_39572_4266# a_39151_4266# a_39477_6258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2043 a_37560_5872# a_38049_5972# a_38257_5972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2044 vdd a_15057_5185# a_14849_5185# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2045 vdd d1 a_3386_3967# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2046 a_41591_1408# a_41848_1218# a_40582_997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2047 a_20101_1437# a_20104_845# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2048 a_6898_7772# a_6685_7772# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2049 a_13774_7905# a_14027_7892# a_13724_7485# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2050 a_5414_5194# a_5414_4912# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2051 a_16351_5020# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2052 a_9422_3955# a_9432_3212# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2053 a_17842_3302# a_17421_3302# a_17743_3302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2054 vdd a_20325_6709# a_20117_6709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2055 a_32304_995# a_32306_896# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2056 a_29602_4651# a_29746_2469# a_29697_2659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2057 a_11052_7567# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2058 a_27381_6943# a_27168_6943# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2059 a_5709_680# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2060 a_10814_1024# a_10816_925# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2061 a_19087_2007# a_19340_1994# a_19037_1587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2062 a_27175_5964# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2063 vdd d1 a_30142_6853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2064 a_30904_5883# a_30914_5140# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2065 a_26912_2926# a_27401_3026# a_27609_3026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2066 a_23276_7322# a_23162_7203# a_23370_7203# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2067 gnd d0 a_41815_6680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2068 a_24636_1187# a_25697_816# a_25652_829# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2069 a_37587_875# a_37594_674# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2070 gnd d3 a_19125_2506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2071 a_29880_8024# a_30941_7653# a_30892_7843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2072 vdd a_30149_5874# a_29941_5874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2073 a_20084_4378# a_20087_3786# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2074 a_36313_837# a_36566_824# a_35297_1195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2075 a_16346_6001# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2076 a_6093_7538# a_5672_7538# a_5404_7368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2077 a_13775_7101# a_14836_6730# a_14787_6920# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2078 a_28589_1424# a_28475_1305# a_28683_1305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2079 gnd d1 a_14032_6911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2080 a_1793_5272# a_1421_4852# a_830_5033# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2081 vdd a_24873_4914# a_24665_4914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2082 a_20101_1437# a_20358_1247# a_19092_1026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2083 a_32793_1095# a_32580_1095# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2084 gnd d0 a_20320_7690# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2085 a_33610_7211# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2086 gnd a_14039_5932# a_13831_5932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2087 a_6973_3294# a_6760_3294# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2088 a_850_1116# a_429_1116# a_153_1016# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2089 a_17822_7219# a_17401_7219# a_17728_7338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2090 a_38074_1074# a_37861_1074# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2091 a_27601_4983# a_27180_4983# a_26904_5165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2092 gnd a_35542_2965# a_35334_2965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2093 a_8344_7456# a_8439_7863# a_8394_7876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2094 vdd a_3391_2986# a_3183_2986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2095 gnd a_4384_7137# a_4176_7137# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2096 a_22914_3847# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2097 a_14823_866# a_15076_853# a_13807_1224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2098 a_17854_1342# a_17799_2370# a_17983_4295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2099 a_32989_3055# a_33793_2874# a_33952_3294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2100 gnd a_3386_3967# a_3178_3967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2101 a_21626_4210# a_22115_4028# a_22323_4028# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2102 a_150_1898# a_155_1512# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2103 a_41578_4172# a_41831_4159# a_40565_3938# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2104 a_21893_5570# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2105 a_39245_1313# a_39136_1313# a_39344_1313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2106 a_11303_1124# a_11090_1124# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2107 a_1813_1355# a_1704_1355# a_1912_1355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2108 a_12120_7240# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2109 a_40557_5895# a_40810_5882# a_40507_5475# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2110 a_11494_4065# a_12298_3884# a_12467_3442# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2111 a_40578_1174# a_41639_803# a_41594_816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2112 a_155_1512# a_636_1682# a_844_1682# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2113 a_605_7974# a_392_7974# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2114 vdd d0 a_4379_8118# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2115 a_21613_7360# a_21611_7146# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2116 a_16579_2084# a_16366_2084# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2117 a_12278_7801# a_12065_7801# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2118 a_30913_4725# a_31166_4712# a_29897_5083# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2119 a_19005_7464# a_19100_7871# a_19051_8061# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2120 a_30913_4725# a_30909_4902# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2121 gnd a_14052_2994# a_13844_2994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2122 vdd d1 a_30174_976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2123 a_16090_1984# a_16092_1885# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2124 a_3126_5133# a_3383_4943# a_3071_5694# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2125 gnd d0 a_20357_832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2126 a_28262_1305# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2127 vdd a_25900_1797# a_25692_1797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2128 a_29917_1166# a_30174_976# a_29862_1727# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2129 a_641_701# a_428_701# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2130 vdd a_24653_6407# a_24445_6407# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2131 gnd a_19328_3954# a_19120_3954# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2132 a_12593_4316# a_12380_4316# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2133 a_33575_3855# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2134 a_22131_672# a_21918_672# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2135 a_40527_1558# a_40622_1965# a_40577_1978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2136 a_25616_8102# a_25869_8089# a_24603_7868# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2137 a_29880_8024# a_30941_7653# a_30896_7666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2138 vdd d0 a_41815_6680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2139 a_11486_6022# a_11065_6022# a_10789_5922# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2140 a_8402_6093# a_8659_5903# a_8356_5496# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2141 a_20088_4201# a_20341_4188# a_19075_3967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2142 a_32287_3936# a_32776_4036# a_32984_4036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2143 a_121_7175# a_610_6993# a_818_6993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2144 a_17755_1342# a_17646_1342# a_17854_1342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2145 gnd d3 a_3163_6436# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2146 a_5903_5012# a_5690_5012# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2147 a_121_6893# a_123_6794# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2148 a_13775_7101# a_14836_6730# a_14791_6743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2149 a_5419_3837# a_5424_3451# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2150 a_817_6578# a_1622_6812# a_1781_7232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2151 gnd a_8652_6882# a_8444_6882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2152 a_19068_5120# a_19325_4930# a_19013_5681# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2153 a_825_6014# a_404_6014# a_128_6196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2154 gnd d1 a_3383_4943# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2155 a_37548_8114# a_38037_7932# a_38245_7932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2156 a_19067_5924# a_19320_5911# a_19017_5504# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2157 a_12353_3323# a_12140_3323# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2158 gnd a_41848_1218# a_41640_1218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2159 a_16092_1885# a_16097_1499# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2160 a_21906_2632# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2161 a_6099_6972# a_6903_6791# a_7062_7211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2162 gnd d3 a_19105_6423# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2163 a_8415_3155# a_8672_2965# a_8360_3716# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2164 vdd d0 a_4415_845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2165 a_27163_7924# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2166 a_17566_6287# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2167 gnd d0 a_25894_3191# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2168 a_4158_1035# a_4415_845# a_3146_1216# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2169 gnd a_20353_2228# a_20145_2228# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2170 a_39233_3273# a_38861_2853# a_38269_2619# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2171 gnd d0 a_31170_4151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2172 a_16775_4044# a_16354_4044# a_16078_3944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2173 a_32772_4597# a_32559_4597# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2174 a_26914_3422# a_27395_3592# a_27603_3592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2175 a_11499_3084# a_11078_3084# a_10802_3266# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2176 a_5429_2258# a_5429_1976# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2177 a_7087_3413# a_6705_3855# a_6113_3621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2178 a_36293_4370# a_36296_3778# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2179 a_6953_7211# a_6740_7211# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2180 a_1471_5272# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2181 a_30909_4902# a_31166_4712# a_29897_5083# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2182 a_6685_7772# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2183 a_37828_6536# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2184 a_12705_228# a_12492_228# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2185 a_18082_4295# a_17986_207# a_15904_140# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2186 a_5397_7853# a_5886_7953# a_6094_7953# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2187 vdd a_3371_6903# a_3163_6903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2188 a_40263_4659# a_40407_2477# a_40362_2490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2189 a_9439_1014# a_9696_824# a_8427_1195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2190 a_17834_5259# a_17779_6287# a_17987_6287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2191 a_3133_3980# a_4191_4201# a_4142_4391# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2192 a_7000_4287# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2193 a_40561_4115# a_40818_3925# a_40515_3518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2194 a_34008_2362# a_33795_2362# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2195 vdd d3 a_3163_6436# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2196 vdd a_30142_6853# a_29934_6853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2197 a_23742_191# a_26624_103# a_26832_103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2198 gnd a_41815_6680# a_41607_6680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2199 gnd a_19125_2506# a_18917_2506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2200 a_39213_7190# a_38841_6770# a_38250_6951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2201 a_11474_7982# a_12278_7801# a_12447_7359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2202 a_28816_6250# a_28395_6250# a_28663_5222# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2203 a_16558_5586# a_16345_5586# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2204 a_39136_1313# a_38923_1313# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2205 a_16338_6565# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2206 a_22111_4589# a_21898_4589# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2207 gnd d2 a_8629_1566# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2208 gnd a_14032_6911# a_13824_6911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2209 a_35276_5916# a_36334_6137# a_36289_6150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2210 vdd d0 a_36555_3199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2211 a_18777_4511# a_19030_4498# a_18095_207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2212 a_32580_1095# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2213 a_21611_6864# a_21613_6765# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2214 a_4138_4952# a_4146_4214# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2215 a_32542_7538# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2216 a_6760_3294# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2217 vdd d3 a_19105_6423# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2218 a_12518_2391# a_12305_2391# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2219 a_24628_2970# a_25686_3191# a_25641_3204# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2220 a_25644_2402# a_25647_1810# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2221 vdd d0 a_31170_4151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2222 a_33988_6279# a_33775_6279# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2223 a_35301_1018# a_36359_1239# a_36310_1429# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2224 a_14811_2826# a_14807_3003# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2225 a_32968_6557# a_32547_6557# a_32281_6389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2226 a_38848_5791# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2227 a_23308_1445# a_22926_1887# a_22334_1653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2228 a_38261_4576# a_39066_4810# a_39225_5230# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2229 vdd d0 a_15065_3228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2230 a_28425_885# a_28212_885# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2231 a_11090_1124# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2232 gnd d0 a_41843_2199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2233 a_37587_1470# a_38068_1640# a_38276_1640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2234 a_392_7974# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2235 a_9402_7872# a_9412_7129# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2236 a_23630_4279# a_23209_4279# a_23535_6271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2237 gnd d0 a_4416_1260# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2238 a_837_2661# a_416_2661# a_150_2493# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2239 a_16366_2084# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2240 a_13806_2028# a_14864_2249# a_14815_2439# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2241 a_12065_7801# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2242 a_6130_680# a_5709_680# a_5443_695# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2243 gnd a_40595_6394# a_40387_6394# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2244 gnd a_20357_832# a_20149_832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2245 a_32976_5993# a_32555_5993# a_32279_5893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2246 a_16065_7376# a_16063_7162# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2247 a_12380_4316# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2248 vdd d1 a_30157_3917# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2249 a_39332_3273# a_38911_3273# a_39233_3273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2250 vdd a_41815_6680# a_41607_6680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2251 a_38264_3600# a_37843_3600# a_37575_3430# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2252 a_11478_6586# a_11057_6586# a_10791_6418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2253 gnd d1 a_30174_976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2254 vdd d1 a_35522_6882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2255 a_27583_7509# a_27162_7509# a_26894_7339# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2256 gnd a_3163_6436# a_2955_6436# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2257 a_5690_5012# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2258 a_14823_866# a_14819_1043# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2259 vdd d2 a_8629_1566# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2260 vdd d1 a_3366_7884# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2261 a_36292_3955# a_36302_3212# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2262 a_24549_7625# a_24653_6874# a_24608_6887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2263 vdd d0 a_15076_853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2264 a_817_6578# a_396_6578# a_123_6794# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2265 a_35265_7072# a_36326_6701# a_36277_6891# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2266 a_3083_3560# a_3178_3967# a_3133_3980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2267 a_20064_8295# a_20321_8105# a_19055_7884# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2268 gnd a_25880_5714# a_25672_5714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2269 a_14819_1043# a_15076_853# a_13807_1224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2270 a_22132_1087# a_21919_1087# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2271 a_13724_7485# a_13819_7892# a_13770_8082# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2272 a_29834_7427# a_29929_7834# a_29884_7847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2273 a_33937_7330# a_33823_7211# a_34031_7211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2274 a_8411_4935# a_9469_5156# a_9420_5346# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2275 a_23107_7764# a_22894_7764# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2276 gnd a_19105_6423# a_18897_6423# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2277 a_27408_2047# a_27195_2047# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2278 a_14792_7158# a_14788_7335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2279 a_9411_6714# a_9407_6891# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2280 a_10796_4842# a_11282_4626# a_11490_4626# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2281 gnd a_25894_3191# a_25686_3191# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2282 vdd d1 a_19308_7871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2283 a_37562_6368# a_37560_6154# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2284 a_21620_5786# a_21625_5400# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2285 a_23303_1326# a_23194_1326# a_23402_1326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2286 a_28420_1866# a_28207_1866# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2287 a_8422_2176# a_9483_1805# a_9434_1995# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2288 vdd d0 a_4416_1260# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2289 gnd a_24881_2957# a_24673_2957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2290 a_16070_5901# a_16072_5802# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2291 gnd d3 a_3183_2519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2292 a_5885_7538# a_5672_7538# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2293 a_24616_5104# a_24873_4914# a_24561_5665# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2294 a_32559_4597# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2295 a_20674_n19# d8 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2296 a_30928_1789# a_30924_1966# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2297 a_138_4453# a_621_4618# a_829_4618# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2298 a_36293_4754# a_36546_4741# a_35277_5112# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2299 a_4921_132# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2300 a_38069_2055# a_37856_2055# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2301 a_33795_2362# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2302 a_19076_3163# a_20137_2792# a_20092_2805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2303 a_29896_5887# a_30149_5874# a_29846_5467# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2304 a_23288_5362# a_22906_5804# a_22314_5570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2305 vdd a_3163_6436# a_2955_6436# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2306 a_16551_6565# a_16338_6565# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2307 a_25643_1987# a_25653_1244# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2308 gnd d0 a_41823_6116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2309 a_39225_5230# a_39116_5230# a_39324_5230# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2310 a_34083_4287# a_33870_4287# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2311 a_39081_1874# a_38868_1874# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2312 a_38054_4991# a_37841_4991# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2313 a_13807_1224# a_14868_853# a_14819_1043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2314 a_17983_4295# a_17586_2370# a_17842_3302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2315 a_36289_6150# a_36285_6327# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2316 a_30908_5706# a_31161_5693# a_29892_6064# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2317 a_21626_3928# a_21628_3829# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2318 a_16085_2864# a_16571_2648# a_16779_2648# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2319 vdd d0 a_25873_6693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2320 a_16072_5802# a_16077_5416# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2321 a_11069_4626# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2322 a_14803_4783# a_15056_4770# a_13787_5141# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2323 a_37394_111# a_39263_178# a_39572_4266# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2324 vdd a_36555_3199# a_36347_3199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2325 a_3113_7897# a_4171_8118# a_4126_8131# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2326 a_21606_8127# a_22095_7945# a_22303_7945# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2327 a_27589_6943# a_28393_6762# a_28552_7182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2328 vdd a_25880_5714# a_25672_5714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2329 a_39263_178# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2330 a_1912_1355# a_1491_1355# a_1818_1474# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2331 a_8411_4935# a_9469_5156# a_9424_5169# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2332 a_40267_4482# a_40387_6394# a_40338_6584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2333 a_22328_3047# a_21907_3047# a_21631_2947# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2334 vdd d0 a_9660_8097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2335 vdd a_19105_6423# a_18897_6423# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2336 a_29897_5083# a_30958_4712# a_30909_4902# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2337 a_40570_2957# a_41628_3178# a_41579_3368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2338 a_9434_1995# a_9444_1252# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2339 a_12305_2391# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2340 a_116_8156# a_116_7874# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2341 a_37575_3430# a_37573_3216# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2342 a_30929_985# a_31186_795# a_29917_1166# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2343 a_23630_4279# a_23534_191# a_23742_191# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2344 a_41554_8266# a_41557_7674# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2345 a_23370_7203# a_22949_7203# a_23276_7322# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2346 a_21887_6964# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2347 a_38841_6770# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2348 a_40503_5652# a_40607_4901# a_40558_5091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2349 a_33785_4831# a_33572_4831# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2350 a_23291_3286# a_22919_2866# a_22327_2632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2351 a_33775_6279# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2352 gnd a_19270_5491# a_19062_5491# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2353 a_20063_7880# a_20073_7137# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2354 a_16771_4605# a_16350_4605# a_16080_4440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2355 a_32787_1661# a_32574_1661# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2356 a_9426_3778# a_9679_3765# a_8410_4136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2357 a_32984_4036# a_32563_4036# a_32287_4218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2358 a_28577_3384# a_28195_3826# a_27603_3592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2359 a_22961_5243# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2360 gnd d0 a_36550_4180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2361 vdd a_15065_3228# a_14857_3228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2362 a_17854_1342# a_17433_1342# a_17760_1461# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2363 a_1629_5833# a_1416_5833# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2364 gnd a_41843_2199# a_41635_2199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2365 a_3071_5694# a_3175_4943# a_3126_5133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2366 a_22112_5004# a_21899_5004# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2367 gnd a_4416_1260# a_4208_1260# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2368 a_26887_7824# a_27376_7924# a_27584_7924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2369 a_36289_4931# a_36546_4741# a_35277_5112# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2370 a_19080_2986# a_20138_3207# a_20089_3397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2371 gnd d2 a_3348_1587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2372 a_14795_6356# a_14798_5764# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2373 vdd d3 a_35334_2498# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2374 a_16358_2648# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2375 a_12459_5399# a_12345_5280# a_12553_5280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2376 a_24623_3951# a_25681_4172# a_25632_4362# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2377 a_12295_4860# a_12082_4860# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2378 a_41595_1231# a_41848_1218# a_40582_997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2379 a_21643_1269# a_21643_987# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2380 vdd d1 a_8664_4922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2381 gnd d0 a_25874_7108# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2382 vdd a_30157_3917# a_29949_3917# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2383 a_34063_1334# a_33642_1334# a_33964_1334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2384 a_11297_1690# a_11084_1690# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2385 gnd d2 a_24806_7435# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2386 a_8402_6093# a_9463_5722# a_9414_5912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2387 vdd d0 a_41823_6116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2388 a_11494_4065# a_11073_4065# a_10797_4247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2389 gnd a_30174_976# a_29966_976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2390 a_24321_4672# a_24465_2490# a_24420_2503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2391 vdd a_35522_6882# a_35314_6882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2392 a_7326_6279# a_7213_4287# a_7421_4287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2393 a_39238_3392# a_38856_3834# a_38265_4015# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2394 a_16085_2864# a_16092_2480# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2395 a_837_2661# a_1642_2895# a_1801_3315# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2396 a_19013_5681# a_19117_4930# a_19068_5120# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2397 a_26933_666# a_27412_651# a_27620_651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2398 a_35292_2176# a_36353_1805# a_36308_1818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2399 gnd a_31149_7653# a_30941_7653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2400 a_1672_7232# a_1459_7232# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2401 a_2045_6300# a_1624_6300# a_1880_7232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2402 a_32767_5578# a_32554_5578# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2403 a_1642_2895# a_1429_2895# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2404 vdd d1 a_3398_2007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2405 a_14799_4960# a_15056_4770# a_13787_5141# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2406 vdd a_3366_7884# a_3158_7884# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2407 a_38868_1874# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2408 a_37580_2237# a_38069_2055# a_38277_2055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2409 vdd d3 a_13844_2527# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2410 a_32964_7953# a_33768_7772# a_33937_7330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2411 a_7326_6279# a_6905_6279# a_7173_5251# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2412 a_6918_3855# a_6705_3855# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2413 a_16755_7961# a_16334_7961# a_16058_7861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2414 a_29897_5083# a_30958_4712# a_30913_4725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2415 a_32304_995# a_32793_1095# a_33001_1095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2416 a_20105_1260# a_20358_1247# a_19092_1026# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2417 a_5416_5408# a_5414_5194# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2418 gnd a_35487_3526# a_35279_3526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2419 a_8360_3716# a_8464_2965# a_8415_3155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2420 a_27401_3026# a_27188_3026# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2421 a_7087_3413# a_6973_3294# a_7181_3294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2422 a_27608_2611# a_27187_2611# a_26914_2827# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2423 a_39061_5791# a_38848_5791# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2424 gnd d4 a_24578_4482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2425 a_16792_1103# a_17596_922# a_17755_1342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2426 a_27195_2047# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2427 a_17987_6287# a_17566_6287# a_17822_7219# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2428 a_26907_4189# a_26907_3907# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2429 vdd d0 a_20337_4749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2430 a_27620_651# a_28425_885# a_28584_1305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2431 a_17584_2882# a_17371_2882# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2432 a_9422_3955# a_9679_3765# a_8410_4136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2433 a_10809_2005# a_11298_2105# a_11506_2105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2434 vdd a_19308_7871# a_19100_7871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2435 a_23535_6271# a_23114_6271# a_23370_7203# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2436 vdd d0 a_36550_4180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2437 a_21606_8127# a_21606_7845# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2438 a_6099_6972# a_5678_6972# a_5402_7154# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2439 a_5922_680# a_5709_680# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2440 a_41562_6693# a_41815_6680# a_40546_7051# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2441 vdd a_4416_1260# a_4208_1260# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2442 a_5672_7538# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2443 a_24623_3951# a_25681_4172# a_25636_4185# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2444 a_7173_5251# a_6752_5251# a_7074_5251# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2445 a_38062_3034# a_37849_3034# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2446 a_18095_207# a_18822_4498# a_18773_4688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2447 gnd d0 a_4379_8118# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2448 vdd d2 a_24806_7435# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2449 a_4130_6735# a_4383_6722# a_3114_7093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2450 a_29889_6866# a_30142_6853# a_29830_7604# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2451 vdd d1 a_40823_2944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2452 a_8402_6093# a_9463_5722# a_9418_5735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2453 a_33835_5251# a_33622_5251# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2454 a_22322_3613# a_21901_3613# a_21633_3443# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2455 a_40561_4115# a_41622_3744# a_41573_3934# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2456 a_39049_7751# a_38836_7751# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2457 a_37573_2934# a_37575_2835# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2458 gnd d1 a_35554_1005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2459 vdd a_40830_1965# a_40622_1965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2460 vdd a_9691_1805# a_9483_1805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2461 vdd a_31149_7653# a_30941_7653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2462 gnd a_41823_6116# a_41615_6116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2463 a_5414_4912# a_5903_5012# a_6111_5012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2464 a_19060_6903# a_20118_7124# a_20069_7314# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2465 vdd a_25873_6693# a_25665_6693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2466 a_26624_103# a_26411_103# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2467 a_625_4057# a_412_4057# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2468 a_24573_3531# a_24668_3938# a_24623_3951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2469 vdd a_35487_3526# a_35279_3526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2470 a_24581_1748# a_24685_997# a_24636_1187# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2471 a_6110_4597# a_6915_4831# a_7074_5251# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2472 a_33587_1895# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2473 gnd d2 a_30099_5454# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2474 a_12345_5280# a_12132_5280# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2475 a_133_5215# a_622_5033# a_830_5033# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2476 vdd d4 a_24578_4482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2477 a_5436_1491# a_5917_1661# a_6125_1661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2478 a_11474_7982# a_11053_7982# a_10777_8164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2479 a_38244_7517# a_37823_7517# a_37555_7347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2480 a_19071_4144# a_20132_3773# a_20083_3963# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2481 gnd d1 a_24856_7855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2482 a_9426_3778# a_9422_3955# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2483 a_32780_2640# a_32567_2640# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2484 a_33572_4831# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2485 a_14802_3984# a_15059_3794# a_13790_4165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2486 a_37575_2835# a_37582_2451# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2487 a_22302_7530# a_21881_7530# a_21608_7746# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2488 a_1622_6812# a_1409_6812# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2489 gnd d4 a_3088_4511# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2490 a_41558_6870# a_41815_6680# a_40546_7051# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2491 a_32574_1661# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2492 a_17735_5259# a_17363_4839# a_16772_5020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2493 a_12303_2903# a_12090_2903# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2494 a_1416_5833# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2495 a_2906_6626# a_3120_5504# a_3071_5694# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2496 a_2140_4308# a_1719_4308# a_2041_4308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2497 a_32286_4813# a_32772_4597# a_32980_4597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2498 a_16786_1669# a_16365_1669# a_16092_1885# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2499 a_28683_1305# a_28628_2333# a_28812_4258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2500 a_40550_6874# a_41608_7095# a_41563_7108# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2501 a_12097_1924# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2502 gnd a_3348_1587# a_3140_1587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2503 a_7067_7330# a_6953_7211# a_7161_7211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2504 a_4126_6912# a_4383_6722# a_3114_7093# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2505 a_8427_1195# a_8684_1005# a_8372_1756# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2506 a_1813_1355# a_1441_935# a_849_701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2507 vdd a_35334_2498# a_35126_2498# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2508 a_22127_2068# a_21914_2068# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2509 a_12082_4860# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2510 a_40561_4115# a_41622_3744# a_41577_3757# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2511 gnd a_25874_7108# a_25666_7108# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2512 a_33982_199# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2513 a_40263_4659# a_40407_2477# a_40358_2667# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2514 vdd d0 a_36530_8097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2515 gnd a_24806_7435# a_24598_7435# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2516 a_130_6410# a_128_6196# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2517 vdd a_41823_6116# a_41615_6116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2518 a_23303_1326# a_22931_906# a_22340_1087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2519 a_11084_1690# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2520 a_9439_2233# a_9435_2410# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2521 a_17358_5820# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2522 a_32760_6557# a_32547_6557# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2523 a_35276_5916# a_35529_5903# a_35226_5496# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2524 a_409_5033# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2525 a_26921_2443# a_26919_2229# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2526 a_19060_6903# a_20118_7124# a_20073_7137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2527 vdd d2 a_3328_5504# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2528 a_38861_2853# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2529 a_32554_5578# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2530 vdd a_3398_2007# a_3190_2007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2531 a_24603_7868# a_25661_8089# a_25616_8102# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2532 a_27388_5964# a_27175_5964# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2533 a_6722_914# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2534 vdd d2 a_30099_5454# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2535 a_6705_3855# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2536 a_37848_2619# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2537 vdd a_13844_2527# a_13636_2527# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2538 a_9414_5912# a_9424_5169# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2539 a_35276_5916# a_36334_6137# a_36285_6327# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2540 a_5417_4218# a_5906_4036# a_6114_4036# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2541 a_19071_4144# a_20132_3773# a_20087_3786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2542 a_16359_3063# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2543 a_30922_3183# a_31175_3170# a_29909_2949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2544 a_16760_6980# a_17564_6799# a_17723_7219# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2545 a_10603_125# a_10182_125# a_10504_125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2546 a_25640_2789# a_25893_2776# a_24624_3147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2547 gnd d1 a_35534_4922# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2548 gnd a_24578_4482# a_24370_4482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2549 a_10182_125# d7 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2550 vdd d4 a_3088_4511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2551 vdd a_20337_4749# a_20129_4749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2552 a_20996_n19# a_31672_96# a_31994_96# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2553 a_17371_2882# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2554 gnd d3 a_24653_6407# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2555 a_32980_4597# a_32559_4597# a_32286_4813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2556 a_10811_2501# a_11290_2669# a_11498_2669# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2557 gnd d1 a_3378_5924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2558 a_3063_7477# a_3316_7464# a_2910_6449# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2559 a_24561_5665# a_24665_4914# a_24616_5104# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2560 a_26924_966# a_27413_1066# a_27621_1066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2561 a_1654_935# a_1441_935# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2562 a_25632_4746# a_25628_4923# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2563 a_38261_4576# a_37840_4576# a_37570_4411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2564 a_29892_6064# a_30953_5693# a_30904_5883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2565 a_32548_6972# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2566 gnd d0 a_15065_3228# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2567 gnd d1 a_30149_5874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2568 a_16058_8143# a_16058_7861# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2569 a_13787_5141# a_14848_4770# a_14799_4960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2570 a_36304_1995# a_36314_1252# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2571 a_6105_5578# a_5684_5578# a_5416_5408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2572 a_20095_2003# a_20352_1813# a_19083_2184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2573 gnd d1 a_14044_4951# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2574 vdd a_24806_7435# a_24598_7435# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2575 gnd a_31187_1210# a_30979_1210# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2576 vdd a_40823_2944# a_40615_2944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2577 a_33622_5251# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2578 a_23742_191# a_23321_191# a_23643_191# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2579 a_11490_4626# a_11069_4626# a_10796_4842# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2580 a_28924_170# a_28815_170# a_26733_103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2581 a_23321_191# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2582 a_38836_7751# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2583 a_23296_3405# a_22914_3847# a_22323_4028# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2584 a_22308_6964# a_21887_6964# a_21611_6864# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2585 a_17834_5259# a_17413_5259# a_17740_5378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2586 gnd a_35554_1005# a_35346_1005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2587 a_39473_4266# a_39076_2341# a_39344_1313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2588 a_16766_5586# a_16345_5586# a_16072_5802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2589 a_29701_2482# a_29899_3497# a_29854_3510# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2590 gnd a_36529_7682# a_36321_7682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2591 a_412_4057# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2592 a_22926_1887# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2593 a_23531_4279# a_23134_2354# a_23390_3286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2594 a_11089_709# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2595 a_21638_2250# a_22127_2068# a_22335_2068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2596 a_41590_2212# a_41843_2199# a_40577_1978# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2597 a_29850_3687# a_29954_2936# a_29905_3126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2598 a_22107_5985# a_21894_5985# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2599 a_22339_672# a_21918_672# a_21645_888# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2600 vdd a_24861_6874# a_24653_6874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2601 a_5431_2472# a_5429_2258# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2602 a_30918_3360# a_31175_3170# a_29909_2949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2603 a_28577_3384# a_28463_3265# a_28671_3265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2604 a_12132_5280# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2605 a_20087_3786# a_20083_3963# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2606 a_29850_3687# a_30107_3497# a_29701_2482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2607 a_12702_4316# a_12305_2391# a_12561_3323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2608 a_25636_2966# a_25893_2776# a_24624_3147# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2609 vdd a_24578_4482# a_24370_4482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2610 gnd a_24856_7855# a_24648_7855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2611 vdd d0 a_4391_6158# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2612 vdd a_36566_824# a_36358_824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2613 gnd d1 a_19333_2973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2614 a_27589_6943# a_27168_6943# a_26892_7125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2615 a_6118_2640# a_5697_2640# a_5424_2856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2616 a_33793_2874# a_33580_2874# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2617 a_128_5914# a_130_5815# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2618 a_33855_1334# a_33642_1334# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2619 a_38911_3273# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2620 a_3059_7654# a_3316_7464# a_2910_6449# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2621 gnd a_19340_1994# a_19132_1994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2622 a_39477_6258# a_39056_6258# a_39312_7190# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2623 a_12090_2903# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2624 a_12474_1363# a_12102_943# a_11510_709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2625 a_12102_943# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2626 a_32299_1976# a_32788_2076# a_32996_2076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2627 a_28552_7182# a_28180_6762# a_27589_6943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2628 a_37555_6752# a_38041_6536# a_38249_6536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2629 a_1637_3876# a_1424_3876# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2630 a_19051_8061# a_20112_7690# a_20067_7703# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2631 a_28663_5222# a_28242_5222# a_28564_5222# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2632 a_33001_1095# a_32580_1095# a_32304_995# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2633 a_13787_5141# a_14848_4770# a_14803_4783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2634 gnd a_9685_3199# a_9477_3199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2635 a_22120_3047# a_21907_3047# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2636 a_23534_191# a_23321_191# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2637 gnd a_8617_3526# a_8409_3526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2638 vdd a_31187_1210# a_30979_1210# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2639 a_33937_7330# a_33555_7772# a_32963_7538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2640 a_4158_2254# a_4154_2431# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2641 a_16060_7762# a_16546_7546# a_16754_7546# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2642 a_37553_6851# a_37555_6752# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2643 a_27167_6528# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2644 a_27396_4007# a_27183_4007# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2645 a_35269_6895# a_35522_6882# a_35210_7633# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2646 a_28815_170# a_28602_170# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2647 a_10791_6418# a_11270_6586# a_11478_6586# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2648 a_37560_6154# a_38049_5972# a_38257_5972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2649 a_12365_1363# a_12152_1363# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2650 a_27381_6943# a_27168_6943# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2651 a_26904_4883# a_27393_4983# a_27601_4983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2652 a_17579_3863# a_17366_3863# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2653 a_3113_7897# a_3366_7884# a_3063_7477# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2654 a_40545_7855# a_41603_8076# a_41554_8266# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2655 vdd a_36529_7682# a_36321_7682# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2656 vdd a_3328_5504# a_3120_5504# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2657 a_27175_5964# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2658 a_20075_5920# a_20085_5177# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2659 a_621_4618# a_408_4618# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2660 a_8419_2978# a_9477_3199# a_9432_3212# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2661 a_24640_1010# a_25698_1231# a_25649_1421# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2662 a_35230_3716# a_35334_2965# a_35289_2978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2663 a_27600_4568# a_28405_4802# a_28564_5222# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2664 a_16787_2084# a_16366_2084# a_16090_1984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2665 a_37841_4991# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2666 a_22340_1087# a_21919_1087# a_21643_1269# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2667 a_26926_1462# a_27407_1632# a_27615_1632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2668 a_13744_3568# a_13997_3555# a_13591_2540# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2669 a_7099_1453# a_6717_1895# a_6125_1661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2670 a_3113_7897# a_4171_8118# a_4122_8308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2671 gnd d2 a_35479_5483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2672 gnd d3 a_8464_2498# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2673 a_37555_6752# a_37562_6368# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2674 a_6965_5251# a_6752_5251# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2675 a_4146_2995# a_4403_2805# a_3134_3176# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2676 a_19055_7884# a_19308_7871# a_19005_7464# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2677 gnd a_35534_4922# a_35326_4922# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2678 a_10802_3266# a_10802_2984# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2679 a_19055_7884# a_20113_8105# a_20064_8295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2680 a_22906_5804# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2681 a_24396_6597# a_24610_5475# a_24561_5665# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2682 a_26909_3808# a_26914_3422# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2683 a_17596_922# a_17383_922# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2684 gnd a_3378_5924# a_3170_5924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2685 gnd d2 a_40760_5462# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2686 a_32289_3837# a_32294_3451# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2687 a_41570_6129# a_41823_6116# a_40557_5895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2688 gnd a_20341_4188# a_20133_4188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2689 a_31994_96# a_31885_96# a_20996_n19# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2690 a_30898_7277# a_31155_7087# a_29889_6866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2691 a_25616_6883# a_25873_6693# a_24604_7064# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2692 a_13567_6634# a_13781_5512# a_13732_5702# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2693 vdd a_8617_3526# a_8409_3526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2694 gnd a_15065_3228# a_14857_3228# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2695 a_22119_2632# a_21906_2632# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2696 a_11486_6022# a_12290_5841# a_12459_5399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2697 a_12498_6308# a_12285_6308# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2698 gnd a_14044_4951# a_13836_4951# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2699 a_36296_3778# a_36292_3955# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2700 vdd d0 a_36567_1239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2701 a_5429_1976# a_5431_1877# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2702 a_605_7974# a_392_7974# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2703 a_33773_6791# a_33560_6791# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2704 gnd a_25889_4172# a_25681_4172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2705 a_21907_3047# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2706 a_38036_7517# a_37823_7517# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2707 a_8340_7633# a_8444_6882# a_8399_6895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2708 gnd a_19320_5911# a_19112_5911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2709 a_32775_3621# a_32562_3621# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2710 a_20100_1022# a_16104_703# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2711 a_33567_5812# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2712 a_34291_4287# a_33870_4287# a_34196_6279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2713 a_40545_7855# a_41603_8076# gnd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2714 a_39054_6770# a_38841_6770# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2715 a_20080_6158# a_20333_6145# a_19067_5924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2716 a_32279_5893# a_32768_5993# a_32976_5993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2717 a_1617_7793# a_1404_7793# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2718 a_24640_1010# a_25698_1231# a_25653_1244# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2719 a_32299_2258# a_32299_1976# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2720 a_32981_5012# a_32560_5012# a_32284_4912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2721 a_10802_3266# a_11291_3084# a_11499_3084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2722 gnd a_9665_7116# a_9457_7116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2723 a_26906_4784# a_26909_4403# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2724 a_1781_7232# a_1672_7232# a_1880_7232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2725 gnd a_8667_3946# a_8459_3946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2726 a_26907_4189# a_27396_4007# a_27604_4007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2727 a_1932_4308# a_1719_4308# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2728 a_13740_3745# a_13997_3555# a_13591_2540# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2729 a_22099_6549# a_21886_6549# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2730 vdd d2 a_35479_5483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2731 vdd d0 a_15059_3794# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2732 vdd d0 a_15077_1268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2733 a_16584_1103# a_16371_1103# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2734 gnd d3 a_13844_2527# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2735 a_7094_1334# a_6985_1334# a_7193_1334# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2736 a_32568_3055# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2737 a_16546_7546# a_16333_7546# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2738 a_16775_4044# a_17579_3863# a_17748_3421# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2739 a_141_2976# a_630_3076# a_838_3076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2740 a_34051_3294# a_33630_3294# a_33957_3413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2741 a_36309_2233# a_36305_2410# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2742 a_5431_1877# a_5436_1491# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2743 a_12077_5841# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2744 a_25628_6142# a_25624_6319# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2745 gnd a_19333_2973# a_19125_2973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2746 a_24396_6597# a_24610_5475# a_24565_5488# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2747 a_25621_7121# a_25874_7108# a_24608_6887# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2748 a_11491_5041# a_11070_5041# a_10794_4941# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2749 a_8407_5112# a_8664_4922# a_8352_5673# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2750 a_33580_2874# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2751 a_24553_7448# a_24806_7435# a_24400_6420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2752 a_41566_6306# a_41823_6116# a_40557_5895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2753 vdd d2 a_40760_5462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2754 a_39225_5230# a_38853_4810# a_38261_4576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2755 a_4146_4214# a_4399_4201# a_3133_3980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2756 a_1692_3315# a_1479_3315# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2757 a_37587_875# a_38073_659# a_38281_659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2758 a_16767_6001# a_16346_6001# a_16070_5901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2759 gnd d0 a_20337_4749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2760 a_38856_3834# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2761 a_38276_1640# a_37855_1640# a_37587_1470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2762 a_13567_6634# a_13781_5512# a_13736_5525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2763 a_37568_3915# a_38057_4015# a_38265_4015# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2764 a_9412_7129# a_9408_7306# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2765 a_1424_3876# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2766 a_7079_5370# a_6697_5812# a_6105_5578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2767 gnd d3 a_8444_6415# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2768 a_27595_5549# a_27174_5549# a_26906_5379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2769 a_30893_8258# a_30896_7666# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2770 a_20100_2241# a_20096_2418# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2771 a_13587_2717# a_13844_2527# a_13492_4709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2772 a_36277_8110# a_36273_8287# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2773 a_29834_7427# a_30087_7414# a_29681_6399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2774 a_6905_6279# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2775 gnd d1 a_35529_5903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2776 a_830_5033# a_409_5033# a_133_5215# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2777 a_22319_4589# a_21898_4589# a_21625_4805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2778 a_25652_829# a_25648_1006# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2779 a_9443_837# a_9439_1014# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2780 vdd a_25889_4172# a_25681_4172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2781 a_27183_4007# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2782 a_27620_651# a_27199_651# a_26926_867# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2783 vdd d1 a_8679_1986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2784 gnd a_19030_4498# a_18822_4498# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2785 a_16754_7546# a_17559_7780# a_17728_7338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2786 a_29909_2949# a_30967_3170# a_30918_3360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2787 a_12152_1363# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2788 a_20076_6335# a_20333_6145# a_19067_5924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2789 a_5397_8135# a_5886_7953# a_6094_7953# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2790 a_24565_5488# a_24660_5895# a_24611_6085# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2791 a_12814_228# a_13541_4519# a_13496_4532# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2792 a_17366_3863# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2793 vref a_116_8156# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2794 gnd a_41830_3744# a_41622_3744# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2795 a_38282_1074# a_39086_893# a_39245_1313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2796 a_9438_1818# a_9434_1995# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2797 vdd a_9665_7116# a_9457_7116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2798 gnd d0 a_15060_4209# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2799 a_6119_3055# a_5698_3055# a_5422_2955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2800 a_155_917# a_162_716# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2801 a_16780_3063# a_16359_3063# a_16083_2963# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2802 a_21918_672# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2803 a_5134_132# a_4921_132# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2804 a_5678_6972# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2805 a_9408_7306# a_9411_6714# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2806 a_38256_5557# a_37835_5557# a_37562_5773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2807 a_7161_7211# a_6740_7211# a_7067_7330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2808 a_7082_3294# a_6710_2874# a_6118_2640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2809 gnd a_31182_2191# a_30974_2191# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2810 vdd d0 a_4410_1826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2811 a_5409_6175# a_5409_5893# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2812 gnd a_8464_2498# a_8256_2498# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2813 a_36273_8287# a_36276_7695# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2814 a_33823_7211# a_33610_7211# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2815 a_23531_4279# a_23422_4279# a_23630_4279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2816 a_6752_5251# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2817 a_5897_5578# a_5684_5578# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2818 a_34192_4287# a_33795_2362# a_34051_3294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2819 a_24549_7625# a_24806_7435# a_24400_6420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2820 a_39104_7190# a_38891_7190# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2821 a_11493_3650# a_12298_3884# a_12467_3442# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2822 a_40566_3134# a_40823_2944# a_40511_3695# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2823 a_10782_7183# a_11271_7001# a_11479_7001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2824 vdd d0 a_25886_5148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2825 a_21901_3613# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2826 a_32294_2856# a_32780_2640# a_32988_2640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2827 vdd d0 a_31162_6108# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2828 a_8414_3959# a_9472_4180# a_9423_4370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2829 vdd d3 a_8444_6415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2830 a_21613_6765# a_22099_6549# a_22307_6549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2831 a_16095_1285# a_16584_1103# a_16792_1103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2832 a_16760_6980# a_16339_6980# a_16063_7162# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2833 a_24631_2168# a_25692_1797# a_25647_1810# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2834 gnd d2 a_8597_7443# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2835 a_19083_2184# a_20144_1813# a_20095_2003# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2836 a_29830_7604# a_30087_7414# a_29681_6399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2837 a_10799_3866# a_11285_3650# a_11493_3650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2838 a_8112_4680# a_8256_2498# a_8211_2511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2839 a_121_6893# a_610_6993# a_818_6993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2840 a_12285_6308# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2841 vdd a_36567_1239# a_36359_1239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2842 a_29909_2949# a_30967_3170# a_30922_3183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2843 a_392_7974# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2844 a_33560_6791# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2845 a_3125_5937# a_4183_6158# a_4138_6171# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2846 a_21618_6167# a_22107_5985# a_22315_5985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2847 vdd a_20321_8105# a_20113_8105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2848 vdd a_41830_3744# a_41622_3744# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2849 a_24603_7868# a_24856_7855# a_24553_7448# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2850 a_37823_7517# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2851 vdd d0 a_9672_6137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2852 a_32562_3621# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2853 a_39324_5230# a_38903_5230# a_39225_5230# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2854 a_143_3472# a_624_3642# a_832_3642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2855 vdd d1 a_35537_3946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2856 a_41594_816# a_41847_803# a_40578_1174# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2857 a_17799_2370# a_17586_2370# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2858 a_1404_7793# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2859 a_21881_7530# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2860 a_20072_6722# a_20325_6709# a_19056_7080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2861 a_32281_6389# a_32760_6557# a_32968_6557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2862 a_9439_2233# a_9692_2220# a_8426_1999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2863 a_23382_5243# a_22961_5243# a_23288_5362# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2864 a_33000_680# a_32579_680# a_32306_896# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2865 a_11058_7001# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2866 vdd a_25869_8089# a_25661_8089# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2867 a_16075_4920# a_16564_5020# a_16772_5020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2868 gnd d2 a_40780_1545# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2869 a_28589_1424# a_28207_1866# a_27615_1632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2870 a_32996_2076# a_32575_2076# a_32299_2258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2871 a_20068_8118# a_21606_8127# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2872 a_21643_987# a_21645_888# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2873 a_15795_140# a_15582_140# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2874 a_16371_1103# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2875 vdd a_15077_1268# a_14869_1268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2876 a_10784_7397# a_11265_7567# a_11473_7567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2877 gnd a_13844_2527# a_13636_2527# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2878 a_28911_4258# a_28490_4258# a_28816_6250# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2879 a_16333_7546# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2880 a_26899_5864# a_27388_5964# a_27596_5964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2881 a_11277_5607# a_11064_5607# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2882 vdd d1 a_14047_3975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2883 a_26926_867# a_26933_666# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2884 gnd d0 a_15040_8126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2885 a_32269_7754# a_32274_7368# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2886 a_429_1116# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2887 a_4131_7150# a_4127_7327# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2888 a_8414_3959# a_9472_4180# a_9427_4193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2889 a_35297_1195# a_36358_824# a_36313_837# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2890 gnd a_20337_4749# a_20129_4749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2891 a_116_7874# a_118_7775# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2892 gnd d2 a_24818_5475# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2893 vdd a_30169_1957# a_29961_1957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2894 vdd d2 a_8597_7443# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2895 a_16759_6565# a_16338_6565# a_16072_6397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2896 a_41557_7674# a_41553_7851# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2897 gnd d0 a_31154_6672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2898 a_616_5599# a_403_5599# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2899 a_6113_3621# a_5692_3621# a_5424_3451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2900 a_39250_1432# a_38868_1874# a_38277_2055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2901 gnd a_8444_6415# a_8236_6415# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2902 a_28671_3265# a_28250_3265# a_28577_3384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2903 a_40491_7612# a_40595_6861# a_40546_7051# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2904 gnd a_31161_5693# a_30953_5693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2905 a_1684_5272# a_1471_5272# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2906 vdd a_25905_816# a_25697_816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2907 a_26914_2827# a_26921_2443# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2908 a_35057_6605# a_35271_5483# a_35222_5673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2909 gnd a_25885_4733# a_25677_4733# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2910 a_4122_8308# a_4379_8118# a_3113_7897# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2911 a_29830_7604# a_29934_6853# a_29889_6866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2912 a_17842_3302# a_17421_3302# a_17748_3421# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2913 a_11290_2669# a_11077_2669# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2914 a_23112_6783# a_22899_6783# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2915 a_14798_5764# a_14794_5941# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2916 a_16566_3629# a_16353_3629# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2917 a_27413_1066# a_27200_1066# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2918 a_8372_1756# a_8476_1005# a_8427_1195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2919 a_9435_2410# a_9692_2220# a_8426_1999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2920 a_30893_8258# a_31150_8068# a_29884_7847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2921 a_4127_7327# a_4130_6735# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2922 gnd d0 a_9664_6701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2923 a_1837_6300# a_1624_6300# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2924 a_32756_7953# a_32543_7953# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2925 a_28388_7743# a_28175_7743# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2926 a_23271_7203# a_23162_7203# a_23370_7203# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2927 a_24400_6420# a_24653_6407# a_24325_4495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2928 a_22328_3047# a_23132_2866# a_23291_3286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2929 gnd d1 a_8647_7863# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2930 vdd d2 a_40780_1545# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2931 a_41570_6129# a_41566_6306# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2932 a_16077_4821# a_16563_4605# a_16771_4605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2933 a_34304_199# a_35031_4490# a_34982_4680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2934 a_6093_7538# a_5672_7538# a_5399_7754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2935 a_5411_5794# a_5416_5408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2936 a_28584_1305# a_28475_1305# a_28683_1305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2937 a_13587_2717# a_13801_1595# a_13756_1608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2938 a_29889_6866# a_30947_7087# a_30902_7100# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2939 a_5890_6557# a_5677_6557# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2940 a_23308_1445# a_22926_1887# a_22335_2068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2941 a_33610_7211# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2942 vdd d1 a_40835_984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2943 vdd d0 a_15040_8126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2944 gnd d2 a_19278_3534# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2945 a_5684_5578# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2946 a_38074_1074# a_37861_1074# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2947 a_850_1116# a_429_1116# a_153_1298# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2948 a_812_7559# a_391_7559# a_123_7389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2949 gnd d0 a_4391_6158# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2950 a_25636_4185# a_25889_4172# a_24623_3951# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2951 a_4142_4775# a_4395_4762# a_3126_5133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2952 a_29901_4906# a_30154_4893# a_29842_5644# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2953 a_23283_5243# a_22911_4823# a_22319_4589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2954 vdd d2 a_24818_5475# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2955 a_32988_2640# a_33793_2874# a_33952_3294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2956 vdd d0 a_31154_6672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2957 vdd a_31162_6108# a_30954_6108# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2958 a_22914_3847# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2959 a_22334_1653# a_21913_1653# a_21645_1483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2960 a_3145_2020# a_4203_2241# a_4154_2431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2961 a_21887_6964# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2962 a_32976_5993# a_32555_5993# a_32279_6175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2963 a_21626_3928# a_22115_4028# a_22323_4028# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2964 a_37587_1470# a_37585_1256# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2965 a_40573_2155# a_41634_1784# a_41585_1974# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2966 vdd a_8444_6415# a_8236_6415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2967 a_41594_816# a_41590_993# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2968 gnd d1 a_40830_1965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2969 gnd d0 a_9692_2220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2970 a_1644_2383# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2971 a_39364_4266# a_39151_4266# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2972 a_26892_7125# a_26892_6843# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2973 a_32286_5408# a_32284_5194# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2974 a_21606_7845# a_21608_7746# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2975 a_32272_7154# a_32272_6872# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2976 a_35057_6605# a_35271_5483# a_35226_5496# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2977 vdd a_25885_4733# a_25677_4733# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2978 a_13756_1608# a_13851_2015# a_13802_2205# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2979 vdd d1 a_14027_7892# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2980 a_33805_914# a_33592_914# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2981 a_637_2097# a_424_2097# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2982 a_35214_7456# a_35467_7443# a_35061_6428# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2983 a_8394_7876# a_9452_8097# a_9407_8110# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2984 a_11302_709# a_11089_709# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2985 a_26887_8106# a_27376_7924# a_27584_7924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2986 a_1649_1916# a_1436_1916# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2987 a_27609_3026# a_27188_3026# a_26912_2926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2988 a_41583_3191# a_41579_3368# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2989 a_12593_4316# a_12380_4316# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2990 vdd a_35537_3946# a_35329_3946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2991 a_22131_672# a_21918_672# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2992 a_10814_1306# a_10814_1024# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2993 a_17586_2370# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2994 a_11486_6022# a_11065_6022# a_10789_6204# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2995 gnd d1 a_24868_5895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2996 a_39230_5349# a_38848_5791# a_38257_5972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2997 a_5697_2640# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2998 a_28651_7182# a_28230_7182# a_28557_7301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2999 a_9431_2797# a_9684_2784# a_8415_3155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3000 a_28572_3265# a_28200_2845# a_27608_2611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3001 gnd a_41811_8076# a_41603_8076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3002 a_22314_5570# a_21893_5570# a_21620_5786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3003 gnd a_8369_4490# a_8161_4490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3004 a_1634_4852# a_1421_4852# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3005 vdd d0 a_31182_2191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3006 a_25636_4185# a_25632_4362# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3007 a_12315_943# a_12102_943# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3008 vdd d2 a_19278_3534# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3009 a_14824_1281# a_14820_1458# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3010 a_17614_7219# a_17401_7219# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3011 a_12353_3323# a_12140_3323# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3012 a_11064_5607# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3013 a_8352_5673# a_8456_4922# a_8407_5112# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3014 a_25632_4362# a_25889_4172# a_24623_3951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3015 a_19037_1587# a_19290_1574# a_18868_2696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3016 a_17346_7780# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3017 vdd a_14047_3975# a_13839_3975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3018 a_14787_8139# a_16058_8143# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3019 a_22094_7530# a_21881_7530# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3020 a_4138_4952# a_4395_4762# a_3126_5133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3021 a_36308_1818# a_36304_1995# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3022 a_35242_1756# a_35346_1005# a_35301_1018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3023 a_41579_3368# a_41582_2776# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3024 a_3145_2020# a_4203_2241# a_4158_2254# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3025 a_34403_199# a_37285_111# a_31994_96# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3026 a_40573_2155# a_41634_1784# a_41589_1797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3027 vdd d0 a_9692_2220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3028 a_39233_3273# a_38861_2853# a_38270_3034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3029 vdd d0 a_36542_6137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3030 gnd a_24818_5475# a_24610_5475# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3031 gnd a_31154_6672# a_30946_6672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3032 a_403_5599# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3033 a_16775_4044# a_16354_4044# a_16078_4226# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3034 a_13756_1608# a_13851_2015# a_13806_2028# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3035 a_7087_3413# a_6705_3855# a_6114_4036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3036 a_6953_7211# a_6740_7211# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3037 a_35210_7633# a_35467_7443# a_35061_6428# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3038 a_6099_6972# a_5678_6972# a_5402_6872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3039 gnd a_13989_5512# a_13781_5512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3040 a_1471_5272# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3041 gnd a_40768_3505# a_40560_3505# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3042 a_6923_2874# a_6710_2874# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3043 a_37585_1256# a_38074_1074# a_38282_1074# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3044 a_16760_6980# a_16339_6980# a_16063_6880# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3045 a_24615_5908# a_25673_6129# a_25628_6142# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3046 a_38054_4991# a_37841_4991# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3047 a_14820_1458# a_14823_866# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3048 vdd a_8647_7863# a_8439_7863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3049 a_29904_3930# a_30157_3917# a_29854_3510# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3050 a_38245_7932# a_39049_7751# a_39218_7309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3051 a_18095_207# a_17986_207# a_15904_140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3052 a_6717_1895# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3053 a_5429_2258# a_5918_2076# a_6126_2076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3054 a_32968_6557# a_33773_6791# a_33932_7211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3055 vdd d1 a_40815_4901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3056 gnd d0 a_36567_1239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3057 a_16353_3629# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3058 a_27200_1066# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3059 a_34008_2362# a_33795_2362# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3060 a_1624_6300# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3061 a_9427_2974# a_9684_2784# a_8415_3155# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3062 vdd a_41811_8076# a_41603_8076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3063 a_28175_7743# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3064 a_26733_103# a_26624_103# a_26832_103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3065 a_32988_2640# a_32567_2640# a_32301_2472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3066 a_116_7874# a_605_7974# a_813_7974# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3067 a_39086_893# a_38873_893# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3068 a_16090_1984# a_16579_2084# a_16787_2084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3069 a_11473_7567# a_12278_7801# a_12447_7359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3070 a_40507_5475# a_40760_5462# a_40338_6584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3071 a_617_6014# a_404_6014# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3072 a_18852_6436# a_19050_7451# a_19001_7641# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3073 a_9424_5169# a_9420_5346# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3074 a_3075_5517# a_3328_5504# a_2906_6626# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3075 a_2045_6300# a_1932_4308# a_2140_4308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3076 vdd a_9697_1239# a_9489_1239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3077 a_19033_1764# a_19290_1574# a_18868_2696# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3078 vdd d1 a_3391_2986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3079 gnd d0 a_15077_1268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3080 a_40511_3695# a_40615_2944# a_40566_3134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3081 a_32542_7538# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3082 gnd a_19278_3534# a_19070_3534# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3083 a_19063_6101# a_20124_5730# a_20075_5920# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3084 a_4146_4214# a_4142_4391# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3085 vdd a_24818_5475# a_24610_5475# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3086 vdd a_31154_6672# a_30946_6672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3087 a_33870_4287# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3088 a_32968_6557# a_32547_6557# a_32274_6773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3089 vdd a_35239_4490# a_35031_4490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3090 a_1806_3434# a_1692_3315# a_1900_3315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3091 gnd d0 a_9684_2784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3092 gnd d0 a_36534_6701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3093 vdd a_13989_5512# a_13781_5512# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3094 a_39151_4266# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3095 a_630_3076# a_417_3076# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3096 a_24569_3708# a_24673_2957# a_24628_2970# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3097 a_9420_5346# a_9423_4754# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3098 a_12303_2903# a_12090_2903# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3099 gnd a_31186_795# a_30978_795# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3100 a_25612_8279# a_25869_8089# a_24603_7868# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3101 a_837_2661# a_416_2661# a_143_2877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3102 a_7421_4287# a_7325_199# a_5243_132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3103 vdd a_14027_7892# a_13819_7892# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3104 a_20084_4378# a_20341_4188# a_19075_3967# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3105 a_33592_914# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3106 a_424_2097# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3107 gnd d0 a_4378_7703# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3108 a_29854_3510# a_29949_3917# a_29904_3930# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3109 a_12097_1924# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3110 a_36285_6327# a_36288_5735# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3111 a_1642_2895# a_1429_2895# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3112 a_29862_1727# a_29966_976# a_29917_1166# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3113 a_13591_2540# a_13844_2527# a_13492_4709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3114 a_24604_7064# a_25665_6693# a_25616_6883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3115 a_37570_4411# a_37568_4197# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3116 a_21628_3829# a_21633_3443# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3117 gnd d1 a_24861_6874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3118 a_40553_6072# a_41614_5701# a_41569_5714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3119 a_29862_1727# a_30119_1537# a_29697_2659# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3120 a_12380_4316# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3121 a_1436_1916# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3122 a_4142_4391# a_4145_3799# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3123 a_6131_1095# a_5710_1095# a_5434_1277# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3124 a_14807_3003# a_15064_2813# a_13795_3184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3125 a_39332_3273# a_38911_3273# a_39238_3392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3126 gnd a_24868_5895# a_24660_5895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3127 a_12814_228# a_13541_4519# a_13492_4709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3128 a_10804_3480# a_10802_3266# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3129 a_40503_5652# a_40760_5462# a_40338_6584# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3130 a_38853_4810# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3131 a_5443_695# a_5922_680# a_6130_680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3132 a_27583_7509# a_27162_7509# a_26889_7725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3133 a_18852_6436# a_19050_7451# a_19005_7464# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3134 gnd a_40748_7422# a_40540_7422# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3135 a_1421_4852# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3136 a_37855_1640# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3137 a_128_6196# a_128_5914# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3138 a_5905_3621# a_5692_3621# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3139 a_17584_2882# a_17371_2882# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3140 a_2252_220# a_1831_220# a_2140_4308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3141 a_12102_943# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3142 vdd a_40615_2477# a_40407_2477# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3143 a_6697_5812# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3144 a_8187_6605# a_8401_5483# a_8352_5673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3145 a_37567_4792# a_38053_4576# a_38261_4576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3146 a_12283_6820# a_12070_6820# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3147 vdd a_19278_3534# a_19070_3534# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3148 a_38281_659# a_37860_659# a_37594_674# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3149 a_17401_7219# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3150 a_19063_6101# a_20124_5730# a_20079_5743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3151 gnd d0 a_31186_795# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3152 a_17378_1903# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3153 vdd d0 a_20345_2792# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3154 a_33932_7211# a_33823_7211# a_34031_7211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3155 a_21898_4589# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3156 a_11285_3650# a_11072_3650# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3157 gnd a_8629_1566# a_8421_1566# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3158 a_21638_2250# a_21638_1968# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3159 a_25632_4746# a_25885_4733# a_24616_5104# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3160 a_36302_3212# a_36555_3199# a_35289_2978# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3161 a_9407_6891# a_9664_6701# a_8395_7072# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3162 a_40263_4659# a_40520_4469# a_39585_178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3163 a_27408_2047# a_27195_2047# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3164 vdd a_3183_2519# a_2975_2519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3165 a_23107_7764# a_22894_7764# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3166 a_16072_5802# a_16558_5586# a_16766_5586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3167 a_27179_4568# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3168 a_2044_220# a_1831_220# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3169 vdd a_36542_6137# a_36334_6137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3170 gnd d0 a_25886_5148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3171 a_10799_4461# a_11282_4626# a_11490_4626# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3172 a_155_917# a_641_701# a_849_701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3173 a_5243_132# a_7112_199# a_7421_4287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3174 a_29884_7847# a_30942_8068# a_30897_8081# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3175 a_5698_3055# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3176 vdd d0 a_9684_2784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3177 a_7112_199# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3178 a_28420_1866# a_28207_1866# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3179 gnd d1 a_24888_1978# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3180 a_27393_4983# a_27180_4983# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3181 a_23422_4279# a_23209_4279# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3182 a_19013_5681# a_19270_5491# a_18848_6613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3183 a_32301_2472# a_32299_2258# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3184 a_6710_2874# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3185 a_8431_1018# a_9489_1239# a_9444_1252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3186 a_12561_3323# a_12518_2391# a_12702_4316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3187 a_5885_7538# a_5672_7538# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3188 gnd d0 a_25900_1797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3189 a_32548_6972# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3190 a_35246_1579# a_35341_1986# a_35292_2176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3191 vdd d0 a_41847_803# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3192 a_11505_1690# a_11084_1690# a_10811_1906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3193 vdd a_40815_4901# a_40607_4901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3194 gnd a_36567_1239# a_36359_1239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3195 a_3125_5937# a_4183_6158# a_4134_6348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3196 a_141_3258# a_141_2976# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3197 a_23182_3286# a_22969_3286# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3198 a_33795_2362# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3199 a_16551_6565# a_16338_6565# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3200 gnd d0 a_9672_6137# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3201 a_23288_5362# a_22906_5804# a_22315_5985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3202 vdd a_40748_7422# a_40540_7422# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3203 a_20085_5177# a_20081_5354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3204 a_18773_4688# a_19030_4498# a_18095_207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3205 a_25616_8102# a_25612_8279# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3206 gnd d0 a_20346_3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3207 a_4157_1839# a_4410_1826# a_3141_2197# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3208 a_16092_2480# a_16571_2648# a_16779_2648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3209 a_404_6014# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3210 a_8187_6605# a_8401_5483# a_8356_5496# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3211 a_609_6578# a_396_6578# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3212 a_41569_5714# a_41565_5891# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3213 a_27588_6528# a_28393_6762# a_28552_7182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3214 a_30910_5317# a_31167_5127# a_29901_4906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3215 vdd a_8629_1566# a_8421_1566# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3216 a_6110_4597# a_5689_4597# a_5419_4432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3217 a_25628_4923# a_25885_4733# a_24616_5104# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3218 gnd a_15077_1268# a_14869_1268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3219 a_37829_6951# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3220 a_22328_3047# a_21907_3047# a_21631_3229# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3221 a_5434_995# a_5436_896# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3222 a_37568_3915# a_37570_3816# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3223 vdd d0 a_41843_2199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3224 gnd d1 a_19325_4930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3225 vdd d0 a_36561_1805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3226 a_21919_1087# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3227 a_23291_3286# a_22919_2866# a_22328_3047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3228 a_38903_5230# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3229 a_33785_4831# a_33572_4831# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3230 a_833_4057# a_1637_3876# a_1806_3434# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3231 a_23402_1326# a_22981_1326# a_23303_1326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3232 a_20081_5354# a_20084_4762# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3233 a_16771_4605# a_16350_4605# a_16077_4821# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3234 a_4141_3976# a_4151_3233# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3235 a_38048_5557# a_37835_5557# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3236 a_28577_3384# a_28195_3826# a_27604_4007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3237 a_32787_1661# a_32574_1661# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3238 a_25612_8279# a_25615_7687# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3239 a_10802_2984# a_10804_2885# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3240 a_27589_6943# a_27168_6943# a_26892_6843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3241 gnd a_36534_6701# a_36326_6701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3242 a_1629_5833# a_1416_5833# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3243 a_22961_5243# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3244 vdd a_3386_3967# a_3178_3967# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3245 a_8356_5496# a_8451_5903# a_8402_6093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3246 a_7322_4287# a_6925_2362# a_7193_1334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3247 a_12090_2903# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3248 a_12333_7240# a_12120_7240# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3249 gnd a_9677_5156# a_9469_5156# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3250 a_22112_5004# a_21899_5004# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3251 a_829_4618# a_408_4618# a_138_4453# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3252 a_13571_6457# a_13769_7472# a_13720_7662# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3253 a_36282_7129# a_36535_7116# a_35269_6895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3254 a_33805_914# a_33592_914# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3255 a_26919_2229# a_27408_2047# a_27616_2047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3256 gnd a_4378_7703# a_4170_7703# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3257 a_22303_7945# a_23107_7764# a_23276_7322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3258 gnd a_8679_1986# a_8471_1986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3259 a_35284_3959# a_35537_3946# a_35234_3539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3260 a_21643_987# a_22132_1087# a_22340_1087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3261 vdd d0 a_15071_1834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3262 a_5411_6389# a_5409_6175# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3263 a_4126_8131# a_4379_8118# a_3113_7897# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3264 a_34063_1334# a_33642_1334# a_33969_1453# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3265 a_28400_5783# a_28187_5783# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3266 a_16104_703# a_16583_688# a_16791_688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3267 a_22340_1087# a_23144_906# a_23303_1326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3268 a_30897_8081# a_31150_8068# a_29884_7847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3269 a_10804_2885# a_10811_2501# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3270 a_24565_5488# a_24818_5475# a_24396_6597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3271 a_35222_5673# a_35326_4922# a_35281_4935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3272 a_14792_7158# a_15045_7145# a_13779_6924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3273 gnd d0 a_25880_5714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3274 a_17371_2882# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3275 a_37585_1256# a_37585_974# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3276 a_1704_1355# a_1491_1355# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3277 a_5692_3621# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3278 a_38868_1874# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3279 a_7326_6279# a_6905_6279# a_7161_7211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3280 vdd d1 a_40810_5882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3281 a_6918_3855# a_6705_3855# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3282 a_13794_3988# a_14047_3975# a_13744_3568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3283 a_32299_1976# a_32301_1877# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3284 a_37580_1955# a_38069_2055# a_38277_2055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3285 a_32963_7538# a_33768_7772# a_33937_7330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3286 a_12070_6820# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3287 vdd a_14009_1595# a_13801_1595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3288 a_5404_6773# a_5890_6557# a_6098_6557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3289 a_33932_7211# a_33560_6791# a_32968_6557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3290 a_13736_5525# a_13989_5512# a_13567_6634# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3291 vdd a_20345_2792# a_20137_2792# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3292 a_13736_5525# a_13831_5932# a_13786_5945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3293 a_11072_3650# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3294 vdd d2 a_24826_3518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3295 a_27401_3026# a_27188_3026# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3296 a_23162_7203# a_22949_7203# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3297 a_29846_5467# a_30099_5454# a_29677_6576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3298 gnd d0 a_4398_3786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3299 a_37565_5173# a_38054_4991# a_38262_4991# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3300 a_27195_2047# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3301 a_1786_7351# a_1404_7793# a_812_7559# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3302 vdd d1 a_30162_2936# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3303 gnd d0 a_20326_7124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3304 a_32776_4036# a_32563_4036# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3305 a_29900_4107# a_30961_3736# a_30912_3926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3306 gnd d0 a_41835_2763# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3307 gnd d1 a_24881_2957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3308 a_3118_6916# a_3371_6903# a_3059_7654# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3309 a_5409_6175# a_5898_5993# a_6106_5993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3310 a_34192_4287# a_34083_4287# a_34291_4287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3311 a_37285_111# a_37072_111# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3312 vdd a_9677_5156# a_9469_5156# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3313 a_27180_4983# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3314 a_8394_7876# a_8647_7863# a_8344_7456# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3315 a_9435_2410# a_9438_1818# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3316 a_13571_6457# a_13769_7472# a_13724_7485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3317 a_36278_7306# a_36535_7116# a_35269_6895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3318 gnd d0 a_20340_3773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3319 a_32301_1877# a_32306_1491# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3320 a_5672_7538# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3321 a_3079_3737# a_3183_2986# a_3138_2999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3322 gnd a_14059_2015# a_13851_2015# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3323 a_7173_5251# a_6752_5251# a_7079_5370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3324 a_17728_7338# a_17346_7780# a_16754_7546# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3325 a_22926_1887# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3326 a_23271_7203# a_22899_6783# a_22308_6964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3327 a_41558_6870# a_41570_6129# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3328 a_21899_5004# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3329 a_19060_6903# a_19313_6890# a_19001_7641# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3330 a_11286_4065# a_11073_4065# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3331 a_8364_3539# a_8459_3946# a_8414_3959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3332 a_30896_7666# a_30892_7843# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3333 a_33835_5251# a_33622_5251# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3334 a_22322_3613# a_21901_3613# a_21628_3829# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3335 a_39069_3834# a_38856_3834# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3336 a_33952_3294# a_33843_3294# a_34051_3294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3337 a_35081_2511# a_35334_2498# a_34982_4680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3338 a_825_6014# a_1629_5833# a_1798_5391# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3339 a_22911_4823# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3340 a_11505_1690# a_12310_1924# a_12479_1482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3341 vdd d0 a_25880_5714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3342 a_24561_5665# a_24818_5475# a_24396_6597# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3343 gnd a_3383_4943# a_3175_4943# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3344 a_14788_7335# a_15045_7145# a_13779_6924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3345 a_10794_5223# a_11283_5041# a_11491_5041# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3346 a_36290_5346# a_36293_4754# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3347 gnd a_20346_3207# a_20138_3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3348 a_21913_1653# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3349 a_25611_7864# a_25621_7121# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3350 a_12140_3323# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3351 a_20887_n19# a_20674_n19# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3352 a_19021_3724# a_19125_2973# a_19080_2986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3353 a_625_4057# a_412_4057# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3354 a_26624_103# a_26411_103# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3355 a_40577_1978# a_40830_1965# a_40527_1558# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3356 a_396_6578# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3357 a_14799_4960# a_14807_4222# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3358 vdd d0 a_4399_4201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3359 a_21625_4805# a_22111_4589# a_22319_4589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3360 a_13732_5702# a_13989_5512# a_13567_6634# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3361 a_11491_5041# a_12295_4860# a_12454_5280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3362 a_19025_3547# a_19120_3954# a_19071_4144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3363 a_29842_5644# a_30099_5454# a_29677_6576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3364 a_2153_220# a_2880_4511# a_2831_4701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3365 a_10811_1906# a_11297_1690# a_11505_1690# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3366 a_16767_6001# a_17571_5820# a_17740_5378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3367 vdd d0 a_4398_3786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3368 vdd a_24673_2490# a_24465_2490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3369 a_610_6993# a_397_6993# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3370 a_133_4933# a_622_5033# a_830_5033# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3371 a_38244_7517# a_37823_7517# a_37550_7733# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3372 a_9443_837# a_9696_824# a_8427_1195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3373 vdd a_41843_2199# a_41635_2199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3374 a_29880_8024# a_30137_7834# a_29834_7427# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3375 vdd d0 a_20326_7124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3376 a_38041_6536# a_37828_6536# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3377 a_30909_6121# a_30905_6298# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3378 gnd a_19325_4930# a_19117_4930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3379 a_29900_4107# a_30961_3736# a_30916_3749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3380 a_11506_2105# a_11085_2105# a_10809_2005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3381 vdd d0 a_41835_2763# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3382 a_36276_7695# a_36272_7872# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3383 a_5409_5893# a_5411_5794# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3384 a_23327_6271# a_23114_6271# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3385 a_33572_4831# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3386 a_5923_1095# a_5710_1095# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3387 a_1622_6812# a_1409_6812# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3388 a_37835_5557# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3389 a_19080_2986# a_20138_3207# a_20093_3220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3390 a_32574_1661# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3391 vdd d2 a_3348_1587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3392 a_13795_3184# a_14856_2813# a_14811_2826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3393 a_6740_7211# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3394 a_24615_5908# a_24868_5895# a_24565_5488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3395 a_13492_4709# a_13749_4519# a_12814_228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3396 vdd d1 a_14052_2994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3397 a_1416_5833# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3398 gnd d0 a_36542_6137# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3399 a_2140_4308# a_1719_4308# a_2045_6300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3400 a_21893_5570# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3401 vdd d0 a_20340_3773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3402 gnd a_8672_2965# a_8464_2965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3403 gnd d1 a_3403_1026# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3404 vdd d2 a_30119_1537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3405 a_12120_7240# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3406 vdd d0 a_25874_7108# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3407 a_16083_3245# a_16572_3063# a_16780_3063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3408 a_35296_1999# a_36354_2220# a_36305_2410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3409 vdd a_14059_2015# a_13851_2015# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3410 a_845_2097# a_424_2097# a_148_2279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3411 a_7062_7211# a_6953_7211# a_7161_7211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3412 a_6119_3055# a_6923_2874# a_7082_3294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3413 vdd a_25881_6129# a_25673_6129# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3414 a_24615_5908# a_25673_6129# a_25624_6319# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3415 a_39245_1313# a_38873_893# a_38282_1074# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3416 a_7325_199# a_7112_199# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3417 a_16780_3063# a_17584_2882# a_17743_3302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3418 a_26926_1462# a_26924_1248# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3419 a_10603_125# a_20887_n19# vout SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3420 a_150_2493# a_148_2279# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3421 a_16345_5586# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3422 gnd d3 a_24673_2490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3423 a_18082_4295# a_17661_4295# a_17987_6287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3424 a_7099_1453# a_6717_1895# a_6126_2076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3425 gnd d0 a_15052_6166# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3426 a_38861_2853# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3427 a_16772_5020# a_16351_5020# a_16075_4920# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3428 a_3059_7654# a_3163_6903# a_3118_6916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3429 a_1491_1355# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3430 a_7074_5251# a_6702_4831# a_6110_4597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3431 a_27600_4568# a_27179_4568# a_26909_4403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3432 a_37848_2619# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3433 a_130_5815# a_135_5429# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3434 a_2153_220# a_2880_4511# a_2835_4524# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3435 a_6705_3855# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3436 a_30922_3183# a_30918_3360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3437 a_5678_6972# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3438 a_16063_6880# a_16552_6980# a_16760_6980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3439 a_5417_3936# a_5906_4036# a_6114_4036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3440 a_6125_1661# a_5704_1661# a_5436_1491# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3441 a_37548_7832# a_37550_7733# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3442 gnd a_9697_1239# a_9489_1239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3443 a_26894_7339# a_26892_7125# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3444 a_35061_6428# a_35314_6415# a_34986_4503# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3445 vdd a_24826_3518# a_24618_3518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3446 a_16359_3063# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3447 a_32274_7368# a_32272_7154# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3448 a_4121_7893# a_4131_7150# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3449 gnd a_4398_3786# a_4190_3786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3450 a_10603_125# a_10182_125# a_5342_132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3451 a_10182_125# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3452 vdd a_30162_2936# a_29954_2936# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3453 a_10782_6901# a_10784_6802# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3454 a_40558_5091# a_40815_4901# a_40503_5652# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3455 a_32563_4036# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3456 gnd a_20326_7124# a_20118_7124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3457 a_17576_4839# a_17363_4839# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3458 gnd a_41835_2763# a_41627_2763# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3459 a_19001_7641# a_19105_6890# a_19060_6903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3460 a_136_4239# a_625_4057# a_833_4057# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3461 a_4154_2431# a_4157_1839# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3462 a_29846_5467# a_29941_5874# a_29892_6064# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3463 a_16578_1669# a_16365_1669# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3464 a_28812_4258# a_28415_2333# a_28683_1305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3465 a_18095_207# a_18822_4498# a_18777_4511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3466 vdd d1 a_3403_1026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3467 a_35296_1999# a_36354_2220# a_36309_2233# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3468 a_38261_4576# a_37840_4576# a_37567_4792# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3469 a_19083_2184# a_19340_1994# a_19037_1587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3470 vdd a_24881_2957# a_24673_2957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3471 a_30918_3360# a_30921_2768# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3472 a_12913_228# a_12492_228# a_12814_228# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3473 vdd d3 a_19125_2506# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3474 a_6105_5578# a_5684_5578# a_5411_5794# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3475 a_29901_4906# a_30959_5127# a_30914_5140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3476 a_5902_4597# a_5689_4597# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3477 a_10797_4247# a_10797_3965# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3478 a_12492_228# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3479 a_3146_1216# a_4207_845# a_4158_1035# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3480 a_33622_5251# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3481 a_11073_4065# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3482 gnd d0 a_9696_824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3483 a_10784_6802# a_10791_6418# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3484 vdd d0 a_15052_6166# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3485 a_3079_3737# a_3336_3547# a_2930_2532# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3486 a_24581_1748# a_24685_997# a_24640_1010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3487 a_29866_1550# a_30119_1537# a_29697_2659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3488 vdd d0 a_20320_7690# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3489 a_39473_4266# a_39076_2341# a_39332_3273# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3490 a_824_5599# a_403_5599# a_135_5429# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3491 a_36277_8110# a_36530_8097# a_35264_7876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3492 a_28816_6250# a_28395_6250# a_28651_7182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3493 a_4130_6735# a_4126_6912# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3494 a_412_4057# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3495 a_11089_709# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3496 a_26894_6744# a_27380_6528# a_27588_6528# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3497 a_21638_1968# a_22127_2068# a_22335_2068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3498 a_35057_6605# a_35314_6415# a_34986_4503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3499 a_28572_3265# a_28463_3265# a_28671_3265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3500 gnd a_40615_2477# a_40407_2477# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3501 a_27187_2611# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3502 vdd a_4398_3786# a_4190_3786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3503 a_35226_5496# a_35479_5483# a_35057_6605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3504 vdd a_20326_7124# a_20118_7124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3505 a_23114_6271# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3506 vdd a_41835_2763# a_41627_2763# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3507 a_11498_2669# a_11077_2669# a_10811_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3508 a_24608_6887# a_24861_6874# a_24549_7625# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3509 a_8406_5916# a_9464_6137# a_9419_6150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3510 gnd a_25901_2212# a_25693_2212# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3511 vdd d1 a_35542_2965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3512 a_26899_6146# a_27388_5964# a_27596_5964# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3513 a_40267_4482# a_40520_4469# a_39585_178# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3514 a_5710_1095# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3515 vdd a_3348_1587# a_3140_1587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3516 a_38911_3273# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3517 gnd a_3183_2519# a_2975_2519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3518 a_33855_1334# a_33642_1334# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3519 vdd a_14052_2994# a_13844_2994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3520 vdd a_31150_8068# a_30942_8068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3521 a_32281_5794# a_32286_5408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3522 vdd a_35549_1986# a_35341_1986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3523 a_29884_7847# a_30942_8068# a_30893_8258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3524 gnd d0 a_41816_7095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3525 gnd a_36542_6137# a_36334_6137# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3526 a_37562_6368# a_38041_6536# a_38249_6536# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3527 gnd a_3403_1026# a_3195_1026# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3528 vdd a_25874_7108# a_25666_7108# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3529 a_28663_5222# a_28242_5222# a_28569_5341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3530 a_13779_6924# a_14837_7145# a_14788_7335# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3531 a_35285_3155# a_36346_2784# a_36297_2974# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3532 a_34986_4503# a_35239_4490# a_34304_199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3533 a_6130_680# a_5709_680# a_5436_896# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3534 a_33937_7330# a_33555_7772# a_32964_7953# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3535 a_13744_3568# a_13839_3975# a_13790_4165# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3536 a_17986_207# a_17773_207# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3537 a_8431_1018# a_9489_1239# a_9440_1429# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3538 gnd d0 a_20321_8105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3539 a_16065_7376# a_16546_7546# a_16754_7546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3540 a_27167_6528# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3541 a_11282_4626# a_11069_4626# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3542 a_26892_6843# a_26894_6744# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3543 a_23127_3847# a_22914_3847# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3544 a_17626_5259# a_17413_5259# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3545 a_12365_1363# a_12152_1363# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3546 a_13790_4165# a_14851_3794# a_14802_3984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3547 vdd d1 a_19328_3954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3548 a_38264_3600# a_37843_3600# a_37570_3816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3549 gnd a_15052_6166# a_14844_6166# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3550 a_22106_5570# a_21893_5570# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3551 a_22303_7945# a_21882_7945# a_21606_8127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3552 a_36305_2410# a_36308_1818# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3553 a_4153_2016# a_4163_1273# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3554 a_25624_6319# a_25627_5727# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3555 a_621_4618# a_408_4618# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3556 a_32756_7953# a_32543_7953# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3557 a_32269_7754# a_32755_7538# a_32963_7538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3558 vdd d3 a_24653_6407# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3559 a_148_1997# a_637_2097# a_845_2097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3560 vdd d0 a_25894_3191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3561 a_25647_1810# a_25900_1797# a_24631_2168# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3562 a_6965_5251# a_6752_5251# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3563 a_35222_5673# a_35479_5483# a_35057_6605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3564 a_4127_7327# a_4384_7137# a_3118_6916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3565 a_30914_5140# a_31167_5127# a_29901_4906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3566 vdd a_25901_2212# a_25693_2212# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3567 a_40565_3938# a_41623_4159# a_41578_4172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3568 a_29916_1970# a_30169_1957# a_29866_1550# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3569 a_16571_2648# a_16358_2648# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3570 a_35260_8053# a_35517_7863# a_35214_7456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3571 a_38257_5972# a_39061_5791# a_39230_5349# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3572 a_20096_2418# a_20099_1826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3573 a_39269_6258# a_39056_6258# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3574 a_17363_4839# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3575 gnd d4 a_29859_4461# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3576 a_22906_5804# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3577 a_8395_7072# a_9456_6701# a_9407_6891# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3578 a_32761_6972# a_32548_6972# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3579 a_28393_6762# a_28180_6762# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3580 a_10816_925# a_10823_724# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3581 a_30928_1789# a_31181_1776# a_29912_2147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3582 a_16365_1669# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3583 a_11266_7982# a_11053_7982# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3584 gnd d1 a_8652_6882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3585 a_21618_5885# a_22107_5985# a_22315_5985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3586 vdd a_3403_1026# a_3195_1026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3587 a_27395_3592# a_27182_3592# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3588 a_41582_2776# a_41578_2953# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3589 a_13779_6924# a_14837_7145# a_14792_7158# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3590 a_28552_7182# a_28443_7182# a_28651_7182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3591 a_29681_6399# a_29934_6386# a_29606_4474# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3592 a_28187_5783# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3593 a_35285_3155# a_36346_2784# a_36301_2797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3594 a_27609_3026# a_28413_2845# a_28572_3265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3595 a_3133_3980# a_4191_4201# a_4146_4214# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3596 a_22119_2632# a_21906_2632# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3597 a_11485_5607# a_12290_5841# a_12459_5399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3598 a_37849_3034# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3599 a_12498_6308# a_12285_6308# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3600 vdd a_19125_2506# a_18917_2506# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3601 a_18848_6613# a_19062_5491# a_19013_5681# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3602 a_21907_3047# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3603 a_23390_3286# a_22969_3286# a_23296_3405# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3604 a_24416_2680# a_24630_1558# a_24585_1571# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3605 a_25641_3204# a_25894_3191# a_24628_2970# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3606 a_40523_1735# a_40627_984# a_40578_1174# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3607 gnd a_19290_1574# a_19082_1574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3608 a_38036_7517# a_37823_7517# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3609 vdd a_15052_6166# a_14844_6166# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3610 vdd a_35529_5903# a_35321_5903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3611 a_850_1116# a_1654_935# a_1813_1355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3612 a_41586_2389# a_41843_2199# a_40577_1978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3613 a_5689_4597# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3614 a_34304_199# a_34195_199# a_34403_199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3615 a_22981_1326# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3616 a_1649_1916# a_1436_1916# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3617 gnd d1 a_40798_7842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3618 a_9423_4754# a_9676_4741# a_8407_5112# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3619 a_32981_5012# a_32560_5012# a_32284_5194# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3620 a_28564_5222# a_28192_4802# a_27600_4568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3621 a_5402_6872# a_5404_6773# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3622 a_26907_3907# a_27396_4007# a_27604_4007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3623 a_3091_1777# a_3195_1026# a_3146_1216# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3624 a_27615_1632# a_27194_1632# a_26926_1462# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3625 a_1932_4308# a_1719_4308# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3626 gnd d0 a_41810_7661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3627 a_39572_4266# a_39476_178# a_37394_111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3628 a_6925_2362# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3629 a_12479_1482# a_12365_1363# a_12573_1363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3630 vdd d1 a_14032_6911# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3631 a_7213_4287# a_7000_4287# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3632 a_16774_3629# a_17579_3863# a_17748_3421# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3633 a_13770_8082# a_14831_7711# a_14782_7901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3634 a_16546_7546# a_16333_7546# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3635 a_39312_7190# a_38891_7190# a_39218_7309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3636 a_20096_2418# a_20353_2228# a_19087_2007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3637 a_16063_7162# a_16552_6980# a_16760_6980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3638 vdd a_14039_5932# a_13831_5932# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3639 gnd d2 a_24826_3518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3640 a_25648_2225# a_25644_2402# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3641 vdd d4 a_29859_4461# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3642 a_41570_4910# a_41578_4172# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3643 a_38841_6770# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3644 vdd a_9685_3199# a_9477_3199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3645 vdd a_35542_2965# a_35334_2965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3646 a_30908_5706# a_30904_5883# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3647 a_11491_5041# a_11070_5041# a_10794_5223# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3648 a_30924_1966# a_31181_1776# a_29912_2147# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3649 vdd a_20357_832# a_20149_832# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3650 a_19033_1764# a_19137_1013# a_19088_1203# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3651 a_17874_4295# a_17661_4295# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3652 gnd a_31169_3736# a_30961_3736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3653 a_1692_3315# a_1479_3315# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3654 a_37594_674# a_38073_659# a_38281_659# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3655 a_29677_6576# a_29934_6386# a_29606_4474# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3656 a_16767_6001# a_16346_6001# a_16070_6183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3657 vdd a_40595_6394# a_40387_6394# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3658 a_143_3472# a_141_3258# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3659 a_32579_680# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3660 a_5404_6773# a_5411_6389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3661 gnd a_41816_7095# a_41608_7095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3662 a_7079_5370# a_6697_5812# a_6106_5993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3663 a_25623_5904# a_25633_5161# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3664 a_32984_4036# a_33788_3855# a_33957_3413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3665 a_16791_688# a_16370_688# a_16097_904# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3666 a_14818_1847# a_15071_1834# a_13802_2205# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3667 a_16339_6980# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3668 a_27595_5549# a_27174_5549# a_26901_5765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3669 gnd a_40760_5462# a_40552_5462# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3670 a_6915_4831# a_6702_4831# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3671 a_16370_688# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3672 a_6905_6279# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3673 a_40553_6072# a_40810_5882# a_40507_5475# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3674 a_21633_3443# a_21631_3229# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3675 a_17596_922# a_17383_922# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3676 a_19005_7464# a_19258_7451# a_18852_6436# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3677 a_12454_5280# a_12345_5280# a_12553_5280# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3678 a_5917_1661# a_5704_1661# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3679 a_19005_7464# a_19100_7871# a_19055_7884# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3680 vdd a_19290_1574# a_19082_1574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3681 a_12295_4860# a_12082_4860# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3682 a_9423_4754# a_9419_4931# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3683 a_24569_3708# a_24826_3518# a_24420_2503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3684 a_20068_8118# a_20064_8295# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3685 a_17413_5259# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3686 a_12152_1363# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3687 a_28443_7182# a_28230_7182# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3688 vdd a_19328_3954# a_19120_3954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3689 a_36288_5735# a_36284_5912# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3690 a_9419_4931# a_9676_4741# a_8407_5112# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3691 a_4151_3233# a_4404_3220# a_3138_2999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3692 a_6119_3055# a_5698_3055# a_5422_3237# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3693 gnd d0 a_20352_1813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3694 a_21633_2848# a_22119_2632# a_22327_2632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3695 a_35265_7072# a_36326_6701# a_36281_6714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3696 a_41582_2776# a_41835_2763# a_40566_3134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3697 vdd d3 a_8464_2498# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3698 a_16780_3063# a_16359_3063# a_16083_3245# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3699 a_3091_1777# a_3195_1026# a_3150_1039# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3700 a_12541_7240# a_12498_6308# a_12706_6308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3701 a_21918_672# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3702 a_5134_132# a_4921_132# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3703 vdd d0 a_41810_7661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3704 a_4145_3799# a_4141_3976# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3705 gnd d3 a_40595_6394# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3706 a_7082_3294# a_6710_2874# a_6119_3055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3707 a_116_8156# a_605_7974# a_813_7974# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3708 a_7193_1334# a_6772_1334# a_7094_1334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3709 a_13770_8082# a_14831_7711# a_14786_7724# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3710 a_838_3076# a_417_3076# a_141_2976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3711 a_118_7775# a_123_7389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3712 vdd a_8652_6882# a_8444_6882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3713 vdd d1 a_3383_4943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3714 vdd a_25894_3191# a_25686_3191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3715 a_29909_2949# a_30162_2936# a_29850_3687# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3716 a_13496_4532# a_13616_6444# a_13567_6634# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3717 a_6752_5251# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3718 a_38250_6951# a_39054_6770# a_39213_7190# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3719 gnd a_3088_4511# a_2880_4511# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3720 vdd a_20341_4188# a_20133_4188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3721 a_37843_3600# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3722 a_8422_2176# a_9483_1805# a_9438_1818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3723 a_812_7559# a_1617_7793# a_1786_7351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3724 a_5897_5578# a_5684_5578# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3725 a_19063_6101# a_19320_5911# a_19017_5504# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3726 a_13756_1608# a_14009_1595# a_13587_2717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3727 a_19033_1764# a_19137_1013# a_19092_1026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3728 a_20092_2805# a_20345_2792# a_19076_3163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3729 a_6094_7953# a_6898_7772# a_7067_7330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3730 a_10782_6901# a_11271_7001# a_11479_7001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3731 a_39056_6258# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3732 a_21901_3613# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3733 vdd a_31169_3736# a_30961_3736# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3734 a_26924_1248# a_26924_966# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3735 a_38265_4015# a_37844_4015# a_37568_3915# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3736 a_21638_1968# a_21640_1869# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3737 a_28180_6762# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3738 a_5434_995# a_5923_1095# a_6131_1095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3739 a_11053_7982# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3740 a_21620_6381# a_22099_6549# a_22307_6549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3741 a_27182_3592# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3742 a_16095_1003# a_16584_1103# a_16792_1103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3743 vdd a_40760_5462# a_40552_5462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3744 a_13496_4532# a_13749_4519# a_12814_228# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3745 a_622_5033# a_409_5033# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3746 gnd d0 a_25889_4172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3747 a_19001_7641# a_19258_7451# a_18852_6436# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3748 gnd d2 a_30119_1537# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3749 a_12285_6308# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3750 a_8356_5496# a_8609_5483# a_8187_6605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3751 gnd d1 a_24876_3938# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3752 gnd a_25881_6129# a_25673_6129# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3753 a_41566_6306# a_41569_5714# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3754 a_30904_5883# a_31161_5693# a_29892_6064# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3755 a_37823_7517# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3756 a_4133_5933# a_4143_5190# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3757 a_4147_3410# a_4404_3220# a_3138_2999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3758 a_10794_4941# a_10796_4842# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3759 a_41578_2953# a_41835_2763# a_40566_3134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3760 vdd a_40520_4469# a_40312_4469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3761 a_37568_4197# a_37568_3915# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3762 a_2926_2709# a_3140_1587# a_3091_1777# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3763 a_636_1682# a_423_1682# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3764 a_1436_1916# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3765 a_2041_4308# a_1644_2383# a_1900_3315# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3766 gnd a_40798_7842# a_40590_7842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3767 a_40267_4482# a_40387_6394# a_40342_6407# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3768 a_26887_8106# a_26887_7824# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3769 a_141_2976# a_143_2877# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3770 a_32267_8135# a_32267_7853# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3771 a_28589_1424# a_28207_1866# a_27616_2047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3772 a_13496_4532# a_13616_6444# a_13571_6457# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3773 a_14806_3807# a_14802_3984# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3774 a_25617_7298# a_25874_7108# a_24608_6887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3775 vdd a_19270_5491# a_19062_5491# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3776 vdd a_3088_4511# a_2880_4511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3777 a_10504_125# a_15582_140# a_15904_140# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3778 vdd a_14032_6911# a_13824_6911# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3779 a_15582_140# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3780 a_12345_5280# a_12132_5280# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3781 a_16333_7546# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3782 a_11277_5607# a_11064_5607# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3783 a_36294_5169# a_36547_5156# a_35281_4935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3784 a_41578_4172# a_41574_4349# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3785 gnd a_24826_3518# a_24618_3518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3786 a_38873_893# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3787 a_1441_935# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3788 a_35296_1999# a_35549_1986# a_35246_1579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3789 a_17378_1903# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3790 a_32780_2640# a_32567_2640# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3791 a_21608_7746# a_21613_7360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3792 a_429_1116# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3793 a_24420_2503# a_24673_2490# a_24321_4672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3794 a_10796_4842# a_10799_4461# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3795 gnd d4 a_35239_4490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3796 a_17661_4295# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3797 a_6717_1895# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3798 a_7062_7211# a_6690_6791# a_6099_6972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3799 a_36308_1818# a_36561_1805# a_35292_2176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3800 a_16759_6565# a_16338_6565# a_16065_6781# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3801 vdd a_19030_4498# a_18822_4498# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3802 vdd d0 a_25889_4172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3803 a_6113_3621# a_5692_3621# a_5419_3837# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3804 a_143_2877# a_150_2493# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3805 a_30909_6121# a_31162_6108# a_29896_5887# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3806 a_14819_2262# a_14815_2439# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3807 a_5910_2640# a_5697_2640# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3808 a_6702_4831# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3809 a_23643_191# a_24370_4482# a_24321_4672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3810 gnd a_4410_1826# a_4202_1826# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3811 a_25615_7687# a_25611_7864# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3812 a_32963_7538# a_32542_7538# a_32274_7368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3813 a_8352_5673# a_8609_5483# a_8187_6605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3814 a_39218_7309# a_39104_7190# a_39312_7190# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3815 a_14804_5198# a_15057_5185# a_13791_4964# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3816 vdd d0 a_15060_4209# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3817 a_17383_922# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3818 a_5704_1661# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3819 a_14819_1043# a_10823_724# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3820 a_11290_2669# a_11077_2669# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3821 a_17564_6799# a_17351_6799# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3822 a_12082_4860# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3823 a_832_3642# a_411_3642# a_143_3472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3824 gnd d0 a_4411_2241# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3825 a_29901_4906# a_30959_5127# a_30910_5317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3826 a_5416_4813# a_5902_4597# a_6110_4597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3827 a_16566_3629# a_16353_3629# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3828 a_27413_1066# a_27200_1066# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3829 vdd d2 a_24838_1558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3830 a_28230_7182# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3831 a_17358_5820# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3832 a_23174_5243# a_22961_5243# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3833 gnd a_20352_1813# a_20144_1813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3834 a_28388_7743# a_28175_7743# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3835 a_3083_3560# a_3336_3547# a_2930_2532# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3836 vdd a_8464_2498# a_8256_2498# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3837 gnd d1 a_24893_997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3838 a_32788_2076# a_32575_2076# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3839 a_22327_2632# a_23132_2866# a_23291_3286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3840 gnd d0 a_20338_5164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3841 a_29912_2147# a_30973_1776# a_30924_1966# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3842 a_14787_8139# a_14783_8316# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3843 a_11473_7567# a_11052_7567# a_10784_7397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3844 a_16080_4440# a_16563_4605# a_16771_4605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3845 gnd d1 a_30169_1957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3846 a_28703_4258# a_28490_4258# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3847 a_5890_6557# a_5677_6557# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3848 a_8406_5916# a_8659_5903# a_8356_5496# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3849 gnd d1 a_14064_1034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3850 a_33800_1895# a_33587_1895# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3851 a_36290_5346# a_36547_5156# a_35281_4935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3852 a_35214_7456# a_35309_7863# a_35260_8053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3853 a_33642_1334# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3854 a_5684_5578# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3855 a_34403_199# a_33982_199# a_34304_199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3856 a_812_7559# a_391_7559# a_118_7775# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3857 a_35260_8053# a_36321_7682# a_36272_7872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3858 a_37829_6951# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3859 a_23283_5243# a_22911_4823# a_22320_5004# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3860 a_3095_1600# a_3190_2007# a_3141_2197# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3861 a_8406_5916# a_9464_6137# a_9415_6327# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3862 a_22334_1653# a_21913_1653# a_21640_1869# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3863 a_28569_5341# a_28187_5783# a_27596_5964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3864 gnd a_36549_3765# a_36341_3765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3865 a_28463_3265# a_28250_3265# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3866 a_9419_6150# a_9415_6327# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3867 a_14783_8316# a_14786_7724# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3868 gnd a_31150_8068# a_30942_8068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3869 a_23643_191# a_24370_4482# a_24325_4495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3870 a_10791_5823# a_11277_5607# a_11485_5607# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3871 a_39364_4266# a_39151_4266# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3872 a_38257_5972# a_37836_5972# a_37560_6154# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3873 a_14800_5375# a_15057_5185# a_13791_4964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3874 a_17634_3302# a_17421_3302# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3875 a_20068_6899# a_20325_6709# a_19056_7080# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3876 vdd d1 a_35554_1005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3877 gnd a_24876_3938# a_24668_3938# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3878 vdd d0 a_4411_2241# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3879 a_16339_6980# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3880 a_11302_709# a_11089_709# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3881 a_19037_1587# a_19132_1994# a_19083_2184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3882 a_27609_3026# a_27188_3026# a_26912_3208# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3883 a_135_5429# a_616_5599# a_824_5599# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3884 a_36288_5735# a_36541_5722# a_35272_6093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3885 gnd a_15059_3794# a_14851_3794# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3886 a_16583_688# a_16370_688# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3887 a_29892_6064# a_30149_5874# a_29846_5467# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3888 vdd d0 a_20338_5164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3889 a_25641_3204# a_25637_3381# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3890 a_35297_1195# a_36358_824# a_36309_1014# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3891 a_29912_2147# a_30973_1776# a_30928_1789# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3892 a_423_1682# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3893 a_22899_6783# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3894 a_37575_2835# a_38061_2619# a_38269_2619# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3895 a_28572_3265# a_28200_2845# a_27609_3026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3896 a_28683_1305# a_28262_1305# a_28584_1305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3897 gnd a_3371_6903# a_3163_6903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3898 a_1634_4852# a_1421_4852# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3899 a_41563_7108# a_41816_7095# a_40550_6874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3900 a_34195_199# a_33982_199# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3901 vdd d1 a_14064_1034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3902 a_34031_7211# a_33988_6279# a_34196_6279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3903 a_33957_3413# a_33575_3855# a_32983_3621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3904 a_11270_6586# a_11057_6586# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3905 a_13786_5945# a_14039_5932# a_13736_5525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3906 a_21645_888# a_22131_672# a_22339_672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3907 a_13802_2205# a_14863_1834# a_14814_2024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3908 a_36293_4754# a_36289_4931# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3909 a_16080_3845# a_16566_3629# a_16774_3629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3910 gnd a_8684_1005# a_8476_1005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3911 a_17614_7219# a_17401_7219# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3912 a_12132_5280# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3913 a_27393_4983# a_27180_4983# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3914 a_35289_2978# a_35542_2965# a_35230_3716# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3915 a_11064_5607# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3916 a_39476_178# a_39263_178# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3917 a_27584_7924# a_28388_7743# a_28557_7301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3918 a_35260_8053# a_36321_7682# a_36276_7695# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3919 a_14798_5764# a_15051_5751# a_13782_6122# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3920 a_2906_6626# a_3120_5504# a_3075_5517# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3921 gnd a_9659_7682# a_9451_7682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3922 a_4131_7150# a_4384_7137# a_3118_6916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3923 vdd d1 a_30154_4893# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3924 a_22307_6549# a_23112_6783# a_23271_7203# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3925 a_10799_4461# a_10797_4247# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3926 a_3133_3980# a_3386_3967# a_3083_3560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3927 a_22323_4028# a_21902_4028# a_21626_3928# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3928 vdd a_41831_4159# a_41623_4159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3929 vdd a_36549_3765# a_36341_3765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3930 gnd d0 a_41827_4720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3931 a_40565_3938# a_41623_4159# a_41574_4349# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3932 a_37394_111# a_37285_111# a_31994_96# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3933 a_32272_6872# a_32761_6972# a_32969_6972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3934 a_25637_3381# a_25640_2789# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3935 a_21882_7945# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3936 a_40507_5475# a_40602_5882# a_40553_6072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3937 a_33780_5812# a_33567_5812# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3938 a_12467_3442# a_12085_3884# a_11493_3650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3939 a_19088_1203# a_20149_832# a_20104_845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3940 a_5414_4912# a_5416_4813# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3941 gnd d0 a_20332_5730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3942 a_37585_974# a_38074_1074# a_38282_1074# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3943 a_6923_2874# a_6710_2874# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3944 a_13799_3007# a_14052_2994# a_13740_3745# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3945 gnd d2 a_35499_1566# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3946 a_3071_5694# a_3175_4943# a_3130_4956# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3947 a_33949_5370# a_33835_5251# a_34043_5251# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3948 a_6985_1334# a_6772_1334# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3949 a_24396_6597# a_24653_6407# a_24325_4495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3950 a_38244_7517# a_39049_7751# a_39218_7309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3951 a_19075_3967# a_19328_3954# a_19025_3547# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3952 a_17351_6799# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3953 a_3075_5517# a_3170_5924# a_3121_6114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3954 a_28815_170# a_28602_170# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3955 a_5429_1976# a_5918_2076# a_6126_2076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3956 a_11278_6022# a_11065_6022# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3957 a_36284_5912# a_36541_5722# a_35272_6093# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3958 a_19075_3967# a_20133_4188# a_20084_4378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3959 gnd d0 a_4403_2805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3960 a_27200_1066# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3961 vdd a_24838_1558# a_24630_1558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3962 a_818_6993# a_397_6993# a_121_6893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3963 a_16353_3629# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3964 a_24416_2680# a_24630_1558# a_24581_1748# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3965 a_20067_7703# a_20063_7880# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3966 a_32781_3055# a_32568_3055# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3967 a_39477_6258# a_39364_4266# a_39572_4266# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3968 a_22335_2068# a_23139_1887# a_23308_1445# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3969 a_28175_7743# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3970 a_12290_5841# a_12077_5841# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3971 gnd d0 a_25869_8089# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3972 vdd d1 a_8659_5903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3973 gnd a_24893_997# a_24685_997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3974 a_32575_2076# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3975 gnd a_20338_5164# a_20130_5164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3976 a_8399_6895# a_8652_6882# a_8340_7633# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3977 a_19013_5681# a_19117_4930# a_19072_4943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3978 a_155_1512# a_153_1298# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3979 a_617_6014# a_404_6014# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3980 a_16070_6183# a_16070_5901# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3981 gnd a_41847_803# a_41639_803# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3982 gnd d2 a_14009_1595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3983 a_11506_2105# a_12310_1924# a_12479_1482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3984 a_28490_4258# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3985 a_19017_5504# a_19112_5911# a_19063_6101# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3986 a_2041_4308# a_1932_4308# a_2140_4308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3987 gnd a_14064_1034# a_13856_1034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3988 a_27199_651# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3989 vdd a_9659_7682# a_9451_7682# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3990 a_14794_5941# a_15051_5751# a_13782_6122# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3991 a_22931_906# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3992 gnd a_15039_7711# a_14831_7711# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3993 a_11291_3084# a_11078_3084# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3994 a_8360_3716# a_8464_2965# a_8419_2978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3995 a_136_4239# a_136_3957# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3996 a_17987_6287# a_17874_4295# a_18082_4295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3997 a_39074_2853# a_38861_2853# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3998 a_29892_6064# a_30953_5693# a_30908_5706# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3999 vdd d0 a_41827_4720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4000 a_20100_2241# a_20353_2228# a_19087_2007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4001 a_20080_6158# a_20076_6335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4002 a_16567_4044# a_16354_4044# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4003 a_123_6794# a_130_6410# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4004 a_27603_3592# a_27182_3592# a_26909_3808# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4005 a_11510_709# a_12315_943# a_12474_1363# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4006 a_38250_6951# a_37829_6951# a_37553_7133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4007 a_28250_3265# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4008 a_1801_3315# a_1692_3315# a_1900_3315# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4009 a_1857_2383# a_1644_2383# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4010 a_17728_7338# a_17614_7219# a_17822_7219# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4011 vdd d0 a_20332_5730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4012 a_39151_4266# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4013 a_16786_1669# a_17591_1903# a_17760_1461# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4014 gnd a_8664_4922# a_8456_4922# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4015 a_630_3076# a_417_3076# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4016 vdd d2 a_35499_1566# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4017 a_21613_6765# a_21620_6381# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4018 a_4157_1839# a_4153_2016# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4019 a_6094_7953# a_5673_7953# a_5397_8135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4020 a_21608_7746# a_22094_7530# a_22302_7530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4021 a_17421_3302# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4022 a_41557_7674# a_41810_7661# a_40541_8032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4023 vdd a_35554_1005# a_35346_1005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4024 a_26906_4784# a_27392_4568# a_27600_4568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4025 a_38891_7190# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4026 a_26909_4403# a_26907_4189# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4027 a_29885_7043# a_30142_6853# a_29830_7604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4028 a_11511_1124# a_11090_1124# a_10814_1024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4029 a_30921_2768# a_30917_2945# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4030 a_24573_3531# a_24826_3518# a_24420_2503# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4031 a_18872_2519# a_19125_2506# a_18773_4688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4032 a_39054_6770# a_38841_6770# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4033 a_16083_3245# a_16083_2963# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4034 gnd d0 a_25906_1231# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4035 vdd a_20338_5164# a_20130_5164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4036 a_10797_3965# a_10799_3866# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4037 a_12447_7359# a_12065_7801# a_11473_7567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4038 a_28608_6250# a_28395_6250# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4039 a_37840_4576# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4040 a_13779_6924# a_14032_6911# a_13720_7662# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4041 a_1421_4852# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4042 a_37565_4891# a_38054_4991# a_38262_4991# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4043 a_6903_6791# a_6690_6791# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4044 a_37570_3816# a_37575_3430# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4045 a_20067_7703# a_20320_7690# a_19051_8061# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4046 a_40578_1174# a_40835_984# a_40523_1735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4047 vdd a_14064_1034# a_13856_1034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4048 gnd d1 a_35549_1986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4049 a_37565_4891# a_37567_4792# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4050 a_5905_3621# a_5692_3621# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4051 a_2140_4308# a_2044_220# a_2252_220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4052 a_6697_5812# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4053 a_29896_5887# a_30954_6108# a_30905_6298# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4054 a_7421_4287# a_7000_4287# a_7326_6279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4055 a_37570_4411# a_38053_4576# a_38261_4576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4056 a_32792_680# a_32579_680# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4057 gnd d0 a_4383_6722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4058 a_5409_5893# a_5898_5993# a_6106_5993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4059 vdd a_25886_5148# a_25678_5148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4060 a_38281_659# a_37860_659# a_37587_875# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4061 vdd a_19340_1994# a_19132_1994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4062 vdd a_15039_7711# a_14831_7711# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4063 a_17401_7219# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4064 a_27180_4983# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4065 a_13791_4964# a_14849_5185# a_14800_5375# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4066 a_24585_1571# a_24680_1978# a_24631_2168# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4067 vdd d1 a_24856_7855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4068 vdd a_30154_4893# a_29946_4893# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4069 a_27179_4568# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4070 a_26906_5379# a_26904_5165# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4071 a_7094_1334# a_6722_914# a_6131_1095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4072 a_23139_1887# a_22926_1887# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4073 a_128_6196# a_617_6014# a_825_6014# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4074 a_39225_5230# a_38853_4810# a_38262_4991# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4075 gnd a_41827_4720# a_41619_4720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4076 a_29862_1727# a_29966_976# a_29921_989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4077 gnd d2 a_13989_5512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4078 a_162_716# a_641_701# a_849_701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4079 a_5698_3055# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4080 a_38276_1640# a_37855_1640# a_37582_1856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4081 a_1459_7232# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4082 a_23422_4279# a_23209_4279# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4083 a_7181_3294# a_6760_3294# a_7087_3413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4084 a_31885_96# a_31672_96# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4085 a_37580_2237# a_37580_1955# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4086 a_629_2661# a_416_2661# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4087 gnd a_36530_8097# a_36322_8097# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4088 a_41553_7851# a_41810_7661# a_40541_8032# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4089 gnd a_20332_5730# a_20124_5730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4090 a_30909_4902# a_30917_4164# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4091 a_6710_2874# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4092 a_37567_4792# a_37570_4411# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4093 a_33843_3294# a_33630_3294# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4094 a_6772_1334# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4095 a_11271_7001# a_11058_7001# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4096 a_32768_5993# a_32555_5993# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4097 a_20104_845# a_20357_832# a_19088_1203# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4098 a_32281_5794# a_32767_5578# a_32975_5578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4099 a_14788_7335# a_14791_6743# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4100 a_11065_6022# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4101 a_38056_3600# a_37843_3600# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4102 gnd a_4403_2805# a_4195_2805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4103 a_39124_3273# a_38911_3273# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4104 vdd d0 a_25906_1231# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4105 a_4139_5367# a_4396_5177# a_3130_4956# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4106 a_2910_6449# a_3163_6436# a_2835_4524# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4107 a_27375_7509# a_27162_7509# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4108 a_610_6993# a_397_6993# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4109 gnd a_40520_4469# a_40312_4469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4110 gnd d2 a_8617_3526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4111 a_404_6014# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4112 a_609_6578# a_396_6578# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4113 vdd d0 a_4383_6722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4114 a_19055_7884# a_20113_8105# a_20068_8118# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4115 a_13791_4964# a_14849_5185# a_14804_5198# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4116 a_25627_5727# a_25623_5904# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4117 a_18852_6436# a_19105_6423# a_18777_4511# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4118 a_24623_3951# a_24876_3938# a_24573_3531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4119 a_39344_1313# a_38923_1313# a_39245_1313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4120 vdd a_41827_4720# a_41619_4720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4121 vdd d2 a_13989_5512# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4122 vdd d1 a_35534_4922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4123 a_16354_4044# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4124 a_32301_2472# a_32780_2640# a_32988_2640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4125 a_832_3642# a_1637_3876# a_1806_3434# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4126 a_30917_4164# a_31170_4151# a_29904_3930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4127 a_23402_1326# a_22981_1326# a_23308_1445# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4128 a_38048_5557# a_37835_5557# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4129 a_11078_3084# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4130 a_1801_3315# a_1429_2895# a_837_2661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4131 a_16779_2648# a_17584_2882# a_17743_3302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4132 a_20099_1826# a_20095_2003# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4133 vdd d1 a_3378_5924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4134 vdd a_20332_5730# a_20124_5730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4135 a_24561_5665# a_24665_4914# a_24620_4927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4136 a_10804_3480# a_11285_3650# a_11493_3650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4137 a_7322_4287# a_6925_2362# a_7181_3294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4138 a_829_4618# a_408_4618# a_135_4834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4139 a_35277_5112# a_36338_4741# a_36289_4931# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4140 a_5424_2856# a_5910_2640# a_6118_2640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4141 vdd d1 a_30149_5874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4142 a_26919_1947# a_27408_2047# a_27616_2047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4143 a_22302_7530# a_23107_7764# a_23276_7322# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4144 gnd d0 a_41822_5701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4145 a_32543_7953# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4146 a_23119_5804# a_22906_5804# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4147 vdd d1 a_14044_4951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4148 a_2906_6626# a_3163_6436# a_2835_4524# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4149 a_13782_6122# a_14843_5751# a_14794_5941# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4150 a_39324_5230# a_38903_5230# a_39230_5349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4151 gnd a_25906_1231# a_25698_1231# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4152 a_17799_2370# a_17586_2370# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4153 gnd d1 a_14039_5932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4154 vdd d2 a_8617_3526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4155 gnd d2 a_24838_1558# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4156 a_28395_6250# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4157 a_16779_2648# a_16358_2648# a_16092_2480# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4158 gnd d0 a_31174_2755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4159 a_6690_6791# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4160 a_22969_3286# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4161 a_36298_3389# a_36555_3199# a_35289_2978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4162 a_32969_6972# a_32548_6972# a_32272_7154# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4163 a_30905_6298# a_30908_5706# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4164 gnd a_31181_1776# a_30973_1776# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4165 a_22303_7945# a_21882_7945# a_21606_7845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4166 a_5692_3621# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4167 a_1704_1355# a_1491_1355# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4168 a_35077_2688# a_35291_1566# a_35242_1756# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4169 a_18848_6613# a_19105_6423# a_18777_4511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4170 a_4142_4391# a_4399_4201# a_3133_3980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4171 a_28816_6250# a_28703_4258# a_28911_4258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4172 a_13740_3745# a_13844_2994# a_13795_3184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4173 a_32996_2076# a_33800_1895# a_33969_1453# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4174 a_29850_3687# a_29954_2936# a_29909_2949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4175 a_5411_6389# a_5890_6557# a_6098_6557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4176 a_23162_7203# a_22949_7203# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4177 a_3134_3176# a_4195_2805# a_4146_2995# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4178 a_23132_2866# a_22919_2866# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4179 vdd a_24856_7855# a_24648_7855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4180 a_16563_4605# a_16350_4605# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4181 a_30913_4341# a_31170_4151# a_29904_3930# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4182 a_32776_4036# a_32563_4036# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4183 a_28408_3826# a_28195_3826# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4184 a_24581_1748# a_24838_1558# a_24416_2680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4185 vdd d1 a_19333_2973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4186 a_23291_3286# a_23182_3286# a_23390_3286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4187 vdd d0 a_25900_1797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4188 a_123_6794# a_609_6578# a_817_6578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4189 gnd d1 a_8667_3946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4190 a_14808_3418# a_15065_3228# a_13799_3007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4191 a_37285_111# a_37072_111# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4192 a_25653_1244# a_25649_1421# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4193 a_4163_1273# a_4416_1260# a_3150_1039# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4194 a_416_2661# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4195 a_27584_7924# a_27163_7924# a_26887_8106# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4196 a_35277_5112# a_36338_4741# a_36293_4754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4197 a_32761_6972# a_32548_6972# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4198 a_12553_5280# a_12132_5280# a_12454_5280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4199 a_33630_3294# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4200 a_25616_8102# a_26887_8106# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4201 a_32555_5993# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4202 a_30897_8081# a_32267_8135# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4203 a_37550_7733# a_38036_7517# a_38244_7517# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4204 a_16063_7162# a_16063_6880# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4205 a_10777_7882# a_10779_7783# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4206 a_13782_6122# a_14843_5751# a_14798_5764# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4207 a_21899_5004# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4208 a_29900_4107# a_30157_3917# a_29854_3510# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4209 vdd d0 a_20346_3207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4210 vdd a_25906_1231# a_25698_1231# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4211 a_11057_6586# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4212 a_11286_4065# a_11073_4065# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4213 a_29921_989# a_30174_976# a_29862_1727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4214 a_35265_7072# a_35522_6882# a_35210_7633# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4215 a_39069_3834# a_38856_3834# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4216 vdd a_31182_2191# a_30974_2191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4217 a_824_5599# a_1629_5833# a_1798_5391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4218 vdd d0 a_31174_2755# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4219 a_27162_7509# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4220 a_37550_7733# a_37555_7347# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4221 a_1837_6300# a_1624_6300# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4222 a_22911_4823# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4223 a_30896_7666# a_31149_7653# a_29880_8024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4224 a_10794_4941# a_11283_5041# a_11491_5041# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4225 vdd a_31181_1776# a_30973_1776# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4226 gnd d0 a_36562_2220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4227 a_3109_8074# a_3366_7884# a_3063_7477# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4228 a_25649_1421# a_25652_829# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4229 a_21913_1653# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4230 a_7118_6279# a_6905_6279# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4231 a_12140_3323# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4232 a_37860_659# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4233 a_38277_2055# a_37856_2055# a_37580_1955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4234 a_396_6578# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4235 gnd d0 a_15064_2813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4236 a_35077_2688# a_35291_1566# a_35246_1579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4237 a_35234_3539# a_35487_3526# a_35081_2511# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4238 a_24635_1991# a_25693_2212# a_25644_2402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4239 a_5886_7953# a_5673_7953# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4240 gnd a_15071_1834# a_14863_1834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4241 a_20088_2982# a_20100_2241# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4242 a_14807_4222# a_14803_4399# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4243 a_17779_6287# a_17566_6287# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4244 a_28584_1305# a_28212_885# a_27621_1066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4245 a_11506_2105# a_11085_2105# a_10809_2287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4246 a_23327_6271# a_23114_6271# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4247 a_38041_6536# a_37828_6536# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4248 a_7434_199# a_8161_4490# a_8112_4680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4249 a_19051_8061# a_19308_7871# a_19005_7464# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4250 vdd a_35534_4922# a_35326_4922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4251 a_29697_2659# a_29911_1537# a_29866_1550# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4252 a_18773_4688# a_18917_2506# a_18868_2696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4253 a_6740_7211# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4254 vdd d1 a_3371_6903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4255 a_40546_7051# a_41607_6680# a_41558_6870# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4256 a_37835_5557# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4257 gnd a_41831_4159# a_41623_4159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4258 a_4159_1450# a_4416_1260# a_3150_1039# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4259 gnd d1 a_40803_6861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4260 vdd a_3378_5924# a_3170_5924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4261 a_13720_7662# a_13824_6911# a_13775_7101# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4262 gnd a_40810_5882# a_40602_5882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4263 a_32976_5993# a_33780_5812# a_33949_5370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4264 a_16083_2963# a_16572_3063# a_16780_3063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4265 a_41590_993# a_41847_803# a_40578_1174# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4266 a_3114_7093# a_4175_6722# a_4126_6912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4267 a_21623_4904# a_21625_4805# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4268 a_6118_2640# a_6923_2874# a_7082_3294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4269 gnd d2 a_30107_3497# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4270 gnd d1 a_8684_1005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4271 gnd a_41822_5701# a_41614_5701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4272 a_25629_5338# a_25886_5148# a_24620_4927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4273 a_22114_3613# a_21901_3613# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4274 vdd d1 a_19313_6890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4275 a_4143_5190# a_4139_5367# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4276 vdd a_14044_4951# a_13836_4951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4277 a_14803_4399# a_14806_3807# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4278 vdd a_30174_976# a_29966_976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4279 a_30892_7843# a_31149_7653# a_29880_8024# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4280 vdd a_19320_5911# a_19112_5911# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4281 vdd d0 a_36562_2220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4282 a_17586_2370# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4283 gnd a_24838_1558# a_24630_1558# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4284 a_32292_3237# a_32781_3055# a_32989_3055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4285 a_8344_7456# a_8597_7443# a_8191_6428# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4286 a_41574_4733# a_41827_4720# a_40558_5091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4287 a_21902_4028# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4288 a_40362_2490# a_40560_3505# a_40511_3695# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4289 a_6935_914# a_6722_914# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4290 gnd a_31174_2755# a_30966_2755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4291 a_135_4834# a_138_4453# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4292 a_35230_3716# a_35487_3526# a_35081_2511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4293 a_7074_5251# a_6702_4831# a_6111_5012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4294 a_6973_3294# a_6760_3294# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4295 a_1491_1355# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4296 a_24635_1991# a_25693_2212# a_25648_2225# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4297 a_27600_4568# a_27179_4568# a_26906_4784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4298 gnd d0 a_4415_845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4299 a_10797_4247# a_11286_4065# a_11494_4065# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4300 vdd a_8667_3946# a_8459_3946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4301 a_6125_1661# a_5704_1661# a_5431_1877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4302 a_21625_4805# a_21628_4424# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4303 a_38265_4015# a_39069_3834# a_39238_3392# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4304 a_9407_8110# a_9403_8287# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4305 a_11266_7982# a_11053_7982# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4306 a_26887_7824# a_26889_7725# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4307 a_37553_7133# a_37553_6851# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4308 a_32267_7853# a_32269_7754# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4309 a_1880_7232# a_1459_7232# a_1781_7232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4310 a_32975_5578# a_32554_5578# a_32286_5408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4311 a_4139_5367# a_4142_4775# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4312 a_22094_7530# a_21881_7530# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4313 vdd d0 a_15072_2249# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4314 a_16350_4605# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4315 a_40546_7051# a_41607_6680# a_41562_6693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4316 vdd a_31161_5693# a_30953_5693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4317 a_17576_4839# a_17363_4839# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4318 a_32563_4036# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4319 a_28195_3826# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4320 a_844_1682# a_423_1682# a_155_1512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4321 a_1900_3315# a_1857_2383# a_2041_4308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4322 vdd a_19333_2973# a_19125_2973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4323 a_136_3957# a_625_4057# a_833_4057# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4324 a_30917_2945# a_30929_2204# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4325 a_2835_4524# a_2955_6436# a_2906_6626# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4326 a_36297_4193# a_36550_4180# a_35284_3959# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4327 vdd a_4415_845# a_4207_845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4328 a_40527_1558# a_40780_1545# a_40358_2667# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4329 a_16578_1669# a_16365_1669# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4330 a_10809_2005# a_10811_1906# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4331 a_28812_4258# a_28415_2333# a_28671_3265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4332 a_18872_2519# a_19070_3534# a_19021_3724# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4333 a_26914_2827# a_27400_2611# a_27608_2611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4334 a_8372_1756# a_8476_1005# a_8431_1018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4335 vdd d1 a_24888_1978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4336 a_3095_1600# a_3348_1587# a_2926_2709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4337 a_3114_7093# a_4175_6722# a_4130_6735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4338 a_35077_2688# a_35334_2498# a_34982_4680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4339 a_32306_896# a_32313_695# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4340 vdd d0 a_9664_6701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4341 a_23370_7203# a_23327_6271# a_23535_6271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4342 a_9403_8287# a_9406_7695# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4343 a_12913_228# a_12492_228# a_12801_4316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4344 vdd a_20346_3207# a_20138_3207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4345 a_12492_228# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4346 a_11073_4065# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4347 a_34304_199# a_35031_4490# a_34986_4503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4348 a_27412_651# a_27199_651# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4349 a_8340_7633# a_8597_7443# a_8191_6428# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4350 a_41570_4910# a_41827_4720# a_40558_5091# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4351 vdd a_31174_2755# a_30966_2755# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4352 a_1624_6300# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4353 a_38270_3034# a_37849_3034# a_37573_2934# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4354 gnd a_36562_2220# a_36354_2220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4355 a_32988_2640# a_32567_2640# a_32294_2856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4356 a_26904_5165# a_26904_4883# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4357 a_29904_3930# a_30962_4151# a_30913_4341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4358 gnd d0 a_36554_2784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4359 a_32284_5194# a_32284_4912# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4360 a_6098_6557# a_6903_6791# a_7062_7211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4361 gnd d0 a_31155_7087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4362 a_6114_4036# a_5693_4036# a_5417_3936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4363 gnd a_15064_2813# a_14856_2813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4364 gnd a_36561_1805# a_36353_1805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4365 gnd d2 a_30087_7414# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4366 a_20068_6899# a_20080_6158# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4367 a_26901_6360# a_27380_6528# a_27588_6528# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4368 a_27187_2611# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4369 a_24624_3147# a_25685_2776# a_25636_2966# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4370 a_5673_7953# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4371 a_17723_7219# a_17351_6799# a_16759_6565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4372 a_24325_4495# a_24578_4482# a_23643_191# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4373 a_41595_1231# a_41591_1408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4374 a_17566_6287# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4375 gnd a_25886_5148# a_25678_5148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4376 a_37585_974# a_37587_875# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4377 a_17646_1342# a_17433_1342# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4378 a_20080_4939# a_20337_4749# a_19068_5120# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4379 a_14802_3984# a_14812_3241# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4380 a_16095_1003# a_16097_904# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4381 a_40342_6407# a_40540_7422# a_40491_7612# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4382 a_23114_6271# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4383 a_32772_4597# a_32559_4597# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4384 a_36293_4370# a_36550_4180# a_35284_3959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4385 gnd a_24888_1978# a_24680_1978# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4386 a_11498_2669# a_11077_2669# a_10804_2885# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4387 a_2835_4524# a_2955_6436# a_2910_6449# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4388 a_40523_1735# a_40780_1545# a_40358_2667# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4389 a_25653_1244# a_25906_1231# a_24640_1010# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4390 a_2910_6449# a_3108_7464# a_3059_7654# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4391 gnd a_40803_6861# a_40595_6861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4392 a_38053_4576# a_37840_4576# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4393 a_18872_2519# a_19070_3534# a_19025_3547# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4394 vdd d0 a_25881_6129# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4395 a_32289_3837# a_32775_3621# a_32983_3621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4396 a_28584_1305# a_28212_885# a_27620_651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4397 a_8207_2688# a_8421_1566# a_8372_1756# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4398 a_28212_885# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4399 a_19083_2184# a_20144_1813# a_20099_1826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4400 a_16072_6397# a_16070_6183# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4401 a_17986_207# a_17773_207# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4402 a_30934_1223# a_31187_1210# a_29921_989# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4403 a_7000_4287# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4404 gnd a_30107_3497# a_29899_3497# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4405 a_14786_7724# a_14782_7901# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4406 a_11282_4626# a_11069_4626# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4407 a_16772_5020# a_17576_4839# a_17735_5259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4408 a_33969_1453# a_33587_1895# a_32995_1661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4409 vdd a_19313_6890# a_19105_6890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4410 a_1880_7232# a_1837_6300# a_2045_6300# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4411 vdd a_8369_4490# a_8161_4490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4412 a_23127_3847# a_22914_3847# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4413 a_16092_1885# a_16578_1669# a_16786_1669# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4414 a_38245_7932# a_37824_7932# a_37548_8114# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4415 a_16558_5586# a_16345_5586# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4416 a_17626_5259# a_17413_5259# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4417 a_35301_1018# a_35554_1005# a_35242_1756# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4418 a_39289_2341# a_39076_2341# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4419 a_29677_6576# a_29891_5454# a_29842_5644# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4420 a_29904_3930# a_30962_4151# a_30917_4164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4421 vdd a_36562_2220# a_36354_2220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4422 vdd d0 a_41836_3178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4423 a_24599_8045# a_24856_7855# a_24553_7448# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4424 a_27596_5964# a_28400_5783# a_28569_5341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4425 vdd d0 a_36554_2784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4426 a_4143_5190# a_4396_5177# a_3130_4956# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4427 a_6722_914# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4428 a_36276_7695# a_36529_7682# a_35260_8053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4429 a_38853_4810# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4430 a_13799_3007# a_14857_3228# a_14812_3241# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4431 a_22335_2068# a_21914_2068# a_21638_1968# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4432 a_40577_1978# a_41635_2199# a_41586_2389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4433 a_3145_2020# a_3398_2007# a_3095_1600# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4434 vdd d2 a_30087_7414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4435 a_6760_3294# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4436 a_37855_1640# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4437 gnd d2 a_19270_5491# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4438 a_32274_7368# a_32755_7538# a_32963_7538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4439 gnd a_4415_845# a_4207_845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4440 a_12518_2391# a_12305_2391# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4441 a_24624_3147# a_25685_2776# a_25640_2789# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4442 a_21628_4424# a_21626_4210# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4443 a_24321_4672# a_24578_4482# a_23643_191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4444 a_11053_7982# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4445 a_10816_1520# a_10814_1306# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4446 vout a_20674_n19# a_10603_125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4447 a_28924_170# a_29651_4461# a_29602_4651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4448 vdd a_15076_853# a_14868_853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4449 a_40342_6407# a_40540_7422# a_40495_7435# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4450 a_38848_5791# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4451 vdd a_15072_2249# a_14864_2249# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4452 a_25649_1421# a_25906_1231# a_24640_1010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4453 a_16571_2648# a_16358_2648# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4454 a_2910_6449# a_3108_7464# a_3063_7477# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4455 a_17363_4839# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4456 vdd a_40768_3505# a_40560_3505# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4457 a_39269_6258# a_39056_6258# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4458 a_2044_220# a_1831_220# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4459 a_16365_1669# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4460 vdd d1 a_24881_2957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4461 a_28393_6762# a_28180_6762# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4462 gnd a_36541_5722# a_36333_5722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4463 a_28455_5222# a_28242_5222# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4464 a_8207_2688# a_8421_1566# a_8376_1579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4465 a_16085_3459# a_16083_3245# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4466 a_32793_1095# a_32580_1095# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4467 a_20064_8295# a_20067_7703# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4468 gnd d1 a_30137_7834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4469 a_8364_3539# a_8617_3526# a_8211_2511# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4470 a_9432_3212# a_9685_3199# a_8419_2978# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4471 a_29917_1166# a_30978_795# a_30929_985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4472 a_27608_2611# a_28413_2845# a_28572_3265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4473 a_33768_7772# a_33555_7772# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4474 a_30930_1400# a_31187_1210# a_29921_989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4475 a_25640_2789# a_25636_2966# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4476 a_16754_7546# a_16333_7546# a_16065_7376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4477 gnd d0 a_31149_7653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4478 a_40491_7612# a_40595_6861# a_40550_6874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4479 a_37849_3034# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4480 a_35210_7633# a_35314_6882# a_35265_7072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4481 vdd a_9672_6137# a_9464_6137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4482 a_844_1682# a_1649_1916# a_1818_1474# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4483 a_36273_8287# a_36530_8097# a_35264_7876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4484 a_11478_6586# a_11057_6586# a_10784_6802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4485 a_38257_5972# a_37836_5972# a_37560_5872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4486 a_40495_7435# a_40590_7842# a_40541_8032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4487 gnd d1 a_19345_1013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4488 gnd d0 a_15044_6730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4489 a_29677_6576# a_29891_5454# a_29846_5467# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4490 a_26919_2229# a_26919_1947# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4491 gnd a_4399_4201# a_4191_4201# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4492 a_38923_1313# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4493 a_3063_7477# a_3158_7884# a_3109_8074# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4494 a_36272_7872# a_36529_7682# a_35260_8053# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4495 a_3071_5694# a_3328_5504# a_2906_6626# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4496 gnd a_15051_5751# a_14843_5751# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4497 a_830_5033# a_1634_4852# a_1793_5272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4498 a_29697_2659# a_29954_2469# a_29602_4651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4499 a_28564_5222# a_28192_4802# a_27601_4983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4500 a_22981_1326# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4501 a_150_1898# a_636_1682# a_844_1682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4502 gnd a_36554_2784# a_36346_2784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4503 a_3109_8074# a_4170_7703# a_4121_7893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4504 gnd d2 a_40768_3505# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4505 a_16579_2084# a_16366_2084# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4506 a_8376_1579# a_8471_1986# a_8422_2176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4507 a_27615_1632# a_27194_1632# a_26921_1848# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4508 vdd d1 a_8647_7863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4509 gnd a_31155_7087# a_30947_7087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4510 a_22132_1087# a_21919_1087# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4511 gnd d0 a_9659_7682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4512 a_13591_2540# a_13789_3555# a_13740_3745# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4513 a_33949_5370# a_33567_5812# a_32975_5578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4514 a_28924_170# a_29651_4461# a_29606_4474# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4515 a_22323_4028# a_23127_3847# a_23296_3405# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4516 a_39585_178# a_39476_178# a_37394_111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4517 a_21640_1869# a_21645_1483# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4518 a_37582_2451# a_37580_2237# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4519 a_6925_2362# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4520 a_17740_5378# a_17626_5259# a_17834_5259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4521 a_12474_1363# a_12365_1363# a_12573_1363# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4522 a_35281_4935# a_35534_4922# a_35222_5673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4523 a_17433_1342# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4524 a_30897_6862# a_30909_6121# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4525 a_21620_5786# a_22106_5570# a_22314_5570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4526 a_23390_3286# a_23347_2354# a_23531_4279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4527 vdd d0 a_36534_6701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4528 a_41569_5714# a_41822_5701# a_40553_6072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4529 a_10789_5922# a_10791_5823# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4530 vdd a_31186_795# a_30978_795# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4531 a_3125_5937# a_3378_5924# a_3075_5517# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4532 a_40557_5895# a_41615_6116# a_41566_6306# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4533 vdd a_36541_5722# a_36333_5722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4534 a_38903_5230# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4535 a_25628_4923# a_25636_4185# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4536 vdd d0 a_4378_7703# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4537 a_8360_3716# a_8617_3526# a_8211_2511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4538 a_24585_1571# a_24838_1558# a_24416_2680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4539 a_32989_3055# a_32568_3055# a_32292_2955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4540 a_24604_7064# a_25665_6693# a_25620_6706# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4541 a_136_3957# a_138_3858# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4542 a_14812_3241# a_15065_3228# a_13799_3007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4543 a_4137_5756# a_4390_5743# a_3121_6114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4544 a_12459_5399# a_12077_5841# a_11485_5607# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4545 a_32983_3621# a_33788_3855# a_33957_3413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4546 vdd d1 a_40830_1965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4547 vdd d0 a_31149_7653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4548 a_32272_7154# a_32761_6972# a_32969_6972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4549 a_21882_7945# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4550 gnd d3 a_29934_6386# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4551 a_6915_4831# a_6702_4831# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4552 a_13791_4964# a_14044_4951# a_13732_5702# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4553 a_33952_3294# a_33580_2874# a_32988_2640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4554 a_4158_1035# a_162_716# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4555 vdd d0 a_15044_6730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4556 vdd d1 a_19345_1013# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4557 a_5917_1661# a_5704_1661# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4558 a_39312_7190# a_39269_6258# a_39477_6258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4559 gnd a_9664_6701# a_9456_6701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4560 a_36277_6891# a_36289_6150# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4561 vdd a_15051_5751# a_14843_5751# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4562 a_17413_5259# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4563 gnd d0 a_4395_4762# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4564 a_1806_3434# a_1424_3876# a_832_3642# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4565 a_34083_4287# a_33870_4287# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4566 a_39076_2341# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4567 a_10777_8164# a_11266_7982# a_11474_7982# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4568 a_19067_5924# a_20125_6145# a_20076_6335# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4569 a_33800_1895# a_33587_1895# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4570 a_10791_5823# a_10796_5437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4571 a_32773_5012# a_32560_5012# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4572 a_26909_3808# a_27395_3592# a_27603_3592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4573 a_3138_2999# a_3391_2986# a_3079_3737# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4574 vdd a_41836_3178# a_41628_3178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4575 a_9412_7129# a_9665_7116# a_8399_6895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4576 a_11499_3084# a_11078_3084# a_10802_2984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4577 a_12801_4316# a_12705_228# a_12913_228# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4578 vdd a_36554_2784# a_36346_2784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4579 vdd d0 a_31186_795# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4580 a_21640_2464# a_22119_2632# a_22327_2632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4581 a_8414_3959# a_8667_3946# a_8364_3539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4582 a_27604_4007# a_27183_4007# a_26907_3907# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4583 a_25643_1987# a_25900_1797# a_24631_2168# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4584 a_12553_5280# a_12498_6308# a_12706_6308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4585 a_41574_4349# a_41577_3757# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4586 vdd d0 a_9659_7682# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4587 a_13591_2540# a_13789_3555# a_13744_3568# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4588 a_30933_808# a_30929_985# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4589 gnd d0 a_9685_3199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4590 a_16083_2963# a_16085_2864# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4591 a_37553_6851# a_38042_6951# a_38250_6951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4592 a_20083_3963# a_20093_3220# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4593 a_7193_1334# a_6772_1334# a_7099_1453# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4594 a_12305_2391# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4595 a_17822_7219# a_17779_6287# a_17987_6287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4596 a_17748_3421# a_17366_3863# a_16774_3629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4597 a_838_3076# a_417_3076# a_141_3258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4598 a_23643_191# a_23534_191# a_23742_191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4599 a_19080_2986# a_19333_2973# a_19021_3724# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
C0 d3 gnd 2.53fF
C1 d2 gnd 5.06fF
C2 a_23643_191# a_23630_4279# 3.90fF
C3 a_34304_199# a_34291_4287# 3.90fF
C4 a_10603_125# a_10504_125# 5.04fF
C5 a_39585_178# a_39572_4266# 3.89fF
C6 d1 vdd 4.27fF
C7 a_7434_199# a_7421_4287# 3.89fF
C8 a_18095_207# a_18082_4295# 3.89fF
C9 vdd gnd 27.04fF
C10 d0 gnd 20.28fF
C11 a_12814_228# a_12801_4316# 3.90fF
C12 d2 vdd 2.14fF
C13 a_2153_220# a_2140_4308# 3.90fF
C14 a_28924_170# a_28911_4258# 3.89fF
C15 a_20996_n19# a_26832_103# 3.01fF
C16 d0 vdd 8.55fF
C17 d1 gnd 10.12fF
C18 gnd SUB 163.97fF
C19 a_37394_111# SUB 3.05fF
C20 vdd SUB 662.53fF
C21 a_31994_96# SUB 6.01fF
C22 d5 SUB 2.75fF
C23 a_34403_199# SUB 4.48fF
C24 a_26733_103# SUB 3.05fF
C25 a_26832_103# SUB 6.47fF
C26 a_20996_n19# SUB 12.03fF
C27 a_23742_191# SUB 4.48fF
C28 a_15904_140# SUB 3.05fF
C29 a_10504_125# SUB 6.01fF
C30 a_10603_125# SUB 12.33fF
C31 a_12913_228# SUB 4.48fF
C32 a_5243_132# SUB 3.05fF
C33 a_5342_132# SUB 6.47fF
C34 a_2252_220# SUB 4.48fF
C35 d0 SUB 82.02fF
C36 a_32313_695# SUB 6.03fF
C37 a_38281_659# SUB 2.20fF
C38 a_26933_666# SUB 6.03fF
C39 d1 SUB 42.64fF
C40 a_40578_1174# SUB 2.33fF
C41 a_38282_1074# SUB 2.33fF
C42 a_33000_680# SUB 2.20fF
C43 a_21652_687# SUB 6.03fF
C44 a_27620_651# SUB 2.20fF
C45 a_35297_1195# SUB 2.33fF
C46 a_40582_997# SUB 2.20fF
C47 a_33001_1095# SUB 2.33fF
C48 a_16104_703# SUB 6.03fF
C49 a_29917_1166# SUB 2.33fF
C50 a_27621_1066# SUB 2.33fF
C51 a_22339_672# SUB 2.20fF
C52 a_10823_724# SUB 6.03fF
C53 a_24636_1187# SUB 2.33fF
C54 a_39245_1313# SUB 2.04fF
C55 a_35301_1018# SUB 2.20fF
C56 d2 SUB 21.48fF
C57 a_33964_1334# SUB 2.04fF
C58 a_29921_989# SUB 2.20fF
C59 a_22340_1087# SUB 2.33fF
C60 a_16791_688# SUB 2.20fF
C61 a_5443_695# SUB 6.03fF
C62 a_19088_1203# SUB 2.33fF
C63 a_28584_1305# SUB 2.04fF
C64 a_24640_1010# SUB 2.20fF
C65 a_16792_1103# SUB 2.33fF
C66 a_11510_709# SUB 2.20fF
C67 a_162_716# SUB 6.03fF
C68 a_6130_680# SUB 2.20fF
C69 a_13807_1224# SUB 2.33fF
C70 a_23303_1326# SUB 2.04fF
C71 a_19092_1026# SUB 2.20fF
C72 a_11511_1124# SUB 2.33fF
C73 a_8427_1195# SUB 2.33fF
C74 a_6131_1095# SUB 2.33fF
C75 a_849_701# SUB 2.20fF
C76 a_3146_1216# SUB 2.33fF
C77 a_17755_1342# SUB 2.04fF
C78 a_13811_1047# SUB 2.20fF
C79 a_12474_1363# SUB 2.04fF
C80 a_8431_1018# SUB 2.20fF
C81 a_7094_1334# SUB 2.04fF
C82 a_3150_1039# SUB 2.20fF
C83 a_1813_1355# SUB 2.04fF
C84 a_38276_1640# SUB 2.20fF
C85 a_40527_1558# SUB 2.04fF
C86 a_40573_2155# SUB 2.33fF
C87 a_38277_2055# SUB 2.33fF
C88 a_32995_1661# SUB 2.20fF
C89 a_35246_1579# SUB 2.04fF
C90 a_27615_1632# SUB 2.20fF
C91 a_35292_2176# SUB 2.33fF
C92 a_32996_2076# SUB 2.33fF
C93 a_29866_1550# SUB 2.04fF
C94 a_29912_2147# SUB 2.33fF
C95 a_27616_2047# SUB 2.33fF
C96 a_22334_1653# SUB 2.20fF
C97 a_24585_1571# SUB 2.04fF
C98 a_24631_2168# SUB 2.33fF
C99 a_40577_1978# SUB 2.20fF
C100 a_39344_1313# SUB 2.78fF
C101 a_35296_1999# SUB 2.20fF
C102 a_22335_2068# SUB 2.33fF
C103 a_16786_1669# SUB 2.20fF
C104 a_19037_1587# SUB 2.04fF
C105 a_19083_2184# SUB 2.33fF
C106 a_29916_1970# SUB 2.20fF
C107 a_16787_2084# SUB 2.33fF
C108 a_11505_1690# SUB 2.20fF
C109 a_13756_1608# SUB 2.04fF
C110 a_6125_1661# SUB 2.20fF
C111 a_13802_2205# SUB 2.33fF
C112 d3 SUB 10.73fF
C113 a_34063_1334# SUB 2.78fF
C114 a_28683_1305# SUB 2.78fF
C115 a_24635_1991# SUB 2.20fF
C116 a_11506_2105# SUB 2.33fF
C117 a_8376_1579# SUB 2.04fF
C118 a_8422_2176# SUB 2.33fF
C119 a_6126_2076# SUB 2.33fF
C120 a_3095_1600# SUB 2.04fF
C121 a_3141_2197# SUB 2.33fF
C122 a_40358_2667# SUB 2.02fF
C123 a_35077_2688# SUB 2.02fF
C124 a_23402_1326# SUB 2.78fF
C125 a_19087_2007# SUB 2.20fF
C126 a_29697_2659# SUB 2.02fF
C127 a_17854_1342# SUB 2.78fF
C128 a_13806_2028# SUB 2.20fF
C129 a_8426_1999# SUB 2.20fF
C130 a_38269_2619# SUB 2.20fF
C131 a_24416_2680# SUB 2.02fF
C132 a_12573_1363# SUB 2.78fF
C133 a_7193_1334# SUB 2.78fF
C134 a_3145_2020# SUB 2.20fF
C135 a_40566_3134# SUB 2.33fF
C136 a_38270_3034# SUB 2.33fF
C137 a_32988_2640# SUB 2.20fF
C138 a_18868_2696# SUB 2.02fF
C139 a_27608_2611# SUB 2.20fF
C140 a_35285_3155# SUB 2.33fF
C141 a_40570_2957# SUB 2.20fF
C142 a_32989_3055# SUB 2.33fF
C143 a_13587_2717# SUB 2.02fF
C144 a_1912_1355# SUB 2.78fF
C145 a_8207_2688# SUB 2.02fF
C146 a_29905_3126# SUB 2.33fF
C147 a_27609_3026# SUB 2.33fF
C148 a_22327_2632# SUB 2.20fF
C149 a_24624_3147# SUB 2.33fF
C150 a_39233_3273# SUB 2.04fF
C151 a_39332_3273# SUB 2.02fF
C152 a_35289_2978# SUB 2.20fF
C153 a_33952_3294# SUB 2.04fF
C154 a_34051_3294# SUB 2.02fF
C155 a_29909_2949# SUB 2.20fF
C156 a_22328_3047# SUB 2.33fF
C157 a_16779_2648# SUB 2.20fF
C158 a_2926_2709# SUB 2.02fF
C159 a_19076_3163# SUB 2.33fF
C160 a_28572_3265# SUB 2.04fF
C161 a_28671_3265# SUB 2.02fF
C162 a_24628_2970# SUB 2.20fF
C163 a_16780_3063# SUB 2.33fF
C164 a_11498_2669# SUB 2.20fF
C165 a_6118_2640# SUB 2.20fF
C166 a_13795_3184# SUB 2.33fF
C167 a_23291_3286# SUB 2.04fF
C168 a_23390_3286# SUB 2.02fF
C169 a_19080_2986# SUB 2.20fF
C170 a_11499_3084# SUB 2.33fF
C171 a_8415_3155# SUB 2.33fF
C172 a_6119_3055# SUB 2.33fF
C173 a_837_2661# SUB 2.20fF
C174 a_3134_3176# SUB 2.33fF
C175 a_40362_2490# SUB 2.78fF
C176 a_17743_3302# SUB 2.04fF
C177 a_17842_3302# SUB 2.02fF
C178 a_13799_3007# SUB 2.20fF
C179 a_35081_2511# SUB 2.78fF
C180 a_29701_2482# SUB 2.78fF
C181 a_12462_3323# SUB 2.04fF
C182 a_12561_3323# SUB 2.02fF
C183 a_8419_2978# SUB 2.20fF
C184 a_7082_3294# SUB 2.04fF
C185 a_7181_3294# SUB 2.02fF
C186 a_3138_2999# SUB 2.20fF
C187 a_1801_3315# SUB 2.04fF
C188 a_1900_3315# SUB 2.02fF
C189 a_38264_3600# SUB 2.20fF
C190 a_24420_2503# SUB 2.78fF
C191 a_40515_3518# SUB 2.04fF
C192 a_40561_4115# SUB 2.33fF
C193 a_38265_4015# SUB 2.33fF
C194 a_32983_3621# SUB 2.20fF
C195 a_18872_2519# SUB 2.78fF
C196 a_35234_3539# SUB 2.04fF
C197 a_27603_3592# SUB 2.20fF
C198 a_35280_4136# SUB 2.33fF
C199 a_32984_4036# SUB 2.33fF
C200 a_29854_3510# SUB 2.04fF
C201 a_13591_2540# SUB 2.78fF
C202 a_8211_2511# SUB 2.78fF
C203 a_29900_4107# SUB 2.33fF
C204 a_27604_4007# SUB 2.33fF
C205 a_22322_3613# SUB 2.20fF
C206 a_24573_3531# SUB 2.04fF
C207 a_24619_4128# SUB 2.33fF
C208 a_40565_3938# SUB 2.20fF
C209 a_39473_4266# SUB 3.86fF
C210 a_39572_4266# SUB 4.80fF
C211 a_35284_3959# SUB 2.20fF
C212 a_22323_4028# SUB 2.33fF
C213 a_16774_3629# SUB 2.20fF
C214 a_2930_2532# SUB 2.78fF
C215 a_19025_3547# SUB 2.04fF
C216 a_19071_4144# SUB 2.33fF
C217 d4 SUB 5.73fF
C218 a_39585_178# SUB 5.58fF
C219 a_40263_4659# SUB 2.93fF
C220 a_34192_4287# SUB 3.86fF
C221 a_34291_4287# SUB 4.80fF
C222 a_29904_3930# SUB 2.20fF
C223 a_28812_4258# SUB 3.86fF
C224 a_28911_4258# SUB 4.80fF
C225 a_16775_4044# SUB 2.33fF
C226 a_11493_3650# SUB 2.20fF
C227 a_13744_3568# SUB 2.04fF
C228 a_6113_3621# SUB 2.20fF
C229 a_13790_4165# SUB 2.33fF
C230 a_24623_3951# SUB 2.20fF
C231 a_34304_199# SUB 5.58fF
C232 a_34982_4680# SUB 2.93fF
C233 a_28924_170# SUB 5.58fF
C234 a_29602_4651# SUB 2.93fF
C235 a_23531_4279# SUB 3.86fF
C236 a_23630_4279# SUB 4.80fF
C237 a_11494_4065# SUB 2.33fF
C238 a_8364_3539# SUB 2.04fF
C239 a_8410_4136# SUB 2.33fF
C240 a_6114_4036# SUB 2.33fF
C241 a_3083_3560# SUB 2.04fF
C242 a_3129_4157# SUB 2.33fF
C243 a_19075_3967# SUB 2.20fF
C244 a_38261_4576# SUB 2.20fF
C245 a_23643_191# SUB 5.58fF
C246 a_24321_4672# SUB 2.93fF
C247 a_17983_4295# SUB 3.86fF
C248 a_18082_4295# SUB 4.80fF
C249 a_13794_3988# SUB 2.20fF
C250 a_833_4057# SUB 2.33fF
C251 a_40558_5091# SUB 2.33fF
C252 a_38262_4991# SUB 2.33fF
C253 a_32980_4597# SUB 2.20fF
C254 a_18095_207# SUB 5.58fF
C255 a_18773_4688# SUB 2.93fF
C256 a_12702_4316# SUB 3.86fF
C257 a_12801_4316# SUB 4.80fF
C258 a_8414_3959# SUB 2.20fF
C259 a_7322_4287# SUB 3.86fF
C260 a_7421_4287# SUB 4.80fF
C261 a_3133_3980# SUB 2.20fF
C262 a_27600_4568# SUB 2.20fF
C263 a_35277_5112# SUB 2.33fF
C264 a_40562_4914# SUB 2.20fF
C265 a_32981_5012# SUB 2.33fF
C266 a_12814_228# SUB 5.58fF
C267 a_13492_4709# SUB 2.93fF
C268 a_7434_199# SUB 5.58fF
C269 a_8112_4680# SUB 2.93fF
C270 a_2041_4308# SUB 3.86fF
C271 a_2140_4308# SUB 4.80fF
C272 a_29897_5083# SUB 2.33fF
C273 a_27601_4983# SUB 2.33fF
C274 a_22319_4589# SUB 2.20fF
C275 a_24616_5104# SUB 2.33fF
C276 a_39225_5230# SUB 2.04fF
C277 a_35281_4935# SUB 2.20fF
C278 a_33944_5251# SUB 2.04fF
C279 a_29901_4906# SUB 2.20fF
C280 a_22320_5004# SUB 2.33fF
C281 a_16771_4605# SUB 2.20fF
C282 a_2153_220# SUB 5.58fF
C283 a_2831_4701# SUB 2.93fF
C284 a_19068_5120# SUB 2.33fF
C285 a_28564_5222# SUB 2.04fF
C286 a_24620_4927# SUB 2.20fF
C287 a_16772_5020# SUB 2.33fF
C288 a_11490_4626# SUB 2.20fF
C289 a_6110_4597# SUB 2.20fF
C290 a_13787_5141# SUB 2.33fF
C291 a_23283_5243# SUB 2.04fF
C292 a_19072_4943# SUB 2.20fF
C293 a_11491_5041# SUB 2.33fF
C294 a_8407_5112# SUB 2.33fF
C295 a_6111_5012# SUB 2.33fF
C296 a_829_4618# SUB 2.20fF
C297 a_3126_5133# SUB 2.33fF
C298 a_17735_5259# SUB 2.04fF
C299 a_13791_4964# SUB 2.20fF
C300 a_12454_5280# SUB 2.04fF
C301 a_8411_4935# SUB 2.20fF
C302 a_7074_5251# SUB 2.04fF
C303 a_3130_4956# SUB 2.20fF
C304 a_1793_5272# SUB 2.04fF
C305 a_38256_5557# SUB 2.20fF
C306 a_40507_5475# SUB 2.04fF
C307 a_40553_6072# SUB 2.33fF
C308 a_38257_5972# SUB 2.33fF
C309 a_32975_5578# SUB 2.20fF
C310 a_35226_5496# SUB 2.04fF
C311 a_27595_5549# SUB 2.20fF
C312 a_35272_6093# SUB 2.33fF
C313 a_32976_5993# SUB 2.33fF
C314 a_29846_5467# SUB 2.04fF
C315 a_29892_6064# SUB 2.33fF
C316 a_27596_5964# SUB 2.33fF
C317 a_22314_5570# SUB 2.20fF
C318 a_24565_5488# SUB 2.04fF
C319 a_24611_6085# SUB 2.33fF
C320 a_40557_5895# SUB 2.20fF
C321 a_39324_5230# SUB 2.78fF
C322 a_39477_6258# SUB 2.93fF
C323 a_35276_5916# SUB 2.20fF
C324 a_22315_5985# SUB 2.33fF
C325 a_16766_5586# SUB 2.20fF
C326 a_19017_5504# SUB 2.04fF
C327 a_19063_6101# SUB 2.33fF
C328 a_29896_5887# SUB 2.20fF
C329 a_16767_6001# SUB 2.33fF
C330 a_11485_5607# SUB 2.20fF
C331 a_13736_5525# SUB 2.04fF
C332 a_6105_5578# SUB 2.20fF
C333 a_13782_6122# SUB 2.33fF
C334 a_34043_5251# SUB 2.78fF
C335 a_34196_6279# SUB 2.93fF
C336 a_28663_5222# SUB 2.78fF
C337 a_28816_6250# SUB 2.93fF
C338 a_24615_5908# SUB 2.20fF
C339 a_11486_6022# SUB 2.33fF
C340 a_8356_5496# SUB 2.04fF
C341 a_8402_6093# SUB 2.33fF
C342 a_6106_5993# SUB 2.33fF
C343 a_3075_5517# SUB 2.04fF
C344 a_3121_6114# SUB 2.33fF
C345 a_40267_4482# SUB 3.86fF
C346 a_40338_6584# SUB 2.02fF
C347 a_34986_4503# SUB 3.86fF
C348 a_35057_6605# SUB 2.02fF
C349 a_23382_5243# SUB 2.78fF
C350 a_23535_6271# SUB 2.93fF
C351 a_19067_5924# SUB 2.20fF
C352 a_29606_4474# SUB 3.86fF
C353 a_29677_6576# SUB 2.02fF
C354 a_17834_5259# SUB 2.78fF
C355 a_17987_6287# SUB 2.93fF
C356 a_13786_5945# SUB 2.20fF
C357 a_8406_5916# SUB 2.20fF
C358 a_38249_6536# SUB 2.20fF
C359 a_24325_4495# SUB 3.86fF
C360 a_24396_6597# SUB 2.02fF
C361 a_12553_5280# SUB 2.78fF
C362 a_12706_6308# SUB 2.93fF
C363 a_7173_5251# SUB 2.78fF
C364 a_7326_6279# SUB 2.93fF
C365 a_3125_5937# SUB 2.20fF
C366 a_40546_7051# SUB 2.33fF
C367 a_38250_6951# SUB 2.33fF
C368 a_32968_6557# SUB 2.20fF
C369 a_18777_4511# SUB 3.86fF
C370 a_18848_6613# SUB 2.02fF
C371 a_27588_6528# SUB 2.20fF
C372 a_35265_7072# SUB 2.33fF
C373 a_40550_6874# SUB 2.20fF
C374 a_32969_6972# SUB 2.33fF
C375 a_13496_4532# SUB 3.86fF
C376 a_13567_6634# SUB 2.02fF
C377 a_1892_5272# SUB 2.78fF
C378 a_2045_6300# SUB 2.93fF
C379 a_8116_4503# SUB 3.86fF
C380 a_8187_6605# SUB 2.02fF
C381 a_29885_7043# SUB 2.33fF
C382 a_27589_6943# SUB 2.33fF
C383 a_22307_6549# SUB 2.20fF
C384 a_24604_7064# SUB 2.33fF
C385 a_39213_7190# SUB 2.04fF
C386 a_39312_7190# SUB 2.02fF
C387 a_35269_6895# SUB 2.20fF
C388 a_33932_7211# SUB 2.04fF
C389 a_34031_7211# SUB 2.02fF
C390 a_29889_6866# SUB 2.20fF
C391 a_22308_6964# SUB 2.33fF
C392 a_16759_6565# SUB 2.20fF
C393 a_2835_4524# SUB 3.86fF
C394 a_2906_6626# SUB 2.02fF
C395 a_19056_7080# SUB 2.33fF
C396 a_28552_7182# SUB 2.04fF
C397 a_28651_7182# SUB 2.02fF
C398 a_24608_6887# SUB 2.20fF
C399 a_16760_6980# SUB 2.33fF
C400 a_11478_6586# SUB 2.20fF
C401 a_6098_6557# SUB 2.20fF
C402 a_13775_7101# SUB 2.33fF
C403 a_23271_7203# SUB 2.04fF
C404 a_23370_7203# SUB 2.02fF
C405 a_19060_6903# SUB 2.20fF
C406 a_11479_7001# SUB 2.33fF
C407 a_8395_7072# SUB 2.33fF
C408 a_6099_6972# SUB 2.33fF
C409 a_3114_7093# SUB 2.33fF
C410 a_40342_6407# SUB 2.78fF
C411 a_17723_7219# SUB 2.04fF
C412 a_17822_7219# SUB 2.02fF
C413 a_13779_6924# SUB 2.20fF
C414 a_35061_6428# SUB 2.78fF
C415 a_29681_6399# SUB 2.78fF
C416 a_12442_7240# SUB 2.04fF
C417 a_12541_7240# SUB 2.02fF
C418 a_8399_6895# SUB 2.20fF
C419 a_818_6993# SUB 2.33fF
C420 a_7062_7211# SUB 2.04fF
C421 a_7161_7211# SUB 2.02fF
C422 a_3118_6916# SUB 2.20fF
C423 a_1781_7232# SUB 2.04fF
C424 a_1880_7232# SUB 2.02fF
C425 a_38244_7517# SUB 2.20fF
C426 a_24400_6420# SUB 2.78fF
C427 a_40495_7435# SUB 2.04fF
C428 a_40541_8032# SUB 2.33fF
C429 a_38245_7932# SUB 2.33fF
C430 a_32963_7538# SUB 2.20fF
C431 a_18852_6436# SUB 2.78fF
C432 a_35214_7456# SUB 2.04fF
C433 a_27583_7509# SUB 2.20fF
C434 a_35260_8053# SUB 2.33fF
C435 a_32964_7953# SUB 2.33fF
C436 a_29834_7427# SUB 2.04fF
C437 a_13571_6457# SUB 2.78fF
C438 a_8191_6428# SUB 2.78fF
C439 a_29880_8024# SUB 2.33fF
C440 a_27584_7924# SUB 2.33fF
C441 a_22302_7530# SUB 2.20fF
C442 a_24553_7448# SUB 2.04fF
C443 a_24599_8045# SUB 2.33fF
C444 a_40545_7855# SUB 2.20fF
C445 a_36277_8110# SUB 2.33fF
C446 a_35264_7876# SUB 2.20fF
C447 a_22303_7945# SUB 2.33fF
C448 a_16754_7546# SUB 2.20fF
C449 a_2910_6449# SUB 2.78fF
C450 a_19005_7464# SUB 2.04fF
C451 a_19051_8061# SUB 2.33fF
C452 a_29884_7847# SUB 2.20fF
C453 a_30897_8081# SUB 2.47fF
C454 a_16755_7961# SUB 2.33fF
C455 a_11473_7567# SUB 2.20fF
C456 a_13724_7485# SUB 2.04fF
C457 a_6093_7538# SUB 2.20fF
C458 a_13770_8082# SUB 2.33fF
C459 a_25616_8102# SUB 2.33fF
C460 a_24603_7868# SUB 2.20fF
C461 a_11474_7982# SUB 2.33fF
C462 a_8344_7456# SUB 2.04fF
C463 a_8390_8053# SUB 2.33fF
C464 a_6094_7953# SUB 2.33fF
C465 a_812_7559# SUB 2.20fF
C466 a_3063_7477# SUB 2.04fF
C467 a_3109_8074# SUB 2.33fF
C468 a_20068_8118# SUB 2.66fF
C469 a_19055_7884# SUB 2.20fF
C470 a_14787_8139# SUB 2.33fF
C471 a_13774_7905# SUB 2.20fF
C472 a_813_7974# SUB 2.33fF
C473 a_8394_7876# SUB 2.20fF
C474 a_4126_8131# SUB 2.33fF
C475 a_3113_7897# SUB 2.20fF
C476 vout gnd 50fF

Vdd vdd 0 dc 1.8
Vsub SUB 0 dc 0
Vin1 vref 0 dc 3.3
Vd0 d0 0 pulse(0 1.8 0 0.1ps 0.1ps 5us 10us)
Vd1 d1 0 pulse(0 1.8 0 0.1ps 0.1ps 10us 20us)
Vd2 d2 0 pulse(0 1.8 0 0.1ps 0.1ps 20us 40us)
Vd3 d3 0 pulse(0 1.8 0 0.1ps 0.1ps 40us 80us)
Vd4 d4 0 pulse(0 1.8 0 0.1ps 0.1ps 80us 160us)
Vd5 d5 0 pulse(0 1.8 0 0.1ps 0.1ps 160us 320us)
Vd6 d6 0 pulse(0 1.8 0 0.1ps 0.1ps 320us 640us)
Vd7 d7 0 pulse(0 1.8 0 0.1ps 0.1ps 640us 1280us)
Vd8 d8 0 pulse(0 1.8 0 0.1ps 0.1ps 1280us 2560us)

.tran 10us 2560us
.control
run
plot V(vout)
.endc
.end
