magic
tech sky130A
timestamp 1616158313
<< nwell >>
rect 278 1592 1089 1742
rect 1290 1411 2101 1561
rect 277 1177 1088 1327
rect 1345 850 2156 1000
rect 283 611 1094 761
rect 1295 430 2106 580
rect 282 196 1093 346
rect 1510 -82 2321 68
rect 290 -368 1101 -218
rect 1302 -549 2113 -399
rect 289 -783 1100 -633
rect 1357 -1110 2168 -960
rect 295 -1349 1106 -1199
rect 1307 -1530 2118 -1380
rect 294 -1764 1105 -1614
<< nmos >>
rect 342 1491 392 1533
rect 555 1491 605 1533
rect 763 1491 813 1533
rect 971 1491 1021 1533
rect 1354 1310 1404 1352
rect 1567 1310 1617 1352
rect 1775 1310 1825 1352
rect 1983 1310 2033 1352
rect 341 1076 391 1118
rect 554 1076 604 1118
rect 762 1076 812 1118
rect 970 1076 1020 1118
rect 1409 749 1459 791
rect 1622 749 1672 791
rect 1830 749 1880 791
rect 2038 749 2088 791
rect 347 510 397 552
rect 560 510 610 552
rect 768 510 818 552
rect 976 510 1026 552
rect 1359 329 1409 371
rect 1572 329 1622 371
rect 1780 329 1830 371
rect 1988 329 2038 371
rect 346 95 396 137
rect 559 95 609 137
rect 767 95 817 137
rect 975 95 1025 137
rect 1574 -183 1624 -141
rect 1787 -183 1837 -141
rect 1995 -183 2045 -141
rect 2203 -183 2253 -141
rect 354 -469 404 -427
rect 567 -469 617 -427
rect 775 -469 825 -427
rect 983 -469 1033 -427
rect 1366 -650 1416 -608
rect 1579 -650 1629 -608
rect 1787 -650 1837 -608
rect 1995 -650 2045 -608
rect 353 -884 403 -842
rect 566 -884 616 -842
rect 774 -884 824 -842
rect 982 -884 1032 -842
rect 1421 -1211 1471 -1169
rect 1634 -1211 1684 -1169
rect 1842 -1211 1892 -1169
rect 2050 -1211 2100 -1169
rect 359 -1450 409 -1408
rect 572 -1450 622 -1408
rect 780 -1450 830 -1408
rect 988 -1450 1038 -1408
rect 1371 -1631 1421 -1589
rect 1584 -1631 1634 -1589
rect 1792 -1631 1842 -1589
rect 2000 -1631 2050 -1589
rect 358 -1865 408 -1823
rect 571 -1865 621 -1823
rect 779 -1865 829 -1823
rect 987 -1865 1037 -1823
<< pmos >>
rect 342 1610 392 1710
rect 555 1610 605 1710
rect 763 1610 813 1710
rect 971 1610 1021 1710
rect 1354 1429 1404 1529
rect 1567 1429 1617 1529
rect 1775 1429 1825 1529
rect 1983 1429 2033 1529
rect 341 1195 391 1295
rect 554 1195 604 1295
rect 762 1195 812 1295
rect 970 1195 1020 1295
rect 1409 868 1459 968
rect 1622 868 1672 968
rect 1830 868 1880 968
rect 2038 868 2088 968
rect 347 629 397 729
rect 560 629 610 729
rect 768 629 818 729
rect 976 629 1026 729
rect 1359 448 1409 548
rect 1572 448 1622 548
rect 1780 448 1830 548
rect 1988 448 2038 548
rect 346 214 396 314
rect 559 214 609 314
rect 767 214 817 314
rect 975 214 1025 314
rect 1574 -64 1624 36
rect 1787 -64 1837 36
rect 1995 -64 2045 36
rect 2203 -64 2253 36
rect 354 -350 404 -250
rect 567 -350 617 -250
rect 775 -350 825 -250
rect 983 -350 1033 -250
rect 1366 -531 1416 -431
rect 1579 -531 1629 -431
rect 1787 -531 1837 -431
rect 1995 -531 2045 -431
rect 353 -765 403 -665
rect 566 -765 616 -665
rect 774 -765 824 -665
rect 982 -765 1032 -665
rect 1421 -1092 1471 -992
rect 1634 -1092 1684 -992
rect 1842 -1092 1892 -992
rect 2050 -1092 2100 -992
rect 359 -1331 409 -1231
rect 572 -1331 622 -1231
rect 780 -1331 830 -1231
rect 988 -1331 1038 -1231
rect 1371 -1512 1421 -1412
rect 1584 -1512 1634 -1412
rect 1792 -1512 1842 -1412
rect 2000 -1512 2050 -1412
rect 358 -1746 408 -1646
rect 571 -1746 621 -1646
rect 779 -1746 829 -1646
rect 987 -1746 1037 -1646
<< ndiff >>
rect 293 1523 342 1533
rect 293 1503 304 1523
rect 324 1503 342 1523
rect 293 1491 342 1503
rect 392 1527 436 1533
rect 392 1507 407 1527
rect 427 1507 436 1527
rect 392 1491 436 1507
rect 506 1523 555 1533
rect 506 1503 517 1523
rect 537 1503 555 1523
rect 506 1491 555 1503
rect 605 1527 649 1533
rect 605 1507 620 1527
rect 640 1507 649 1527
rect 605 1491 649 1507
rect 714 1523 763 1533
rect 714 1503 725 1523
rect 745 1503 763 1523
rect 714 1491 763 1503
rect 813 1527 857 1533
rect 813 1507 828 1527
rect 848 1507 857 1527
rect 813 1491 857 1507
rect 927 1527 971 1533
rect 927 1507 936 1527
rect 956 1507 971 1527
rect 927 1491 971 1507
rect 1021 1523 1070 1533
rect 1021 1503 1039 1523
rect 1059 1503 1070 1523
rect 1021 1491 1070 1503
rect 1305 1342 1354 1352
rect 1305 1322 1316 1342
rect 1336 1322 1354 1342
rect 1305 1310 1354 1322
rect 1404 1346 1448 1352
rect 1404 1326 1419 1346
rect 1439 1326 1448 1346
rect 1404 1310 1448 1326
rect 1518 1342 1567 1352
rect 1518 1322 1529 1342
rect 1549 1322 1567 1342
rect 1518 1310 1567 1322
rect 1617 1346 1661 1352
rect 1617 1326 1632 1346
rect 1652 1326 1661 1346
rect 1617 1310 1661 1326
rect 1726 1342 1775 1352
rect 1726 1322 1737 1342
rect 1757 1322 1775 1342
rect 1726 1310 1775 1322
rect 1825 1346 1869 1352
rect 1825 1326 1840 1346
rect 1860 1326 1869 1346
rect 1825 1310 1869 1326
rect 1939 1346 1983 1352
rect 1939 1326 1948 1346
rect 1968 1326 1983 1346
rect 1939 1310 1983 1326
rect 2033 1342 2082 1352
rect 2033 1322 2051 1342
rect 2071 1322 2082 1342
rect 2033 1310 2082 1322
rect 292 1108 341 1118
rect 292 1088 303 1108
rect 323 1088 341 1108
rect 292 1076 341 1088
rect 391 1112 435 1118
rect 391 1092 406 1112
rect 426 1092 435 1112
rect 391 1076 435 1092
rect 505 1108 554 1118
rect 505 1088 516 1108
rect 536 1088 554 1108
rect 505 1076 554 1088
rect 604 1112 648 1118
rect 604 1092 619 1112
rect 639 1092 648 1112
rect 604 1076 648 1092
rect 713 1108 762 1118
rect 713 1088 724 1108
rect 744 1088 762 1108
rect 713 1076 762 1088
rect 812 1112 856 1118
rect 812 1092 827 1112
rect 847 1092 856 1112
rect 812 1076 856 1092
rect 926 1112 970 1118
rect 926 1092 935 1112
rect 955 1092 970 1112
rect 926 1076 970 1092
rect 1020 1108 1069 1118
rect 1020 1088 1038 1108
rect 1058 1088 1069 1108
rect 1020 1076 1069 1088
rect 1360 781 1409 791
rect 1360 761 1371 781
rect 1391 761 1409 781
rect 1360 749 1409 761
rect 1459 785 1503 791
rect 1459 765 1474 785
rect 1494 765 1503 785
rect 1459 749 1503 765
rect 1573 781 1622 791
rect 1573 761 1584 781
rect 1604 761 1622 781
rect 1573 749 1622 761
rect 1672 785 1716 791
rect 1672 765 1687 785
rect 1707 765 1716 785
rect 1672 749 1716 765
rect 1781 781 1830 791
rect 1781 761 1792 781
rect 1812 761 1830 781
rect 1781 749 1830 761
rect 1880 785 1924 791
rect 1880 765 1895 785
rect 1915 765 1924 785
rect 1880 749 1924 765
rect 1994 785 2038 791
rect 1994 765 2003 785
rect 2023 765 2038 785
rect 1994 749 2038 765
rect 2088 781 2137 791
rect 2088 761 2106 781
rect 2126 761 2137 781
rect 2088 749 2137 761
rect 298 542 347 552
rect 298 522 309 542
rect 329 522 347 542
rect 298 510 347 522
rect 397 546 441 552
rect 397 526 412 546
rect 432 526 441 546
rect 397 510 441 526
rect 511 542 560 552
rect 511 522 522 542
rect 542 522 560 542
rect 511 510 560 522
rect 610 546 654 552
rect 610 526 625 546
rect 645 526 654 546
rect 610 510 654 526
rect 719 542 768 552
rect 719 522 730 542
rect 750 522 768 542
rect 719 510 768 522
rect 818 546 862 552
rect 818 526 833 546
rect 853 526 862 546
rect 818 510 862 526
rect 932 546 976 552
rect 932 526 941 546
rect 961 526 976 546
rect 932 510 976 526
rect 1026 542 1075 552
rect 1026 522 1044 542
rect 1064 522 1075 542
rect 1026 510 1075 522
rect 1310 361 1359 371
rect 1310 341 1321 361
rect 1341 341 1359 361
rect 1310 329 1359 341
rect 1409 365 1453 371
rect 1409 345 1424 365
rect 1444 345 1453 365
rect 1409 329 1453 345
rect 1523 361 1572 371
rect 1523 341 1534 361
rect 1554 341 1572 361
rect 1523 329 1572 341
rect 1622 365 1666 371
rect 1622 345 1637 365
rect 1657 345 1666 365
rect 1622 329 1666 345
rect 1731 361 1780 371
rect 1731 341 1742 361
rect 1762 341 1780 361
rect 1731 329 1780 341
rect 1830 365 1874 371
rect 1830 345 1845 365
rect 1865 345 1874 365
rect 1830 329 1874 345
rect 1944 365 1988 371
rect 1944 345 1953 365
rect 1973 345 1988 365
rect 1944 329 1988 345
rect 2038 361 2087 371
rect 2038 341 2056 361
rect 2076 341 2087 361
rect 2038 329 2087 341
rect 297 127 346 137
rect 297 107 308 127
rect 328 107 346 127
rect 297 95 346 107
rect 396 131 440 137
rect 396 111 411 131
rect 431 111 440 131
rect 396 95 440 111
rect 510 127 559 137
rect 510 107 521 127
rect 541 107 559 127
rect 510 95 559 107
rect 609 131 653 137
rect 609 111 624 131
rect 644 111 653 131
rect 609 95 653 111
rect 718 127 767 137
rect 718 107 729 127
rect 749 107 767 127
rect 718 95 767 107
rect 817 131 861 137
rect 817 111 832 131
rect 852 111 861 131
rect 817 95 861 111
rect 931 131 975 137
rect 931 111 940 131
rect 960 111 975 131
rect 931 95 975 111
rect 1025 127 1074 137
rect 1025 107 1043 127
rect 1063 107 1074 127
rect 1025 95 1074 107
rect 1525 -151 1574 -141
rect 1525 -171 1536 -151
rect 1556 -171 1574 -151
rect 1525 -183 1574 -171
rect 1624 -147 1668 -141
rect 1624 -167 1639 -147
rect 1659 -167 1668 -147
rect 1624 -183 1668 -167
rect 1738 -151 1787 -141
rect 1738 -171 1749 -151
rect 1769 -171 1787 -151
rect 1738 -183 1787 -171
rect 1837 -147 1881 -141
rect 1837 -167 1852 -147
rect 1872 -167 1881 -147
rect 1837 -183 1881 -167
rect 1946 -151 1995 -141
rect 1946 -171 1957 -151
rect 1977 -171 1995 -151
rect 1946 -183 1995 -171
rect 2045 -147 2089 -141
rect 2045 -167 2060 -147
rect 2080 -167 2089 -147
rect 2045 -183 2089 -167
rect 2159 -147 2203 -141
rect 2159 -167 2168 -147
rect 2188 -167 2203 -147
rect 2159 -183 2203 -167
rect 2253 -151 2302 -141
rect 2253 -171 2271 -151
rect 2291 -171 2302 -151
rect 2253 -183 2302 -171
rect 305 -437 354 -427
rect 305 -457 316 -437
rect 336 -457 354 -437
rect 305 -469 354 -457
rect 404 -433 448 -427
rect 404 -453 419 -433
rect 439 -453 448 -433
rect 404 -469 448 -453
rect 518 -437 567 -427
rect 518 -457 529 -437
rect 549 -457 567 -437
rect 518 -469 567 -457
rect 617 -433 661 -427
rect 617 -453 632 -433
rect 652 -453 661 -433
rect 617 -469 661 -453
rect 726 -437 775 -427
rect 726 -457 737 -437
rect 757 -457 775 -437
rect 726 -469 775 -457
rect 825 -433 869 -427
rect 825 -453 840 -433
rect 860 -453 869 -433
rect 825 -469 869 -453
rect 939 -433 983 -427
rect 939 -453 948 -433
rect 968 -453 983 -433
rect 939 -469 983 -453
rect 1033 -437 1082 -427
rect 1033 -457 1051 -437
rect 1071 -457 1082 -437
rect 1033 -469 1082 -457
rect 1317 -618 1366 -608
rect 1317 -638 1328 -618
rect 1348 -638 1366 -618
rect 1317 -650 1366 -638
rect 1416 -614 1460 -608
rect 1416 -634 1431 -614
rect 1451 -634 1460 -614
rect 1416 -650 1460 -634
rect 1530 -618 1579 -608
rect 1530 -638 1541 -618
rect 1561 -638 1579 -618
rect 1530 -650 1579 -638
rect 1629 -614 1673 -608
rect 1629 -634 1644 -614
rect 1664 -634 1673 -614
rect 1629 -650 1673 -634
rect 1738 -618 1787 -608
rect 1738 -638 1749 -618
rect 1769 -638 1787 -618
rect 1738 -650 1787 -638
rect 1837 -614 1881 -608
rect 1837 -634 1852 -614
rect 1872 -634 1881 -614
rect 1837 -650 1881 -634
rect 1951 -614 1995 -608
rect 1951 -634 1960 -614
rect 1980 -634 1995 -614
rect 1951 -650 1995 -634
rect 2045 -618 2094 -608
rect 2045 -638 2063 -618
rect 2083 -638 2094 -618
rect 2045 -650 2094 -638
rect 304 -852 353 -842
rect 304 -872 315 -852
rect 335 -872 353 -852
rect 304 -884 353 -872
rect 403 -848 447 -842
rect 403 -868 418 -848
rect 438 -868 447 -848
rect 403 -884 447 -868
rect 517 -852 566 -842
rect 517 -872 528 -852
rect 548 -872 566 -852
rect 517 -884 566 -872
rect 616 -848 660 -842
rect 616 -868 631 -848
rect 651 -868 660 -848
rect 616 -884 660 -868
rect 725 -852 774 -842
rect 725 -872 736 -852
rect 756 -872 774 -852
rect 725 -884 774 -872
rect 824 -848 868 -842
rect 824 -868 839 -848
rect 859 -868 868 -848
rect 824 -884 868 -868
rect 938 -848 982 -842
rect 938 -868 947 -848
rect 967 -868 982 -848
rect 938 -884 982 -868
rect 1032 -852 1081 -842
rect 1032 -872 1050 -852
rect 1070 -872 1081 -852
rect 1032 -884 1081 -872
rect 1372 -1179 1421 -1169
rect 1372 -1199 1383 -1179
rect 1403 -1199 1421 -1179
rect 1372 -1211 1421 -1199
rect 1471 -1175 1515 -1169
rect 1471 -1195 1486 -1175
rect 1506 -1195 1515 -1175
rect 1471 -1211 1515 -1195
rect 1585 -1179 1634 -1169
rect 1585 -1199 1596 -1179
rect 1616 -1199 1634 -1179
rect 1585 -1211 1634 -1199
rect 1684 -1175 1728 -1169
rect 1684 -1195 1699 -1175
rect 1719 -1195 1728 -1175
rect 1684 -1211 1728 -1195
rect 1793 -1179 1842 -1169
rect 1793 -1199 1804 -1179
rect 1824 -1199 1842 -1179
rect 1793 -1211 1842 -1199
rect 1892 -1175 1936 -1169
rect 1892 -1195 1907 -1175
rect 1927 -1195 1936 -1175
rect 1892 -1211 1936 -1195
rect 2006 -1175 2050 -1169
rect 2006 -1195 2015 -1175
rect 2035 -1195 2050 -1175
rect 2006 -1211 2050 -1195
rect 2100 -1179 2149 -1169
rect 2100 -1199 2118 -1179
rect 2138 -1199 2149 -1179
rect 2100 -1211 2149 -1199
rect 310 -1418 359 -1408
rect 310 -1438 321 -1418
rect 341 -1438 359 -1418
rect 310 -1450 359 -1438
rect 409 -1414 453 -1408
rect 409 -1434 424 -1414
rect 444 -1434 453 -1414
rect 409 -1450 453 -1434
rect 523 -1418 572 -1408
rect 523 -1438 534 -1418
rect 554 -1438 572 -1418
rect 523 -1450 572 -1438
rect 622 -1414 666 -1408
rect 622 -1434 637 -1414
rect 657 -1434 666 -1414
rect 622 -1450 666 -1434
rect 731 -1418 780 -1408
rect 731 -1438 742 -1418
rect 762 -1438 780 -1418
rect 731 -1450 780 -1438
rect 830 -1414 874 -1408
rect 830 -1434 845 -1414
rect 865 -1434 874 -1414
rect 830 -1450 874 -1434
rect 944 -1414 988 -1408
rect 944 -1434 953 -1414
rect 973 -1434 988 -1414
rect 944 -1450 988 -1434
rect 1038 -1418 1087 -1408
rect 1038 -1438 1056 -1418
rect 1076 -1438 1087 -1418
rect 1038 -1450 1087 -1438
rect 1322 -1599 1371 -1589
rect 1322 -1619 1333 -1599
rect 1353 -1619 1371 -1599
rect 1322 -1631 1371 -1619
rect 1421 -1595 1465 -1589
rect 1421 -1615 1436 -1595
rect 1456 -1615 1465 -1595
rect 1421 -1631 1465 -1615
rect 1535 -1599 1584 -1589
rect 1535 -1619 1546 -1599
rect 1566 -1619 1584 -1599
rect 1535 -1631 1584 -1619
rect 1634 -1595 1678 -1589
rect 1634 -1615 1649 -1595
rect 1669 -1615 1678 -1595
rect 1634 -1631 1678 -1615
rect 1743 -1599 1792 -1589
rect 1743 -1619 1754 -1599
rect 1774 -1619 1792 -1599
rect 1743 -1631 1792 -1619
rect 1842 -1595 1886 -1589
rect 1842 -1615 1857 -1595
rect 1877 -1615 1886 -1595
rect 1842 -1631 1886 -1615
rect 1956 -1595 2000 -1589
rect 1956 -1615 1965 -1595
rect 1985 -1615 2000 -1595
rect 1956 -1631 2000 -1615
rect 2050 -1599 2099 -1589
rect 2050 -1619 2068 -1599
rect 2088 -1619 2099 -1599
rect 2050 -1631 2099 -1619
rect 309 -1833 358 -1823
rect 309 -1853 320 -1833
rect 340 -1853 358 -1833
rect 309 -1865 358 -1853
rect 408 -1829 452 -1823
rect 408 -1849 423 -1829
rect 443 -1849 452 -1829
rect 408 -1865 452 -1849
rect 522 -1833 571 -1823
rect 522 -1853 533 -1833
rect 553 -1853 571 -1833
rect 522 -1865 571 -1853
rect 621 -1829 665 -1823
rect 621 -1849 636 -1829
rect 656 -1849 665 -1829
rect 621 -1865 665 -1849
rect 730 -1833 779 -1823
rect 730 -1853 741 -1833
rect 761 -1853 779 -1833
rect 730 -1865 779 -1853
rect 829 -1829 873 -1823
rect 829 -1849 844 -1829
rect 864 -1849 873 -1829
rect 829 -1865 873 -1849
rect 943 -1829 987 -1823
rect 943 -1849 952 -1829
rect 972 -1849 987 -1829
rect 943 -1865 987 -1849
rect 1037 -1833 1086 -1823
rect 1037 -1853 1055 -1833
rect 1075 -1853 1086 -1833
rect 1037 -1865 1086 -1853
<< pdiff >>
rect 298 1672 342 1710
rect 298 1652 310 1672
rect 330 1652 342 1672
rect 298 1610 342 1652
rect 392 1672 434 1710
rect 392 1652 406 1672
rect 426 1652 434 1672
rect 392 1610 434 1652
rect 511 1672 555 1710
rect 511 1652 523 1672
rect 543 1652 555 1672
rect 511 1610 555 1652
rect 605 1672 647 1710
rect 605 1652 619 1672
rect 639 1652 647 1672
rect 605 1610 647 1652
rect 719 1672 763 1710
rect 719 1652 731 1672
rect 751 1652 763 1672
rect 719 1610 763 1652
rect 813 1672 855 1710
rect 813 1652 827 1672
rect 847 1652 855 1672
rect 813 1610 855 1652
rect 929 1672 971 1710
rect 929 1652 937 1672
rect 957 1652 971 1672
rect 929 1610 971 1652
rect 1021 1679 1066 1710
rect 1021 1672 1065 1679
rect 1021 1652 1033 1672
rect 1053 1652 1065 1672
rect 1021 1610 1065 1652
rect 1310 1491 1354 1529
rect 1310 1471 1322 1491
rect 1342 1471 1354 1491
rect 1310 1429 1354 1471
rect 1404 1491 1446 1529
rect 1404 1471 1418 1491
rect 1438 1471 1446 1491
rect 1404 1429 1446 1471
rect 1523 1491 1567 1529
rect 1523 1471 1535 1491
rect 1555 1471 1567 1491
rect 1523 1429 1567 1471
rect 1617 1491 1659 1529
rect 1617 1471 1631 1491
rect 1651 1471 1659 1491
rect 1617 1429 1659 1471
rect 1731 1491 1775 1529
rect 1731 1471 1743 1491
rect 1763 1471 1775 1491
rect 1731 1429 1775 1471
rect 1825 1491 1867 1529
rect 1825 1471 1839 1491
rect 1859 1471 1867 1491
rect 1825 1429 1867 1471
rect 1941 1491 1983 1529
rect 1941 1471 1949 1491
rect 1969 1471 1983 1491
rect 1941 1429 1983 1471
rect 2033 1498 2078 1529
rect 2033 1491 2077 1498
rect 2033 1471 2045 1491
rect 2065 1471 2077 1491
rect 2033 1429 2077 1471
rect 297 1257 341 1295
rect 297 1237 309 1257
rect 329 1237 341 1257
rect 297 1195 341 1237
rect 391 1257 433 1295
rect 391 1237 405 1257
rect 425 1237 433 1257
rect 391 1195 433 1237
rect 510 1257 554 1295
rect 510 1237 522 1257
rect 542 1237 554 1257
rect 510 1195 554 1237
rect 604 1257 646 1295
rect 604 1237 618 1257
rect 638 1237 646 1257
rect 604 1195 646 1237
rect 718 1257 762 1295
rect 718 1237 730 1257
rect 750 1237 762 1257
rect 718 1195 762 1237
rect 812 1257 854 1295
rect 812 1237 826 1257
rect 846 1237 854 1257
rect 812 1195 854 1237
rect 928 1257 970 1295
rect 928 1237 936 1257
rect 956 1237 970 1257
rect 928 1195 970 1237
rect 1020 1264 1065 1295
rect 1020 1257 1064 1264
rect 1020 1237 1032 1257
rect 1052 1237 1064 1257
rect 1020 1195 1064 1237
rect 1365 930 1409 968
rect 1365 910 1377 930
rect 1397 910 1409 930
rect 1365 868 1409 910
rect 1459 930 1501 968
rect 1459 910 1473 930
rect 1493 910 1501 930
rect 1459 868 1501 910
rect 1578 930 1622 968
rect 1578 910 1590 930
rect 1610 910 1622 930
rect 1578 868 1622 910
rect 1672 930 1714 968
rect 1672 910 1686 930
rect 1706 910 1714 930
rect 1672 868 1714 910
rect 1786 930 1830 968
rect 1786 910 1798 930
rect 1818 910 1830 930
rect 1786 868 1830 910
rect 1880 930 1922 968
rect 1880 910 1894 930
rect 1914 910 1922 930
rect 1880 868 1922 910
rect 1996 930 2038 968
rect 1996 910 2004 930
rect 2024 910 2038 930
rect 1996 868 2038 910
rect 2088 937 2133 968
rect 2088 930 2132 937
rect 2088 910 2100 930
rect 2120 910 2132 930
rect 2088 868 2132 910
rect 303 691 347 729
rect 303 671 315 691
rect 335 671 347 691
rect 303 629 347 671
rect 397 691 439 729
rect 397 671 411 691
rect 431 671 439 691
rect 397 629 439 671
rect 516 691 560 729
rect 516 671 528 691
rect 548 671 560 691
rect 516 629 560 671
rect 610 691 652 729
rect 610 671 624 691
rect 644 671 652 691
rect 610 629 652 671
rect 724 691 768 729
rect 724 671 736 691
rect 756 671 768 691
rect 724 629 768 671
rect 818 691 860 729
rect 818 671 832 691
rect 852 671 860 691
rect 818 629 860 671
rect 934 691 976 729
rect 934 671 942 691
rect 962 671 976 691
rect 934 629 976 671
rect 1026 698 1071 729
rect 1026 691 1070 698
rect 1026 671 1038 691
rect 1058 671 1070 691
rect 1026 629 1070 671
rect 1315 510 1359 548
rect 1315 490 1327 510
rect 1347 490 1359 510
rect 1315 448 1359 490
rect 1409 510 1451 548
rect 1409 490 1423 510
rect 1443 490 1451 510
rect 1409 448 1451 490
rect 1528 510 1572 548
rect 1528 490 1540 510
rect 1560 490 1572 510
rect 1528 448 1572 490
rect 1622 510 1664 548
rect 1622 490 1636 510
rect 1656 490 1664 510
rect 1622 448 1664 490
rect 1736 510 1780 548
rect 1736 490 1748 510
rect 1768 490 1780 510
rect 1736 448 1780 490
rect 1830 510 1872 548
rect 1830 490 1844 510
rect 1864 490 1872 510
rect 1830 448 1872 490
rect 1946 510 1988 548
rect 1946 490 1954 510
rect 1974 490 1988 510
rect 1946 448 1988 490
rect 2038 517 2083 548
rect 2038 510 2082 517
rect 2038 490 2050 510
rect 2070 490 2082 510
rect 2038 448 2082 490
rect 302 276 346 314
rect 302 256 314 276
rect 334 256 346 276
rect 302 214 346 256
rect 396 276 438 314
rect 396 256 410 276
rect 430 256 438 276
rect 396 214 438 256
rect 515 276 559 314
rect 515 256 527 276
rect 547 256 559 276
rect 515 214 559 256
rect 609 276 651 314
rect 609 256 623 276
rect 643 256 651 276
rect 609 214 651 256
rect 723 276 767 314
rect 723 256 735 276
rect 755 256 767 276
rect 723 214 767 256
rect 817 276 859 314
rect 817 256 831 276
rect 851 256 859 276
rect 817 214 859 256
rect 933 276 975 314
rect 933 256 941 276
rect 961 256 975 276
rect 933 214 975 256
rect 1025 283 1070 314
rect 1025 276 1069 283
rect 1025 256 1037 276
rect 1057 256 1069 276
rect 1025 214 1069 256
rect 1530 -2 1574 36
rect 1530 -22 1542 -2
rect 1562 -22 1574 -2
rect 1530 -64 1574 -22
rect 1624 -2 1666 36
rect 1624 -22 1638 -2
rect 1658 -22 1666 -2
rect 1624 -64 1666 -22
rect 1743 -2 1787 36
rect 1743 -22 1755 -2
rect 1775 -22 1787 -2
rect 1743 -64 1787 -22
rect 1837 -2 1879 36
rect 1837 -22 1851 -2
rect 1871 -22 1879 -2
rect 1837 -64 1879 -22
rect 1951 -2 1995 36
rect 1951 -22 1963 -2
rect 1983 -22 1995 -2
rect 1951 -64 1995 -22
rect 2045 -2 2087 36
rect 2045 -22 2059 -2
rect 2079 -22 2087 -2
rect 2045 -64 2087 -22
rect 2161 -2 2203 36
rect 2161 -22 2169 -2
rect 2189 -22 2203 -2
rect 2161 -64 2203 -22
rect 2253 5 2298 36
rect 2253 -2 2297 5
rect 2253 -22 2265 -2
rect 2285 -22 2297 -2
rect 2253 -64 2297 -22
rect 310 -288 354 -250
rect 310 -308 322 -288
rect 342 -308 354 -288
rect 310 -350 354 -308
rect 404 -288 446 -250
rect 404 -308 418 -288
rect 438 -308 446 -288
rect 404 -350 446 -308
rect 523 -288 567 -250
rect 523 -308 535 -288
rect 555 -308 567 -288
rect 523 -350 567 -308
rect 617 -288 659 -250
rect 617 -308 631 -288
rect 651 -308 659 -288
rect 617 -350 659 -308
rect 731 -288 775 -250
rect 731 -308 743 -288
rect 763 -308 775 -288
rect 731 -350 775 -308
rect 825 -288 867 -250
rect 825 -308 839 -288
rect 859 -308 867 -288
rect 825 -350 867 -308
rect 941 -288 983 -250
rect 941 -308 949 -288
rect 969 -308 983 -288
rect 941 -350 983 -308
rect 1033 -281 1078 -250
rect 1033 -288 1077 -281
rect 1033 -308 1045 -288
rect 1065 -308 1077 -288
rect 1033 -350 1077 -308
rect 1322 -469 1366 -431
rect 1322 -489 1334 -469
rect 1354 -489 1366 -469
rect 1322 -531 1366 -489
rect 1416 -469 1458 -431
rect 1416 -489 1430 -469
rect 1450 -489 1458 -469
rect 1416 -531 1458 -489
rect 1535 -469 1579 -431
rect 1535 -489 1547 -469
rect 1567 -489 1579 -469
rect 1535 -531 1579 -489
rect 1629 -469 1671 -431
rect 1629 -489 1643 -469
rect 1663 -489 1671 -469
rect 1629 -531 1671 -489
rect 1743 -469 1787 -431
rect 1743 -489 1755 -469
rect 1775 -489 1787 -469
rect 1743 -531 1787 -489
rect 1837 -469 1879 -431
rect 1837 -489 1851 -469
rect 1871 -489 1879 -469
rect 1837 -531 1879 -489
rect 1953 -469 1995 -431
rect 1953 -489 1961 -469
rect 1981 -489 1995 -469
rect 1953 -531 1995 -489
rect 2045 -462 2090 -431
rect 2045 -469 2089 -462
rect 2045 -489 2057 -469
rect 2077 -489 2089 -469
rect 2045 -531 2089 -489
rect 309 -703 353 -665
rect 309 -723 321 -703
rect 341 -723 353 -703
rect 309 -765 353 -723
rect 403 -703 445 -665
rect 403 -723 417 -703
rect 437 -723 445 -703
rect 403 -765 445 -723
rect 522 -703 566 -665
rect 522 -723 534 -703
rect 554 -723 566 -703
rect 522 -765 566 -723
rect 616 -703 658 -665
rect 616 -723 630 -703
rect 650 -723 658 -703
rect 616 -765 658 -723
rect 730 -703 774 -665
rect 730 -723 742 -703
rect 762 -723 774 -703
rect 730 -765 774 -723
rect 824 -703 866 -665
rect 824 -723 838 -703
rect 858 -723 866 -703
rect 824 -765 866 -723
rect 940 -703 982 -665
rect 940 -723 948 -703
rect 968 -723 982 -703
rect 940 -765 982 -723
rect 1032 -696 1077 -665
rect 1032 -703 1076 -696
rect 1032 -723 1044 -703
rect 1064 -723 1076 -703
rect 1032 -765 1076 -723
rect 1377 -1030 1421 -992
rect 1377 -1050 1389 -1030
rect 1409 -1050 1421 -1030
rect 1377 -1092 1421 -1050
rect 1471 -1030 1513 -992
rect 1471 -1050 1485 -1030
rect 1505 -1050 1513 -1030
rect 1471 -1092 1513 -1050
rect 1590 -1030 1634 -992
rect 1590 -1050 1602 -1030
rect 1622 -1050 1634 -1030
rect 1590 -1092 1634 -1050
rect 1684 -1030 1726 -992
rect 1684 -1050 1698 -1030
rect 1718 -1050 1726 -1030
rect 1684 -1092 1726 -1050
rect 1798 -1030 1842 -992
rect 1798 -1050 1810 -1030
rect 1830 -1050 1842 -1030
rect 1798 -1092 1842 -1050
rect 1892 -1030 1934 -992
rect 1892 -1050 1906 -1030
rect 1926 -1050 1934 -1030
rect 1892 -1092 1934 -1050
rect 2008 -1030 2050 -992
rect 2008 -1050 2016 -1030
rect 2036 -1050 2050 -1030
rect 2008 -1092 2050 -1050
rect 2100 -1023 2145 -992
rect 2100 -1030 2144 -1023
rect 2100 -1050 2112 -1030
rect 2132 -1050 2144 -1030
rect 2100 -1092 2144 -1050
rect 315 -1269 359 -1231
rect 315 -1289 327 -1269
rect 347 -1289 359 -1269
rect 315 -1331 359 -1289
rect 409 -1269 451 -1231
rect 409 -1289 423 -1269
rect 443 -1289 451 -1269
rect 409 -1331 451 -1289
rect 528 -1269 572 -1231
rect 528 -1289 540 -1269
rect 560 -1289 572 -1269
rect 528 -1331 572 -1289
rect 622 -1269 664 -1231
rect 622 -1289 636 -1269
rect 656 -1289 664 -1269
rect 622 -1331 664 -1289
rect 736 -1269 780 -1231
rect 736 -1289 748 -1269
rect 768 -1289 780 -1269
rect 736 -1331 780 -1289
rect 830 -1269 872 -1231
rect 830 -1289 844 -1269
rect 864 -1289 872 -1269
rect 830 -1331 872 -1289
rect 946 -1269 988 -1231
rect 946 -1289 954 -1269
rect 974 -1289 988 -1269
rect 946 -1331 988 -1289
rect 1038 -1262 1083 -1231
rect 1038 -1269 1082 -1262
rect 1038 -1289 1050 -1269
rect 1070 -1289 1082 -1269
rect 1038 -1331 1082 -1289
rect 1327 -1450 1371 -1412
rect 1327 -1470 1339 -1450
rect 1359 -1470 1371 -1450
rect 1327 -1512 1371 -1470
rect 1421 -1450 1463 -1412
rect 1421 -1470 1435 -1450
rect 1455 -1470 1463 -1450
rect 1421 -1512 1463 -1470
rect 1540 -1450 1584 -1412
rect 1540 -1470 1552 -1450
rect 1572 -1470 1584 -1450
rect 1540 -1512 1584 -1470
rect 1634 -1450 1676 -1412
rect 1634 -1470 1648 -1450
rect 1668 -1470 1676 -1450
rect 1634 -1512 1676 -1470
rect 1748 -1450 1792 -1412
rect 1748 -1470 1760 -1450
rect 1780 -1470 1792 -1450
rect 1748 -1512 1792 -1470
rect 1842 -1450 1884 -1412
rect 1842 -1470 1856 -1450
rect 1876 -1470 1884 -1450
rect 1842 -1512 1884 -1470
rect 1958 -1450 2000 -1412
rect 1958 -1470 1966 -1450
rect 1986 -1470 2000 -1450
rect 1958 -1512 2000 -1470
rect 2050 -1443 2095 -1412
rect 2050 -1450 2094 -1443
rect 2050 -1470 2062 -1450
rect 2082 -1470 2094 -1450
rect 2050 -1512 2094 -1470
rect 314 -1684 358 -1646
rect 314 -1704 326 -1684
rect 346 -1704 358 -1684
rect 314 -1746 358 -1704
rect 408 -1684 450 -1646
rect 408 -1704 422 -1684
rect 442 -1704 450 -1684
rect 408 -1746 450 -1704
rect 527 -1684 571 -1646
rect 527 -1704 539 -1684
rect 559 -1704 571 -1684
rect 527 -1746 571 -1704
rect 621 -1684 663 -1646
rect 621 -1704 635 -1684
rect 655 -1704 663 -1684
rect 621 -1746 663 -1704
rect 735 -1684 779 -1646
rect 735 -1704 747 -1684
rect 767 -1704 779 -1684
rect 735 -1746 779 -1704
rect 829 -1684 871 -1646
rect 829 -1704 843 -1684
rect 863 -1704 871 -1684
rect 829 -1746 871 -1704
rect 945 -1684 987 -1646
rect 945 -1704 953 -1684
rect 973 -1704 987 -1684
rect 945 -1746 987 -1704
rect 1037 -1677 1082 -1646
rect 1037 -1684 1081 -1677
rect 1037 -1704 1049 -1684
rect 1069 -1704 1081 -1684
rect 1037 -1746 1081 -1704
<< ndiffc >>
rect 118 1887 136 1905
rect 120 1788 138 1806
rect 116 1673 134 1691
rect 118 1574 136 1592
rect 304 1503 324 1523
rect 407 1507 427 1527
rect 517 1503 537 1523
rect 620 1507 640 1527
rect 725 1503 745 1523
rect 828 1507 848 1527
rect 936 1507 956 1527
rect 1039 1503 1059 1523
rect 116 1391 134 1409
rect 1316 1322 1336 1342
rect 1419 1326 1439 1346
rect 1529 1322 1549 1342
rect 1632 1326 1652 1346
rect 1737 1322 1757 1342
rect 1840 1326 1860 1346
rect 1948 1326 1968 1346
rect 2051 1322 2071 1342
rect 118 1292 136 1310
rect 123 1190 141 1208
rect 125 1091 143 1109
rect 303 1088 323 1108
rect 406 1092 426 1112
rect 516 1088 536 1108
rect 619 1092 639 1112
rect 724 1088 744 1108
rect 827 1092 847 1112
rect 935 1092 955 1112
rect 1038 1088 1058 1108
rect 123 906 141 924
rect 125 807 143 825
rect 1371 761 1391 781
rect 1474 765 1494 785
rect 1584 761 1604 781
rect 1687 765 1707 785
rect 1792 761 1812 781
rect 1895 765 1915 785
rect 2003 765 2023 785
rect 2106 761 2126 781
rect 121 692 139 710
rect 123 593 141 611
rect 309 522 329 542
rect 412 526 432 546
rect 522 522 542 542
rect 625 526 645 546
rect 730 522 750 542
rect 833 526 853 546
rect 941 526 961 546
rect 1044 522 1064 542
rect 121 410 139 428
rect 1321 341 1341 361
rect 1424 345 1444 365
rect 1534 341 1554 361
rect 1637 345 1657 365
rect 1742 341 1762 361
rect 1845 345 1865 365
rect 1953 345 1973 365
rect 2056 341 2076 361
rect 123 311 141 329
rect 128 209 146 227
rect 130 110 148 128
rect 308 107 328 127
rect 411 111 431 131
rect 521 107 541 127
rect 624 111 644 131
rect 729 107 749 127
rect 832 111 852 131
rect 940 111 960 131
rect 1043 107 1063 127
rect 130 -73 148 -55
rect 132 -172 150 -154
rect 1536 -171 1556 -151
rect 1639 -167 1659 -147
rect 1749 -171 1769 -151
rect 1852 -167 1872 -147
rect 1957 -171 1977 -151
rect 2060 -167 2080 -147
rect 2168 -167 2188 -147
rect 2271 -171 2291 -151
rect 128 -287 146 -269
rect 130 -386 148 -368
rect 316 -457 336 -437
rect 419 -453 439 -433
rect 529 -457 549 -437
rect 632 -453 652 -433
rect 737 -457 757 -437
rect 840 -453 860 -433
rect 948 -453 968 -433
rect 1051 -457 1071 -437
rect 128 -569 146 -551
rect 1328 -638 1348 -618
rect 1431 -634 1451 -614
rect 1541 -638 1561 -618
rect 1644 -634 1664 -614
rect 1749 -638 1769 -618
rect 1852 -634 1872 -614
rect 1960 -634 1980 -614
rect 2063 -638 2083 -618
rect 130 -668 148 -650
rect 135 -770 153 -752
rect 137 -869 155 -851
rect 315 -872 335 -852
rect 418 -868 438 -848
rect 528 -872 548 -852
rect 631 -868 651 -848
rect 736 -872 756 -852
rect 839 -868 859 -848
rect 947 -868 967 -848
rect 1050 -872 1070 -852
rect 135 -1054 153 -1036
rect 137 -1153 155 -1135
rect 1383 -1199 1403 -1179
rect 1486 -1195 1506 -1175
rect 1596 -1199 1616 -1179
rect 1699 -1195 1719 -1175
rect 1804 -1199 1824 -1179
rect 1907 -1195 1927 -1175
rect 2015 -1195 2035 -1175
rect 2118 -1199 2138 -1179
rect 133 -1268 151 -1250
rect 135 -1367 153 -1349
rect 321 -1438 341 -1418
rect 424 -1434 444 -1414
rect 534 -1438 554 -1418
rect 637 -1434 657 -1414
rect 742 -1438 762 -1418
rect 845 -1434 865 -1414
rect 953 -1434 973 -1414
rect 1056 -1438 1076 -1418
rect 133 -1550 151 -1532
rect 1333 -1619 1353 -1599
rect 1436 -1615 1456 -1595
rect 1546 -1619 1566 -1599
rect 1649 -1615 1669 -1595
rect 1754 -1619 1774 -1599
rect 1857 -1615 1877 -1595
rect 1965 -1615 1985 -1595
rect 2068 -1619 2088 -1599
rect 135 -1649 153 -1631
rect 140 -1751 158 -1733
rect 142 -1850 160 -1832
rect 320 -1853 340 -1833
rect 423 -1849 443 -1829
rect 533 -1853 553 -1833
rect 636 -1849 656 -1829
rect 741 -1853 761 -1833
rect 844 -1849 864 -1829
rect 952 -1849 972 -1829
rect 1055 -1853 1075 -1833
<< pdiffc >>
rect 310 1652 330 1672
rect 406 1652 426 1672
rect 523 1652 543 1672
rect 619 1652 639 1672
rect 731 1652 751 1672
rect 827 1652 847 1672
rect 937 1652 957 1672
rect 1033 1652 1053 1672
rect 1322 1471 1342 1491
rect 1418 1471 1438 1491
rect 1535 1471 1555 1491
rect 1631 1471 1651 1491
rect 1743 1471 1763 1491
rect 1839 1471 1859 1491
rect 1949 1471 1969 1491
rect 2045 1471 2065 1491
rect 309 1237 329 1257
rect 405 1237 425 1257
rect 522 1237 542 1257
rect 618 1237 638 1257
rect 730 1237 750 1257
rect 826 1237 846 1257
rect 936 1237 956 1257
rect 1032 1237 1052 1257
rect 1377 910 1397 930
rect 1473 910 1493 930
rect 1590 910 1610 930
rect 1686 910 1706 930
rect 1798 910 1818 930
rect 1894 910 1914 930
rect 2004 910 2024 930
rect 2100 910 2120 930
rect 315 671 335 691
rect 411 671 431 691
rect 528 671 548 691
rect 624 671 644 691
rect 736 671 756 691
rect 832 671 852 691
rect 942 671 962 691
rect 1038 671 1058 691
rect 1327 490 1347 510
rect 1423 490 1443 510
rect 1540 490 1560 510
rect 1636 490 1656 510
rect 1748 490 1768 510
rect 1844 490 1864 510
rect 1954 490 1974 510
rect 2050 490 2070 510
rect 314 256 334 276
rect 410 256 430 276
rect 527 256 547 276
rect 623 256 643 276
rect 735 256 755 276
rect 831 256 851 276
rect 941 256 961 276
rect 1037 256 1057 276
rect 1542 -22 1562 -2
rect 1638 -22 1658 -2
rect 1755 -22 1775 -2
rect 1851 -22 1871 -2
rect 1963 -22 1983 -2
rect 2059 -22 2079 -2
rect 2169 -22 2189 -2
rect 2265 -22 2285 -2
rect 322 -308 342 -288
rect 418 -308 438 -288
rect 535 -308 555 -288
rect 631 -308 651 -288
rect 743 -308 763 -288
rect 839 -308 859 -288
rect 949 -308 969 -288
rect 1045 -308 1065 -288
rect 1334 -489 1354 -469
rect 1430 -489 1450 -469
rect 1547 -489 1567 -469
rect 1643 -489 1663 -469
rect 1755 -489 1775 -469
rect 1851 -489 1871 -469
rect 1961 -489 1981 -469
rect 2057 -489 2077 -469
rect 321 -723 341 -703
rect 417 -723 437 -703
rect 534 -723 554 -703
rect 630 -723 650 -703
rect 742 -723 762 -703
rect 838 -723 858 -703
rect 948 -723 968 -703
rect 1044 -723 1064 -703
rect 1389 -1050 1409 -1030
rect 1485 -1050 1505 -1030
rect 1602 -1050 1622 -1030
rect 1698 -1050 1718 -1030
rect 1810 -1050 1830 -1030
rect 1906 -1050 1926 -1030
rect 2016 -1050 2036 -1030
rect 2112 -1050 2132 -1030
rect 327 -1289 347 -1269
rect 423 -1289 443 -1269
rect 540 -1289 560 -1269
rect 636 -1289 656 -1269
rect 748 -1289 768 -1269
rect 844 -1289 864 -1269
rect 954 -1289 974 -1269
rect 1050 -1289 1070 -1269
rect 1339 -1470 1359 -1450
rect 1435 -1470 1455 -1450
rect 1552 -1470 1572 -1450
rect 1648 -1470 1668 -1450
rect 1760 -1470 1780 -1450
rect 1856 -1470 1876 -1450
rect 1966 -1470 1986 -1450
rect 2062 -1470 2082 -1450
rect 326 -1704 346 -1684
rect 422 -1704 442 -1684
rect 539 -1704 559 -1684
rect 635 -1704 655 -1684
rect 747 -1704 767 -1684
rect 843 -1704 863 -1684
rect 953 -1704 973 -1684
rect 1049 -1704 1069 -1684
<< poly >>
rect 342 1710 392 1723
rect 555 1710 605 1723
rect 763 1710 813 1723
rect 971 1710 1021 1723
rect 342 1582 392 1610
rect 342 1562 355 1582
rect 375 1562 392 1582
rect 342 1533 392 1562
rect 555 1581 605 1610
rect 555 1557 566 1581
rect 590 1557 605 1581
rect 555 1533 605 1557
rect 763 1586 813 1610
rect 763 1562 775 1586
rect 799 1562 813 1586
rect 763 1533 813 1562
rect 971 1584 1021 1610
rect 971 1558 989 1584
rect 1015 1558 1021 1584
rect 971 1533 1021 1558
rect 1354 1529 1404 1542
rect 1567 1529 1617 1542
rect 1775 1529 1825 1542
rect 1983 1529 2033 1542
rect 342 1475 392 1491
rect 555 1475 605 1491
rect 763 1475 813 1491
rect 971 1475 1021 1491
rect 1354 1401 1404 1429
rect 1354 1381 1367 1401
rect 1387 1381 1404 1401
rect 1354 1352 1404 1381
rect 1567 1400 1617 1429
rect 1567 1376 1578 1400
rect 1602 1376 1617 1400
rect 1567 1352 1617 1376
rect 1775 1405 1825 1429
rect 1775 1381 1787 1405
rect 1811 1381 1825 1405
rect 1775 1352 1825 1381
rect 1983 1403 2033 1429
rect 1983 1377 2001 1403
rect 2027 1377 2033 1403
rect 1983 1352 2033 1377
rect 341 1295 391 1308
rect 554 1295 604 1308
rect 762 1295 812 1308
rect 970 1295 1020 1308
rect 1354 1294 1404 1310
rect 1567 1294 1617 1310
rect 1775 1294 1825 1310
rect 1983 1294 2033 1310
rect 341 1167 391 1195
rect 341 1147 354 1167
rect 374 1147 391 1167
rect 341 1118 391 1147
rect 554 1166 604 1195
rect 554 1142 565 1166
rect 589 1142 604 1166
rect 554 1118 604 1142
rect 762 1171 812 1195
rect 762 1147 774 1171
rect 798 1147 812 1171
rect 762 1118 812 1147
rect 970 1169 1020 1195
rect 970 1143 988 1169
rect 1014 1143 1020 1169
rect 970 1118 1020 1143
rect 341 1060 391 1076
rect 554 1060 604 1076
rect 762 1060 812 1076
rect 970 1060 1020 1076
rect 1409 968 1459 981
rect 1622 968 1672 981
rect 1830 968 1880 981
rect 2038 968 2088 981
rect 1409 840 1459 868
rect 1409 820 1422 840
rect 1442 820 1459 840
rect 1409 791 1459 820
rect 1622 839 1672 868
rect 1622 815 1633 839
rect 1657 815 1672 839
rect 1622 791 1672 815
rect 1830 844 1880 868
rect 1830 820 1842 844
rect 1866 820 1880 844
rect 1830 791 1880 820
rect 2038 842 2088 868
rect 2038 816 2056 842
rect 2082 816 2088 842
rect 2038 791 2088 816
rect 347 729 397 742
rect 560 729 610 742
rect 768 729 818 742
rect 976 729 1026 742
rect 1409 733 1459 749
rect 1622 733 1672 749
rect 1830 733 1880 749
rect 2038 733 2088 749
rect 347 601 397 629
rect 347 581 360 601
rect 380 581 397 601
rect 347 552 397 581
rect 560 600 610 629
rect 560 576 571 600
rect 595 576 610 600
rect 560 552 610 576
rect 768 605 818 629
rect 768 581 780 605
rect 804 581 818 605
rect 768 552 818 581
rect 976 603 1026 629
rect 976 577 994 603
rect 1020 577 1026 603
rect 976 552 1026 577
rect 1359 548 1409 561
rect 1572 548 1622 561
rect 1780 548 1830 561
rect 1988 548 2038 561
rect 347 494 397 510
rect 560 494 610 510
rect 768 494 818 510
rect 976 494 1026 510
rect 1359 420 1409 448
rect 1359 400 1372 420
rect 1392 400 1409 420
rect 1359 371 1409 400
rect 1572 419 1622 448
rect 1572 395 1583 419
rect 1607 395 1622 419
rect 1572 371 1622 395
rect 1780 424 1830 448
rect 1780 400 1792 424
rect 1816 400 1830 424
rect 1780 371 1830 400
rect 1988 422 2038 448
rect 1988 396 2006 422
rect 2032 396 2038 422
rect 1988 371 2038 396
rect 346 314 396 327
rect 559 314 609 327
rect 767 314 817 327
rect 975 314 1025 327
rect 1359 313 1409 329
rect 1572 313 1622 329
rect 1780 313 1830 329
rect 1988 313 2038 329
rect 346 186 396 214
rect 346 166 359 186
rect 379 166 396 186
rect 346 137 396 166
rect 559 185 609 214
rect 559 161 570 185
rect 594 161 609 185
rect 559 137 609 161
rect 767 190 817 214
rect 767 166 779 190
rect 803 166 817 190
rect 767 137 817 166
rect 975 188 1025 214
rect 975 162 993 188
rect 1019 162 1025 188
rect 975 137 1025 162
rect 346 79 396 95
rect 559 79 609 95
rect 767 79 817 95
rect 975 79 1025 95
rect 1574 36 1624 49
rect 1787 36 1837 49
rect 1995 36 2045 49
rect 2203 36 2253 49
rect 1574 -92 1624 -64
rect 1574 -112 1587 -92
rect 1607 -112 1624 -92
rect 1574 -141 1624 -112
rect 1787 -93 1837 -64
rect 1787 -117 1798 -93
rect 1822 -117 1837 -93
rect 1787 -141 1837 -117
rect 1995 -88 2045 -64
rect 1995 -112 2007 -88
rect 2031 -112 2045 -88
rect 1995 -141 2045 -112
rect 2203 -90 2253 -64
rect 2203 -116 2221 -90
rect 2247 -116 2253 -90
rect 2203 -141 2253 -116
rect 1574 -199 1624 -183
rect 1787 -199 1837 -183
rect 1995 -199 2045 -183
rect 2203 -199 2253 -183
rect 354 -250 404 -237
rect 567 -250 617 -237
rect 775 -250 825 -237
rect 983 -250 1033 -237
rect 354 -378 404 -350
rect 354 -398 367 -378
rect 387 -398 404 -378
rect 354 -427 404 -398
rect 567 -379 617 -350
rect 567 -403 578 -379
rect 602 -403 617 -379
rect 567 -427 617 -403
rect 775 -374 825 -350
rect 775 -398 787 -374
rect 811 -398 825 -374
rect 775 -427 825 -398
rect 983 -376 1033 -350
rect 983 -402 1001 -376
rect 1027 -402 1033 -376
rect 983 -427 1033 -402
rect 1366 -431 1416 -418
rect 1579 -431 1629 -418
rect 1787 -431 1837 -418
rect 1995 -431 2045 -418
rect 354 -485 404 -469
rect 567 -485 617 -469
rect 775 -485 825 -469
rect 983 -485 1033 -469
rect 1366 -559 1416 -531
rect 1366 -579 1379 -559
rect 1399 -579 1416 -559
rect 1366 -608 1416 -579
rect 1579 -560 1629 -531
rect 1579 -584 1590 -560
rect 1614 -584 1629 -560
rect 1579 -608 1629 -584
rect 1787 -555 1837 -531
rect 1787 -579 1799 -555
rect 1823 -579 1837 -555
rect 1787 -608 1837 -579
rect 1995 -557 2045 -531
rect 1995 -583 2013 -557
rect 2039 -583 2045 -557
rect 1995 -608 2045 -583
rect 353 -665 403 -652
rect 566 -665 616 -652
rect 774 -665 824 -652
rect 982 -665 1032 -652
rect 1366 -666 1416 -650
rect 1579 -666 1629 -650
rect 1787 -666 1837 -650
rect 1995 -666 2045 -650
rect 353 -793 403 -765
rect 353 -813 366 -793
rect 386 -813 403 -793
rect 353 -842 403 -813
rect 566 -794 616 -765
rect 566 -818 577 -794
rect 601 -818 616 -794
rect 566 -842 616 -818
rect 774 -789 824 -765
rect 774 -813 786 -789
rect 810 -813 824 -789
rect 774 -842 824 -813
rect 982 -791 1032 -765
rect 982 -817 1000 -791
rect 1026 -817 1032 -791
rect 982 -842 1032 -817
rect 353 -900 403 -884
rect 566 -900 616 -884
rect 774 -900 824 -884
rect 982 -900 1032 -884
rect 1421 -992 1471 -979
rect 1634 -992 1684 -979
rect 1842 -992 1892 -979
rect 2050 -992 2100 -979
rect 1421 -1120 1471 -1092
rect 1421 -1140 1434 -1120
rect 1454 -1140 1471 -1120
rect 1421 -1169 1471 -1140
rect 1634 -1121 1684 -1092
rect 1634 -1145 1645 -1121
rect 1669 -1145 1684 -1121
rect 1634 -1169 1684 -1145
rect 1842 -1116 1892 -1092
rect 1842 -1140 1854 -1116
rect 1878 -1140 1892 -1116
rect 1842 -1169 1892 -1140
rect 2050 -1118 2100 -1092
rect 2050 -1144 2068 -1118
rect 2094 -1144 2100 -1118
rect 2050 -1169 2100 -1144
rect 359 -1231 409 -1218
rect 572 -1231 622 -1218
rect 780 -1231 830 -1218
rect 988 -1231 1038 -1218
rect 1421 -1227 1471 -1211
rect 1634 -1227 1684 -1211
rect 1842 -1227 1892 -1211
rect 2050 -1227 2100 -1211
rect 359 -1359 409 -1331
rect 359 -1379 372 -1359
rect 392 -1379 409 -1359
rect 359 -1408 409 -1379
rect 572 -1360 622 -1331
rect 572 -1384 583 -1360
rect 607 -1384 622 -1360
rect 572 -1408 622 -1384
rect 780 -1355 830 -1331
rect 780 -1379 792 -1355
rect 816 -1379 830 -1355
rect 780 -1408 830 -1379
rect 988 -1357 1038 -1331
rect 988 -1383 1006 -1357
rect 1032 -1383 1038 -1357
rect 988 -1408 1038 -1383
rect 1371 -1412 1421 -1399
rect 1584 -1412 1634 -1399
rect 1792 -1412 1842 -1399
rect 2000 -1412 2050 -1399
rect 359 -1466 409 -1450
rect 572 -1466 622 -1450
rect 780 -1466 830 -1450
rect 988 -1466 1038 -1450
rect 1371 -1540 1421 -1512
rect 1371 -1560 1384 -1540
rect 1404 -1560 1421 -1540
rect 1371 -1589 1421 -1560
rect 1584 -1541 1634 -1512
rect 1584 -1565 1595 -1541
rect 1619 -1565 1634 -1541
rect 1584 -1589 1634 -1565
rect 1792 -1536 1842 -1512
rect 1792 -1560 1804 -1536
rect 1828 -1560 1842 -1536
rect 1792 -1589 1842 -1560
rect 2000 -1538 2050 -1512
rect 2000 -1564 2018 -1538
rect 2044 -1564 2050 -1538
rect 2000 -1589 2050 -1564
rect 358 -1646 408 -1633
rect 571 -1646 621 -1633
rect 779 -1646 829 -1633
rect 987 -1646 1037 -1633
rect 1371 -1647 1421 -1631
rect 1584 -1647 1634 -1631
rect 1792 -1647 1842 -1631
rect 2000 -1647 2050 -1631
rect 358 -1774 408 -1746
rect 358 -1794 371 -1774
rect 391 -1794 408 -1774
rect 358 -1823 408 -1794
rect 571 -1775 621 -1746
rect 571 -1799 582 -1775
rect 606 -1799 621 -1775
rect 571 -1823 621 -1799
rect 779 -1770 829 -1746
rect 779 -1794 791 -1770
rect 815 -1794 829 -1770
rect 779 -1823 829 -1794
rect 987 -1772 1037 -1746
rect 987 -1798 1005 -1772
rect 1031 -1798 1037 -1772
rect 987 -1823 1037 -1798
rect 358 -1881 408 -1865
rect 571 -1881 621 -1865
rect 779 -1881 829 -1865
rect 987 -1881 1037 -1865
<< polycont >>
rect 355 1562 375 1582
rect 566 1557 590 1581
rect 775 1562 799 1586
rect 989 1558 1015 1584
rect 1367 1381 1387 1401
rect 1578 1376 1602 1400
rect 1787 1381 1811 1405
rect 2001 1377 2027 1403
rect 354 1147 374 1167
rect 565 1142 589 1166
rect 774 1147 798 1171
rect 988 1143 1014 1169
rect 1422 820 1442 840
rect 1633 815 1657 839
rect 1842 820 1866 844
rect 2056 816 2082 842
rect 360 581 380 601
rect 571 576 595 600
rect 780 581 804 605
rect 994 577 1020 603
rect 1372 400 1392 420
rect 1583 395 1607 419
rect 1792 400 1816 424
rect 2006 396 2032 422
rect 359 166 379 186
rect 570 161 594 185
rect 779 166 803 190
rect 993 162 1019 188
rect 1587 -112 1607 -92
rect 1798 -117 1822 -93
rect 2007 -112 2031 -88
rect 2221 -116 2247 -90
rect 367 -398 387 -378
rect 578 -403 602 -379
rect 787 -398 811 -374
rect 1001 -402 1027 -376
rect 1379 -579 1399 -559
rect 1590 -584 1614 -560
rect 1799 -579 1823 -555
rect 2013 -583 2039 -557
rect 366 -813 386 -793
rect 577 -818 601 -794
rect 786 -813 810 -789
rect 1000 -817 1026 -791
rect 1434 -1140 1454 -1120
rect 1645 -1145 1669 -1121
rect 1854 -1140 1878 -1116
rect 2068 -1144 2094 -1118
rect 372 -1379 392 -1359
rect 583 -1384 607 -1360
rect 792 -1379 816 -1355
rect 1006 -1383 1032 -1357
rect 1384 -1560 1404 -1540
rect 1595 -1565 1619 -1541
rect 1804 -1560 1828 -1536
rect 2018 -1564 2044 -1538
rect 371 -1794 391 -1774
rect 582 -1799 606 -1775
rect 791 -1794 815 -1770
rect 1005 -1798 1031 -1772
<< ndiffres >>
rect 97 1905 154 1924
rect 97 1902 118 1905
rect 3 1887 118 1902
rect 136 1887 154 1905
rect 3 1864 154 1887
rect 3 1828 45 1864
rect 2 1827 102 1828
rect 2 1806 158 1827
rect 2 1788 120 1806
rect 138 1788 158 1806
rect 2 1784 158 1788
rect 97 1768 158 1784
rect 95 1691 152 1710
rect 95 1688 116 1691
rect 1 1673 116 1688
rect 134 1673 152 1691
rect 1 1650 152 1673
rect 1 1614 43 1650
rect 0 1613 100 1614
rect 0 1592 156 1613
rect 0 1574 118 1592
rect 136 1574 156 1592
rect 0 1570 156 1574
rect 95 1554 156 1570
rect 95 1409 152 1428
rect 95 1406 116 1409
rect 1 1391 116 1406
rect 134 1391 152 1409
rect 1 1368 152 1391
rect 1 1332 43 1368
rect 0 1331 100 1332
rect 0 1310 156 1331
rect 0 1292 118 1310
rect 136 1292 156 1310
rect 0 1288 156 1292
rect 95 1272 156 1288
rect 102 1208 159 1227
rect 102 1205 123 1208
rect 8 1190 123 1205
rect 141 1190 159 1208
rect 8 1167 159 1190
rect 8 1131 50 1167
rect 7 1130 107 1131
rect 7 1109 163 1130
rect 7 1091 125 1109
rect 143 1091 163 1109
rect 7 1087 163 1091
rect 102 1071 163 1087
rect 102 924 159 943
rect 102 921 123 924
rect 8 906 123 921
rect 141 906 159 924
rect 8 883 159 906
rect 8 847 50 883
rect 7 846 107 847
rect 7 825 163 846
rect 7 807 125 825
rect 143 807 163 825
rect 7 803 163 807
rect 102 787 163 803
rect 100 710 157 729
rect 100 707 121 710
rect 6 692 121 707
rect 139 692 157 710
rect 6 669 157 692
rect 6 633 48 669
rect 5 632 105 633
rect 5 611 161 632
rect 5 593 123 611
rect 141 593 161 611
rect 5 589 161 593
rect 100 573 161 589
rect 100 428 157 447
rect 100 425 121 428
rect 6 410 121 425
rect 139 410 157 428
rect 6 387 157 410
rect 6 351 48 387
rect 5 350 105 351
rect 5 329 161 350
rect 5 311 123 329
rect 141 311 161 329
rect 5 307 161 311
rect 100 291 161 307
rect 107 227 164 246
rect 107 224 128 227
rect 13 209 128 224
rect 146 209 164 227
rect 13 186 164 209
rect 13 150 55 186
rect 12 149 112 150
rect 12 128 168 149
rect 12 110 130 128
rect 148 110 168 128
rect 12 106 168 110
rect 107 90 168 106
rect 109 -55 166 -36
rect 109 -58 130 -55
rect 15 -73 130 -58
rect 148 -73 166 -55
rect 15 -96 166 -73
rect 15 -132 57 -96
rect 14 -133 114 -132
rect 14 -154 170 -133
rect 14 -172 132 -154
rect 150 -172 170 -154
rect 14 -176 170 -172
rect 109 -192 170 -176
rect 107 -269 164 -250
rect 107 -272 128 -269
rect 13 -287 128 -272
rect 146 -287 164 -269
rect 13 -310 164 -287
rect 13 -346 55 -310
rect 12 -347 112 -346
rect 12 -368 168 -347
rect 12 -386 130 -368
rect 148 -386 168 -368
rect 12 -390 168 -386
rect 107 -406 168 -390
rect 107 -551 164 -532
rect 107 -554 128 -551
rect 13 -569 128 -554
rect 146 -569 164 -551
rect 13 -592 164 -569
rect 13 -628 55 -592
rect 12 -629 112 -628
rect 12 -650 168 -629
rect 12 -668 130 -650
rect 148 -668 168 -650
rect 12 -672 168 -668
rect 107 -688 168 -672
rect 114 -752 171 -733
rect 114 -755 135 -752
rect 20 -770 135 -755
rect 153 -770 171 -752
rect 20 -793 171 -770
rect 20 -829 62 -793
rect 19 -830 119 -829
rect 19 -851 175 -830
rect 19 -869 137 -851
rect 155 -869 175 -851
rect 19 -873 175 -869
rect 114 -889 175 -873
rect 114 -1036 171 -1017
rect 114 -1039 135 -1036
rect 20 -1054 135 -1039
rect 153 -1054 171 -1036
rect 20 -1077 171 -1054
rect 20 -1113 62 -1077
rect 19 -1114 119 -1113
rect 19 -1135 175 -1114
rect 19 -1153 137 -1135
rect 155 -1153 175 -1135
rect 19 -1157 175 -1153
rect 114 -1173 175 -1157
rect 112 -1250 169 -1231
rect 112 -1253 133 -1250
rect 18 -1268 133 -1253
rect 151 -1268 169 -1250
rect 18 -1291 169 -1268
rect 18 -1327 60 -1291
rect 17 -1328 117 -1327
rect 17 -1349 173 -1328
rect 17 -1367 135 -1349
rect 153 -1367 173 -1349
rect 17 -1371 173 -1367
rect 112 -1387 173 -1371
rect 112 -1532 169 -1513
rect 112 -1535 133 -1532
rect 18 -1550 133 -1535
rect 151 -1550 169 -1532
rect 18 -1573 169 -1550
rect 18 -1609 60 -1573
rect 17 -1610 117 -1609
rect 17 -1631 173 -1610
rect 17 -1649 135 -1631
rect 153 -1649 173 -1631
rect 17 -1653 173 -1649
rect 112 -1669 173 -1653
rect 119 -1733 176 -1714
rect 119 -1736 140 -1733
rect 25 -1751 140 -1736
rect 158 -1751 176 -1733
rect 25 -1774 176 -1751
rect 25 -1810 67 -1774
rect 24 -1811 124 -1810
rect 24 -1832 180 -1811
rect 24 -1850 142 -1832
rect 160 -1850 180 -1832
rect 24 -1854 180 -1850
rect 119 -1870 180 -1854
<< locali >>
rect 110 1914 145 1962
rect 108 1905 145 1914
rect 108 1887 118 1905
rect 136 1887 145 1905
rect 108 1877 145 1887
rect 111 1813 148 1815
rect 111 1812 759 1813
rect 110 1806 759 1812
rect 110 1788 120 1806
rect 138 1792 759 1806
rect 138 1788 148 1792
rect 589 1791 759 1792
rect 110 1778 148 1788
rect 110 1700 145 1778
rect 722 1768 759 1791
rect 106 1691 145 1700
rect 106 1673 116 1691
rect 134 1673 145 1691
rect 106 1667 145 1673
rect 301 1743 551 1767
rect 301 1672 338 1743
rect 453 1682 484 1683
rect 106 1663 143 1667
rect 301 1652 310 1672
rect 330 1652 338 1672
rect 301 1642 338 1652
rect 397 1672 484 1682
rect 397 1652 406 1672
rect 426 1652 484 1672
rect 397 1643 484 1652
rect 397 1642 434 1643
rect 109 1592 146 1601
rect 107 1574 118 1592
rect 136 1574 146 1592
rect 453 1590 484 1643
rect 514 1672 551 1743
rect 722 1748 1115 1768
rect 1135 1748 1138 1768
rect 722 1743 1138 1748
rect 722 1742 1063 1743
rect 666 1682 697 1683
rect 514 1652 523 1672
rect 543 1652 551 1672
rect 514 1642 551 1652
rect 610 1675 697 1682
rect 610 1672 671 1675
rect 610 1652 619 1672
rect 639 1655 671 1672
rect 692 1655 697 1675
rect 639 1652 697 1655
rect 610 1645 697 1652
rect 722 1672 759 1742
rect 1025 1741 1062 1742
rect 874 1682 910 1683
rect 722 1652 731 1672
rect 751 1652 759 1672
rect 610 1643 666 1645
rect 610 1642 647 1643
rect 722 1642 759 1652
rect 818 1672 966 1682
rect 1066 1679 1162 1681
rect 818 1652 827 1672
rect 847 1652 937 1672
rect 957 1652 966 1672
rect 818 1643 966 1652
rect 1024 1672 1162 1679
rect 1024 1652 1033 1672
rect 1053 1652 1162 1672
rect 1024 1643 1162 1652
rect 818 1642 855 1643
rect 874 1591 910 1643
rect 929 1642 966 1643
rect 1025 1642 1062 1643
rect 345 1589 386 1590
rect 107 1425 146 1574
rect 237 1582 386 1589
rect 237 1562 355 1582
rect 375 1562 386 1582
rect 237 1554 386 1562
rect 453 1586 812 1590
rect 453 1581 775 1586
rect 453 1557 566 1581
rect 590 1562 775 1581
rect 799 1562 812 1586
rect 590 1557 812 1562
rect 453 1554 812 1557
rect 874 1554 909 1591
rect 977 1588 1077 1591
rect 977 1584 1044 1588
rect 977 1558 989 1584
rect 1015 1562 1044 1584
rect 1070 1562 1077 1588
rect 1015 1558 1077 1562
rect 977 1554 1077 1558
rect 453 1533 484 1554
rect 874 1533 910 1554
rect 296 1532 333 1533
rect 295 1523 333 1532
rect 295 1503 304 1523
rect 324 1503 333 1523
rect 295 1495 333 1503
rect 399 1527 484 1533
rect 509 1532 546 1533
rect 399 1507 407 1527
rect 427 1507 484 1527
rect 399 1499 484 1507
rect 508 1523 546 1532
rect 508 1503 517 1523
rect 537 1503 546 1523
rect 399 1498 435 1499
rect 508 1495 546 1503
rect 612 1527 697 1533
rect 717 1532 754 1533
rect 612 1507 620 1527
rect 640 1526 697 1527
rect 640 1507 669 1526
rect 612 1506 669 1507
rect 690 1506 697 1526
rect 612 1499 697 1506
rect 716 1523 754 1532
rect 716 1503 725 1523
rect 745 1503 754 1523
rect 612 1498 648 1499
rect 716 1495 754 1503
rect 820 1528 964 1533
rect 820 1527 885 1528
rect 820 1507 828 1527
rect 848 1507 885 1527
rect 907 1527 964 1528
rect 907 1507 936 1527
rect 956 1507 964 1527
rect 820 1499 964 1507
rect 820 1498 856 1499
rect 928 1498 964 1499
rect 1030 1532 1067 1533
rect 1030 1531 1068 1532
rect 1030 1523 1094 1531
rect 1030 1503 1039 1523
rect 1059 1509 1094 1523
rect 1114 1509 1117 1529
rect 1059 1504 1117 1509
rect 1059 1503 1094 1504
rect 296 1466 333 1495
rect 297 1464 333 1466
rect 509 1464 546 1495
rect 297 1442 546 1464
rect 717 1463 754 1495
rect 1030 1491 1094 1503
rect 1134 1465 1161 1643
rect 993 1463 1161 1465
rect 717 1437 1161 1463
rect 1313 1562 1563 1586
rect 1313 1491 1350 1562
rect 1465 1501 1496 1502
rect 1313 1471 1322 1491
rect 1342 1471 1350 1491
rect 1313 1461 1350 1471
rect 1409 1491 1496 1501
rect 1409 1471 1418 1491
rect 1438 1471 1496 1491
rect 1409 1462 1496 1471
rect 1409 1461 1446 1462
rect 717 1427 739 1437
rect 993 1436 1161 1437
rect 677 1425 739 1427
rect 107 1418 739 1425
rect 106 1409 739 1418
rect 1465 1409 1496 1462
rect 1526 1491 1563 1562
rect 1734 1567 2127 1587
rect 2147 1567 2150 1587
rect 1734 1562 2150 1567
rect 1734 1561 2075 1562
rect 1678 1501 1709 1502
rect 1526 1471 1535 1491
rect 1555 1471 1563 1491
rect 1526 1461 1563 1471
rect 1622 1494 1709 1501
rect 1622 1491 1683 1494
rect 1622 1471 1631 1491
rect 1651 1474 1683 1491
rect 1704 1474 1709 1494
rect 1651 1471 1709 1474
rect 1622 1464 1709 1471
rect 1734 1491 1771 1561
rect 2037 1560 2074 1561
rect 1886 1501 1922 1502
rect 1734 1471 1743 1491
rect 1763 1471 1771 1491
rect 1622 1462 1678 1464
rect 1622 1461 1659 1462
rect 1734 1461 1771 1471
rect 1830 1491 1978 1501
rect 2078 1498 2174 1500
rect 1830 1471 1839 1491
rect 1859 1471 1949 1491
rect 1969 1471 1978 1491
rect 1830 1462 1978 1471
rect 2036 1491 2174 1498
rect 2036 1471 2045 1491
rect 2065 1471 2174 1491
rect 2036 1462 2174 1471
rect 1830 1461 1867 1462
rect 1886 1410 1922 1462
rect 1941 1461 1978 1462
rect 2037 1461 2074 1462
rect 106 1391 116 1409
rect 134 1408 739 1409
rect 1357 1408 1398 1409
rect 134 1403 155 1408
rect 134 1391 146 1403
rect 1249 1401 1398 1408
rect 106 1383 146 1391
rect 189 1390 215 1391
rect 106 1381 143 1383
rect 189 1372 743 1390
rect 1249 1381 1367 1401
rect 1387 1381 1398 1401
rect 1249 1373 1398 1381
rect 1465 1405 1824 1409
rect 1465 1400 1787 1405
rect 1465 1376 1578 1400
rect 1602 1381 1787 1400
rect 1811 1381 1824 1405
rect 1602 1376 1824 1381
rect 1465 1373 1824 1376
rect 1886 1373 1921 1410
rect 1989 1407 2089 1410
rect 1989 1403 2056 1407
rect 1989 1377 2001 1403
rect 2027 1381 2056 1403
rect 2082 1381 2089 1407
rect 2027 1377 2089 1381
rect 1989 1373 2089 1377
rect 109 1313 146 1319
rect 189 1313 215 1372
rect 722 1353 743 1372
rect 109 1310 215 1313
rect 109 1292 118 1310
rect 136 1296 215 1310
rect 300 1328 550 1352
rect 136 1294 212 1296
rect 136 1292 146 1294
rect 109 1282 146 1292
rect 114 1217 145 1282
rect 300 1257 337 1328
rect 452 1267 483 1268
rect 300 1237 309 1257
rect 329 1237 337 1257
rect 300 1227 337 1237
rect 396 1257 483 1267
rect 396 1237 405 1257
rect 425 1237 483 1257
rect 396 1228 483 1237
rect 396 1227 433 1228
rect 113 1208 150 1217
rect 113 1190 123 1208
rect 141 1190 150 1208
rect 113 1180 150 1190
rect 452 1175 483 1228
rect 513 1257 550 1328
rect 721 1333 1114 1353
rect 1134 1333 1137 1353
rect 1465 1352 1496 1373
rect 1886 1352 1922 1373
rect 1308 1351 1345 1352
rect 721 1328 1137 1333
rect 1307 1342 1345 1351
rect 721 1327 1062 1328
rect 665 1267 696 1268
rect 513 1237 522 1257
rect 542 1237 550 1257
rect 513 1227 550 1237
rect 609 1260 696 1267
rect 609 1257 670 1260
rect 609 1237 618 1257
rect 638 1240 670 1257
rect 691 1240 696 1260
rect 638 1237 696 1240
rect 609 1230 696 1237
rect 721 1257 758 1327
rect 1024 1326 1061 1327
rect 1307 1322 1316 1342
rect 1336 1322 1345 1342
rect 1307 1314 1345 1322
rect 1411 1346 1496 1352
rect 1521 1351 1558 1352
rect 1411 1326 1419 1346
rect 1439 1326 1496 1346
rect 1411 1318 1496 1326
rect 1520 1342 1558 1351
rect 1520 1322 1529 1342
rect 1549 1322 1558 1342
rect 1411 1317 1447 1318
rect 1520 1314 1558 1322
rect 1624 1346 1709 1352
rect 1729 1351 1766 1352
rect 1624 1326 1632 1346
rect 1652 1345 1709 1346
rect 1652 1326 1681 1345
rect 1624 1325 1681 1326
rect 1702 1325 1709 1345
rect 1624 1318 1709 1325
rect 1728 1342 1766 1351
rect 1728 1322 1737 1342
rect 1757 1322 1766 1342
rect 1624 1317 1660 1318
rect 1728 1314 1766 1322
rect 1832 1346 1976 1352
rect 1832 1326 1840 1346
rect 1860 1326 1892 1346
rect 1916 1326 1948 1346
rect 1968 1326 1976 1346
rect 1832 1318 1976 1326
rect 1832 1317 1868 1318
rect 1940 1317 1976 1318
rect 2042 1351 2079 1352
rect 2042 1350 2080 1351
rect 2042 1342 2106 1350
rect 2042 1322 2051 1342
rect 2071 1328 2106 1342
rect 2126 1328 2129 1348
rect 2071 1323 2129 1328
rect 2071 1322 2106 1323
rect 1308 1285 1345 1314
rect 1309 1283 1345 1285
rect 1521 1283 1558 1314
rect 873 1267 909 1268
rect 721 1237 730 1257
rect 750 1237 758 1257
rect 609 1228 665 1230
rect 609 1227 646 1228
rect 721 1227 758 1237
rect 817 1257 965 1267
rect 1065 1264 1161 1266
rect 817 1237 826 1257
rect 846 1237 936 1257
rect 956 1237 965 1257
rect 817 1228 965 1237
rect 1023 1257 1161 1264
rect 1309 1261 1558 1283
rect 1729 1282 1766 1314
rect 2042 1310 2106 1322
rect 2146 1284 2173 1462
rect 2005 1282 2173 1284
rect 1729 1278 2173 1282
rect 1023 1237 1032 1257
rect 1052 1237 1161 1257
rect 1729 1259 1778 1278
rect 1798 1259 2173 1278
rect 1729 1256 2173 1259
rect 2005 1255 2173 1256
rect 1023 1228 1161 1237
rect 817 1227 854 1228
rect 873 1176 909 1228
rect 928 1227 965 1228
rect 1024 1227 1061 1228
rect 344 1174 385 1175
rect 236 1167 385 1174
rect 236 1147 354 1167
rect 374 1147 385 1167
rect 236 1139 385 1147
rect 452 1171 811 1175
rect 452 1166 774 1171
rect 452 1142 565 1166
rect 589 1147 774 1166
rect 798 1147 811 1171
rect 589 1142 811 1147
rect 452 1139 811 1142
rect 873 1139 908 1176
rect 976 1173 1076 1176
rect 976 1169 1043 1173
rect 976 1143 988 1169
rect 1014 1147 1043 1169
rect 1069 1147 1076 1173
rect 1014 1143 1076 1147
rect 976 1139 1076 1143
rect 452 1118 483 1139
rect 873 1118 909 1139
rect 116 1109 153 1118
rect 295 1117 332 1118
rect 116 1091 125 1109
rect 143 1091 153 1109
rect 116 1081 153 1091
rect 117 1046 153 1081
rect 294 1108 332 1117
rect 294 1088 303 1108
rect 323 1088 332 1108
rect 294 1080 332 1088
rect 398 1112 483 1118
rect 508 1117 545 1118
rect 398 1092 406 1112
rect 426 1092 483 1112
rect 398 1084 483 1092
rect 507 1108 545 1117
rect 507 1088 516 1108
rect 536 1088 545 1108
rect 398 1083 434 1084
rect 507 1080 545 1088
rect 611 1112 696 1118
rect 716 1117 753 1118
rect 611 1092 619 1112
rect 639 1111 696 1112
rect 639 1092 668 1111
rect 611 1091 668 1092
rect 689 1091 696 1111
rect 611 1084 696 1091
rect 715 1108 753 1117
rect 715 1088 724 1108
rect 744 1088 753 1108
rect 611 1083 647 1084
rect 715 1080 753 1088
rect 819 1112 963 1118
rect 819 1092 827 1112
rect 847 1111 935 1112
rect 847 1092 875 1111
rect 819 1090 875 1092
rect 897 1092 935 1111
rect 955 1092 963 1112
rect 897 1090 963 1092
rect 819 1084 963 1090
rect 819 1083 855 1084
rect 927 1083 963 1084
rect 1029 1117 1066 1118
rect 1029 1116 1067 1117
rect 1029 1108 1093 1116
rect 1029 1088 1038 1108
rect 1058 1094 1093 1108
rect 1113 1094 1116 1114
rect 1058 1089 1116 1094
rect 1058 1088 1093 1089
rect 295 1051 332 1080
rect 115 1005 153 1046
rect 296 1049 332 1051
rect 508 1049 545 1080
rect 296 1027 545 1049
rect 716 1048 753 1080
rect 1029 1076 1093 1088
rect 1133 1050 1160 1228
rect 992 1048 1160 1050
rect 716 1022 1160 1048
rect 717 1005 741 1022
rect 992 1021 1160 1022
rect 115 987 742 1005
rect 1368 1001 1618 1025
rect 115 981 153 987
rect 115 957 152 981
rect 115 933 150 957
rect 113 924 150 933
rect 113 906 123 924
rect 141 906 150 924
rect 113 896 150 906
rect 1368 930 1405 1001
rect 1520 940 1551 941
rect 1368 910 1377 930
rect 1397 910 1405 930
rect 1368 900 1405 910
rect 1464 930 1551 940
rect 1464 910 1473 930
rect 1493 910 1551 930
rect 1464 901 1551 910
rect 1464 900 1501 901
rect 1520 848 1551 901
rect 1581 930 1618 1001
rect 1789 1006 2182 1026
rect 2202 1006 2205 1026
rect 1789 1001 2205 1006
rect 1789 1000 2130 1001
rect 1733 940 1764 941
rect 1581 910 1590 930
rect 1610 910 1618 930
rect 1581 900 1618 910
rect 1677 933 1764 940
rect 1677 930 1738 933
rect 1677 910 1686 930
rect 1706 913 1738 930
rect 1759 913 1764 933
rect 1706 910 1764 913
rect 1677 903 1764 910
rect 1789 930 1826 1000
rect 2092 999 2129 1000
rect 1941 940 1977 941
rect 1789 910 1798 930
rect 1818 910 1826 930
rect 1677 901 1733 903
rect 1677 900 1714 901
rect 1789 900 1826 910
rect 1885 930 2033 940
rect 2133 937 2229 939
rect 1885 910 1894 930
rect 1914 910 2004 930
rect 2024 910 2033 930
rect 1885 901 2033 910
rect 2091 930 2229 937
rect 2091 910 2100 930
rect 2120 910 2229 930
rect 2091 901 2229 910
rect 1885 900 1922 901
rect 1941 849 1977 901
rect 1996 900 2033 901
rect 2092 900 2129 901
rect 1412 847 1453 848
rect 1304 840 1453 847
rect 116 832 153 834
rect 116 831 764 832
rect 115 825 764 831
rect 115 807 125 825
rect 143 811 764 825
rect 1304 820 1422 840
rect 1442 820 1453 840
rect 1304 812 1453 820
rect 1520 844 1879 848
rect 1520 839 1842 844
rect 1520 815 1633 839
rect 1657 820 1842 839
rect 1866 820 1879 844
rect 1657 815 1879 820
rect 1520 812 1879 815
rect 1941 812 1976 849
rect 2044 846 2144 849
rect 2044 842 2111 846
rect 2044 816 2056 842
rect 2082 820 2111 842
rect 2137 820 2144 846
rect 2082 816 2144 820
rect 2044 812 2144 816
rect 143 807 153 811
rect 594 810 764 811
rect 115 797 153 807
rect 115 719 150 797
rect 727 787 764 810
rect 1520 791 1551 812
rect 1941 791 1977 812
rect 1363 790 1400 791
rect 111 710 150 719
rect 111 692 121 710
rect 139 692 150 710
rect 111 686 150 692
rect 306 762 556 786
rect 306 691 343 762
rect 458 701 489 702
rect 111 682 148 686
rect 306 671 315 691
rect 335 671 343 691
rect 306 661 343 671
rect 402 691 489 701
rect 402 671 411 691
rect 431 671 489 691
rect 402 662 489 671
rect 402 661 439 662
rect 114 611 151 620
rect 112 593 123 611
rect 141 593 151 611
rect 458 609 489 662
rect 519 691 556 762
rect 727 767 1120 787
rect 1140 767 1143 787
rect 727 762 1143 767
rect 1362 781 1400 790
rect 727 761 1068 762
rect 1362 761 1371 781
rect 1391 761 1400 781
rect 671 701 702 702
rect 519 671 528 691
rect 548 671 556 691
rect 519 661 556 671
rect 615 694 702 701
rect 615 691 676 694
rect 615 671 624 691
rect 644 674 676 691
rect 697 674 702 694
rect 644 671 702 674
rect 615 664 702 671
rect 727 691 764 761
rect 1030 760 1067 761
rect 1362 753 1400 761
rect 1466 785 1551 791
rect 1576 790 1613 791
rect 1466 765 1474 785
rect 1494 765 1551 785
rect 1466 757 1551 765
rect 1575 781 1613 790
rect 1575 761 1584 781
rect 1604 761 1613 781
rect 1466 756 1502 757
rect 1575 753 1613 761
rect 1679 785 1764 791
rect 1784 790 1821 791
rect 1679 765 1687 785
rect 1707 784 1764 785
rect 1707 765 1736 784
rect 1679 764 1736 765
rect 1757 764 1764 784
rect 1679 757 1764 764
rect 1783 781 1821 790
rect 1783 761 1792 781
rect 1812 761 1821 781
rect 1679 756 1715 757
rect 1783 753 1821 761
rect 1887 785 2031 791
rect 1887 765 1895 785
rect 1915 783 2003 785
rect 1915 766 1951 783
rect 1975 766 2003 783
rect 1915 765 2003 766
rect 2023 765 2031 785
rect 1887 757 2031 765
rect 1887 756 1923 757
rect 1995 756 2031 757
rect 2097 790 2134 791
rect 2097 789 2135 790
rect 2097 781 2161 789
rect 2097 761 2106 781
rect 2126 767 2161 781
rect 2181 767 2184 787
rect 2126 762 2184 767
rect 2126 761 2161 762
rect 1363 724 1400 753
rect 1364 722 1400 724
rect 1576 722 1613 753
rect 879 701 915 702
rect 727 671 736 691
rect 756 671 764 691
rect 615 662 671 664
rect 615 661 652 662
rect 727 661 764 671
rect 823 691 971 701
rect 1364 700 1613 722
rect 1784 721 1821 753
rect 2097 749 2161 761
rect 2201 723 2228 901
rect 2060 721 2228 723
rect 1784 710 2228 721
rect 1071 698 1167 700
rect 823 671 832 691
rect 852 671 942 691
rect 962 671 971 691
rect 823 662 971 671
rect 1029 691 1167 698
rect 1784 695 2230 710
rect 2060 694 2230 695
rect 1029 671 1038 691
rect 1058 671 1167 691
rect 1029 662 1167 671
rect 823 661 860 662
rect 879 610 915 662
rect 934 661 971 662
rect 1030 661 1067 662
rect 350 608 391 609
rect 112 444 151 593
rect 242 601 391 608
rect 242 581 360 601
rect 380 581 391 601
rect 242 573 391 581
rect 458 605 817 609
rect 458 600 780 605
rect 458 576 571 600
rect 595 581 780 600
rect 804 581 817 605
rect 595 576 817 581
rect 458 573 817 576
rect 879 573 914 610
rect 982 607 1082 610
rect 982 603 1049 607
rect 982 577 994 603
rect 1020 581 1049 603
rect 1075 581 1082 607
rect 1020 577 1082 581
rect 982 573 1082 577
rect 458 552 489 573
rect 879 552 915 573
rect 301 551 338 552
rect 300 542 338 551
rect 300 522 309 542
rect 329 522 338 542
rect 300 514 338 522
rect 404 546 489 552
rect 514 551 551 552
rect 404 526 412 546
rect 432 526 489 546
rect 404 518 489 526
rect 513 542 551 551
rect 513 522 522 542
rect 542 522 551 542
rect 404 517 440 518
rect 513 514 551 522
rect 617 546 702 552
rect 722 551 759 552
rect 617 526 625 546
rect 645 545 702 546
rect 645 526 674 545
rect 617 525 674 526
rect 695 525 702 545
rect 617 518 702 525
rect 721 542 759 551
rect 721 522 730 542
rect 750 522 759 542
rect 617 517 653 518
rect 721 514 759 522
rect 825 547 969 552
rect 825 546 890 547
rect 825 526 833 546
rect 853 526 890 546
rect 912 546 969 547
rect 912 526 941 546
rect 961 526 969 546
rect 825 518 969 526
rect 825 517 861 518
rect 933 517 969 518
rect 1035 551 1072 552
rect 1035 550 1073 551
rect 1035 542 1099 550
rect 1035 522 1044 542
rect 1064 528 1099 542
rect 1119 528 1122 548
rect 1064 523 1122 528
rect 1064 522 1099 523
rect 301 485 338 514
rect 302 483 338 485
rect 514 483 551 514
rect 302 461 551 483
rect 722 482 759 514
rect 1035 510 1099 522
rect 1139 484 1166 662
rect 998 482 1166 484
rect 722 456 1166 482
rect 1318 581 1568 605
rect 1318 510 1355 581
rect 1470 520 1501 521
rect 1318 490 1327 510
rect 1347 490 1355 510
rect 1318 480 1355 490
rect 1414 510 1501 520
rect 1414 490 1423 510
rect 1443 490 1501 510
rect 1414 481 1501 490
rect 1414 480 1451 481
rect 722 446 744 456
rect 998 455 1166 456
rect 682 444 744 446
rect 112 437 744 444
rect 111 428 744 437
rect 1470 428 1501 481
rect 1531 510 1568 581
rect 1739 586 2132 606
rect 2152 586 2155 606
rect 1739 581 2155 586
rect 1739 580 2080 581
rect 1683 520 1714 521
rect 1531 490 1540 510
rect 1560 490 1568 510
rect 1531 480 1568 490
rect 1627 513 1714 520
rect 1627 510 1688 513
rect 1627 490 1636 510
rect 1656 493 1688 510
rect 1709 493 1714 513
rect 1656 490 1714 493
rect 1627 483 1714 490
rect 1739 510 1776 580
rect 2042 579 2079 580
rect 1891 520 1927 521
rect 1739 490 1748 510
rect 1768 490 1776 510
rect 1627 481 1683 483
rect 1627 480 1664 481
rect 1739 480 1776 490
rect 1835 510 1983 520
rect 2083 517 2179 519
rect 1835 490 1844 510
rect 1864 490 1954 510
rect 1974 490 1983 510
rect 1835 481 1983 490
rect 2041 510 2179 517
rect 2041 490 2050 510
rect 2070 490 2179 510
rect 2041 481 2179 490
rect 1835 480 1872 481
rect 1891 429 1927 481
rect 1946 480 1983 481
rect 2042 480 2079 481
rect 111 410 121 428
rect 139 427 744 428
rect 1362 427 1403 428
rect 139 422 160 427
rect 139 410 151 422
rect 1254 420 1403 427
rect 111 402 151 410
rect 194 409 220 410
rect 111 400 148 402
rect 194 391 748 409
rect 1254 400 1372 420
rect 1392 400 1403 420
rect 1254 392 1403 400
rect 1470 424 1829 428
rect 1470 419 1792 424
rect 1470 395 1583 419
rect 1607 400 1792 419
rect 1816 400 1829 424
rect 1607 395 1829 400
rect 1470 392 1829 395
rect 1891 392 1926 429
rect 1994 426 2094 429
rect 1994 422 2061 426
rect 1994 396 2006 422
rect 2032 400 2061 422
rect 2087 400 2094 426
rect 2032 396 2094 400
rect 1994 392 2094 396
rect 114 332 151 338
rect 194 332 220 391
rect 727 372 748 391
rect 114 329 220 332
rect 114 311 123 329
rect 141 315 220 329
rect 305 347 555 371
rect 141 313 217 315
rect 141 311 151 313
rect 114 301 151 311
rect 119 236 150 301
rect 305 276 342 347
rect 457 286 488 287
rect 305 256 314 276
rect 334 256 342 276
rect 305 246 342 256
rect 401 276 488 286
rect 401 256 410 276
rect 430 256 488 276
rect 401 247 488 256
rect 401 246 438 247
rect 118 227 155 236
rect 118 209 128 227
rect 146 209 155 227
rect 118 199 155 209
rect 457 194 488 247
rect 518 276 555 347
rect 726 352 1119 372
rect 1139 352 1142 372
rect 1470 371 1501 392
rect 1891 371 1927 392
rect 1313 370 1350 371
rect 726 347 1142 352
rect 1312 361 1350 370
rect 726 346 1067 347
rect 670 286 701 287
rect 518 256 527 276
rect 547 256 555 276
rect 518 246 555 256
rect 614 279 701 286
rect 614 276 675 279
rect 614 256 623 276
rect 643 259 675 276
rect 696 259 701 279
rect 643 256 701 259
rect 614 249 701 256
rect 726 276 763 346
rect 1029 345 1066 346
rect 1312 341 1321 361
rect 1341 341 1350 361
rect 1312 333 1350 341
rect 1416 365 1501 371
rect 1526 370 1563 371
rect 1416 345 1424 365
rect 1444 345 1501 365
rect 1416 337 1501 345
rect 1525 361 1563 370
rect 1525 341 1534 361
rect 1554 341 1563 361
rect 1416 336 1452 337
rect 1525 333 1563 341
rect 1629 365 1714 371
rect 1734 370 1771 371
rect 1629 345 1637 365
rect 1657 364 1714 365
rect 1657 345 1686 364
rect 1629 344 1686 345
rect 1707 344 1714 364
rect 1629 337 1714 344
rect 1733 361 1771 370
rect 1733 341 1742 361
rect 1762 341 1771 361
rect 1629 336 1665 337
rect 1733 333 1771 341
rect 1837 366 1981 371
rect 1837 365 1896 366
rect 1837 345 1845 365
rect 1865 346 1896 365
rect 1920 365 1981 366
rect 1920 346 1953 365
rect 1865 345 1953 346
rect 1973 345 1981 365
rect 1837 337 1981 345
rect 1837 336 1873 337
rect 1945 336 1981 337
rect 2047 370 2084 371
rect 2047 369 2085 370
rect 2047 361 2111 369
rect 2047 341 2056 361
rect 2076 347 2111 361
rect 2131 347 2134 367
rect 2076 342 2134 347
rect 2076 341 2111 342
rect 1313 304 1350 333
rect 1314 302 1350 304
rect 1526 302 1563 333
rect 878 286 914 287
rect 726 256 735 276
rect 755 256 763 276
rect 614 247 670 249
rect 614 246 651 247
rect 726 246 763 256
rect 822 276 970 286
rect 1070 283 1166 285
rect 822 256 831 276
rect 851 256 941 276
rect 961 256 970 276
rect 822 247 970 256
rect 1028 276 1166 283
rect 1314 280 1563 302
rect 1734 301 1771 333
rect 2047 329 2111 341
rect 2151 303 2178 481
rect 2010 301 2178 303
rect 1734 297 2178 301
rect 1028 256 1037 276
rect 1057 256 1166 276
rect 1734 278 1783 297
rect 1803 278 2178 297
rect 1734 275 2178 278
rect 2010 274 2178 275
rect 2199 300 2230 694
rect 2199 274 2204 300
rect 2223 274 2230 300
rect 2199 271 2230 274
rect 1028 247 1166 256
rect 822 246 859 247
rect 878 195 914 247
rect 933 246 970 247
rect 1029 246 1066 247
rect 349 193 390 194
rect 241 186 390 193
rect 241 166 359 186
rect 379 166 390 186
rect 241 158 390 166
rect 457 190 816 194
rect 457 185 779 190
rect 457 161 570 185
rect 594 166 779 185
rect 803 166 816 190
rect 594 161 816 166
rect 457 158 816 161
rect 878 158 913 195
rect 981 192 1081 195
rect 981 188 1048 192
rect 981 162 993 188
rect 1019 166 1048 188
rect 1074 166 1081 192
rect 1019 162 1081 166
rect 981 158 1081 162
rect 457 137 488 158
rect 878 137 914 158
rect 121 128 158 137
rect 300 136 337 137
rect 121 110 130 128
rect 148 110 158 128
rect 121 100 158 110
rect 122 65 158 100
rect 299 127 337 136
rect 299 107 308 127
rect 328 107 337 127
rect 299 99 337 107
rect 403 131 488 137
rect 513 136 550 137
rect 403 111 411 131
rect 431 111 488 131
rect 403 103 488 111
rect 512 127 550 136
rect 512 107 521 127
rect 541 107 550 127
rect 403 102 439 103
rect 512 99 550 107
rect 616 131 701 137
rect 721 136 758 137
rect 616 111 624 131
rect 644 130 701 131
rect 644 111 673 130
rect 616 110 673 111
rect 694 110 701 130
rect 616 103 701 110
rect 720 127 758 136
rect 720 107 729 127
rect 749 107 758 127
rect 616 102 652 103
rect 720 99 758 107
rect 824 131 968 137
rect 824 111 832 131
rect 852 130 940 131
rect 852 111 880 130
rect 824 109 880 111
rect 902 111 940 130
rect 960 111 968 131
rect 902 109 968 111
rect 824 103 968 109
rect 824 102 860 103
rect 932 102 968 103
rect 1034 136 1071 137
rect 1034 135 1072 136
rect 1034 127 1098 135
rect 1034 107 1043 127
rect 1063 113 1098 127
rect 1118 113 1121 133
rect 1063 108 1121 113
rect 1063 107 1098 108
rect 300 70 337 99
rect 120 24 158 65
rect 301 68 337 70
rect 513 68 550 99
rect 301 46 550 68
rect 721 67 758 99
rect 1034 95 1098 107
rect 1138 69 1165 247
rect 997 67 1165 69
rect 721 41 1165 67
rect 722 24 746 41
rect 997 40 1165 41
rect 1533 69 1783 93
rect 120 6 747 24
rect 120 0 158 6
rect 122 -46 157 0
rect 1533 -2 1570 69
rect 1685 8 1716 9
rect 1533 -22 1542 -2
rect 1562 -22 1570 -2
rect 1533 -32 1570 -22
rect 1629 -2 1716 8
rect 1629 -22 1638 -2
rect 1658 -22 1716 -2
rect 1629 -31 1716 -22
rect 1629 -32 1666 -31
rect 120 -55 157 -46
rect 120 -73 130 -55
rect 148 -73 157 -55
rect 120 -83 157 -73
rect 1685 -84 1716 -31
rect 1746 -2 1783 69
rect 1954 74 2347 94
rect 2367 74 2370 94
rect 1954 69 2370 74
rect 1954 68 2295 69
rect 1898 8 1929 9
rect 1746 -22 1755 -2
rect 1775 -22 1783 -2
rect 1746 -32 1783 -22
rect 1842 1 1929 8
rect 1842 -2 1903 1
rect 1842 -22 1851 -2
rect 1871 -19 1903 -2
rect 1924 -19 1929 1
rect 1871 -22 1929 -19
rect 1842 -29 1929 -22
rect 1954 -2 1991 68
rect 2257 67 2294 68
rect 2106 8 2142 9
rect 1954 -22 1963 -2
rect 1983 -22 1991 -2
rect 1842 -31 1898 -29
rect 1842 -32 1879 -31
rect 1954 -32 1991 -22
rect 2050 -2 2198 8
rect 2298 5 2394 7
rect 2050 -22 2059 -2
rect 2079 -22 2169 -2
rect 2189 -22 2198 -2
rect 2050 -31 2198 -22
rect 2256 -2 2394 5
rect 2256 -22 2265 -2
rect 2285 -22 2394 -2
rect 2256 -31 2394 -22
rect 2050 -32 2087 -31
rect 2106 -83 2142 -31
rect 2161 -32 2198 -31
rect 2257 -32 2294 -31
rect 1577 -85 1618 -84
rect 1469 -92 1618 -85
rect 1469 -112 1587 -92
rect 1607 -112 1618 -92
rect 1469 -120 1618 -112
rect 1685 -88 2044 -84
rect 1685 -93 2007 -88
rect 1685 -117 1798 -93
rect 1822 -112 2007 -93
rect 2031 -112 2044 -88
rect 1822 -117 2044 -112
rect 1685 -120 2044 -117
rect 2106 -120 2141 -83
rect 2209 -86 2309 -83
rect 2209 -90 2276 -86
rect 2209 -116 2221 -90
rect 2247 -112 2276 -90
rect 2302 -112 2309 -86
rect 2247 -116 2309 -112
rect 2209 -120 2309 -116
rect 1685 -141 1716 -120
rect 2106 -141 2142 -120
rect 1528 -142 1565 -141
rect 123 -147 160 -145
rect 123 -148 771 -147
rect 122 -154 771 -148
rect 122 -172 132 -154
rect 150 -168 771 -154
rect 150 -172 160 -168
rect 601 -169 771 -168
rect 122 -182 160 -172
rect 122 -260 157 -182
rect 734 -192 771 -169
rect 1527 -151 1565 -142
rect 1527 -171 1536 -151
rect 1556 -171 1565 -151
rect 1527 -179 1565 -171
rect 1631 -147 1716 -141
rect 1741 -142 1778 -141
rect 1631 -167 1639 -147
rect 1659 -167 1716 -147
rect 1631 -175 1716 -167
rect 1740 -151 1778 -142
rect 1740 -171 1749 -151
rect 1769 -171 1778 -151
rect 1631 -176 1667 -175
rect 1740 -179 1778 -171
rect 1844 -147 1929 -141
rect 1949 -142 1986 -141
rect 1844 -167 1852 -147
rect 1872 -148 1929 -147
rect 1872 -167 1901 -148
rect 1844 -168 1901 -167
rect 1922 -168 1929 -148
rect 1844 -175 1929 -168
rect 1948 -151 1986 -142
rect 1948 -171 1957 -151
rect 1977 -171 1986 -151
rect 1844 -176 1880 -175
rect 1948 -179 1986 -171
rect 2052 -147 2196 -141
rect 2052 -167 2060 -147
rect 2080 -167 2168 -147
rect 2188 -167 2196 -147
rect 2052 -175 2196 -167
rect 2052 -176 2088 -175
rect 2160 -176 2196 -175
rect 2262 -142 2299 -141
rect 2262 -143 2300 -142
rect 2262 -151 2326 -143
rect 2262 -171 2271 -151
rect 2291 -165 2326 -151
rect 2346 -165 2349 -145
rect 2291 -170 2349 -165
rect 2291 -171 2326 -170
rect 118 -269 157 -260
rect 118 -287 128 -269
rect 146 -287 157 -269
rect 118 -293 157 -287
rect 313 -217 563 -193
rect 313 -288 350 -217
rect 465 -278 496 -277
rect 118 -297 155 -293
rect 313 -308 322 -288
rect 342 -308 350 -288
rect 313 -318 350 -308
rect 409 -288 496 -278
rect 409 -308 418 -288
rect 438 -308 496 -288
rect 409 -317 496 -308
rect 409 -318 446 -317
rect 121 -368 158 -359
rect 119 -386 130 -368
rect 148 -386 158 -368
rect 465 -370 496 -317
rect 526 -288 563 -217
rect 734 -212 1127 -192
rect 1147 -212 1150 -192
rect 1528 -208 1565 -179
rect 734 -217 1150 -212
rect 1529 -210 1565 -208
rect 1741 -210 1778 -179
rect 734 -218 1075 -217
rect 678 -278 709 -277
rect 526 -308 535 -288
rect 555 -308 563 -288
rect 526 -318 563 -308
rect 622 -285 709 -278
rect 622 -288 683 -285
rect 622 -308 631 -288
rect 651 -305 683 -288
rect 704 -305 709 -285
rect 651 -308 709 -305
rect 622 -315 709 -308
rect 734 -288 771 -218
rect 1037 -219 1074 -218
rect 1529 -232 1778 -210
rect 1949 -211 1986 -179
rect 2262 -183 2326 -171
rect 2366 -209 2393 -31
rect 2225 -211 2393 -209
rect 1949 -237 2393 -211
rect 2225 -238 2393 -237
rect 886 -278 922 -277
rect 734 -308 743 -288
rect 763 -308 771 -288
rect 622 -317 678 -315
rect 622 -318 659 -317
rect 734 -318 771 -308
rect 830 -288 978 -278
rect 1078 -281 1174 -279
rect 830 -308 839 -288
rect 859 -308 949 -288
rect 969 -308 978 -288
rect 830 -317 978 -308
rect 1036 -288 1174 -281
rect 1036 -308 1045 -288
rect 1065 -308 1174 -288
rect 1036 -317 1174 -308
rect 830 -318 867 -317
rect 886 -369 922 -317
rect 941 -318 978 -317
rect 1037 -318 1074 -317
rect 357 -371 398 -370
rect 119 -535 158 -386
rect 249 -378 398 -371
rect 249 -398 367 -378
rect 387 -398 398 -378
rect 249 -406 398 -398
rect 465 -374 824 -370
rect 465 -379 787 -374
rect 465 -403 578 -379
rect 602 -398 787 -379
rect 811 -398 824 -374
rect 602 -403 824 -398
rect 465 -406 824 -403
rect 886 -406 921 -369
rect 989 -372 1089 -369
rect 989 -376 1056 -372
rect 989 -402 1001 -376
rect 1027 -398 1056 -376
rect 1082 -398 1089 -372
rect 1027 -402 1089 -398
rect 989 -406 1089 -402
rect 465 -427 496 -406
rect 886 -427 922 -406
rect 308 -428 345 -427
rect 307 -437 345 -428
rect 307 -457 316 -437
rect 336 -457 345 -437
rect 307 -465 345 -457
rect 411 -433 496 -427
rect 521 -428 558 -427
rect 411 -453 419 -433
rect 439 -453 496 -433
rect 411 -461 496 -453
rect 520 -437 558 -428
rect 520 -457 529 -437
rect 549 -457 558 -437
rect 411 -462 447 -461
rect 520 -465 558 -457
rect 624 -433 709 -427
rect 729 -428 766 -427
rect 624 -453 632 -433
rect 652 -434 709 -433
rect 652 -453 681 -434
rect 624 -454 681 -453
rect 702 -454 709 -434
rect 624 -461 709 -454
rect 728 -437 766 -428
rect 728 -457 737 -437
rect 757 -457 766 -437
rect 624 -462 660 -461
rect 728 -465 766 -457
rect 832 -432 976 -427
rect 832 -433 897 -432
rect 832 -453 840 -433
rect 860 -453 897 -433
rect 919 -433 976 -432
rect 919 -453 948 -433
rect 968 -453 976 -433
rect 832 -461 976 -453
rect 832 -462 868 -461
rect 940 -462 976 -461
rect 1042 -428 1079 -427
rect 1042 -429 1080 -428
rect 1042 -437 1106 -429
rect 1042 -457 1051 -437
rect 1071 -451 1106 -437
rect 1126 -451 1129 -431
rect 1071 -456 1129 -451
rect 1071 -457 1106 -456
rect 308 -494 345 -465
rect 309 -496 345 -494
rect 521 -496 558 -465
rect 309 -518 558 -496
rect 729 -497 766 -465
rect 1042 -469 1106 -457
rect 1146 -495 1173 -317
rect 1005 -497 1173 -495
rect 729 -523 1173 -497
rect 1325 -398 1575 -374
rect 1325 -469 1362 -398
rect 1477 -459 1508 -458
rect 1325 -489 1334 -469
rect 1354 -489 1362 -469
rect 1325 -499 1362 -489
rect 1421 -469 1508 -459
rect 1421 -489 1430 -469
rect 1450 -489 1508 -469
rect 1421 -498 1508 -489
rect 1421 -499 1458 -498
rect 729 -533 751 -523
rect 1005 -524 1173 -523
rect 689 -535 751 -533
rect 119 -542 751 -535
rect 118 -551 751 -542
rect 1477 -551 1508 -498
rect 1538 -469 1575 -398
rect 1746 -393 2139 -373
rect 2159 -393 2162 -373
rect 1746 -398 2162 -393
rect 1746 -399 2087 -398
rect 1690 -459 1721 -458
rect 1538 -489 1547 -469
rect 1567 -489 1575 -469
rect 1538 -499 1575 -489
rect 1634 -466 1721 -459
rect 1634 -469 1695 -466
rect 1634 -489 1643 -469
rect 1663 -486 1695 -469
rect 1716 -486 1721 -466
rect 1663 -489 1721 -486
rect 1634 -496 1721 -489
rect 1746 -469 1783 -399
rect 2049 -400 2086 -399
rect 1898 -459 1934 -458
rect 1746 -489 1755 -469
rect 1775 -489 1783 -469
rect 1634 -498 1690 -496
rect 1634 -499 1671 -498
rect 1746 -499 1783 -489
rect 1842 -469 1990 -459
rect 2090 -462 2186 -460
rect 1842 -489 1851 -469
rect 1871 -489 1961 -469
rect 1981 -489 1990 -469
rect 1842 -498 1990 -489
rect 2048 -469 2186 -462
rect 2048 -489 2057 -469
rect 2077 -489 2186 -469
rect 2048 -498 2186 -489
rect 1842 -499 1879 -498
rect 1898 -550 1934 -498
rect 1953 -499 1990 -498
rect 2049 -499 2086 -498
rect 118 -569 128 -551
rect 146 -552 751 -551
rect 1369 -552 1410 -551
rect 146 -557 167 -552
rect 146 -569 158 -557
rect 1261 -559 1410 -552
rect 118 -577 158 -569
rect 201 -570 227 -569
rect 118 -579 155 -577
rect 201 -588 755 -570
rect 1261 -579 1379 -559
rect 1399 -579 1410 -559
rect 1261 -587 1410 -579
rect 1477 -555 1836 -551
rect 1477 -560 1799 -555
rect 1477 -584 1590 -560
rect 1614 -579 1799 -560
rect 1823 -579 1836 -555
rect 1614 -584 1836 -579
rect 1477 -587 1836 -584
rect 1898 -587 1933 -550
rect 2001 -553 2101 -550
rect 2001 -557 2068 -553
rect 2001 -583 2013 -557
rect 2039 -579 2068 -557
rect 2094 -579 2101 -553
rect 2039 -583 2101 -579
rect 2001 -587 2101 -583
rect 121 -647 158 -641
rect 201 -647 227 -588
rect 734 -607 755 -588
rect 121 -650 227 -647
rect 121 -668 130 -650
rect 148 -664 227 -650
rect 312 -632 562 -608
rect 148 -666 224 -664
rect 148 -668 158 -666
rect 121 -678 158 -668
rect 126 -743 157 -678
rect 312 -703 349 -632
rect 464 -693 495 -692
rect 312 -723 321 -703
rect 341 -723 349 -703
rect 312 -733 349 -723
rect 408 -703 495 -693
rect 408 -723 417 -703
rect 437 -723 495 -703
rect 408 -732 495 -723
rect 408 -733 445 -732
rect 125 -752 162 -743
rect 125 -770 135 -752
rect 153 -770 162 -752
rect 125 -780 162 -770
rect 464 -785 495 -732
rect 525 -703 562 -632
rect 733 -627 1126 -607
rect 1146 -627 1149 -607
rect 1477 -608 1508 -587
rect 1898 -608 1934 -587
rect 1320 -609 1357 -608
rect 733 -632 1149 -627
rect 1319 -618 1357 -609
rect 733 -633 1074 -632
rect 677 -693 708 -692
rect 525 -723 534 -703
rect 554 -723 562 -703
rect 525 -733 562 -723
rect 621 -700 708 -693
rect 621 -703 682 -700
rect 621 -723 630 -703
rect 650 -720 682 -703
rect 703 -720 708 -700
rect 650 -723 708 -720
rect 621 -730 708 -723
rect 733 -703 770 -633
rect 1036 -634 1073 -633
rect 1319 -638 1328 -618
rect 1348 -638 1357 -618
rect 1319 -646 1357 -638
rect 1423 -614 1508 -608
rect 1533 -609 1570 -608
rect 1423 -634 1431 -614
rect 1451 -634 1508 -614
rect 1423 -642 1508 -634
rect 1532 -618 1570 -609
rect 1532 -638 1541 -618
rect 1561 -638 1570 -618
rect 1423 -643 1459 -642
rect 1532 -646 1570 -638
rect 1636 -614 1721 -608
rect 1741 -609 1778 -608
rect 1636 -634 1644 -614
rect 1664 -615 1721 -614
rect 1664 -634 1693 -615
rect 1636 -635 1693 -634
rect 1714 -635 1721 -615
rect 1636 -642 1721 -635
rect 1740 -618 1778 -609
rect 1740 -638 1749 -618
rect 1769 -638 1778 -618
rect 1636 -643 1672 -642
rect 1740 -646 1778 -638
rect 1844 -614 1988 -608
rect 1844 -634 1852 -614
rect 1872 -634 1904 -614
rect 1928 -634 1960 -614
rect 1980 -634 1988 -614
rect 1844 -642 1988 -634
rect 1844 -643 1880 -642
rect 1952 -643 1988 -642
rect 2054 -609 2091 -608
rect 2054 -610 2092 -609
rect 2054 -618 2118 -610
rect 2054 -638 2063 -618
rect 2083 -632 2118 -618
rect 2138 -632 2141 -612
rect 2083 -637 2141 -632
rect 2083 -638 2118 -637
rect 1320 -675 1357 -646
rect 1321 -677 1357 -675
rect 1533 -677 1570 -646
rect 885 -693 921 -692
rect 733 -723 742 -703
rect 762 -723 770 -703
rect 621 -732 677 -730
rect 621 -733 658 -732
rect 733 -733 770 -723
rect 829 -703 977 -693
rect 1077 -696 1173 -694
rect 829 -723 838 -703
rect 858 -723 948 -703
rect 968 -723 977 -703
rect 829 -732 977 -723
rect 1035 -703 1173 -696
rect 1321 -699 1570 -677
rect 1741 -678 1778 -646
rect 2054 -650 2118 -638
rect 2158 -676 2185 -498
rect 2017 -678 2185 -676
rect 1741 -682 2185 -678
rect 1035 -723 1044 -703
rect 1064 -723 1173 -703
rect 1741 -701 1790 -682
rect 1810 -701 2185 -682
rect 1741 -704 2185 -701
rect 2017 -705 2185 -704
rect 1035 -732 1173 -723
rect 829 -733 866 -732
rect 885 -784 921 -732
rect 940 -733 977 -732
rect 1036 -733 1073 -732
rect 356 -786 397 -785
rect 248 -793 397 -786
rect 248 -813 366 -793
rect 386 -813 397 -793
rect 248 -821 397 -813
rect 464 -789 823 -785
rect 464 -794 786 -789
rect 464 -818 577 -794
rect 601 -813 786 -794
rect 810 -813 823 -789
rect 601 -818 823 -813
rect 464 -821 823 -818
rect 885 -821 920 -784
rect 988 -787 1088 -784
rect 988 -791 1055 -787
rect 988 -817 1000 -791
rect 1026 -813 1055 -791
rect 1081 -813 1088 -787
rect 1026 -817 1088 -813
rect 988 -821 1088 -817
rect 464 -842 495 -821
rect 885 -842 921 -821
rect 128 -851 165 -842
rect 307 -843 344 -842
rect 128 -869 137 -851
rect 155 -869 165 -851
rect 128 -879 165 -869
rect 129 -914 165 -879
rect 306 -852 344 -843
rect 306 -872 315 -852
rect 335 -872 344 -852
rect 306 -880 344 -872
rect 410 -848 495 -842
rect 520 -843 557 -842
rect 410 -868 418 -848
rect 438 -868 495 -848
rect 410 -876 495 -868
rect 519 -852 557 -843
rect 519 -872 528 -852
rect 548 -872 557 -852
rect 410 -877 446 -876
rect 519 -880 557 -872
rect 623 -848 708 -842
rect 728 -843 765 -842
rect 623 -868 631 -848
rect 651 -849 708 -848
rect 651 -868 680 -849
rect 623 -869 680 -868
rect 701 -869 708 -849
rect 623 -876 708 -869
rect 727 -852 765 -843
rect 727 -872 736 -852
rect 756 -872 765 -852
rect 623 -877 659 -876
rect 727 -880 765 -872
rect 831 -848 975 -842
rect 831 -868 839 -848
rect 859 -849 947 -848
rect 859 -868 887 -849
rect 831 -870 887 -868
rect 909 -868 947 -849
rect 967 -868 975 -848
rect 909 -870 975 -868
rect 831 -876 975 -870
rect 831 -877 867 -876
rect 939 -877 975 -876
rect 1041 -843 1078 -842
rect 1041 -844 1079 -843
rect 1041 -852 1105 -844
rect 1041 -872 1050 -852
rect 1070 -866 1105 -852
rect 1125 -866 1128 -846
rect 1070 -871 1128 -866
rect 1070 -872 1105 -871
rect 307 -909 344 -880
rect 127 -955 165 -914
rect 308 -911 344 -909
rect 520 -911 557 -880
rect 308 -933 557 -911
rect 728 -912 765 -880
rect 1041 -884 1105 -872
rect 1145 -910 1172 -732
rect 1004 -912 1172 -910
rect 728 -938 1172 -912
rect 729 -955 753 -938
rect 1004 -939 1172 -938
rect 127 -973 754 -955
rect 1380 -959 1630 -935
rect 127 -979 165 -973
rect 127 -1003 164 -979
rect 127 -1027 162 -1003
rect 125 -1036 162 -1027
rect 125 -1054 135 -1036
rect 153 -1054 162 -1036
rect 125 -1064 162 -1054
rect 1380 -1030 1417 -959
rect 1532 -1020 1563 -1019
rect 1380 -1050 1389 -1030
rect 1409 -1050 1417 -1030
rect 1380 -1060 1417 -1050
rect 1476 -1030 1563 -1020
rect 1476 -1050 1485 -1030
rect 1505 -1050 1563 -1030
rect 1476 -1059 1563 -1050
rect 1476 -1060 1513 -1059
rect 1532 -1112 1563 -1059
rect 1593 -1030 1630 -959
rect 1801 -954 2194 -934
rect 2214 -954 2217 -934
rect 1801 -959 2217 -954
rect 1801 -960 2142 -959
rect 1745 -1020 1776 -1019
rect 1593 -1050 1602 -1030
rect 1622 -1050 1630 -1030
rect 1593 -1060 1630 -1050
rect 1689 -1027 1776 -1020
rect 1689 -1030 1750 -1027
rect 1689 -1050 1698 -1030
rect 1718 -1047 1750 -1030
rect 1771 -1047 1776 -1027
rect 1718 -1050 1776 -1047
rect 1689 -1057 1776 -1050
rect 1801 -1030 1838 -960
rect 2104 -961 2141 -960
rect 1953 -1020 1989 -1019
rect 1801 -1050 1810 -1030
rect 1830 -1050 1838 -1030
rect 1689 -1059 1745 -1057
rect 1689 -1060 1726 -1059
rect 1801 -1060 1838 -1050
rect 1897 -1030 2045 -1020
rect 2145 -1023 2241 -1021
rect 1897 -1050 1906 -1030
rect 1926 -1050 2016 -1030
rect 2036 -1050 2045 -1030
rect 1897 -1059 2045 -1050
rect 2103 -1030 2241 -1023
rect 2103 -1050 2112 -1030
rect 2132 -1050 2241 -1030
rect 2103 -1059 2241 -1050
rect 1897 -1060 1934 -1059
rect 1953 -1111 1989 -1059
rect 2008 -1060 2045 -1059
rect 2104 -1060 2141 -1059
rect 1424 -1113 1465 -1112
rect 1316 -1120 1465 -1113
rect 128 -1128 165 -1126
rect 128 -1129 776 -1128
rect 127 -1135 776 -1129
rect 127 -1153 137 -1135
rect 155 -1149 776 -1135
rect 1316 -1140 1434 -1120
rect 1454 -1140 1465 -1120
rect 1316 -1148 1465 -1140
rect 1532 -1116 1891 -1112
rect 1532 -1121 1854 -1116
rect 1532 -1145 1645 -1121
rect 1669 -1140 1854 -1121
rect 1878 -1140 1891 -1116
rect 1669 -1145 1891 -1140
rect 1532 -1148 1891 -1145
rect 1953 -1148 1988 -1111
rect 2056 -1114 2156 -1111
rect 2056 -1118 2123 -1114
rect 2056 -1144 2068 -1118
rect 2094 -1140 2123 -1118
rect 2149 -1140 2156 -1114
rect 2094 -1144 2156 -1140
rect 2056 -1148 2156 -1144
rect 155 -1153 165 -1149
rect 606 -1150 776 -1149
rect 127 -1163 165 -1153
rect 127 -1241 162 -1163
rect 739 -1173 776 -1150
rect 1532 -1169 1563 -1148
rect 1953 -1169 1989 -1148
rect 1375 -1170 1412 -1169
rect 123 -1250 162 -1241
rect 123 -1268 133 -1250
rect 151 -1268 162 -1250
rect 123 -1274 162 -1268
rect 318 -1198 568 -1174
rect 318 -1269 355 -1198
rect 470 -1259 501 -1258
rect 123 -1278 160 -1274
rect 318 -1289 327 -1269
rect 347 -1289 355 -1269
rect 318 -1299 355 -1289
rect 414 -1269 501 -1259
rect 414 -1289 423 -1269
rect 443 -1289 501 -1269
rect 414 -1298 501 -1289
rect 414 -1299 451 -1298
rect 126 -1349 163 -1340
rect 124 -1367 135 -1349
rect 153 -1367 163 -1349
rect 470 -1351 501 -1298
rect 531 -1269 568 -1198
rect 739 -1193 1132 -1173
rect 1152 -1193 1155 -1173
rect 739 -1198 1155 -1193
rect 1374 -1179 1412 -1170
rect 739 -1199 1080 -1198
rect 1374 -1199 1383 -1179
rect 1403 -1199 1412 -1179
rect 683 -1259 714 -1258
rect 531 -1289 540 -1269
rect 560 -1289 568 -1269
rect 531 -1299 568 -1289
rect 627 -1266 714 -1259
rect 627 -1269 688 -1266
rect 627 -1289 636 -1269
rect 656 -1286 688 -1269
rect 709 -1286 714 -1266
rect 656 -1289 714 -1286
rect 627 -1296 714 -1289
rect 739 -1269 776 -1199
rect 1042 -1200 1079 -1199
rect 1374 -1207 1412 -1199
rect 1478 -1175 1563 -1169
rect 1588 -1170 1625 -1169
rect 1478 -1195 1486 -1175
rect 1506 -1195 1563 -1175
rect 1478 -1203 1563 -1195
rect 1587 -1179 1625 -1170
rect 1587 -1199 1596 -1179
rect 1616 -1199 1625 -1179
rect 1478 -1204 1514 -1203
rect 1587 -1207 1625 -1199
rect 1691 -1175 1776 -1169
rect 1796 -1170 1833 -1169
rect 1691 -1195 1699 -1175
rect 1719 -1176 1776 -1175
rect 1719 -1195 1748 -1176
rect 1691 -1196 1748 -1195
rect 1769 -1196 1776 -1176
rect 1691 -1203 1776 -1196
rect 1795 -1179 1833 -1170
rect 1795 -1199 1804 -1179
rect 1824 -1199 1833 -1179
rect 1691 -1204 1727 -1203
rect 1795 -1207 1833 -1199
rect 1899 -1175 2043 -1169
rect 1899 -1195 1907 -1175
rect 1927 -1176 2015 -1175
rect 1927 -1195 1960 -1176
rect 1983 -1195 2015 -1176
rect 2035 -1195 2043 -1175
rect 1899 -1203 2043 -1195
rect 1899 -1204 1935 -1203
rect 2007 -1204 2043 -1203
rect 2109 -1170 2146 -1169
rect 2109 -1171 2147 -1170
rect 2109 -1179 2173 -1171
rect 2109 -1199 2118 -1179
rect 2138 -1193 2173 -1179
rect 2193 -1193 2196 -1173
rect 2138 -1198 2196 -1193
rect 2138 -1199 2173 -1198
rect 1375 -1236 1412 -1207
rect 1376 -1238 1412 -1236
rect 1588 -1238 1625 -1207
rect 891 -1259 927 -1258
rect 739 -1289 748 -1269
rect 768 -1289 776 -1269
rect 627 -1298 683 -1296
rect 627 -1299 664 -1298
rect 739 -1299 776 -1289
rect 835 -1269 983 -1259
rect 1376 -1260 1625 -1238
rect 1796 -1239 1833 -1207
rect 2109 -1211 2173 -1199
rect 2213 -1237 2240 -1059
rect 2072 -1239 2240 -1237
rect 1796 -1250 2240 -1239
rect 2303 -1239 2333 -238
rect 2303 -1244 2335 -1239
rect 1083 -1262 1179 -1260
rect 835 -1289 844 -1269
rect 864 -1289 954 -1269
rect 974 -1289 983 -1269
rect 835 -1298 983 -1289
rect 1041 -1269 1179 -1262
rect 1796 -1265 2242 -1250
rect 2072 -1266 2242 -1265
rect 1041 -1289 1050 -1269
rect 1070 -1289 1179 -1269
rect 1041 -1298 1179 -1289
rect 835 -1299 872 -1298
rect 891 -1350 927 -1298
rect 946 -1299 983 -1298
rect 1042 -1299 1079 -1298
rect 362 -1352 403 -1351
rect 124 -1516 163 -1367
rect 254 -1359 403 -1352
rect 254 -1379 372 -1359
rect 392 -1379 403 -1359
rect 254 -1387 403 -1379
rect 470 -1355 829 -1351
rect 470 -1360 792 -1355
rect 470 -1384 583 -1360
rect 607 -1379 792 -1360
rect 816 -1379 829 -1355
rect 607 -1384 829 -1379
rect 470 -1387 829 -1384
rect 891 -1387 926 -1350
rect 994 -1353 1094 -1350
rect 994 -1357 1061 -1353
rect 994 -1383 1006 -1357
rect 1032 -1379 1061 -1357
rect 1087 -1379 1094 -1353
rect 1032 -1383 1094 -1379
rect 994 -1387 1094 -1383
rect 470 -1408 501 -1387
rect 891 -1408 927 -1387
rect 313 -1409 350 -1408
rect 312 -1418 350 -1409
rect 312 -1438 321 -1418
rect 341 -1438 350 -1418
rect 312 -1446 350 -1438
rect 416 -1414 501 -1408
rect 526 -1409 563 -1408
rect 416 -1434 424 -1414
rect 444 -1434 501 -1414
rect 416 -1442 501 -1434
rect 525 -1418 563 -1409
rect 525 -1438 534 -1418
rect 554 -1438 563 -1418
rect 416 -1443 452 -1442
rect 525 -1446 563 -1438
rect 629 -1414 714 -1408
rect 734 -1409 771 -1408
rect 629 -1434 637 -1414
rect 657 -1415 714 -1414
rect 657 -1434 686 -1415
rect 629 -1435 686 -1434
rect 707 -1435 714 -1415
rect 629 -1442 714 -1435
rect 733 -1418 771 -1409
rect 733 -1438 742 -1418
rect 762 -1438 771 -1418
rect 629 -1443 665 -1442
rect 733 -1446 771 -1438
rect 837 -1413 981 -1408
rect 837 -1414 902 -1413
rect 837 -1434 845 -1414
rect 865 -1434 902 -1414
rect 924 -1414 981 -1413
rect 924 -1434 953 -1414
rect 973 -1434 981 -1414
rect 837 -1442 981 -1434
rect 837 -1443 873 -1442
rect 945 -1443 981 -1442
rect 1047 -1409 1084 -1408
rect 1047 -1410 1085 -1409
rect 1047 -1418 1111 -1410
rect 1047 -1438 1056 -1418
rect 1076 -1432 1111 -1418
rect 1131 -1432 1134 -1412
rect 1076 -1437 1134 -1432
rect 1076 -1438 1111 -1437
rect 313 -1475 350 -1446
rect 314 -1477 350 -1475
rect 526 -1477 563 -1446
rect 314 -1499 563 -1477
rect 734 -1478 771 -1446
rect 1047 -1450 1111 -1438
rect 1151 -1476 1178 -1298
rect 1010 -1478 1178 -1476
rect 734 -1504 1178 -1478
rect 1330 -1379 1580 -1355
rect 1330 -1450 1367 -1379
rect 1482 -1440 1513 -1439
rect 1330 -1470 1339 -1450
rect 1359 -1470 1367 -1450
rect 1330 -1480 1367 -1470
rect 1426 -1450 1513 -1440
rect 1426 -1470 1435 -1450
rect 1455 -1470 1513 -1450
rect 1426 -1479 1513 -1470
rect 1426 -1480 1463 -1479
rect 734 -1514 756 -1504
rect 1010 -1505 1178 -1504
rect 694 -1516 756 -1514
rect 124 -1523 756 -1516
rect 123 -1532 756 -1523
rect 1482 -1532 1513 -1479
rect 1543 -1450 1580 -1379
rect 1751 -1374 2144 -1354
rect 2164 -1374 2167 -1354
rect 1751 -1379 2167 -1374
rect 1751 -1380 2092 -1379
rect 1695 -1440 1726 -1439
rect 1543 -1470 1552 -1450
rect 1572 -1470 1580 -1450
rect 1543 -1480 1580 -1470
rect 1639 -1447 1726 -1440
rect 1639 -1450 1700 -1447
rect 1639 -1470 1648 -1450
rect 1668 -1467 1700 -1450
rect 1721 -1467 1726 -1447
rect 1668 -1470 1726 -1467
rect 1639 -1477 1726 -1470
rect 1751 -1450 1788 -1380
rect 2054 -1381 2091 -1380
rect 1903 -1440 1939 -1439
rect 1751 -1470 1760 -1450
rect 1780 -1470 1788 -1450
rect 1639 -1479 1695 -1477
rect 1639 -1480 1676 -1479
rect 1751 -1480 1788 -1470
rect 1847 -1450 1995 -1440
rect 2095 -1443 2191 -1441
rect 1847 -1470 1856 -1450
rect 1876 -1470 1966 -1450
rect 1986 -1470 1995 -1450
rect 1847 -1479 1995 -1470
rect 2053 -1450 2191 -1443
rect 2053 -1470 2062 -1450
rect 2082 -1470 2191 -1450
rect 2053 -1479 2191 -1470
rect 1847 -1480 1884 -1479
rect 1903 -1531 1939 -1479
rect 1958 -1480 1995 -1479
rect 2054 -1480 2091 -1479
rect 123 -1550 133 -1532
rect 151 -1533 756 -1532
rect 1374 -1533 1415 -1532
rect 151 -1538 172 -1533
rect 151 -1550 163 -1538
rect 1266 -1540 1415 -1533
rect 123 -1558 163 -1550
rect 206 -1551 232 -1550
rect 123 -1560 160 -1558
rect 206 -1569 760 -1551
rect 1266 -1560 1384 -1540
rect 1404 -1560 1415 -1540
rect 1266 -1568 1415 -1560
rect 1482 -1536 1841 -1532
rect 1482 -1541 1804 -1536
rect 1482 -1565 1595 -1541
rect 1619 -1560 1804 -1541
rect 1828 -1560 1841 -1536
rect 1619 -1565 1841 -1560
rect 1482 -1568 1841 -1565
rect 1903 -1568 1938 -1531
rect 2006 -1534 2106 -1531
rect 2006 -1538 2073 -1534
rect 2006 -1564 2018 -1538
rect 2044 -1560 2073 -1538
rect 2099 -1560 2106 -1534
rect 2044 -1564 2106 -1560
rect 2006 -1568 2106 -1564
rect 126 -1628 163 -1622
rect 206 -1628 232 -1569
rect 739 -1588 760 -1569
rect 126 -1631 232 -1628
rect 126 -1649 135 -1631
rect 153 -1645 232 -1631
rect 317 -1613 567 -1589
rect 153 -1647 229 -1645
rect 153 -1649 163 -1647
rect 126 -1659 163 -1649
rect 131 -1724 162 -1659
rect 317 -1684 354 -1613
rect 469 -1674 500 -1673
rect 317 -1704 326 -1684
rect 346 -1704 354 -1684
rect 317 -1714 354 -1704
rect 413 -1684 500 -1674
rect 413 -1704 422 -1684
rect 442 -1704 500 -1684
rect 413 -1713 500 -1704
rect 413 -1714 450 -1713
rect 130 -1733 167 -1724
rect 130 -1751 140 -1733
rect 158 -1751 167 -1733
rect 130 -1761 167 -1751
rect 469 -1766 500 -1713
rect 530 -1684 567 -1613
rect 738 -1608 1131 -1588
rect 1151 -1608 1154 -1588
rect 1482 -1589 1513 -1568
rect 1903 -1589 1939 -1568
rect 1325 -1590 1362 -1589
rect 738 -1613 1154 -1608
rect 1324 -1599 1362 -1590
rect 738 -1614 1079 -1613
rect 682 -1674 713 -1673
rect 530 -1704 539 -1684
rect 559 -1704 567 -1684
rect 530 -1714 567 -1704
rect 626 -1681 713 -1674
rect 626 -1684 687 -1681
rect 626 -1704 635 -1684
rect 655 -1701 687 -1684
rect 708 -1701 713 -1681
rect 655 -1704 713 -1701
rect 626 -1711 713 -1704
rect 738 -1684 775 -1614
rect 1041 -1615 1078 -1614
rect 1324 -1619 1333 -1599
rect 1353 -1619 1362 -1599
rect 1324 -1627 1362 -1619
rect 1428 -1595 1513 -1589
rect 1538 -1590 1575 -1589
rect 1428 -1615 1436 -1595
rect 1456 -1615 1513 -1595
rect 1428 -1623 1513 -1615
rect 1537 -1599 1575 -1590
rect 1537 -1619 1546 -1599
rect 1566 -1619 1575 -1599
rect 1428 -1624 1464 -1623
rect 1537 -1627 1575 -1619
rect 1641 -1595 1726 -1589
rect 1746 -1590 1783 -1589
rect 1641 -1615 1649 -1595
rect 1669 -1596 1726 -1595
rect 1669 -1615 1698 -1596
rect 1641 -1616 1698 -1615
rect 1719 -1616 1726 -1596
rect 1641 -1623 1726 -1616
rect 1745 -1599 1783 -1590
rect 1745 -1619 1754 -1599
rect 1774 -1619 1783 -1599
rect 1641 -1624 1677 -1623
rect 1745 -1627 1783 -1619
rect 1849 -1594 1993 -1589
rect 1849 -1595 1908 -1594
rect 1849 -1615 1857 -1595
rect 1877 -1614 1908 -1595
rect 1932 -1595 1993 -1594
rect 1932 -1614 1965 -1595
rect 1877 -1615 1965 -1614
rect 1985 -1615 1993 -1595
rect 1849 -1623 1993 -1615
rect 1849 -1624 1885 -1623
rect 1957 -1624 1993 -1623
rect 2059 -1590 2096 -1589
rect 2059 -1591 2097 -1590
rect 2059 -1599 2123 -1591
rect 2059 -1619 2068 -1599
rect 2088 -1613 2123 -1599
rect 2143 -1613 2146 -1593
rect 2088 -1618 2146 -1613
rect 2088 -1619 2123 -1618
rect 1325 -1656 1362 -1627
rect 1326 -1658 1362 -1656
rect 1538 -1658 1575 -1627
rect 890 -1674 926 -1673
rect 738 -1704 747 -1684
rect 767 -1704 775 -1684
rect 626 -1713 682 -1711
rect 626 -1714 663 -1713
rect 738 -1714 775 -1704
rect 834 -1684 982 -1674
rect 1082 -1677 1178 -1675
rect 834 -1704 843 -1684
rect 863 -1704 953 -1684
rect 973 -1704 982 -1684
rect 834 -1713 982 -1704
rect 1040 -1684 1178 -1677
rect 1326 -1680 1575 -1658
rect 1746 -1659 1783 -1627
rect 2059 -1631 2123 -1619
rect 2163 -1657 2190 -1479
rect 2022 -1659 2190 -1657
rect 1746 -1663 2190 -1659
rect 1040 -1704 1049 -1684
rect 1069 -1704 1178 -1684
rect 1746 -1682 1795 -1663
rect 1815 -1682 2190 -1663
rect 1746 -1685 2190 -1682
rect 2022 -1686 2190 -1685
rect 2211 -1660 2242 -1266
rect 2303 -1262 2308 -1244
rect 2328 -1262 2335 -1244
rect 2303 -1267 2335 -1262
rect 2306 -1269 2335 -1267
rect 2211 -1686 2216 -1660
rect 2235 -1686 2242 -1660
rect 2211 -1689 2242 -1686
rect 1040 -1713 1178 -1704
rect 834 -1714 871 -1713
rect 890 -1765 926 -1713
rect 945 -1714 982 -1713
rect 1041 -1714 1078 -1713
rect 361 -1767 402 -1766
rect 253 -1774 402 -1767
rect 253 -1794 371 -1774
rect 391 -1794 402 -1774
rect 253 -1802 402 -1794
rect 469 -1770 828 -1766
rect 469 -1775 791 -1770
rect 469 -1799 582 -1775
rect 606 -1794 791 -1775
rect 815 -1794 828 -1770
rect 606 -1799 828 -1794
rect 469 -1802 828 -1799
rect 890 -1802 925 -1765
rect 993 -1768 1093 -1765
rect 993 -1772 1060 -1768
rect 993 -1798 1005 -1772
rect 1031 -1794 1060 -1772
rect 1086 -1794 1093 -1768
rect 1031 -1798 1093 -1794
rect 993 -1802 1093 -1798
rect 469 -1823 500 -1802
rect 890 -1823 926 -1802
rect 133 -1832 170 -1823
rect 312 -1824 349 -1823
rect 133 -1850 142 -1832
rect 160 -1850 170 -1832
rect 133 -1860 170 -1850
rect 134 -1895 170 -1860
rect 311 -1833 349 -1824
rect 311 -1853 320 -1833
rect 340 -1853 349 -1833
rect 311 -1861 349 -1853
rect 415 -1829 500 -1823
rect 525 -1824 562 -1823
rect 415 -1849 423 -1829
rect 443 -1849 500 -1829
rect 415 -1857 500 -1849
rect 524 -1833 562 -1824
rect 524 -1853 533 -1833
rect 553 -1853 562 -1833
rect 415 -1858 451 -1857
rect 524 -1861 562 -1853
rect 628 -1829 713 -1823
rect 733 -1824 770 -1823
rect 628 -1849 636 -1829
rect 656 -1830 713 -1829
rect 656 -1849 685 -1830
rect 628 -1850 685 -1849
rect 706 -1850 713 -1830
rect 628 -1857 713 -1850
rect 732 -1833 770 -1824
rect 732 -1853 741 -1833
rect 761 -1853 770 -1833
rect 628 -1858 664 -1857
rect 732 -1861 770 -1853
rect 836 -1829 980 -1823
rect 836 -1849 844 -1829
rect 864 -1830 952 -1829
rect 864 -1849 892 -1830
rect 836 -1851 892 -1849
rect 914 -1849 952 -1830
rect 972 -1849 980 -1829
rect 914 -1851 980 -1849
rect 836 -1857 980 -1851
rect 836 -1858 872 -1857
rect 944 -1858 980 -1857
rect 1046 -1824 1083 -1823
rect 1046 -1825 1084 -1824
rect 1046 -1833 1110 -1825
rect 1046 -1853 1055 -1833
rect 1075 -1847 1110 -1833
rect 1130 -1847 1133 -1827
rect 1075 -1852 1133 -1847
rect 1075 -1853 1110 -1852
rect 312 -1890 349 -1861
rect 132 -1936 170 -1895
rect 313 -1892 349 -1890
rect 525 -1892 562 -1861
rect 313 -1914 562 -1892
rect 733 -1893 770 -1861
rect 1046 -1865 1110 -1853
rect 1150 -1891 1177 -1713
rect 1009 -1893 1177 -1891
rect 733 -1919 1177 -1893
rect 734 -1936 758 -1919
rect 1009 -1920 1177 -1919
rect 132 -1954 759 -1936
rect 132 -1960 170 -1954
<< viali >>
rect 1115 1748 1135 1768
rect 671 1655 692 1675
rect 1044 1562 1070 1588
rect 669 1506 690 1526
rect 885 1507 907 1528
rect 1094 1509 1114 1529
rect 2127 1567 2147 1587
rect 1683 1474 1704 1494
rect 2056 1381 2082 1407
rect 1114 1333 1134 1353
rect 670 1240 691 1260
rect 1681 1325 1702 1345
rect 1892 1326 1916 1346
rect 2106 1328 2126 1348
rect 1778 1259 1798 1278
rect 1043 1147 1069 1173
rect 668 1091 689 1111
rect 875 1090 897 1111
rect 1093 1094 1113 1114
rect 2182 1006 2202 1026
rect 1738 913 1759 933
rect 2111 820 2137 846
rect 1120 767 1140 787
rect 676 674 697 694
rect 1736 764 1757 784
rect 1951 766 1975 783
rect 2161 767 2181 787
rect 1049 581 1075 607
rect 674 525 695 545
rect 890 526 912 547
rect 1099 528 1119 548
rect 2132 586 2152 606
rect 1688 493 1709 513
rect 2061 400 2087 426
rect 1119 352 1139 372
rect 675 259 696 279
rect 1686 344 1707 364
rect 1896 346 1920 366
rect 2111 347 2131 367
rect 1783 278 1803 297
rect 2204 274 2223 300
rect 1048 166 1074 192
rect 673 110 694 130
rect 880 109 902 130
rect 1098 113 1118 133
rect 2347 74 2367 94
rect 1903 -19 1924 1
rect 2276 -112 2302 -86
rect 1901 -168 1922 -148
rect 2326 -165 2346 -145
rect 1127 -212 1147 -192
rect 683 -305 704 -285
rect 1056 -398 1082 -372
rect 681 -454 702 -434
rect 897 -453 919 -432
rect 1106 -451 1126 -431
rect 2139 -393 2159 -373
rect 1695 -486 1716 -466
rect 2068 -579 2094 -553
rect 1126 -627 1146 -607
rect 682 -720 703 -700
rect 1693 -635 1714 -615
rect 1904 -634 1928 -614
rect 2118 -632 2138 -612
rect 1790 -701 1810 -682
rect 1055 -813 1081 -787
rect 680 -869 701 -849
rect 887 -870 909 -849
rect 1105 -866 1125 -846
rect 2194 -954 2214 -934
rect 1750 -1047 1771 -1027
rect 2123 -1140 2149 -1114
rect 1132 -1193 1152 -1173
rect 688 -1286 709 -1266
rect 1748 -1196 1769 -1176
rect 1960 -1195 1983 -1176
rect 2173 -1193 2193 -1173
rect 1061 -1379 1087 -1353
rect 686 -1435 707 -1415
rect 902 -1434 924 -1413
rect 1111 -1432 1131 -1412
rect 2144 -1374 2164 -1354
rect 1700 -1467 1721 -1447
rect 2073 -1560 2099 -1534
rect 1131 -1608 1151 -1588
rect 687 -1701 708 -1681
rect 1698 -1616 1719 -1596
rect 1908 -1614 1932 -1594
rect 2123 -1613 2143 -1593
rect 1795 -1682 1815 -1663
rect 2308 -1262 2328 -1244
rect 2216 -1686 2235 -1660
rect 1060 -1794 1086 -1768
rect 685 -1850 706 -1830
rect 892 -1851 914 -1830
rect 1110 -1847 1130 -1827
<< metal1 >>
rect 1111 1773 1143 1774
rect 1108 1768 1143 1773
rect 1108 1748 1115 1768
rect 1135 1748 1143 1768
rect 1108 1740 1143 1748
rect 664 1675 696 1682
rect 664 1655 671 1675
rect 692 1655 696 1675
rect 664 1590 696 1655
rect 1034 1590 1074 1591
rect 664 1588 1076 1590
rect 664 1562 1044 1588
rect 1070 1562 1076 1588
rect 664 1554 1076 1562
rect 664 1526 696 1554
rect 1109 1534 1143 1740
rect 664 1506 669 1526
rect 690 1506 696 1526
rect 664 1499 696 1506
rect 873 1528 913 1533
rect 873 1507 885 1528
rect 907 1507 913 1528
rect 873 1495 913 1507
rect 1087 1529 1143 1534
rect 1087 1509 1094 1529
rect 1114 1509 1143 1529
rect 1087 1502 1143 1509
rect 1200 1603 2157 1622
rect 1087 1501 1122 1502
rect 879 1463 907 1495
rect 1200 1463 1231 1603
rect 2120 1587 2155 1603
rect 2120 1567 2127 1587
rect 2147 1567 2155 1587
rect 2120 1559 2155 1567
rect 879 1432 1231 1463
rect 1676 1494 1708 1501
rect 1676 1474 1683 1494
rect 1704 1474 1708 1494
rect 1676 1409 1708 1474
rect 2046 1409 2086 1410
rect 1676 1407 2088 1409
rect 1676 1381 2056 1407
rect 2082 1381 2088 1407
rect 1676 1373 2088 1381
rect 1110 1358 1142 1359
rect 1107 1353 1142 1358
rect 1107 1333 1114 1353
rect 1134 1333 1142 1353
rect 1107 1325 1142 1333
rect 663 1260 695 1267
rect 663 1240 670 1260
rect 691 1240 695 1260
rect 663 1175 695 1240
rect 1033 1175 1073 1176
rect 663 1173 1075 1175
rect 663 1147 1043 1173
rect 1069 1147 1075 1173
rect 663 1139 1075 1147
rect 663 1111 695 1139
rect 663 1091 668 1111
rect 689 1091 695 1111
rect 663 1084 695 1091
rect 863 1111 913 1120
rect 1108 1119 1142 1325
rect 1676 1345 1708 1373
rect 1676 1325 1681 1345
rect 1702 1325 1708 1345
rect 1676 1318 1708 1325
rect 1883 1346 1925 1354
rect 2121 1353 2155 1559
rect 1883 1326 1892 1346
rect 1916 1326 1925 1346
rect 1883 1314 1925 1326
rect 2099 1348 2155 1353
rect 2099 1328 2106 1348
rect 2126 1328 2155 1348
rect 2099 1321 2155 1328
rect 2099 1320 2134 1321
rect 1885 1285 1920 1314
rect 1885 1284 2195 1285
rect 1770 1278 1806 1282
rect 1770 1259 1778 1278
rect 1798 1259 1806 1278
rect 1770 1256 1806 1259
rect 1771 1228 1805 1256
rect 1885 1250 2212 1284
rect 863 1090 875 1111
rect 897 1090 913 1111
rect 863 1082 913 1090
rect 1086 1114 1142 1119
rect 1086 1094 1093 1114
rect 1113 1094 1142 1114
rect 1086 1087 1142 1094
rect 1243 1200 1806 1228
rect 1086 1086 1121 1087
rect 868 1049 909 1082
rect 1243 1049 1283 1200
rect 868 1020 1283 1049
rect 2172 1026 2212 1250
rect 868 1019 1277 1020
rect 2172 1006 2182 1026
rect 2202 1006 2212 1026
rect 2172 996 2212 1006
rect 1731 933 1763 940
rect 1731 913 1738 933
rect 1759 913 1763 933
rect 1731 848 1763 913
rect 2101 848 2141 849
rect 1731 846 2143 848
rect 1731 820 2111 846
rect 2137 820 2143 846
rect 1731 812 2143 820
rect 1116 792 1148 793
rect 1113 787 1148 792
rect 1113 767 1120 787
rect 1140 767 1148 787
rect 1113 759 1148 767
rect 669 694 701 701
rect 669 674 676 694
rect 697 674 701 694
rect 669 609 701 674
rect 1039 609 1079 610
rect 669 607 1081 609
rect 669 581 1049 607
rect 1075 581 1081 607
rect 669 573 1081 581
rect 669 545 701 573
rect 1114 553 1148 759
rect 1731 784 1763 812
rect 1731 764 1736 784
rect 1757 764 1763 784
rect 1731 757 1763 764
rect 1942 783 1980 795
rect 2176 792 2210 996
rect 1942 766 1951 783
rect 1975 766 1980 783
rect 1942 723 1980 766
rect 2154 787 2210 792
rect 2154 767 2161 787
rect 2181 767 2210 787
rect 2154 760 2210 767
rect 2154 759 2189 760
rect 2288 723 2372 728
rect 1942 694 2372 723
rect 669 525 674 545
rect 695 525 701 545
rect 669 518 701 525
rect 878 547 918 552
rect 878 526 890 547
rect 912 526 918 547
rect 878 514 918 526
rect 1092 548 1148 553
rect 1092 528 1099 548
rect 1119 528 1148 548
rect 1092 521 1148 528
rect 1205 622 2162 641
rect 1092 520 1127 521
rect 884 482 912 514
rect 1205 482 1236 622
rect 2125 606 2160 622
rect 2125 586 2132 606
rect 2152 586 2160 606
rect 2125 578 2160 586
rect 884 451 1236 482
rect 1681 513 1713 520
rect 1681 493 1688 513
rect 1709 493 1713 513
rect 1681 428 1713 493
rect 2051 428 2091 429
rect 1681 426 2093 428
rect 1681 400 2061 426
rect 2087 400 2093 426
rect 1681 392 2093 400
rect 1115 377 1147 378
rect 1112 372 1147 377
rect 1112 352 1119 372
rect 1139 352 1147 372
rect 1112 344 1147 352
rect 668 279 700 286
rect 668 259 675 279
rect 696 259 700 279
rect 668 194 700 259
rect 1038 194 1078 195
rect 668 192 1080 194
rect 668 166 1048 192
rect 1074 166 1080 192
rect 668 158 1080 166
rect 668 130 700 158
rect 668 110 673 130
rect 694 110 700 130
rect 668 103 700 110
rect 868 130 918 139
rect 1113 138 1147 344
rect 1681 364 1713 392
rect 1681 344 1686 364
rect 1707 344 1713 364
rect 1886 366 1928 375
rect 2126 372 2160 578
rect 1886 352 1896 366
rect 1681 337 1713 344
rect 1885 346 1896 352
rect 1920 346 1928 366
rect 1885 335 1928 346
rect 2104 367 2160 372
rect 2104 347 2111 367
rect 2131 347 2160 367
rect 2104 340 2160 347
rect 2104 339 2139 340
rect 1885 305 1925 335
rect 1775 297 1811 301
rect 1775 278 1783 297
rect 1803 278 1811 297
rect 1775 275 1811 278
rect 1885 300 2232 305
rect 1776 247 1810 275
rect 1885 274 2204 300
rect 2223 274 2232 300
rect 1885 270 2232 274
rect 868 109 880 130
rect 902 109 918 130
rect 868 101 918 109
rect 1091 133 1147 138
rect 1091 113 1098 133
rect 1118 113 1147 133
rect 1091 106 1147 113
rect 1248 219 1811 247
rect 1091 105 1126 106
rect 873 68 914 101
rect 1248 68 1288 219
rect 2337 100 2372 694
rect 2337 94 2375 100
rect 2337 74 2347 94
rect 2367 74 2375 94
rect 2337 72 2375 74
rect 873 39 1288 68
rect 2340 66 2375 72
rect 873 38 1282 39
rect 1896 1 1928 8
rect 1896 -19 1903 1
rect 1924 -19 1928 1
rect 1896 -84 1928 -19
rect 2266 -84 2306 -83
rect 1896 -86 2308 -84
rect 1896 -112 2276 -86
rect 2302 -112 2308 -86
rect 1896 -120 2308 -112
rect 1896 -148 1928 -120
rect 2341 -140 2375 66
rect 1896 -168 1901 -148
rect 1922 -168 1928 -148
rect 1896 -175 1928 -168
rect 2319 -145 2375 -140
rect 2319 -165 2326 -145
rect 2346 -165 2375 -145
rect 2319 -172 2375 -165
rect 2319 -173 2354 -172
rect 1123 -187 1155 -186
rect 1120 -192 1155 -187
rect 1120 -212 1127 -192
rect 1147 -212 1155 -192
rect 1120 -220 1155 -212
rect 676 -285 708 -278
rect 676 -305 683 -285
rect 704 -305 708 -285
rect 676 -370 708 -305
rect 1046 -370 1086 -369
rect 676 -372 1088 -370
rect 676 -398 1056 -372
rect 1082 -398 1088 -372
rect 676 -406 1088 -398
rect 676 -434 708 -406
rect 1121 -426 1155 -220
rect 676 -454 681 -434
rect 702 -454 708 -434
rect 676 -461 708 -454
rect 885 -432 925 -427
rect 885 -453 897 -432
rect 919 -453 925 -432
rect 885 -465 925 -453
rect 1099 -431 1155 -426
rect 1099 -451 1106 -431
rect 1126 -451 1155 -431
rect 1099 -458 1155 -451
rect 1212 -357 2169 -338
rect 1099 -459 1134 -458
rect 891 -497 919 -465
rect 1212 -497 1243 -357
rect 2132 -373 2167 -357
rect 2132 -393 2139 -373
rect 2159 -393 2167 -373
rect 2132 -401 2167 -393
rect 891 -528 1243 -497
rect 1688 -466 1720 -459
rect 1688 -486 1695 -466
rect 1716 -486 1720 -466
rect 1688 -551 1720 -486
rect 2058 -551 2098 -550
rect 1688 -553 2100 -551
rect 1688 -579 2068 -553
rect 2094 -579 2100 -553
rect 1688 -587 2100 -579
rect 1122 -602 1154 -601
rect 1119 -607 1154 -602
rect 1119 -627 1126 -607
rect 1146 -627 1154 -607
rect 1119 -635 1154 -627
rect 675 -700 707 -693
rect 675 -720 682 -700
rect 703 -720 707 -700
rect 675 -785 707 -720
rect 1045 -785 1085 -784
rect 675 -787 1087 -785
rect 675 -813 1055 -787
rect 1081 -813 1087 -787
rect 675 -821 1087 -813
rect 675 -849 707 -821
rect 675 -869 680 -849
rect 701 -869 707 -849
rect 675 -876 707 -869
rect 875 -849 925 -840
rect 1120 -841 1154 -635
rect 1688 -615 1720 -587
rect 1688 -635 1693 -615
rect 1714 -635 1720 -615
rect 1688 -642 1720 -635
rect 1895 -614 1937 -606
rect 2133 -607 2167 -401
rect 1895 -634 1904 -614
rect 1928 -634 1937 -614
rect 1895 -646 1937 -634
rect 2111 -612 2167 -607
rect 2111 -632 2118 -612
rect 2138 -632 2167 -612
rect 2111 -639 2167 -632
rect 2111 -640 2146 -639
rect 1897 -675 1932 -646
rect 1897 -676 2207 -675
rect 1782 -682 1818 -678
rect 1782 -701 1790 -682
rect 1810 -701 1818 -682
rect 1782 -704 1818 -701
rect 1783 -732 1817 -704
rect 1897 -710 2224 -676
rect 875 -870 887 -849
rect 909 -870 925 -849
rect 875 -878 925 -870
rect 1098 -846 1154 -841
rect 1098 -866 1105 -846
rect 1125 -866 1154 -846
rect 1098 -873 1154 -866
rect 1255 -760 1818 -732
rect 1098 -874 1133 -873
rect 880 -911 921 -878
rect 1255 -911 1295 -760
rect 880 -940 1295 -911
rect 2184 -934 2224 -710
rect 880 -941 1289 -940
rect 2184 -954 2194 -934
rect 2214 -954 2224 -934
rect 2184 -964 2224 -954
rect 1743 -1027 1775 -1020
rect 1743 -1047 1750 -1027
rect 1771 -1047 1775 -1027
rect 1743 -1112 1775 -1047
rect 2113 -1112 2153 -1111
rect 1743 -1114 2155 -1112
rect 1743 -1140 2123 -1114
rect 2149 -1140 2155 -1114
rect 1743 -1148 2155 -1140
rect 1128 -1168 1160 -1167
rect 1125 -1173 1160 -1168
rect 1125 -1193 1132 -1173
rect 1152 -1193 1160 -1173
rect 1125 -1201 1160 -1193
rect 681 -1266 713 -1259
rect 681 -1286 688 -1266
rect 709 -1286 713 -1266
rect 681 -1351 713 -1286
rect 1051 -1351 1091 -1350
rect 681 -1353 1093 -1351
rect 681 -1379 1061 -1353
rect 1087 -1379 1093 -1353
rect 681 -1387 1093 -1379
rect 681 -1415 713 -1387
rect 1126 -1407 1160 -1201
rect 1743 -1176 1775 -1148
rect 2188 -1168 2222 -964
rect 1743 -1196 1748 -1176
rect 1769 -1196 1775 -1176
rect 1743 -1203 1775 -1196
rect 1954 -1176 1991 -1170
rect 1954 -1195 1960 -1176
rect 1983 -1195 1991 -1176
rect 1954 -1200 1991 -1195
rect 2166 -1173 2222 -1168
rect 2166 -1193 2173 -1173
rect 2193 -1193 2222 -1173
rect 2166 -1200 2222 -1193
rect 1962 -1237 1986 -1200
rect 2166 -1201 2201 -1200
rect 1962 -1239 2330 -1237
rect 1962 -1244 2335 -1239
rect 1962 -1262 2308 -1244
rect 2328 -1262 2335 -1244
rect 1962 -1267 2335 -1262
rect 2306 -1269 2335 -1267
rect 681 -1435 686 -1415
rect 707 -1435 713 -1415
rect 681 -1442 713 -1435
rect 890 -1413 930 -1408
rect 890 -1434 902 -1413
rect 924 -1434 930 -1413
rect 890 -1446 930 -1434
rect 1104 -1412 1160 -1407
rect 1104 -1432 1111 -1412
rect 1131 -1432 1160 -1412
rect 1104 -1439 1160 -1432
rect 1217 -1338 2174 -1319
rect 1104 -1440 1139 -1439
rect 896 -1478 924 -1446
rect 1217 -1478 1248 -1338
rect 2137 -1354 2172 -1338
rect 2137 -1374 2144 -1354
rect 2164 -1374 2172 -1354
rect 2137 -1382 2172 -1374
rect 896 -1509 1248 -1478
rect 1693 -1447 1725 -1440
rect 1693 -1467 1700 -1447
rect 1721 -1467 1725 -1447
rect 1693 -1532 1725 -1467
rect 2063 -1532 2103 -1531
rect 1693 -1534 2105 -1532
rect 1693 -1560 2073 -1534
rect 2099 -1560 2105 -1534
rect 1693 -1568 2105 -1560
rect 1127 -1583 1159 -1582
rect 1124 -1588 1159 -1583
rect 1124 -1608 1131 -1588
rect 1151 -1608 1159 -1588
rect 1124 -1616 1159 -1608
rect 680 -1681 712 -1674
rect 680 -1701 687 -1681
rect 708 -1701 712 -1681
rect 680 -1766 712 -1701
rect 1050 -1766 1090 -1765
rect 680 -1768 1092 -1766
rect 680 -1794 1060 -1768
rect 1086 -1794 1092 -1768
rect 680 -1802 1092 -1794
rect 680 -1830 712 -1802
rect 680 -1850 685 -1830
rect 706 -1850 712 -1830
rect 680 -1857 712 -1850
rect 880 -1830 930 -1821
rect 1125 -1822 1159 -1616
rect 1693 -1596 1725 -1568
rect 1693 -1616 1698 -1596
rect 1719 -1616 1725 -1596
rect 1898 -1594 1940 -1585
rect 2138 -1588 2172 -1382
rect 1898 -1608 1908 -1594
rect 1693 -1623 1725 -1616
rect 1897 -1614 1908 -1608
rect 1932 -1614 1940 -1594
rect 1897 -1625 1940 -1614
rect 2116 -1593 2172 -1588
rect 2116 -1613 2123 -1593
rect 2143 -1613 2172 -1593
rect 2116 -1620 2172 -1613
rect 2116 -1621 2151 -1620
rect 1897 -1655 1937 -1625
rect 1787 -1663 1823 -1659
rect 1787 -1682 1795 -1663
rect 1815 -1682 1823 -1663
rect 1787 -1685 1823 -1682
rect 1897 -1660 2244 -1655
rect 1788 -1713 1822 -1685
rect 1897 -1686 2216 -1660
rect 2235 -1686 2244 -1660
rect 1897 -1690 2244 -1686
rect 880 -1851 892 -1830
rect 914 -1851 930 -1830
rect 880 -1859 930 -1851
rect 1103 -1827 1159 -1822
rect 1103 -1847 1110 -1827
rect 1130 -1847 1159 -1827
rect 1103 -1854 1159 -1847
rect 1260 -1741 1823 -1713
rect 1103 -1855 1138 -1854
rect 885 -1892 926 -1859
rect 1260 -1892 1300 -1741
rect 885 -1921 1300 -1892
rect 885 -1922 1294 -1921
<< labels >>
rlabel locali 304 1752 333 1758 1 vdd
rlabel locali 517 1749 546 1755 1 vdd
rlabel locali 250 1564 272 1579 1 d0
rlabel nwell 671 1719 694 1722 1 vdd
rlabel locali 301 1453 330 1459 1 gnd
rlabel locali 514 1453 543 1459 1 gnd
rlabel space 611 1448 640 1457 1 gnd
rlabel locali 303 1337 332 1343 1 vdd
rlabel locali 516 1334 545 1340 1 vdd
rlabel locali 249 1149 271 1164 1 d0
rlabel nwell 670 1304 693 1307 1 vdd
rlabel locali 300 1038 329 1044 1 gnd
rlabel locali 513 1038 542 1044 1 gnd
rlabel space 610 1033 639 1042 1 gnd
rlabel locali 1316 1571 1345 1577 1 vdd
rlabel locali 1529 1568 1558 1574 1 vdd
rlabel nwell 1683 1538 1706 1541 1 vdd
rlabel locali 1313 1272 1342 1278 1 gnd
rlabel locali 1526 1272 1555 1278 1 gnd
rlabel space 1623 1267 1652 1276 1 gnd
rlabel locali 1254 1382 1301 1403 1 d1
rlabel locali 116 1944 141 1953 1 vref
rlabel locali 309 771 338 777 1 vdd
rlabel locali 522 768 551 774 1 vdd
rlabel locali 255 583 277 598 1 d0
rlabel nwell 676 738 699 741 1 vdd
rlabel locali 306 472 335 478 1 gnd
rlabel locali 519 472 548 478 1 gnd
rlabel space 616 467 645 476 1 gnd
rlabel locali 308 356 337 362 1 vdd
rlabel locali 521 353 550 359 1 vdd
rlabel locali 254 168 276 183 1 d0
rlabel nwell 675 323 698 326 1 vdd
rlabel locali 305 57 334 63 1 gnd
rlabel locali 518 57 547 63 1 gnd
rlabel locali 1321 590 1350 596 1 vdd
rlabel locali 1534 587 1563 593 1 vdd
rlabel nwell 1688 557 1711 560 1 vdd
rlabel locali 1318 291 1347 297 1 gnd
rlabel locali 1531 291 1560 297 1 gnd
rlabel space 1628 286 1657 295 1 gnd
rlabel locali 1259 401 1306 422 1 d1
rlabel locali 1371 1010 1400 1016 1 vdd
rlabel locali 1584 1007 1613 1013 1 vdd
rlabel nwell 1738 977 1761 980 1 vdd
rlabel locali 1368 711 1397 717 1 gnd
rlabel locali 1581 711 1610 717 1 gnd
rlabel space 1678 706 1707 715 1 gnd
rlabel locali 1314 822 1337 837 1 d2
rlabel space 615 52 644 61 1 gnd
rlabel locali 1326 -1138 1349 -1123 1 d2
rlabel space 1690 -1254 1719 -1245 1 gnd
rlabel locali 1593 -1249 1622 -1243 1 gnd
rlabel locali 1380 -1249 1409 -1243 1 gnd
rlabel nwell 1750 -983 1773 -980 1 vdd
rlabel locali 1596 -953 1625 -947 1 vdd
rlabel locali 1383 -950 1412 -944 1 vdd
rlabel locali 138 -1952 165 -1939 1 gnd
rlabel locali 1271 -1559 1318 -1538 1 d1
rlabel space 1640 -1674 1669 -1665 1 gnd
rlabel locali 1543 -1669 1572 -1663 1 gnd
rlabel locali 1330 -1669 1359 -1663 1 gnd
rlabel nwell 1700 -1403 1723 -1400 1 vdd
rlabel locali 1546 -1373 1575 -1367 1 vdd
rlabel locali 1333 -1370 1362 -1364 1 vdd
rlabel space 627 -1908 656 -1899 1 gnd
rlabel locali 530 -1903 559 -1897 1 gnd
rlabel locali 317 -1903 346 -1897 1 gnd
rlabel nwell 687 -1637 710 -1634 1 vdd
rlabel locali 266 -1792 288 -1777 1 d0
rlabel locali 533 -1607 562 -1601 1 vdd
rlabel locali 320 -1604 349 -1598 1 vdd
rlabel space 628 -1493 657 -1484 1 gnd
rlabel locali 531 -1488 560 -1482 1 gnd
rlabel locali 318 -1488 347 -1482 1 gnd
rlabel nwell 688 -1222 711 -1219 1 vdd
rlabel locali 267 -1377 289 -1362 1 d0
rlabel locali 534 -1192 563 -1186 1 vdd
rlabel locali 321 -1189 350 -1183 1 vdd
rlabel locali 1266 -578 1313 -557 1 d1
rlabel space 1635 -693 1664 -684 1 gnd
rlabel locali 1538 -688 1567 -682 1 gnd
rlabel locali 1325 -688 1354 -682 1 gnd
rlabel nwell 1695 -422 1718 -419 1 vdd
rlabel locali 1541 -392 1570 -386 1 vdd
rlabel locali 1328 -389 1357 -383 1 vdd
rlabel space 622 -927 651 -918 1 gnd
rlabel locali 525 -922 554 -916 1 gnd
rlabel locali 312 -922 341 -916 1 gnd
rlabel nwell 682 -656 705 -653 1 vdd
rlabel locali 261 -811 283 -796 1 d0
rlabel locali 528 -626 557 -620 1 vdd
rlabel locali 315 -623 344 -617 1 vdd
rlabel space 623 -512 652 -503 1 gnd
rlabel locali 526 -507 555 -501 1 gnd
rlabel locali 313 -507 342 -501 1 gnd
rlabel nwell 683 -241 706 -238 1 vdd
rlabel locali 262 -396 284 -381 1 d0
rlabel locali 529 -211 558 -205 1 vdd
rlabel locali 316 -208 345 -202 1 vdd
rlabel locali 1536 78 1565 84 1 vdd
rlabel locali 1749 75 1778 81 1 vdd
rlabel locali 2112 -75 2134 -60 1 vout
rlabel nwell 1903 45 1926 48 1 vdd
rlabel locali 1533 -221 1562 -215 1 gnd
rlabel locali 1746 -221 1775 -215 1 gnd
rlabel space 1843 -226 1872 -217 1 gnd
rlabel locali 1474 -112 1506 -93 1 d3
<< end >>
