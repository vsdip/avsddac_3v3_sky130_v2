* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******* SkyWater sky130 model library *********

* Typical corner (tt)
.lib tt
* MOSFET
.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice"
* Mismatch parameters
.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice"
* All models
.include "all.spice"
.endl


* Slow-Fast corner (sf)
.lib sf
* MOSFET
.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__sf.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__sf.corner.spice"
* Mismatch parameters
.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice"
* All models
.include "all.spice"
.endl


* Fast-Fast corner (ff)
.lib ff
* MOSFET
.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__ff.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__ff.corner.spice"
* Mismatch parameters
.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice"
* All models
.include "all.spice"
.endl


* Slow-Slow corner (ss)
.lib ss
* MOSFET
.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__ss.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__ss.corner.spice"
* Mismatch parameters
.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice"
* All models
.include "all.spice"
.endl


* Fast-Slow corner (fs)
.lib fs
* MOSFET
.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__fs.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__fs.corner.spice"
* Mismatch parameters
.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice"
* All models
.include "all.spice"
.endl
