* SPICE3 file created from 8bit_DAC.ext - technology: sky130A

.option scale=10000u

X0 gnd a_40764_12735# a_40556_12735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1 vdd d0 a_20139_11965# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2 a_984_9065# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X3 a_40508_8511# a_41605_8317# a_41560_8330# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X4 a_22657_8384# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X5 gnd d0 a_41812_12731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X6 a_981_7471# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X7 a_30848_9192# a_30852_8336# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8 a_40512_8334# a_40765_8321# a_39061_9191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X9 a_22869_12798# a_22656_12798# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X10 a_11692_8380# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X11 a_12953_9055# a_12740_9055# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X12 a_11690_3051# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X13 a_25150_3818# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X14 a_32955_2478# a_33576_2370# a_33784_2370# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X15 a_22246_7804# a_22870_8384# a_23078_8384# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X16 a_18839_9783# a_19932_10445# a_19883_10635# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X17 a_41557_6736# a_41553_6913# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X18 a_1194_6792# a_981_6792# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X19 a_9178_11305# a_9431_11292# a_8126_11486# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X20 a_11689_6786# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X21 vdd a_31105_9002# a_30897_9002# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X22 a_39022_10459# a_39109_11968# a_39064_11981# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X23 a_24126_10506# a_23705_10506# a_23078_10510# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X24 a_34412_13467# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X25 a_8131_8342# a_9224_9004# a_9179_9017# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X26 gnd a_19089_6729# a_18881_6729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X27 a_25151_12793# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X28 gnd d2 a_28609_11974# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X29 a_9173_3954# a_9177_3009# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X30 vdd a_40764_12735# a_40556_12735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X31 gnd a_31103_2315# a_30895_2315# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X32 vdd d0 a_41812_12731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X33 a_30847_12159# a_30851_11303# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X34 a_14650_11344# a_14229_11344# a_14556_11463# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X35 a_19886_11978# a_19882_12155# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X36 a_30851_11982# a_31104_11969# a_29803_11307# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X37 a_8125_2511# a_9222_2317# a_9173_2507# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X38 a_40508_8511# a_40765_8321# a_39061_9191# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X39 vdd d0 a_20138_3758# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X40 gnd a_9432_10451# a_9224_10451# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X41 a_9178_13431# a_9174_13608# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X42 a_12953_10502# a_12740_10502# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X43 a_39016_4628# a_39108_2993# a_39059_3183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X44 a_33365_10504# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X45 a_982_2378# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X46 a_14184_6781# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X47 a_13160_12022# a_12739_12022# a_12112_12026# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X48 a_41560_9009# a_41813_8996# a_40512_8334# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X49 a_18839_9783# a_19932_10445# a_19887_10458# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X50 a_32956_12900# a_33577_12792# a_33785_12792# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X51 a_22867_6022# a_22654_6022# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X52 a_40507_12925# a_41604_12731# a_41555_12921# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X53 a_24124_3051# a_23703_3051# a_23076_2376# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X54 a_23075_7469# a_22654_7469# a_22246_7548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X55 gnd d0 a_41811_3756# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X56 a_11904_12794# a_11691_12794# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X57 a_11902_6018# a_11689_6018# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X58 a_576_8494# a_1197_8386# a_1405_8386# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X59 a_9177_4456# a_9430_4443# a_8129_3781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X60 a_25194_11348# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X61 a_3477_3820# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X62 a_19883_10635# a_19887_9779# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X63 vdd a_31103_2315# a_30895_2315# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X64 a_33783_5337# a_34623_6012# a_34831_6012# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X65 a_1402_5345# a_981_5345# a_573_5453# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X66 a_18837_3775# a_19090_3762# a_17390_3008# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X67 a_6683_11989# a_6936_11976# a_6641_10467# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X68 a_14398_3814# a_14185_3814# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X69 a_30845_6919# a_30849_5974# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X70 a_33786_8378# a_33365_8378# a_32957_8486# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X71 gnd d0 a_20139_11286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X72 a_36115_11342# a_35902_11342# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X73 vdd a_9432_10451# a_9224_10451# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X74 gnd a_40763_3760# a_40555_3760# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X75 a_33783_6784# a_33362_6784# a_32954_6351# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X76 vdd a_19091_12737# a_18883_12737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X77 gnd a_41812_13410# a_41604_13410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X78 a_28314_10465# a_28401_11974# a_28352_12164# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X79 vdd a_30056_11294# a_29848_11294# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X80 a_29802_2332# a_30895_2994# a_30846_3184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X81 a_11283_13552# a_11904_13473# a_12112_13473# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X82 a_9172_6921# a_9176_5976# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X83 a_40507_12925# a_41604_12731# a_41559_12744# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X84 vdd d0 a_41811_3756# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X85 a_32956_11708# a_32956_11453# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X86 a_573_7806# a_573_7550# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X87 gnd a_27499_7417# a_27291_7417# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X88 vdd d1 a_40764_11288# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X89 gnd a_20140_8998# a_19932_8998# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X90 a_16277_7603# a_17392_4440# a_17343_4630# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X91 a_41558_2322# a_41811_2309# a_40506_2503# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X92 a_573_7155# a_1194_7471# a_1402_7471# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X93 a_11905_9827# a_11692_9827# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X94 a_9173_4633# a_9430_4443# a_8129_3781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X95 a_32957_9392# a_32957_9136# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X96 a_14440_5336# a_14227_5336# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X97 a_30849_6742# a_31102_6729# a_29797_6923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X98 a_22248_11459# a_22869_11351# a_23077_11351# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X99 a_18833_3952# a_19090_3762# a_17390_3008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X100 a_34834_10500# a_36073_9820# a_36224_11342# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X101 a_13160_13469# a_14399_12789# a_14556_11463# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X102 a_29800_8517# a_30897_8323# a_30848_8513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X103 vdd d0 a_20139_11286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X104 vdd a_40763_3760# a_40555_3760# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X105 vdd a_20138_3758# a_19930_3758# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X106 a_1402_7471# a_2242_7467# a_2450_7467# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X107 a_39059_3183# a_40555_2313# a_40506_2503# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X108 a_25149_6785# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X109 a_12952_13469# a_12739_13469# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X110 vdd a_41812_13410# a_41604_13410# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X111 gnd d1 a_40762_5280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X112 a_18832_6919# a_19929_6725# a_19880_6915# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X113 a_576_9144# a_576_8749# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X114 a_11282_3130# a_11903_3051# a_12111_3051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X115 a_11281_6894# a_11902_6786# a_12110_6786# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X116 a_22654_6022# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X117 a_1405_9065# a_984_9065# a_576_8749# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X118 a_14400_9822# a_14187_9822# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X119 a_574_4188# a_574_3933# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X120 a_16277_7603# a_17392_4440# a_17347_4453# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X121 a_983_12032# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X122 a_30846_3184# a_31103_2994# a_29802_2332# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X123 gnd a_28608_2999# a_28400_2999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X124 a_32955_4831# a_33575_5337# a_33783_5337# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X125 a_1194_6024# a_981_6024# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X126 a_11691_13473# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X127 a_11281_7544# a_11281_7149# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X128 a_1404_12800# a_983_12800# a_575_12908# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X129 a_33578_9057# a_33365_9057# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X130 a_1404_12800# a_2244_13475# a_2452_13475# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X131 a_33575_7463# a_33362_7463# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X132 a_39060_12158# a_40556_11288# a_40511_11301# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X133 a_29800_8517# a_30897_8323# a_30852_8336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X134 a_2450_6020# a_2029_6020# a_1402_5345# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X135 a_14185_3814# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X136 a_39059_3183# a_40555_2313# a_40510_2326# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X137 a_22247_4186# a_22868_4502# a_23076_4502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X138 a_22656_11351# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X139 a_28350_6156# a_29846_5286# a_29797_5476# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X140 a_41557_5968# a_41553_6145# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X141 vdd d1 a_40762_5280# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X142 a_18832_6919# a_19929_6725# a_19884_6738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X143 a_5353_4506# a_4932_4506# a_5008_8377# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X144 a_40510_2326# a_41603_2988# a_41554_3178# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X145 a_23078_9063# a_23918_9059# a_24126_9059# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X146 a_22657_9831# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X147 a_30847_11480# a_30852_10462# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X148 a_11692_9827# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X149 a_32956_11708# a_33577_12024# a_33785_12024# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X150 a_1403_2378# a_982_2378# a_576_2387# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X151 a_24123_6018# a_23702_6018# a_23075_6022# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X152 a_9178_11305# a_9174_11482# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X153 vdd d1 a_8381_5288# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X154 a_11904_12026# a_11691_12026# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X155 a_34413_10500# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X156 a_1197_9833# a_984_9833# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X157 a_19881_4627# a_20138_4437# a_18837_3775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X158 vdd d0 a_20140_8319# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X159 a_23916_3051# a_23703_3051# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X160 a_22867_7469# a_22654_7469# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X161 a_573_6103# a_1194_6024# a_1402_6024# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X162 a_33576_2370# a_33363_2370# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X163 vdd d1 a_8382_3768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X164 a_40508_8511# a_41605_8317# a_41556_8507# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X165 a_32955_3384# a_32955_3128# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X166 a_28350_6156# a_29846_5286# a_29801_5299# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X167 a_32957_9136# a_33578_9057# a_33786_9057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X168 a_12740_10502# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X169 gnd d1 a_19089_5282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X170 a_12113_9059# a_12953_9055# a_13161_9055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X171 a_33783_6016# a_33362_6016# a_32954_6095# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X172 a_30851_13429# a_31104_13416# a_29803_12754# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X173 a_575_11716# a_1196_12032# a_1404_12032# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X174 a_17345_10638# a_17602_10448# a_16281_7426# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X175 a_17390_3008# a_18882_3762# a_18833_3952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X176 a_13158_6014# a_12737_6014# a_12110_6018# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X177 a_22870_9063# a_22657_9063# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X178 vdd a_17643_2995# a_17435_2995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X179 a_12112_11347# a_11691_11347# a_11284_10841# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X180 a_982_3825# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X181 vdd d2 a_6935_3001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X182 vdd d2 a_17644_11970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X183 a_33365_9057# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X184 a_9174_12929# a_9431_12739# a_8126_12933# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X185 a_36222_5334# a_35858_3812# a_34832_3045# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X186 gnd a_9430_2996# a_9222_2996# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X187 a_33362_7463# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X188 a_19882_12155# a_20139_11965# a_18838_11303# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X189 a_576_10196# a_576_9941# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X190 a_30845_7598# a_30849_6742# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X191 a_33786_8378# a_34626_9053# a_34834_9053# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X192 a_29803_11307# a_30896_11969# a_30851_11982# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X193 a_576_9941# a_1197_9833# a_1405_9833# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X194 vdd a_9431_11292# a_9223_11292# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X195 vdd d1 a_19089_5282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X196 a_8130_11309# a_9223_11971# a_9174_12161# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X197 gnd d2 a_17643_2995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X198 gnd d0 a_20138_3758# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X199 a_9172_7600# a_9176_6744# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X200 a_30851_13429# a_30847_13606# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X201 a_1404_12032# a_2244_12028# a_2452_12028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X202 a_11284_10585# a_11905_10506# a_12113_10506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X203 a_1402_6792# a_981_6792# a_573_6900# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X204 a_1195_3057# a_982_3057# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X205 gnd d0 a_31102_5961# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X206 a_30847_13606# a_31104_13416# a_29803_12754# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X207 a_17390_3008# a_18882_3762# a_18837_3775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X208 a_41560_9009# a_41556_9186# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X209 a_33786_9825# a_33365_9825# a_32957_9933# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X210 gnd d0 a_20139_12733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X211 a_11015_219# a_15640_4500# a_15962_4500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X212 a_29800_8517# a_30057_8327# a_28353_9197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X213 a_36321_5334# a_35900_5334# a_36222_5334# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X214 a_11281_5702# a_11902_6018# a_12110_6018# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X215 a_29802_3779# a_30895_4441# a_30846_4631# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X216 a_22246_7548# a_22246_7153# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X217 a_30852_9015# a_31105_9002# a_29804_8340# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X218 a_19880_6147# a_20137_5957# a_18836_5295# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X219 a_575_13163# a_575_12908# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X220 a_22654_7469# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X221 a_23703_3051# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X222 a_34833_12020# a_34412_12020# a_33785_11345# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X223 vdd a_39317_11968# a_39109_11968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X224 a_41558_3769# a_41811_3756# a_40506_3950# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X225 a_33363_2370# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X226 a_33785_13471# a_33364_13471# a_32956_13155# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X227 a_36072_12787# a_35859_12787# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X228 a_17349_10461# a_17436_11970# a_17391_11983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X229 gnd d3 a_6892_4446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X230 a_34623_6012# a_34410_6012# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X231 gnd a_19091_12737# a_18883_12737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X232 a_2243_3053# a_2030_3053# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X233 a_11281_5447# a_11282_4833# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X234 a_39016_4628# a_39273_4438# a_37950_7601# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X235 a_36321_5334# a_37181_8369# a_37389_8369# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X236 a_30849_6742# a_30845_6919# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X237 vdd d0 a_20139_12733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X238 a_32956_11453# a_32957_10839# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X239 a_18835_9960# a_19932_9766# a_19883_9956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X240 gnd d0 a_31105_9770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X241 a_37526_4498# a_37313_4498# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X242 a_34624_4492# a_34411_4492# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X243 a_2450_7467# a_2029_7467# a_1402_7471# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X244 a_3942_11350# a_3521_11350# a_3843_11350# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X245 a_29802_3779# a_30895_4441# a_30850_4454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X246 a_23075_6790# a_22654_6790# a_22246_6357# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X247 a_25613_5340# a_25192_5340# a_25519_5459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X248 a_6639_4459# a_6726_5968# a_6677_6158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X249 a_9176_6744# a_9172_6921# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X250 vdd a_6935_3001# a_6727_3001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X251 a_12111_3051# a_11690_3051# a_11282_3130# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X252 a_14554_5455# a_14184_6781# a_13158_6014# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X253 a_11692_10506# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X254 a_19884_5291# a_19880_5468# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X255 a_26473_8375# a_26260_8375# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X256 a_23917_13473# a_23704_13473# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X257 a_41556_9186# a_41560_8330# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X258 a_1405_9833# a_2245_10508# a_2453_10508# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X259 a_41554_3946# a_41811_3756# a_40506_3950# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X260 a_27026_4504# a_32579_217# a_21652_206# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X261 a_32954_7542# a_32954_7147# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X262 a_19886_11299# a_20139_11286# a_18834_11480# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X263 a_32954_6351# a_33575_6784# a_33783_6784# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X264 vdd d3 a_6892_4446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X265 a_29799_11484# a_30896_11290# a_30847_11480# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X266 a_33784_3049# a_33363_3049# a_32955_2733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X267 gnd a_20138_3758# a_19930_3758# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X268 vdd d0 a_9431_11971# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X269 a_6677_6158# a_8173_5288# a_8128_5301# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X270 a_575_12908# a_575_12367# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X271 a_13159_3047# a_12738_3047# a_12111_2372# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X272 a_23915_6018# a_23702_6018# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X273 a_41554_3946# a_41558_3001# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X274 vdd d0 a_9430_2317# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X275 gnd a_31102_5961# a_30894_5961# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X276 a_18835_9960# a_19932_9766# a_19887_9779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X277 vdd d0 a_31105_9770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X278 a_36224_11342# a_36115_11342# a_36323_11342# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X279 a_8128_5301# a_9221_5963# a_9172_6153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X280 a_23077_12030# a_22656_12030# a_22248_11714# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X281 a_9175_8515# a_9176_7423# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X282 a_14442_11344# a_14229_11344# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X283 a_6682_3014# a_8174_3768# a_8129_3781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X284 a_39020_4451# a_39107_5960# a_39062_5973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X285 a_3848_11469# a_3478_12795# a_2452_12028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X286 a_28354_5979# a_29846_6733# a_29797_6923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X287 vdd d1 a_40762_6727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X288 a_19883_9188# a_20140_8998# a_18839_8336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X289 gnd a_17645_9003# a_17437_9003# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X290 gnd a_20140_10445# a_19932_10445# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X291 a_40510_3773# a_41603_4435# a_41554_4625# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X292 a_25364_12793# a_25151_12793# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X293 a_40509_5293# a_40762_5280# a_39058_6150# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X294 gnd d0 a_41810_7402# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X295 a_19882_11476# a_20139_11286# a_18834_11480# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X296 a_34832_3045# a_34411_3045# a_33784_3049# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X297 a_1403_3825# a_982_3825# a_574_3392# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X298 a_22247_4837# a_22867_5343# a_23075_5343# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X299 a_41559_11976# a_41812_11963# a_40511_11301# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X300 a_21330_206# d7 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X301 a_34410_6012# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X302 gnd a_6892_4446# a_6684_4446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X303 gnd d2 a_28607_5966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X304 a_25365_9826# a_25152_9826# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X305 a_30848_9960# a_30852_9015# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X306 gnd a_41811_2988# a_41603_2988# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X307 gnd a_31105_9770# a_30897_9770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X308 a_33576_3817# a_33363_3817# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X309 a_34411_4492# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X310 a_37313_4498# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X311 a_28354_5979# a_29846_6733# a_29801_6746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X312 a_8127_9966# a_9224_9772# a_9175_9962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X313 a_29801_5299# a_30894_5961# a_30849_5974# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X314 vdd a_20140_10445# a_19932_10445# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X315 a_40510_3773# a_41603_4435# a_41558_4448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X316 a_13161_9055# a_12740_9055# a_12113_9059# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X317 a_11284_9394# a_11284_9138# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X318 a_19883_8509# a_19884_7417# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X319 a_26260_8375# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X320 a_28352_12164# a_29848_11294# a_29803_11307# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X321 a_40505_5470# a_40762_5280# a_39058_6150# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X322 a_2032_9061# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X323 a_35902_11342# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X324 a_30851_11303# a_30847_11480# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X325 a_19880_5468# a_20137_5278# a_18832_5472# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X326 a_574_2741# a_574_2486# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X327 a_19885_4450# a_20138_4437# a_18837_3775# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X328 gnd d0 a_20140_8319# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X329 a_12739_13469# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X330 a_15853_4500# a_15640_4500# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X331 vdd a_31104_11290# a_30896_11290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X332 vdd a_6892_4446# a_6684_4446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X333 gnd d1 a_8382_3768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X334 a_12110_5339# a_11689_5339# a_11282_4833# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X335 a_33364_13471# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X336 a_23917_12026# a_23704_12026# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X337 a_28352_12164# a_28609_11974# a_28314_10465# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X338 a_23702_6018# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X339 vdd a_40764_11288# a_40556_11288# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X340 a_36071_3812# a_35858_3812# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X341 gnd a_9430_4443# a_9222_4443# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X342 a_22246_5451# a_22247_4837# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X343 gnd d0 a_9431_11292# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X344 a_22869_13477# a_22656_13477# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X345 a_39018_10636# a_39110_9001# a_39065_9014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X346 vdd a_31105_9770# a_30897_9770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X347 a_32957_9933# a_32957_9392# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X348 a_33577_11345# a_33364_11345# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X349 a_8127_9966# a_9224_9772# a_9179_9785# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X350 a_17349_10461# a_17602_10448# a_16281_7426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X351 gnd a_19090_3762# a_18882_3762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X352 vdd d1 a_19089_6729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X353 a_16281_7426# a_16534_7413# a_15962_4500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X354 a_22249_9142# a_22870_9063# a_23078_9063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X355 a_34833_13467# a_34412_13467# a_33785_13471# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X356 a_8131_9789# a_8384_9776# a_6684_9022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X357 a_19881_4627# a_19885_3771# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X358 a_11689_7465# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X359 a_25521_11467# a_25151_12793# a_24125_13473# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X360 a_11284_8743# a_11905_9059# a_12113_9059# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X361 a_11283_12105# a_11283_11710# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X362 a_34623_7459# a_34410_7459# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X363 a_32955_3925# a_33576_3817# a_33784_3817# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X364 a_1195_4504# a_982_4504# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X365 a_23075_6022# a_22654_6022# a_22246_6101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X366 a_9178_12752# a_9431_12739# a_8126_12933# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X367 gnd d0 a_31104_11969# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X368 vdd a_28607_5966# a_28399_5966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X369 a_30849_5974# a_30845_6151# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X370 a_33786_10504# a_33365_10504# a_32957_10188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X371 a_22867_6790# a_22654_6790# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X372 a_4587_8377# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X373 a_6678_3191# a_6935_3001# a_6635_4636# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X374 vdd a_9430_4443# a_9222_4443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X375 a_1196_11353# a_983_11353# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X376 a_11903_3051# a_11690_3051# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X377 a_25152_9826# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X378 a_14648_5336# a_14227_5336# a_14549_5336# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X379 a_9176_5976# a_9172_6153# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X380 a_15508_8371# a_15295_8371# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X381 a_35858_3812# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X382 a_574_4583# a_574_4188# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X383 a_16277_7603# a_16534_7413# a_15962_4500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X384 vdd a_19090_3762# a_18882_3762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X385 a_33363_3817# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X386 gnd d1 a_30055_3766# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X387 a_11282_3927# a_11282_3386# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X388 a_12737_7461# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X389 a_8130_12756# a_9223_13418# a_9178_13431# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X390 a_36229_11461# a_35859_12787# a_34833_12020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X391 a_22870_10510# a_22657_10510# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X392 a_8127_9966# a_8384_9776# a_6684_9022# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X393 a_29804_8340# a_30057_8327# a_28353_9197# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X394 a_37954_7424# a_39067_10446# a_39018_10636# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X395 a_40509_5293# a_41602_5955# a_41557_5968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X396 a_25615_11348# a_25194_11348# a_25521_11467# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X397 a_29797_5476# a_30894_5282# a_30845_5472# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X398 a_2029_6020# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X399 a_17390_3008# a_17643_2995# a_17343_4630# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X400 vdd d0 a_31102_7408# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X401 vdd d0 a_41811_2309# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X402 a_18838_11303# a_19931_11965# a_19882_12155# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X403 a_22247_2484# a_22868_2376# a_23076_2376# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X404 a_23918_10506# a_23705_10506# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X405 a_18838_11303# a_19091_11290# a_17387_12160# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X406 a_23078_9831# a_22657_9831# a_22249_9939# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X407 a_575_12111# a_575_11716# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X408 a_1405_10512# a_984_10512# a_576_10196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X409 a_19885_3771# a_19881_3948# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X410 a_24125_12026# a_23704_12026# a_23077_12030# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X411 a_14551_11344# a_14187_9822# a_13161_10502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X412 a_32579_217# a_32366_217# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X413 a_22246_7804# a_22246_7548# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X414 a_23077_13477# a_22656_13477# a_22248_13556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X415 a_35900_5334# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X416 a_984_8386# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X417 a_10693_219# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X418 a_29803_11307# a_30056_11294# a_28352_12164# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X419 a_39020_4451# a_39273_4438# a_37950_7601# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X420 gnd d4 a_38207_7411# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X421 a_30850_3775# a_31103_3762# a_29798_3956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X422 vdd d1 a_30055_3766# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X423 a_28312_4457# a_28399_5966# a_28354_5979# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X424 a_19886_12746# a_20139_12733# a_18834_12927# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X425 a_37954_7424# a_39067_10446# a_39022_10459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X426 a_1402_6024# a_2242_6020# a_2450_6020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X427 a_12952_12022# a_12739_12022# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X428 a_39065_9014# a_40557_9768# a_40512_9781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X429 a_29797_5476# a_30894_5282# a_30849_5295# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X430 a_33364_12024# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X431 a_4932_4506# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X432 a_9174_12161# a_9178_11305# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X433 a_37181_8369# a_36968_8369# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X434 a_22249_9398# a_22249_9142# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X435 a_3479_9828# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X436 a_34410_7459# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X437 a_8128_6748# a_9221_7410# a_9172_7600# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X438 a_16281_7426# a_17394_10448# a_17349_10461# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X439 a_981_7471# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X440 vdd d0 a_9432_9004# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X441 a_22654_6790# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X442 a_32956_12900# a_32956_12359# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X443 a_22247_4186# a_22247_3931# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X444 vdd a_9429_5963# a_9221_5963# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X445 a_12953_9055# a_12740_9055# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X446 a_11690_3051# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X447 a_36224_11342# a_35860_9820# a_34834_10500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X448 a_575_11716# a_575_11461# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X449 vdd d4 a_38207_7411# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X450 a_12950_7461# a_12737_7461# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X451 a_8126_11486# a_8383_11296# a_6679_12166# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X452 a_30846_3952# a_31103_3762# a_29798_3956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X453 a_19882_12923# a_20139_12733# a_18834_12927# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X454 gnd d0 a_9430_2317# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X455 a_34832_4492# a_34411_4492# a_33784_4496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X456 a_15295_8371# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X457 gnd d2 a_28610_9007# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X458 vdd a_17644_11970# a_17436_11970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X459 a_3690_3820# a_3477_3820# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X460 vdd d2 a_17642_5962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X461 gnd a_41812_13410# a_40511_12748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X462 a_29799_12931# a_30896_12737# a_30851_12750# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X463 gnd a_30055_3766# a_29847_3766# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X464 a_23076_3055# a_22655_3055# a_22247_2739# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X465 gnd d2 a_39316_2993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X466 a_6682_3014# a_8174_3768# a_8125_3958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X467 a_13158_6014# a_14397_6781# a_14554_5455# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X468 gnd d0 a_20137_7404# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X469 a_11902_5339# a_11689_5339# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X470 gnd d1 a_40762_6727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X471 vdd a_31102_7408# a_30894_7408# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X472 a_40505_5470# a_41602_5276# a_41553_5466# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X473 gnd a_41811_4435# a_41603_4435# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X474 a_8128_6748# a_9221_7410# a_9176_7423# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X475 vdd a_6936_11976# a_6728_11976# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X476 a_12737_6014# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X477 a_1404_13479# a_983_13479# a_575_13163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X478 a_32957_9136# a_32957_8741# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X479 a_40505_6917# a_40762_6727# a_39062_5973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X480 a_12738_4494# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X481 a_33365_10504# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X482 a_26681_8375# a_26818_4504# a_27026_4504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X483 a_11284_10190# a_11284_9935# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X484 a_32955_4180# a_32955_3925# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X485 a_22867_6022# a_22654_6022# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X486 gnd a_38207_7411# a_37999_7411# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X487 a_41555_13600# a_41812_13410# a_40511_12748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X488 vdd a_30055_3766# a_29847_3766# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X489 a_24124_3051# a_23703_3051# a_23076_3055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X490 a_41557_7415# a_41810_7402# a_40509_6740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X491 a_22247_3931# a_22247_3390# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X492 a_34834_10500# a_34413_10500# a_33786_10504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X493 vdd a_41811_4435# a_41603_4435# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X494 a_40505_5470# a_41602_5276# a_41557_5289# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X495 gnd d3 a_6894_10454# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X496 a_573_6900# a_1194_6792# a_1402_6792# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X497 a_28354_5979# a_28607_5966# a_28312_4457# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X498 gnd d2 a_6937_9009# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X499 a_19884_5291# a_20137_5278# a_18832_5472# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X500 a_574_2486# a_576_2387# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X501 a_14398_3814# a_14185_3814# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X502 a_19887_8332# a_19883_8509# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X503 vdd a_9432_9004# a_9224_9004# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X504 a_15716_8371# a_15853_4500# a_11015_219# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X505 a_17345_10638# a_17437_9003# a_17392_9016# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X506 a_24125_13473# a_25364_12793# a_25521_11467# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X507 a_36227_5453# a_36113_5334# a_36321_5334# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X508 a_28314_10465# a_28567_10452# a_27246_7430# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X509 a_11282_3130# a_11282_2735# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X510 vdd a_38207_7411# a_37999_7411# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X511 a_11283_13157# a_11904_13473# a_12112_13473# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X512 a_30850_4454# a_30846_4631# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X513 gnd a_9429_5284# a_9221_5284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X514 gnd d0 a_31104_13416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X515 a_5353_4506# a_10906_219# a_11114_219# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X516 a_981_6024# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X517 a_25405_5340# a_25192_5340# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X518 gnd a_39316_2993# a_39108_2993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X519 gnd d0 a_20138_2311# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X520 a_9177_4456# a_9173_4633# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X521 gnd d1 a_19089_6729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X522 gnd a_20137_7404# a_19929_7404# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X523 a_1196_12800# a_983_12800# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X524 vdd d0 a_9431_12739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X525 a_983_11353# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X526 vdd d3 a_6894_10454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X527 a_19885_3003# a_19881_3180# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X528 a_14440_5336# a_14227_5336# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X529 a_22249_10845# a_22869_11351# a_23077_11351# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X530 a_1194_5345# a_981_5345# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X531 a_32688_217# a_37313_4498# a_37635_4498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X532 a_33578_8378# a_33365_8378# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X533 a_23078_10510# a_22657_10510# a_22249_10589# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X534 a_18837_2328# a_19930_2990# a_19881_3180# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X535 a_34412_12020# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X536 a_28310_10642# a_28567_10452# a_27246_7430# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X537 a_1402_6792# a_2242_7467# a_2450_7467# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X538 a_18838_12750# a_19931_13412# a_19882_13602# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X539 a_22247_3931# a_22868_3823# a_23076_3823# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X540 vdd a_9429_5284# a_9221_5284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X541 vdd d0 a_31104_13416# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X542 a_11282_2735# a_11903_3051# a_12111_3051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X543 a_13159_4494# a_14398_3814# a_14549_5336# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X544 a_22654_6022# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X545 a_1405_9065# a_984_9065# a_576_9144# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X546 a_3843_11350# a_3479_9828# a_2453_9061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X547 a_11283_13552# a_11283_13157# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X548 a_1402_7471# a_981_7471# a_573_7155# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X549 vdd d0 a_20138_2311# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X550 vdd d0 a_41813_8996# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X551 a_984_9833# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X552 a_8130_12756# a_9223_13418# a_9174_13608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X553 a_11282_2735# a_11282_2480# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X554 a_3521_11350# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X555 a_1405_9065# a_2245_9061# a_2453_9061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X556 vdd a_41810_5955# a_41602_5955# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X557 a_11691_13473# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X558 a_32956_11453# a_33577_11345# a_33785_11345# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X559 a_29803_12754# a_30056_12741# a_28356_11987# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X560 gnd a_6937_9009# a_6729_9009# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X561 a_11904_11347# a_11691_11347# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X562 a_33575_7463# a_33362_7463# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X563 a_11284_8488# a_11905_8380# a_12113_8380# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X564 a_14185_3814# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X565 a_29797_6923# a_30894_6729# a_30849_6742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X566 a_9176_5976# a_9429_5963# a_8128_5301# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X567 a_19881_3180# a_19885_2324# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X568 a_22868_3055# a_22655_3055# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X569 a_5254_4506# a_5618_7419# a_5573_7432# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X570 a_18838_12750# a_19931_13412# a_19886_13425# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X571 a_22248_12906# a_22248_12365# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X572 a_22656_11351# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X573 a_18834_12927# a_19091_12737# a_17391_11983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X574 vdd a_20140_8998# a_19932_8998# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X575 a_18836_5295# a_19089_5282# a_17385_6152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X576 a_18837_2328# a_19090_2315# a_17386_3185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X577 a_41554_2499# a_41811_2309# a_40506_2503# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X578 a_6635_4636# a_6727_3001# a_6678_3191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X579 a_23078_8384# a_23918_9059# a_24126_9059# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X580 a_22657_9831# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X581 gnd a_40763_2313# a_40555_2313# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X582 a_25192_5340# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X583 a_23075_7469# a_23915_7465# a_24123_7465# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X584 a_33783_5337# a_33362_5337# a_32955_4831# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X585 a_34831_7459# a_36070_6779# a_36227_5453# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X586 vdd a_19091_11290# a_18883_11290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X587 gnd a_20138_2311# a_19930_2311# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X588 a_575_11461# a_1196_11353# a_1404_11353# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X589 a_1403_2378# a_982_2378# a_574_2486# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X590 a_2243_4500# a_2030_4500# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X591 a_39065_9014# a_40557_9768# a_40508_9958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X592 a_11283_12105# a_11904_12026# a_12112_12026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X593 a_29799_12931# a_30056_12741# a_28356_11987# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X594 a_18835_8513# a_19932_8319# a_19887_8332# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X595 a_27026_4504# a_26605_4504# a_26927_4504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X596 a_32957_10839# a_32957_10583# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X597 a_23076_4502# a_22655_4502# a_22247_4186# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X598 a_25362_6785# a_25149_6785# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X599 a_33365_8378# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X600 gnd a_39275_10446# a_39067_10446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X601 a_23916_3051# a_23703_3051# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X602 a_573_5708# a_1194_6024# a_1402_6024# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X603 a_12740_9055# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X604 a_16281_7426# a_17394_10448# a_17345_10638# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X605 a_9173_3186# a_9430_2996# a_8129_2334# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X606 a_11281_5702# a_11281_5447# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X607 a_30847_12159# a_31104_11969# a_29803_11307# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X608 a_12111_4498# a_11690_4498# a_11282_4577# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X609 a_32957_8741# a_33578_9057# a_33786_9057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X610 a_2245_9061# a_2032_9061# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X611 a_40505_6917# a_41602_6723# a_41553_6913# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X612 a_18832_5472# a_19089_5282# a_17385_6152# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X613 a_32954_7542# a_33575_7463# a_33783_7463# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X614 a_18833_2505# a_19090_2315# a_17386_3185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X615 a_12113_8380# a_12953_9055# a_13161_9055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X616 a_12110_7465# a_12950_7461# a_13158_7461# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X617 vdd a_28608_2999# a_28400_2999# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X618 vdd a_40763_2313# a_40555_2313# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X619 a_2451_4500# a_3690_3820# a_3841_5342# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X620 vdd a_20138_2311# a_19930_2311# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X621 vdd a_41813_8996# a_41605_8996# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X622 a_22870_9063# a_22657_9063# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X623 a_29799_12931# a_30896_12737# a_30847_12927# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X624 a_12112_11347# a_11691_11347# a_11283_11455# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X625 a_11281_5447# a_11902_5339# a_12110_5339# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X626 gnd a_41810_5276# a_41602_5276# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X627 a_35860_9820# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X628 vdd a_39275_10446# a_39067_10446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X629 a_36222_5334# a_35858_3812# a_34832_4492# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X630 a_30850_2328# a_30846_2505# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X631 a_33362_7463# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X632 a_3519_5342# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X633 a_28357_9020# a_28610_9007# a_28310_10642# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X634 a_39061_9191# a_39318_9001# a_39018_10636# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X635 a_17385_6152# a_17642_5962# a_17347_4453# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X636 a_576_9400# a_1197_9833# a_1405_9833# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X637 a_22655_3055# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X638 a_40510_2326# a_41603_2988# a_41558_3001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X639 a_40505_6917# a_41602_6723# a_41557_6736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X640 a_11691_12026# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X641 a_40509_6740# a_40762_6727# a_39062_5973# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X642 a_1404_11353# a_2244_12028# a_2452_12028# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X643 a_33575_6016# a_33362_6016# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X644 a_11284_10190# a_11905_10506# a_12113_10506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X645 a_19884_6738# a_20137_6725# a_18832_6919# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X646 a_1195_3057# a_982_3057# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X647 a_32957_2379# a_33576_2370# a_33784_2370# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X648 a_3689_6787# a_3476_6787# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X649 a_12739_12022# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X650 a_30848_8513# a_30849_7421# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X651 a_22246_6357# a_22867_6790# a_23075_6790# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X652 a_9179_9785# a_9175_9962# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X653 gnd d1 a_8382_2321# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X654 a_36321_5334# a_35900_5334# a_36227_5453# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X655 a_22247_2739# a_22247_2484# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X656 a_3848_11469# a_3734_11350# a_3942_11350# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X657 a_33576_4496# a_33363_4496# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X658 a_2451_3053# a_2030_3053# a_1403_2378# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X659 vdd a_41810_5276# a_41602_5276# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X660 a_22869_12030# a_22656_12030# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X661 gnd a_9429_6731# a_9221_6731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X662 a_12111_2372# a_11690_2372# a_11284_2381# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X663 a_34834_9053# a_34413_9053# a_33786_8378# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X664 a_23703_3051# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X665 a_30848_10639# a_30852_9783# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X666 a_33785_13471# a_33364_13471# a_32956_13550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X667 a_983_12800# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X668 gnd a_20139_11965# a_19931_11965# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X669 a_34623_6012# a_34410_6012# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X670 a_1197_8386# a_984_8386# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X671 a_30851_11303# a_31104_11290# a_29799_11484# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X672 a_19881_3180# a_20138_2990# a_18837_2328# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X673 a_29801_5299# a_30054_5286# a_28350_6156# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X674 a_19880_6915# a_20137_6725# a_18832_6919# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X675 a_30846_4631# a_30850_3775# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X676 a_6684_9022# a_6937_9009# a_6637_10644# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X677 a_33578_9825# a_33365_9825# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X678 vdd d1 a_8382_2321# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X679 a_9173_4633# a_9177_3777# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X680 vdd a_9429_6731# a_9221_6731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X681 a_11692_10506# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X682 a_19887_9779# a_19883_9956# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X683 a_574_3136# a_1195_3057# a_1403_3057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X684 gnd d0 a_9431_12739# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X685 a_39064_11981# a_39317_11968# a_39022_10459# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X686 gnd d0 a_9429_5963# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X687 a_23077_13477# a_23917_13473# a_24125_13473# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X688 a_22248_12109# a_22248_11714# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X689 vdd a_41812_11963# a_41604_11963# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X690 a_17386_3185# a_18882_2315# a_18833_2505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X691 vdd d2 a_39315_5960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X692 a_32688_217# a_32579_217# a_21652_206# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X693 a_8127_8519# a_8384_8329# a_6680_9199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X694 a_33784_3049# a_33363_3049# a_32955_3128# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X695 a_29797_5476# a_30054_5286# a_28350_6156# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X696 a_9174_11482# a_9431_11292# a_8126_11486# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X697 a_9179_9017# a_9432_9004# a_8131_8342# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X698 a_36073_9820# a_35860_9820# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X699 a_13159_3047# a_12738_3047# a_12111_3051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X700 a_37389_8369# a_36968_8369# a_36321_5334# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X701 a_33362_6016# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X702 a_17391_11983# a_17644_11970# a_17349_10461# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X703 a_27242_7607# a_28357_4444# a_28308_4634# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X704 a_3476_6787# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X705 a_18837_3775# a_19930_4437# a_19885_4450# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X706 a_9176_7423# a_9429_7410# a_8128_6748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X707 a_22868_4502# a_22655_4502# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X708 a_33363_4496# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X709 a_11903_4498# a_11690_4498# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X710 a_2450_6020# a_3689_6787# a_3846_5461# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X711 a_2452_13475# a_2031_13475# a_1404_12800# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X712 a_573_7155# a_573_6900# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X713 a_9178_13431# a_11283_13552# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X714 a_17386_3185# a_18882_2315# a_18837_2328# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X715 a_37635_4498# a_37526_4498# a_32688_217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X716 vdd d1 a_30055_2319# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X717 a_33784_4496# a_34624_4492# a_34832_4492# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X718 vdd a_31105_10449# a_30897_10449# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X719 gnd d0 a_9432_9772# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X720 a_34834_9053# a_36073_9820# a_36224_11342# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X721 a_28308_4634# a_28400_2999# a_28351_3189# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X722 a_39016_4628# a_39108_2993# a_39063_3006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X723 a_575_12908# a_1196_12800# a_1404_12800# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X724 a_3841_5342# a_3477_3820# a_2451_3053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X725 a_1403_3825# a_982_3825# a_574_3933# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X726 a_29797_6923# a_30894_6729# a_30845_6919# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X727 a_41556_9186# a_41813_8996# a_40512_8334# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X728 gnd d0 a_31103_2994# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X729 a_21330_206# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X730 a_34410_6012# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X731 a_5254_4506# a_5618_7419# a_5569_7609# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X732 a_23704_13473# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X733 a_32956_12359# a_32956_12103# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X734 a_22248_11714# a_22248_11459# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X735 gnd d1 a_30056_11294# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X736 a_25365_9826# a_25152_9826# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X737 a_18838_12750# a_19091_12737# a_17391_11983# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X738 a_11284_10585# a_11284_10190# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X739 a_32955_4575# a_32955_4180# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X740 a_27242_7607# a_28357_4444# a_28312_4457# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X741 a_33365_9825# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X742 a_33364_12792# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X743 gnd d3 a_17600_4440# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X744 a_9172_7600# a_9429_7410# a_8128_6748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X745 a_33785_12024# a_33364_12024# a_32956_11708# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X746 a_18832_6919# a_19089_6729# a_17389_5975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X747 a_3940_5342# a_3519_5342# a_3841_5342# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X748 vdd d0 a_9432_9772# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X749 gnd d0 a_31105_8323# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X750 a_18835_8513# a_19932_8319# a_19883_8509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X751 vdd a_8382_3768# a_8174_3768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X752 vdd a_39315_5960# a_39107_5960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X753 a_17347_4453# a_17434_5962# a_17385_6152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X754 a_34624_3045# a_34411_3045# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X755 a_2450_6020# a_2029_6020# a_1402_6024# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X756 a_29802_2332# a_30895_2994# a_30850_3007# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X757 a_23075_5343# a_22654_5343# a_22247_4837# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X758 gnd a_41812_11284# a_41604_11284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X759 a_6678_3191# a_8174_2321# a_8125_2511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X760 a_12739_13469# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X761 a_12112_12794# a_11691_12794# a_11283_12902# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X762 a_41558_4448# a_41554_4625# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X763 a_17387_12160# a_18883_11290# a_18834_11480# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X764 a_12110_5339# a_11689_5339# a_11281_5447# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X765 gnd a_41810_6723# a_41602_6723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X766 a_23917_12026# a_23704_12026# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X767 a_9179_9017# a_9175_9194# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X768 a_22869_13477# a_22656_13477# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X769 a_1404_12032# a_983_12032# a_575_11716# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X770 vdd d3 a_17600_4440# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X771 a_33577_11345# a_33364_11345# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X772 gnd d1 a_40763_3760# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X773 a_11903_2372# a_11690_2372# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X774 a_6679_12166# a_8175_11296# a_8126_11486# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X775 a_19887_9779# a_20140_9766# a_18835_9960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X776 a_22655_4502# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X777 a_22249_8747# a_22870_9063# a_23078_9063# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X778 a_3691_12795# a_3478_12795# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X779 a_11689_7465# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X780 a_24126_10506# a_25365_9826# a_25516_11348# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X781 a_11690_4498# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X782 vdd d0 a_31105_8323# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X783 a_19887_10458# a_20140_10445# a_18839_9783# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X784 a_32955_3384# a_33576_3817# a_33784_3817# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X785 a_1195_4504# a_982_4504# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X786 vdd a_30055_2319# a_29847_2319# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X787 gnd a_9432_9772# a_9224_9772# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X788 a_25519_5459# a_25149_6785# a_24123_7465# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X789 vdd d2 a_28609_11974# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X790 vdd a_41812_11284# a_41604_11284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X791 a_6678_3191# a_8174_2321# a_8129_2334# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X792 a_14186_12789# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X793 gnd a_31103_2994# a_30895_2994# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X794 a_2451_4500# a_2030_4500# a_1403_3825# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X795 vdd a_41811_2988# a_41603_2988# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X796 a_33786_10504# a_33365_10504# a_32957_10583# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X797 vdd a_41810_6723# a_41602_6723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X798 a_8129_2334# a_9222_2996# a_9173_3186# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X799 a_1196_11353# a_983_11353# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X800 a_23077_12798# a_22656_12798# a_22248_12365# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X801 a_14648_5336# a_14227_5336# a_14554_5455# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X802 gnd d0 a_41810_5955# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X803 a_25152_9826# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X804 a_28355_3012# a_29847_3766# a_29798_3956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X805 vdd d1 a_40763_3760# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X806 a_15508_8371# a_15295_8371# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X807 a_19883_9956# a_20140_9766# a_18835_9960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X808 gnd a_28609_11974# a_28401_11974# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X809 a_35858_3812# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X810 gnd a_20139_13412# a_19931_13412# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X811 a_12113_9059# a_11692_9059# a_11284_8743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X812 a_19882_12923# a_19886_11978# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X813 a_22247_2484# a_22249_2385# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X814 a_29801_6746# a_30054_6733# a_28354_5979# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X815 a_6639_4459# a_6726_5968# a_6681_5981# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X816 a_19883_10635# a_20140_10445# a_18839_9783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X817 vdd a_9432_9772# a_9224_9772# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X818 a_22249_2385# a_22868_2376# a_23076_2376# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X819 a_24124_4498# a_23703_4498# a_23076_4502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X820 gnd a_31105_8323# a_30897_8323# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X821 a_23078_10510# a_23918_10506# a_24126_10506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X822 a_34411_3045# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X823 a_19880_6915# a_19884_5970# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X824 a_8127_8519# a_9224_8325# a_9175_8515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X825 a_1405_10512# a_984_10512# a_576_10591# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X826 gnd d2 a_28608_2999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X827 a_32579_217# a_32366_217# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X828 a_6679_12166# a_6936_11976# a_6641_10467# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X829 gnd d3 a_28567_10452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X830 a_35900_5334# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X831 a_574_4583# a_1195_4504# a_1403_4504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X832 a_28355_3012# a_29847_3766# a_29802_3779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X833 a_981_6792# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X834 gnd d0 a_9429_7410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X835 a_28314_10465# a_28401_11974# a_28356_11987# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X836 a_3846_5461# a_3476_6787# a_2450_7467# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X837 gnd d1 a_19090_3762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X838 gnd d0 a_41813_9764# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X839 a_11690_2372# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X840 vdd a_20139_13412# a_19931_13412# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X841 a_11015_219# a_15640_4500# a_15716_8371# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X842 a_33784_4496# a_33363_4496# a_32955_4575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X843 a_30847_12927# a_31104_12737# a_29799_12931# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X844 a_29797_6923# a_30054_6733# a_28354_5979# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X845 a_33364_12024# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X846 a_4932_4506# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X847 a_37181_8369# a_36968_8369# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X848 a_13159_4494# a_12738_4494# a_12111_4498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X849 a_3479_9828# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X850 a_9177_3009# a_9173_3186# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X851 a_14650_11344# a_15508_8371# a_15716_8371# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X852 vdd a_31105_8323# a_30897_8323# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X853 a_2453_10508# a_2032_10508# a_1405_9833# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X854 gnd d1 a_8383_11296# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X855 a_18839_9783# a_19092_9770# a_17392_9016# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X856 a_32955_2478# a_32957_2379# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X857 a_30849_7421# a_31102_7408# a_29801_6746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X858 a_8127_8519# a_9224_8325# a_9179_8338# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X859 gnd a_19090_2315# a_18882_2315# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X860 a_34833_12020# a_34412_12020# a_33785_12024# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X861 vdd d3 a_28567_10452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X862 a_11281_6097# a_11281_5702# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X863 a_8131_8342# a_8384_8329# a_6680_9199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X864 a_11689_6018# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X865 a_29804_8340# a_30897_9002# a_30848_9192# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X866 vdd d0 a_9429_7410# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X867 a_22248_12365# a_22869_12798# a_23077_12798# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X868 a_23705_10506# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X869 vdd d1 a_19090_3762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X870 a_12950_7461# a_12737_7461# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X871 vdd d0 a_41813_9764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X872 a_36323_11342# a_35902_11342# a_36224_11342# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X873 a_15295_8371# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X874 a_40511_11301# a_40764_11288# a_39060_12158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X875 a_18836_6742# a_19929_7404# a_19880_7594# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X876 a_34626_10500# a_34413_10500# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X877 gnd d0 a_31103_4441# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X878 a_18837_3775# a_19930_4437# a_19881_4627# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X879 a_3942_11350# a_3521_11350# a_3848_11469# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X880 a_23076_3055# a_22655_3055# a_22247_3134# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X881 a_22867_5343# a_22654_5343# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X882 a_25514_5340# a_25150_3818# a_24124_3051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X883 vdd a_9430_2996# a_9222_2996# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X884 gnd d1 a_30056_12741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X885 a_11902_5339# a_11689_5339# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X886 a_11282_4182# a_11903_4498# a_12111_4498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X887 a_39062_5973# a_39315_5960# a_39020_4451# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X888 a_18835_9960# a_19092_9770# a_17392_9016# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X889 a_36968_8369# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X890 a_30846_3184# a_30850_2328# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X891 vdd a_19090_2315# a_18882_2315# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X892 a_9177_3777# a_9430_3764# a_8125_3958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X893 vdd d2 a_17643_2995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X894 gnd d1 a_30055_2319# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X895 a_12737_6014# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X896 vdd a_40765_9768# a_40557_9768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X897 a_1404_13479# a_983_13479# a_575_13558# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X898 gnd a_31105_10449# a_30897_10449# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X899 a_39061_9191# a_40557_8321# a_40508_8511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X900 a_9173_3186# a_9177_2330# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X901 gnd d0 a_41813_10443# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X902 a_41556_8507# a_41557_7415# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X903 a_26927_4504# a_26818_4504# a_27026_4504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X904 a_11284_9935# a_11905_9827# a_12113_9827# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X905 a_33784_2370# a_33363_2370# a_32957_2379# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X906 a_23078_8384# a_22657_8384# a_22249_8492# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X907 gnd a_41813_9764# a_41605_9764# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X908 gnd a_41812_12731# a_41604_12731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X909 vdd d0 a_31103_4441# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X910 a_11283_12902# a_11904_12794# a_12112_12794# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X911 a_23077_12030# a_22656_12030# a_22248_12109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X912 a_30848_9192# a_31105_9002# a_29804_8340# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X913 gnd a_28610_9007# a_28402_9007# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X914 a_22656_12798# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X915 a_12110_6786# a_11689_6786# a_11281_6894# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X916 vdd d1 a_30056_12741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X917 a_18836_6742# a_19089_6729# a_17389_5975# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X918 a_41553_6913# a_41557_5968# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X919 a_9173_3954# a_9430_3764# a_8125_3958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X920 a_33577_12792# a_33364_12792# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X921 a_30850_2328# a_31103_2315# a_29798_2509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X922 a_15640_4500# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X923 a_6683_11989# a_8175_12743# a_8126_12933# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X924 a_14187_9822# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X925 gnd a_8382_3768# a_8174_3768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X926 a_17347_4453# a_17600_4440# a_16277_7603# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X927 a_39061_9191# a_40557_8321# a_40512_8334# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X928 vdd d0 a_31104_11969# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X929 vdd d4 a_27499_7417# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X930 vdd d0 a_41813_10443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X931 a_41554_4625# a_41558_3769# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X932 a_36222_5334# a_36113_5334# a_36321_5334# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X933 vdd d2 a_28610_9007# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X934 a_11905_9059# a_11692_9059# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X935 a_573_5708# a_573_5453# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X936 a_40512_8334# a_41605_8996# a_41556_9186# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X937 a_1403_3057# a_2243_3053# a_2451_3053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X938 vdd a_41813_9764# a_41605_9764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X939 vdd a_41812_12731# a_41604_12731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X940 gnd a_9431_11971# a_9223_11971# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X941 a_23916_4498# a_23703_4498# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X942 a_11015_219# a_10906_219# a_11114_219# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X943 a_981_6024# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X944 a_34625_13467# a_34412_13467# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X945 a_17391_11983# a_18883_12737# a_18838_12750# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X946 a_11282_2480# a_11903_2372# a_12111_2372# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X947 gnd a_31103_4441# a_30895_4441# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X948 a_22654_5343# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X949 a_6639_4459# a_6892_4446# a_5569_7609# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X950 a_1405_8386# a_984_8386# a_573_7806# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X951 a_40512_9781# a_41605_10443# a_41556_10633# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X952 a_8129_3781# a_9222_4443# a_9173_4633# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X953 a_19882_13602# a_19886_12746# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X954 a_983_11353# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X955 a_12950_6014# a_12737_6014# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X956 a_30846_2505# a_31103_2315# a_29798_2509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X957 a_4800_8377# a_4587_8377# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X958 a_6683_11989# a_8175_12743# a_8130_12756# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X959 a_1194_5345# a_981_5345# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X960 a_11691_12794# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X961 a_17343_4630# a_17600_4440# a_16277_7603# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X962 a_29799_11484# a_30896_11290# a_30851_11303# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X963 gnd a_30055_2319# a_29847_2319# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X964 a_19880_7594# a_19884_6738# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X965 a_40510_3773# a_40763_3760# a_39063_3006# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X966 a_33578_8378# a_33365_8378# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X967 a_12951_4494# a_12738_4494# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X968 a_15853_4500# a_15640_4500# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X969 a_22246_6101# a_22246_5706# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X970 gnd d0 a_20137_5957# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X971 a_33575_6784# a_33362_6784# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X972 a_32954_7798# a_32954_7542# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X973 a_8130_11309# a_9223_11971# a_9178_11984# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X974 a_22247_3390# a_22868_3823# a_23076_3823# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X975 a_34833_12020# a_36072_12787# a_36229_11461# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X976 a_2244_13475# a_2031_13475# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X977 a_13159_3047# a_14398_3814# a_14549_5336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X978 a_14399_12789# a_14186_12789# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X979 a_17392_9016# a_18884_9770# a_18835_9960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X980 vdd d0 a_31102_5961# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X981 a_3843_11350# a_3479_9828# a_2453_10508# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X982 vdd a_31103_4441# a_30895_4441# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X983 a_6635_4636# a_6892_4446# a_5569_7609# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X984 vdd a_17645_9003# a_17437_9003# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X985 a_40512_9781# a_41605_10443# a_41560_10456# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X986 a_40506_2503# a_41603_2309# a_41554_2499# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X987 a_1402_7471# a_981_7471# a_573_7550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X988 a_8129_3781# a_9222_4443# a_9177_4456# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X989 a_25407_11348# a_25194_11348# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X990 a_984_9833# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X991 vdd d2 a_6937_9009# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X992 a_12738_3047# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X993 vdd d0 a_41810_7402# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X994 a_22246_7548# a_22867_7469# a_23075_7469# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X995 a_1405_8386# a_2245_9061# a_2453_9061# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X996 a_574_3392# a_574_3136# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X997 a_32957_10839# a_33577_11345# a_33785_11345# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X998 a_41557_5968# a_41810_5955# a_40509_5293# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X999 gnd a_8383_11296# a_8175_11296# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1000 a_25519_5459# a_25405_5340# a_25613_5340# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1001 a_11904_11347# a_11691_11347# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1002 a_40506_3950# a_40763_3760# a_39063_3006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1003 a_12113_10506# a_12953_10502# a_13161_10502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1004 a_19881_3948# a_20138_3758# a_18833_3952# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1005 a_6641_10467# a_6894_10454# a_5573_7432# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1006 gnd d2 a_17645_9003# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1007 a_22868_3055# a_22655_3055# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1008 a_2452_12028# a_3691_12795# a_3848_11469# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1009 gnd d0 a_31104_11290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1010 a_573_5453# a_1194_5345# a_1402_5345# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1011 a_11692_9059# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1012 gnd d1 a_8383_12743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1013 a_12111_3819# a_11690_3819# a_11282_3386# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1014 a_32957_8486# a_33578_8378# a_33786_8378# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1015 a_1197_9065# a_984_9065# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1016 a_17392_9016# a_18884_9770# a_18839_9783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1017 a_23703_4498# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1018 a_11284_8488# a_11281_7800# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1019 a_30852_9783# a_30848_9960# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1020 a_28355_3012# a_28608_2999# a_28308_4634# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1021 a_23075_6790# a_23915_7465# a_24123_7465# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1022 a_33783_5337# a_33362_5337# a_32954_5445# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1023 a_34831_6012# a_36070_6779# a_36227_5453# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1024 a_576_10847# a_1196_11353# a_1404_11353# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1025 a_30851_12750# a_31104_12737# a_29799_12931# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1026 a_35859_12787# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1027 gnd d2 a_39317_11968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1028 a_22870_8384# a_22657_8384# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1029 a_11283_11710# a_11904_12026# a_12112_12026# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1030 a_27026_4504# a_26605_4504# a_26681_8375# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1031 a_40511_12748# a_40764_12735# a_39064_11981# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1032 a_41560_9777# a_41813_9764# a_40508_9958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1033 a_23076_4502# a_22655_4502# a_22247_4581# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1034 a_33365_8378# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1035 a_6637_10644# a_6894_10454# a_5573_7432# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1036 gnd a_20137_5957# a_19929_5957# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1037 a_12740_9055# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1038 a_33362_6784# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1039 vdd d0 a_9431_11292# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1040 a_11902_6786# a_11689_6786# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1041 a_2245_9061# a_2032_9061# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1042 vdd d1 a_8383_12743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1043 a_982_3057# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1044 a_32954_7147# a_33575_7463# a_33783_7463# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1045 a_8126_11486# a_9223_11292# a_9174_11482# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1046 a_24126_9059# a_23705_9059# a_23078_8384# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1047 a_12110_6786# a_12950_7461# a_13158_7461# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1048 vdd a_31102_5961# a_30894_5961# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1049 a_22246_7153# a_22246_6898# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1050 a_3478_12795# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1051 a_8128_5301# a_9221_5963# a_9176_5976# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1052 gnd d2 a_6936_11976# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1053 gnd d0 a_31102_5282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1054 a_1402_5345# a_2242_6020# a_2450_6020# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1055 a_26927_4504# a_27291_7417# a_27246_7430# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1056 a_1195_2378# a_982_2378# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1057 vdd a_6937_9009# a_6729_9009# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1058 a_11282_4833# a_11902_5339# a_12110_5339# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1059 a_41553_7592# a_41557_6736# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1060 a_40507_12925# a_40764_12735# a_39064_11981# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1061 a_29798_3956# a_30895_3762# a_30846_3952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1062 a_30845_5472# a_30850_4454# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1063 a_41556_9954# a_41813_9764# a_40508_9958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1064 a_1402_6024# a_981_6024# a_573_5708# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1065 a_19886_13425# a_22248_13556# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1066 a_3519_5342# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1067 gnd a_40765_9768# a_40557_9768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1068 a_12112_13473# a_12952_13469# a_13160_13469# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1069 a_33786_9057# a_33365_9057# a_32957_8741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1070 a_9179_10464# a_9432_10451# a_8131_9789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1071 a_11691_12026# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1072 gnd a_20140_9766# a_19932_9766# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1073 a_22655_3055# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1074 a_41555_12153# a_41812_11963# a_40511_11301# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1075 a_19883_9956# a_19887_9011# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1076 a_33785_12792# a_33364_12792# a_32956_12359# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1077 a_33575_6016# a_33362_6016# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1078 vdd d2 a_28607_5966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1079 a_12739_12022# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1080 a_22249_10589# a_22249_10194# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1081 a_3690_3820# a_3477_3820# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1082 a_17386_3185# a_17643_2995# a_17343_4630# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1083 vdd d0 a_31102_5282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1084 a_24123_6018# a_25362_6785# a_25519_5459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1085 a_5008_8377# a_5145_4506# a_5353_4506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1086 a_41560_8330# a_41556_8507# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1087 a_18834_11480# a_19091_11290# a_17387_12160# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1088 a_32954_7147# a_32954_6892# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1089 a_2451_3053# a_2030_3053# a_1403_3057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1090 a_1403_4504# a_2243_4500# a_2451_4500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1091 a_29798_3956# a_30895_3762# a_30850_3775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1092 a_22657_8384# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1093 a_33786_10504# a_34626_10500# a_34834_10500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1094 a_12111_2372# a_11690_2372# a_11282_2480# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1095 a_34834_9053# a_34413_9053# a_33786_9057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1096 a_6641_10467# a_6728_11976# a_6679_12166# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1097 a_23075_6022# a_23915_6018# a_24123_6018# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1098 a_9175_10641# a_9432_10451# a_8131_9789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1099 a_1405_9833# a_984_9833# a_576_9400# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1100 vdd a_20140_9766# a_19932_9766# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1101 gnd d4 a_27499_7417# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1102 a_575_12367# a_575_12111# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1103 a_29799_11484# a_30056_11294# a_28352_12164# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1104 gnd d0 a_20140_8998# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1105 a_12112_13473# a_11691_13473# a_11283_13157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1106 a_41558_3001# a_41554_3178# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1107 a_1194_6792# a_981_6792# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1108 a_23076_4502# a_23916_4498# a_24124_4498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1109 a_573_5453# a_574_4839# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1110 a_2245_10508# a_2032_10508# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1111 a_22249_8492# a_22246_7804# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1112 a_33578_9825# a_33365_9825# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1113 a_36113_5334# a_35900_5334# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1114 gnd a_31102_5282# a_30894_5282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1115 a_17391_11983# a_18883_12737# a_18834_12927# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1116 a_8124_5478# a_9221_5284# a_9172_5474# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1117 a_32954_6095# a_33575_6016# a_33783_6016# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1118 a_23077_11351# a_22656_11351# a_22249_10845# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1119 a_32956_12103# a_32956_11708# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1120 gnd d0 a_20140_10445# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1121 a_28353_9197# a_28610_9007# a_28310_10642# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1122 vdd a_9431_13418# a_9223_13418# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1123 a_574_2741# a_1195_3057# a_1403_3057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1124 gnd d3 a_28565_4444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1125 a_12110_6018# a_12950_6014# a_13158_6014# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1126 a_14556_11463# a_14186_12789# a_13160_12022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1127 a_19883_8509# a_20140_8319# a_18835_8513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1128 a_23077_12798# a_23917_13473# a_24125_13473# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1129 a_11903_3819# a_11690_3819# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1130 a_3942_11350# a_4800_8377# a_5008_8377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1131 a_40506_3950# a_41603_3756# a_41554_3946# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1132 a_32955_4575# a_33576_4496# a_33784_4496# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1133 a_5145_4506# a_4932_4506# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1134 a_19884_5970# a_19880_6147# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1135 gnd d1 a_8384_9776# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1136 a_12111_4498# a_12951_4494# a_13159_4494# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1137 a_15962_4500# a_15853_4500# a_11015_219# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1138 a_32956_12359# a_33577_12792# a_33785_12792# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1139 a_37950_7601# a_39065_4438# a_39020_4451# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1140 a_30852_9015# a_30848_9192# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1141 a_41559_11297# a_41812_11284# a_40507_11478# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1142 a_37389_8369# a_36968_8369# a_36323_11342# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1143 gnd a_8383_12743# a_8175_12743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1144 a_33362_6016# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1145 a_11904_12794# a_11691_12794# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1146 vdd d2 a_39316_2993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1147 a_22249_10589# a_22870_10510# a_23078_10510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1148 vdd d0 a_20137_7404# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1149 vdd a_31102_5282# a_30894_5282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1150 a_573_7806# a_1197_8386# a_1405_8386# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1151 gnd a_41811_2309# a_41603_2309# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1152 a_22868_4502# a_22655_4502# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1153 a_25405_5340# a_25192_5340# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1154 a_8124_5478# a_9221_5284# a_9176_5297# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1155 vdd d0 a_20140_10445# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1156 a_41554_3178# a_41558_2322# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1157 a_14397_6781# a_14184_6781# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1158 a_1196_12800# a_983_12800# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1159 a_28351_3189# a_29847_2319# a_29802_2332# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1160 vdd d3 a_28565_4444# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1161 a_8128_5301# a_8381_5288# a_6677_6158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1162 a_32957_9933# a_33578_9825# a_33786_9825# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1163 a_2452_13475# a_2031_13475# a_1404_13479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1164 a_40506_3950# a_41603_3756# a_41558_3769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1165 a_33785_13471# a_34625_13467# a_34833_13467# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1166 a_18838_11303# a_19931_11965# a_19886_11978# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1167 a_23918_9059# a_23705_9059# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1168 vdd d3 a_17602_10448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1169 vdd d1 a_8384_9776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1170 a_33783_6784# a_33362_6784# a_32954_6892# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1171 a_33576_3049# a_33363_3049# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1172 a_576_9941# a_576_9400# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1173 a_19885_3771# a_20138_3758# a_18833_3952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1174 a_22870_9831# a_22657_9831# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1175 a_6680_9199# a_6937_9009# a_6637_10644# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1176 a_41555_11474# a_41812_11284# a_40507_11478# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1177 a_24124_4498# a_25363_3818# a_25514_5340# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1178 a_41553_7592# a_41810_7402# a_40509_6740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1179 a_23704_13473# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1180 vdd a_8383_12743# a_8175_12743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1181 a_30849_5974# a_31102_5961# a_29801_5299# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1182 a_10906_219# a_10693_219# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1183 a_33365_9825# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1184 gnd d1 a_30057_9774# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1185 vdd d0 a_31104_12737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1186 gnd a_9430_3764# a_9222_3764# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1187 a_22869_12798# a_22656_12798# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1188 a_33785_12024# a_33364_12024# a_32956_12103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1189 a_982_4504# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1190 a_17392_9016# a_17645_9003# a_17345_10638# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1191 vdd d0 a_41813_8317# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1192 gnd a_28565_4444# a_28357_4444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1193 a_39058_6150# a_40554_5280# a_40505_5470# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1194 a_3940_5342# a_3519_5342# a_3846_5461# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1195 a_22249_8492# a_22870_8384# a_23078_8384# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1196 a_13160_12022# a_14399_12789# a_14556_11463# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1197 a_22657_10510# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1198 a_11689_6786# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1199 a_11690_3819# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1200 a_34624_3045# a_34411_3045# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1201 a_36070_6779# a_35857_6779# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1202 a_11281_7800# a_11905_8380# a_12113_8380# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1203 gnd a_41555_13600# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1204 a_25521_11467# a_25407_11348# a_25615_11348# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1205 a_25149_6785# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1206 a_26681_8375# a_26260_8375# a_25613_5340# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1207 a_1195_3825# a_982_3825# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1208 a_23075_5343# a_22654_5343# a_22246_5451# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1209 a_11114_219# a_21543_206# vout gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1210 a_30846_3952# a_30850_3007# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1211 a_25151_12793# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1212 a_11281_6353# a_11902_6786# a_12110_6786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1213 a_23077_12030# a_23917_12026# a_24125_12026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1214 vdd a_39316_2993# a_39108_2993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1215 vdd d1 a_30057_9774# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1216 a_22248_13556# a_22869_13477# a_23077_13477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1217 a_1404_12032# a_983_12032# a_575_12111# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1218 vdd a_20137_7404# a_19929_7404# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1219 a_30852_9783# a_31105_9770# a_29800_9964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1220 vdd a_9430_3764# a_9222_3764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1221 a_11282_3386# a_11282_3130# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1222 a_11903_2372# a_11690_2372# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1223 a_19881_2501# a_11284_2381# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1224 a_22655_4502# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1225 a_25192_5340# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1226 gnd d0 a_9430_2996# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1227 gnd a_17600_4440# a_17392_4440# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1228 a_26927_4504# a_27291_7417# a_27242_7607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1229 a_14184_6781# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1230 a_24126_9059# a_25365_9826# a_25516_11348# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1231 vdd a_28565_4444# a_28357_4444# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1232 a_39058_6150# a_40554_5280# a_40509_5293# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1233 a_8126_12933# a_9223_12739# a_9178_12752# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1234 a_28308_4634# a_28400_2999# a_28355_3012# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1235 a_14554_5455# a_14440_5336# a_14648_5336# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1236 a_18837_2328# a_19930_2990# a_19885_3003# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1237 a_23705_9059# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1238 vdd d0 a_31102_6729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1239 a_18834_11480# a_19931_11286# a_19882_11476# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1240 a_33363_3049# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1241 a_2031_13475# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1242 a_2452_12028# a_2031_12028# a_1404_11353# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1243 a_12113_10506# a_11692_10506# a_11284_10190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1244 a_33784_3049# a_34624_3045# a_34832_3045# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1245 a_9173_2507# a_9430_2317# a_8125_2511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1246 gnd a_17642_5962# a_17434_5962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1247 a_2242_7467# a_2029_7467# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1248 a_30848_9960# a_31105_9770# a_29800_9964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1249 a_32957_10188# a_32957_9933# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1250 gnd d0 a_9432_8325# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1251 gnd a_8382_2321# a_8174_2321# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1252 a_5008_8377# a_4587_8377# a_3940_5342# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1253 gnd a_30057_9774# a_29849_9774# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1254 a_15962_4500# a_16326_7413# a_16277_7603# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1255 a_23078_9063# a_22657_9063# a_22249_8747# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1256 a_2451_3053# a_3690_3820# a_3841_5342# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1257 vdd a_17600_4440# a_17392_4440# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1258 gnd d2 a_39318_9001# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1259 a_6684_9022# a_8176_9776# a_8127_9966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1260 a_574_3933# a_574_3392# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1261 a_23704_12026# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1262 a_12113_9059# a_11692_9059# a_11284_9138# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1263 vdd a_41813_8317# a_41605_8317# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1264 a_22656_13477# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1265 a_33784_3817# a_33363_3817# a_32955_3384# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1266 a_12110_7465# a_11689_7465# a_11281_7149# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1267 a_9174_12929# a_9178_11984# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1268 a_22249_10845# a_22249_10589# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1269 a_33364_11345# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1270 a_23078_9831# a_23918_10506# a_24126_10506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1271 a_28350_6156# a_28607_5966# a_28312_4457# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1272 a_39060_12158# a_39317_11968# a_39022_10459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1273 a_34411_3045# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1274 a_22246_5706# a_22246_5451# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1275 a_34625_12020# a_34412_12020# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1276 a_18834_11480# a_19931_11286# a_19886_11299# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1277 a_33577_13471# a_33364_13471# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1278 a_8124_6925# a_9221_6731# a_9172_6921# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1279 a_6635_4636# a_6727_3001# a_6682_3014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1280 a_574_4188# a_1195_4504# a_1403_4504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1281 a_19885_4450# a_19881_4627# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1282 vdd d0 a_9432_8325# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1283 a_41560_9777# a_41556_9954# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1284 vdd a_8382_2321# a_8174_2321# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1285 gnd a_31104_11969# a_30896_11969# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1286 vdd a_30057_9774# a_29849_9774# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1287 a_15962_4500# a_16326_7413# a_16281_7426# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1288 a_3734_11350# a_3521_11350# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1289 a_6684_9022# a_8176_9776# a_8131_9789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1290 a_11690_2372# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1291 gnd d0 a_41812_11963# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1292 a_3843_11350# a_3734_11350# a_3942_11350# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1293 a_17343_4630# a_17435_2995# a_17386_3185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1294 a_41559_12744# a_41812_12731# a_40507_12925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1295 a_23076_2376# a_22655_2376# a_22249_2385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1296 a_14648_5336# a_15508_8371# a_15716_8371# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1297 a_22869_12030# a_22656_12030# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1298 a_14229_11344# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1299 gnd a_9431_13418# a_9223_13418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1300 a_2453_10508# a_2032_10508# a_1405_10512# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1301 gnd d0 a_20138_2990# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1302 gnd d1 a_40763_2313# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1303 vdd a_31102_6729# a_30894_6729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1304 a_11282_3927# a_11903_3819# a_12111_3819# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1305 a_19887_8332# a_20140_8319# a_18835_8513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1306 gnd a_41811_3756# a_41603_3756# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1307 a_8124_6925# a_9221_6731# a_9176_6744# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1308 a_573_6900# a_573_6359# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1309 a_34831_7459# a_34410_7459# a_33783_6784# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1310 a_11689_6018# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1311 a_22246_6101# a_22867_6022# a_23075_6022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1312 a_983_12800# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1313 a_8128_6748# a_8381_6735# a_6681_5981# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1314 a_23705_10506# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1315 gnd a_9432_8325# a_9224_8325# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1316 a_36323_11342# a_35902_11342# a_36229_11461# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1317 a_37950_7601# a_39065_4438# a_39016_4628# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1318 a_19886_13425# a_19882_13602# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1319 a_32956_13550# a_32956_13155# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1320 a_22247_3390# a_22247_3134# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1321 a_41559_11297# a_41555_11474# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1322 gnd a_39318_9001# a_39110_9001# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1323 a_22867_5343# a_22654_5343# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1324 a_41555_12921# a_41812_12731# a_40507_12925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1325 a_25514_5340# a_25150_3818# a_24124_4498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1326 a_19884_7417# a_19880_7594# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1327 a_28351_3189# a_29847_2319# a_29798_2509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1328 vdd d2 a_28608_2999# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1329 vdd d1 a_40763_2313# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1330 a_36968_8369# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1331 vdd a_41811_3756# a_41603_3756# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1332 a_40511_11301# a_41604_11963# a_41555_12153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1333 gnd d0 a_41811_2988# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1334 gnd d3 a_17602_10448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1335 a_8124_6925# a_8381_6735# a_6681_5981# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1336 a_9172_6153# a_9429_5963# a_8128_5301# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1337 a_27242_7607# a_27499_7417# a_26927_4504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1338 a_576_8749# a_576_8494# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1339 a_22249_9939# a_22870_9831# a_23078_9831# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1340 a_14227_5336# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1341 a_36073_9820# a_35860_9820# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1342 vdd a_9432_8325# a_9224_8325# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1343 a_13161_10502# a_14400_9822# a_14551_11344# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1344 a_11284_9394# a_11905_9827# a_12113_9827# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1345 a_34624_4492# a_34411_4492# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1346 a_29802_3779# a_30055_3766# a_28355_3012# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1347 gnd d0 a_31104_12737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1348 a_14554_5455# a_14184_6781# a_13158_7461# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1349 a_30845_7598# a_31102_7408# a_29801_6746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1350 a_981_5345# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1351 a_29804_9787# a_30897_10449# a_30852_10462# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1352 gnd a_20138_2990# a_19930_2990# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1353 gnd d1 a_19090_2315# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1354 gnd d0 a_41813_8317# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1355 a_14187_9822# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1356 a_30847_11480# a_31104_11290# a_29799_11484# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1357 gnd d0 a_9430_4443# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1358 a_575_12367# a_1196_12800# a_1404_12800# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1359 a_2030_3053# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1360 a_3841_5342# a_3477_3820# a_2451_4500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1361 a_14556_11463# a_14442_11344# a_14650_11344# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1362 a_2032_10508# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1363 a_39062_5973# a_40554_6727# a_40509_6740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1364 a_11283_13157# a_11283_12902# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1365 a_40507_11478# a_40764_11288# a_39060_12158# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1366 a_11905_9059# a_11692_9059# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1367 a_574_3136# a_574_2741# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1368 a_1403_2378# a_2243_3053# a_2451_3053# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1369 a_41556_8507# a_41813_8317# a_40508_8511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1370 a_18839_8336# a_19092_8323# a_17388_9193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1371 a_37954_7424# a_38207_7411# a_37635_4498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1372 a_11902_7465# a_11689_7465# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1373 a_29798_3956# a_30055_3766# a_28355_3012# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1374 a_40509_6740# a_41602_7402# a_41553_7592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1375 a_3848_11469# a_3478_12795# a_2452_13475# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1376 gnd a_40765_8321# a_40557_8321# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1377 a_18834_12927# a_19931_12733# a_19882_12923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1378 a_12112_12026# a_12952_12022# a_13160_12022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1379 a_34625_13467# a_34412_13467# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1380 a_11284_2381# a_11903_2372# a_12111_2372# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1381 a_22654_5343# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1382 a_25364_12793# a_25151_12793# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1383 vdd d1 a_19090_2315# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1384 a_1402_6792# a_981_6792# a_573_6359# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1385 a_9174_13608# a_9178_12752# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1386 a_12950_6014# a_12737_6014# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1387 a_8126_12933# a_9223_12739# a_9174_12929# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1388 vout a_21330_206# a_21652_206# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1389 a_19885_2324# a_19881_2501# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1390 a_4800_8377# a_4587_8377# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1391 a_18836_5295# a_19929_5957# a_19880_6147# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1392 vdd d0 a_9430_4443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1393 gnd d0 a_9432_10451# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1394 gnd d0 a_31102_6729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1395 a_9175_9194# a_9432_9004# a_8131_8342# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1396 a_33578_10504# a_33365_10504# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1397 a_22248_12365# a_22248_12109# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1398 gnd a_6894_10454# a_6686_10454# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1399 a_18835_8513# a_19092_8323# a_17388_9193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1400 a_37950_7601# a_38207_7411# a_37635_4498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1401 a_9176_5297# a_9429_5284# a_8124_5478# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1402 a_9177_2330# a_9430_2317# a_8125_2511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1403 a_22868_2376# a_22655_2376# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1404 a_2244_13475# a_2031_13475# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1405 a_34411_4492# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1406 vdd a_40765_8321# a_40557_8321# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1407 vdd a_28610_9007# a_28402_9007# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1408 a_18834_12927# a_19931_12733# a_19886_12746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1409 a_36072_12787# a_35859_12787# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1410 vdd a_20140_8319# a_19932_8319# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1411 a_39063_3006# a_39316_2993# a_39016_4628# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1412 a_9179_10464# a_9175_10641# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1413 a_41557_7415# a_41553_7592# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1414 a_19884_7417# a_20137_7404# a_18836_6742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1415 a_25407_11348# a_25194_11348# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1416 a_12738_3047# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1417 a_22246_7153# a_22867_7469# a_23075_7469# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1418 a_23076_3055# a_23916_3051# a_24124_3051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1419 vdd a_17602_10448# a_17394_10448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1420 gnd a_31104_13416# a_30896_13416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1421 gnd a_41813_8317# a_41605_8317# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1422 a_37526_4498# a_37313_4498# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1423 a_1197_10512# a_984_10512# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1424 vdd d0 a_9432_10451# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1425 vdd d0 a_31103_2994# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1426 a_30847_12927# a_30851_11982# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1427 a_11283_11455# a_11904_11347# a_12112_11347# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1428 a_19886_11299# a_19882_11476# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1429 gnd d0 a_41812_13410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1430 vdd d1 a_30056_11294# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1431 a_12113_9827# a_12953_10502# a_13161_10502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1432 a_22657_9063# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1433 a_9178_12752# a_9174_12929# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1434 vdd a_6894_10454# a_6686_10454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1435 a_2451_4500# a_2030_4500# a_1403_4504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1436 a_23076_3823# a_22655_3823# a_22247_3390# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1437 a_9172_5474# a_9429_5284# a_8124_5478# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1438 vdd a_20139_11965# a_19931_11965# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1439 a_574_4839# a_1194_5345# a_1402_5345# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1440 a_11692_9059# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1441 a_14549_5336# a_14185_3814# a_13159_3047# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1442 gnd a_8381_5288# a_8173_5288# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1443 a_12111_3819# a_11690_3819# a_11282_3927# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1444 a_32954_7798# a_33578_8378# a_33786_8378# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1445 a_1197_9065# a_984_9065# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1446 a_3692_9828# a_3479_9828# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1447 gnd d2 a_6934_5968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1448 a_32954_6892# a_33575_6784# a_33783_6784# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1449 a_1194_7471# a_981_7471# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1450 a_9178_11984# a_9431_11971# a_8130_11309# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1451 a_2453_9061# a_2032_9061# a_1405_8386# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1452 vdd a_31104_13416# a_30896_13416# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1453 a_12113_8380# a_11692_8380# a_11281_7800# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1454 vdd d0 a_9429_5963# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1455 a_17387_12160# a_18883_11290# a_18838_11303# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1456 vdd d0 a_41812_13410# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1457 gnd a_31102_6729# a_30894_6729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1458 a_21652_206# a_32366_217# a_32688_217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1459 a_32366_217# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1460 vdd d0 a_20138_4437# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1461 a_32954_5445# a_32955_4831# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1462 a_982_3057# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1463 a_6679_12166# a_8175_11296# a_8130_11309# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1464 a_40506_2503# a_41603_2309# a_41558_2322# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1465 a_33785_12024# a_34625_12020# a_34833_12020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1466 a_11691_11347# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1467 a_22655_2376# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1468 a_24126_9059# a_23705_9059# a_23078_9063# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1469 a_36229_11461# a_35859_12787# a_34833_13467# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1470 a_17387_12160# a_17644_11970# a_17349_10461# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1471 a_32956_13550# a_33577_13471# a_33785_13471# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1472 a_40510_2326# a_40763_2313# a_39059_3183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1473 vdd d1 a_8384_8329# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1474 a_40511_12748# a_41604_13410# a_41555_13600# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1475 a_24123_7465# a_23702_7465# a_23075_6790# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1476 a_12951_3047# a_12738_3047# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1477 gnd d0 a_41811_4435# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1478 a_11904_13473# a_11691_13473# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1479 a_33575_5337# a_33362_5337# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1480 a_36227_5453# a_35857_6779# a_34831_6012# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1481 a_19885_2324# a_20138_2311# a_18833_2505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1482 a_1195_2378# a_982_2378# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1483 a_25615_11348# a_26473_8375# a_26681_8375# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1484 a_576_9144# a_1197_9065# a_1405_9065# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1485 a_26818_4504# a_26605_4504# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1486 a_30851_13429# a_32956_13550# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1487 a_2244_12028# a_2031_12028# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1488 a_37313_4498# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1489 a_17388_9193# a_18884_8323# a_18835_8513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1490 a_1196_13479# a_983_13479# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1491 vdd a_31103_2994# a_30895_2994# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1492 a_1402_6024# a_981_6024# a_573_6103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1493 a_22869_11351# a_22656_11351# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1494 a_8129_2334# a_9222_2996# a_9177_3009# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1495 a_984_8386# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1496 a_12112_12794# a_12952_13469# a_13160_13469# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1497 a_33786_9057# a_33365_9057# a_32957_9136# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1498 gnd d0 a_20139_11965# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1499 a_13161_10502# a_12740_10502# a_12113_9827# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1500 gnd d1 a_19091_11290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1501 a_33783_7463# a_33362_7463# a_32954_7147# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1502 a_27246_7430# a_27499_7417# a_26927_4504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1503 a_576_8494# a_573_7806# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1504 a_21543_206# a_21330_206# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1505 a_32957_10583# a_32957_10188# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1506 a_29801_6746# a_30894_7408# a_30845_7598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1507 a_13158_7461# a_12737_7461# a_12110_6786# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1508 a_40511_12748# a_41604_13410# gnd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1509 gnd a_20139_11286# a_19931_11286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1510 a_28351_3189# a_28608_2999# a_28308_4634# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1511 a_40506_2503# a_40763_2313# a_39059_3183# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1512 gnd a_6934_5968# a_6726_5968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1513 vdd d0 a_41811_4435# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1514 a_19881_2501# a_20138_2311# a_18833_2505# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1515 a_2030_4500# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1516 a_34626_10500# a_34413_10500# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1517 a_5254_4506# a_5145_4506# a_5353_4506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1518 a_41558_3001# a_41811_2988# a_40510_2326# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1519 a_11282_4182# a_11282_3927# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1520 a_11281_6894# a_11281_6353# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1521 a_29804_9787# a_30897_10449# a_30848_10639# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1522 vdd d1 a_30057_8327# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1523 a_17388_9193# a_18884_8323# a_18839_8336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1524 a_22248_12109# a_22869_12030# a_23077_12030# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1525 vdd a_9430_2317# a_9222_2317# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1526 a_28310_10642# a_28402_9007# a_28353_9197# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1527 a_574_2486# a_1195_2378# a_1403_2378# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1528 a_23075_5343# a_23915_6018# a_24123_6018# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1529 a_17347_4453# a_17434_5962# a_17389_5975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1530 a_1405_9833# a_984_9833# a_576_9941# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1531 gnd d0 a_9429_5284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1532 gnd d0 a_31105_9002# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1533 a_18839_8336# a_19932_8998# a_19883_9188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1534 a_25521_11467# a_25151_12793# a_24125_12026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1535 a_41557_5289# a_41553_5466# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1536 vdd d0 a_20137_5957# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1537 a_27246_7430# a_28359_10452# a_28310_10642# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1538 vdd a_20138_4437# a_19930_4437# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1539 a_39062_5973# a_40554_6727# a_40505_6917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1540 a_12112_13473# a_11691_13473# a_11283_13552# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1541 a_30846_2505# a_22249_2385# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1542 vdd a_20139_11286# a_19931_11286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1543 a_33784_2370# a_33363_2370# a_32955_2478# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1544 a_11281_7544# a_11902_7465# a_12110_7465# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1545 a_41560_8330# a_41813_8317# a_40508_8511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1546 a_2245_10508# a_2032_10508# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1547 gnd a_41810_7402# a_41602_7402# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1548 a_23075_6790# a_22654_6790# a_22246_6898# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1549 a_9173_2507# a_576_2387# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1550 a_33362_5337# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1551 a_36113_5334# a_35900_5334# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1552 vdd d1 a_8383_11296# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1553 vdd d3 a_39273_4438# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1554 a_18833_3952# a_19930_3758# a_19885_3771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1555 a_32954_5700# a_33575_6016# a_33783_6016# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1556 a_9176_6744# a_9429_6731# a_8124_6925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1557 a_23077_11351# a_22656_11351# a_22248_11459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1558 a_2242_6020# a_2029_6020# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1559 a_22868_3823# a_22655_3823# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1560 a_26605_4504# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1561 a_12110_5339# a_12950_6014# a_13158_6014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1562 a_9178_11984# a_9174_12161# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1563 a_34626_9053# a_34413_9053# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1564 a_3940_5342# a_4800_8377# a_5008_8377# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1565 a_30847_13606# a_30851_12750# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1566 a_11903_3819# a_11690_3819# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1567 a_15640_4500# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1568 vdd d0 a_9429_5284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1569 a_29804_8340# a_30897_9002# a_30852_9015# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1570 a_5145_4506# a_4932_4506# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1571 a_13160_13469# a_12739_13469# a_12112_12794# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1572 a_27246_7430# a_28359_10452# a_28314_10465# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1573 a_12738_4494# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1574 a_22656_12030# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1575 a_34832_4492# a_36071_3812# a_36222_5334# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1576 a_18836_6742# a_19929_7404# a_19884_7417# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1577 a_29798_2509# a_30895_2315# a_30846_2505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1578 a_984_10512# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1579 a_6637_10644# a_6729_9009# a_6680_9199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1580 vdd d0 a_41810_5955# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1581 a_11905_8380# a_11692_8380# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1582 a_41555_12153# a_41559_11297# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1583 vdd a_28609_11974# a_28401_11974# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1584 gnd a_20140_8319# a_19932_8319# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1585 a_9175_10641# a_9179_9785# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1586 a_9172_6921# a_9429_6731# a_8124_6925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1587 a_573_6359# a_1194_6792# a_1402_6792# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1588 a_33783_7463# a_34623_7459# a_34831_7459# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1589 a_11283_11710# a_11283_11455# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1590 a_1403_3057# a_982_3057# a_574_2741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1591 a_30852_10462# a_30848_10639# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1592 a_33785_11345# a_33364_11345# a_32957_10839# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1593 gnd a_8381_6735# a_8173_6735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1594 a_32957_9392# a_33578_9825# a_33786_9825# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1595 vdd a_30057_8327# a_29849_8327# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1596 vdd d2 a_39317_11968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1597 gnd a_17602_10448# a_17394_10448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1598 a_6680_9199# a_8176_8329# a_8131_8342# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1599 a_33785_12792# a_34625_13467# a_34833_13467# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1600 a_23918_9059# a_23705_9059# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1601 vdd d0 a_20140_8998# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1602 a_24125_12026# a_25364_12793# a_25521_11467# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1603 a_23915_7465# a_23702_7465# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1604 gnd a_31105_9002# a_30897_9002# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1605 a_33576_3049# a_33363_3049# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1606 a_573_6359# a_573_6103# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1607 vdd a_20137_5957# a_19929_5957# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1608 a_22870_9831# a_22657_9831# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1609 a_8131_8342# a_9224_9004# a_9175_9194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1610 a_29798_2509# a_30895_2315# a_30850_2328# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1611 a_30851_12750# a_30847_12927# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1612 a_24124_3051# a_25363_3818# a_25514_5340# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1613 a_28357_9020# a_29849_9774# a_29800_9964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1614 vdd d1 a_40765_9768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1615 a_32955_3925# a_32955_3384# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1616 a_10906_219# a_10693_219# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1617 a_32957_10583# a_33578_10504# a_33786_10504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1618 a_2453_10508# a_3692_9828# a_3843_11350# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1619 a_34831_6012# a_34410_6012# a_33783_5337# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1620 a_1404_11353# a_983_11353# a_576_10847# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1621 a_11905_10506# a_11692_10506# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1622 vdd a_39273_4438# a_39065_4438# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1623 a_12112_12026# a_11691_12026# a_11283_11710# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1624 a_982_4504# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1625 a_22246_6898# a_22246_6357# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1626 vdd a_8381_6735# a_8173_6735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1627 a_22655_3823# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1628 a_34832_4492# a_34411_4492# a_33784_3817# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1629 a_32688_217# a_37313_4498# a_37389_8369# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1630 a_9174_13608# a_9431_13418# a_8130_12756# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1631 a_34413_9053# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1632 a_11690_3819# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1633 a_22246_6898# a_22867_6790# a_23075_6790# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1634 a_39022_10459# a_39275_10446# a_37954_7424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1635 a_25514_5340# a_25405_5340# a_25613_5340# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1636 a_36070_6779# a_35857_6779# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1637 a_6681_5981# a_6934_5968# a_6639_4459# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1638 a_25516_11348# a_25407_11348# a_25615_11348# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1639 a_1195_3825# a_982_3825# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1640 a_13158_7461# a_14397_6781# a_14554_5455# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1641 a_26681_8375# a_26260_8375# a_25615_11348# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1642 a_40512_8334# a_41605_8996# a_41560_9009# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1643 a_21652_206# a_21543_206# vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1644 vdd d0 a_20137_5278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1645 gnd d0 a_20138_4437# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1646 a_28357_9020# a_29849_9774# a_29804_9787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1647 a_576_10591# a_1197_10512# a_1405_10512# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1648 a_983_13479# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1649 a_23077_11351# a_23917_12026# a_24125_12026# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1650 gnd d1 a_19092_9770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1651 vdd a_41811_2309# a_41603_2309# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1652 a_11692_8380# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1653 a_9179_8338# a_9175_8515# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1654 a_22248_13161# a_22869_13477# a_23077_13477# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1655 a_32955_3128# a_33576_3049# a_33784_3049# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1656 a_576_10591# a_576_10196# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1657 a_8124_5478# a_8381_5288# a_6677_6158# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1658 a_30849_7421# a_30845_7598# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1659 gnd d1 a_8384_8329# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1660 gnd d0 a_41810_5276# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1661 gnd d0 a_20139_13412# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1662 a_12111_3051# a_12951_3047# a_13159_3047# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1663 a_3732_5342# a_3519_5342# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1664 gnd a_30056_11294# a_29848_11294# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1665 a_14549_5336# a_14440_5336# a_14648_5336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1666 a_9176_7423# a_9172_7600# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1667 gnd a_20139_12733# a_19931_12733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1668 a_41556_9954# a_41560_9009# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1669 a_8125_3958# a_8382_3768# a_6682_3014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1670 gnd d4 a_16534_7413# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1671 a_39018_10636# a_39275_10446# a_37954_7424# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1672 a_39058_6150# a_39315_5960# a_39020_4451# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1673 a_32954_6892# a_32954_6351# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1674 a_23705_9059# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1675 a_22867_6790# a_22654_6790# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1676 a_23702_7465# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1677 a_41558_4448# a_41811_4435# a_40510_3773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1678 a_33363_3049# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1679 a_35857_6779# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1680 a_2031_13475# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1681 gnd a_40762_5280# a_40554_5280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1682 a_2452_12028# a_2031_12028# a_1404_12032# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1683 vdd d1 a_19092_9770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1684 a_12113_10506# a_11692_10506# a_11284_10585# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1685 a_33784_2370# a_34624_3045# a_34832_3045# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1686 a_2242_7467# a_2029_7467# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1687 a_574_3933# a_1195_3825# a_1403_3825# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1688 a_575_13558# a_575_13163# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1689 vdd d0 a_41810_5276# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1690 vdd d0 a_20139_13412# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1691 gnd d0 a_9429_6731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1692 a_5008_8377# a_4587_8377# a_3942_11350# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1693 vdd d1 a_19091_12737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1694 a_23078_9063# a_22657_9063# a_22249_9142# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1695 a_25516_11348# a_25152_9826# a_24126_9059# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1696 vdd a_20139_12733# a_19931_12733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1697 a_23704_12026# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1698 vdd a_8383_11296# a_8175_11296# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1699 a_33784_3817# a_33363_3817# a_32955_3925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1700 vdd d4 a_16534_7413# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1701 a_22656_13477# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1702 a_29798_2509# a_30055_2319# a_28351_3189# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1703 a_12110_7465# a_11689_7465# a_11281_7544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1704 a_25362_6785# a_25149_6785# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1705 a_33364_11345# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1706 a_9179_9785# a_9432_9772# a_8127_9966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1707 gnd d2 a_17644_11970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1708 gnd d1 a_30057_8327# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1709 vdd d2 a_17645_9003# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1710 vdd d0 a_31104_11290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1711 gnd a_9430_2317# a_9222_2317# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1712 a_19882_12155# a_19886_11299# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1713 a_22247_3134# a_22247_2739# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1714 a_41554_4625# a_41811_4435# a_40510_3773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1715 a_3477_3820# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1716 a_41555_11474# a_41560_10456# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1717 a_33577_13471# a_33364_13471# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1718 a_30850_3007# a_31103_2994# a_29802_2332# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1719 vdd a_40762_5280# a_40554_5280# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1720 a_32957_8741# a_32957_8486# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1721 a_19886_11978# a_20139_11965# a_18838_11303# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1722 vdd a_20137_5278# a_19929_5278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1723 gnd a_20138_4437# a_19930_4437# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1724 a_575_13558# a_1196_13479# a_1404_13479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1725 a_11689_5339# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1726 a_19880_6147# a_19884_5291# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1727 gnd a_19092_9770# a_18884_9770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1728 a_22248_13161# a_22248_12906# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1729 vdd d0 a_9429_6731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1730 a_2029_7467# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1731 vdd a_9431_11971# a_9223_11971# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1732 a_11114_219# a_10693_219# a_11015_219# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1733 a_18833_3952# a_19930_3758# a_19881_3948# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1734 gnd d3 a_39273_4438# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1735 a_1403_3825# a_2243_4500# a_2451_4500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1736 gnd d0 a_31103_3762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1737 a_24125_13473# a_23704_13473# a_23077_12798# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1738 a_39022_10459# a_39109_11968# a_39060_12158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1739 a_9175_9962# a_9432_9772# a_8127_9966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1740 a_23076_2376# a_22655_2376# a_22247_2484# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1741 a_30852_8336# a_31105_8323# a_29800_8517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1742 a_14229_11344# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1743 gnd a_16534_7413# a_16326_7413# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1744 a_9177_2330# a_9173_2507# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1745 gnd a_8384_9776# a_8176_9776# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1746 a_33786_9825# a_34626_10500# a_34834_10500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1747 a_11282_3386# a_11903_3819# a_12111_3819# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1748 a_22654_6790# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1749 a_30851_11982# a_30847_12159# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1750 a_34831_7459# a_34410_7459# a_33783_7463# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1751 a_1403_4504# a_982_4504# a_574_4188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1752 a_22246_5706# a_22867_6022# a_23075_6022# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1753 a_8126_11486# a_9223_11292# a_9178_11305# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1754 a_32955_3128# a_32955_2733# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1755 a_17349_10461# a_17436_11970# a_17387_12160# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1756 vdd a_19092_9770# a_18884_9770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1757 a_3689_6787# a_3476_6787# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1758 a_574_4839# a_574_4583# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1759 gnd a_28567_10452# a_28359_10452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1760 a_33576_4496# a_33363_4496# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1761 a_2031_12028# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1762 vdd d0 a_31103_3762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1763 a_15716_8371# a_15295_8371# a_14648_5336# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1764 a_30848_8513# a_31105_8323# a_29800_8517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1765 a_11283_11455# a_11284_10841# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1766 vdd a_16534_7413# a_16326_7413# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1767 a_30848_10639# a_31105_10449# a_29804_9787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1768 vdd a_8384_9776# a_8176_9776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1769 gnd a_30057_8327# a_29849_8327# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1770 vdd d4 a_5826_7419# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1771 a_41553_6145# a_41810_5955# a_40509_5293# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1772 a_1404_12800# a_983_12800# a_575_12367# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1773 a_11284_9935# a_11284_9394# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1774 a_6680_9199# a_8176_8329# a_8127_8519# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1775 gnd a_17643_2995# a_17435_2995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1776 a_30849_5295# a_30845_5472# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1777 gnd d2 a_6935_3001# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1778 a_12110_6018# a_11689_6018# a_11281_5702# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1779 a_22249_9398# a_22870_9831# a_23078_9831# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1780 a_14227_5336# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1781 a_9176_5297# a_9172_5474# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1782 a_13161_9055# a_14400_9822# a_14551_11344# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1783 gnd d0 a_9431_11971# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1784 gnd d1 a_40765_9768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1785 a_22249_10194# a_22870_10510# a_23078_10510# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1786 vdd a_28567_10452# a_28359_10452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1787 a_33577_12024# a_33364_12024# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1788 a_32955_2733# a_32955_2478# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1789 a_12111_4498# a_11690_4498# a_11282_4182# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1790 a_17385_6152# a_18881_5282# a_18832_5472# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1791 a_25363_3818# a_25150_3818# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1792 gnd a_9431_11292# a_9223_11292# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1793 a_11282_4577# a_11282_4182# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1794 gnd a_39273_4438# a_39065_4438# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1795 a_39020_4451# a_39107_5960# a_39058_6150# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1796 gnd a_31103_3762# a_30895_3762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1797 a_981_5345# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1798 a_8125_3958# a_9222_3764# a_9173_3954# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1799 a_40508_9958# a_40765_9768# a_39065_9014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1800 a_9178_13431# a_9431_13418# a_8130_12756# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1801 gnd d0 a_41810_6723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1802 a_575_11461# a_576_10847# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1803 a_34413_10500# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1804 a_41554_2499# a_32957_2379# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1805 a_41553_6145# a_41557_5289# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1806 a_2030_3053# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1807 gnd a_30056_12741# a_29848_12741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1808 a_14551_11344# a_14442_11344# a_14650_11344# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1809 a_2032_10508# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1810 gnd d0 a_20137_5278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1811 a_3476_6787# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1812 a_1196_12032# a_983_12032# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1813 a_12113_9827# a_11692_9827# a_11284_9394# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1814 a_33576_2370# a_33363_2370# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1815 a_11902_7465# a_11689_7465# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1816 a_12112_11347# a_12952_12022# a_13160_12022# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1817 a_33363_4496# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1818 a_17385_6152# a_18881_5282# a_18836_5295# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1819 a_19882_11476# a_19887_10458# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1820 vdd d2 a_6936_11976# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1821 gnd a_41813_10443# a_41605_10443# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1822 vdd a_31103_3762# a_30895_3762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1823 a_33784_3817# a_34624_4492# a_34832_4492# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1824 a_3846_5461# a_3732_5342# a_3940_5342# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1825 a_29801_5299# a_30894_5961# a_30845_6151# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1826 a_11281_6353# a_11281_6097# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1827 vout a_21330_206# a_11114_219# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1828 a_8125_3958# a_9222_3764# a_9177_3777# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1829 a_19880_5468# a_19885_4450# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1830 a_576_10847# a_576_10591# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1831 a_22657_10510# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1832 vdd d0 a_41811_2988# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1833 a_22247_3134# a_22868_3055# a_23076_3055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1834 vdd d0 a_41810_6723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1835 vdd a_5826_7419# a_5618_7419# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1836 a_8129_3781# a_8382_3768# a_6682_3014# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1837 a_32954_5700# a_32954_5445# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1838 vdd a_30056_12741# a_29848_12741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1839 a_41557_5289# a_41810_5276# a_40505_5470# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1840 a_33578_10504# a_33365_10504# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1841 gnd a_6935_3001# a_6727_3001# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1842 a_984_9065# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1843 a_33364_12792# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1844 a_22868_2376# a_22655_2376# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1845 a_28356_11987# a_28609_11974# a_28314_10465# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1846 vdd a_31104_11969# a_30896_11969# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1847 a_30850_4454# a_31103_4441# a_29802_3779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1848 vdd a_40762_6727# a_40554_6727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1849 a_19886_13425# a_20139_13412# a_18838_12750# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1850 a_5569_7609# a_6684_4446# a_6635_4636# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1851 a_1197_8386# a_984_8386# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1852 a_25150_3818# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1853 gnd d1 a_19091_12737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1854 vdd a_41813_10443# a_41605_10443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1855 vref a_575_13558# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1856 a_23076_2376# a_23916_3051# a_24124_3051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1857 a_29800_9964# a_30897_9770# a_30848_9960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1858 a_24126_10506# a_23705_10506# a_23078_9831# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1859 a_29802_2332# a_30055_2319# a_28351_3189# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1860 a_1197_10512# a_984_10512# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1861 a_34412_13467# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1862 a_11284_10841# a_11904_11347# a_12112_11347# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1863 a_39063_3006# a_40555_3760# a_40506_3950# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1864 gnd d1 a_40764_11288# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1865 a_22249_9939# a_22249_9398# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1866 a_41553_5466# a_41810_5276# a_40505_5470# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1867 a_6641_10467# a_6728_11976# a_6683_11989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1868 a_32957_8486# a_32954_7798# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1869 a_22657_9063# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1870 gnd a_28607_5966# a_28399_5966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1871 a_14650_11344# a_14229_11344# a_14551_11344# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1872 a_23076_3823# a_22655_3823# a_22247_3931# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1873 a_33363_2370# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1874 gnd a_20137_5278# a_19929_5278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1875 a_14549_5336# a_14185_3814# a_13159_4494# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1876 a_12953_10502# a_12740_10502# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1877 a_30846_4631# a_31103_4441# a_29802_3779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1878 a_19882_13602# a_20139_13412# a_18838_12750# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1879 a_3692_9828# a_3479_9828# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1880 a_17388_9193# a_17645_9003# a_17345_10638# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1881 a_982_2378# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1882 a_5569_7609# a_6684_4446# a_6639_4459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1883 a_1194_7471# a_981_7471# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1884 a_3691_12795# a_3478_12795# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1885 a_13160_12022# a_12739_12022# a_12112_11347# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1886 a_23075_7469# a_22654_7469# a_22246_7153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1887 a_2453_9061# a_2032_9061# a_1405_9065# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1888 a_22247_4581# a_22247_4186# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1889 a_41555_12921# a_41559_11976# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1890 a_11284_9138# a_11284_8743# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1891 a_29800_9964# a_30897_9770# a_30852_9783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1892 a_11902_6018# a_11689_6018# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1893 a_40509_5293# a_41602_5955# a_41553_6145# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1894 a_14186_12789# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1895 a_25613_5340# a_25192_5340# a_25514_5340# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1896 a_39063_3006# a_40555_3760# a_40510_3773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1897 a_34625_12020# a_34412_12020# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1898 a_25194_11348# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1899 a_33783_6016# a_34623_6012# a_34831_6012# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1900 a_11903_4498# a_11690_4498# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1901 a_21652_206# a_32366_217# a_27026_4504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1902 a_1402_5345# a_981_5345# a_574_4839# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1903 a_23077_12798# a_22656_12798# a_22248_12906# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1904 a_2450_7467# a_3689_6787# a_3846_5461# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1905 a_29803_11307# a_30896_11969# a_30847_12159# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1906 a_22249_10194# a_22249_9939# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1907 a_32366_217# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1908 a_19887_9011# a_19883_9188# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1909 a_11282_2480# a_11284_2381# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1910 a_37389_8369# a_37526_4498# a_32688_217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1911 a_28352_12164# a_29848_11294# a_29799_11484# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1912 a_36115_11342# a_35902_11342# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1913 a_30850_3775# a_30846_3952# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1914 a_33786_8378# a_33365_8378# a_32954_7798# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1915 a_22655_2376# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1916 a_11691_11347# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1917 vdd d0 a_9430_2996# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1918 a_9175_9194# a_9179_8338# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1919 a_39060_12158# a_40556_11288# a_40507_11478# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1920 a_32956_13155# a_33577_13471# a_33785_13471# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1921 a_3734_11350# a_3521_11350# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1922 a_24123_7465# a_23702_7465# a_23075_7469# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1923 a_12951_3047# a_12738_3047# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1924 a_33575_5337# a_33362_5337# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1925 a_11904_13473# a_11691_13473# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1926 gnd a_31104_11290# a_30896_11290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1927 a_9177_3777# a_9173_3954# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1928 a_36227_5453# a_35857_6779# a_34831_7459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1929 a_41553_5466# a_41558_4448# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1930 a_28312_4457# a_28399_5966# a_28350_6156# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1931 a_25613_5340# a_26473_8375# a_26681_8375# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1932 a_576_8749# a_1197_9065# a_1405_9065# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1933 a_22246_6357# a_22246_6101# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1934 a_2244_12028# a_2031_12028# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1935 a_26818_4504# a_26605_4504# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1936 a_11905_9827# a_11692_9827# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1937 a_573_7550# a_1194_7471# a_1402_7471# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1938 a_39018_10636# a_39110_9001# a_39061_9191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1939 a_1196_13479# a_983_13479# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1940 a_30852_10462# a_31105_10449# a_29804_9787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1941 a_40508_9958# a_41605_9764# a_41556_9954# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1942 gnd d4 a_5826_7419# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1943 a_22869_11351# a_22656_11351# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1944 a_19884_5970# a_20137_5957# a_18836_5295# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1945 a_11284_8743# a_11284_8488# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1946 vdd a_8381_5288# a_8173_5288# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1947 a_981_6792# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1948 gnd a_39317_11968# a_39109_11968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1949 a_13161_10502# a_12740_10502# a_12113_10506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1950 gnd d1 a_8381_5288# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1951 a_33783_7463# a_33362_7463# a_32954_7542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1952 a_21543_206# a_21330_206# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1953 vdd d2 a_39318_9001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1954 a_13158_7461# a_12737_7461# a_12110_7465# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1955 a_12952_13469# a_12739_13469# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1956 a_30845_6151# a_31102_5961# a_29801_5299# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1957 gnd a_9429_5963# a_9221_5963# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1958 a_5569_7609# a_5826_7419# a_5254_4506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1959 a_11283_12902# a_11283_12361# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1960 a_12112_12794# a_11691_12794# a_11283_12361# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1961 a_19883_9188# a_19887_8332# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1962 gnd a_19089_5282# a_18881_5282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1963 gnd a_17644_11970# a_17436_11970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1964 a_14400_9822# a_14187_9822# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1965 gnd d2 a_17642_5962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1966 a_28353_9197# a_29849_8327# a_29804_8340# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1967 a_6682_3014# a_6935_3001# a_6635_4636# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1968 gnd d0 a_20137_6725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1969 vdd d0 a_9431_13418# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1970 a_983_12032# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1971 gnd d3 a_39275_10446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1972 a_40508_9958# a_41605_9764# a_41560_9777# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1973 a_32954_5445# a_33575_5337# a_33783_5337# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1974 a_1194_6024# a_981_6024# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1975 a_17389_5975# a_18881_6729# a_18836_6742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1976 vdd a_9431_12739# a_9223_12739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1977 a_576_2387# a_1195_2378# a_1403_2378# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1978 a_32954_6351# a_32954_6095# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1979 a_40512_9781# a_40765_9768# a_39065_9014# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1980 gnd a_6936_11976# a_6728_11976# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1981 a_11282_4833# a_11282_4577# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1982 a_18836_5295# a_19929_5957# a_19884_5970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1983 a_33578_9057# a_33365_9057# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1984 a_19881_3948# a_19885_3003# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1985 a_11690_4498# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1986 a_1404_13479# a_2244_13475# a_2452_13475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1987 a_22247_4581# a_22868_4502# a_23076_4502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1988 a_25519_5459# a_25149_6785# a_24123_6018# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1989 a_22248_13556# a_22248_13161# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1990 a_41558_2322# a_41554_2499# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1991 a_11281_7149# a_11902_7465# a_12110_7465# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1992 a_17343_4630# a_17435_2995# a_17390_3008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1993 a_5353_4506# a_4932_4506# a_5254_4506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1994 a_41557_6736# a_41810_6723# a_40505_6917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1995 a_33362_5337# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1996 vdd a_19089_5282# a_18881_5282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1997 vdd d0 a_20138_2990# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1998 gnd d1 a_30054_5286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1999 a_573_6103# a_573_5708# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2000 vdd d0 a_20137_6725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2001 vdd d3 a_39275_10446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2002 a_22249_9142# a_22249_8747# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2003 a_22868_3823# a_22655_3823# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2004 a_26605_4504# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2005 a_11692_9827# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2006 a_32956_12103# a_33577_12024# a_33785_12024# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2007 a_24123_6018# a_23702_6018# a_23075_5343# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2008 a_34626_9053# a_34413_9053# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2009 a_11904_12026# a_11691_12026# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2010 a_1197_9833# a_984_9833# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2011 gnd a_5826_7419# a_5618_7419# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2012 a_576_9400# a_576_9144# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2013 a_29801_6746# a_30894_7408# a_30849_7421# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2014 a_13160_13469# a_12739_13469# a_12112_13473# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2015 a_22867_7469# a_22654_7469# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2016 a_34832_3045# a_36071_3812# a_36222_5334# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2017 a_24124_4498# a_23703_4498# a_23076_3823# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2018 vdd a_39318_9001# a_39110_9001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2019 a_984_10512# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2020 vdd a_17642_5962# a_17434_5962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2021 a_30852_8336# a_30848_8513# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2022 a_11283_12361# a_11904_12794# a_12112_12794# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2023 a_41554_3178# a_41811_2988# a_40510_2326# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2024 gnd d1 a_40764_12735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2025 a_41553_6913# a_41810_6723# a_40505_6917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2026 a_12740_10502# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2027 vdd d2 a_6934_5968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2028 a_11281_7800# a_11281_7544# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2029 vdd d1 a_30054_5286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2030 a_30849_5295# a_31102_5282# a_29797_5476# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2031 gnd d0 a_9432_9004# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2032 gnd a_40762_6727# a_40554_6727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2033 a_33783_6016# a_33362_6016# a_32954_5700# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2034 a_33783_6784# a_34623_7459# a_34831_7459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2035 a_575_12111# a_1196_12032# a_1404_12032# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2036 gnd a_20137_6725# a_19929_6725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2037 a_28310_10642# a_28402_9007# a_28357_9020# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2038 a_41555_13600# a_41559_12744# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2039 a_1403_3057# a_982_3057# a_574_3136# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2040 a_13158_6014# a_12737_6014# a_12110_5339# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2041 a_3846_5461# a_3476_6787# a_2450_6020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2042 a_33785_11345# a_33364_11345# a_32956_11453# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2043 a_22870_10510# a_22657_10510# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2044 a_37635_4498# a_37999_7411# a_37950_7601# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2045 a_8130_11309# a_8383_11296# a_6679_12166# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2046 a_18839_8336# a_19932_8998# a_19887_9011# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2047 a_982_3825# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2048 a_2029_6020# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2049 a_33784_4496# a_33363_4496# a_32955_4180# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2050 a_5573_7432# a_6686_10454# a_6637_10644# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2051 a_30850_3007# a_30846_3184# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2052 a_30845_6151# a_30849_5295# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2053 a_33365_9057# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2054 a_13159_4494# a_12738_4494# a_12111_3819# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2055 a_23915_7465# a_23702_7465# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2056 a_22249_8747# a_22249_8492# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2057 a_18833_2505# a_19930_2311# a_19881_2501# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2058 a_33786_9057# a_34626_9053# a_34834_9053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2059 a_9172_6153# a_9176_5297# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2060 vdd d1 a_40764_12735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2061 a_30845_5472# a_31102_5282# a_29797_5476# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2062 a_32957_10188# a_33578_10504# a_33786_10504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2063 a_2453_9061# a_3692_9828# a_3843_11350# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2064 a_1405_8386# a_984_8386# a_576_8494# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2065 a_34831_6012# a_34410_6012# a_33783_6016# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2066 a_41560_10456# a_41556_10633# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2067 a_11905_10506# a_11692_10506# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2068 gnd a_30054_5286# a_29846_5286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2069 a_22248_12906# a_22869_12798# a_23077_12798# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2070 a_1404_11353# a_983_11353# a_575_11461# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2071 vdd a_20138_2990# a_19930_2990# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2072 vdd a_20137_6725# a_19929_6725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2073 a_29803_12754# a_30896_13416# a_30847_13606# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2074 a_28356_11987# a_29848_12741# a_29799_12931# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2075 a_12112_12026# a_11691_12026# a_11283_12105# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2076 a_6677_6158# a_8173_5288# a_8124_5478# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2077 a_37635_4498# a_37999_7411# a_37954_7424# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2078 a_33786_9825# a_33365_9825# a_32957_9392# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2079 vdd d0 a_41812_11963# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2080 a_22655_3823# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2081 a_11691_12794# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2082 a_39064_11981# a_40556_12735# a_40507_12925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2083 a_11281_6097# a_11902_6018# a_12110_6018# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2084 gnd a_41810_5955# a_41602_5955# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2085 a_34413_9053# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2086 a_5573_7432# a_6686_10454# a_6641_10467# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2087 a_12951_4494# a_12738_4494# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2088 a_33575_6784# a_33362_6784# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2089 a_22247_4837# a_22247_4581# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2090 a_18832_5472# a_19929_5278# a_19884_5291# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2091 a_41559_12744# a_41555_12921# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2092 a_18833_2505# a_19930_2311# a_19885_2324# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2093 a_11282_4577# a_11903_4498# a_12111_4498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2094 a_6637_10644# a_6729_9009# a_6684_9022# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2095 a_40509_6740# a_41602_7402# a_41557_7415# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2096 a_19887_9011# a_20140_8998# a_18839_8336# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2097 a_22654_7469# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2098 vdd a_8384_8329# a_8176_8329# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2099 a_576_10196# a_1197_10512# a_1405_10512# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2100 a_983_13479# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2101 a_32955_2733# a_33576_3049# a_33784_3049# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2102 vdd a_6934_5968# a_6726_5968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2103 a_2243_3053# a_2030_3053# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2104 vdd a_30054_5286# a_29846_5286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2105 gnd a_9432_9004# a_9224_9004# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2106 a_36224_11342# a_35860_9820# a_34834_9053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2107 a_29803_12754# a_30896_13416# a_30851_13429# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2108 a_12111_2372# a_12951_3047# a_13159_3047# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2109 a_36323_11342# a_37181_8369# a_37389_8369# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2110 a_28356_11987# a_29848_12741# a_29803_12754# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2111 a_17345_10638# a_17437_9003# a_17388_9193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2112 gnd d1 a_8381_6735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2113 a_28312_4457# a_28565_4444# a_27242_7607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2114 a_3732_5342# a_3519_5342# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2115 a_39064_11981# a_40556_12735# a_40511_12748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2116 vdd d0 a_31105_10449# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2117 a_23078_8384# a_22657_8384# a_22246_7804# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2118 a_2450_7467# a_2029_7467# a_1402_6792# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2119 gnd a_9429_7410# a_9221_7410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2120 gnd d0 a_20140_9766# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2121 gnd d1 a_40765_8321# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2122 a_22248_11459# a_22249_10845# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2123 a_12113_8380# a_11692_8380# a_11284_8488# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2124 vdd a_31104_12737# a_30896_12737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2125 a_12111_3051# a_11690_3051# a_11282_2735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2126 a_32954_6095# a_32954_5700# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2127 a_26473_8375# a_26260_8375# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2128 a_22656_12798# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2129 a_12110_6786# a_11689_6786# a_11281_6353# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2130 a_8131_9789# a_9224_10451# a_9175_10641# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2131 a_23702_7465# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2132 a_23917_13473# a_23704_13473# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2133 a_35857_6779# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2134 a_40511_11301# a_41604_11963# a_41559_11976# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2135 a_1405_10512# a_2245_10508# a_2453_10508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2136 a_32955_4831# a_32955_4575# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2137 a_11284_10841# a_11284_10585# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2138 a_33577_12792# a_33364_12792# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2139 a_39059_3183# a_39316_2993# a_39016_4628# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2140 a_33785_11345# a_34625_12020# a_34833_12020# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2141 a_19880_7594# a_20137_7404# a_18836_6742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2142 a_574_3392# a_1195_3825# a_1403_3825# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2143 a_23915_6018# a_23702_6018# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2144 a_5573_7432# a_5826_7419# a_5254_4506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2145 vdd d1 a_8381_6735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2146 a_22870_8384# a_22657_8384# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2147 a_25516_11348# a_25152_9826# a_24126_10506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2148 a_28308_4634# a_28565_4444# a_27242_7607# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2149 a_36229_11461# a_36115_11342# a_36323_11342# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2150 vdd a_9429_7410# a_9221_7410# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2151 a_28353_9197# a_29849_8327# a_29800_8517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2152 a_14442_11344# a_14229_11344# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2153 gnd a_40764_11288# a_40556_11288# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2154 vdd d1 a_40765_8321# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2155 vdd d0 a_20140_9766# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2156 a_23916_4498# a_23703_4498# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2157 gnd d0 a_9431_13418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2158 gnd d0 a_41812_11284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2159 a_34834_10500# a_34413_10500# a_33786_9825# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2160 a_8131_9789# a_9224_10451# a_9179_10464# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2161 a_33362_6784# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2162 vdd a_19089_6729# a_18881_6729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2163 gnd d1 a_30054_6733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2164 a_17389_5975# a_18881_6729# a_18832_6919# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2165 a_11281_7149# a_11281_6894# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2166 gnd d0 a_41813_8996# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2167 gnd a_9431_12739# a_9223_12739# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2168 a_32956_13155# a_32956_12900# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2169 a_8125_2511# a_9222_2317# a_9177_2330# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2170 a_17389_5975# a_17642_5962# a_17347_4453# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2171 a_34832_3045# a_34411_3045# a_33784_2370# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2172 a_575_13163# a_1196_13479# a_1404_13479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2173 a_11689_5339# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2174 a_22246_5451# a_22867_5343# a_23075_5343# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2175 a_8129_2334# a_8382_2321# a_6678_3191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2176 a_29804_9787# a_30057_9774# a_28357_9020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2177 a_2029_7467# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2178 a_2030_4500# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2179 a_11114_219# a_10693_219# a_5353_4506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2180 a_33576_3817# a_33363_3817# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2181 a_34833_13467# a_36072_12787# a_36229_11461# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2182 gnd d1 a_19092_8323# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2183 vdd d0 a_41812_11284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2184 a_24125_13473# a_23704_13473# a_23077_13477# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2185 a_14399_12789# a_14186_12789# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2186 a_22248_11714# a_22869_12030# a_23077_12030# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2187 a_9172_5474# a_9177_4456# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2188 a_13161_9055# a_12740_9055# a_12113_8380# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2189 vdd d1 a_30054_6733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2190 a_26260_8375# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2191 a_19887_10458# a_19883_10635# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2192 a_2032_9061# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2193 gnd a_19091_11290# a_18883_11290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2194 a_35902_11342# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2195 a_41558_3769# a_41554_3946# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2196 a_1403_4504# a_982_4504# a_574_4583# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2197 a_33785_12792# a_33364_12792# a_32956_12900# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2198 gnd d0 a_31102_7408# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2199 a_40507_11478# a_41604_11284# a_41555_11474# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2200 a_8130_12756# a_8383_12743# a_6683_11989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2201 a_8125_2511# a_8382_2321# a_6678_3191# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2202 gnd d0 a_41811_2309# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2203 a_573_7550# a_573_7155# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2204 a_29800_9964# a_30057_9774# a_28357_9020# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2205 a_34412_12020# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2206 a_23078_10510# a_22657_10510# a_22249_10194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2207 a_33364_13471# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2208 a_23702_6018# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2209 a_36071_3812# a_35858_3812# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2210 a_9177_3009# a_9430_2996# a_8129_2334# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2211 a_2452_13475# a_3691_12795# a_3848_11469# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2212 a_19886_12746# a_19882_12923# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2213 a_2031_12028# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2214 vdd a_27499_7417# a_27291_7417# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2215 vdd d1 a_19092_8323# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2216 a_15716_8371# a_15295_8371# a_14650_11344# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2217 a_2242_6020# a_2029_6020# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2218 a_41559_11976# a_41555_12153# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2219 a_23703_4498# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2220 a_34833_13467# a_34412_13467# a_33785_12792# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2221 a_30845_6919# a_31102_6729# a_29797_6923# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2222 a_19884_6738# a_19880_6915# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2223 a_3521_11350# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2224 a_41560_10456# a_41813_10443# a_40512_9781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2225 vdd d1 a_19091_11290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2226 a_11284_9138# a_11905_9059# a_12113_9059# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2227 gnd a_30054_6733# a_29846_6733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2228 a_34623_7459# a_34410_7459# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2229 gnd a_41813_8996# a_41605_8996# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2230 a_6677_6158# a_6934_5968# a_6639_4459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2231 gnd a_41812_11963# a_41604_11963# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2232 a_23075_6022# a_22654_6022# a_22246_5706# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2233 a_35859_12787# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2234 gnd d2 a_39315_5960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2235 a_6681_5981# a_8173_6735# a_8124_6925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2236 a_40507_11478# a_41604_11284# a_41559_11297# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2237 a_23076_3823# a_23916_4498# a_24124_4498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2238 a_8126_12933# a_8383_12743# a_6683_11989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2239 a_22656_12030# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2240 gnd d0 a_9430_3764# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2241 a_12110_6018# a_11689_6018# a_11281_6097# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2242 a_9179_8338# a_9432_8325# a_8127_8519# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2243 a_4587_8377# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2244 a_11905_8380# a_11692_8380# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2245 a_39065_9014# a_39318_9001# a_39018_10636# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2246 a_33577_12024# a_33364_12024# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2247 a_11903_3051# a_11690_3051# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2248 a_11902_6786# a_11689_6786# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2249 a_9174_12161# a_9431_11971# a_8130_11309# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2250 a_41556_10633# a_41560_9777# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2251 a_25363_3818# a_25150_3818# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2252 a_9175_9962# a_9179_9017# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2253 a_33363_3817# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2254 a_12737_7461# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2255 a_14556_11463# a_14186_12789# a_13160_13469# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2256 gnd a_19092_8323# a_18884_8323# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2257 a_41556_10633# a_41813_10443# a_40512_9781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2258 vdd d0 a_31105_9002# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2259 a_32955_4180# a_33576_4496# a_33784_4496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2260 a_3478_12795# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2261 a_25615_11348# a_25194_11348# a_25516_11348# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2262 a_2243_4500# a_2030_4500# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2263 vdd a_30054_6733# a_29846_6733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2264 a_12111_3819# a_12951_4494# a_13159_4494# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2265 a_6681_5981# a_8173_6735# a_8128_6748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2266 a_23918_10506# a_23705_10506# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2267 a_18832_5472# a_19929_5278# a_19880_5468# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2268 a_23078_9831# a_22657_9831# a_22249_9398# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2269 vdd d0 a_9430_3764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2270 gnd d0 a_31103_2315# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2271 vdd a_41810_7402# a_41602_7402# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2272 gnd a_31102_7408# a_30894_7408# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2273 a_9175_8515# a_9432_8325# a_8127_8519# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2274 a_24125_12026# a_23704_12026# a_23077_11351# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2275 a_14551_11344# a_14187_9822# a_13161_9055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2276 a_12113_9827# a_11692_9827# a_11284_9935# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2277 a_23077_13477# a_22656_13477# a_22248_13161# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2278 a_1196_12032# a_983_12032# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2279 gnd a_8384_8329# a_8176_8329# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2280 a_11283_12361# a_11283_12105# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2281 a_10693_219# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2282 a_14397_6781# a_14184_6781# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2283 a_9174_11482# a_9179_10464# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2284 vdd a_19092_8323# a_18884_8323# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2285 a_19885_3003# a_20138_2990# a_18837_2328# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2286 a_3841_5342# a_3732_5342# a_3940_5342# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2287 gnd d0 a_31105_10449# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2288 a_12952_12022# a_12739_12022# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2289 a_22247_2739# a_22868_3055# a_23076_3055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2290 a_24123_7465# a_25362_6785# a_25519_5459# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2291 gnd a_31104_12737# a_30896_12737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2292 a_34410_7459# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2293 gnd a_39315_5960# a_39107_5960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X2294 vdd d0 a_31103_2315# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2295 a_35860_9820# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
C0 d2 d1 23.33fF
C1 d1 d0 26.82fF
C2 d5 d4 24.94fF
C3 d2 d3 31.17fF
C4 d3 d4 28.04fF
C5 d2 vdd 20.62fF
C6 d0 vdd 42.34fF
C7 d3 d5 6.33fF
C8 d1 vdd 37.50fF
C9 d3 vdd 22.44fF
C10 a_21652_206# gnd 12.30fF
C11 d7 gnd 23.31fF
C12 a_11114_219# gnd 12.71fF
C13 d6 gnd 43.69fF
C14 a_41554_2499# gnd 2.27fF
C15 a_40506_2503# gnd 2.80fF
C16 a_32957_2379# gnd 17.59fF
C17 a_30846_2505# gnd 2.27fF
C18 a_29798_2509# gnd 2.80fF
C19 a_32955_2478# gnd 2.28fF
C20 a_22249_2385# gnd 17.59fF
C21 a_19881_2501# gnd 2.27fF
C22 a_18833_2505# gnd 2.80fF
C23 a_22247_2484# gnd 2.28fF
C24 a_11284_2381# gnd 17.59fF
C25 a_9173_2507# gnd 2.27fF
C26 a_8125_2511# gnd 2.80fF
C27 a_11282_2480# gnd 2.28fF
C28 a_576_2387# gnd 17.59fF
C29 a_574_2486# gnd 2.28fF
C30 a_41558_2322# gnd 3.17fF
C31 a_30850_2328# gnd 3.17fF
C32 a_19885_2324# gnd 3.17fF
C33 a_9177_2330# gnd 3.17fF
C34 a_40510_2326# gnd 3.33fF
C35 a_41554_3178# gnd 2.33fF
C36 a_39059_3183# gnd 4.37fF
C37 a_33784_2370# gnd 3.33fF
C38 a_32955_2733# gnd 3.17fF
C39 a_33784_3049# gnd 2.80fF
C40 a_29802_2332# gnd 3.33fF
C41 a_30846_3184# gnd 2.33fF
C42 a_28351_3189# gnd 4.37fF
C43 a_23076_2376# gnd 3.33fF
C44 a_32955_3128# gnd 2.27fF
C45 a_22247_2739# gnd 3.17fF
C46 a_23076_3055# gnd 2.80fF
C47 a_18837_2328# gnd 3.33fF
C48 a_19881_3180# gnd 2.33fF
C49 a_17386_3185# gnd 4.37fF
C50 a_12111_2372# gnd 3.33fF
C51 a_22247_3134# gnd 2.27fF
C52 a_11282_2735# gnd 3.17fF
C53 a_12111_3051# gnd 2.80fF
C54 a_8129_2334# gnd 3.33fF
C55 a_9173_3186# gnd 2.33fF
C56 a_6678_3191# gnd 4.37fF
C57 a_1403_2378# gnd 3.33fF
C58 a_11282_3130# gnd 2.27fF
C59 a_574_2741# gnd 3.17fF
C60 a_1403_3057# gnd 2.80fF
C61 a_574_3136# gnd 2.27fF
C62 a_41558_3001# gnd 3.43fF
C63 a_30850_3007# gnd 3.43fF
C64 a_19885_3003# gnd 3.43fF
C65 a_9177_3009# gnd 3.43fF
C66 a_41554_3946# gnd 2.27fF
C67 a_39063_3006# gnd 3.43fF
C68 a_40506_3950# gnd 2.80fF
C69 a_34832_3045# gnd 3.16fF
C70 a_32955_3384# gnd 3.43fF
C71 a_30846_3952# gnd 2.27fF
C72 a_28355_3012# gnd 3.43fF
C73 a_29798_3956# gnd 2.80fF
C74 a_24124_3051# gnd 3.16fF
C75 a_32955_3925# gnd 2.33fF
C76 a_22247_3390# gnd 3.43fF
C77 a_19881_3948# gnd 2.27fF
C78 a_17390_3008# gnd 3.43fF
C79 a_18833_3952# gnd 2.80fF
C80 a_13159_3047# gnd 3.16fF
C81 a_22247_3931# gnd 2.33fF
C82 a_11282_3386# gnd 3.43fF
C83 a_9173_3954# gnd 2.27fF
C84 a_6682_3014# gnd 3.43fF
C85 a_8125_3958# gnd 2.80fF
C86 a_2451_3053# gnd 3.16fF
C87 a_11282_3927# gnd 2.33fF
C88 a_574_3392# gnd 3.43fF
C89 a_574_3933# gnd 2.33fF
C90 a_41558_3769# gnd 3.17fF
C91 a_30850_3775# gnd 3.17fF
C92 a_19885_3771# gnd 3.17fF
C93 a_9177_3777# gnd 3.17fF
C94 a_40510_3773# gnd 3.33fF
C95 a_41554_4625# gnd 2.33fF
C96 a_39016_4628# gnd 3.27fF
C97 a_32688_217# gnd 10.85fF
C98 a_33784_3817# gnd 3.33fF
C99 a_34832_4492# gnd 3.64fF
C100 a_32955_4180# gnd 3.17fF
C101 a_33784_4496# gnd 2.80fF
C102 a_29802_3779# gnd 3.33fF
C103 a_30846_4631# gnd 2.33fF
C104 a_28308_4634# gnd 3.27fF
C105 a_32955_4575# gnd 2.27fF
C106 a_27026_4504# gnd 11.63fF
C107 a_23076_3823# gnd 3.33fF
C108 a_24124_4498# gnd 3.64fF
C109 a_22247_4186# gnd 3.17fF
C110 a_23076_4502# gnd 2.80fF
C111 a_18837_3775# gnd 3.33fF
C112 a_19881_4627# gnd 2.33fF
C113 a_17343_4630# gnd 3.27fF
C114 a_22247_4581# gnd 2.27fF
C115 a_11015_219# gnd 10.85fF
C116 a_12111_3819# gnd 3.33fF
C117 a_13159_4494# gnd 3.64fF
C118 a_11282_4182# gnd 3.17fF
C119 a_12111_4498# gnd 2.80fF
C120 a_8129_3781# gnd 3.33fF
C121 a_9173_4633# gnd 2.33fF
C122 a_6635_4636# gnd 3.27fF
C123 a_11282_4577# gnd 2.27fF
C124 a_5353_4506# gnd 11.63fF
C125 a_1403_3825# gnd 3.33fF
C126 a_2451_4500# gnd 3.64fF
C127 d5 gnd 84.36fF
C128 a_574_4188# gnd 3.17fF
C129 a_1403_4504# gnd 2.80fF
C130 a_574_4583# gnd 2.27fF
C131 a_41558_4448# gnd 3.52fF
C132 a_30850_4454# gnd 3.52fF
C133 a_19885_4450# gnd 3.52fF
C134 a_9177_4456# gnd 3.52fF
C135 a_41553_5466# gnd 2.27fF
C136 a_40505_5470# gnd 2.80fF
C137 a_36222_5334# gnd 3.19fF
C138 a_32955_4831# gnd 3.52fF
C139 a_30845_5472# gnd 2.27fF
C140 a_29797_5476# gnd 2.80fF
C141 a_25514_5340# gnd 3.19fF
C142 a_32954_5445# gnd 2.33fF
C143 a_22247_4837# gnd 3.52fF
C144 a_19880_5468# gnd 2.27fF
C145 a_18832_5472# gnd 2.80fF
C146 a_14549_5336# gnd 3.19fF
C147 a_22246_5451# gnd 2.33fF
C148 a_11282_4833# gnd 3.52fF
C149 a_9172_5474# gnd 2.27fF
C150 a_8124_5478# gnd 2.80fF
C151 a_3841_5342# gnd 3.19fF
C152 a_11281_5447# gnd 2.33fF
C153 a_574_4839# gnd 3.52fF
C154 a_573_5453# gnd 2.33fF
C155 a_41557_5289# gnd 3.17fF
C156 a_30849_5295# gnd 3.17fF
C157 a_19884_5291# gnd 3.17fF
C158 a_9176_5297# gnd 3.17fF
C159 a_40509_5293# gnd 3.33fF
C160 a_41553_6145# gnd 2.33fF
C161 a_39020_4451# gnd 3.19fF
C162 a_39058_6150# gnd 3.65fF
C163 a_33783_5337# gnd 3.33fF
C164 a_32954_5700# gnd 3.17fF
C165 a_33783_6016# gnd 2.80fF
C166 a_29801_5299# gnd 3.33fF
C167 a_30845_6151# gnd 2.33fF
C168 a_28312_4457# gnd 3.19fF
C169 a_28350_6156# gnd 3.65fF
C170 a_23075_5343# gnd 3.33fF
C171 a_32954_6095# gnd 2.27fF
C172 a_22246_5706# gnd 3.17fF
C173 a_23075_6022# gnd 2.80fF
C174 a_18836_5295# gnd 3.33fF
C175 a_19880_6147# gnd 2.33fF
C176 a_17347_4453# gnd 3.19fF
C177 a_17385_6152# gnd 3.65fF
C178 a_12110_5339# gnd 3.33fF
C179 a_22246_6101# gnd 2.27fF
C180 a_11281_5702# gnd 3.17fF
C181 a_12110_6018# gnd 2.80fF
C182 a_8128_5301# gnd 3.33fF
C183 a_9172_6153# gnd 2.33fF
C184 a_6639_4459# gnd 3.19fF
C185 a_6677_6158# gnd 3.65fF
C186 a_1402_5345# gnd 3.33fF
C187 a_11281_6097# gnd 2.27fF
C188 a_573_5708# gnd 3.17fF
C189 a_1402_6024# gnd 2.80fF
C190 a_573_6103# gnd 2.27fF
C191 a_41557_5968# gnd 3.43fF
C192 a_30849_5974# gnd 3.43fF
C193 a_19884_5970# gnd 3.43fF
C194 a_9176_5976# gnd 3.43fF
C195 a_41553_6913# gnd 2.27fF
C196 a_39062_5973# gnd 3.20fF
C197 a_40505_6917# gnd 2.80fF
C198 a_34831_6012# gnd 3.43fF
C199 a_36227_5453# gnd 3.27fF
C200 a_32954_6351# gnd 3.43fF
C201 a_30845_6919# gnd 2.27fF
C202 a_28354_5979# gnd 3.20fF
C203 a_29797_6923# gnd 2.80fF
C204 a_24123_6018# gnd 3.43fF
C205 a_25519_5459# gnd 3.27fF
C206 a_32954_6892# gnd 2.33fF
C207 a_22246_6357# gnd 3.43fF
C208 a_19880_6915# gnd 2.27fF
C209 a_17389_5975# gnd 3.20fF
C210 a_18832_6919# gnd 2.80fF
C211 a_13158_6014# gnd 3.43fF
C212 a_14554_5455# gnd 3.27fF
C213 a_22246_6898# gnd 2.33fF
C214 a_11281_6353# gnd 3.43fF
C215 a_9172_6921# gnd 2.27fF
C216 a_6681_5981# gnd 3.20fF
C217 a_8124_6925# gnd 2.80fF
C218 a_2450_6020# gnd 3.43fF
C219 a_3846_5461# gnd 3.27fF
C220 a_11281_6894# gnd 2.33fF
C221 a_573_6359# gnd 3.43fF
C222 a_573_6900# gnd 2.33fF
C223 a_41557_6736# gnd 3.17fF
C224 a_30849_6742# gnd 3.17fF
C225 a_19884_6738# gnd 3.17fF
C226 a_9176_6744# gnd 3.17fF
C227 a_40509_6740# gnd 3.33fF
C228 a_41553_7592# gnd 2.33fF
C229 a_37635_4498# gnd 4.30fF
C230 a_37950_7601# gnd 7.03fF
C231 a_33783_6784# gnd 3.33fF
C232 a_34831_7459# gnd 4.35fF
C233 a_32954_7147# gnd 3.17fF
C234 a_33783_7463# gnd 2.80fF
C235 a_29801_6746# gnd 3.33fF
C236 a_30845_7598# gnd 2.33fF
C237 a_26927_4504# gnd 4.30fF
C238 a_27242_7607# gnd 7.03fF
C239 a_23075_6790# gnd 3.33fF
C240 a_24123_7465# gnd 4.35fF
C241 a_32954_7542# gnd 2.27fF
C242 a_22246_7153# gnd 3.17fF
C243 a_23075_7469# gnd 2.80fF
C244 a_18836_6742# gnd 3.33fF
C245 a_19880_7594# gnd 2.33fF
C246 a_15962_4500# gnd 4.30fF
C247 a_16277_7603# gnd 7.03fF
C248 a_12110_6786# gnd 3.33fF
C249 a_13158_7461# gnd 4.35fF
C250 a_22246_7548# gnd 2.27fF
C251 a_11281_7149# gnd 3.17fF
C252 a_12110_7465# gnd 2.80fF
C253 a_8128_6748# gnd 3.33fF
C254 a_9172_7600# gnd 2.33fF
C255 a_5254_4506# gnd 4.30fF
C256 a_5569_7609# gnd 7.03fF
C257 a_1402_6792# gnd 3.33fF
C258 a_2450_7467# gnd 4.35fF
C259 a_11281_7544# gnd 2.27fF
C260 a_573_7155# gnd 3.17fF
C261 a_1402_7471# gnd 2.80fF
C262 a_573_7550# gnd 2.27fF
C263 a_41557_7415# gnd 3.62fF
C264 a_30849_7421# gnd 3.62fF
C265 a_19884_7417# gnd 3.62fF
C266 a_9176_7423# gnd 3.62fF
C267 a_41556_8507# gnd 2.27fF
C268 a_40508_8511# gnd 2.80fF
C269 a_36321_5334# gnd 4.97fF
C270 a_37389_8369# gnd 4.72fF
C271 a_32954_7798# gnd 3.62fF
C272 a_30848_8513# gnd 2.27fF
C273 a_29800_8517# gnd 2.80fF
C274 a_25613_5340# gnd 4.97fF
C275 a_26681_8375# gnd 4.72fF
C276 a_32957_8486# gnd 2.33fF
C277 a_22246_7804# gnd 3.62fF
C278 a_19883_8509# gnd 2.27fF
C279 a_18835_8513# gnd 2.80fF
C280 a_14648_5336# gnd 4.97fF
C281 a_15716_8371# gnd 4.72fF
C282 a_22249_8492# gnd 2.33fF
C283 a_11281_7800# gnd 3.62fF
C284 a_9175_8515# gnd 2.27fF
C285 a_8127_8519# gnd 2.80fF
C286 a_3940_5342# gnd 4.97fF
C287 a_5008_8377# gnd 4.72fF
C288 a_11284_8488# gnd 2.33fF
C289 d4 gnd 107.15fF
C290 a_573_7806# gnd 3.62fF
C291 a_576_8494# gnd 2.33fF
C292 a_41560_8330# gnd 3.17fF
C293 a_30852_8336# gnd 3.17fF
C294 a_19887_8332# gnd 3.17fF
C295 a_9179_8338# gnd 3.17fF
C296 a_40512_8334# gnd 3.33fF
C297 a_41556_9186# gnd 2.33fF
C298 a_39061_9191# gnd 4.35fF
C299 a_33786_8378# gnd 3.33fF
C300 a_32957_8741# gnd 3.17fF
C301 a_33786_9057# gnd 2.80fF
C302 a_29804_8340# gnd 3.33fF
C303 a_30848_9192# gnd 2.33fF
C304 a_28353_9197# gnd 4.35fF
C305 a_23078_8384# gnd 3.33fF
C306 a_32957_9136# gnd 2.27fF
C307 a_22249_8747# gnd 3.17fF
C308 a_23078_9063# gnd 2.80fF
C309 a_18839_8336# gnd 3.33fF
C310 a_19883_9188# gnd 2.33fF
C311 a_17388_9193# gnd 4.35fF
C312 a_12113_8380# gnd 3.33fF
C313 a_22249_9142# gnd 2.27fF
C314 a_11284_8743# gnd 3.17fF
C315 a_12113_9059# gnd 2.80fF
C316 a_8131_8342# gnd 3.33fF
C317 a_9175_9194# gnd 2.33fF
C318 a_6680_9199# gnd 4.35fF
C319 a_1405_8386# gnd 3.33fF
C320 a_11284_9138# gnd 2.27fF
C321 a_576_8749# gnd 3.17fF
C322 a_1405_9065# gnd 2.80fF
C323 a_576_9144# gnd 2.27fF
C324 a_41560_9009# gnd 3.43fF
C325 a_30852_9015# gnd 3.43fF
C326 a_19887_9011# gnd 3.43fF
C327 a_9179_9017# gnd 3.43fF
C328 a_41556_9954# gnd 2.27fF
C329 a_39065_9014# gnd 3.43fF
C330 a_40508_9958# gnd 2.80fF
C331 a_34834_9053# gnd 3.20fF
C332 a_32957_9392# gnd 3.43fF
C333 a_30848_9960# gnd 2.27fF
C334 a_28357_9020# gnd 3.43fF
C335 a_29800_9964# gnd 2.80fF
C336 a_24126_9059# gnd 3.20fF
C337 a_32957_9933# gnd 2.33fF
C338 a_22249_9398# gnd 3.43fF
C339 a_19883_9956# gnd 2.27fF
C340 a_17392_9016# gnd 3.43fF
C341 a_18835_9960# gnd 2.80fF
C342 a_13161_9055# gnd 3.20fF
C343 a_22249_9939# gnd 2.33fF
C344 a_11284_9394# gnd 3.43fF
C345 a_9175_9962# gnd 2.27fF
C346 a_6684_9022# gnd 3.43fF
C347 a_8127_9966# gnd 2.80fF
C348 a_2453_9061# gnd 3.20fF
C349 a_11284_9935# gnd 2.33fF
C350 a_576_9400# gnd 3.43fF
C351 a_576_9941# gnd 2.33fF
C352 a_41560_9777# gnd 3.17fF
C353 a_30852_9783# gnd 3.17fF
C354 a_19887_9779# gnd 3.17fF
C355 a_9179_9785# gnd 3.17fF
C356 a_40512_9781# gnd 3.33fF
C357 a_41556_10633# gnd 2.33fF
C358 a_37954_7424# gnd 4.90fF
C359 a_39018_10636# gnd 3.27fF
C360 a_33786_9825# gnd 3.33fF
C361 a_34834_10500# gnd 3.65fF
C362 a_32957_10188# gnd 3.17fF
C363 a_33786_10504# gnd 2.80fF
C364 a_29804_9787# gnd 3.33fF
C365 a_30848_10639# gnd 2.33fF
C366 a_27246_7430# gnd 4.90fF
C367 a_28310_10642# gnd 3.27fF
C368 a_23078_9831# gnd 3.33fF
C369 a_24126_10506# gnd 3.65fF
C370 a_32957_10583# gnd 2.27fF
C371 a_22249_10194# gnd 3.17fF
C372 a_23078_10510# gnd 2.80fF
C373 a_18839_9783# gnd 3.33fF
C374 a_19883_10635# gnd 2.33fF
C375 a_16281_7426# gnd 4.90fF
C376 a_17345_10638# gnd 3.27fF
C377 a_12113_9827# gnd 3.33fF
C378 a_13161_10502# gnd 3.65fF
C379 a_22249_10589# gnd 2.27fF
C380 a_11284_10190# gnd 3.17fF
C381 a_12113_10506# gnd 2.80fF
C382 a_8131_9789# gnd 3.33fF
C383 a_9175_10641# gnd 2.33fF
C384 a_5573_7432# gnd 4.90fF
C385 a_6637_10644# gnd 3.27fF
C386 a_1405_9833# gnd 3.33fF
C387 a_2453_10508# gnd 3.65fF
C388 a_11284_10585# gnd 2.27fF
C389 a_576_10196# gnd 3.17fF
C390 a_1405_10512# gnd 2.80fF
C391 a_576_10591# gnd 2.27fF
C392 a_41560_10456# gnd 3.52fF
C393 a_30852_10462# gnd 3.52fF
C394 a_19887_10458# gnd 3.52fF
C395 a_9179_10464# gnd 3.52fF
C396 a_41555_11474# gnd 2.27fF
C397 a_40507_11478# gnd 2.80fF
C398 a_36224_11342# gnd 3.19fF
C399 a_36323_11342# gnd 7.02fF
C400 a_32957_10839# gnd 3.52fF
C401 a_30847_11480# gnd 2.27fF
C402 a_29799_11484# gnd 2.80fF
C403 a_25516_11348# gnd 3.19fF
C404 a_25615_11348# gnd 7.02fF
C405 a_32956_11453# gnd 2.33fF
C406 a_22249_10845# gnd 3.52fF
C407 a_19882_11476# gnd 2.27fF
C408 a_18834_11480# gnd 2.80fF
C409 a_14551_11344# gnd 3.19fF
C410 a_14650_11344# gnd 7.02fF
C411 a_22248_11459# gnd 2.33fF
C412 a_11284_10841# gnd 3.52fF
C413 a_9174_11482# gnd 2.27fF
C414 a_8126_11486# gnd 2.80fF
C415 a_3843_11350# gnd 3.19fF
C416 a_3942_11350# gnd 7.02fF
C417 a_11283_11455# gnd 2.33fF
C418 d3 gnd 207.02fF
C419 a_576_10847# gnd 3.52fF
C420 a_575_11461# gnd 2.33fF
C421 a_41559_11297# gnd 3.17fF
C422 a_30851_11303# gnd 3.17fF
C423 a_19886_11299# gnd 3.17fF
C424 a_9178_11305# gnd 3.17fF
C425 a_40511_11301# gnd 3.33fF
C426 a_41555_12153# gnd 2.33fF
C427 a_39022_10459# gnd 3.19fF
C428 a_39060_12158# gnd 3.73fF
C429 a_33785_11345# gnd 3.33fF
C430 a_32956_11708# gnd 3.17fF
C431 a_33785_12024# gnd 2.80fF
C432 a_29803_11307# gnd 3.33fF
C433 a_30847_12159# gnd 2.33fF
C434 a_28314_10465# gnd 3.19fF
C435 a_28352_12164# gnd 3.73fF
C436 a_23077_11351# gnd 3.33fF
C437 a_32956_12103# gnd 2.27fF
C438 a_22248_11714# gnd 3.17fF
C439 a_23077_12030# gnd 2.80fF
C440 a_18838_11303# gnd 3.33fF
C441 a_19882_12155# gnd 2.33fF
C442 a_17349_10461# gnd 3.19fF
C443 a_17387_12160# gnd 3.73fF
C444 a_12112_11347# gnd 3.33fF
C445 a_22248_12109# gnd 2.27fF
C446 a_11283_11710# gnd 3.17fF
C447 a_12112_12026# gnd 2.80fF
C448 a_8130_11309# gnd 3.33fF
C449 a_9174_12161# gnd 2.33fF
C450 a_6641_10467# gnd 3.19fF
C451 a_6679_12166# gnd 3.73fF
C452 a_1404_11353# gnd 3.33fF
C453 a_11283_12105# gnd 2.27fF
C454 a_575_11716# gnd 3.17fF
C455 a_1404_12032# gnd 2.80fF
C456 a_575_12111# gnd 2.27fF
C457 a_41559_11976# gnd 3.43fF
C458 a_30851_11982# gnd 3.43fF
C459 a_19886_11978# gnd 3.43fF
C460 a_9178_11984# gnd 3.43fF
C461 a_41555_12921# gnd 2.27fF
C462 a_39064_11981# gnd 3.35fF
C463 a_40507_12925# gnd 2.80fF
C464 a_34833_12020# gnd 3.43fF
C465 a_36229_11461# gnd 3.27fF
C466 a_32956_12359# gnd 3.43fF
C467 a_30847_12927# gnd 2.27fF
C468 a_28356_11987# gnd 3.35fF
C469 a_29799_12931# gnd 2.80fF
C470 a_24125_12026# gnd 3.43fF
C471 a_25521_11467# gnd 3.27fF
C472 a_32956_12900# gnd 2.33fF
C473 a_22248_12365# gnd 3.43fF
C474 a_19882_12923# gnd 2.27fF
C475 a_17391_11983# gnd 3.35fF
C476 a_18834_12927# gnd 2.80fF
C477 a_13160_12022# gnd 3.43fF
C478 a_14556_11463# gnd 3.27fF
C479 a_22248_12906# gnd 2.33fF
C480 a_11283_12361# gnd 3.43fF
C481 a_9174_12929# gnd 2.27fF
C482 a_6683_11989# gnd 3.35fF
C483 a_8126_12933# gnd 2.80fF
C484 a_2452_12028# gnd 3.43fF
C485 a_3848_11469# gnd 3.27fF
C486 a_11283_12902# gnd 2.33fF
C487 d2 gnd 211.93fF
C488 a_575_12367# gnd 3.43fF
C489 a_575_12908# gnd 2.33fF
C490 a_41559_12744# gnd 3.17fF
C491 a_30851_12750# gnd 3.17fF
C492 a_19886_12746# gnd 3.17fF
C493 a_9178_12752# gnd 3.17fF
C494 a_40511_12748# gnd 3.40fF
C495 a_41555_13600# gnd 2.73fF
C496 a_33785_12792# gnd 3.33fF
C497 a_34833_13467# gnd 4.35fF
C498 a_32956_13155# gnd 3.17fF
C499 a_33785_13471# gnd 2.80fF
C500 a_29803_12754# gnd 3.33fF
C501 a_30847_13606# gnd 2.33fF
C502 a_23077_12798# gnd 3.33fF
C503 a_24125_13473# gnd 4.35fF
C504 a_32956_13550# gnd 2.27fF
C505 a_22248_13161# gnd 3.17fF
C506 a_23077_13477# gnd 2.80fF
C507 a_18838_12750# gnd 3.33fF
C508 a_19882_13602# gnd 2.33fF
C509 a_12112_12794# gnd 3.33fF
C510 a_13160_13469# gnd 4.35fF
C511 a_22248_13556# gnd 2.27fF
C512 a_11283_13157# gnd 3.17fF
C513 a_12112_13473# gnd 2.80fF
C514 a_8130_12756# gnd 3.33fF
C515 a_9174_13608# gnd 2.33fF
C516 a_1404_12800# gnd 3.33fF
C517 a_2452_13475# gnd 4.35fF
C518 a_11283_13552# gnd 2.27fF
C519 d1 gnd 247.46fF
C520 a_575_13163# gnd 3.17fF
C521 a_1404_13479# gnd 2.80fF
C522 d0 gnd 307.27fF
C523 a_575_13558# gnd 2.27fF
C524 a_30851_13429# gnd 4.89fF
C525 a_19886_13425# gnd 5.08fF
C526 a_9178_13431# gnd 4.89fF
C527 vdd gnd 1304.67fF
