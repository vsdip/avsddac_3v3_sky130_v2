magic
tech sky130A
timestamp 1633145158
<< nwell >>
rect 41 201 852 425
<< nmos >>
rect 105 100 155 142
rect 318 100 368 142
rect 526 100 576 142
rect 734 100 784 142
<< pmos >>
rect 105 219 155 319
rect 318 219 368 319
rect 526 219 576 319
rect 734 219 784 319
<< ndiff >>
rect 56 132 105 142
rect 56 112 67 132
rect 87 112 105 132
rect 56 100 105 112
rect 155 136 199 142
rect 155 116 170 136
rect 190 116 199 136
rect 155 100 199 116
rect 269 132 318 142
rect 269 112 280 132
rect 300 112 318 132
rect 269 100 318 112
rect 368 136 412 142
rect 368 116 383 136
rect 403 116 412 136
rect 368 100 412 116
rect 477 132 526 142
rect 477 112 488 132
rect 508 112 526 132
rect 477 100 526 112
rect 576 136 620 142
rect 576 116 591 136
rect 611 116 620 136
rect 576 100 620 116
rect 690 136 734 142
rect 690 116 699 136
rect 719 116 734 136
rect 690 100 734 116
rect 784 132 833 142
rect 784 112 802 132
rect 822 112 833 132
rect 784 100 833 112
<< pdiff >>
rect 61 281 105 319
rect 61 261 73 281
rect 93 261 105 281
rect 61 219 105 261
rect 155 281 197 319
rect 155 261 169 281
rect 189 261 197 281
rect 155 219 197 261
rect 274 281 318 319
rect 274 261 286 281
rect 306 261 318 281
rect 274 219 318 261
rect 368 281 410 319
rect 368 261 382 281
rect 402 261 410 281
rect 368 219 410 261
rect 482 281 526 319
rect 482 261 494 281
rect 514 261 526 281
rect 482 219 526 261
rect 576 281 618 319
rect 576 261 590 281
rect 610 261 618 281
rect 576 219 618 261
rect 692 281 734 319
rect 692 261 700 281
rect 720 261 734 281
rect 692 219 734 261
rect 784 288 829 319
rect 784 281 828 288
rect 784 261 796 281
rect 816 261 828 281
rect 784 219 828 261
<< ndiffc >>
rect 67 112 87 132
rect 170 116 190 136
rect 280 112 300 132
rect 383 116 403 136
rect 488 112 508 132
rect 591 116 611 136
rect 699 116 719 136
rect 802 112 822 132
<< pdiffc >>
rect 73 261 93 281
rect 169 261 189 281
rect 286 261 306 281
rect 382 261 402 281
rect 494 261 514 281
rect 590 261 610 281
rect 700 261 720 281
rect 796 261 816 281
<< psubdiff >>
rect 141 45 252 59
rect 141 15 182 45
rect 210 15 252 45
rect 141 0 252 15
<< nsubdiff >>
rect 142 392 252 406
rect 142 362 185 392
rect 213 362 252 392
rect 142 347 252 362
<< psubdiffcont >>
rect 182 15 210 45
<< nsubdiffcont >>
rect 185 362 213 392
<< poly >>
rect 105 319 155 332
rect 318 319 368 332
rect 526 319 576 332
rect 734 319 784 332
rect 105 191 155 219
rect 105 171 118 191
rect 138 171 155 191
rect 105 142 155 171
rect 318 190 368 219
rect 318 166 329 190
rect 353 166 368 190
rect 318 142 368 166
rect 526 195 576 219
rect 526 171 538 195
rect 562 171 576 195
rect 526 142 576 171
rect 734 193 784 219
rect 734 167 752 193
rect 778 167 784 193
rect 734 142 784 167
rect 105 84 155 100
rect 318 84 368 100
rect 526 84 576 100
rect 734 84 784 100
<< polycont >>
rect 118 171 138 191
rect 329 166 353 190
rect 538 171 562 195
rect 752 167 778 193
<< locali >>
rect 485 429 878 449
rect 898 429 901 449
rect 485 424 901 429
rect 485 423 826 424
rect 142 392 252 406
rect 142 389 185 392
rect 142 384 146 389
rect 64 362 146 384
rect 175 362 185 389
rect 213 365 220 392
rect 249 384 252 392
rect 249 365 314 384
rect 213 362 314 365
rect 64 360 314 362
rect 64 281 101 360
rect 142 347 252 360
rect 216 291 247 292
rect 64 261 73 281
rect 93 261 101 281
rect 64 251 101 261
rect 160 281 247 291
rect 160 261 169 281
rect 189 261 247 281
rect 160 252 247 261
rect 160 251 197 252
rect 216 199 247 252
rect 277 281 314 360
rect 429 291 460 292
rect 277 261 286 281
rect 306 261 314 281
rect 277 251 314 261
rect 373 284 460 291
rect 373 281 434 284
rect 373 261 382 281
rect 402 264 434 281
rect 455 264 460 284
rect 402 261 460 264
rect 373 254 460 261
rect 485 281 522 423
rect 788 422 825 423
rect 637 291 673 292
rect 485 261 494 281
rect 514 261 522 281
rect 373 252 429 254
rect 373 251 410 252
rect 485 251 522 261
rect 581 281 729 291
rect 829 288 925 290
rect 581 261 590 281
rect 610 261 700 281
rect 720 261 729 281
rect 581 255 729 261
rect 581 252 645 255
rect 581 251 618 252
rect 637 225 645 252
rect 666 252 729 255
rect 787 281 925 288
rect 787 261 796 281
rect 816 261 925 281
rect 787 252 925 261
rect 666 225 673 252
rect 692 251 729 252
rect 788 251 825 252
rect 637 200 673 225
rect 108 198 149 199
rect 0 191 149 198
rect 0 171 118 191
rect 138 171 149 191
rect 0 163 149 171
rect 216 195 575 199
rect 216 190 538 195
rect 216 166 329 190
rect 353 171 538 190
rect 562 171 575 195
rect 353 166 575 171
rect 216 163 575 166
rect 637 163 672 200
rect 740 197 840 200
rect 740 193 807 197
rect 740 167 752 193
rect 778 171 807 193
rect 833 171 840 197
rect 778 167 840 171
rect 740 163 840 167
rect 216 142 247 163
rect 637 142 673 163
rect 59 141 96 142
rect 58 132 96 141
rect 58 112 67 132
rect 87 112 96 132
rect 58 104 96 112
rect 162 136 247 142
rect 272 141 309 142
rect 162 116 170 136
rect 190 116 247 136
rect 162 108 247 116
rect 271 132 309 141
rect 271 112 280 132
rect 300 112 309 132
rect 162 107 198 108
rect 271 104 309 112
rect 375 136 460 142
rect 480 141 517 142
rect 375 116 383 136
rect 403 135 460 136
rect 403 116 432 135
rect 375 115 432 116
rect 453 115 460 135
rect 375 108 460 115
rect 479 132 517 141
rect 479 112 488 132
rect 508 112 517 132
rect 375 107 411 108
rect 479 104 517 112
rect 583 136 727 142
rect 583 116 591 136
rect 611 116 699 136
rect 719 116 727 136
rect 583 108 727 116
rect 583 107 619 108
rect 691 107 727 108
rect 793 141 830 142
rect 793 140 831 141
rect 793 132 857 140
rect 793 112 802 132
rect 822 118 857 132
rect 877 118 880 138
rect 822 113 880 118
rect 822 112 857 113
rect 59 75 96 104
rect 60 73 96 75
rect 272 73 309 104
rect 60 51 309 73
rect 141 45 252 51
rect 141 37 182 45
rect 141 17 149 37
rect 168 17 182 37
rect 141 15 182 17
rect 210 37 252 45
rect 210 17 226 37
rect 245 17 252 37
rect 210 15 252 17
rect 141 0 252 15
rect 480 -17 517 104
rect 793 100 857 112
rect 897 -15 924 252
rect 756 -17 924 -15
rect 480 -43 924 -17
rect 756 -44 924 -43
<< viali >>
rect 878 429 898 449
rect 146 362 175 389
rect 220 365 249 392
rect 434 264 455 284
rect 645 225 666 255
rect 807 171 833 197
rect 432 115 453 135
rect 857 118 877 138
rect 149 17 168 37
rect 226 17 245 37
<< metal1 >>
rect 49 393 252 406
rect 49 360 73 393
rect 109 392 252 393
rect 109 389 220 392
rect 109 362 146 389
rect 175 365 220 389
rect 249 365 252 392
rect 175 362 252 365
rect 109 360 252 362
rect 49 347 252 360
rect 49 346 150 347
rect 427 284 459 291
rect 427 264 434 284
rect 455 264 459 284
rect 427 199 459 264
rect 639 255 670 481
rect 874 454 906 455
rect 871 449 906 454
rect 871 429 878 449
rect 898 429 906 449
rect 871 421 906 429
rect 639 225 645 255
rect 666 225 670 255
rect 639 217 670 225
rect 797 199 837 200
rect 427 197 839 199
rect 427 171 807 197
rect 833 171 839 197
rect 427 163 839 171
rect 427 135 459 163
rect 872 143 906 421
rect 427 115 432 135
rect 453 115 459 135
rect 427 108 459 115
rect 850 138 906 143
rect 850 118 857 138
rect 877 118 906 138
rect 850 111 906 118
rect 850 110 885 111
rect 141 37 252 59
rect 141 17 149 37
rect 168 17 226 37
rect 245 17 252 37
rect 141 0 252 17
<< via1 >>
rect 73 360 109 393
<< metal2 >>
rect 50 393 136 406
rect 50 360 73 393
rect 109 360 136 393
rect 50 348 136 360
<< end >>
