magic
tech sky130A
timestamp 1620560744
<< nwell >>
rect 318 982 645 1056
rect 318 832 1129 982
rect 1256 738 1583 812
rect 1256 588 2067 738
rect 317 428 644 502
rect 317 278 1128 428
rect 1397 146 1724 220
rect 1397 -4 2208 146
rect 319 -121 646 -47
rect 319 -271 1130 -121
rect 1257 -365 1584 -291
rect 1257 -515 2068 -365
rect 318 -675 645 -601
rect 318 -825 1129 -675
<< nmos >>
rect 382 731 432 773
rect 595 731 645 773
rect 803 731 853 773
rect 1011 731 1061 773
rect 1320 487 1370 529
rect 1533 487 1583 529
rect 1741 487 1791 529
rect 1949 487 1999 529
rect 381 177 431 219
rect 594 177 644 219
rect 802 177 852 219
rect 1010 177 1060 219
rect 1461 -105 1511 -63
rect 1674 -105 1724 -63
rect 1882 -105 1932 -63
rect 2090 -105 2140 -63
rect 383 -372 433 -330
rect 596 -372 646 -330
rect 804 -372 854 -330
rect 1012 -372 1062 -330
rect 1321 -616 1371 -574
rect 1534 -616 1584 -574
rect 1742 -616 1792 -574
rect 1950 -616 2000 -574
rect 382 -926 432 -884
rect 595 -926 645 -884
rect 803 -926 853 -884
rect 1011 -926 1061 -884
<< pmos >>
rect 382 850 432 950
rect 595 850 645 950
rect 803 850 853 950
rect 1011 850 1061 950
rect 1320 606 1370 706
rect 1533 606 1583 706
rect 1741 606 1791 706
rect 1949 606 1999 706
rect 381 296 431 396
rect 594 296 644 396
rect 802 296 852 396
rect 1010 296 1060 396
rect 1461 14 1511 114
rect 1674 14 1724 114
rect 1882 14 1932 114
rect 2090 14 2140 114
rect 383 -253 433 -153
rect 596 -253 646 -153
rect 804 -253 854 -153
rect 1012 -253 1062 -153
rect 1321 -497 1371 -397
rect 1534 -497 1584 -397
rect 1742 -497 1792 -397
rect 1950 -497 2000 -397
rect 382 -807 432 -707
rect 595 -807 645 -707
rect 803 -807 853 -707
rect 1011 -807 1061 -707
<< ndiff >>
rect 333 763 382 773
rect 333 743 344 763
rect 364 743 382 763
rect 333 731 382 743
rect 432 767 476 773
rect 432 747 447 767
rect 467 747 476 767
rect 432 731 476 747
rect 546 763 595 773
rect 546 743 557 763
rect 577 743 595 763
rect 546 731 595 743
rect 645 767 689 773
rect 645 747 660 767
rect 680 747 689 767
rect 645 731 689 747
rect 754 763 803 773
rect 754 743 765 763
rect 785 743 803 763
rect 754 731 803 743
rect 853 767 897 773
rect 853 747 868 767
rect 888 747 897 767
rect 853 731 897 747
rect 967 767 1011 773
rect 967 747 976 767
rect 996 747 1011 767
rect 967 731 1011 747
rect 1061 763 1110 773
rect 1061 743 1079 763
rect 1099 743 1110 763
rect 1061 731 1110 743
rect 1271 519 1320 529
rect 1271 499 1282 519
rect 1302 499 1320 519
rect 1271 487 1320 499
rect 1370 523 1414 529
rect 1370 503 1385 523
rect 1405 503 1414 523
rect 1370 487 1414 503
rect 1484 519 1533 529
rect 1484 499 1495 519
rect 1515 499 1533 519
rect 1484 487 1533 499
rect 1583 523 1627 529
rect 1583 503 1598 523
rect 1618 503 1627 523
rect 1583 487 1627 503
rect 1692 519 1741 529
rect 1692 499 1703 519
rect 1723 499 1741 519
rect 1692 487 1741 499
rect 1791 523 1835 529
rect 1791 503 1806 523
rect 1826 503 1835 523
rect 1791 487 1835 503
rect 1905 523 1949 529
rect 1905 503 1914 523
rect 1934 503 1949 523
rect 1905 487 1949 503
rect 1999 519 2048 529
rect 1999 499 2017 519
rect 2037 499 2048 519
rect 1999 487 2048 499
rect 332 209 381 219
rect 332 189 343 209
rect 363 189 381 209
rect 332 177 381 189
rect 431 213 475 219
rect 431 193 446 213
rect 466 193 475 213
rect 431 177 475 193
rect 545 209 594 219
rect 545 189 556 209
rect 576 189 594 209
rect 545 177 594 189
rect 644 213 688 219
rect 644 193 659 213
rect 679 193 688 213
rect 644 177 688 193
rect 753 209 802 219
rect 753 189 764 209
rect 784 189 802 209
rect 753 177 802 189
rect 852 213 896 219
rect 852 193 867 213
rect 887 193 896 213
rect 852 177 896 193
rect 966 213 1010 219
rect 966 193 975 213
rect 995 193 1010 213
rect 966 177 1010 193
rect 1060 209 1109 219
rect 1060 189 1078 209
rect 1098 189 1109 209
rect 1060 177 1109 189
rect 1412 -73 1461 -63
rect 1412 -93 1423 -73
rect 1443 -93 1461 -73
rect 1412 -105 1461 -93
rect 1511 -69 1555 -63
rect 1511 -89 1526 -69
rect 1546 -89 1555 -69
rect 1511 -105 1555 -89
rect 1625 -73 1674 -63
rect 1625 -93 1636 -73
rect 1656 -93 1674 -73
rect 1625 -105 1674 -93
rect 1724 -69 1768 -63
rect 1724 -89 1739 -69
rect 1759 -89 1768 -69
rect 1724 -105 1768 -89
rect 1833 -73 1882 -63
rect 1833 -93 1844 -73
rect 1864 -93 1882 -73
rect 1833 -105 1882 -93
rect 1932 -69 1976 -63
rect 1932 -89 1947 -69
rect 1967 -89 1976 -69
rect 1932 -105 1976 -89
rect 2046 -69 2090 -63
rect 2046 -89 2055 -69
rect 2075 -89 2090 -69
rect 2046 -105 2090 -89
rect 2140 -73 2189 -63
rect 2140 -93 2158 -73
rect 2178 -93 2189 -73
rect 2140 -105 2189 -93
rect 334 -340 383 -330
rect 334 -360 345 -340
rect 365 -360 383 -340
rect 334 -372 383 -360
rect 433 -336 477 -330
rect 433 -356 448 -336
rect 468 -356 477 -336
rect 433 -372 477 -356
rect 547 -340 596 -330
rect 547 -360 558 -340
rect 578 -360 596 -340
rect 547 -372 596 -360
rect 646 -336 690 -330
rect 646 -356 661 -336
rect 681 -356 690 -336
rect 646 -372 690 -356
rect 755 -340 804 -330
rect 755 -360 766 -340
rect 786 -360 804 -340
rect 755 -372 804 -360
rect 854 -336 898 -330
rect 854 -356 869 -336
rect 889 -356 898 -336
rect 854 -372 898 -356
rect 968 -336 1012 -330
rect 968 -356 977 -336
rect 997 -356 1012 -336
rect 968 -372 1012 -356
rect 1062 -340 1111 -330
rect 1062 -360 1080 -340
rect 1100 -360 1111 -340
rect 1062 -372 1111 -360
rect 1272 -584 1321 -574
rect 1272 -604 1283 -584
rect 1303 -604 1321 -584
rect 1272 -616 1321 -604
rect 1371 -580 1415 -574
rect 1371 -600 1386 -580
rect 1406 -600 1415 -580
rect 1371 -616 1415 -600
rect 1485 -584 1534 -574
rect 1485 -604 1496 -584
rect 1516 -604 1534 -584
rect 1485 -616 1534 -604
rect 1584 -580 1628 -574
rect 1584 -600 1599 -580
rect 1619 -600 1628 -580
rect 1584 -616 1628 -600
rect 1693 -584 1742 -574
rect 1693 -604 1704 -584
rect 1724 -604 1742 -584
rect 1693 -616 1742 -604
rect 1792 -580 1836 -574
rect 1792 -600 1807 -580
rect 1827 -600 1836 -580
rect 1792 -616 1836 -600
rect 1906 -580 1950 -574
rect 1906 -600 1915 -580
rect 1935 -600 1950 -580
rect 1906 -616 1950 -600
rect 2000 -584 2049 -574
rect 2000 -604 2018 -584
rect 2038 -604 2049 -584
rect 2000 -616 2049 -604
rect 333 -894 382 -884
rect 333 -914 344 -894
rect 364 -914 382 -894
rect 333 -926 382 -914
rect 432 -890 476 -884
rect 432 -910 447 -890
rect 467 -910 476 -890
rect 432 -926 476 -910
rect 546 -894 595 -884
rect 546 -914 557 -894
rect 577 -914 595 -894
rect 546 -926 595 -914
rect 645 -890 689 -884
rect 645 -910 660 -890
rect 680 -910 689 -890
rect 645 -926 689 -910
rect 754 -894 803 -884
rect 754 -914 765 -894
rect 785 -914 803 -894
rect 754 -926 803 -914
rect 853 -890 897 -884
rect 853 -910 868 -890
rect 888 -910 897 -890
rect 853 -926 897 -910
rect 967 -890 1011 -884
rect 967 -910 976 -890
rect 996 -910 1011 -890
rect 967 -926 1011 -910
rect 1061 -894 1110 -884
rect 1061 -914 1079 -894
rect 1099 -914 1110 -894
rect 1061 -926 1110 -914
<< pdiff >>
rect 338 912 382 950
rect 338 892 350 912
rect 370 892 382 912
rect 338 850 382 892
rect 432 912 474 950
rect 432 892 446 912
rect 466 892 474 912
rect 432 850 474 892
rect 551 912 595 950
rect 551 892 563 912
rect 583 892 595 912
rect 551 850 595 892
rect 645 912 687 950
rect 645 892 659 912
rect 679 892 687 912
rect 645 850 687 892
rect 759 912 803 950
rect 759 892 771 912
rect 791 892 803 912
rect 759 850 803 892
rect 853 912 895 950
rect 853 892 867 912
rect 887 892 895 912
rect 853 850 895 892
rect 969 912 1011 950
rect 969 892 977 912
rect 997 892 1011 912
rect 969 850 1011 892
rect 1061 919 1106 950
rect 1061 912 1105 919
rect 1061 892 1073 912
rect 1093 892 1105 912
rect 1061 850 1105 892
rect 1276 668 1320 706
rect 1276 648 1288 668
rect 1308 648 1320 668
rect 1276 606 1320 648
rect 1370 668 1412 706
rect 1370 648 1384 668
rect 1404 648 1412 668
rect 1370 606 1412 648
rect 1489 668 1533 706
rect 1489 648 1501 668
rect 1521 648 1533 668
rect 1489 606 1533 648
rect 1583 668 1625 706
rect 1583 648 1597 668
rect 1617 648 1625 668
rect 1583 606 1625 648
rect 1697 668 1741 706
rect 1697 648 1709 668
rect 1729 648 1741 668
rect 1697 606 1741 648
rect 1791 668 1833 706
rect 1791 648 1805 668
rect 1825 648 1833 668
rect 1791 606 1833 648
rect 1907 668 1949 706
rect 1907 648 1915 668
rect 1935 648 1949 668
rect 1907 606 1949 648
rect 1999 675 2044 706
rect 1999 668 2043 675
rect 1999 648 2011 668
rect 2031 648 2043 668
rect 1999 606 2043 648
rect 337 358 381 396
rect 337 338 349 358
rect 369 338 381 358
rect 337 296 381 338
rect 431 358 473 396
rect 431 338 445 358
rect 465 338 473 358
rect 431 296 473 338
rect 550 358 594 396
rect 550 338 562 358
rect 582 338 594 358
rect 550 296 594 338
rect 644 358 686 396
rect 644 338 658 358
rect 678 338 686 358
rect 644 296 686 338
rect 758 358 802 396
rect 758 338 770 358
rect 790 338 802 358
rect 758 296 802 338
rect 852 358 894 396
rect 852 338 866 358
rect 886 338 894 358
rect 852 296 894 338
rect 968 358 1010 396
rect 968 338 976 358
rect 996 338 1010 358
rect 968 296 1010 338
rect 1060 365 1105 396
rect 1060 358 1104 365
rect 1060 338 1072 358
rect 1092 338 1104 358
rect 1060 296 1104 338
rect 1417 76 1461 114
rect 1417 56 1429 76
rect 1449 56 1461 76
rect 1417 14 1461 56
rect 1511 76 1553 114
rect 1511 56 1525 76
rect 1545 56 1553 76
rect 1511 14 1553 56
rect 1630 76 1674 114
rect 1630 56 1642 76
rect 1662 56 1674 76
rect 1630 14 1674 56
rect 1724 76 1766 114
rect 1724 56 1738 76
rect 1758 56 1766 76
rect 1724 14 1766 56
rect 1838 76 1882 114
rect 1838 56 1850 76
rect 1870 56 1882 76
rect 1838 14 1882 56
rect 1932 76 1974 114
rect 1932 56 1946 76
rect 1966 56 1974 76
rect 1932 14 1974 56
rect 2048 76 2090 114
rect 2048 56 2056 76
rect 2076 56 2090 76
rect 2048 14 2090 56
rect 2140 83 2185 114
rect 2140 76 2184 83
rect 2140 56 2152 76
rect 2172 56 2184 76
rect 2140 14 2184 56
rect 339 -191 383 -153
rect 339 -211 351 -191
rect 371 -211 383 -191
rect 339 -253 383 -211
rect 433 -191 475 -153
rect 433 -211 447 -191
rect 467 -211 475 -191
rect 433 -253 475 -211
rect 552 -191 596 -153
rect 552 -211 564 -191
rect 584 -211 596 -191
rect 552 -253 596 -211
rect 646 -191 688 -153
rect 646 -211 660 -191
rect 680 -211 688 -191
rect 646 -253 688 -211
rect 760 -191 804 -153
rect 760 -211 772 -191
rect 792 -211 804 -191
rect 760 -253 804 -211
rect 854 -191 896 -153
rect 854 -211 868 -191
rect 888 -211 896 -191
rect 854 -253 896 -211
rect 970 -191 1012 -153
rect 970 -211 978 -191
rect 998 -211 1012 -191
rect 970 -253 1012 -211
rect 1062 -184 1107 -153
rect 1062 -191 1106 -184
rect 1062 -211 1074 -191
rect 1094 -211 1106 -191
rect 1062 -253 1106 -211
rect 1277 -435 1321 -397
rect 1277 -455 1289 -435
rect 1309 -455 1321 -435
rect 1277 -497 1321 -455
rect 1371 -435 1413 -397
rect 1371 -455 1385 -435
rect 1405 -455 1413 -435
rect 1371 -497 1413 -455
rect 1490 -435 1534 -397
rect 1490 -455 1502 -435
rect 1522 -455 1534 -435
rect 1490 -497 1534 -455
rect 1584 -435 1626 -397
rect 1584 -455 1598 -435
rect 1618 -455 1626 -435
rect 1584 -497 1626 -455
rect 1698 -435 1742 -397
rect 1698 -455 1710 -435
rect 1730 -455 1742 -435
rect 1698 -497 1742 -455
rect 1792 -435 1834 -397
rect 1792 -455 1806 -435
rect 1826 -455 1834 -435
rect 1792 -497 1834 -455
rect 1908 -435 1950 -397
rect 1908 -455 1916 -435
rect 1936 -455 1950 -435
rect 1908 -497 1950 -455
rect 2000 -428 2045 -397
rect 2000 -435 2044 -428
rect 2000 -455 2012 -435
rect 2032 -455 2044 -435
rect 2000 -497 2044 -455
rect 338 -745 382 -707
rect 338 -765 350 -745
rect 370 -765 382 -745
rect 338 -807 382 -765
rect 432 -745 474 -707
rect 432 -765 446 -745
rect 466 -765 474 -745
rect 432 -807 474 -765
rect 551 -745 595 -707
rect 551 -765 563 -745
rect 583 -765 595 -745
rect 551 -807 595 -765
rect 645 -745 687 -707
rect 645 -765 659 -745
rect 679 -765 687 -745
rect 645 -807 687 -765
rect 759 -745 803 -707
rect 759 -765 771 -745
rect 791 -765 803 -745
rect 759 -807 803 -765
rect 853 -745 895 -707
rect 853 -765 867 -745
rect 887 -765 895 -745
rect 853 -807 895 -765
rect 969 -745 1011 -707
rect 969 -765 977 -745
rect 997 -765 1011 -745
rect 969 -807 1011 -765
rect 1061 -738 1106 -707
rect 1061 -745 1105 -738
rect 1061 -765 1073 -745
rect 1093 -765 1105 -745
rect 1061 -807 1105 -765
<< ndiffc >>
rect 116 1028 134 1046
rect 118 929 136 947
rect 116 841 134 859
rect 118 742 136 760
rect 344 743 364 763
rect 447 747 467 767
rect 557 743 577 763
rect 660 747 680 767
rect 765 743 785 763
rect 868 747 888 767
rect 976 747 996 767
rect 1079 743 1099 763
rect 116 612 134 630
rect 118 513 136 531
rect 1282 499 1302 519
rect 1385 503 1405 523
rect 1495 499 1515 519
rect 1598 503 1618 523
rect 1703 499 1723 519
rect 1806 503 1826 523
rect 1914 503 1934 523
rect 2017 499 2037 519
rect 116 382 134 400
rect 118 283 136 301
rect 343 189 363 209
rect 446 193 466 213
rect 556 189 576 209
rect 659 193 679 213
rect 764 189 784 209
rect 867 193 887 213
rect 975 193 995 213
rect 1078 189 1098 209
rect 117 -75 135 -57
rect 1423 -93 1443 -73
rect 1526 -89 1546 -69
rect 1636 -93 1656 -73
rect 1739 -89 1759 -69
rect 1844 -93 1864 -73
rect 1947 -89 1967 -69
rect 2055 -89 2075 -69
rect 2158 -93 2178 -73
rect 119 -174 137 -156
rect 117 -262 135 -244
rect 119 -361 137 -343
rect 345 -360 365 -340
rect 448 -356 468 -336
rect 558 -360 578 -340
rect 661 -356 681 -336
rect 766 -360 786 -340
rect 869 -356 889 -336
rect 977 -356 997 -336
rect 1080 -360 1100 -340
rect 117 -491 135 -473
rect 119 -590 137 -572
rect 1283 -604 1303 -584
rect 1386 -600 1406 -580
rect 1496 -604 1516 -584
rect 1599 -600 1619 -580
rect 1704 -604 1724 -584
rect 1807 -600 1827 -580
rect 1915 -600 1935 -580
rect 2018 -604 2038 -584
rect 117 -721 135 -703
rect 119 -820 137 -802
rect 344 -914 364 -894
rect 447 -910 467 -890
rect 557 -914 577 -894
rect 660 -910 680 -890
rect 765 -914 785 -894
rect 868 -910 888 -890
rect 976 -910 996 -890
rect 1079 -914 1099 -894
<< pdiffc >>
rect 350 892 370 912
rect 446 892 466 912
rect 563 892 583 912
rect 659 892 679 912
rect 771 892 791 912
rect 867 892 887 912
rect 977 892 997 912
rect 1073 892 1093 912
rect 1288 648 1308 668
rect 1384 648 1404 668
rect 1501 648 1521 668
rect 1597 648 1617 668
rect 1709 648 1729 668
rect 1805 648 1825 668
rect 1915 648 1935 668
rect 2011 648 2031 668
rect 349 338 369 358
rect 445 338 465 358
rect 562 338 582 358
rect 658 338 678 358
rect 770 338 790 358
rect 866 338 886 358
rect 976 338 996 358
rect 1072 338 1092 358
rect 1429 56 1449 76
rect 1525 56 1545 76
rect 1642 56 1662 76
rect 1738 56 1758 76
rect 1850 56 1870 76
rect 1946 56 1966 76
rect 2056 56 2076 76
rect 2152 56 2172 76
rect 351 -211 371 -191
rect 447 -211 467 -191
rect 564 -211 584 -191
rect 660 -211 680 -191
rect 772 -211 792 -191
rect 868 -211 888 -191
rect 978 -211 998 -191
rect 1074 -211 1094 -191
rect 1289 -455 1309 -435
rect 1385 -455 1405 -435
rect 1502 -455 1522 -435
rect 1598 -455 1618 -435
rect 1710 -455 1730 -435
rect 1806 -455 1826 -435
rect 1916 -455 1936 -435
rect 2012 -455 2032 -435
rect 350 -765 370 -745
rect 446 -765 466 -745
rect 563 -765 583 -745
rect 659 -765 679 -745
rect 771 -765 791 -745
rect 867 -765 887 -745
rect 977 -765 997 -745
rect 1073 -765 1093 -745
<< psubdiff >>
rect 418 676 529 690
rect 418 646 459 676
rect 487 646 529 676
rect 418 631 529 646
rect 1356 432 1467 446
rect 1356 402 1397 432
rect 1425 402 1467 432
rect 1356 387 1467 402
rect 417 122 528 136
rect 417 92 458 122
rect 486 92 528 122
rect 417 77 528 92
rect 1497 -160 1608 -146
rect 1497 -190 1538 -160
rect 1566 -190 1608 -160
rect 1497 -205 1608 -190
rect 419 -427 530 -413
rect 419 -457 460 -427
rect 488 -457 530 -427
rect 419 -472 530 -457
rect 1357 -671 1468 -657
rect 1357 -701 1398 -671
rect 1426 -701 1468 -671
rect 1357 -716 1468 -701
rect 418 -981 529 -967
rect 418 -1011 459 -981
rect 487 -1011 529 -981
rect 418 -1026 529 -1011
<< nsubdiff >>
rect 419 1023 529 1037
rect 419 993 462 1023
rect 490 993 529 1023
rect 419 978 529 993
rect 1357 779 1467 793
rect 1357 749 1400 779
rect 1428 749 1467 779
rect 1357 734 1467 749
rect 418 469 528 483
rect 418 439 461 469
rect 489 439 528 469
rect 418 424 528 439
rect 1498 187 1608 201
rect 1498 157 1541 187
rect 1569 157 1608 187
rect 1498 142 1608 157
rect 420 -80 530 -66
rect 420 -110 463 -80
rect 491 -110 530 -80
rect 420 -125 530 -110
rect 1358 -324 1468 -310
rect 1358 -354 1401 -324
rect 1429 -354 1468 -324
rect 1358 -369 1468 -354
rect 419 -634 529 -620
rect 419 -664 462 -634
rect 490 -664 529 -634
rect 419 -679 529 -664
<< psubdiffcont >>
rect 459 646 487 676
rect 1397 402 1425 432
rect 458 92 486 122
rect 1538 -190 1566 -160
rect 460 -457 488 -427
rect 1398 -701 1426 -671
rect 459 -1011 487 -981
<< nsubdiffcont >>
rect 462 993 490 1023
rect 1400 749 1428 779
rect 461 439 489 469
rect 1541 157 1569 187
rect 463 -110 491 -80
rect 1401 -354 1429 -324
rect 462 -664 490 -634
<< poly >>
rect 382 950 432 963
rect 595 950 645 963
rect 803 950 853 963
rect 1011 950 1061 963
rect 382 822 432 850
rect 382 802 395 822
rect 415 802 432 822
rect 382 773 432 802
rect 595 821 645 850
rect 595 797 606 821
rect 630 797 645 821
rect 595 773 645 797
rect 803 826 853 850
rect 803 802 815 826
rect 839 802 853 826
rect 803 773 853 802
rect 1011 824 1061 850
rect 1011 798 1029 824
rect 1055 798 1061 824
rect 1011 773 1061 798
rect 382 715 432 731
rect 595 715 645 731
rect 803 715 853 731
rect 1011 715 1061 731
rect 1320 706 1370 719
rect 1533 706 1583 719
rect 1741 706 1791 719
rect 1949 706 1999 719
rect 1320 578 1370 606
rect 1320 558 1333 578
rect 1353 558 1370 578
rect 1320 529 1370 558
rect 1533 577 1583 606
rect 1533 553 1544 577
rect 1568 553 1583 577
rect 1533 529 1583 553
rect 1741 582 1791 606
rect 1741 558 1753 582
rect 1777 558 1791 582
rect 1741 529 1791 558
rect 1949 580 1999 606
rect 1949 554 1967 580
rect 1993 554 1999 580
rect 1949 529 1999 554
rect 1320 471 1370 487
rect 1533 471 1583 487
rect 1741 471 1791 487
rect 1949 471 1999 487
rect 381 396 431 409
rect 594 396 644 409
rect 802 396 852 409
rect 1010 396 1060 409
rect 381 268 431 296
rect 381 248 394 268
rect 414 248 431 268
rect 381 219 431 248
rect 594 267 644 296
rect 594 243 605 267
rect 629 243 644 267
rect 594 219 644 243
rect 802 272 852 296
rect 802 248 814 272
rect 838 248 852 272
rect 802 219 852 248
rect 1010 270 1060 296
rect 1010 244 1028 270
rect 1054 244 1060 270
rect 1010 219 1060 244
rect 381 161 431 177
rect 594 161 644 177
rect 802 161 852 177
rect 1010 161 1060 177
rect 1461 114 1511 127
rect 1674 114 1724 127
rect 1882 114 1932 127
rect 2090 114 2140 127
rect 1461 -14 1511 14
rect 1461 -34 1474 -14
rect 1494 -34 1511 -14
rect 1461 -63 1511 -34
rect 1674 -15 1724 14
rect 1674 -39 1685 -15
rect 1709 -39 1724 -15
rect 1674 -63 1724 -39
rect 1882 -10 1932 14
rect 1882 -34 1894 -10
rect 1918 -34 1932 -10
rect 1882 -63 1932 -34
rect 2090 -12 2140 14
rect 2090 -38 2108 -12
rect 2134 -38 2140 -12
rect 2090 -63 2140 -38
rect 1461 -121 1511 -105
rect 1674 -121 1724 -105
rect 1882 -121 1932 -105
rect 2090 -121 2140 -105
rect 383 -153 433 -140
rect 596 -153 646 -140
rect 804 -153 854 -140
rect 1012 -153 1062 -140
rect 383 -281 433 -253
rect 383 -301 396 -281
rect 416 -301 433 -281
rect 383 -330 433 -301
rect 596 -282 646 -253
rect 596 -306 607 -282
rect 631 -306 646 -282
rect 596 -330 646 -306
rect 804 -277 854 -253
rect 804 -301 816 -277
rect 840 -301 854 -277
rect 804 -330 854 -301
rect 1012 -279 1062 -253
rect 1012 -305 1030 -279
rect 1056 -305 1062 -279
rect 1012 -330 1062 -305
rect 383 -388 433 -372
rect 596 -388 646 -372
rect 804 -388 854 -372
rect 1012 -388 1062 -372
rect 1321 -397 1371 -384
rect 1534 -397 1584 -384
rect 1742 -397 1792 -384
rect 1950 -397 2000 -384
rect 1321 -525 1371 -497
rect 1321 -545 1334 -525
rect 1354 -545 1371 -525
rect 1321 -574 1371 -545
rect 1534 -526 1584 -497
rect 1534 -550 1545 -526
rect 1569 -550 1584 -526
rect 1534 -574 1584 -550
rect 1742 -521 1792 -497
rect 1742 -545 1754 -521
rect 1778 -545 1792 -521
rect 1742 -574 1792 -545
rect 1950 -523 2000 -497
rect 1950 -549 1968 -523
rect 1994 -549 2000 -523
rect 1950 -574 2000 -549
rect 1321 -632 1371 -616
rect 1534 -632 1584 -616
rect 1742 -632 1792 -616
rect 1950 -632 2000 -616
rect 382 -707 432 -694
rect 595 -707 645 -694
rect 803 -707 853 -694
rect 1011 -707 1061 -694
rect 382 -835 432 -807
rect 382 -855 395 -835
rect 415 -855 432 -835
rect 382 -884 432 -855
rect 595 -836 645 -807
rect 595 -860 606 -836
rect 630 -860 645 -836
rect 595 -884 645 -860
rect 803 -831 853 -807
rect 803 -855 815 -831
rect 839 -855 853 -831
rect 803 -884 853 -855
rect 1011 -833 1061 -807
rect 1011 -859 1029 -833
rect 1055 -859 1061 -833
rect 1011 -884 1061 -859
rect 382 -942 432 -926
rect 595 -942 645 -926
rect 803 -942 853 -926
rect 1011 -942 1061 -926
<< polycont >>
rect 395 802 415 822
rect 606 797 630 821
rect 815 802 839 826
rect 1029 798 1055 824
rect 1333 558 1353 578
rect 1544 553 1568 577
rect 1753 558 1777 582
rect 1967 554 1993 580
rect 394 248 414 268
rect 605 243 629 267
rect 814 248 838 272
rect 1028 244 1054 270
rect 1474 -34 1494 -14
rect 1685 -39 1709 -15
rect 1894 -34 1918 -10
rect 2108 -38 2134 -12
rect 396 -301 416 -281
rect 607 -306 631 -282
rect 816 -301 840 -277
rect 1030 -305 1056 -279
rect 1334 -545 1354 -525
rect 1545 -550 1569 -526
rect 1754 -545 1778 -521
rect 1968 -549 1994 -523
rect 395 -855 415 -835
rect 606 -860 630 -836
rect 815 -855 839 -831
rect 1029 -859 1055 -833
<< ndiffres >>
rect 95 1046 152 1065
rect 95 1043 116 1046
rect 1 1028 116 1043
rect 134 1028 152 1046
rect 1 1005 152 1028
rect 1 969 43 1005
rect 0 968 100 969
rect 0 947 156 968
rect 0 929 118 947
rect 136 929 156 947
rect 0 925 156 929
rect 95 909 156 925
rect 95 859 152 878
rect 95 856 116 859
rect 1 841 116 856
rect 134 841 152 859
rect 1 818 152 841
rect 1 782 43 818
rect 0 781 100 782
rect 0 760 156 781
rect 0 742 118 760
rect 136 742 156 760
rect 0 738 156 742
rect 95 722 156 738
rect 95 630 152 649
rect 95 627 116 630
rect 1 612 116 627
rect 134 612 152 630
rect 1 589 152 612
rect 1 553 43 589
rect 0 552 100 553
rect 0 531 156 552
rect 0 513 118 531
rect 136 513 156 531
rect 0 509 156 513
rect 95 493 156 509
rect 95 400 152 419
rect 95 397 116 400
rect 1 382 116 397
rect 134 382 152 400
rect 1 359 152 382
rect 1 323 43 359
rect 0 322 100 323
rect 0 301 156 322
rect 0 283 118 301
rect 136 283 156 301
rect 0 279 156 283
rect 95 263 156 279
rect 96 -57 153 -38
rect 96 -60 117 -57
rect 2 -75 117 -60
rect 135 -75 153 -57
rect 2 -98 153 -75
rect 2 -134 44 -98
rect 1 -135 101 -134
rect 1 -156 157 -135
rect 1 -174 119 -156
rect 137 -174 157 -156
rect 1 -178 157 -174
rect 96 -194 157 -178
rect 96 -244 153 -225
rect 96 -247 117 -244
rect 2 -262 117 -247
rect 135 -262 153 -244
rect 2 -285 153 -262
rect 2 -321 44 -285
rect 1 -322 101 -321
rect 1 -343 157 -322
rect 1 -361 119 -343
rect 137 -361 157 -343
rect 1 -365 157 -361
rect 96 -381 157 -365
rect 96 -473 153 -454
rect 96 -476 117 -473
rect 2 -491 117 -476
rect 135 -491 153 -473
rect 2 -514 153 -491
rect 2 -550 44 -514
rect 1 -551 101 -550
rect 1 -572 157 -551
rect 1 -590 119 -572
rect 137 -590 157 -572
rect 1 -594 157 -590
rect 96 -610 157 -594
rect 96 -703 153 -684
rect 96 -706 117 -703
rect 2 -721 117 -706
rect 135 -721 153 -703
rect 2 -744 153 -721
rect 2 -780 44 -744
rect 1 -781 101 -780
rect 1 -802 157 -781
rect 1 -820 119 -802
rect 137 -820 157 -802
rect 1 -824 157 -820
rect 96 -840 157 -824
<< locali >>
rect 105 1048 144 1105
rect 105 1046 153 1048
rect 105 1028 116 1046
rect 134 1028 153 1046
rect 105 1019 153 1028
rect 106 1018 153 1019
rect 419 1023 529 1037
rect 419 1020 462 1023
rect 419 1015 423 1020
rect 341 993 423 1015
rect 452 993 462 1020
rect 490 996 497 1023
rect 526 1015 529 1023
rect 526 996 591 1015
rect 490 993 591 996
rect 341 991 591 993
rect 109 955 146 956
rect 105 952 146 955
rect 105 947 147 952
rect 105 929 118 947
rect 136 929 147 947
rect 105 915 147 929
rect 185 915 232 919
rect 105 909 232 915
rect 105 880 193 909
rect 222 880 232 909
rect 341 912 378 991
rect 419 978 529 991
rect 493 922 524 923
rect 341 892 350 912
rect 370 892 378 912
rect 341 882 378 892
rect 437 912 524 922
rect 437 892 446 912
rect 466 892 524 912
rect 437 883 524 892
rect 437 882 474 883
rect 105 876 232 880
rect 105 859 144 876
rect 185 875 232 876
rect 105 841 116 859
rect 134 841 144 859
rect 105 832 144 841
rect 106 831 143 832
rect 493 830 524 883
rect 554 912 591 991
rect 762 988 1155 1008
rect 1175 988 1178 1008
rect 762 983 1178 988
rect 762 982 1103 983
rect 706 922 737 923
rect 554 892 563 912
rect 583 892 591 912
rect 554 882 591 892
rect 650 915 737 922
rect 650 912 711 915
rect 650 892 659 912
rect 679 895 711 912
rect 732 895 737 915
rect 679 892 737 895
rect 650 885 737 892
rect 762 912 799 982
rect 1065 981 1102 982
rect 914 922 950 923
rect 762 892 771 912
rect 791 892 799 912
rect 650 883 706 885
rect 650 882 687 883
rect 762 882 799 892
rect 858 912 1006 922
rect 1106 919 1202 921
rect 858 892 867 912
rect 887 892 977 912
rect 997 892 1006 912
rect 858 883 1006 892
rect 1064 912 1202 919
rect 1064 892 1073 912
rect 1093 892 1202 912
rect 1064 883 1202 892
rect 858 882 895 883
rect 914 831 950 883
rect 969 882 1006 883
rect 1065 882 1102 883
rect 385 829 426 830
rect 277 822 426 829
rect 277 802 395 822
rect 415 802 426 822
rect 277 794 426 802
rect 493 826 852 830
rect 493 821 815 826
rect 493 797 606 821
rect 630 802 815 821
rect 839 802 852 826
rect 630 797 852 802
rect 493 794 852 797
rect 914 794 949 831
rect 1017 828 1117 831
rect 1017 824 1084 828
rect 1017 798 1029 824
rect 1055 802 1084 824
rect 1110 802 1117 828
rect 1055 798 1117 802
rect 1017 794 1117 798
rect 493 773 524 794
rect 914 773 950 794
rect 336 772 373 773
rect 110 769 144 770
rect 109 760 146 769
rect 109 742 118 760
rect 136 742 146 760
rect 109 732 146 742
rect 335 763 373 772
rect 335 743 344 763
rect 364 743 373 763
rect 335 735 373 743
rect 439 767 524 773
rect 549 772 586 773
rect 439 747 447 767
rect 467 747 524 767
rect 439 739 524 747
rect 548 763 586 772
rect 548 743 557 763
rect 577 743 586 763
rect 439 738 475 739
rect 548 735 586 743
rect 652 767 737 773
rect 757 772 794 773
rect 652 747 660 767
rect 680 766 737 767
rect 680 747 709 766
rect 652 746 709 747
rect 730 746 737 766
rect 652 739 737 746
rect 756 763 794 772
rect 756 743 765 763
rect 785 743 794 763
rect 652 738 688 739
rect 756 735 794 743
rect 860 767 1004 773
rect 860 747 868 767
rect 888 766 976 767
rect 888 747 919 766
rect 860 746 919 747
rect 944 747 976 766
rect 996 747 1004 767
rect 944 746 1004 747
rect 860 739 1004 746
rect 860 738 896 739
rect 968 738 1004 739
rect 1070 772 1107 773
rect 1070 771 1108 772
rect 1070 763 1134 771
rect 1070 743 1079 763
rect 1099 749 1134 763
rect 1154 749 1157 769
rect 1099 744 1157 749
rect 1099 743 1134 744
rect 110 704 144 732
rect 336 706 373 735
rect 337 704 373 706
rect 549 704 586 735
rect 110 703 282 704
rect 110 671 296 703
rect 337 682 586 704
rect 757 703 794 735
rect 1070 731 1134 743
rect 1174 705 1201 883
rect 1357 779 1467 793
rect 1357 776 1400 779
rect 1357 771 1361 776
rect 1033 703 1201 705
rect 757 697 1201 703
rect 110 639 144 671
rect 106 630 144 639
rect 106 612 116 630
rect 134 612 144 630
rect 106 606 144 612
rect 262 608 296 671
rect 418 676 529 682
rect 418 668 459 676
rect 418 648 426 668
rect 445 648 459 668
rect 418 646 459 648
rect 487 668 529 676
rect 487 648 503 668
rect 522 648 529 668
rect 487 646 529 648
rect 418 631 529 646
rect 756 677 1201 697
rect 756 608 794 677
rect 1033 676 1201 677
rect 1279 749 1361 771
rect 1390 749 1400 776
rect 1428 752 1435 779
rect 1464 771 1467 779
rect 1464 752 1529 771
rect 1428 749 1529 752
rect 1279 747 1529 749
rect 1279 668 1316 747
rect 1357 734 1467 747
rect 1431 678 1462 679
rect 1279 648 1288 668
rect 1308 648 1316 668
rect 1279 638 1316 648
rect 1375 668 1462 678
rect 1375 648 1384 668
rect 1404 648 1462 668
rect 1375 639 1462 648
rect 1375 638 1412 639
rect 106 602 143 606
rect 262 597 794 608
rect 261 581 794 597
rect 1431 586 1462 639
rect 1492 668 1529 747
rect 1700 744 2093 764
rect 2113 744 2116 764
rect 1700 739 2116 744
rect 1700 738 2041 739
rect 1644 678 1675 679
rect 1492 648 1501 668
rect 1521 648 1529 668
rect 1492 638 1529 648
rect 1588 671 1675 678
rect 1588 668 1649 671
rect 1588 648 1597 668
rect 1617 651 1649 668
rect 1670 651 1675 671
rect 1617 648 1675 651
rect 1588 641 1675 648
rect 1700 668 1737 738
rect 2003 737 2040 738
rect 1852 678 1888 679
rect 1700 648 1709 668
rect 1729 648 1737 668
rect 1588 639 1644 641
rect 1588 638 1625 639
rect 1700 638 1737 648
rect 1796 668 1944 678
rect 2044 675 2140 677
rect 1796 648 1805 668
rect 1825 648 1915 668
rect 1935 648 1944 668
rect 1796 639 1944 648
rect 2002 668 2140 675
rect 2002 648 2011 668
rect 2031 648 2140 668
rect 2002 639 2140 648
rect 1796 638 1833 639
rect 1852 587 1888 639
rect 1907 638 1944 639
rect 2003 638 2040 639
rect 1323 585 1364 586
rect 261 580 775 581
rect 1215 578 1364 585
rect 1215 558 1333 578
rect 1353 558 1364 578
rect 1215 550 1364 558
rect 1431 582 1790 586
rect 1431 577 1753 582
rect 1431 553 1544 577
rect 1568 558 1753 577
rect 1777 558 1790 582
rect 1568 553 1790 558
rect 1431 550 1790 553
rect 1852 550 1887 587
rect 1955 584 2055 587
rect 1955 580 2022 584
rect 1955 554 1967 580
rect 1993 558 2022 580
rect 2048 558 2055 584
rect 1993 554 2055 558
rect 1955 550 2055 554
rect 109 539 146 540
rect 107 531 147 539
rect 107 513 118 531
rect 136 513 147 531
rect 1431 529 1462 550
rect 1852 529 1888 550
rect 1274 528 1311 529
rect 107 465 147 513
rect 1273 519 1311 528
rect 1273 499 1282 519
rect 1302 499 1311 519
rect 1273 491 1311 499
rect 1377 523 1462 529
rect 1487 528 1524 529
rect 1377 503 1385 523
rect 1405 503 1462 523
rect 1377 495 1462 503
rect 1486 519 1524 528
rect 1486 499 1495 519
rect 1515 499 1524 519
rect 1377 494 1413 495
rect 1486 491 1524 499
rect 1590 523 1675 529
rect 1695 528 1732 529
rect 1590 503 1598 523
rect 1618 522 1675 523
rect 1618 503 1647 522
rect 1590 502 1647 503
rect 1668 502 1675 522
rect 1590 495 1675 502
rect 1694 519 1732 528
rect 1694 499 1703 519
rect 1723 499 1732 519
rect 1590 494 1626 495
rect 1694 491 1732 499
rect 1798 523 1942 529
rect 1798 503 1806 523
rect 1826 506 1862 523
rect 1882 506 1914 523
rect 1826 503 1914 506
rect 1934 503 1942 523
rect 1798 495 1942 503
rect 1798 494 1834 495
rect 1906 494 1942 495
rect 2008 528 2045 529
rect 2008 527 2046 528
rect 2008 519 2072 527
rect 2008 499 2017 519
rect 2037 505 2072 519
rect 2092 505 2095 525
rect 2037 500 2095 505
rect 2037 499 2072 500
rect 418 469 528 483
rect 418 466 461 469
rect 107 458 232 465
rect 418 461 422 466
rect 107 439 199 458
rect 224 439 232 458
rect 107 429 232 439
rect 340 439 422 461
rect 451 439 461 466
rect 489 442 496 469
rect 525 461 528 469
rect 1274 462 1311 491
rect 525 442 590 461
rect 1275 460 1311 462
rect 1487 460 1524 491
rect 1695 464 1732 491
rect 2008 487 2072 499
rect 489 439 590 442
rect 340 437 590 439
rect 107 409 147 429
rect 106 400 147 409
rect 106 382 116 400
rect 134 382 147 400
rect 106 373 147 382
rect 106 372 143 373
rect 340 358 377 437
rect 418 424 528 437
rect 492 368 523 369
rect 340 338 349 358
rect 369 338 377 358
rect 340 328 377 338
rect 436 358 523 368
rect 436 338 445 358
rect 465 338 523 358
rect 436 329 523 338
rect 436 328 473 329
rect 109 306 146 310
rect 106 301 146 306
rect 106 283 118 301
rect 136 283 146 301
rect 106 103 146 283
rect 492 276 523 329
rect 553 358 590 437
rect 761 434 1154 454
rect 1174 434 1177 454
rect 1275 438 1524 460
rect 1693 459 1734 464
rect 2112 461 2139 639
rect 1971 459 2139 461
rect 1693 453 2139 459
rect 761 429 1177 434
rect 1356 432 1467 438
rect 761 428 1102 429
rect 705 368 736 369
rect 553 338 562 358
rect 582 338 590 358
rect 553 328 590 338
rect 649 361 736 368
rect 649 358 710 361
rect 649 338 658 358
rect 678 341 710 358
rect 731 341 736 361
rect 678 338 736 341
rect 649 331 736 338
rect 761 358 798 428
rect 1064 427 1101 428
rect 1356 424 1397 432
rect 1356 404 1364 424
rect 1383 404 1397 424
rect 1356 402 1397 404
rect 1425 424 1467 432
rect 1425 404 1441 424
rect 1460 404 1467 424
rect 1693 431 1699 453
rect 1725 433 2139 453
rect 1725 431 1734 433
rect 1971 432 2139 433
rect 1693 422 1734 431
rect 1425 402 1467 404
rect 1356 387 1467 402
rect 913 368 949 369
rect 761 338 770 358
rect 790 338 798 358
rect 649 329 705 331
rect 649 328 686 329
rect 761 328 798 338
rect 857 358 1005 368
rect 1105 365 1201 367
rect 857 338 866 358
rect 886 338 976 358
rect 996 338 1005 358
rect 857 329 1005 338
rect 1063 358 1201 365
rect 1063 338 1072 358
rect 1092 338 1201 358
rect 1063 329 1201 338
rect 857 328 894 329
rect 913 277 949 329
rect 968 328 1005 329
rect 1064 328 1101 329
rect 384 275 425 276
rect 276 268 425 275
rect 276 248 394 268
rect 414 248 425 268
rect 276 240 425 248
rect 492 272 851 276
rect 492 267 814 272
rect 492 243 605 267
rect 629 248 814 267
rect 838 248 851 272
rect 629 243 851 248
rect 492 240 851 243
rect 913 240 948 277
rect 1016 274 1116 277
rect 1016 270 1083 274
rect 1016 244 1028 270
rect 1054 248 1083 270
rect 1109 248 1116 274
rect 1054 244 1116 248
rect 1016 240 1116 244
rect 492 219 523 240
rect 913 219 949 240
rect 335 218 372 219
rect 334 209 372 218
rect 334 189 343 209
rect 363 189 372 209
rect 334 181 372 189
rect 438 213 523 219
rect 548 218 585 219
rect 438 193 446 213
rect 466 193 523 213
rect 438 185 523 193
rect 547 209 585 218
rect 547 189 556 209
rect 576 189 585 209
rect 438 184 474 185
rect 547 181 585 189
rect 651 213 736 219
rect 756 218 793 219
rect 651 193 659 213
rect 679 212 736 213
rect 679 193 708 212
rect 651 192 708 193
rect 729 192 736 212
rect 651 185 736 192
rect 755 209 793 218
rect 755 189 764 209
rect 784 189 793 209
rect 651 184 687 185
rect 755 181 793 189
rect 859 213 1003 219
rect 859 193 867 213
rect 887 210 975 213
rect 887 193 918 210
rect 859 190 918 193
rect 941 193 975 210
rect 995 193 1003 213
rect 941 190 1003 193
rect 859 185 1003 190
rect 859 184 895 185
rect 967 184 1003 185
rect 1069 218 1106 219
rect 1069 217 1107 218
rect 1069 209 1133 217
rect 1069 189 1078 209
rect 1098 195 1133 209
rect 1153 195 1156 215
rect 1098 190 1156 195
rect 1098 189 1133 190
rect 335 152 372 181
rect 336 150 372 152
rect 548 150 585 181
rect 336 128 585 150
rect 756 149 793 181
rect 1069 177 1133 189
rect 1173 151 1200 329
rect 1498 187 1608 201
rect 1498 184 1541 187
rect 1498 179 1502 184
rect 1032 149 1200 151
rect 756 146 1200 149
rect 417 122 528 128
rect 417 114 458 122
rect 106 59 145 103
rect 417 94 425 114
rect 444 94 458 114
rect 417 92 458 94
rect 486 114 528 122
rect 486 94 502 114
rect 521 94 528 114
rect 486 92 528 94
rect 417 77 528 92
rect 754 123 1200 146
rect 106 35 146 59
rect 446 35 493 37
rect 754 35 792 123
rect 1032 122 1200 123
rect 1420 157 1502 179
rect 1531 157 1541 184
rect 1569 160 1576 187
rect 1605 179 1608 187
rect 1605 160 1670 179
rect 1569 157 1670 160
rect 1420 155 1670 157
rect 1420 76 1457 155
rect 1498 142 1608 155
rect 1572 86 1603 87
rect 1420 56 1429 76
rect 1449 56 1457 76
rect 1420 46 1457 56
rect 1516 76 1603 86
rect 1516 56 1525 76
rect 1545 56 1603 76
rect 1516 47 1603 56
rect 1516 46 1553 47
rect 106 2 792 35
rect 106 -55 145 2
rect 754 0 792 2
rect 1572 -6 1603 47
rect 1633 76 1670 155
rect 1841 168 2234 172
rect 1841 151 1860 168
rect 1880 152 2234 168
rect 2254 152 2257 172
rect 1880 151 2257 152
rect 1841 147 2257 151
rect 1841 146 2182 147
rect 1785 86 1816 87
rect 1633 56 1642 76
rect 1662 56 1670 76
rect 1633 46 1670 56
rect 1729 79 1816 86
rect 1729 76 1790 79
rect 1729 56 1738 76
rect 1758 59 1790 76
rect 1811 59 1816 79
rect 1758 56 1816 59
rect 1729 49 1816 56
rect 1841 76 1878 146
rect 2144 145 2181 146
rect 1993 86 2029 87
rect 1841 56 1850 76
rect 1870 56 1878 76
rect 1729 47 1785 49
rect 1729 46 1766 47
rect 1841 46 1878 56
rect 1937 76 2085 86
rect 2185 83 2281 85
rect 1937 56 1946 76
rect 1966 56 2056 76
rect 2076 56 2085 76
rect 1937 47 2085 56
rect 2143 76 2281 83
rect 2143 56 2152 76
rect 2172 56 2281 76
rect 2143 47 2281 56
rect 1937 46 1974 47
rect 1993 -5 2029 47
rect 2048 46 2085 47
rect 2144 46 2181 47
rect 1464 -7 1505 -6
rect 1356 -14 1505 -7
rect 1356 -34 1474 -14
rect 1494 -34 1505 -14
rect 1356 -42 1505 -34
rect 1572 -10 1931 -6
rect 1572 -15 1894 -10
rect 1572 -39 1685 -15
rect 1709 -34 1894 -15
rect 1918 -34 1931 -10
rect 1709 -39 1931 -34
rect 1572 -42 1931 -39
rect 1993 -42 2028 -5
rect 2096 -8 2196 -5
rect 2096 -12 2163 -8
rect 2096 -38 2108 -12
rect 2134 -34 2163 -12
rect 2189 -34 2196 -8
rect 2134 -38 2196 -34
rect 2096 -42 2196 -38
rect 106 -57 154 -55
rect 106 -75 117 -57
rect 135 -75 154 -57
rect 1572 -63 1603 -42
rect 1993 -63 2029 -42
rect 1415 -64 1452 -63
rect 106 -84 154 -75
rect 107 -85 154 -84
rect 420 -80 530 -66
rect 420 -83 463 -80
rect 420 -88 424 -83
rect 342 -110 424 -88
rect 453 -110 463 -83
rect 491 -107 498 -80
rect 527 -88 530 -80
rect 1414 -73 1452 -64
rect 527 -107 592 -88
rect 1414 -93 1423 -73
rect 1443 -93 1452 -73
rect 491 -110 592 -107
rect 342 -112 592 -110
rect 110 -148 147 -147
rect 106 -151 147 -148
rect 106 -156 148 -151
rect 106 -174 119 -156
rect 137 -174 148 -156
rect 106 -188 148 -174
rect 186 -188 233 -184
rect 106 -194 233 -188
rect 106 -223 194 -194
rect 223 -223 233 -194
rect 342 -191 379 -112
rect 420 -125 530 -112
rect 494 -181 525 -180
rect 342 -211 351 -191
rect 371 -211 379 -191
rect 342 -221 379 -211
rect 438 -191 525 -181
rect 438 -211 447 -191
rect 467 -211 525 -191
rect 438 -220 525 -211
rect 438 -221 475 -220
rect 106 -227 233 -223
rect 106 -244 145 -227
rect 186 -228 233 -227
rect 106 -262 117 -244
rect 135 -262 145 -244
rect 106 -271 145 -262
rect 107 -272 144 -271
rect 494 -273 525 -220
rect 555 -191 592 -112
rect 763 -115 1156 -95
rect 1176 -115 1179 -95
rect 1414 -101 1452 -93
rect 1518 -69 1603 -63
rect 1628 -64 1665 -63
rect 1518 -89 1526 -69
rect 1546 -89 1603 -69
rect 1518 -97 1603 -89
rect 1627 -73 1665 -64
rect 1627 -93 1636 -73
rect 1656 -93 1665 -73
rect 1518 -98 1554 -97
rect 1627 -101 1665 -93
rect 1731 -69 1816 -63
rect 1836 -64 1873 -63
rect 1731 -89 1739 -69
rect 1759 -70 1816 -69
rect 1759 -89 1788 -70
rect 1731 -90 1788 -89
rect 1809 -90 1816 -70
rect 1731 -97 1816 -90
rect 1835 -73 1873 -64
rect 1835 -93 1844 -73
rect 1864 -93 1873 -73
rect 1731 -98 1767 -97
rect 1835 -101 1873 -93
rect 1939 -69 2083 -63
rect 1939 -89 1947 -69
rect 1967 -89 2055 -69
rect 2075 -89 2083 -69
rect 1939 -97 2083 -89
rect 1939 -98 1975 -97
rect 2047 -98 2083 -97
rect 2149 -64 2186 -63
rect 2149 -65 2187 -64
rect 2149 -73 2213 -65
rect 2149 -93 2158 -73
rect 2178 -87 2213 -73
rect 2233 -87 2236 -67
rect 2178 -92 2236 -87
rect 2178 -93 2213 -92
rect 763 -120 1179 -115
rect 763 -121 1104 -120
rect 707 -181 738 -180
rect 555 -211 564 -191
rect 584 -211 592 -191
rect 555 -221 592 -211
rect 651 -188 738 -181
rect 651 -191 712 -188
rect 651 -211 660 -191
rect 680 -208 712 -191
rect 733 -208 738 -188
rect 680 -211 738 -208
rect 651 -218 738 -211
rect 763 -191 800 -121
rect 1066 -122 1103 -121
rect 1415 -130 1452 -101
rect 1416 -132 1452 -130
rect 1628 -132 1665 -101
rect 1416 -154 1665 -132
rect 1836 -133 1873 -101
rect 2149 -105 2213 -93
rect 2253 -131 2280 47
rect 2112 -133 2280 -131
rect 1833 -140 2280 -133
rect 1497 -160 1608 -154
rect 1497 -168 1538 -160
rect 915 -181 951 -180
rect 763 -211 772 -191
rect 792 -211 800 -191
rect 651 -220 707 -218
rect 651 -221 688 -220
rect 763 -221 800 -211
rect 859 -191 1007 -181
rect 1107 -184 1203 -182
rect 859 -211 868 -191
rect 888 -211 978 -191
rect 998 -211 1007 -191
rect 859 -220 1007 -211
rect 1065 -191 1203 -184
rect 1065 -211 1074 -191
rect 1094 -211 1203 -191
rect 1497 -188 1505 -168
rect 1524 -188 1538 -168
rect 1497 -190 1538 -188
rect 1566 -168 1608 -160
rect 1566 -188 1582 -168
rect 1601 -188 1608 -168
rect 1833 -167 1858 -140
rect 1889 -159 2280 -140
rect 1889 -167 1938 -159
rect 2112 -160 2280 -159
rect 1833 -169 1938 -167
rect 1566 -190 1608 -188
rect 1497 -205 1608 -190
rect 1065 -220 1203 -211
rect 859 -221 896 -220
rect 915 -272 951 -220
rect 970 -221 1007 -220
rect 1066 -221 1103 -220
rect 386 -274 427 -273
rect 278 -281 427 -274
rect 278 -301 396 -281
rect 416 -301 427 -281
rect 278 -309 427 -301
rect 494 -277 853 -273
rect 494 -282 816 -277
rect 494 -306 607 -282
rect 631 -301 816 -282
rect 840 -301 853 -277
rect 631 -306 853 -301
rect 494 -309 853 -306
rect 915 -309 950 -272
rect 1018 -275 1118 -272
rect 1018 -279 1085 -275
rect 1018 -305 1030 -279
rect 1056 -301 1085 -279
rect 1111 -301 1118 -275
rect 1056 -305 1118 -301
rect 1018 -309 1118 -305
rect 494 -330 525 -309
rect 915 -330 951 -309
rect 337 -331 374 -330
rect 111 -334 145 -333
rect 110 -343 147 -334
rect 110 -361 119 -343
rect 137 -361 147 -343
rect 110 -371 147 -361
rect 336 -340 374 -331
rect 336 -360 345 -340
rect 365 -360 374 -340
rect 336 -368 374 -360
rect 440 -336 525 -330
rect 550 -331 587 -330
rect 440 -356 448 -336
rect 468 -356 525 -336
rect 440 -364 525 -356
rect 549 -340 587 -331
rect 549 -360 558 -340
rect 578 -360 587 -340
rect 440 -365 476 -364
rect 549 -368 587 -360
rect 653 -336 738 -330
rect 758 -331 795 -330
rect 653 -356 661 -336
rect 681 -337 738 -336
rect 681 -356 710 -337
rect 653 -357 710 -356
rect 731 -357 738 -337
rect 653 -364 738 -357
rect 757 -340 795 -331
rect 757 -360 766 -340
rect 786 -360 795 -340
rect 653 -365 689 -364
rect 757 -368 795 -360
rect 861 -336 1005 -330
rect 861 -356 869 -336
rect 889 -337 977 -336
rect 889 -356 920 -337
rect 861 -357 920 -356
rect 945 -356 977 -337
rect 997 -356 1005 -336
rect 945 -357 1005 -356
rect 861 -364 1005 -357
rect 861 -365 897 -364
rect 969 -365 1005 -364
rect 1071 -331 1108 -330
rect 1071 -332 1109 -331
rect 1071 -340 1135 -332
rect 1071 -360 1080 -340
rect 1100 -354 1135 -340
rect 1155 -354 1158 -334
rect 1100 -359 1158 -354
rect 1100 -360 1135 -359
rect 111 -399 145 -371
rect 337 -397 374 -368
rect 338 -399 374 -397
rect 550 -399 587 -368
rect 111 -400 283 -399
rect 111 -432 297 -400
rect 338 -421 587 -399
rect 758 -400 795 -368
rect 1071 -372 1135 -360
rect 1175 -398 1202 -220
rect 1358 -324 1468 -310
rect 1358 -327 1401 -324
rect 1358 -332 1362 -327
rect 1034 -400 1202 -398
rect 758 -406 1202 -400
rect 111 -464 145 -432
rect 107 -473 145 -464
rect 107 -491 117 -473
rect 135 -491 145 -473
rect 107 -497 145 -491
rect 263 -495 297 -432
rect 419 -427 530 -421
rect 419 -435 460 -427
rect 419 -455 427 -435
rect 446 -455 460 -435
rect 419 -457 460 -455
rect 488 -435 530 -427
rect 488 -455 504 -435
rect 523 -455 530 -435
rect 488 -457 530 -455
rect 419 -472 530 -457
rect 757 -426 1202 -406
rect 757 -495 795 -426
rect 1034 -427 1202 -426
rect 1280 -354 1362 -332
rect 1391 -354 1401 -327
rect 1429 -351 1436 -324
rect 1465 -332 1468 -324
rect 1465 -351 1530 -332
rect 1429 -354 1530 -351
rect 1280 -356 1530 -354
rect 1280 -435 1317 -356
rect 1358 -369 1468 -356
rect 1432 -425 1463 -424
rect 1280 -455 1289 -435
rect 1309 -455 1317 -435
rect 1280 -465 1317 -455
rect 1376 -435 1463 -425
rect 1376 -455 1385 -435
rect 1405 -455 1463 -435
rect 1376 -464 1463 -455
rect 1376 -465 1413 -464
rect 107 -501 144 -497
rect 263 -506 795 -495
rect 262 -522 795 -506
rect 1432 -517 1463 -464
rect 1493 -435 1530 -356
rect 1701 -346 2094 -339
rect 1701 -363 1709 -346
rect 1741 -359 2094 -346
rect 2114 -359 2117 -339
rect 1741 -363 2117 -359
rect 1701 -364 2117 -363
rect 1701 -365 2042 -364
rect 1645 -425 1676 -424
rect 1493 -455 1502 -435
rect 1522 -455 1530 -435
rect 1493 -465 1530 -455
rect 1589 -432 1676 -425
rect 1589 -435 1650 -432
rect 1589 -455 1598 -435
rect 1618 -452 1650 -435
rect 1671 -452 1676 -432
rect 1618 -455 1676 -452
rect 1589 -462 1676 -455
rect 1701 -435 1738 -365
rect 2004 -366 2041 -365
rect 1853 -425 1889 -424
rect 1701 -455 1710 -435
rect 1730 -455 1738 -435
rect 1589 -464 1645 -462
rect 1589 -465 1626 -464
rect 1701 -465 1738 -455
rect 1797 -435 1945 -425
rect 2045 -428 2141 -426
rect 1797 -455 1806 -435
rect 1826 -440 1916 -435
rect 1826 -455 1861 -440
rect 1797 -464 1861 -455
rect 1797 -465 1834 -464
rect 1853 -481 1861 -464
rect 1882 -455 1916 -440
rect 1936 -455 1945 -435
rect 1882 -464 1945 -455
rect 2003 -435 2141 -428
rect 2003 -455 2012 -435
rect 2032 -455 2141 -435
rect 2003 -464 2141 -455
rect 1882 -481 1889 -464
rect 1908 -465 1945 -464
rect 2004 -465 2041 -464
rect 1853 -516 1889 -481
rect 1324 -518 1365 -517
rect 262 -523 776 -522
rect 1216 -525 1365 -518
rect 1216 -545 1334 -525
rect 1354 -545 1365 -525
rect 1216 -553 1365 -545
rect 1432 -521 1791 -517
rect 1432 -526 1754 -521
rect 1432 -550 1545 -526
rect 1569 -545 1754 -526
rect 1778 -545 1791 -521
rect 1569 -550 1791 -545
rect 1432 -553 1791 -550
rect 1853 -553 1888 -516
rect 1956 -519 2056 -516
rect 1956 -523 2023 -519
rect 1956 -549 1968 -523
rect 1994 -545 2023 -523
rect 2049 -545 2056 -519
rect 1994 -549 2056 -545
rect 1956 -553 2056 -549
rect 110 -564 147 -563
rect 108 -572 148 -564
rect 108 -590 119 -572
rect 137 -590 148 -572
rect 1432 -574 1463 -553
rect 1853 -574 1889 -553
rect 1275 -575 1312 -574
rect 108 -638 148 -590
rect 1274 -584 1312 -575
rect 1274 -604 1283 -584
rect 1303 -604 1312 -584
rect 1274 -612 1312 -604
rect 1378 -580 1463 -574
rect 1488 -575 1525 -574
rect 1378 -600 1386 -580
rect 1406 -600 1463 -580
rect 1378 -608 1463 -600
rect 1487 -584 1525 -575
rect 1487 -604 1496 -584
rect 1516 -604 1525 -584
rect 1378 -609 1414 -608
rect 1487 -612 1525 -604
rect 1591 -580 1676 -574
rect 1696 -575 1733 -574
rect 1591 -600 1599 -580
rect 1619 -581 1676 -580
rect 1619 -600 1648 -581
rect 1591 -601 1648 -600
rect 1669 -601 1676 -581
rect 1591 -608 1676 -601
rect 1695 -584 1733 -575
rect 1695 -604 1704 -584
rect 1724 -604 1733 -584
rect 1591 -609 1627 -608
rect 1695 -612 1733 -604
rect 1799 -580 1943 -574
rect 1799 -600 1807 -580
rect 1827 -600 1915 -580
rect 1935 -600 1943 -580
rect 1799 -608 1943 -600
rect 1799 -609 1835 -608
rect 1907 -609 1943 -608
rect 2009 -575 2046 -574
rect 2009 -576 2047 -575
rect 2009 -584 2073 -576
rect 2009 -604 2018 -584
rect 2038 -598 2073 -584
rect 2093 -598 2096 -578
rect 2038 -603 2096 -598
rect 2038 -604 2073 -603
rect 419 -634 529 -620
rect 419 -637 462 -634
rect 108 -645 233 -638
rect 419 -642 423 -637
rect 108 -664 200 -645
rect 225 -664 233 -645
rect 108 -674 233 -664
rect 341 -664 423 -642
rect 452 -664 462 -637
rect 490 -661 497 -634
rect 526 -642 529 -634
rect 1275 -641 1312 -612
rect 526 -661 591 -642
rect 1276 -643 1312 -641
rect 1488 -643 1525 -612
rect 1696 -639 1733 -612
rect 2009 -616 2073 -604
rect 490 -664 591 -661
rect 341 -666 591 -664
rect 108 -694 148 -674
rect 107 -703 148 -694
rect 107 -721 117 -703
rect 135 -721 148 -703
rect 107 -730 148 -721
rect 107 -731 144 -730
rect 341 -745 378 -666
rect 419 -679 529 -666
rect 493 -735 524 -734
rect 341 -765 350 -745
rect 370 -765 378 -745
rect 341 -775 378 -765
rect 437 -745 524 -735
rect 437 -765 446 -745
rect 466 -765 524 -745
rect 437 -774 524 -765
rect 437 -775 474 -774
rect 110 -797 147 -793
rect 107 -802 147 -797
rect 107 -820 119 -802
rect 137 -820 147 -802
rect 107 -1000 147 -820
rect 493 -827 524 -774
rect 554 -745 591 -666
rect 762 -669 1155 -649
rect 1175 -669 1178 -649
rect 1276 -665 1525 -643
rect 1694 -644 1735 -639
rect 2113 -642 2140 -464
rect 1972 -644 2140 -642
rect 1694 -650 2140 -644
rect 762 -674 1178 -669
rect 1357 -671 1468 -665
rect 762 -675 1103 -674
rect 706 -735 737 -734
rect 554 -765 563 -745
rect 583 -765 591 -745
rect 554 -775 591 -765
rect 650 -742 737 -735
rect 650 -745 711 -742
rect 650 -765 659 -745
rect 679 -762 711 -745
rect 732 -762 737 -742
rect 679 -765 737 -762
rect 650 -772 737 -765
rect 762 -745 799 -675
rect 1065 -676 1102 -675
rect 1357 -679 1398 -671
rect 1357 -699 1365 -679
rect 1384 -699 1398 -679
rect 1357 -701 1398 -699
rect 1426 -679 1468 -671
rect 1426 -699 1442 -679
rect 1461 -699 1468 -679
rect 1694 -672 1700 -650
rect 1726 -670 2140 -650
rect 1726 -672 1735 -670
rect 1972 -671 2140 -670
rect 1694 -681 1735 -672
rect 1426 -701 1468 -699
rect 1357 -716 1468 -701
rect 914 -735 950 -734
rect 762 -765 771 -745
rect 791 -765 799 -745
rect 650 -774 706 -772
rect 650 -775 687 -774
rect 762 -775 799 -765
rect 858 -745 1006 -735
rect 1106 -738 1202 -736
rect 858 -765 867 -745
rect 887 -765 977 -745
rect 997 -765 1006 -745
rect 858 -774 1006 -765
rect 1064 -745 1202 -738
rect 1064 -765 1073 -745
rect 1093 -765 1202 -745
rect 1064 -774 1202 -765
rect 858 -775 895 -774
rect 914 -826 950 -774
rect 969 -775 1006 -774
rect 1065 -775 1102 -774
rect 385 -828 426 -827
rect 277 -835 426 -828
rect 277 -855 395 -835
rect 415 -855 426 -835
rect 277 -863 426 -855
rect 493 -831 852 -827
rect 493 -836 815 -831
rect 493 -860 606 -836
rect 630 -855 815 -836
rect 839 -855 852 -831
rect 630 -860 852 -855
rect 493 -863 852 -860
rect 914 -863 949 -826
rect 1017 -829 1117 -826
rect 1017 -833 1084 -829
rect 1017 -859 1029 -833
rect 1055 -855 1084 -833
rect 1110 -855 1117 -829
rect 1055 -859 1117 -855
rect 1017 -863 1117 -859
rect 493 -884 524 -863
rect 914 -884 950 -863
rect 336 -885 373 -884
rect 335 -894 373 -885
rect 335 -914 344 -894
rect 364 -914 373 -894
rect 335 -922 373 -914
rect 439 -890 524 -884
rect 549 -885 586 -884
rect 439 -910 447 -890
rect 467 -910 524 -890
rect 439 -918 524 -910
rect 548 -894 586 -885
rect 548 -914 557 -894
rect 577 -914 586 -894
rect 439 -919 475 -918
rect 548 -922 586 -914
rect 652 -890 737 -884
rect 757 -885 794 -884
rect 652 -910 660 -890
rect 680 -891 737 -890
rect 680 -910 709 -891
rect 652 -911 709 -910
rect 730 -911 737 -891
rect 652 -918 737 -911
rect 756 -894 794 -885
rect 756 -914 765 -894
rect 785 -914 794 -894
rect 652 -919 688 -918
rect 756 -922 794 -914
rect 860 -890 1004 -884
rect 860 -910 868 -890
rect 888 -893 976 -890
rect 888 -910 919 -893
rect 860 -913 919 -910
rect 942 -910 976 -893
rect 996 -910 1004 -890
rect 942 -913 1004 -910
rect 860 -918 1004 -913
rect 860 -919 896 -918
rect 968 -919 1004 -918
rect 1070 -885 1107 -884
rect 1070 -886 1108 -885
rect 1070 -894 1134 -886
rect 1070 -914 1079 -894
rect 1099 -908 1134 -894
rect 1154 -908 1157 -888
rect 1099 -913 1157 -908
rect 1099 -914 1134 -913
rect 336 -951 373 -922
rect 337 -953 373 -951
rect 549 -953 586 -922
rect 337 -975 586 -953
rect 757 -954 794 -922
rect 1070 -926 1134 -914
rect 1174 -952 1201 -774
rect 1033 -954 1201 -952
rect 757 -957 1201 -954
rect 418 -981 529 -975
rect 418 -989 459 -981
rect 107 -1044 146 -1000
rect 418 -1009 426 -989
rect 445 -1009 459 -989
rect 418 -1011 459 -1009
rect 487 -989 529 -981
rect 487 -1009 503 -989
rect 522 -1009 529 -989
rect 487 -1010 529 -1009
rect 755 -980 1201 -957
rect 487 -1011 530 -1010
rect 107 -1068 147 -1044
rect 418 -1050 530 -1011
rect 447 -1068 494 -1050
rect 755 -1068 793 -980
rect 1033 -981 1201 -980
rect 107 -1101 793 -1068
rect 755 -1103 793 -1101
<< viali >>
rect 423 993 452 1020
rect 497 996 526 1023
rect 193 880 222 909
rect 1155 988 1175 1008
rect 711 895 732 915
rect 1084 802 1110 828
rect 709 746 730 766
rect 919 746 944 766
rect 1134 749 1154 769
rect 426 648 445 668
rect 503 648 522 668
rect 1361 749 1390 776
rect 1435 752 1464 779
rect 2093 744 2113 764
rect 1649 651 1670 671
rect 2022 558 2048 584
rect 1647 502 1668 522
rect 1862 506 1882 523
rect 2072 505 2092 525
rect 199 439 224 458
rect 422 439 451 466
rect 496 442 525 469
rect 1154 434 1174 454
rect 710 341 731 361
rect 1364 404 1383 424
rect 1441 404 1460 424
rect 1699 431 1725 453
rect 1083 248 1109 274
rect 708 192 729 212
rect 918 190 941 210
rect 1133 195 1153 215
rect 425 94 444 114
rect 502 94 521 114
rect 1502 157 1531 184
rect 1576 160 1605 187
rect 1860 151 1880 168
rect 2234 152 2254 172
rect 1790 59 1811 79
rect 2163 -34 2189 -8
rect 424 -110 453 -83
rect 498 -107 527 -80
rect 194 -223 223 -194
rect 1156 -115 1176 -95
rect 1788 -90 1809 -70
rect 2213 -87 2233 -67
rect 712 -208 733 -188
rect 1505 -188 1524 -168
rect 1582 -188 1601 -168
rect 1858 -167 1889 -140
rect 1085 -301 1111 -275
rect 710 -357 731 -337
rect 920 -357 945 -337
rect 1135 -354 1155 -334
rect 427 -455 446 -435
rect 504 -455 523 -435
rect 1362 -354 1391 -327
rect 1436 -351 1465 -324
rect 1709 -363 1741 -346
rect 2094 -359 2114 -339
rect 1650 -452 1671 -432
rect 1861 -481 1882 -440
rect 2023 -545 2049 -519
rect 1648 -601 1669 -581
rect 2073 -598 2093 -578
rect 200 -664 225 -645
rect 423 -664 452 -637
rect 497 -661 526 -634
rect 1155 -669 1175 -649
rect 711 -762 732 -742
rect 1365 -699 1384 -679
rect 1442 -699 1461 -679
rect 1700 -672 1726 -650
rect 1084 -855 1110 -829
rect 709 -911 730 -891
rect 919 -913 942 -893
rect 1134 -908 1154 -888
rect 426 -1009 445 -989
rect 503 -1009 522 -989
<< metal1 >>
rect 1150 1091 1185 1093
rect 186 1088 1185 1091
rect 185 1064 1185 1088
rect 185 909 233 1064
rect 419 1023 529 1037
rect 419 1020 497 1023
rect 419 993 423 1020
rect 452 996 497 1020
rect 526 996 529 1023
rect 1150 1013 1185 1064
rect 452 993 529 996
rect 419 978 529 993
rect 1148 1008 1185 1013
rect 1148 988 1155 1008
rect 1175 988 1185 1008
rect 1148 981 1185 988
rect 1148 980 1183 981
rect 185 880 193 909
rect 222 880 233 909
rect 185 875 233 880
rect 704 915 736 922
rect 704 895 711 915
rect 732 895 736 915
rect 704 830 736 895
rect 1074 830 1114 831
rect 704 828 1116 830
rect 704 802 1084 828
rect 1110 802 1116 828
rect 704 794 1116 802
rect 704 766 736 794
rect 1149 774 1183 980
rect 2087 847 2121 848
rect 1218 812 2122 847
rect 704 746 709 766
rect 730 746 736 766
rect 704 739 736 746
rect 911 766 950 772
rect 911 746 919 766
rect 944 746 950 766
rect 911 739 950 746
rect 1127 769 1183 774
rect 1127 749 1134 769
rect 1154 749 1183 769
rect 1127 742 1183 749
rect 1127 741 1162 742
rect 919 693 950 739
rect 418 668 529 690
rect 418 648 426 668
rect 445 648 503 668
rect 522 648 529 668
rect 918 676 950 693
rect 1219 676 1256 812
rect 1357 779 1467 793
rect 1357 776 1435 779
rect 1357 749 1361 776
rect 1390 752 1435 776
rect 1464 752 1467 779
rect 2087 769 2121 812
rect 1390 749 1467 752
rect 1357 734 1467 749
rect 2086 764 2121 769
rect 2086 744 2093 764
rect 2113 744 2121 764
rect 2086 736 2121 744
rect 918 663 1256 676
rect 418 631 529 648
rect 919 644 1256 663
rect 1198 643 1256 644
rect 1642 671 1674 678
rect 1642 651 1649 671
rect 1670 651 1674 671
rect 1642 586 1674 651
rect 2012 586 2052 587
rect 1642 584 2054 586
rect 1642 558 2022 584
rect 2048 558 2054 584
rect 1642 550 2054 558
rect 188 511 1184 537
rect 1642 522 1674 550
rect 190 458 232 511
rect 190 439 199 458
rect 224 439 232 458
rect 190 429 232 439
rect 418 469 528 483
rect 418 466 496 469
rect 418 439 422 466
rect 451 442 496 466
rect 525 442 528 469
rect 1148 459 1182 511
rect 1642 502 1647 522
rect 1668 502 1674 522
rect 1642 495 1674 502
rect 1852 523 1890 533
rect 2087 530 2121 736
rect 1852 506 1862 523
rect 1882 506 1890 523
rect 1693 463 1734 464
rect 451 439 528 442
rect 418 424 528 439
rect 1147 454 1182 459
rect 1147 434 1154 454
rect 1174 434 1182 454
rect 1692 453 1734 463
rect 1147 426 1182 434
rect 703 361 735 368
rect 703 341 710 361
rect 731 341 735 361
rect 703 276 735 341
rect 1073 276 1113 277
rect 703 274 1115 276
rect 703 248 1083 274
rect 1109 248 1115 274
rect 703 240 1115 248
rect 703 212 735 240
rect 1148 220 1182 426
rect 1356 424 1467 446
rect 1356 404 1364 424
rect 1383 404 1441 424
rect 1460 404 1467 424
rect 1356 387 1467 404
rect 1692 431 1699 453
rect 1725 431 1734 453
rect 1692 422 1734 431
rect 909 217 952 219
rect 703 192 708 212
rect 729 192 735 212
rect 703 185 735 192
rect 908 210 952 217
rect 908 190 918 210
rect 941 190 952 210
rect 908 186 952 190
rect 1126 215 1182 220
rect 1126 195 1133 215
rect 1153 195 1182 215
rect 1126 188 1182 195
rect 1238 356 1271 357
rect 1692 356 1729 422
rect 1238 327 1729 356
rect 1126 187 1161 188
rect 417 114 528 136
rect 417 94 425 114
rect 444 94 502 114
rect 521 94 528 114
rect 417 77 528 94
rect 908 105 950 186
rect 1238 107 1271 327
rect 1692 325 1729 327
rect 1498 187 1608 201
rect 1498 184 1576 187
rect 1498 157 1502 184
rect 1531 160 1576 184
rect 1605 160 1608 187
rect 1531 157 1608 160
rect 1498 142 1608 157
rect 1852 168 1890 506
rect 2065 525 2121 530
rect 2065 505 2072 525
rect 2092 505 2121 525
rect 2065 498 2121 505
rect 2065 497 2100 498
rect 2230 177 2262 178
rect 1852 151 1860 168
rect 1880 151 1890 168
rect 1852 145 1890 151
rect 2227 172 2262 177
rect 2227 152 2234 172
rect 2254 152 2262 172
rect 2227 144 2262 152
rect 1210 105 1271 107
rect 908 76 1271 105
rect 1783 79 1815 86
rect 908 74 1210 76
rect 1783 59 1790 79
rect 1811 59 1815 79
rect 1783 -6 1815 59
rect 2153 -6 2193 -5
rect 1783 -8 2195 -6
rect 1151 -12 1186 -10
rect 187 -15 1186 -12
rect 186 -39 1186 -15
rect 186 -194 234 -39
rect 420 -80 530 -66
rect 420 -83 498 -80
rect 420 -110 424 -83
rect 453 -107 498 -83
rect 527 -107 530 -80
rect 1151 -90 1186 -39
rect 453 -110 530 -107
rect 420 -125 530 -110
rect 1149 -95 1186 -90
rect 1149 -115 1156 -95
rect 1176 -115 1186 -95
rect 1783 -34 2163 -8
rect 2189 -34 2195 -8
rect 1783 -42 2195 -34
rect 1783 -70 1815 -42
rect 2228 -62 2262 144
rect 1783 -90 1788 -70
rect 1809 -90 1815 -70
rect 1783 -97 1815 -90
rect 2206 -67 2262 -62
rect 2206 -87 2213 -67
rect 2233 -87 2262 -67
rect 2206 -94 2262 -87
rect 2206 -95 2241 -94
rect 1149 -122 1186 -115
rect 1149 -123 1184 -122
rect 186 -223 194 -194
rect 223 -223 234 -194
rect 186 -228 234 -223
rect 705 -188 737 -181
rect 705 -208 712 -188
rect 733 -208 737 -188
rect 705 -273 737 -208
rect 1075 -273 1115 -272
rect 705 -275 1117 -273
rect 705 -301 1085 -275
rect 1111 -301 1117 -275
rect 705 -309 1117 -301
rect 705 -337 737 -309
rect 1150 -329 1184 -123
rect 1854 -140 1893 -133
rect 1497 -168 1608 -146
rect 1497 -188 1505 -168
rect 1524 -188 1582 -168
rect 1601 -188 1608 -168
rect 1497 -205 1608 -188
rect 1854 -167 1858 -140
rect 1889 -167 1893 -140
rect 1701 -256 1754 -252
rect 1219 -291 1754 -256
rect 705 -357 710 -337
rect 731 -357 737 -337
rect 705 -364 737 -357
rect 912 -337 951 -331
rect 912 -357 920 -337
rect 945 -357 951 -337
rect 912 -364 951 -357
rect 1128 -334 1184 -329
rect 1128 -354 1135 -334
rect 1155 -354 1184 -334
rect 1128 -361 1184 -354
rect 1128 -362 1163 -361
rect 920 -410 951 -364
rect 419 -435 530 -413
rect 419 -455 427 -435
rect 446 -455 504 -435
rect 523 -455 530 -435
rect 919 -427 951 -410
rect 1220 -427 1257 -291
rect 1358 -324 1468 -310
rect 1358 -327 1436 -324
rect 1358 -354 1362 -327
rect 1391 -351 1436 -327
rect 1465 -351 1468 -324
rect 1391 -354 1468 -351
rect 1358 -369 1468 -354
rect 1700 -338 1754 -291
rect 1700 -346 1753 -338
rect 1700 -363 1709 -346
rect 1741 -363 1753 -346
rect 1700 -366 1753 -363
rect 919 -440 1257 -427
rect 419 -472 530 -455
rect 920 -459 1257 -440
rect 1199 -460 1257 -459
rect 1643 -432 1675 -425
rect 1643 -452 1650 -432
rect 1671 -452 1675 -432
rect 1643 -517 1675 -452
rect 1854 -440 1893 -167
rect 2089 -338 2123 -327
rect 2087 -339 2123 -338
rect 2087 -359 2094 -339
rect 2114 -359 2123 -339
rect 2087 -367 2123 -359
rect 1854 -481 1861 -440
rect 1882 -481 1893 -440
rect 1854 -496 1893 -481
rect 2013 -517 2053 -516
rect 1643 -519 2055 -517
rect 1643 -545 2023 -519
rect 2049 -545 2055 -519
rect 1643 -553 2055 -545
rect 189 -592 1185 -566
rect 1643 -581 1675 -553
rect 2088 -573 2122 -367
rect 191 -645 233 -592
rect 191 -664 200 -645
rect 225 -664 233 -645
rect 191 -674 233 -664
rect 419 -634 529 -620
rect 419 -637 497 -634
rect 419 -664 423 -637
rect 452 -661 497 -637
rect 526 -661 529 -634
rect 1149 -644 1183 -592
rect 1643 -601 1648 -581
rect 1669 -601 1675 -581
rect 1643 -608 1675 -601
rect 2066 -578 2122 -573
rect 2066 -598 2073 -578
rect 2093 -598 2122 -578
rect 2066 -605 2122 -598
rect 2066 -606 2101 -605
rect 1694 -640 1735 -639
rect 452 -664 529 -661
rect 419 -679 529 -664
rect 1148 -649 1183 -644
rect 1148 -669 1155 -649
rect 1175 -669 1183 -649
rect 1693 -650 1735 -640
rect 1148 -677 1183 -669
rect 704 -742 736 -735
rect 704 -762 711 -742
rect 732 -762 736 -742
rect 704 -827 736 -762
rect 1074 -827 1114 -826
rect 704 -829 1116 -827
rect 704 -855 1084 -829
rect 1110 -855 1116 -829
rect 704 -863 1116 -855
rect 704 -891 736 -863
rect 1149 -883 1183 -677
rect 1357 -679 1468 -657
rect 1357 -699 1365 -679
rect 1384 -699 1442 -679
rect 1461 -699 1468 -679
rect 1357 -716 1468 -699
rect 1693 -672 1700 -650
rect 1726 -672 1735 -650
rect 1693 -681 1735 -672
rect 910 -886 953 -884
rect 704 -911 709 -891
rect 730 -911 736 -891
rect 704 -918 736 -911
rect 909 -893 953 -886
rect 909 -913 919 -893
rect 942 -913 953 -893
rect 909 -917 953 -913
rect 1127 -888 1183 -883
rect 1127 -908 1134 -888
rect 1154 -908 1183 -888
rect 1127 -915 1183 -908
rect 1239 -747 1272 -746
rect 1693 -747 1730 -681
rect 1239 -776 1730 -747
rect 1127 -916 1162 -915
rect 418 -989 529 -967
rect 418 -1009 426 -989
rect 445 -1009 503 -989
rect 522 -1009 529 -989
rect 418 -1026 529 -1009
rect 909 -998 951 -917
rect 1239 -996 1272 -776
rect 1693 -778 1730 -776
rect 1211 -998 1272 -996
rect 909 -1027 1272 -998
rect 909 -1029 1211 -1027
<< labels >>
rlabel locali 290 804 312 819 1 d0
rlabel metal1 459 1027 487 1032 1 vdd
rlabel metal1 456 634 490 640 1 gnd
rlabel locali 1227 556 1255 577 1 d1
rlabel metal1 1394 390 1428 396 1 gnd
rlabel metal1 1397 783 1425 788 1 vdd
rlabel locali 289 250 311 265 1 d0
rlabel metal1 458 473 486 478 1 vdd
rlabel metal1 455 80 489 86 1 gnd
rlabel locali 110 1089 138 1097 1 vref
rlabel locali 291 -299 313 -284 1 d0
rlabel metal1 460 -76 488 -71 1 vdd
rlabel metal1 457 -469 491 -463 1 gnd
rlabel locali 1228 -547 1256 -526 1 d1
rlabel metal1 1395 -713 1429 -707 1 gnd
rlabel metal1 1398 -320 1426 -315 1 vdd
rlabel locali 290 -853 312 -838 1 d0
rlabel metal1 459 -630 487 -625 1 vdd
rlabel metal1 456 -1023 490 -1017 1 gnd
rlabel locali 1999 3 2021 18 1 vout
rlabel metal1 1538 191 1566 196 1 vdd
rlabel metal1 1535 -202 1569 -196 1 gnd
rlabel locali 1366 -37 1387 -18 1 d2
<< end >>
