magic
tech sky130A
timestamp 1620567396
<< nwell >>
rect 318 9238 645 9312
rect 5374 9279 5701 9353
rect 318 9088 1129 9238
rect 1256 8994 1583 9068
rect 3801 9018 4612 9168
rect 5374 9129 6185 9279
rect 10349 9243 10676 9317
rect 15405 9284 15732 9358
rect 1256 8844 2067 8994
rect 4285 8944 4612 9018
rect 6312 9035 6639 9109
rect 8857 9059 9668 9209
rect 10349 9093 11160 9243
rect 6312 8885 7123 9035
rect 9341 8985 9668 9059
rect 11287 8999 11614 9073
rect 13832 9023 14643 9173
rect 15405 9134 16216 9284
rect 317 8684 644 8758
rect 2862 8708 3673 8858
rect 317 8534 1128 8684
rect 3346 8634 3673 8708
rect 5373 8725 5700 8799
rect 7918 8749 8729 8899
rect 11287 8849 12098 8999
rect 14316 8949 14643 9023
rect 16343 9040 16670 9114
rect 18888 9064 19699 9214
rect 16343 8890 17154 9040
rect 19372 8990 19699 9064
rect 1397 8402 1724 8476
rect 3800 8464 4611 8614
rect 5373 8575 6184 8725
rect 8402 8675 8729 8749
rect 10348 8689 10675 8763
rect 12893 8713 13704 8863
rect 1397 8252 2208 8402
rect 4284 8390 4611 8464
rect 6453 8443 6780 8517
rect 8856 8505 9667 8655
rect 10348 8539 11159 8689
rect 13377 8639 13704 8713
rect 15404 8730 15731 8804
rect 17949 8754 18760 8904
rect 319 8135 646 8209
rect 2722 8197 3533 8347
rect 6453 8293 7264 8443
rect 9340 8431 9667 8505
rect 11428 8407 11755 8481
rect 13831 8469 14642 8619
rect 15404 8580 16215 8730
rect 18433 8680 18760 8754
rect 319 7985 1130 8135
rect 3206 8123 3533 8197
rect 5375 8176 5702 8250
rect 7778 8238 8589 8388
rect 11428 8257 12239 8407
rect 14315 8395 14642 8469
rect 16484 8448 16811 8522
rect 18887 8510 19698 8660
rect 1257 7891 1584 7965
rect 3802 7915 4613 8065
rect 5375 8026 6186 8176
rect 8262 8164 8589 8238
rect 10350 8140 10677 8214
rect 12753 8202 13564 8352
rect 16484 8298 17295 8448
rect 19371 8436 19698 8510
rect 1257 7741 2068 7891
rect 4286 7841 4613 7915
rect 6313 7932 6640 8006
rect 8858 7956 9669 8106
rect 10350 7990 11161 8140
rect 13237 8128 13564 8202
rect 15406 8181 15733 8255
rect 17809 8243 18620 8393
rect 6313 7782 7124 7932
rect 9342 7882 9669 7956
rect 11288 7896 11615 7970
rect 13833 7920 14644 8070
rect 15406 8031 16217 8181
rect 18293 8169 18620 8243
rect 318 7581 645 7655
rect 2863 7605 3674 7755
rect 318 7431 1129 7581
rect 3347 7531 3674 7605
rect 5374 7622 5701 7696
rect 7919 7646 8730 7796
rect 11288 7746 12099 7896
rect 14317 7846 14644 7920
rect 16344 7937 16671 8011
rect 18889 7961 19700 8111
rect 16344 7787 17155 7937
rect 19373 7887 19700 7961
rect 1367 7312 1694 7386
rect 3801 7361 4612 7511
rect 5374 7472 6185 7622
rect 8403 7572 8730 7646
rect 10349 7586 10676 7660
rect 12894 7610 13705 7760
rect 1367 7162 2178 7312
rect 4285 7287 4612 7361
rect 6423 7353 6750 7427
rect 8857 7402 9668 7552
rect 10349 7436 11160 7586
rect 13378 7536 13705 7610
rect 15405 7627 15732 7701
rect 17950 7651 18761 7801
rect 319 7032 646 7106
rect 2753 7081 3564 7231
rect 6423 7203 7234 7353
rect 9341 7328 9668 7402
rect 11398 7317 11725 7391
rect 13832 7366 14643 7516
rect 15405 7477 16216 7627
rect 18434 7577 18761 7651
rect 319 6882 1130 7032
rect 3237 7007 3564 7081
rect 5375 7073 5702 7147
rect 7809 7122 8620 7272
rect 11398 7167 12209 7317
rect 14316 7292 14643 7366
rect 16454 7358 16781 7432
rect 18888 7407 19699 7557
rect 1257 6788 1584 6862
rect 3802 6812 4613 6962
rect 5375 6923 6186 7073
rect 8293 7048 8620 7122
rect 10350 7037 10677 7111
rect 12784 7086 13595 7236
rect 16454 7208 17265 7358
rect 19372 7333 19699 7407
rect 1257 6638 2068 6788
rect 4286 6738 4613 6812
rect 6313 6829 6640 6903
rect 8858 6853 9669 7003
rect 10350 6887 11161 7037
rect 13268 7012 13595 7086
rect 15406 7078 15733 7152
rect 17840 7127 18651 7277
rect 6313 6679 7124 6829
rect 9342 6779 9669 6853
rect 11288 6793 11615 6867
rect 13833 6817 14644 6967
rect 15406 6928 16217 7078
rect 18324 7053 18651 7127
rect 318 6478 645 6552
rect 2863 6502 3674 6652
rect 318 6328 1129 6478
rect 3347 6428 3674 6502
rect 5374 6519 5701 6593
rect 7919 6543 8730 6693
rect 11288 6643 12099 6793
rect 14317 6743 14644 6817
rect 16344 6834 16671 6908
rect 18889 6858 19700 7008
rect 16344 6684 17155 6834
rect 19373 6784 19700 6858
rect 1398 6196 1725 6270
rect 3801 6258 4612 6408
rect 5374 6369 6185 6519
rect 8403 6469 8730 6543
rect 10349 6483 10676 6557
rect 12894 6507 13705 6657
rect 1398 6046 2209 6196
rect 4285 6184 4612 6258
rect 6454 6237 6781 6311
rect 8857 6299 9668 6449
rect 10349 6333 11160 6483
rect 13378 6433 13705 6507
rect 15405 6524 15732 6598
rect 17950 6548 18761 6698
rect 320 5929 647 6003
rect 2723 5991 3534 6141
rect 6454 6087 7265 6237
rect 9341 6225 9668 6299
rect 11429 6201 11756 6275
rect 13832 6263 14643 6413
rect 15405 6374 16216 6524
rect 18434 6474 18761 6548
rect 320 5779 1131 5929
rect 3207 5917 3534 5991
rect 5376 5970 5703 6044
rect 7779 6032 8590 6182
rect 11429 6051 12240 6201
rect 14316 6189 14643 6263
rect 16485 6242 16812 6316
rect 18888 6304 19699 6454
rect 1258 5685 1585 5759
rect 3803 5709 4614 5859
rect 5376 5820 6187 5970
rect 8263 5958 8590 6032
rect 10351 5934 10678 6008
rect 12754 5996 13565 6146
rect 16485 6092 17296 6242
rect 19372 6230 19699 6304
rect 1258 5535 2069 5685
rect 4287 5635 4614 5709
rect 6314 5726 6641 5800
rect 8859 5750 9670 5900
rect 10351 5784 11162 5934
rect 13238 5922 13565 5996
rect 15407 5975 15734 6049
rect 17810 6037 18621 6187
rect 6314 5576 7125 5726
rect 9343 5676 9670 5750
rect 11289 5690 11616 5764
rect 13834 5714 14645 5864
rect 15407 5825 16218 5975
rect 18294 5963 18621 6037
rect 319 5375 646 5449
rect 2864 5399 3675 5549
rect 319 5225 1130 5375
rect 3348 5325 3675 5399
rect 5375 5416 5702 5490
rect 7920 5440 8731 5590
rect 11289 5540 12100 5690
rect 14318 5640 14645 5714
rect 16345 5731 16672 5805
rect 18890 5755 19701 5905
rect 16345 5581 17156 5731
rect 19374 5681 19701 5755
rect 1367 5112 1694 5186
rect 3802 5155 4613 5305
rect 5375 5266 6186 5416
rect 8404 5366 8731 5440
rect 10350 5380 10677 5454
rect 12895 5404 13706 5554
rect 1367 4962 2178 5112
rect 4286 5081 4613 5155
rect 6423 5153 6750 5227
rect 8858 5196 9669 5346
rect 10350 5230 11161 5380
rect 13379 5330 13706 5404
rect 15406 5421 15733 5495
rect 17951 5445 18762 5595
rect 320 4826 647 4900
rect 2755 4869 3566 5019
rect 6423 5003 7234 5153
rect 9342 5122 9669 5196
rect 11398 5117 11725 5191
rect 13833 5160 14644 5310
rect 15406 5271 16217 5421
rect 18435 5371 18762 5445
rect 320 4676 1131 4826
rect 3239 4795 3566 4869
rect 5376 4867 5703 4941
rect 7811 4910 8622 5060
rect 11398 4967 12209 5117
rect 14317 5086 14644 5160
rect 16454 5158 16781 5232
rect 18889 5201 19700 5351
rect 1258 4582 1585 4656
rect 3803 4606 4614 4756
rect 5376 4717 6187 4867
rect 8295 4836 8622 4910
rect 10351 4831 10678 4905
rect 12786 4874 13597 5024
rect 16454 5008 17265 5158
rect 19373 5127 19700 5201
rect 1258 4432 2069 4582
rect 4287 4532 4614 4606
rect 6314 4623 6641 4697
rect 8859 4647 9670 4797
rect 10351 4681 11162 4831
rect 13270 4800 13597 4874
rect 15407 4872 15734 4946
rect 17842 4915 18653 5065
rect 6314 4473 7125 4623
rect 9343 4573 9670 4647
rect 11289 4587 11616 4661
rect 13834 4611 14645 4761
rect 15407 4722 16218 4872
rect 18326 4841 18653 4915
rect 319 4272 646 4346
rect 2864 4296 3675 4446
rect 319 4122 1130 4272
rect 3348 4222 3675 4296
rect 5375 4313 5702 4387
rect 7920 4337 8731 4487
rect 11289 4437 12100 4587
rect 14318 4537 14645 4611
rect 16345 4628 16672 4702
rect 18890 4652 19701 4802
rect 16345 4478 17156 4628
rect 19374 4578 19701 4652
rect 1399 3990 1726 4064
rect 3802 4052 4613 4202
rect 5375 4163 6186 4313
rect 8404 4263 8731 4337
rect 10350 4277 10677 4351
rect 12895 4301 13706 4451
rect 1399 3840 2210 3990
rect 4286 3978 4613 4052
rect 6455 4031 6782 4105
rect 8858 4093 9669 4243
rect 10350 4127 11161 4277
rect 13379 4227 13706 4301
rect 15406 4318 15733 4392
rect 17951 4342 18762 4492
rect 321 3723 648 3797
rect 2724 3785 3535 3935
rect 6455 3881 7266 4031
rect 9342 4019 9669 4093
rect 11430 3995 11757 4069
rect 13833 4057 14644 4207
rect 15406 4168 16217 4318
rect 18435 4268 18762 4342
rect 321 3573 1132 3723
rect 3208 3711 3535 3785
rect 5377 3764 5704 3838
rect 7780 3826 8591 3976
rect 11430 3845 12241 3995
rect 14317 3983 14644 4057
rect 16486 4036 16813 4110
rect 18889 4098 19700 4248
rect 1259 3479 1586 3553
rect 3804 3503 4615 3653
rect 5377 3614 6188 3764
rect 8264 3752 8591 3826
rect 10352 3728 10679 3802
rect 12755 3790 13566 3940
rect 16486 3886 17297 4036
rect 19373 4024 19700 4098
rect 1259 3329 2070 3479
rect 4288 3429 4615 3503
rect 6315 3520 6642 3594
rect 8860 3544 9671 3694
rect 10352 3578 11163 3728
rect 13239 3716 13566 3790
rect 15408 3769 15735 3843
rect 17811 3831 18622 3981
rect 6315 3370 7126 3520
rect 9344 3470 9671 3544
rect 11290 3484 11617 3558
rect 13835 3508 14646 3658
rect 15408 3619 16219 3769
rect 18295 3757 18622 3831
rect 320 3169 647 3243
rect 2865 3193 3676 3343
rect 320 3019 1131 3169
rect 3349 3119 3676 3193
rect 5376 3210 5703 3284
rect 7921 3234 8732 3384
rect 11290 3334 12101 3484
rect 14319 3434 14646 3508
rect 16346 3525 16673 3599
rect 18891 3549 19702 3699
rect 16346 3375 17157 3525
rect 19375 3475 19702 3549
rect 1369 2900 1696 2974
rect 3803 2949 4614 3099
rect 5376 3060 6187 3210
rect 8405 3160 8732 3234
rect 10351 3174 10678 3248
rect 12896 3198 13707 3348
rect 1369 2750 2180 2900
rect 4287 2875 4614 2949
rect 6425 2941 6752 3015
rect 8859 2990 9670 3140
rect 10351 3024 11162 3174
rect 13380 3124 13707 3198
rect 15407 3215 15734 3289
rect 17952 3239 18763 3389
rect 321 2620 648 2694
rect 2755 2669 3566 2819
rect 6425 2791 7236 2941
rect 9343 2916 9670 2990
rect 11400 2905 11727 2979
rect 13834 2954 14645 3104
rect 15407 3065 16218 3215
rect 18436 3165 18763 3239
rect 321 2470 1132 2620
rect 3239 2595 3566 2669
rect 5377 2661 5704 2735
rect 7811 2710 8622 2860
rect 11400 2755 12211 2905
rect 14318 2880 14645 2954
rect 16456 2946 16783 3020
rect 18890 2995 19701 3145
rect 1259 2376 1586 2450
rect 3804 2400 4615 2550
rect 5377 2511 6188 2661
rect 8295 2636 8622 2710
rect 10352 2625 10679 2699
rect 12786 2674 13597 2824
rect 16456 2796 17267 2946
rect 19374 2921 19701 2995
rect 1259 2226 2070 2376
rect 4288 2326 4615 2400
rect 6315 2417 6642 2491
rect 8860 2441 9671 2591
rect 10352 2475 11163 2625
rect 13270 2600 13597 2674
rect 15408 2666 15735 2740
rect 17842 2715 18653 2865
rect 6315 2267 7126 2417
rect 9344 2367 9671 2441
rect 11290 2381 11617 2455
rect 13835 2405 14646 2555
rect 15408 2516 16219 2666
rect 18326 2641 18653 2715
rect 320 2066 647 2140
rect 2865 2090 3676 2240
rect 320 1916 1131 2066
rect 3349 2016 3676 2090
rect 5376 2107 5703 2181
rect 7921 2131 8732 2281
rect 11290 2231 12101 2381
rect 14319 2331 14646 2405
rect 16346 2422 16673 2496
rect 18891 2446 19702 2596
rect 16346 2272 17157 2422
rect 19375 2372 19702 2446
rect 1400 1784 1727 1858
rect 3803 1846 4614 1996
rect 5376 1957 6187 2107
rect 8405 2057 8732 2131
rect 10351 2071 10678 2145
rect 12896 2095 13707 2245
rect 1400 1634 2211 1784
rect 4287 1772 4614 1846
rect 6456 1825 6783 1899
rect 8859 1887 9670 2037
rect 10351 1921 11162 2071
rect 13380 2021 13707 2095
rect 15407 2112 15734 2186
rect 17952 2136 18763 2286
rect 322 1517 649 1591
rect 2725 1579 3536 1729
rect 6456 1675 7267 1825
rect 9343 1813 9670 1887
rect 11431 1789 11758 1863
rect 13834 1851 14645 2001
rect 15407 1962 16218 2112
rect 18436 2062 18763 2136
rect 322 1367 1133 1517
rect 3209 1505 3536 1579
rect 5378 1558 5705 1632
rect 7781 1620 8592 1770
rect 11431 1639 12242 1789
rect 14318 1777 14645 1851
rect 16487 1830 16814 1904
rect 18890 1892 19701 2042
rect 1260 1273 1587 1347
rect 3805 1297 4616 1447
rect 5378 1408 6189 1558
rect 8265 1546 8592 1620
rect 10353 1522 10680 1596
rect 12756 1584 13567 1734
rect 16487 1680 17298 1830
rect 19374 1818 19701 1892
rect 1260 1123 2071 1273
rect 4289 1223 4616 1297
rect 6316 1314 6643 1388
rect 8861 1338 9672 1488
rect 10353 1372 11164 1522
rect 13240 1510 13567 1584
rect 15409 1563 15736 1637
rect 17812 1625 18623 1775
rect 6316 1164 7127 1314
rect 9345 1264 9672 1338
rect 11291 1278 11618 1352
rect 13836 1302 14647 1452
rect 15409 1413 16220 1563
rect 18296 1551 18623 1625
rect 321 963 648 1037
rect 2866 987 3677 1137
rect 321 813 1132 963
rect 3350 913 3677 987
rect 5377 1004 5704 1078
rect 7922 1028 8733 1178
rect 11291 1128 12102 1278
rect 14320 1228 14647 1302
rect 16347 1319 16674 1393
rect 18892 1343 19703 1493
rect 16347 1169 17158 1319
rect 19376 1269 19703 1343
rect 3804 743 4615 893
rect 5377 854 6188 1004
rect 8406 954 8733 1028
rect 10352 968 10679 1042
rect 12897 992 13708 1142
rect 8860 784 9671 934
rect 10352 818 11163 968
rect 13381 918 13708 992
rect 15408 1009 15735 1083
rect 17953 1033 18764 1183
rect 4288 669 4615 743
rect 9344 710 9671 784
rect 13835 748 14646 898
rect 15408 859 16219 1009
rect 18437 959 18764 1033
rect 18891 789 19702 939
rect 14319 674 14646 748
rect 19375 715 19702 789
rect 1568 404 1895 478
rect 1568 254 2379 404
rect 4518 384 4845 458
rect 6624 445 6951 519
rect 4518 234 5329 384
rect 6624 295 7435 445
rect 11599 409 11926 483
rect 9452 268 9779 342
rect 9452 118 10263 268
rect 11599 259 12410 409
rect 14549 389 14876 463
rect 16655 450 16982 524
rect 14549 239 15360 389
rect 16655 300 17466 450
<< nmos >>
rect 3869 9227 3919 9269
rect 4077 9227 4127 9269
rect 4285 9227 4335 9269
rect 4498 9227 4548 9269
rect 8925 9268 8975 9310
rect 9133 9268 9183 9310
rect 9341 9268 9391 9310
rect 9554 9268 9604 9310
rect 382 8987 432 9029
rect 595 8987 645 9029
rect 803 8987 853 9029
rect 1011 8987 1061 9029
rect 13900 9232 13950 9274
rect 14108 9232 14158 9274
rect 14316 9232 14366 9274
rect 14529 9232 14579 9274
rect 18956 9273 19006 9315
rect 19164 9273 19214 9315
rect 19372 9273 19422 9315
rect 19585 9273 19635 9315
rect 5438 9028 5488 9070
rect 5651 9028 5701 9070
rect 5859 9028 5909 9070
rect 6067 9028 6117 9070
rect 2930 8917 2980 8959
rect 3138 8917 3188 8959
rect 3346 8917 3396 8959
rect 3559 8917 3609 8959
rect 1320 8743 1370 8785
rect 1533 8743 1583 8785
rect 1741 8743 1791 8785
rect 1949 8743 1999 8785
rect 7986 8958 8036 9000
rect 8194 8958 8244 9000
rect 8402 8958 8452 9000
rect 8615 8958 8665 9000
rect 10413 8992 10463 9034
rect 10626 8992 10676 9034
rect 10834 8992 10884 9034
rect 11042 8992 11092 9034
rect 15469 9033 15519 9075
rect 15682 9033 15732 9075
rect 15890 9033 15940 9075
rect 16098 9033 16148 9075
rect 6376 8784 6426 8826
rect 6589 8784 6639 8826
rect 6797 8784 6847 8826
rect 7005 8784 7055 8826
rect 12961 8922 13011 8964
rect 13169 8922 13219 8964
rect 13377 8922 13427 8964
rect 13590 8922 13640 8964
rect 3868 8673 3918 8715
rect 4076 8673 4126 8715
rect 4284 8673 4334 8715
rect 4497 8673 4547 8715
rect 8924 8714 8974 8756
rect 9132 8714 9182 8756
rect 9340 8714 9390 8756
rect 9553 8714 9603 8756
rect 11351 8748 11401 8790
rect 11564 8748 11614 8790
rect 11772 8748 11822 8790
rect 11980 8748 12030 8790
rect 18017 8963 18067 9005
rect 18225 8963 18275 9005
rect 18433 8963 18483 9005
rect 18646 8963 18696 9005
rect 16407 8789 16457 8831
rect 16620 8789 16670 8831
rect 16828 8789 16878 8831
rect 17036 8789 17086 8831
rect 13899 8678 13949 8720
rect 14107 8678 14157 8720
rect 14315 8678 14365 8720
rect 14528 8678 14578 8720
rect 381 8433 431 8475
rect 594 8433 644 8475
rect 802 8433 852 8475
rect 1010 8433 1060 8475
rect 2790 8406 2840 8448
rect 2998 8406 3048 8448
rect 3206 8406 3256 8448
rect 3419 8406 3469 8448
rect 5437 8474 5487 8516
rect 5650 8474 5700 8516
rect 5858 8474 5908 8516
rect 6066 8474 6116 8516
rect 7846 8447 7896 8489
rect 8054 8447 8104 8489
rect 8262 8447 8312 8489
rect 8475 8447 8525 8489
rect 18955 8719 19005 8761
rect 19163 8719 19213 8761
rect 19371 8719 19421 8761
rect 19584 8719 19634 8761
rect 10412 8438 10462 8480
rect 10625 8438 10675 8480
rect 10833 8438 10883 8480
rect 11041 8438 11091 8480
rect 12821 8411 12871 8453
rect 13029 8411 13079 8453
rect 13237 8411 13287 8453
rect 13450 8411 13500 8453
rect 15468 8479 15518 8521
rect 15681 8479 15731 8521
rect 15889 8479 15939 8521
rect 16097 8479 16147 8521
rect 17877 8452 17927 8494
rect 18085 8452 18135 8494
rect 18293 8452 18343 8494
rect 18506 8452 18556 8494
rect 1461 8151 1511 8193
rect 1674 8151 1724 8193
rect 1882 8151 1932 8193
rect 2090 8151 2140 8193
rect 3870 8124 3920 8166
rect 4078 8124 4128 8166
rect 4286 8124 4336 8166
rect 4499 8124 4549 8166
rect 6517 8192 6567 8234
rect 6730 8192 6780 8234
rect 6938 8192 6988 8234
rect 7146 8192 7196 8234
rect 8926 8165 8976 8207
rect 9134 8165 9184 8207
rect 9342 8165 9392 8207
rect 9555 8165 9605 8207
rect 383 7884 433 7926
rect 596 7884 646 7926
rect 804 7884 854 7926
rect 1012 7884 1062 7926
rect 11492 8156 11542 8198
rect 11705 8156 11755 8198
rect 11913 8156 11963 8198
rect 12121 8156 12171 8198
rect 13901 8129 13951 8171
rect 14109 8129 14159 8171
rect 14317 8129 14367 8171
rect 14530 8129 14580 8171
rect 16548 8197 16598 8239
rect 16761 8197 16811 8239
rect 16969 8197 17019 8239
rect 17177 8197 17227 8239
rect 18957 8170 19007 8212
rect 19165 8170 19215 8212
rect 19373 8170 19423 8212
rect 19586 8170 19636 8212
rect 5439 7925 5489 7967
rect 5652 7925 5702 7967
rect 5860 7925 5910 7967
rect 6068 7925 6118 7967
rect 2931 7814 2981 7856
rect 3139 7814 3189 7856
rect 3347 7814 3397 7856
rect 3560 7814 3610 7856
rect 1321 7640 1371 7682
rect 1534 7640 1584 7682
rect 1742 7640 1792 7682
rect 1950 7640 2000 7682
rect 7987 7855 8037 7897
rect 8195 7855 8245 7897
rect 8403 7855 8453 7897
rect 8616 7855 8666 7897
rect 10414 7889 10464 7931
rect 10627 7889 10677 7931
rect 10835 7889 10885 7931
rect 11043 7889 11093 7931
rect 15470 7930 15520 7972
rect 15683 7930 15733 7972
rect 15891 7930 15941 7972
rect 16099 7930 16149 7972
rect 6377 7681 6427 7723
rect 6590 7681 6640 7723
rect 6798 7681 6848 7723
rect 7006 7681 7056 7723
rect 12962 7819 13012 7861
rect 13170 7819 13220 7861
rect 13378 7819 13428 7861
rect 13591 7819 13641 7861
rect 3869 7570 3919 7612
rect 4077 7570 4127 7612
rect 4285 7570 4335 7612
rect 4498 7570 4548 7612
rect 8925 7611 8975 7653
rect 9133 7611 9183 7653
rect 9341 7611 9391 7653
rect 9554 7611 9604 7653
rect 11352 7645 11402 7687
rect 11565 7645 11615 7687
rect 11773 7645 11823 7687
rect 11981 7645 12031 7687
rect 18018 7860 18068 7902
rect 18226 7860 18276 7902
rect 18434 7860 18484 7902
rect 18647 7860 18697 7902
rect 16408 7686 16458 7728
rect 16621 7686 16671 7728
rect 16829 7686 16879 7728
rect 17037 7686 17087 7728
rect 13900 7575 13950 7617
rect 14108 7575 14158 7617
rect 14316 7575 14366 7617
rect 14529 7575 14579 7617
rect 382 7330 432 7372
rect 595 7330 645 7372
rect 803 7330 853 7372
rect 1011 7330 1061 7372
rect 2821 7290 2871 7332
rect 3029 7290 3079 7332
rect 3237 7290 3287 7332
rect 3450 7290 3500 7332
rect 5438 7371 5488 7413
rect 5651 7371 5701 7413
rect 5859 7371 5909 7413
rect 6067 7371 6117 7413
rect 7877 7331 7927 7373
rect 8085 7331 8135 7373
rect 8293 7331 8343 7373
rect 8506 7331 8556 7373
rect 18956 7616 19006 7658
rect 19164 7616 19214 7658
rect 19372 7616 19422 7658
rect 19585 7616 19635 7658
rect 10413 7335 10463 7377
rect 10626 7335 10676 7377
rect 10834 7335 10884 7377
rect 11042 7335 11092 7377
rect 12852 7295 12902 7337
rect 13060 7295 13110 7337
rect 13268 7295 13318 7337
rect 13481 7295 13531 7337
rect 15469 7376 15519 7418
rect 15682 7376 15732 7418
rect 15890 7376 15940 7418
rect 16098 7376 16148 7418
rect 17908 7336 17958 7378
rect 18116 7336 18166 7378
rect 18324 7336 18374 7378
rect 18537 7336 18587 7378
rect 1431 7061 1481 7103
rect 1644 7061 1694 7103
rect 1852 7061 1902 7103
rect 2060 7061 2110 7103
rect 3870 7021 3920 7063
rect 4078 7021 4128 7063
rect 4286 7021 4336 7063
rect 4499 7021 4549 7063
rect 6487 7102 6537 7144
rect 6700 7102 6750 7144
rect 6908 7102 6958 7144
rect 7116 7102 7166 7144
rect 8926 7062 8976 7104
rect 9134 7062 9184 7104
rect 9342 7062 9392 7104
rect 9555 7062 9605 7104
rect 383 6781 433 6823
rect 596 6781 646 6823
rect 804 6781 854 6823
rect 1012 6781 1062 6823
rect 11462 7066 11512 7108
rect 11675 7066 11725 7108
rect 11883 7066 11933 7108
rect 12091 7066 12141 7108
rect 13901 7026 13951 7068
rect 14109 7026 14159 7068
rect 14317 7026 14367 7068
rect 14530 7026 14580 7068
rect 16518 7107 16568 7149
rect 16731 7107 16781 7149
rect 16939 7107 16989 7149
rect 17147 7107 17197 7149
rect 18957 7067 19007 7109
rect 19165 7067 19215 7109
rect 19373 7067 19423 7109
rect 19586 7067 19636 7109
rect 5439 6822 5489 6864
rect 5652 6822 5702 6864
rect 5860 6822 5910 6864
rect 6068 6822 6118 6864
rect 2931 6711 2981 6753
rect 3139 6711 3189 6753
rect 3347 6711 3397 6753
rect 3560 6711 3610 6753
rect 1321 6537 1371 6579
rect 1534 6537 1584 6579
rect 1742 6537 1792 6579
rect 1950 6537 2000 6579
rect 7987 6752 8037 6794
rect 8195 6752 8245 6794
rect 8403 6752 8453 6794
rect 8616 6752 8666 6794
rect 10414 6786 10464 6828
rect 10627 6786 10677 6828
rect 10835 6786 10885 6828
rect 11043 6786 11093 6828
rect 15470 6827 15520 6869
rect 15683 6827 15733 6869
rect 15891 6827 15941 6869
rect 16099 6827 16149 6869
rect 6377 6578 6427 6620
rect 6590 6578 6640 6620
rect 6798 6578 6848 6620
rect 7006 6578 7056 6620
rect 12962 6716 13012 6758
rect 13170 6716 13220 6758
rect 13378 6716 13428 6758
rect 13591 6716 13641 6758
rect 3869 6467 3919 6509
rect 4077 6467 4127 6509
rect 4285 6467 4335 6509
rect 4498 6467 4548 6509
rect 8925 6508 8975 6550
rect 9133 6508 9183 6550
rect 9341 6508 9391 6550
rect 9554 6508 9604 6550
rect 11352 6542 11402 6584
rect 11565 6542 11615 6584
rect 11773 6542 11823 6584
rect 11981 6542 12031 6584
rect 18018 6757 18068 6799
rect 18226 6757 18276 6799
rect 18434 6757 18484 6799
rect 18647 6757 18697 6799
rect 16408 6583 16458 6625
rect 16621 6583 16671 6625
rect 16829 6583 16879 6625
rect 17037 6583 17087 6625
rect 13900 6472 13950 6514
rect 14108 6472 14158 6514
rect 14316 6472 14366 6514
rect 14529 6472 14579 6514
rect 382 6227 432 6269
rect 595 6227 645 6269
rect 803 6227 853 6269
rect 1011 6227 1061 6269
rect 2791 6200 2841 6242
rect 2999 6200 3049 6242
rect 3207 6200 3257 6242
rect 3420 6200 3470 6242
rect 5438 6268 5488 6310
rect 5651 6268 5701 6310
rect 5859 6268 5909 6310
rect 6067 6268 6117 6310
rect 7847 6241 7897 6283
rect 8055 6241 8105 6283
rect 8263 6241 8313 6283
rect 8476 6241 8526 6283
rect 18956 6513 19006 6555
rect 19164 6513 19214 6555
rect 19372 6513 19422 6555
rect 19585 6513 19635 6555
rect 10413 6232 10463 6274
rect 10626 6232 10676 6274
rect 10834 6232 10884 6274
rect 11042 6232 11092 6274
rect 12822 6205 12872 6247
rect 13030 6205 13080 6247
rect 13238 6205 13288 6247
rect 13451 6205 13501 6247
rect 15469 6273 15519 6315
rect 15682 6273 15732 6315
rect 15890 6273 15940 6315
rect 16098 6273 16148 6315
rect 17878 6246 17928 6288
rect 18086 6246 18136 6288
rect 18294 6246 18344 6288
rect 18507 6246 18557 6288
rect 1462 5945 1512 5987
rect 1675 5945 1725 5987
rect 1883 5945 1933 5987
rect 2091 5945 2141 5987
rect 3871 5918 3921 5960
rect 4079 5918 4129 5960
rect 4287 5918 4337 5960
rect 4500 5918 4550 5960
rect 6518 5986 6568 6028
rect 6731 5986 6781 6028
rect 6939 5986 6989 6028
rect 7147 5986 7197 6028
rect 8927 5959 8977 6001
rect 9135 5959 9185 6001
rect 9343 5959 9393 6001
rect 9556 5959 9606 6001
rect 384 5678 434 5720
rect 597 5678 647 5720
rect 805 5678 855 5720
rect 1013 5678 1063 5720
rect 11493 5950 11543 5992
rect 11706 5950 11756 5992
rect 11914 5950 11964 5992
rect 12122 5950 12172 5992
rect 13902 5923 13952 5965
rect 14110 5923 14160 5965
rect 14318 5923 14368 5965
rect 14531 5923 14581 5965
rect 16549 5991 16599 6033
rect 16762 5991 16812 6033
rect 16970 5991 17020 6033
rect 17178 5991 17228 6033
rect 18958 5964 19008 6006
rect 19166 5964 19216 6006
rect 19374 5964 19424 6006
rect 19587 5964 19637 6006
rect 5440 5719 5490 5761
rect 5653 5719 5703 5761
rect 5861 5719 5911 5761
rect 6069 5719 6119 5761
rect 2932 5608 2982 5650
rect 3140 5608 3190 5650
rect 3348 5608 3398 5650
rect 3561 5608 3611 5650
rect 1322 5434 1372 5476
rect 1535 5434 1585 5476
rect 1743 5434 1793 5476
rect 1951 5434 2001 5476
rect 7988 5649 8038 5691
rect 8196 5649 8246 5691
rect 8404 5649 8454 5691
rect 8617 5649 8667 5691
rect 10415 5683 10465 5725
rect 10628 5683 10678 5725
rect 10836 5683 10886 5725
rect 11044 5683 11094 5725
rect 15471 5724 15521 5766
rect 15684 5724 15734 5766
rect 15892 5724 15942 5766
rect 16100 5724 16150 5766
rect 6378 5475 6428 5517
rect 6591 5475 6641 5517
rect 6799 5475 6849 5517
rect 7007 5475 7057 5517
rect 12963 5613 13013 5655
rect 13171 5613 13221 5655
rect 13379 5613 13429 5655
rect 13592 5613 13642 5655
rect 3870 5364 3920 5406
rect 4078 5364 4128 5406
rect 4286 5364 4336 5406
rect 4499 5364 4549 5406
rect 8926 5405 8976 5447
rect 9134 5405 9184 5447
rect 9342 5405 9392 5447
rect 9555 5405 9605 5447
rect 11353 5439 11403 5481
rect 11566 5439 11616 5481
rect 11774 5439 11824 5481
rect 11982 5439 12032 5481
rect 18019 5654 18069 5696
rect 18227 5654 18277 5696
rect 18435 5654 18485 5696
rect 18648 5654 18698 5696
rect 16409 5480 16459 5522
rect 16622 5480 16672 5522
rect 16830 5480 16880 5522
rect 17038 5480 17088 5522
rect 13901 5369 13951 5411
rect 14109 5369 14159 5411
rect 14317 5369 14367 5411
rect 14530 5369 14580 5411
rect 383 5124 433 5166
rect 596 5124 646 5166
rect 804 5124 854 5166
rect 1012 5124 1062 5166
rect 2823 5078 2873 5120
rect 3031 5078 3081 5120
rect 3239 5078 3289 5120
rect 3452 5078 3502 5120
rect 5439 5165 5489 5207
rect 5652 5165 5702 5207
rect 5860 5165 5910 5207
rect 6068 5165 6118 5207
rect 7879 5119 7929 5161
rect 8087 5119 8137 5161
rect 8295 5119 8345 5161
rect 8508 5119 8558 5161
rect 18957 5410 19007 5452
rect 19165 5410 19215 5452
rect 19373 5410 19423 5452
rect 19586 5410 19636 5452
rect 10414 5129 10464 5171
rect 10627 5129 10677 5171
rect 10835 5129 10885 5171
rect 11043 5129 11093 5171
rect 1431 4861 1481 4903
rect 1644 4861 1694 4903
rect 1852 4861 1902 4903
rect 2060 4861 2110 4903
rect 3871 4815 3921 4857
rect 4079 4815 4129 4857
rect 4287 4815 4337 4857
rect 4500 4815 4550 4857
rect 6487 4902 6537 4944
rect 6700 4902 6750 4944
rect 6908 4902 6958 4944
rect 7116 4902 7166 4944
rect 12854 5083 12904 5125
rect 13062 5083 13112 5125
rect 13270 5083 13320 5125
rect 13483 5083 13533 5125
rect 15470 5170 15520 5212
rect 15683 5170 15733 5212
rect 15891 5170 15941 5212
rect 16099 5170 16149 5212
rect 17910 5124 17960 5166
rect 18118 5124 18168 5166
rect 18326 5124 18376 5166
rect 18539 5124 18589 5166
rect 8927 4856 8977 4898
rect 9135 4856 9185 4898
rect 9343 4856 9393 4898
rect 9556 4856 9606 4898
rect 384 4575 434 4617
rect 597 4575 647 4617
rect 805 4575 855 4617
rect 1013 4575 1063 4617
rect 11462 4866 11512 4908
rect 11675 4866 11725 4908
rect 11883 4866 11933 4908
rect 12091 4866 12141 4908
rect 13902 4820 13952 4862
rect 14110 4820 14160 4862
rect 14318 4820 14368 4862
rect 14531 4820 14581 4862
rect 16518 4907 16568 4949
rect 16731 4907 16781 4949
rect 16939 4907 16989 4949
rect 17147 4907 17197 4949
rect 18958 4861 19008 4903
rect 19166 4861 19216 4903
rect 19374 4861 19424 4903
rect 19587 4861 19637 4903
rect 5440 4616 5490 4658
rect 5653 4616 5703 4658
rect 5861 4616 5911 4658
rect 6069 4616 6119 4658
rect 2932 4505 2982 4547
rect 3140 4505 3190 4547
rect 3348 4505 3398 4547
rect 3561 4505 3611 4547
rect 1322 4331 1372 4373
rect 1535 4331 1585 4373
rect 1743 4331 1793 4373
rect 1951 4331 2001 4373
rect 7988 4546 8038 4588
rect 8196 4546 8246 4588
rect 8404 4546 8454 4588
rect 8617 4546 8667 4588
rect 10415 4580 10465 4622
rect 10628 4580 10678 4622
rect 10836 4580 10886 4622
rect 11044 4580 11094 4622
rect 15471 4621 15521 4663
rect 15684 4621 15734 4663
rect 15892 4621 15942 4663
rect 16100 4621 16150 4663
rect 6378 4372 6428 4414
rect 6591 4372 6641 4414
rect 6799 4372 6849 4414
rect 7007 4372 7057 4414
rect 12963 4510 13013 4552
rect 13171 4510 13221 4552
rect 13379 4510 13429 4552
rect 13592 4510 13642 4552
rect 3870 4261 3920 4303
rect 4078 4261 4128 4303
rect 4286 4261 4336 4303
rect 4499 4261 4549 4303
rect 8926 4302 8976 4344
rect 9134 4302 9184 4344
rect 9342 4302 9392 4344
rect 9555 4302 9605 4344
rect 11353 4336 11403 4378
rect 11566 4336 11616 4378
rect 11774 4336 11824 4378
rect 11982 4336 12032 4378
rect 18019 4551 18069 4593
rect 18227 4551 18277 4593
rect 18435 4551 18485 4593
rect 18648 4551 18698 4593
rect 16409 4377 16459 4419
rect 16622 4377 16672 4419
rect 16830 4377 16880 4419
rect 17038 4377 17088 4419
rect 13901 4266 13951 4308
rect 14109 4266 14159 4308
rect 14317 4266 14367 4308
rect 14530 4266 14580 4308
rect 383 4021 433 4063
rect 596 4021 646 4063
rect 804 4021 854 4063
rect 1012 4021 1062 4063
rect 2792 3994 2842 4036
rect 3000 3994 3050 4036
rect 3208 3994 3258 4036
rect 3421 3994 3471 4036
rect 5439 4062 5489 4104
rect 5652 4062 5702 4104
rect 5860 4062 5910 4104
rect 6068 4062 6118 4104
rect 7848 4035 7898 4077
rect 8056 4035 8106 4077
rect 8264 4035 8314 4077
rect 8477 4035 8527 4077
rect 18957 4307 19007 4349
rect 19165 4307 19215 4349
rect 19373 4307 19423 4349
rect 19586 4307 19636 4349
rect 10414 4026 10464 4068
rect 10627 4026 10677 4068
rect 10835 4026 10885 4068
rect 11043 4026 11093 4068
rect 12823 3999 12873 4041
rect 13031 3999 13081 4041
rect 13239 3999 13289 4041
rect 13452 3999 13502 4041
rect 15470 4067 15520 4109
rect 15683 4067 15733 4109
rect 15891 4067 15941 4109
rect 16099 4067 16149 4109
rect 17879 4040 17929 4082
rect 18087 4040 18137 4082
rect 18295 4040 18345 4082
rect 18508 4040 18558 4082
rect 1463 3739 1513 3781
rect 1676 3739 1726 3781
rect 1884 3739 1934 3781
rect 2092 3739 2142 3781
rect 3872 3712 3922 3754
rect 4080 3712 4130 3754
rect 4288 3712 4338 3754
rect 4501 3712 4551 3754
rect 6519 3780 6569 3822
rect 6732 3780 6782 3822
rect 6940 3780 6990 3822
rect 7148 3780 7198 3822
rect 8928 3753 8978 3795
rect 9136 3753 9186 3795
rect 9344 3753 9394 3795
rect 9557 3753 9607 3795
rect 385 3472 435 3514
rect 598 3472 648 3514
rect 806 3472 856 3514
rect 1014 3472 1064 3514
rect 11494 3744 11544 3786
rect 11707 3744 11757 3786
rect 11915 3744 11965 3786
rect 12123 3744 12173 3786
rect 13903 3717 13953 3759
rect 14111 3717 14161 3759
rect 14319 3717 14369 3759
rect 14532 3717 14582 3759
rect 16550 3785 16600 3827
rect 16763 3785 16813 3827
rect 16971 3785 17021 3827
rect 17179 3785 17229 3827
rect 18959 3758 19009 3800
rect 19167 3758 19217 3800
rect 19375 3758 19425 3800
rect 19588 3758 19638 3800
rect 5441 3513 5491 3555
rect 5654 3513 5704 3555
rect 5862 3513 5912 3555
rect 6070 3513 6120 3555
rect 2933 3402 2983 3444
rect 3141 3402 3191 3444
rect 3349 3402 3399 3444
rect 3562 3402 3612 3444
rect 1323 3228 1373 3270
rect 1536 3228 1586 3270
rect 1744 3228 1794 3270
rect 1952 3228 2002 3270
rect 7989 3443 8039 3485
rect 8197 3443 8247 3485
rect 8405 3443 8455 3485
rect 8618 3443 8668 3485
rect 10416 3477 10466 3519
rect 10629 3477 10679 3519
rect 10837 3477 10887 3519
rect 11045 3477 11095 3519
rect 15472 3518 15522 3560
rect 15685 3518 15735 3560
rect 15893 3518 15943 3560
rect 16101 3518 16151 3560
rect 6379 3269 6429 3311
rect 6592 3269 6642 3311
rect 6800 3269 6850 3311
rect 7008 3269 7058 3311
rect 12964 3407 13014 3449
rect 13172 3407 13222 3449
rect 13380 3407 13430 3449
rect 13593 3407 13643 3449
rect 3871 3158 3921 3200
rect 4079 3158 4129 3200
rect 4287 3158 4337 3200
rect 4500 3158 4550 3200
rect 8927 3199 8977 3241
rect 9135 3199 9185 3241
rect 9343 3199 9393 3241
rect 9556 3199 9606 3241
rect 11354 3233 11404 3275
rect 11567 3233 11617 3275
rect 11775 3233 11825 3275
rect 11983 3233 12033 3275
rect 18020 3448 18070 3490
rect 18228 3448 18278 3490
rect 18436 3448 18486 3490
rect 18649 3448 18699 3490
rect 16410 3274 16460 3316
rect 16623 3274 16673 3316
rect 16831 3274 16881 3316
rect 17039 3274 17089 3316
rect 13902 3163 13952 3205
rect 14110 3163 14160 3205
rect 14318 3163 14368 3205
rect 14531 3163 14581 3205
rect 384 2918 434 2960
rect 597 2918 647 2960
rect 805 2918 855 2960
rect 1013 2918 1063 2960
rect 2823 2878 2873 2920
rect 3031 2878 3081 2920
rect 3239 2878 3289 2920
rect 3452 2878 3502 2920
rect 5440 2959 5490 3001
rect 5653 2959 5703 3001
rect 5861 2959 5911 3001
rect 6069 2959 6119 3001
rect 7879 2919 7929 2961
rect 8087 2919 8137 2961
rect 8295 2919 8345 2961
rect 8508 2919 8558 2961
rect 18958 3204 19008 3246
rect 19166 3204 19216 3246
rect 19374 3204 19424 3246
rect 19587 3204 19637 3246
rect 10415 2923 10465 2965
rect 10628 2923 10678 2965
rect 10836 2923 10886 2965
rect 11044 2923 11094 2965
rect 12854 2883 12904 2925
rect 13062 2883 13112 2925
rect 13270 2883 13320 2925
rect 13483 2883 13533 2925
rect 15471 2964 15521 3006
rect 15684 2964 15734 3006
rect 15892 2964 15942 3006
rect 16100 2964 16150 3006
rect 17910 2924 17960 2966
rect 18118 2924 18168 2966
rect 18326 2924 18376 2966
rect 18539 2924 18589 2966
rect 1433 2649 1483 2691
rect 1646 2649 1696 2691
rect 1854 2649 1904 2691
rect 2062 2649 2112 2691
rect 3872 2609 3922 2651
rect 4080 2609 4130 2651
rect 4288 2609 4338 2651
rect 4501 2609 4551 2651
rect 6489 2690 6539 2732
rect 6702 2690 6752 2732
rect 6910 2690 6960 2732
rect 7118 2690 7168 2732
rect 8928 2650 8978 2692
rect 9136 2650 9186 2692
rect 9344 2650 9394 2692
rect 9557 2650 9607 2692
rect 385 2369 435 2411
rect 598 2369 648 2411
rect 806 2369 856 2411
rect 1014 2369 1064 2411
rect 11464 2654 11514 2696
rect 11677 2654 11727 2696
rect 11885 2654 11935 2696
rect 12093 2654 12143 2696
rect 13903 2614 13953 2656
rect 14111 2614 14161 2656
rect 14319 2614 14369 2656
rect 14532 2614 14582 2656
rect 16520 2695 16570 2737
rect 16733 2695 16783 2737
rect 16941 2695 16991 2737
rect 17149 2695 17199 2737
rect 18959 2655 19009 2697
rect 19167 2655 19217 2697
rect 19375 2655 19425 2697
rect 19588 2655 19638 2697
rect 5441 2410 5491 2452
rect 5654 2410 5704 2452
rect 5862 2410 5912 2452
rect 6070 2410 6120 2452
rect 2933 2299 2983 2341
rect 3141 2299 3191 2341
rect 3349 2299 3399 2341
rect 3562 2299 3612 2341
rect 1323 2125 1373 2167
rect 1536 2125 1586 2167
rect 1744 2125 1794 2167
rect 1952 2125 2002 2167
rect 7989 2340 8039 2382
rect 8197 2340 8247 2382
rect 8405 2340 8455 2382
rect 8618 2340 8668 2382
rect 10416 2374 10466 2416
rect 10629 2374 10679 2416
rect 10837 2374 10887 2416
rect 11045 2374 11095 2416
rect 15472 2415 15522 2457
rect 15685 2415 15735 2457
rect 15893 2415 15943 2457
rect 16101 2415 16151 2457
rect 6379 2166 6429 2208
rect 6592 2166 6642 2208
rect 6800 2166 6850 2208
rect 7008 2166 7058 2208
rect 12964 2304 13014 2346
rect 13172 2304 13222 2346
rect 13380 2304 13430 2346
rect 13593 2304 13643 2346
rect 3871 2055 3921 2097
rect 4079 2055 4129 2097
rect 4287 2055 4337 2097
rect 4500 2055 4550 2097
rect 8927 2096 8977 2138
rect 9135 2096 9185 2138
rect 9343 2096 9393 2138
rect 9556 2096 9606 2138
rect 11354 2130 11404 2172
rect 11567 2130 11617 2172
rect 11775 2130 11825 2172
rect 11983 2130 12033 2172
rect 18020 2345 18070 2387
rect 18228 2345 18278 2387
rect 18436 2345 18486 2387
rect 18649 2345 18699 2387
rect 16410 2171 16460 2213
rect 16623 2171 16673 2213
rect 16831 2171 16881 2213
rect 17039 2171 17089 2213
rect 13902 2060 13952 2102
rect 14110 2060 14160 2102
rect 14318 2060 14368 2102
rect 14531 2060 14581 2102
rect 384 1815 434 1857
rect 597 1815 647 1857
rect 805 1815 855 1857
rect 1013 1815 1063 1857
rect 2793 1788 2843 1830
rect 3001 1788 3051 1830
rect 3209 1788 3259 1830
rect 3422 1788 3472 1830
rect 5440 1856 5490 1898
rect 5653 1856 5703 1898
rect 5861 1856 5911 1898
rect 6069 1856 6119 1898
rect 7849 1829 7899 1871
rect 8057 1829 8107 1871
rect 8265 1829 8315 1871
rect 8478 1829 8528 1871
rect 18958 2101 19008 2143
rect 19166 2101 19216 2143
rect 19374 2101 19424 2143
rect 19587 2101 19637 2143
rect 10415 1820 10465 1862
rect 10628 1820 10678 1862
rect 10836 1820 10886 1862
rect 11044 1820 11094 1862
rect 12824 1793 12874 1835
rect 13032 1793 13082 1835
rect 13240 1793 13290 1835
rect 13453 1793 13503 1835
rect 15471 1861 15521 1903
rect 15684 1861 15734 1903
rect 15892 1861 15942 1903
rect 16100 1861 16150 1903
rect 17880 1834 17930 1876
rect 18088 1834 18138 1876
rect 18296 1834 18346 1876
rect 18509 1834 18559 1876
rect 1464 1533 1514 1575
rect 1677 1533 1727 1575
rect 1885 1533 1935 1575
rect 2093 1533 2143 1575
rect 3873 1506 3923 1548
rect 4081 1506 4131 1548
rect 4289 1506 4339 1548
rect 4502 1506 4552 1548
rect 6520 1574 6570 1616
rect 6733 1574 6783 1616
rect 6941 1574 6991 1616
rect 7149 1574 7199 1616
rect 8929 1547 8979 1589
rect 9137 1547 9187 1589
rect 9345 1547 9395 1589
rect 9558 1547 9608 1589
rect 386 1266 436 1308
rect 599 1266 649 1308
rect 807 1266 857 1308
rect 1015 1266 1065 1308
rect 11495 1538 11545 1580
rect 11708 1538 11758 1580
rect 11916 1538 11966 1580
rect 12124 1538 12174 1580
rect 13904 1511 13954 1553
rect 14112 1511 14162 1553
rect 14320 1511 14370 1553
rect 14533 1511 14583 1553
rect 16551 1579 16601 1621
rect 16764 1579 16814 1621
rect 16972 1579 17022 1621
rect 17180 1579 17230 1621
rect 18960 1552 19010 1594
rect 19168 1552 19218 1594
rect 19376 1552 19426 1594
rect 19589 1552 19639 1594
rect 5442 1307 5492 1349
rect 5655 1307 5705 1349
rect 5863 1307 5913 1349
rect 6071 1307 6121 1349
rect 2934 1196 2984 1238
rect 3142 1196 3192 1238
rect 3350 1196 3400 1238
rect 3563 1196 3613 1238
rect 1324 1022 1374 1064
rect 1537 1022 1587 1064
rect 1745 1022 1795 1064
rect 1953 1022 2003 1064
rect 7990 1237 8040 1279
rect 8198 1237 8248 1279
rect 8406 1237 8456 1279
rect 8619 1237 8669 1279
rect 10417 1271 10467 1313
rect 10630 1271 10680 1313
rect 10838 1271 10888 1313
rect 11046 1271 11096 1313
rect 15473 1312 15523 1354
rect 15686 1312 15736 1354
rect 15894 1312 15944 1354
rect 16102 1312 16152 1354
rect 6380 1063 6430 1105
rect 6593 1063 6643 1105
rect 6801 1063 6851 1105
rect 7009 1063 7059 1105
rect 12965 1201 13015 1243
rect 13173 1201 13223 1243
rect 13381 1201 13431 1243
rect 13594 1201 13644 1243
rect 3872 952 3922 994
rect 4080 952 4130 994
rect 4288 952 4338 994
rect 4501 952 4551 994
rect 8928 993 8978 1035
rect 9136 993 9186 1035
rect 9344 993 9394 1035
rect 9557 993 9607 1035
rect 11355 1027 11405 1069
rect 11568 1027 11618 1069
rect 11776 1027 11826 1069
rect 11984 1027 12034 1069
rect 18021 1242 18071 1284
rect 18229 1242 18279 1284
rect 18437 1242 18487 1284
rect 18650 1242 18700 1284
rect 16411 1068 16461 1110
rect 16624 1068 16674 1110
rect 16832 1068 16882 1110
rect 17040 1068 17090 1110
rect 13903 957 13953 999
rect 14111 957 14161 999
rect 14319 957 14369 999
rect 14532 957 14582 999
rect 385 712 435 754
rect 598 712 648 754
rect 806 712 856 754
rect 1014 712 1064 754
rect 5441 753 5491 795
rect 5654 753 5704 795
rect 5862 753 5912 795
rect 6070 753 6120 795
rect 18959 998 19009 1040
rect 19167 998 19217 1040
rect 19375 998 19425 1040
rect 19588 998 19638 1040
rect 10416 717 10466 759
rect 10629 717 10679 759
rect 10837 717 10887 759
rect 11045 717 11095 759
rect 15472 758 15522 800
rect 15685 758 15735 800
rect 15893 758 15943 800
rect 16101 758 16151 800
rect 1632 153 1682 195
rect 1845 153 1895 195
rect 2053 153 2103 195
rect 2261 153 2311 195
rect 6688 194 6738 236
rect 6901 194 6951 236
rect 7109 194 7159 236
rect 7317 194 7367 236
rect 4582 133 4632 175
rect 4795 133 4845 175
rect 5003 133 5053 175
rect 5211 133 5261 175
rect 11663 158 11713 200
rect 11876 158 11926 200
rect 12084 158 12134 200
rect 12292 158 12342 200
rect 16719 199 16769 241
rect 16932 199 16982 241
rect 17140 199 17190 241
rect 17348 199 17398 241
rect 14613 138 14663 180
rect 14826 138 14876 180
rect 15034 138 15084 180
rect 15242 138 15292 180
rect 9516 17 9566 59
rect 9729 17 9779 59
rect 9937 17 9987 59
rect 10145 17 10195 59
<< pmos >>
rect 382 9106 432 9206
rect 595 9106 645 9206
rect 803 9106 853 9206
rect 1011 9106 1061 9206
rect 3869 9050 3919 9150
rect 4077 9050 4127 9150
rect 4285 9050 4335 9150
rect 4498 9050 4548 9150
rect 5438 9147 5488 9247
rect 5651 9147 5701 9247
rect 5859 9147 5909 9247
rect 6067 9147 6117 9247
rect 8925 9091 8975 9191
rect 9133 9091 9183 9191
rect 9341 9091 9391 9191
rect 9554 9091 9604 9191
rect 10413 9111 10463 9211
rect 10626 9111 10676 9211
rect 10834 9111 10884 9211
rect 11042 9111 11092 9211
rect 1320 8862 1370 8962
rect 1533 8862 1583 8962
rect 1741 8862 1791 8962
rect 1949 8862 1999 8962
rect 2930 8740 2980 8840
rect 3138 8740 3188 8840
rect 3346 8740 3396 8840
rect 3559 8740 3609 8840
rect 6376 8903 6426 9003
rect 6589 8903 6639 9003
rect 6797 8903 6847 9003
rect 7005 8903 7055 9003
rect 13900 9055 13950 9155
rect 14108 9055 14158 9155
rect 14316 9055 14366 9155
rect 14529 9055 14579 9155
rect 15469 9152 15519 9252
rect 15682 9152 15732 9252
rect 15890 9152 15940 9252
rect 16098 9152 16148 9252
rect 18956 9096 19006 9196
rect 19164 9096 19214 9196
rect 19372 9096 19422 9196
rect 19585 9096 19635 9196
rect 7986 8781 8036 8881
rect 8194 8781 8244 8881
rect 8402 8781 8452 8881
rect 8615 8781 8665 8881
rect 11351 8867 11401 8967
rect 11564 8867 11614 8967
rect 11772 8867 11822 8967
rect 11980 8867 12030 8967
rect 381 8552 431 8652
rect 594 8552 644 8652
rect 802 8552 852 8652
rect 1010 8552 1060 8652
rect 3868 8496 3918 8596
rect 4076 8496 4126 8596
rect 4284 8496 4334 8596
rect 4497 8496 4547 8596
rect 5437 8593 5487 8693
rect 5650 8593 5700 8693
rect 5858 8593 5908 8693
rect 6066 8593 6116 8693
rect 12961 8745 13011 8845
rect 13169 8745 13219 8845
rect 13377 8745 13427 8845
rect 13590 8745 13640 8845
rect 16407 8908 16457 9008
rect 16620 8908 16670 9008
rect 16828 8908 16878 9008
rect 17036 8908 17086 9008
rect 18017 8786 18067 8886
rect 18225 8786 18275 8886
rect 18433 8786 18483 8886
rect 18646 8786 18696 8886
rect 8924 8537 8974 8637
rect 9132 8537 9182 8637
rect 9340 8537 9390 8637
rect 9553 8537 9603 8637
rect 10412 8557 10462 8657
rect 10625 8557 10675 8657
rect 10833 8557 10883 8657
rect 11041 8557 11091 8657
rect 13899 8501 13949 8601
rect 14107 8501 14157 8601
rect 14315 8501 14365 8601
rect 14528 8501 14578 8601
rect 15468 8598 15518 8698
rect 15681 8598 15731 8698
rect 15889 8598 15939 8698
rect 16097 8598 16147 8698
rect 18955 8542 19005 8642
rect 19163 8542 19213 8642
rect 19371 8542 19421 8642
rect 19584 8542 19634 8642
rect 1461 8270 1511 8370
rect 1674 8270 1724 8370
rect 1882 8270 1932 8370
rect 2090 8270 2140 8370
rect 2790 8229 2840 8329
rect 2998 8229 3048 8329
rect 3206 8229 3256 8329
rect 3419 8229 3469 8329
rect 6517 8311 6567 8411
rect 6730 8311 6780 8411
rect 6938 8311 6988 8411
rect 7146 8311 7196 8411
rect 7846 8270 7896 8370
rect 8054 8270 8104 8370
rect 8262 8270 8312 8370
rect 8475 8270 8525 8370
rect 11492 8275 11542 8375
rect 11705 8275 11755 8375
rect 11913 8275 11963 8375
rect 12121 8275 12171 8375
rect 12821 8234 12871 8334
rect 13029 8234 13079 8334
rect 13237 8234 13287 8334
rect 13450 8234 13500 8334
rect 16548 8316 16598 8416
rect 16761 8316 16811 8416
rect 16969 8316 17019 8416
rect 17177 8316 17227 8416
rect 17877 8275 17927 8375
rect 18085 8275 18135 8375
rect 18293 8275 18343 8375
rect 18506 8275 18556 8375
rect 383 8003 433 8103
rect 596 8003 646 8103
rect 804 8003 854 8103
rect 1012 8003 1062 8103
rect 3870 7947 3920 8047
rect 4078 7947 4128 8047
rect 4286 7947 4336 8047
rect 4499 7947 4549 8047
rect 5439 8044 5489 8144
rect 5652 8044 5702 8144
rect 5860 8044 5910 8144
rect 6068 8044 6118 8144
rect 8926 7988 8976 8088
rect 9134 7988 9184 8088
rect 9342 7988 9392 8088
rect 9555 7988 9605 8088
rect 10414 8008 10464 8108
rect 10627 8008 10677 8108
rect 10835 8008 10885 8108
rect 11043 8008 11093 8108
rect 1321 7759 1371 7859
rect 1534 7759 1584 7859
rect 1742 7759 1792 7859
rect 1950 7759 2000 7859
rect 2931 7637 2981 7737
rect 3139 7637 3189 7737
rect 3347 7637 3397 7737
rect 3560 7637 3610 7737
rect 6377 7800 6427 7900
rect 6590 7800 6640 7900
rect 6798 7800 6848 7900
rect 7006 7800 7056 7900
rect 13901 7952 13951 8052
rect 14109 7952 14159 8052
rect 14317 7952 14367 8052
rect 14530 7952 14580 8052
rect 15470 8049 15520 8149
rect 15683 8049 15733 8149
rect 15891 8049 15941 8149
rect 16099 8049 16149 8149
rect 18957 7993 19007 8093
rect 19165 7993 19215 8093
rect 19373 7993 19423 8093
rect 19586 7993 19636 8093
rect 7987 7678 8037 7778
rect 8195 7678 8245 7778
rect 8403 7678 8453 7778
rect 8616 7678 8666 7778
rect 11352 7764 11402 7864
rect 11565 7764 11615 7864
rect 11773 7764 11823 7864
rect 11981 7764 12031 7864
rect 382 7449 432 7549
rect 595 7449 645 7549
rect 803 7449 853 7549
rect 1011 7449 1061 7549
rect 3869 7393 3919 7493
rect 4077 7393 4127 7493
rect 4285 7393 4335 7493
rect 4498 7393 4548 7493
rect 5438 7490 5488 7590
rect 5651 7490 5701 7590
rect 5859 7490 5909 7590
rect 6067 7490 6117 7590
rect 12962 7642 13012 7742
rect 13170 7642 13220 7742
rect 13378 7642 13428 7742
rect 13591 7642 13641 7742
rect 16408 7805 16458 7905
rect 16621 7805 16671 7905
rect 16829 7805 16879 7905
rect 17037 7805 17087 7905
rect 18018 7683 18068 7783
rect 18226 7683 18276 7783
rect 18434 7683 18484 7783
rect 18647 7683 18697 7783
rect 8925 7434 8975 7534
rect 9133 7434 9183 7534
rect 9341 7434 9391 7534
rect 9554 7434 9604 7534
rect 10413 7454 10463 7554
rect 10626 7454 10676 7554
rect 10834 7454 10884 7554
rect 11042 7454 11092 7554
rect 13900 7398 13950 7498
rect 14108 7398 14158 7498
rect 14316 7398 14366 7498
rect 14529 7398 14579 7498
rect 15469 7495 15519 7595
rect 15682 7495 15732 7595
rect 15890 7495 15940 7595
rect 16098 7495 16148 7595
rect 18956 7439 19006 7539
rect 19164 7439 19214 7539
rect 19372 7439 19422 7539
rect 19585 7439 19635 7539
rect 1431 7180 1481 7280
rect 1644 7180 1694 7280
rect 1852 7180 1902 7280
rect 2060 7180 2110 7280
rect 6487 7221 6537 7321
rect 6700 7221 6750 7321
rect 6908 7221 6958 7321
rect 7116 7221 7166 7321
rect 2821 7113 2871 7213
rect 3029 7113 3079 7213
rect 3237 7113 3287 7213
rect 3450 7113 3500 7213
rect 7877 7154 7927 7254
rect 8085 7154 8135 7254
rect 8293 7154 8343 7254
rect 8506 7154 8556 7254
rect 11462 7185 11512 7285
rect 11675 7185 11725 7285
rect 11883 7185 11933 7285
rect 12091 7185 12141 7285
rect 16518 7226 16568 7326
rect 16731 7226 16781 7326
rect 16939 7226 16989 7326
rect 17147 7226 17197 7326
rect 12852 7118 12902 7218
rect 13060 7118 13110 7218
rect 13268 7118 13318 7218
rect 13481 7118 13531 7218
rect 17908 7159 17958 7259
rect 18116 7159 18166 7259
rect 18324 7159 18374 7259
rect 18537 7159 18587 7259
rect 383 6900 433 7000
rect 596 6900 646 7000
rect 804 6900 854 7000
rect 1012 6900 1062 7000
rect 3870 6844 3920 6944
rect 4078 6844 4128 6944
rect 4286 6844 4336 6944
rect 4499 6844 4549 6944
rect 5439 6941 5489 7041
rect 5652 6941 5702 7041
rect 5860 6941 5910 7041
rect 6068 6941 6118 7041
rect 8926 6885 8976 6985
rect 9134 6885 9184 6985
rect 9342 6885 9392 6985
rect 9555 6885 9605 6985
rect 10414 6905 10464 7005
rect 10627 6905 10677 7005
rect 10835 6905 10885 7005
rect 11043 6905 11093 7005
rect 1321 6656 1371 6756
rect 1534 6656 1584 6756
rect 1742 6656 1792 6756
rect 1950 6656 2000 6756
rect 2931 6534 2981 6634
rect 3139 6534 3189 6634
rect 3347 6534 3397 6634
rect 3560 6534 3610 6634
rect 6377 6697 6427 6797
rect 6590 6697 6640 6797
rect 6798 6697 6848 6797
rect 7006 6697 7056 6797
rect 13901 6849 13951 6949
rect 14109 6849 14159 6949
rect 14317 6849 14367 6949
rect 14530 6849 14580 6949
rect 15470 6946 15520 7046
rect 15683 6946 15733 7046
rect 15891 6946 15941 7046
rect 16099 6946 16149 7046
rect 18957 6890 19007 6990
rect 19165 6890 19215 6990
rect 19373 6890 19423 6990
rect 19586 6890 19636 6990
rect 7987 6575 8037 6675
rect 8195 6575 8245 6675
rect 8403 6575 8453 6675
rect 8616 6575 8666 6675
rect 11352 6661 11402 6761
rect 11565 6661 11615 6761
rect 11773 6661 11823 6761
rect 11981 6661 12031 6761
rect 382 6346 432 6446
rect 595 6346 645 6446
rect 803 6346 853 6446
rect 1011 6346 1061 6446
rect 3869 6290 3919 6390
rect 4077 6290 4127 6390
rect 4285 6290 4335 6390
rect 4498 6290 4548 6390
rect 5438 6387 5488 6487
rect 5651 6387 5701 6487
rect 5859 6387 5909 6487
rect 6067 6387 6117 6487
rect 12962 6539 13012 6639
rect 13170 6539 13220 6639
rect 13378 6539 13428 6639
rect 13591 6539 13641 6639
rect 16408 6702 16458 6802
rect 16621 6702 16671 6802
rect 16829 6702 16879 6802
rect 17037 6702 17087 6802
rect 18018 6580 18068 6680
rect 18226 6580 18276 6680
rect 18434 6580 18484 6680
rect 18647 6580 18697 6680
rect 8925 6331 8975 6431
rect 9133 6331 9183 6431
rect 9341 6331 9391 6431
rect 9554 6331 9604 6431
rect 10413 6351 10463 6451
rect 10626 6351 10676 6451
rect 10834 6351 10884 6451
rect 11042 6351 11092 6451
rect 13900 6295 13950 6395
rect 14108 6295 14158 6395
rect 14316 6295 14366 6395
rect 14529 6295 14579 6395
rect 15469 6392 15519 6492
rect 15682 6392 15732 6492
rect 15890 6392 15940 6492
rect 16098 6392 16148 6492
rect 18956 6336 19006 6436
rect 19164 6336 19214 6436
rect 19372 6336 19422 6436
rect 19585 6336 19635 6436
rect 1462 6064 1512 6164
rect 1675 6064 1725 6164
rect 1883 6064 1933 6164
rect 2091 6064 2141 6164
rect 2791 6023 2841 6123
rect 2999 6023 3049 6123
rect 3207 6023 3257 6123
rect 3420 6023 3470 6123
rect 6518 6105 6568 6205
rect 6731 6105 6781 6205
rect 6939 6105 6989 6205
rect 7147 6105 7197 6205
rect 7847 6064 7897 6164
rect 8055 6064 8105 6164
rect 8263 6064 8313 6164
rect 8476 6064 8526 6164
rect 11493 6069 11543 6169
rect 11706 6069 11756 6169
rect 11914 6069 11964 6169
rect 12122 6069 12172 6169
rect 12822 6028 12872 6128
rect 13030 6028 13080 6128
rect 13238 6028 13288 6128
rect 13451 6028 13501 6128
rect 16549 6110 16599 6210
rect 16762 6110 16812 6210
rect 16970 6110 17020 6210
rect 17178 6110 17228 6210
rect 17878 6069 17928 6169
rect 18086 6069 18136 6169
rect 18294 6069 18344 6169
rect 18507 6069 18557 6169
rect 384 5797 434 5897
rect 597 5797 647 5897
rect 805 5797 855 5897
rect 1013 5797 1063 5897
rect 3871 5741 3921 5841
rect 4079 5741 4129 5841
rect 4287 5741 4337 5841
rect 4500 5741 4550 5841
rect 5440 5838 5490 5938
rect 5653 5838 5703 5938
rect 5861 5838 5911 5938
rect 6069 5838 6119 5938
rect 8927 5782 8977 5882
rect 9135 5782 9185 5882
rect 9343 5782 9393 5882
rect 9556 5782 9606 5882
rect 10415 5802 10465 5902
rect 10628 5802 10678 5902
rect 10836 5802 10886 5902
rect 11044 5802 11094 5902
rect 1322 5553 1372 5653
rect 1535 5553 1585 5653
rect 1743 5553 1793 5653
rect 1951 5553 2001 5653
rect 2932 5431 2982 5531
rect 3140 5431 3190 5531
rect 3348 5431 3398 5531
rect 3561 5431 3611 5531
rect 6378 5594 6428 5694
rect 6591 5594 6641 5694
rect 6799 5594 6849 5694
rect 7007 5594 7057 5694
rect 13902 5746 13952 5846
rect 14110 5746 14160 5846
rect 14318 5746 14368 5846
rect 14531 5746 14581 5846
rect 15471 5843 15521 5943
rect 15684 5843 15734 5943
rect 15892 5843 15942 5943
rect 16100 5843 16150 5943
rect 18958 5787 19008 5887
rect 19166 5787 19216 5887
rect 19374 5787 19424 5887
rect 19587 5787 19637 5887
rect 7988 5472 8038 5572
rect 8196 5472 8246 5572
rect 8404 5472 8454 5572
rect 8617 5472 8667 5572
rect 11353 5558 11403 5658
rect 11566 5558 11616 5658
rect 11774 5558 11824 5658
rect 11982 5558 12032 5658
rect 383 5243 433 5343
rect 596 5243 646 5343
rect 804 5243 854 5343
rect 1012 5243 1062 5343
rect 3870 5187 3920 5287
rect 4078 5187 4128 5287
rect 4286 5187 4336 5287
rect 4499 5187 4549 5287
rect 5439 5284 5489 5384
rect 5652 5284 5702 5384
rect 5860 5284 5910 5384
rect 6068 5284 6118 5384
rect 12963 5436 13013 5536
rect 13171 5436 13221 5536
rect 13379 5436 13429 5536
rect 13592 5436 13642 5536
rect 16409 5599 16459 5699
rect 16622 5599 16672 5699
rect 16830 5599 16880 5699
rect 17038 5599 17088 5699
rect 18019 5477 18069 5577
rect 18227 5477 18277 5577
rect 18435 5477 18485 5577
rect 18648 5477 18698 5577
rect 8926 5228 8976 5328
rect 9134 5228 9184 5328
rect 9342 5228 9392 5328
rect 9555 5228 9605 5328
rect 10414 5248 10464 5348
rect 10627 5248 10677 5348
rect 10835 5248 10885 5348
rect 11043 5248 11093 5348
rect 1431 4980 1481 5080
rect 1644 4980 1694 5080
rect 1852 4980 1902 5080
rect 2060 4980 2110 5080
rect 6487 5021 6537 5121
rect 6700 5021 6750 5121
rect 6908 5021 6958 5121
rect 7116 5021 7166 5121
rect 13901 5192 13951 5292
rect 14109 5192 14159 5292
rect 14317 5192 14367 5292
rect 14530 5192 14580 5292
rect 15470 5289 15520 5389
rect 15683 5289 15733 5389
rect 15891 5289 15941 5389
rect 16099 5289 16149 5389
rect 18957 5233 19007 5333
rect 19165 5233 19215 5333
rect 19373 5233 19423 5333
rect 19586 5233 19636 5333
rect 2823 4901 2873 5001
rect 3031 4901 3081 5001
rect 3239 4901 3289 5001
rect 3452 4901 3502 5001
rect 7879 4942 7929 5042
rect 8087 4942 8137 5042
rect 8295 4942 8345 5042
rect 8508 4942 8558 5042
rect 11462 4985 11512 5085
rect 11675 4985 11725 5085
rect 11883 4985 11933 5085
rect 12091 4985 12141 5085
rect 16518 5026 16568 5126
rect 16731 5026 16781 5126
rect 16939 5026 16989 5126
rect 17147 5026 17197 5126
rect 384 4694 434 4794
rect 597 4694 647 4794
rect 805 4694 855 4794
rect 1013 4694 1063 4794
rect 3871 4638 3921 4738
rect 4079 4638 4129 4738
rect 4287 4638 4337 4738
rect 4500 4638 4550 4738
rect 5440 4735 5490 4835
rect 5653 4735 5703 4835
rect 5861 4735 5911 4835
rect 6069 4735 6119 4835
rect 12854 4906 12904 5006
rect 13062 4906 13112 5006
rect 13270 4906 13320 5006
rect 13483 4906 13533 5006
rect 17910 4947 17960 5047
rect 18118 4947 18168 5047
rect 18326 4947 18376 5047
rect 18539 4947 18589 5047
rect 8927 4679 8977 4779
rect 9135 4679 9185 4779
rect 9343 4679 9393 4779
rect 9556 4679 9606 4779
rect 10415 4699 10465 4799
rect 10628 4699 10678 4799
rect 10836 4699 10886 4799
rect 11044 4699 11094 4799
rect 1322 4450 1372 4550
rect 1535 4450 1585 4550
rect 1743 4450 1793 4550
rect 1951 4450 2001 4550
rect 2932 4328 2982 4428
rect 3140 4328 3190 4428
rect 3348 4328 3398 4428
rect 3561 4328 3611 4428
rect 6378 4491 6428 4591
rect 6591 4491 6641 4591
rect 6799 4491 6849 4591
rect 7007 4491 7057 4591
rect 13902 4643 13952 4743
rect 14110 4643 14160 4743
rect 14318 4643 14368 4743
rect 14531 4643 14581 4743
rect 15471 4740 15521 4840
rect 15684 4740 15734 4840
rect 15892 4740 15942 4840
rect 16100 4740 16150 4840
rect 18958 4684 19008 4784
rect 19166 4684 19216 4784
rect 19374 4684 19424 4784
rect 19587 4684 19637 4784
rect 7988 4369 8038 4469
rect 8196 4369 8246 4469
rect 8404 4369 8454 4469
rect 8617 4369 8667 4469
rect 11353 4455 11403 4555
rect 11566 4455 11616 4555
rect 11774 4455 11824 4555
rect 11982 4455 12032 4555
rect 383 4140 433 4240
rect 596 4140 646 4240
rect 804 4140 854 4240
rect 1012 4140 1062 4240
rect 3870 4084 3920 4184
rect 4078 4084 4128 4184
rect 4286 4084 4336 4184
rect 4499 4084 4549 4184
rect 5439 4181 5489 4281
rect 5652 4181 5702 4281
rect 5860 4181 5910 4281
rect 6068 4181 6118 4281
rect 12963 4333 13013 4433
rect 13171 4333 13221 4433
rect 13379 4333 13429 4433
rect 13592 4333 13642 4433
rect 16409 4496 16459 4596
rect 16622 4496 16672 4596
rect 16830 4496 16880 4596
rect 17038 4496 17088 4596
rect 18019 4374 18069 4474
rect 18227 4374 18277 4474
rect 18435 4374 18485 4474
rect 18648 4374 18698 4474
rect 8926 4125 8976 4225
rect 9134 4125 9184 4225
rect 9342 4125 9392 4225
rect 9555 4125 9605 4225
rect 10414 4145 10464 4245
rect 10627 4145 10677 4245
rect 10835 4145 10885 4245
rect 11043 4145 11093 4245
rect 13901 4089 13951 4189
rect 14109 4089 14159 4189
rect 14317 4089 14367 4189
rect 14530 4089 14580 4189
rect 15470 4186 15520 4286
rect 15683 4186 15733 4286
rect 15891 4186 15941 4286
rect 16099 4186 16149 4286
rect 18957 4130 19007 4230
rect 19165 4130 19215 4230
rect 19373 4130 19423 4230
rect 19586 4130 19636 4230
rect 1463 3858 1513 3958
rect 1676 3858 1726 3958
rect 1884 3858 1934 3958
rect 2092 3858 2142 3958
rect 2792 3817 2842 3917
rect 3000 3817 3050 3917
rect 3208 3817 3258 3917
rect 3421 3817 3471 3917
rect 6519 3899 6569 3999
rect 6732 3899 6782 3999
rect 6940 3899 6990 3999
rect 7148 3899 7198 3999
rect 7848 3858 7898 3958
rect 8056 3858 8106 3958
rect 8264 3858 8314 3958
rect 8477 3858 8527 3958
rect 11494 3863 11544 3963
rect 11707 3863 11757 3963
rect 11915 3863 11965 3963
rect 12123 3863 12173 3963
rect 12823 3822 12873 3922
rect 13031 3822 13081 3922
rect 13239 3822 13289 3922
rect 13452 3822 13502 3922
rect 16550 3904 16600 4004
rect 16763 3904 16813 4004
rect 16971 3904 17021 4004
rect 17179 3904 17229 4004
rect 17879 3863 17929 3963
rect 18087 3863 18137 3963
rect 18295 3863 18345 3963
rect 18508 3863 18558 3963
rect 385 3591 435 3691
rect 598 3591 648 3691
rect 806 3591 856 3691
rect 1014 3591 1064 3691
rect 3872 3535 3922 3635
rect 4080 3535 4130 3635
rect 4288 3535 4338 3635
rect 4501 3535 4551 3635
rect 5441 3632 5491 3732
rect 5654 3632 5704 3732
rect 5862 3632 5912 3732
rect 6070 3632 6120 3732
rect 8928 3576 8978 3676
rect 9136 3576 9186 3676
rect 9344 3576 9394 3676
rect 9557 3576 9607 3676
rect 10416 3596 10466 3696
rect 10629 3596 10679 3696
rect 10837 3596 10887 3696
rect 11045 3596 11095 3696
rect 1323 3347 1373 3447
rect 1536 3347 1586 3447
rect 1744 3347 1794 3447
rect 1952 3347 2002 3447
rect 2933 3225 2983 3325
rect 3141 3225 3191 3325
rect 3349 3225 3399 3325
rect 3562 3225 3612 3325
rect 6379 3388 6429 3488
rect 6592 3388 6642 3488
rect 6800 3388 6850 3488
rect 7008 3388 7058 3488
rect 13903 3540 13953 3640
rect 14111 3540 14161 3640
rect 14319 3540 14369 3640
rect 14532 3540 14582 3640
rect 15472 3637 15522 3737
rect 15685 3637 15735 3737
rect 15893 3637 15943 3737
rect 16101 3637 16151 3737
rect 18959 3581 19009 3681
rect 19167 3581 19217 3681
rect 19375 3581 19425 3681
rect 19588 3581 19638 3681
rect 7989 3266 8039 3366
rect 8197 3266 8247 3366
rect 8405 3266 8455 3366
rect 8618 3266 8668 3366
rect 11354 3352 11404 3452
rect 11567 3352 11617 3452
rect 11775 3352 11825 3452
rect 11983 3352 12033 3452
rect 384 3037 434 3137
rect 597 3037 647 3137
rect 805 3037 855 3137
rect 1013 3037 1063 3137
rect 3871 2981 3921 3081
rect 4079 2981 4129 3081
rect 4287 2981 4337 3081
rect 4500 2981 4550 3081
rect 5440 3078 5490 3178
rect 5653 3078 5703 3178
rect 5861 3078 5911 3178
rect 6069 3078 6119 3178
rect 12964 3230 13014 3330
rect 13172 3230 13222 3330
rect 13380 3230 13430 3330
rect 13593 3230 13643 3330
rect 16410 3393 16460 3493
rect 16623 3393 16673 3493
rect 16831 3393 16881 3493
rect 17039 3393 17089 3493
rect 18020 3271 18070 3371
rect 18228 3271 18278 3371
rect 18436 3271 18486 3371
rect 18649 3271 18699 3371
rect 8927 3022 8977 3122
rect 9135 3022 9185 3122
rect 9343 3022 9393 3122
rect 9556 3022 9606 3122
rect 10415 3042 10465 3142
rect 10628 3042 10678 3142
rect 10836 3042 10886 3142
rect 11044 3042 11094 3142
rect 13902 2986 13952 3086
rect 14110 2986 14160 3086
rect 14318 2986 14368 3086
rect 14531 2986 14581 3086
rect 15471 3083 15521 3183
rect 15684 3083 15734 3183
rect 15892 3083 15942 3183
rect 16100 3083 16150 3183
rect 18958 3027 19008 3127
rect 19166 3027 19216 3127
rect 19374 3027 19424 3127
rect 19587 3027 19637 3127
rect 1433 2768 1483 2868
rect 1646 2768 1696 2868
rect 1854 2768 1904 2868
rect 2062 2768 2112 2868
rect 6489 2809 6539 2909
rect 6702 2809 6752 2909
rect 6910 2809 6960 2909
rect 7118 2809 7168 2909
rect 2823 2701 2873 2801
rect 3031 2701 3081 2801
rect 3239 2701 3289 2801
rect 3452 2701 3502 2801
rect 7879 2742 7929 2842
rect 8087 2742 8137 2842
rect 8295 2742 8345 2842
rect 8508 2742 8558 2842
rect 11464 2773 11514 2873
rect 11677 2773 11727 2873
rect 11885 2773 11935 2873
rect 12093 2773 12143 2873
rect 16520 2814 16570 2914
rect 16733 2814 16783 2914
rect 16941 2814 16991 2914
rect 17149 2814 17199 2914
rect 12854 2706 12904 2806
rect 13062 2706 13112 2806
rect 13270 2706 13320 2806
rect 13483 2706 13533 2806
rect 17910 2747 17960 2847
rect 18118 2747 18168 2847
rect 18326 2747 18376 2847
rect 18539 2747 18589 2847
rect 385 2488 435 2588
rect 598 2488 648 2588
rect 806 2488 856 2588
rect 1014 2488 1064 2588
rect 3872 2432 3922 2532
rect 4080 2432 4130 2532
rect 4288 2432 4338 2532
rect 4501 2432 4551 2532
rect 5441 2529 5491 2629
rect 5654 2529 5704 2629
rect 5862 2529 5912 2629
rect 6070 2529 6120 2629
rect 8928 2473 8978 2573
rect 9136 2473 9186 2573
rect 9344 2473 9394 2573
rect 9557 2473 9607 2573
rect 10416 2493 10466 2593
rect 10629 2493 10679 2593
rect 10837 2493 10887 2593
rect 11045 2493 11095 2593
rect 1323 2244 1373 2344
rect 1536 2244 1586 2344
rect 1744 2244 1794 2344
rect 1952 2244 2002 2344
rect 2933 2122 2983 2222
rect 3141 2122 3191 2222
rect 3349 2122 3399 2222
rect 3562 2122 3612 2222
rect 6379 2285 6429 2385
rect 6592 2285 6642 2385
rect 6800 2285 6850 2385
rect 7008 2285 7058 2385
rect 13903 2437 13953 2537
rect 14111 2437 14161 2537
rect 14319 2437 14369 2537
rect 14532 2437 14582 2537
rect 15472 2534 15522 2634
rect 15685 2534 15735 2634
rect 15893 2534 15943 2634
rect 16101 2534 16151 2634
rect 18959 2478 19009 2578
rect 19167 2478 19217 2578
rect 19375 2478 19425 2578
rect 19588 2478 19638 2578
rect 7989 2163 8039 2263
rect 8197 2163 8247 2263
rect 8405 2163 8455 2263
rect 8618 2163 8668 2263
rect 11354 2249 11404 2349
rect 11567 2249 11617 2349
rect 11775 2249 11825 2349
rect 11983 2249 12033 2349
rect 384 1934 434 2034
rect 597 1934 647 2034
rect 805 1934 855 2034
rect 1013 1934 1063 2034
rect 3871 1878 3921 1978
rect 4079 1878 4129 1978
rect 4287 1878 4337 1978
rect 4500 1878 4550 1978
rect 5440 1975 5490 2075
rect 5653 1975 5703 2075
rect 5861 1975 5911 2075
rect 6069 1975 6119 2075
rect 12964 2127 13014 2227
rect 13172 2127 13222 2227
rect 13380 2127 13430 2227
rect 13593 2127 13643 2227
rect 16410 2290 16460 2390
rect 16623 2290 16673 2390
rect 16831 2290 16881 2390
rect 17039 2290 17089 2390
rect 18020 2168 18070 2268
rect 18228 2168 18278 2268
rect 18436 2168 18486 2268
rect 18649 2168 18699 2268
rect 8927 1919 8977 2019
rect 9135 1919 9185 2019
rect 9343 1919 9393 2019
rect 9556 1919 9606 2019
rect 10415 1939 10465 2039
rect 10628 1939 10678 2039
rect 10836 1939 10886 2039
rect 11044 1939 11094 2039
rect 13902 1883 13952 1983
rect 14110 1883 14160 1983
rect 14318 1883 14368 1983
rect 14531 1883 14581 1983
rect 15471 1980 15521 2080
rect 15684 1980 15734 2080
rect 15892 1980 15942 2080
rect 16100 1980 16150 2080
rect 18958 1924 19008 2024
rect 19166 1924 19216 2024
rect 19374 1924 19424 2024
rect 19587 1924 19637 2024
rect 1464 1652 1514 1752
rect 1677 1652 1727 1752
rect 1885 1652 1935 1752
rect 2093 1652 2143 1752
rect 2793 1611 2843 1711
rect 3001 1611 3051 1711
rect 3209 1611 3259 1711
rect 3422 1611 3472 1711
rect 6520 1693 6570 1793
rect 6733 1693 6783 1793
rect 6941 1693 6991 1793
rect 7149 1693 7199 1793
rect 7849 1652 7899 1752
rect 8057 1652 8107 1752
rect 8265 1652 8315 1752
rect 8478 1652 8528 1752
rect 11495 1657 11545 1757
rect 11708 1657 11758 1757
rect 11916 1657 11966 1757
rect 12124 1657 12174 1757
rect 12824 1616 12874 1716
rect 13032 1616 13082 1716
rect 13240 1616 13290 1716
rect 13453 1616 13503 1716
rect 16551 1698 16601 1798
rect 16764 1698 16814 1798
rect 16972 1698 17022 1798
rect 17180 1698 17230 1798
rect 17880 1657 17930 1757
rect 18088 1657 18138 1757
rect 18296 1657 18346 1757
rect 18509 1657 18559 1757
rect 386 1385 436 1485
rect 599 1385 649 1485
rect 807 1385 857 1485
rect 1015 1385 1065 1485
rect 3873 1329 3923 1429
rect 4081 1329 4131 1429
rect 4289 1329 4339 1429
rect 4502 1329 4552 1429
rect 5442 1426 5492 1526
rect 5655 1426 5705 1526
rect 5863 1426 5913 1526
rect 6071 1426 6121 1526
rect 8929 1370 8979 1470
rect 9137 1370 9187 1470
rect 9345 1370 9395 1470
rect 9558 1370 9608 1470
rect 10417 1390 10467 1490
rect 10630 1390 10680 1490
rect 10838 1390 10888 1490
rect 11046 1390 11096 1490
rect 1324 1141 1374 1241
rect 1537 1141 1587 1241
rect 1745 1141 1795 1241
rect 1953 1141 2003 1241
rect 2934 1019 2984 1119
rect 3142 1019 3192 1119
rect 3350 1019 3400 1119
rect 3563 1019 3613 1119
rect 6380 1182 6430 1282
rect 6593 1182 6643 1282
rect 6801 1182 6851 1282
rect 7009 1182 7059 1282
rect 13904 1334 13954 1434
rect 14112 1334 14162 1434
rect 14320 1334 14370 1434
rect 14533 1334 14583 1434
rect 15473 1431 15523 1531
rect 15686 1431 15736 1531
rect 15894 1431 15944 1531
rect 16102 1431 16152 1531
rect 18960 1375 19010 1475
rect 19168 1375 19218 1475
rect 19376 1375 19426 1475
rect 19589 1375 19639 1475
rect 7990 1060 8040 1160
rect 8198 1060 8248 1160
rect 8406 1060 8456 1160
rect 8619 1060 8669 1160
rect 11355 1146 11405 1246
rect 11568 1146 11618 1246
rect 11776 1146 11826 1246
rect 11984 1146 12034 1246
rect 385 831 435 931
rect 598 831 648 931
rect 806 831 856 931
rect 1014 831 1064 931
rect 3872 775 3922 875
rect 4080 775 4130 875
rect 4288 775 4338 875
rect 4501 775 4551 875
rect 5441 872 5491 972
rect 5654 872 5704 972
rect 5862 872 5912 972
rect 6070 872 6120 972
rect 12965 1024 13015 1124
rect 13173 1024 13223 1124
rect 13381 1024 13431 1124
rect 13594 1024 13644 1124
rect 16411 1187 16461 1287
rect 16624 1187 16674 1287
rect 16832 1187 16882 1287
rect 17040 1187 17090 1287
rect 18021 1065 18071 1165
rect 18229 1065 18279 1165
rect 18437 1065 18487 1165
rect 18650 1065 18700 1165
rect 8928 816 8978 916
rect 9136 816 9186 916
rect 9344 816 9394 916
rect 9557 816 9607 916
rect 10416 836 10466 936
rect 10629 836 10679 936
rect 10837 836 10887 936
rect 11045 836 11095 936
rect 13903 780 13953 880
rect 14111 780 14161 880
rect 14319 780 14369 880
rect 14532 780 14582 880
rect 15472 877 15522 977
rect 15685 877 15735 977
rect 15893 877 15943 977
rect 16101 877 16151 977
rect 18959 821 19009 921
rect 19167 821 19217 921
rect 19375 821 19425 921
rect 19588 821 19638 921
rect 1632 272 1682 372
rect 1845 272 1895 372
rect 2053 272 2103 372
rect 2261 272 2311 372
rect 4582 252 4632 352
rect 4795 252 4845 352
rect 5003 252 5053 352
rect 5211 252 5261 352
rect 6688 313 6738 413
rect 6901 313 6951 413
rect 7109 313 7159 413
rect 7317 313 7367 413
rect 11663 277 11713 377
rect 11876 277 11926 377
rect 12084 277 12134 377
rect 12292 277 12342 377
rect 9516 136 9566 236
rect 9729 136 9779 236
rect 9937 136 9987 236
rect 10145 136 10195 236
rect 14613 257 14663 357
rect 14826 257 14876 357
rect 15034 257 15084 357
rect 15242 257 15292 357
rect 16719 318 16769 418
rect 16932 318 16982 418
rect 17140 318 17190 418
rect 17348 318 17398 418
<< ndiff >>
rect 3820 9257 3869 9269
rect 3820 9237 3831 9257
rect 3851 9237 3869 9257
rect 3820 9227 3869 9237
rect 3919 9253 3963 9269
rect 3919 9233 3934 9253
rect 3954 9233 3963 9253
rect 3919 9227 3963 9233
rect 4033 9253 4077 9269
rect 4033 9233 4042 9253
rect 4062 9233 4077 9253
rect 4033 9227 4077 9233
rect 4127 9257 4176 9269
rect 4127 9237 4145 9257
rect 4165 9237 4176 9257
rect 4127 9227 4176 9237
rect 4241 9253 4285 9269
rect 4241 9233 4250 9253
rect 4270 9233 4285 9253
rect 4241 9227 4285 9233
rect 4335 9257 4384 9269
rect 4335 9237 4353 9257
rect 4373 9237 4384 9257
rect 4335 9227 4384 9237
rect 4454 9253 4498 9269
rect 4454 9233 4463 9253
rect 4483 9233 4498 9253
rect 4454 9227 4498 9233
rect 4548 9257 4597 9269
rect 8876 9298 8925 9310
rect 8876 9278 8887 9298
rect 8907 9278 8925 9298
rect 8876 9268 8925 9278
rect 8975 9294 9019 9310
rect 8975 9274 8990 9294
rect 9010 9274 9019 9294
rect 8975 9268 9019 9274
rect 9089 9294 9133 9310
rect 9089 9274 9098 9294
rect 9118 9274 9133 9294
rect 9089 9268 9133 9274
rect 9183 9298 9232 9310
rect 9183 9278 9201 9298
rect 9221 9278 9232 9298
rect 9183 9268 9232 9278
rect 9297 9294 9341 9310
rect 9297 9274 9306 9294
rect 9326 9274 9341 9294
rect 9297 9268 9341 9274
rect 9391 9298 9440 9310
rect 9391 9278 9409 9298
rect 9429 9278 9440 9298
rect 9391 9268 9440 9278
rect 9510 9294 9554 9310
rect 9510 9274 9519 9294
rect 9539 9274 9554 9294
rect 9510 9268 9554 9274
rect 9604 9298 9653 9310
rect 9604 9278 9622 9298
rect 9642 9278 9653 9298
rect 9604 9268 9653 9278
rect 4548 9237 4566 9257
rect 4586 9237 4597 9257
rect 4548 9227 4597 9237
rect 333 9019 382 9029
rect 333 8999 344 9019
rect 364 8999 382 9019
rect 333 8987 382 8999
rect 432 9023 476 9029
rect 432 9003 447 9023
rect 467 9003 476 9023
rect 432 8987 476 9003
rect 546 9019 595 9029
rect 546 8999 557 9019
rect 577 8999 595 9019
rect 546 8987 595 8999
rect 645 9023 689 9029
rect 645 9003 660 9023
rect 680 9003 689 9023
rect 645 8987 689 9003
rect 754 9019 803 9029
rect 754 8999 765 9019
rect 785 8999 803 9019
rect 754 8987 803 8999
rect 853 9023 897 9029
rect 853 9003 868 9023
rect 888 9003 897 9023
rect 853 8987 897 9003
rect 967 9023 1011 9029
rect 967 9003 976 9023
rect 996 9003 1011 9023
rect 967 8987 1011 9003
rect 1061 9019 1110 9029
rect 1061 8999 1079 9019
rect 1099 8999 1110 9019
rect 1061 8987 1110 8999
rect 13851 9262 13900 9274
rect 13851 9242 13862 9262
rect 13882 9242 13900 9262
rect 13851 9232 13900 9242
rect 13950 9258 13994 9274
rect 13950 9238 13965 9258
rect 13985 9238 13994 9258
rect 13950 9232 13994 9238
rect 14064 9258 14108 9274
rect 14064 9238 14073 9258
rect 14093 9238 14108 9258
rect 14064 9232 14108 9238
rect 14158 9262 14207 9274
rect 14158 9242 14176 9262
rect 14196 9242 14207 9262
rect 14158 9232 14207 9242
rect 14272 9258 14316 9274
rect 14272 9238 14281 9258
rect 14301 9238 14316 9258
rect 14272 9232 14316 9238
rect 14366 9262 14415 9274
rect 14366 9242 14384 9262
rect 14404 9242 14415 9262
rect 14366 9232 14415 9242
rect 14485 9258 14529 9274
rect 14485 9238 14494 9258
rect 14514 9238 14529 9258
rect 14485 9232 14529 9238
rect 14579 9262 14628 9274
rect 18907 9303 18956 9315
rect 18907 9283 18918 9303
rect 18938 9283 18956 9303
rect 18907 9273 18956 9283
rect 19006 9299 19050 9315
rect 19006 9279 19021 9299
rect 19041 9279 19050 9299
rect 19006 9273 19050 9279
rect 19120 9299 19164 9315
rect 19120 9279 19129 9299
rect 19149 9279 19164 9299
rect 19120 9273 19164 9279
rect 19214 9303 19263 9315
rect 19214 9283 19232 9303
rect 19252 9283 19263 9303
rect 19214 9273 19263 9283
rect 19328 9299 19372 9315
rect 19328 9279 19337 9299
rect 19357 9279 19372 9299
rect 19328 9273 19372 9279
rect 19422 9303 19471 9315
rect 19422 9283 19440 9303
rect 19460 9283 19471 9303
rect 19422 9273 19471 9283
rect 19541 9299 19585 9315
rect 19541 9279 19550 9299
rect 19570 9279 19585 9299
rect 19541 9273 19585 9279
rect 19635 9303 19684 9315
rect 19635 9283 19653 9303
rect 19673 9283 19684 9303
rect 19635 9273 19684 9283
rect 14579 9242 14597 9262
rect 14617 9242 14628 9262
rect 14579 9232 14628 9242
rect 5389 9060 5438 9070
rect 5389 9040 5400 9060
rect 5420 9040 5438 9060
rect 5389 9028 5438 9040
rect 5488 9064 5532 9070
rect 5488 9044 5503 9064
rect 5523 9044 5532 9064
rect 5488 9028 5532 9044
rect 5602 9060 5651 9070
rect 5602 9040 5613 9060
rect 5633 9040 5651 9060
rect 5602 9028 5651 9040
rect 5701 9064 5745 9070
rect 5701 9044 5716 9064
rect 5736 9044 5745 9064
rect 5701 9028 5745 9044
rect 5810 9060 5859 9070
rect 5810 9040 5821 9060
rect 5841 9040 5859 9060
rect 5810 9028 5859 9040
rect 5909 9064 5953 9070
rect 5909 9044 5924 9064
rect 5944 9044 5953 9064
rect 5909 9028 5953 9044
rect 6023 9064 6067 9070
rect 6023 9044 6032 9064
rect 6052 9044 6067 9064
rect 6023 9028 6067 9044
rect 6117 9060 6166 9070
rect 6117 9040 6135 9060
rect 6155 9040 6166 9060
rect 6117 9028 6166 9040
rect 2881 8947 2930 8959
rect 2881 8927 2892 8947
rect 2912 8927 2930 8947
rect 2881 8917 2930 8927
rect 2980 8943 3024 8959
rect 2980 8923 2995 8943
rect 3015 8923 3024 8943
rect 2980 8917 3024 8923
rect 3094 8943 3138 8959
rect 3094 8923 3103 8943
rect 3123 8923 3138 8943
rect 3094 8917 3138 8923
rect 3188 8947 3237 8959
rect 3188 8927 3206 8947
rect 3226 8927 3237 8947
rect 3188 8917 3237 8927
rect 3302 8943 3346 8959
rect 3302 8923 3311 8943
rect 3331 8923 3346 8943
rect 3302 8917 3346 8923
rect 3396 8947 3445 8959
rect 3396 8927 3414 8947
rect 3434 8927 3445 8947
rect 3396 8917 3445 8927
rect 3515 8943 3559 8959
rect 3515 8923 3524 8943
rect 3544 8923 3559 8943
rect 3515 8917 3559 8923
rect 3609 8947 3658 8959
rect 3609 8927 3627 8947
rect 3647 8927 3658 8947
rect 3609 8917 3658 8927
rect 1271 8775 1320 8785
rect 1271 8755 1282 8775
rect 1302 8755 1320 8775
rect 1271 8743 1320 8755
rect 1370 8779 1414 8785
rect 1370 8759 1385 8779
rect 1405 8759 1414 8779
rect 1370 8743 1414 8759
rect 1484 8775 1533 8785
rect 1484 8755 1495 8775
rect 1515 8755 1533 8775
rect 1484 8743 1533 8755
rect 1583 8779 1627 8785
rect 1583 8759 1598 8779
rect 1618 8759 1627 8779
rect 1583 8743 1627 8759
rect 1692 8775 1741 8785
rect 1692 8755 1703 8775
rect 1723 8755 1741 8775
rect 1692 8743 1741 8755
rect 1791 8779 1835 8785
rect 1791 8759 1806 8779
rect 1826 8759 1835 8779
rect 1791 8743 1835 8759
rect 1905 8779 1949 8785
rect 1905 8759 1914 8779
rect 1934 8759 1949 8779
rect 1905 8743 1949 8759
rect 1999 8775 2048 8785
rect 1999 8755 2017 8775
rect 2037 8755 2048 8775
rect 1999 8743 2048 8755
rect 7937 8988 7986 9000
rect 7937 8968 7948 8988
rect 7968 8968 7986 8988
rect 7937 8958 7986 8968
rect 8036 8984 8080 9000
rect 8036 8964 8051 8984
rect 8071 8964 8080 8984
rect 8036 8958 8080 8964
rect 8150 8984 8194 9000
rect 8150 8964 8159 8984
rect 8179 8964 8194 8984
rect 8150 8958 8194 8964
rect 8244 8988 8293 9000
rect 8244 8968 8262 8988
rect 8282 8968 8293 8988
rect 8244 8958 8293 8968
rect 8358 8984 8402 9000
rect 8358 8964 8367 8984
rect 8387 8964 8402 8984
rect 8358 8958 8402 8964
rect 8452 8988 8501 9000
rect 8452 8968 8470 8988
rect 8490 8968 8501 8988
rect 8452 8958 8501 8968
rect 8571 8984 8615 9000
rect 8571 8964 8580 8984
rect 8600 8964 8615 8984
rect 8571 8958 8615 8964
rect 8665 8988 8714 9000
rect 8665 8968 8683 8988
rect 8703 8968 8714 8988
rect 8665 8958 8714 8968
rect 10364 9024 10413 9034
rect 10364 9004 10375 9024
rect 10395 9004 10413 9024
rect 10364 8992 10413 9004
rect 10463 9028 10507 9034
rect 10463 9008 10478 9028
rect 10498 9008 10507 9028
rect 10463 8992 10507 9008
rect 10577 9024 10626 9034
rect 10577 9004 10588 9024
rect 10608 9004 10626 9024
rect 10577 8992 10626 9004
rect 10676 9028 10720 9034
rect 10676 9008 10691 9028
rect 10711 9008 10720 9028
rect 10676 8992 10720 9008
rect 10785 9024 10834 9034
rect 10785 9004 10796 9024
rect 10816 9004 10834 9024
rect 10785 8992 10834 9004
rect 10884 9028 10928 9034
rect 10884 9008 10899 9028
rect 10919 9008 10928 9028
rect 10884 8992 10928 9008
rect 10998 9028 11042 9034
rect 10998 9008 11007 9028
rect 11027 9008 11042 9028
rect 10998 8992 11042 9008
rect 11092 9024 11141 9034
rect 11092 9004 11110 9024
rect 11130 9004 11141 9024
rect 11092 8992 11141 9004
rect 15420 9065 15469 9075
rect 15420 9045 15431 9065
rect 15451 9045 15469 9065
rect 15420 9033 15469 9045
rect 15519 9069 15563 9075
rect 15519 9049 15534 9069
rect 15554 9049 15563 9069
rect 15519 9033 15563 9049
rect 15633 9065 15682 9075
rect 15633 9045 15644 9065
rect 15664 9045 15682 9065
rect 15633 9033 15682 9045
rect 15732 9069 15776 9075
rect 15732 9049 15747 9069
rect 15767 9049 15776 9069
rect 15732 9033 15776 9049
rect 15841 9065 15890 9075
rect 15841 9045 15852 9065
rect 15872 9045 15890 9065
rect 15841 9033 15890 9045
rect 15940 9069 15984 9075
rect 15940 9049 15955 9069
rect 15975 9049 15984 9069
rect 15940 9033 15984 9049
rect 16054 9069 16098 9075
rect 16054 9049 16063 9069
rect 16083 9049 16098 9069
rect 16054 9033 16098 9049
rect 16148 9065 16197 9075
rect 16148 9045 16166 9065
rect 16186 9045 16197 9065
rect 16148 9033 16197 9045
rect 6327 8816 6376 8826
rect 6327 8796 6338 8816
rect 6358 8796 6376 8816
rect 6327 8784 6376 8796
rect 6426 8820 6470 8826
rect 6426 8800 6441 8820
rect 6461 8800 6470 8820
rect 6426 8784 6470 8800
rect 6540 8816 6589 8826
rect 6540 8796 6551 8816
rect 6571 8796 6589 8816
rect 6540 8784 6589 8796
rect 6639 8820 6683 8826
rect 6639 8800 6654 8820
rect 6674 8800 6683 8820
rect 6639 8784 6683 8800
rect 6748 8816 6797 8826
rect 6748 8796 6759 8816
rect 6779 8796 6797 8816
rect 6748 8784 6797 8796
rect 6847 8820 6891 8826
rect 6847 8800 6862 8820
rect 6882 8800 6891 8820
rect 6847 8784 6891 8800
rect 6961 8820 7005 8826
rect 6961 8800 6970 8820
rect 6990 8800 7005 8820
rect 6961 8784 7005 8800
rect 7055 8816 7104 8826
rect 7055 8796 7073 8816
rect 7093 8796 7104 8816
rect 7055 8784 7104 8796
rect 12912 8952 12961 8964
rect 12912 8932 12923 8952
rect 12943 8932 12961 8952
rect 12912 8922 12961 8932
rect 13011 8948 13055 8964
rect 13011 8928 13026 8948
rect 13046 8928 13055 8948
rect 13011 8922 13055 8928
rect 13125 8948 13169 8964
rect 13125 8928 13134 8948
rect 13154 8928 13169 8948
rect 13125 8922 13169 8928
rect 13219 8952 13268 8964
rect 13219 8932 13237 8952
rect 13257 8932 13268 8952
rect 13219 8922 13268 8932
rect 13333 8948 13377 8964
rect 13333 8928 13342 8948
rect 13362 8928 13377 8948
rect 13333 8922 13377 8928
rect 13427 8952 13476 8964
rect 13427 8932 13445 8952
rect 13465 8932 13476 8952
rect 13427 8922 13476 8932
rect 13546 8948 13590 8964
rect 13546 8928 13555 8948
rect 13575 8928 13590 8948
rect 13546 8922 13590 8928
rect 13640 8952 13689 8964
rect 13640 8932 13658 8952
rect 13678 8932 13689 8952
rect 13640 8922 13689 8932
rect 3819 8703 3868 8715
rect 3819 8683 3830 8703
rect 3850 8683 3868 8703
rect 3819 8673 3868 8683
rect 3918 8699 3962 8715
rect 3918 8679 3933 8699
rect 3953 8679 3962 8699
rect 3918 8673 3962 8679
rect 4032 8699 4076 8715
rect 4032 8679 4041 8699
rect 4061 8679 4076 8699
rect 4032 8673 4076 8679
rect 4126 8703 4175 8715
rect 4126 8683 4144 8703
rect 4164 8683 4175 8703
rect 4126 8673 4175 8683
rect 4240 8699 4284 8715
rect 4240 8679 4249 8699
rect 4269 8679 4284 8699
rect 4240 8673 4284 8679
rect 4334 8703 4383 8715
rect 4334 8683 4352 8703
rect 4372 8683 4383 8703
rect 4334 8673 4383 8683
rect 4453 8699 4497 8715
rect 4453 8679 4462 8699
rect 4482 8679 4497 8699
rect 4453 8673 4497 8679
rect 4547 8703 4596 8715
rect 4547 8683 4565 8703
rect 4585 8683 4596 8703
rect 4547 8673 4596 8683
rect 8875 8744 8924 8756
rect 8875 8724 8886 8744
rect 8906 8724 8924 8744
rect 8875 8714 8924 8724
rect 8974 8740 9018 8756
rect 8974 8720 8989 8740
rect 9009 8720 9018 8740
rect 8974 8714 9018 8720
rect 9088 8740 9132 8756
rect 9088 8720 9097 8740
rect 9117 8720 9132 8740
rect 9088 8714 9132 8720
rect 9182 8744 9231 8756
rect 9182 8724 9200 8744
rect 9220 8724 9231 8744
rect 9182 8714 9231 8724
rect 9296 8740 9340 8756
rect 9296 8720 9305 8740
rect 9325 8720 9340 8740
rect 9296 8714 9340 8720
rect 9390 8744 9439 8756
rect 9390 8724 9408 8744
rect 9428 8724 9439 8744
rect 9390 8714 9439 8724
rect 9509 8740 9553 8756
rect 9509 8720 9518 8740
rect 9538 8720 9553 8740
rect 9509 8714 9553 8720
rect 9603 8744 9652 8756
rect 9603 8724 9621 8744
rect 9641 8724 9652 8744
rect 9603 8714 9652 8724
rect 11302 8780 11351 8790
rect 11302 8760 11313 8780
rect 11333 8760 11351 8780
rect 11302 8748 11351 8760
rect 11401 8784 11445 8790
rect 11401 8764 11416 8784
rect 11436 8764 11445 8784
rect 11401 8748 11445 8764
rect 11515 8780 11564 8790
rect 11515 8760 11526 8780
rect 11546 8760 11564 8780
rect 11515 8748 11564 8760
rect 11614 8784 11658 8790
rect 11614 8764 11629 8784
rect 11649 8764 11658 8784
rect 11614 8748 11658 8764
rect 11723 8780 11772 8790
rect 11723 8760 11734 8780
rect 11754 8760 11772 8780
rect 11723 8748 11772 8760
rect 11822 8784 11866 8790
rect 11822 8764 11837 8784
rect 11857 8764 11866 8784
rect 11822 8748 11866 8764
rect 11936 8784 11980 8790
rect 11936 8764 11945 8784
rect 11965 8764 11980 8784
rect 11936 8748 11980 8764
rect 12030 8780 12079 8790
rect 12030 8760 12048 8780
rect 12068 8760 12079 8780
rect 12030 8748 12079 8760
rect 17968 8993 18017 9005
rect 17968 8973 17979 8993
rect 17999 8973 18017 8993
rect 17968 8963 18017 8973
rect 18067 8989 18111 9005
rect 18067 8969 18082 8989
rect 18102 8969 18111 8989
rect 18067 8963 18111 8969
rect 18181 8989 18225 9005
rect 18181 8969 18190 8989
rect 18210 8969 18225 8989
rect 18181 8963 18225 8969
rect 18275 8993 18324 9005
rect 18275 8973 18293 8993
rect 18313 8973 18324 8993
rect 18275 8963 18324 8973
rect 18389 8989 18433 9005
rect 18389 8969 18398 8989
rect 18418 8969 18433 8989
rect 18389 8963 18433 8969
rect 18483 8993 18532 9005
rect 18483 8973 18501 8993
rect 18521 8973 18532 8993
rect 18483 8963 18532 8973
rect 18602 8989 18646 9005
rect 18602 8969 18611 8989
rect 18631 8969 18646 8989
rect 18602 8963 18646 8969
rect 18696 8993 18745 9005
rect 18696 8973 18714 8993
rect 18734 8973 18745 8993
rect 18696 8963 18745 8973
rect 16358 8821 16407 8831
rect 16358 8801 16369 8821
rect 16389 8801 16407 8821
rect 16358 8789 16407 8801
rect 16457 8825 16501 8831
rect 16457 8805 16472 8825
rect 16492 8805 16501 8825
rect 16457 8789 16501 8805
rect 16571 8821 16620 8831
rect 16571 8801 16582 8821
rect 16602 8801 16620 8821
rect 16571 8789 16620 8801
rect 16670 8825 16714 8831
rect 16670 8805 16685 8825
rect 16705 8805 16714 8825
rect 16670 8789 16714 8805
rect 16779 8821 16828 8831
rect 16779 8801 16790 8821
rect 16810 8801 16828 8821
rect 16779 8789 16828 8801
rect 16878 8825 16922 8831
rect 16878 8805 16893 8825
rect 16913 8805 16922 8825
rect 16878 8789 16922 8805
rect 16992 8825 17036 8831
rect 16992 8805 17001 8825
rect 17021 8805 17036 8825
rect 16992 8789 17036 8805
rect 17086 8821 17135 8831
rect 17086 8801 17104 8821
rect 17124 8801 17135 8821
rect 17086 8789 17135 8801
rect 13850 8708 13899 8720
rect 13850 8688 13861 8708
rect 13881 8688 13899 8708
rect 13850 8678 13899 8688
rect 13949 8704 13993 8720
rect 13949 8684 13964 8704
rect 13984 8684 13993 8704
rect 13949 8678 13993 8684
rect 14063 8704 14107 8720
rect 14063 8684 14072 8704
rect 14092 8684 14107 8704
rect 14063 8678 14107 8684
rect 14157 8708 14206 8720
rect 14157 8688 14175 8708
rect 14195 8688 14206 8708
rect 14157 8678 14206 8688
rect 14271 8704 14315 8720
rect 14271 8684 14280 8704
rect 14300 8684 14315 8704
rect 14271 8678 14315 8684
rect 14365 8708 14414 8720
rect 14365 8688 14383 8708
rect 14403 8688 14414 8708
rect 14365 8678 14414 8688
rect 14484 8704 14528 8720
rect 14484 8684 14493 8704
rect 14513 8684 14528 8704
rect 14484 8678 14528 8684
rect 14578 8708 14627 8720
rect 14578 8688 14596 8708
rect 14616 8688 14627 8708
rect 14578 8678 14627 8688
rect 5388 8506 5437 8516
rect 5388 8486 5399 8506
rect 5419 8486 5437 8506
rect 332 8465 381 8475
rect 332 8445 343 8465
rect 363 8445 381 8465
rect 332 8433 381 8445
rect 431 8469 475 8475
rect 431 8449 446 8469
rect 466 8449 475 8469
rect 431 8433 475 8449
rect 545 8465 594 8475
rect 545 8445 556 8465
rect 576 8445 594 8465
rect 545 8433 594 8445
rect 644 8469 688 8475
rect 644 8449 659 8469
rect 679 8449 688 8469
rect 644 8433 688 8449
rect 753 8465 802 8475
rect 753 8445 764 8465
rect 784 8445 802 8465
rect 753 8433 802 8445
rect 852 8469 896 8475
rect 852 8449 867 8469
rect 887 8449 896 8469
rect 852 8433 896 8449
rect 966 8469 1010 8475
rect 966 8449 975 8469
rect 995 8449 1010 8469
rect 966 8433 1010 8449
rect 1060 8465 1109 8475
rect 1060 8445 1078 8465
rect 1098 8445 1109 8465
rect 1060 8433 1109 8445
rect 2741 8436 2790 8448
rect 2741 8416 2752 8436
rect 2772 8416 2790 8436
rect 2741 8406 2790 8416
rect 2840 8432 2884 8448
rect 2840 8412 2855 8432
rect 2875 8412 2884 8432
rect 2840 8406 2884 8412
rect 2954 8432 2998 8448
rect 2954 8412 2963 8432
rect 2983 8412 2998 8432
rect 2954 8406 2998 8412
rect 3048 8436 3097 8448
rect 3048 8416 3066 8436
rect 3086 8416 3097 8436
rect 3048 8406 3097 8416
rect 3162 8432 3206 8448
rect 3162 8412 3171 8432
rect 3191 8412 3206 8432
rect 3162 8406 3206 8412
rect 3256 8436 3305 8448
rect 3256 8416 3274 8436
rect 3294 8416 3305 8436
rect 3256 8406 3305 8416
rect 3375 8432 3419 8448
rect 3375 8412 3384 8432
rect 3404 8412 3419 8432
rect 3375 8406 3419 8412
rect 3469 8436 3518 8448
rect 3469 8416 3487 8436
rect 3507 8416 3518 8436
rect 3469 8406 3518 8416
rect 5388 8474 5437 8486
rect 5487 8510 5531 8516
rect 5487 8490 5502 8510
rect 5522 8490 5531 8510
rect 5487 8474 5531 8490
rect 5601 8506 5650 8516
rect 5601 8486 5612 8506
rect 5632 8486 5650 8506
rect 5601 8474 5650 8486
rect 5700 8510 5744 8516
rect 5700 8490 5715 8510
rect 5735 8490 5744 8510
rect 5700 8474 5744 8490
rect 5809 8506 5858 8516
rect 5809 8486 5820 8506
rect 5840 8486 5858 8506
rect 5809 8474 5858 8486
rect 5908 8510 5952 8516
rect 5908 8490 5923 8510
rect 5943 8490 5952 8510
rect 5908 8474 5952 8490
rect 6022 8510 6066 8516
rect 6022 8490 6031 8510
rect 6051 8490 6066 8510
rect 6022 8474 6066 8490
rect 6116 8506 6165 8516
rect 6116 8486 6134 8506
rect 6154 8486 6165 8506
rect 6116 8474 6165 8486
rect 7797 8477 7846 8489
rect 7797 8457 7808 8477
rect 7828 8457 7846 8477
rect 7797 8447 7846 8457
rect 7896 8473 7940 8489
rect 7896 8453 7911 8473
rect 7931 8453 7940 8473
rect 7896 8447 7940 8453
rect 8010 8473 8054 8489
rect 8010 8453 8019 8473
rect 8039 8453 8054 8473
rect 8010 8447 8054 8453
rect 8104 8477 8153 8489
rect 8104 8457 8122 8477
rect 8142 8457 8153 8477
rect 8104 8447 8153 8457
rect 8218 8473 8262 8489
rect 8218 8453 8227 8473
rect 8247 8453 8262 8473
rect 8218 8447 8262 8453
rect 8312 8477 8361 8489
rect 8312 8457 8330 8477
rect 8350 8457 8361 8477
rect 8312 8447 8361 8457
rect 8431 8473 8475 8489
rect 8431 8453 8440 8473
rect 8460 8453 8475 8473
rect 8431 8447 8475 8453
rect 8525 8477 8574 8489
rect 8525 8457 8543 8477
rect 8563 8457 8574 8477
rect 8525 8447 8574 8457
rect 18906 8749 18955 8761
rect 18906 8729 18917 8749
rect 18937 8729 18955 8749
rect 18906 8719 18955 8729
rect 19005 8745 19049 8761
rect 19005 8725 19020 8745
rect 19040 8725 19049 8745
rect 19005 8719 19049 8725
rect 19119 8745 19163 8761
rect 19119 8725 19128 8745
rect 19148 8725 19163 8745
rect 19119 8719 19163 8725
rect 19213 8749 19262 8761
rect 19213 8729 19231 8749
rect 19251 8729 19262 8749
rect 19213 8719 19262 8729
rect 19327 8745 19371 8761
rect 19327 8725 19336 8745
rect 19356 8725 19371 8745
rect 19327 8719 19371 8725
rect 19421 8749 19470 8761
rect 19421 8729 19439 8749
rect 19459 8729 19470 8749
rect 19421 8719 19470 8729
rect 19540 8745 19584 8761
rect 19540 8725 19549 8745
rect 19569 8725 19584 8745
rect 19540 8719 19584 8725
rect 19634 8749 19683 8761
rect 19634 8729 19652 8749
rect 19672 8729 19683 8749
rect 19634 8719 19683 8729
rect 15419 8511 15468 8521
rect 15419 8491 15430 8511
rect 15450 8491 15468 8511
rect 10363 8470 10412 8480
rect 10363 8450 10374 8470
rect 10394 8450 10412 8470
rect 10363 8438 10412 8450
rect 10462 8474 10506 8480
rect 10462 8454 10477 8474
rect 10497 8454 10506 8474
rect 10462 8438 10506 8454
rect 10576 8470 10625 8480
rect 10576 8450 10587 8470
rect 10607 8450 10625 8470
rect 10576 8438 10625 8450
rect 10675 8474 10719 8480
rect 10675 8454 10690 8474
rect 10710 8454 10719 8474
rect 10675 8438 10719 8454
rect 10784 8470 10833 8480
rect 10784 8450 10795 8470
rect 10815 8450 10833 8470
rect 10784 8438 10833 8450
rect 10883 8474 10927 8480
rect 10883 8454 10898 8474
rect 10918 8454 10927 8474
rect 10883 8438 10927 8454
rect 10997 8474 11041 8480
rect 10997 8454 11006 8474
rect 11026 8454 11041 8474
rect 10997 8438 11041 8454
rect 11091 8470 11140 8480
rect 11091 8450 11109 8470
rect 11129 8450 11140 8470
rect 11091 8438 11140 8450
rect 12772 8441 12821 8453
rect 12772 8421 12783 8441
rect 12803 8421 12821 8441
rect 12772 8411 12821 8421
rect 12871 8437 12915 8453
rect 12871 8417 12886 8437
rect 12906 8417 12915 8437
rect 12871 8411 12915 8417
rect 12985 8437 13029 8453
rect 12985 8417 12994 8437
rect 13014 8417 13029 8437
rect 12985 8411 13029 8417
rect 13079 8441 13128 8453
rect 13079 8421 13097 8441
rect 13117 8421 13128 8441
rect 13079 8411 13128 8421
rect 13193 8437 13237 8453
rect 13193 8417 13202 8437
rect 13222 8417 13237 8437
rect 13193 8411 13237 8417
rect 13287 8441 13336 8453
rect 13287 8421 13305 8441
rect 13325 8421 13336 8441
rect 13287 8411 13336 8421
rect 13406 8437 13450 8453
rect 13406 8417 13415 8437
rect 13435 8417 13450 8437
rect 13406 8411 13450 8417
rect 13500 8441 13549 8453
rect 13500 8421 13518 8441
rect 13538 8421 13549 8441
rect 13500 8411 13549 8421
rect 15419 8479 15468 8491
rect 15518 8515 15562 8521
rect 15518 8495 15533 8515
rect 15553 8495 15562 8515
rect 15518 8479 15562 8495
rect 15632 8511 15681 8521
rect 15632 8491 15643 8511
rect 15663 8491 15681 8511
rect 15632 8479 15681 8491
rect 15731 8515 15775 8521
rect 15731 8495 15746 8515
rect 15766 8495 15775 8515
rect 15731 8479 15775 8495
rect 15840 8511 15889 8521
rect 15840 8491 15851 8511
rect 15871 8491 15889 8511
rect 15840 8479 15889 8491
rect 15939 8515 15983 8521
rect 15939 8495 15954 8515
rect 15974 8495 15983 8515
rect 15939 8479 15983 8495
rect 16053 8515 16097 8521
rect 16053 8495 16062 8515
rect 16082 8495 16097 8515
rect 16053 8479 16097 8495
rect 16147 8511 16196 8521
rect 16147 8491 16165 8511
rect 16185 8491 16196 8511
rect 16147 8479 16196 8491
rect 17828 8482 17877 8494
rect 17828 8462 17839 8482
rect 17859 8462 17877 8482
rect 17828 8452 17877 8462
rect 17927 8478 17971 8494
rect 17927 8458 17942 8478
rect 17962 8458 17971 8478
rect 17927 8452 17971 8458
rect 18041 8478 18085 8494
rect 18041 8458 18050 8478
rect 18070 8458 18085 8478
rect 18041 8452 18085 8458
rect 18135 8482 18184 8494
rect 18135 8462 18153 8482
rect 18173 8462 18184 8482
rect 18135 8452 18184 8462
rect 18249 8478 18293 8494
rect 18249 8458 18258 8478
rect 18278 8458 18293 8478
rect 18249 8452 18293 8458
rect 18343 8482 18392 8494
rect 18343 8462 18361 8482
rect 18381 8462 18392 8482
rect 18343 8452 18392 8462
rect 18462 8478 18506 8494
rect 18462 8458 18471 8478
rect 18491 8458 18506 8478
rect 18462 8452 18506 8458
rect 18556 8482 18605 8494
rect 18556 8462 18574 8482
rect 18594 8462 18605 8482
rect 18556 8452 18605 8462
rect 1412 8183 1461 8193
rect 1412 8163 1423 8183
rect 1443 8163 1461 8183
rect 1412 8151 1461 8163
rect 1511 8187 1555 8193
rect 1511 8167 1526 8187
rect 1546 8167 1555 8187
rect 1511 8151 1555 8167
rect 1625 8183 1674 8193
rect 1625 8163 1636 8183
rect 1656 8163 1674 8183
rect 1625 8151 1674 8163
rect 1724 8187 1768 8193
rect 1724 8167 1739 8187
rect 1759 8167 1768 8187
rect 1724 8151 1768 8167
rect 1833 8183 1882 8193
rect 1833 8163 1844 8183
rect 1864 8163 1882 8183
rect 1833 8151 1882 8163
rect 1932 8187 1976 8193
rect 1932 8167 1947 8187
rect 1967 8167 1976 8187
rect 1932 8151 1976 8167
rect 2046 8187 2090 8193
rect 2046 8167 2055 8187
rect 2075 8167 2090 8187
rect 2046 8151 2090 8167
rect 2140 8183 2189 8193
rect 2140 8163 2158 8183
rect 2178 8163 2189 8183
rect 2140 8151 2189 8163
rect 3821 8154 3870 8166
rect 3821 8134 3832 8154
rect 3852 8134 3870 8154
rect 3821 8124 3870 8134
rect 3920 8150 3964 8166
rect 3920 8130 3935 8150
rect 3955 8130 3964 8150
rect 3920 8124 3964 8130
rect 4034 8150 4078 8166
rect 4034 8130 4043 8150
rect 4063 8130 4078 8150
rect 4034 8124 4078 8130
rect 4128 8154 4177 8166
rect 4128 8134 4146 8154
rect 4166 8134 4177 8154
rect 4128 8124 4177 8134
rect 4242 8150 4286 8166
rect 4242 8130 4251 8150
rect 4271 8130 4286 8150
rect 4242 8124 4286 8130
rect 4336 8154 4385 8166
rect 4336 8134 4354 8154
rect 4374 8134 4385 8154
rect 4336 8124 4385 8134
rect 4455 8150 4499 8166
rect 4455 8130 4464 8150
rect 4484 8130 4499 8150
rect 4455 8124 4499 8130
rect 4549 8154 4598 8166
rect 6468 8224 6517 8234
rect 6468 8204 6479 8224
rect 6499 8204 6517 8224
rect 6468 8192 6517 8204
rect 6567 8228 6611 8234
rect 6567 8208 6582 8228
rect 6602 8208 6611 8228
rect 6567 8192 6611 8208
rect 6681 8224 6730 8234
rect 6681 8204 6692 8224
rect 6712 8204 6730 8224
rect 6681 8192 6730 8204
rect 6780 8228 6824 8234
rect 6780 8208 6795 8228
rect 6815 8208 6824 8228
rect 6780 8192 6824 8208
rect 6889 8224 6938 8234
rect 6889 8204 6900 8224
rect 6920 8204 6938 8224
rect 6889 8192 6938 8204
rect 6988 8228 7032 8234
rect 6988 8208 7003 8228
rect 7023 8208 7032 8228
rect 6988 8192 7032 8208
rect 7102 8228 7146 8234
rect 7102 8208 7111 8228
rect 7131 8208 7146 8228
rect 7102 8192 7146 8208
rect 7196 8224 7245 8234
rect 7196 8204 7214 8224
rect 7234 8204 7245 8224
rect 7196 8192 7245 8204
rect 8877 8195 8926 8207
rect 8877 8175 8888 8195
rect 8908 8175 8926 8195
rect 8877 8165 8926 8175
rect 8976 8191 9020 8207
rect 8976 8171 8991 8191
rect 9011 8171 9020 8191
rect 8976 8165 9020 8171
rect 9090 8191 9134 8207
rect 9090 8171 9099 8191
rect 9119 8171 9134 8191
rect 9090 8165 9134 8171
rect 9184 8195 9233 8207
rect 9184 8175 9202 8195
rect 9222 8175 9233 8195
rect 9184 8165 9233 8175
rect 9298 8191 9342 8207
rect 9298 8171 9307 8191
rect 9327 8171 9342 8191
rect 9298 8165 9342 8171
rect 9392 8195 9441 8207
rect 9392 8175 9410 8195
rect 9430 8175 9441 8195
rect 9392 8165 9441 8175
rect 9511 8191 9555 8207
rect 9511 8171 9520 8191
rect 9540 8171 9555 8191
rect 9511 8165 9555 8171
rect 9605 8195 9654 8207
rect 9605 8175 9623 8195
rect 9643 8175 9654 8195
rect 9605 8165 9654 8175
rect 4549 8134 4567 8154
rect 4587 8134 4598 8154
rect 4549 8124 4598 8134
rect 334 7916 383 7926
rect 334 7896 345 7916
rect 365 7896 383 7916
rect 334 7884 383 7896
rect 433 7920 477 7926
rect 433 7900 448 7920
rect 468 7900 477 7920
rect 433 7884 477 7900
rect 547 7916 596 7926
rect 547 7896 558 7916
rect 578 7896 596 7916
rect 547 7884 596 7896
rect 646 7920 690 7926
rect 646 7900 661 7920
rect 681 7900 690 7920
rect 646 7884 690 7900
rect 755 7916 804 7926
rect 755 7896 766 7916
rect 786 7896 804 7916
rect 755 7884 804 7896
rect 854 7920 898 7926
rect 854 7900 869 7920
rect 889 7900 898 7920
rect 854 7884 898 7900
rect 968 7920 1012 7926
rect 968 7900 977 7920
rect 997 7900 1012 7920
rect 968 7884 1012 7900
rect 1062 7916 1111 7926
rect 1062 7896 1080 7916
rect 1100 7896 1111 7916
rect 1062 7884 1111 7896
rect 11443 8188 11492 8198
rect 11443 8168 11454 8188
rect 11474 8168 11492 8188
rect 11443 8156 11492 8168
rect 11542 8192 11586 8198
rect 11542 8172 11557 8192
rect 11577 8172 11586 8192
rect 11542 8156 11586 8172
rect 11656 8188 11705 8198
rect 11656 8168 11667 8188
rect 11687 8168 11705 8188
rect 11656 8156 11705 8168
rect 11755 8192 11799 8198
rect 11755 8172 11770 8192
rect 11790 8172 11799 8192
rect 11755 8156 11799 8172
rect 11864 8188 11913 8198
rect 11864 8168 11875 8188
rect 11895 8168 11913 8188
rect 11864 8156 11913 8168
rect 11963 8192 12007 8198
rect 11963 8172 11978 8192
rect 11998 8172 12007 8192
rect 11963 8156 12007 8172
rect 12077 8192 12121 8198
rect 12077 8172 12086 8192
rect 12106 8172 12121 8192
rect 12077 8156 12121 8172
rect 12171 8188 12220 8198
rect 12171 8168 12189 8188
rect 12209 8168 12220 8188
rect 12171 8156 12220 8168
rect 13852 8159 13901 8171
rect 13852 8139 13863 8159
rect 13883 8139 13901 8159
rect 13852 8129 13901 8139
rect 13951 8155 13995 8171
rect 13951 8135 13966 8155
rect 13986 8135 13995 8155
rect 13951 8129 13995 8135
rect 14065 8155 14109 8171
rect 14065 8135 14074 8155
rect 14094 8135 14109 8155
rect 14065 8129 14109 8135
rect 14159 8159 14208 8171
rect 14159 8139 14177 8159
rect 14197 8139 14208 8159
rect 14159 8129 14208 8139
rect 14273 8155 14317 8171
rect 14273 8135 14282 8155
rect 14302 8135 14317 8155
rect 14273 8129 14317 8135
rect 14367 8159 14416 8171
rect 14367 8139 14385 8159
rect 14405 8139 14416 8159
rect 14367 8129 14416 8139
rect 14486 8155 14530 8171
rect 14486 8135 14495 8155
rect 14515 8135 14530 8155
rect 14486 8129 14530 8135
rect 14580 8159 14629 8171
rect 16499 8229 16548 8239
rect 16499 8209 16510 8229
rect 16530 8209 16548 8229
rect 16499 8197 16548 8209
rect 16598 8233 16642 8239
rect 16598 8213 16613 8233
rect 16633 8213 16642 8233
rect 16598 8197 16642 8213
rect 16712 8229 16761 8239
rect 16712 8209 16723 8229
rect 16743 8209 16761 8229
rect 16712 8197 16761 8209
rect 16811 8233 16855 8239
rect 16811 8213 16826 8233
rect 16846 8213 16855 8233
rect 16811 8197 16855 8213
rect 16920 8229 16969 8239
rect 16920 8209 16931 8229
rect 16951 8209 16969 8229
rect 16920 8197 16969 8209
rect 17019 8233 17063 8239
rect 17019 8213 17034 8233
rect 17054 8213 17063 8233
rect 17019 8197 17063 8213
rect 17133 8233 17177 8239
rect 17133 8213 17142 8233
rect 17162 8213 17177 8233
rect 17133 8197 17177 8213
rect 17227 8229 17276 8239
rect 17227 8209 17245 8229
rect 17265 8209 17276 8229
rect 17227 8197 17276 8209
rect 18908 8200 18957 8212
rect 18908 8180 18919 8200
rect 18939 8180 18957 8200
rect 18908 8170 18957 8180
rect 19007 8196 19051 8212
rect 19007 8176 19022 8196
rect 19042 8176 19051 8196
rect 19007 8170 19051 8176
rect 19121 8196 19165 8212
rect 19121 8176 19130 8196
rect 19150 8176 19165 8196
rect 19121 8170 19165 8176
rect 19215 8200 19264 8212
rect 19215 8180 19233 8200
rect 19253 8180 19264 8200
rect 19215 8170 19264 8180
rect 19329 8196 19373 8212
rect 19329 8176 19338 8196
rect 19358 8176 19373 8196
rect 19329 8170 19373 8176
rect 19423 8200 19472 8212
rect 19423 8180 19441 8200
rect 19461 8180 19472 8200
rect 19423 8170 19472 8180
rect 19542 8196 19586 8212
rect 19542 8176 19551 8196
rect 19571 8176 19586 8196
rect 19542 8170 19586 8176
rect 19636 8200 19685 8212
rect 19636 8180 19654 8200
rect 19674 8180 19685 8200
rect 19636 8170 19685 8180
rect 14580 8139 14598 8159
rect 14618 8139 14629 8159
rect 14580 8129 14629 8139
rect 5390 7957 5439 7967
rect 5390 7937 5401 7957
rect 5421 7937 5439 7957
rect 5390 7925 5439 7937
rect 5489 7961 5533 7967
rect 5489 7941 5504 7961
rect 5524 7941 5533 7961
rect 5489 7925 5533 7941
rect 5603 7957 5652 7967
rect 5603 7937 5614 7957
rect 5634 7937 5652 7957
rect 5603 7925 5652 7937
rect 5702 7961 5746 7967
rect 5702 7941 5717 7961
rect 5737 7941 5746 7961
rect 5702 7925 5746 7941
rect 5811 7957 5860 7967
rect 5811 7937 5822 7957
rect 5842 7937 5860 7957
rect 5811 7925 5860 7937
rect 5910 7961 5954 7967
rect 5910 7941 5925 7961
rect 5945 7941 5954 7961
rect 5910 7925 5954 7941
rect 6024 7961 6068 7967
rect 6024 7941 6033 7961
rect 6053 7941 6068 7961
rect 6024 7925 6068 7941
rect 6118 7957 6167 7967
rect 6118 7937 6136 7957
rect 6156 7937 6167 7957
rect 6118 7925 6167 7937
rect 2882 7844 2931 7856
rect 2882 7824 2893 7844
rect 2913 7824 2931 7844
rect 2882 7814 2931 7824
rect 2981 7840 3025 7856
rect 2981 7820 2996 7840
rect 3016 7820 3025 7840
rect 2981 7814 3025 7820
rect 3095 7840 3139 7856
rect 3095 7820 3104 7840
rect 3124 7820 3139 7840
rect 3095 7814 3139 7820
rect 3189 7844 3238 7856
rect 3189 7824 3207 7844
rect 3227 7824 3238 7844
rect 3189 7814 3238 7824
rect 3303 7840 3347 7856
rect 3303 7820 3312 7840
rect 3332 7820 3347 7840
rect 3303 7814 3347 7820
rect 3397 7844 3446 7856
rect 3397 7824 3415 7844
rect 3435 7824 3446 7844
rect 3397 7814 3446 7824
rect 3516 7840 3560 7856
rect 3516 7820 3525 7840
rect 3545 7820 3560 7840
rect 3516 7814 3560 7820
rect 3610 7844 3659 7856
rect 3610 7824 3628 7844
rect 3648 7824 3659 7844
rect 3610 7814 3659 7824
rect 1272 7672 1321 7682
rect 1272 7652 1283 7672
rect 1303 7652 1321 7672
rect 1272 7640 1321 7652
rect 1371 7676 1415 7682
rect 1371 7656 1386 7676
rect 1406 7656 1415 7676
rect 1371 7640 1415 7656
rect 1485 7672 1534 7682
rect 1485 7652 1496 7672
rect 1516 7652 1534 7672
rect 1485 7640 1534 7652
rect 1584 7676 1628 7682
rect 1584 7656 1599 7676
rect 1619 7656 1628 7676
rect 1584 7640 1628 7656
rect 1693 7672 1742 7682
rect 1693 7652 1704 7672
rect 1724 7652 1742 7672
rect 1693 7640 1742 7652
rect 1792 7676 1836 7682
rect 1792 7656 1807 7676
rect 1827 7656 1836 7676
rect 1792 7640 1836 7656
rect 1906 7676 1950 7682
rect 1906 7656 1915 7676
rect 1935 7656 1950 7676
rect 1906 7640 1950 7656
rect 2000 7672 2049 7682
rect 2000 7652 2018 7672
rect 2038 7652 2049 7672
rect 2000 7640 2049 7652
rect 7938 7885 7987 7897
rect 7938 7865 7949 7885
rect 7969 7865 7987 7885
rect 7938 7855 7987 7865
rect 8037 7881 8081 7897
rect 8037 7861 8052 7881
rect 8072 7861 8081 7881
rect 8037 7855 8081 7861
rect 8151 7881 8195 7897
rect 8151 7861 8160 7881
rect 8180 7861 8195 7881
rect 8151 7855 8195 7861
rect 8245 7885 8294 7897
rect 8245 7865 8263 7885
rect 8283 7865 8294 7885
rect 8245 7855 8294 7865
rect 8359 7881 8403 7897
rect 8359 7861 8368 7881
rect 8388 7861 8403 7881
rect 8359 7855 8403 7861
rect 8453 7885 8502 7897
rect 8453 7865 8471 7885
rect 8491 7865 8502 7885
rect 8453 7855 8502 7865
rect 8572 7881 8616 7897
rect 8572 7861 8581 7881
rect 8601 7861 8616 7881
rect 8572 7855 8616 7861
rect 8666 7885 8715 7897
rect 8666 7865 8684 7885
rect 8704 7865 8715 7885
rect 8666 7855 8715 7865
rect 10365 7921 10414 7931
rect 10365 7901 10376 7921
rect 10396 7901 10414 7921
rect 10365 7889 10414 7901
rect 10464 7925 10508 7931
rect 10464 7905 10479 7925
rect 10499 7905 10508 7925
rect 10464 7889 10508 7905
rect 10578 7921 10627 7931
rect 10578 7901 10589 7921
rect 10609 7901 10627 7921
rect 10578 7889 10627 7901
rect 10677 7925 10721 7931
rect 10677 7905 10692 7925
rect 10712 7905 10721 7925
rect 10677 7889 10721 7905
rect 10786 7921 10835 7931
rect 10786 7901 10797 7921
rect 10817 7901 10835 7921
rect 10786 7889 10835 7901
rect 10885 7925 10929 7931
rect 10885 7905 10900 7925
rect 10920 7905 10929 7925
rect 10885 7889 10929 7905
rect 10999 7925 11043 7931
rect 10999 7905 11008 7925
rect 11028 7905 11043 7925
rect 10999 7889 11043 7905
rect 11093 7921 11142 7931
rect 11093 7901 11111 7921
rect 11131 7901 11142 7921
rect 11093 7889 11142 7901
rect 15421 7962 15470 7972
rect 15421 7942 15432 7962
rect 15452 7942 15470 7962
rect 15421 7930 15470 7942
rect 15520 7966 15564 7972
rect 15520 7946 15535 7966
rect 15555 7946 15564 7966
rect 15520 7930 15564 7946
rect 15634 7962 15683 7972
rect 15634 7942 15645 7962
rect 15665 7942 15683 7962
rect 15634 7930 15683 7942
rect 15733 7966 15777 7972
rect 15733 7946 15748 7966
rect 15768 7946 15777 7966
rect 15733 7930 15777 7946
rect 15842 7962 15891 7972
rect 15842 7942 15853 7962
rect 15873 7942 15891 7962
rect 15842 7930 15891 7942
rect 15941 7966 15985 7972
rect 15941 7946 15956 7966
rect 15976 7946 15985 7966
rect 15941 7930 15985 7946
rect 16055 7966 16099 7972
rect 16055 7946 16064 7966
rect 16084 7946 16099 7966
rect 16055 7930 16099 7946
rect 16149 7962 16198 7972
rect 16149 7942 16167 7962
rect 16187 7942 16198 7962
rect 16149 7930 16198 7942
rect 6328 7713 6377 7723
rect 6328 7693 6339 7713
rect 6359 7693 6377 7713
rect 6328 7681 6377 7693
rect 6427 7717 6471 7723
rect 6427 7697 6442 7717
rect 6462 7697 6471 7717
rect 6427 7681 6471 7697
rect 6541 7713 6590 7723
rect 6541 7693 6552 7713
rect 6572 7693 6590 7713
rect 6541 7681 6590 7693
rect 6640 7717 6684 7723
rect 6640 7697 6655 7717
rect 6675 7697 6684 7717
rect 6640 7681 6684 7697
rect 6749 7713 6798 7723
rect 6749 7693 6760 7713
rect 6780 7693 6798 7713
rect 6749 7681 6798 7693
rect 6848 7717 6892 7723
rect 6848 7697 6863 7717
rect 6883 7697 6892 7717
rect 6848 7681 6892 7697
rect 6962 7717 7006 7723
rect 6962 7697 6971 7717
rect 6991 7697 7006 7717
rect 6962 7681 7006 7697
rect 7056 7713 7105 7723
rect 7056 7693 7074 7713
rect 7094 7693 7105 7713
rect 7056 7681 7105 7693
rect 12913 7849 12962 7861
rect 12913 7829 12924 7849
rect 12944 7829 12962 7849
rect 12913 7819 12962 7829
rect 13012 7845 13056 7861
rect 13012 7825 13027 7845
rect 13047 7825 13056 7845
rect 13012 7819 13056 7825
rect 13126 7845 13170 7861
rect 13126 7825 13135 7845
rect 13155 7825 13170 7845
rect 13126 7819 13170 7825
rect 13220 7849 13269 7861
rect 13220 7829 13238 7849
rect 13258 7829 13269 7849
rect 13220 7819 13269 7829
rect 13334 7845 13378 7861
rect 13334 7825 13343 7845
rect 13363 7825 13378 7845
rect 13334 7819 13378 7825
rect 13428 7849 13477 7861
rect 13428 7829 13446 7849
rect 13466 7829 13477 7849
rect 13428 7819 13477 7829
rect 13547 7845 13591 7861
rect 13547 7825 13556 7845
rect 13576 7825 13591 7845
rect 13547 7819 13591 7825
rect 13641 7849 13690 7861
rect 13641 7829 13659 7849
rect 13679 7829 13690 7849
rect 13641 7819 13690 7829
rect 3820 7600 3869 7612
rect 3820 7580 3831 7600
rect 3851 7580 3869 7600
rect 3820 7570 3869 7580
rect 3919 7596 3963 7612
rect 3919 7576 3934 7596
rect 3954 7576 3963 7596
rect 3919 7570 3963 7576
rect 4033 7596 4077 7612
rect 4033 7576 4042 7596
rect 4062 7576 4077 7596
rect 4033 7570 4077 7576
rect 4127 7600 4176 7612
rect 4127 7580 4145 7600
rect 4165 7580 4176 7600
rect 4127 7570 4176 7580
rect 4241 7596 4285 7612
rect 4241 7576 4250 7596
rect 4270 7576 4285 7596
rect 4241 7570 4285 7576
rect 4335 7600 4384 7612
rect 4335 7580 4353 7600
rect 4373 7580 4384 7600
rect 4335 7570 4384 7580
rect 4454 7596 4498 7612
rect 4454 7576 4463 7596
rect 4483 7576 4498 7596
rect 4454 7570 4498 7576
rect 4548 7600 4597 7612
rect 4548 7580 4566 7600
rect 4586 7580 4597 7600
rect 4548 7570 4597 7580
rect 8876 7641 8925 7653
rect 8876 7621 8887 7641
rect 8907 7621 8925 7641
rect 8876 7611 8925 7621
rect 8975 7637 9019 7653
rect 8975 7617 8990 7637
rect 9010 7617 9019 7637
rect 8975 7611 9019 7617
rect 9089 7637 9133 7653
rect 9089 7617 9098 7637
rect 9118 7617 9133 7637
rect 9089 7611 9133 7617
rect 9183 7641 9232 7653
rect 9183 7621 9201 7641
rect 9221 7621 9232 7641
rect 9183 7611 9232 7621
rect 9297 7637 9341 7653
rect 9297 7617 9306 7637
rect 9326 7617 9341 7637
rect 9297 7611 9341 7617
rect 9391 7641 9440 7653
rect 9391 7621 9409 7641
rect 9429 7621 9440 7641
rect 9391 7611 9440 7621
rect 9510 7637 9554 7653
rect 9510 7617 9519 7637
rect 9539 7617 9554 7637
rect 9510 7611 9554 7617
rect 9604 7641 9653 7653
rect 9604 7621 9622 7641
rect 9642 7621 9653 7641
rect 9604 7611 9653 7621
rect 11303 7677 11352 7687
rect 11303 7657 11314 7677
rect 11334 7657 11352 7677
rect 11303 7645 11352 7657
rect 11402 7681 11446 7687
rect 11402 7661 11417 7681
rect 11437 7661 11446 7681
rect 11402 7645 11446 7661
rect 11516 7677 11565 7687
rect 11516 7657 11527 7677
rect 11547 7657 11565 7677
rect 11516 7645 11565 7657
rect 11615 7681 11659 7687
rect 11615 7661 11630 7681
rect 11650 7661 11659 7681
rect 11615 7645 11659 7661
rect 11724 7677 11773 7687
rect 11724 7657 11735 7677
rect 11755 7657 11773 7677
rect 11724 7645 11773 7657
rect 11823 7681 11867 7687
rect 11823 7661 11838 7681
rect 11858 7661 11867 7681
rect 11823 7645 11867 7661
rect 11937 7681 11981 7687
rect 11937 7661 11946 7681
rect 11966 7661 11981 7681
rect 11937 7645 11981 7661
rect 12031 7677 12080 7687
rect 12031 7657 12049 7677
rect 12069 7657 12080 7677
rect 12031 7645 12080 7657
rect 17969 7890 18018 7902
rect 17969 7870 17980 7890
rect 18000 7870 18018 7890
rect 17969 7860 18018 7870
rect 18068 7886 18112 7902
rect 18068 7866 18083 7886
rect 18103 7866 18112 7886
rect 18068 7860 18112 7866
rect 18182 7886 18226 7902
rect 18182 7866 18191 7886
rect 18211 7866 18226 7886
rect 18182 7860 18226 7866
rect 18276 7890 18325 7902
rect 18276 7870 18294 7890
rect 18314 7870 18325 7890
rect 18276 7860 18325 7870
rect 18390 7886 18434 7902
rect 18390 7866 18399 7886
rect 18419 7866 18434 7886
rect 18390 7860 18434 7866
rect 18484 7890 18533 7902
rect 18484 7870 18502 7890
rect 18522 7870 18533 7890
rect 18484 7860 18533 7870
rect 18603 7886 18647 7902
rect 18603 7866 18612 7886
rect 18632 7866 18647 7886
rect 18603 7860 18647 7866
rect 18697 7890 18746 7902
rect 18697 7870 18715 7890
rect 18735 7870 18746 7890
rect 18697 7860 18746 7870
rect 16359 7718 16408 7728
rect 16359 7698 16370 7718
rect 16390 7698 16408 7718
rect 16359 7686 16408 7698
rect 16458 7722 16502 7728
rect 16458 7702 16473 7722
rect 16493 7702 16502 7722
rect 16458 7686 16502 7702
rect 16572 7718 16621 7728
rect 16572 7698 16583 7718
rect 16603 7698 16621 7718
rect 16572 7686 16621 7698
rect 16671 7722 16715 7728
rect 16671 7702 16686 7722
rect 16706 7702 16715 7722
rect 16671 7686 16715 7702
rect 16780 7718 16829 7728
rect 16780 7698 16791 7718
rect 16811 7698 16829 7718
rect 16780 7686 16829 7698
rect 16879 7722 16923 7728
rect 16879 7702 16894 7722
rect 16914 7702 16923 7722
rect 16879 7686 16923 7702
rect 16993 7722 17037 7728
rect 16993 7702 17002 7722
rect 17022 7702 17037 7722
rect 16993 7686 17037 7702
rect 17087 7718 17136 7728
rect 17087 7698 17105 7718
rect 17125 7698 17136 7718
rect 17087 7686 17136 7698
rect 13851 7605 13900 7617
rect 13851 7585 13862 7605
rect 13882 7585 13900 7605
rect 13851 7575 13900 7585
rect 13950 7601 13994 7617
rect 13950 7581 13965 7601
rect 13985 7581 13994 7601
rect 13950 7575 13994 7581
rect 14064 7601 14108 7617
rect 14064 7581 14073 7601
rect 14093 7581 14108 7601
rect 14064 7575 14108 7581
rect 14158 7605 14207 7617
rect 14158 7585 14176 7605
rect 14196 7585 14207 7605
rect 14158 7575 14207 7585
rect 14272 7601 14316 7617
rect 14272 7581 14281 7601
rect 14301 7581 14316 7601
rect 14272 7575 14316 7581
rect 14366 7605 14415 7617
rect 14366 7585 14384 7605
rect 14404 7585 14415 7605
rect 14366 7575 14415 7585
rect 14485 7601 14529 7617
rect 14485 7581 14494 7601
rect 14514 7581 14529 7601
rect 14485 7575 14529 7581
rect 14579 7605 14628 7617
rect 14579 7585 14597 7605
rect 14617 7585 14628 7605
rect 14579 7575 14628 7585
rect 5389 7403 5438 7413
rect 5389 7383 5400 7403
rect 5420 7383 5438 7403
rect 333 7362 382 7372
rect 333 7342 344 7362
rect 364 7342 382 7362
rect 333 7330 382 7342
rect 432 7366 476 7372
rect 432 7346 447 7366
rect 467 7346 476 7366
rect 432 7330 476 7346
rect 546 7362 595 7372
rect 546 7342 557 7362
rect 577 7342 595 7362
rect 546 7330 595 7342
rect 645 7366 689 7372
rect 645 7346 660 7366
rect 680 7346 689 7366
rect 645 7330 689 7346
rect 754 7362 803 7372
rect 754 7342 765 7362
rect 785 7342 803 7362
rect 754 7330 803 7342
rect 853 7366 897 7372
rect 853 7346 868 7366
rect 888 7346 897 7366
rect 853 7330 897 7346
rect 967 7366 1011 7372
rect 967 7346 976 7366
rect 996 7346 1011 7366
rect 967 7330 1011 7346
rect 1061 7362 1110 7372
rect 1061 7342 1079 7362
rect 1099 7342 1110 7362
rect 1061 7330 1110 7342
rect 2772 7320 2821 7332
rect 2772 7300 2783 7320
rect 2803 7300 2821 7320
rect 2772 7290 2821 7300
rect 2871 7316 2915 7332
rect 2871 7296 2886 7316
rect 2906 7296 2915 7316
rect 2871 7290 2915 7296
rect 2985 7316 3029 7332
rect 2985 7296 2994 7316
rect 3014 7296 3029 7316
rect 2985 7290 3029 7296
rect 3079 7320 3128 7332
rect 3079 7300 3097 7320
rect 3117 7300 3128 7320
rect 3079 7290 3128 7300
rect 3193 7316 3237 7332
rect 3193 7296 3202 7316
rect 3222 7296 3237 7316
rect 3193 7290 3237 7296
rect 3287 7320 3336 7332
rect 3287 7300 3305 7320
rect 3325 7300 3336 7320
rect 3287 7290 3336 7300
rect 3406 7316 3450 7332
rect 3406 7296 3415 7316
rect 3435 7296 3450 7316
rect 3406 7290 3450 7296
rect 3500 7320 3549 7332
rect 3500 7300 3518 7320
rect 3538 7300 3549 7320
rect 5389 7371 5438 7383
rect 5488 7407 5532 7413
rect 5488 7387 5503 7407
rect 5523 7387 5532 7407
rect 5488 7371 5532 7387
rect 5602 7403 5651 7413
rect 5602 7383 5613 7403
rect 5633 7383 5651 7403
rect 5602 7371 5651 7383
rect 5701 7407 5745 7413
rect 5701 7387 5716 7407
rect 5736 7387 5745 7407
rect 5701 7371 5745 7387
rect 5810 7403 5859 7413
rect 5810 7383 5821 7403
rect 5841 7383 5859 7403
rect 5810 7371 5859 7383
rect 5909 7407 5953 7413
rect 5909 7387 5924 7407
rect 5944 7387 5953 7407
rect 5909 7371 5953 7387
rect 6023 7407 6067 7413
rect 6023 7387 6032 7407
rect 6052 7387 6067 7407
rect 6023 7371 6067 7387
rect 6117 7403 6166 7413
rect 6117 7383 6135 7403
rect 6155 7383 6166 7403
rect 6117 7371 6166 7383
rect 7828 7361 7877 7373
rect 7828 7341 7839 7361
rect 7859 7341 7877 7361
rect 3500 7290 3549 7300
rect 7828 7331 7877 7341
rect 7927 7357 7971 7373
rect 7927 7337 7942 7357
rect 7962 7337 7971 7357
rect 7927 7331 7971 7337
rect 8041 7357 8085 7373
rect 8041 7337 8050 7357
rect 8070 7337 8085 7357
rect 8041 7331 8085 7337
rect 8135 7361 8184 7373
rect 8135 7341 8153 7361
rect 8173 7341 8184 7361
rect 8135 7331 8184 7341
rect 8249 7357 8293 7373
rect 8249 7337 8258 7357
rect 8278 7337 8293 7357
rect 8249 7331 8293 7337
rect 8343 7361 8392 7373
rect 8343 7341 8361 7361
rect 8381 7341 8392 7361
rect 8343 7331 8392 7341
rect 8462 7357 8506 7373
rect 8462 7337 8471 7357
rect 8491 7337 8506 7357
rect 8462 7331 8506 7337
rect 8556 7361 8605 7373
rect 8556 7341 8574 7361
rect 8594 7341 8605 7361
rect 18907 7646 18956 7658
rect 18907 7626 18918 7646
rect 18938 7626 18956 7646
rect 18907 7616 18956 7626
rect 19006 7642 19050 7658
rect 19006 7622 19021 7642
rect 19041 7622 19050 7642
rect 19006 7616 19050 7622
rect 19120 7642 19164 7658
rect 19120 7622 19129 7642
rect 19149 7622 19164 7642
rect 19120 7616 19164 7622
rect 19214 7646 19263 7658
rect 19214 7626 19232 7646
rect 19252 7626 19263 7646
rect 19214 7616 19263 7626
rect 19328 7642 19372 7658
rect 19328 7622 19337 7642
rect 19357 7622 19372 7642
rect 19328 7616 19372 7622
rect 19422 7646 19471 7658
rect 19422 7626 19440 7646
rect 19460 7626 19471 7646
rect 19422 7616 19471 7626
rect 19541 7642 19585 7658
rect 19541 7622 19550 7642
rect 19570 7622 19585 7642
rect 19541 7616 19585 7622
rect 19635 7646 19684 7658
rect 19635 7626 19653 7646
rect 19673 7626 19684 7646
rect 19635 7616 19684 7626
rect 15420 7408 15469 7418
rect 15420 7388 15431 7408
rect 15451 7388 15469 7408
rect 8556 7331 8605 7341
rect 10364 7367 10413 7377
rect 10364 7347 10375 7367
rect 10395 7347 10413 7367
rect 10364 7335 10413 7347
rect 10463 7371 10507 7377
rect 10463 7351 10478 7371
rect 10498 7351 10507 7371
rect 10463 7335 10507 7351
rect 10577 7367 10626 7377
rect 10577 7347 10588 7367
rect 10608 7347 10626 7367
rect 10577 7335 10626 7347
rect 10676 7371 10720 7377
rect 10676 7351 10691 7371
rect 10711 7351 10720 7371
rect 10676 7335 10720 7351
rect 10785 7367 10834 7377
rect 10785 7347 10796 7367
rect 10816 7347 10834 7367
rect 10785 7335 10834 7347
rect 10884 7371 10928 7377
rect 10884 7351 10899 7371
rect 10919 7351 10928 7371
rect 10884 7335 10928 7351
rect 10998 7371 11042 7377
rect 10998 7351 11007 7371
rect 11027 7351 11042 7371
rect 10998 7335 11042 7351
rect 11092 7367 11141 7377
rect 11092 7347 11110 7367
rect 11130 7347 11141 7367
rect 11092 7335 11141 7347
rect 12803 7325 12852 7337
rect 12803 7305 12814 7325
rect 12834 7305 12852 7325
rect 12803 7295 12852 7305
rect 12902 7321 12946 7337
rect 12902 7301 12917 7321
rect 12937 7301 12946 7321
rect 12902 7295 12946 7301
rect 13016 7321 13060 7337
rect 13016 7301 13025 7321
rect 13045 7301 13060 7321
rect 13016 7295 13060 7301
rect 13110 7325 13159 7337
rect 13110 7305 13128 7325
rect 13148 7305 13159 7325
rect 13110 7295 13159 7305
rect 13224 7321 13268 7337
rect 13224 7301 13233 7321
rect 13253 7301 13268 7321
rect 13224 7295 13268 7301
rect 13318 7325 13367 7337
rect 13318 7305 13336 7325
rect 13356 7305 13367 7325
rect 13318 7295 13367 7305
rect 13437 7321 13481 7337
rect 13437 7301 13446 7321
rect 13466 7301 13481 7321
rect 13437 7295 13481 7301
rect 13531 7325 13580 7337
rect 13531 7305 13549 7325
rect 13569 7305 13580 7325
rect 15420 7376 15469 7388
rect 15519 7412 15563 7418
rect 15519 7392 15534 7412
rect 15554 7392 15563 7412
rect 15519 7376 15563 7392
rect 15633 7408 15682 7418
rect 15633 7388 15644 7408
rect 15664 7388 15682 7408
rect 15633 7376 15682 7388
rect 15732 7412 15776 7418
rect 15732 7392 15747 7412
rect 15767 7392 15776 7412
rect 15732 7376 15776 7392
rect 15841 7408 15890 7418
rect 15841 7388 15852 7408
rect 15872 7388 15890 7408
rect 15841 7376 15890 7388
rect 15940 7412 15984 7418
rect 15940 7392 15955 7412
rect 15975 7392 15984 7412
rect 15940 7376 15984 7392
rect 16054 7412 16098 7418
rect 16054 7392 16063 7412
rect 16083 7392 16098 7412
rect 16054 7376 16098 7392
rect 16148 7408 16197 7418
rect 16148 7388 16166 7408
rect 16186 7388 16197 7408
rect 16148 7376 16197 7388
rect 17859 7366 17908 7378
rect 17859 7346 17870 7366
rect 17890 7346 17908 7366
rect 13531 7295 13580 7305
rect 17859 7336 17908 7346
rect 17958 7362 18002 7378
rect 17958 7342 17973 7362
rect 17993 7342 18002 7362
rect 17958 7336 18002 7342
rect 18072 7362 18116 7378
rect 18072 7342 18081 7362
rect 18101 7342 18116 7362
rect 18072 7336 18116 7342
rect 18166 7366 18215 7378
rect 18166 7346 18184 7366
rect 18204 7346 18215 7366
rect 18166 7336 18215 7346
rect 18280 7362 18324 7378
rect 18280 7342 18289 7362
rect 18309 7342 18324 7362
rect 18280 7336 18324 7342
rect 18374 7366 18423 7378
rect 18374 7346 18392 7366
rect 18412 7346 18423 7366
rect 18374 7336 18423 7346
rect 18493 7362 18537 7378
rect 18493 7342 18502 7362
rect 18522 7342 18537 7362
rect 18493 7336 18537 7342
rect 18587 7366 18636 7378
rect 18587 7346 18605 7366
rect 18625 7346 18636 7366
rect 18587 7336 18636 7346
rect 1382 7093 1431 7103
rect 1382 7073 1393 7093
rect 1413 7073 1431 7093
rect 1382 7061 1431 7073
rect 1481 7097 1525 7103
rect 1481 7077 1496 7097
rect 1516 7077 1525 7097
rect 1481 7061 1525 7077
rect 1595 7093 1644 7103
rect 1595 7073 1606 7093
rect 1626 7073 1644 7093
rect 1595 7061 1644 7073
rect 1694 7097 1738 7103
rect 1694 7077 1709 7097
rect 1729 7077 1738 7097
rect 1694 7061 1738 7077
rect 1803 7093 1852 7103
rect 1803 7073 1814 7093
rect 1834 7073 1852 7093
rect 1803 7061 1852 7073
rect 1902 7097 1946 7103
rect 1902 7077 1917 7097
rect 1937 7077 1946 7097
rect 1902 7061 1946 7077
rect 2016 7097 2060 7103
rect 2016 7077 2025 7097
rect 2045 7077 2060 7097
rect 2016 7061 2060 7077
rect 2110 7093 2159 7103
rect 6438 7134 6487 7144
rect 2110 7073 2128 7093
rect 2148 7073 2159 7093
rect 2110 7061 2159 7073
rect 3821 7051 3870 7063
rect 3821 7031 3832 7051
rect 3852 7031 3870 7051
rect 3821 7021 3870 7031
rect 3920 7047 3964 7063
rect 3920 7027 3935 7047
rect 3955 7027 3964 7047
rect 3920 7021 3964 7027
rect 4034 7047 4078 7063
rect 4034 7027 4043 7047
rect 4063 7027 4078 7047
rect 4034 7021 4078 7027
rect 4128 7051 4177 7063
rect 4128 7031 4146 7051
rect 4166 7031 4177 7051
rect 4128 7021 4177 7031
rect 4242 7047 4286 7063
rect 4242 7027 4251 7047
rect 4271 7027 4286 7047
rect 4242 7021 4286 7027
rect 4336 7051 4385 7063
rect 4336 7031 4354 7051
rect 4374 7031 4385 7051
rect 4336 7021 4385 7031
rect 4455 7047 4499 7063
rect 4455 7027 4464 7047
rect 4484 7027 4499 7047
rect 4455 7021 4499 7027
rect 4549 7051 4598 7063
rect 6438 7114 6449 7134
rect 6469 7114 6487 7134
rect 6438 7102 6487 7114
rect 6537 7138 6581 7144
rect 6537 7118 6552 7138
rect 6572 7118 6581 7138
rect 6537 7102 6581 7118
rect 6651 7134 6700 7144
rect 6651 7114 6662 7134
rect 6682 7114 6700 7134
rect 6651 7102 6700 7114
rect 6750 7138 6794 7144
rect 6750 7118 6765 7138
rect 6785 7118 6794 7138
rect 6750 7102 6794 7118
rect 6859 7134 6908 7144
rect 6859 7114 6870 7134
rect 6890 7114 6908 7134
rect 6859 7102 6908 7114
rect 6958 7138 7002 7144
rect 6958 7118 6973 7138
rect 6993 7118 7002 7138
rect 6958 7102 7002 7118
rect 7072 7138 7116 7144
rect 7072 7118 7081 7138
rect 7101 7118 7116 7138
rect 7072 7102 7116 7118
rect 7166 7134 7215 7144
rect 7166 7114 7184 7134
rect 7204 7114 7215 7134
rect 7166 7102 7215 7114
rect 8877 7092 8926 7104
rect 8877 7072 8888 7092
rect 8908 7072 8926 7092
rect 8877 7062 8926 7072
rect 8976 7088 9020 7104
rect 8976 7068 8991 7088
rect 9011 7068 9020 7088
rect 8976 7062 9020 7068
rect 9090 7088 9134 7104
rect 9090 7068 9099 7088
rect 9119 7068 9134 7088
rect 9090 7062 9134 7068
rect 9184 7092 9233 7104
rect 9184 7072 9202 7092
rect 9222 7072 9233 7092
rect 9184 7062 9233 7072
rect 9298 7088 9342 7104
rect 9298 7068 9307 7088
rect 9327 7068 9342 7088
rect 9298 7062 9342 7068
rect 9392 7092 9441 7104
rect 9392 7072 9410 7092
rect 9430 7072 9441 7092
rect 9392 7062 9441 7072
rect 9511 7088 9555 7104
rect 9511 7068 9520 7088
rect 9540 7068 9555 7088
rect 9511 7062 9555 7068
rect 9605 7092 9654 7104
rect 9605 7072 9623 7092
rect 9643 7072 9654 7092
rect 9605 7062 9654 7072
rect 11413 7098 11462 7108
rect 4549 7031 4567 7051
rect 4587 7031 4598 7051
rect 4549 7021 4598 7031
rect 334 6813 383 6823
rect 334 6793 345 6813
rect 365 6793 383 6813
rect 334 6781 383 6793
rect 433 6817 477 6823
rect 433 6797 448 6817
rect 468 6797 477 6817
rect 433 6781 477 6797
rect 547 6813 596 6823
rect 547 6793 558 6813
rect 578 6793 596 6813
rect 547 6781 596 6793
rect 646 6817 690 6823
rect 646 6797 661 6817
rect 681 6797 690 6817
rect 646 6781 690 6797
rect 755 6813 804 6823
rect 755 6793 766 6813
rect 786 6793 804 6813
rect 755 6781 804 6793
rect 854 6817 898 6823
rect 854 6797 869 6817
rect 889 6797 898 6817
rect 854 6781 898 6797
rect 968 6817 1012 6823
rect 968 6797 977 6817
rect 997 6797 1012 6817
rect 968 6781 1012 6797
rect 1062 6813 1111 6823
rect 1062 6793 1080 6813
rect 1100 6793 1111 6813
rect 1062 6781 1111 6793
rect 11413 7078 11424 7098
rect 11444 7078 11462 7098
rect 11413 7066 11462 7078
rect 11512 7102 11556 7108
rect 11512 7082 11527 7102
rect 11547 7082 11556 7102
rect 11512 7066 11556 7082
rect 11626 7098 11675 7108
rect 11626 7078 11637 7098
rect 11657 7078 11675 7098
rect 11626 7066 11675 7078
rect 11725 7102 11769 7108
rect 11725 7082 11740 7102
rect 11760 7082 11769 7102
rect 11725 7066 11769 7082
rect 11834 7098 11883 7108
rect 11834 7078 11845 7098
rect 11865 7078 11883 7098
rect 11834 7066 11883 7078
rect 11933 7102 11977 7108
rect 11933 7082 11948 7102
rect 11968 7082 11977 7102
rect 11933 7066 11977 7082
rect 12047 7102 12091 7108
rect 12047 7082 12056 7102
rect 12076 7082 12091 7102
rect 12047 7066 12091 7082
rect 12141 7098 12190 7108
rect 16469 7139 16518 7149
rect 12141 7078 12159 7098
rect 12179 7078 12190 7098
rect 12141 7066 12190 7078
rect 13852 7056 13901 7068
rect 13852 7036 13863 7056
rect 13883 7036 13901 7056
rect 13852 7026 13901 7036
rect 13951 7052 13995 7068
rect 13951 7032 13966 7052
rect 13986 7032 13995 7052
rect 13951 7026 13995 7032
rect 14065 7052 14109 7068
rect 14065 7032 14074 7052
rect 14094 7032 14109 7052
rect 14065 7026 14109 7032
rect 14159 7056 14208 7068
rect 14159 7036 14177 7056
rect 14197 7036 14208 7056
rect 14159 7026 14208 7036
rect 14273 7052 14317 7068
rect 14273 7032 14282 7052
rect 14302 7032 14317 7052
rect 14273 7026 14317 7032
rect 14367 7056 14416 7068
rect 14367 7036 14385 7056
rect 14405 7036 14416 7056
rect 14367 7026 14416 7036
rect 14486 7052 14530 7068
rect 14486 7032 14495 7052
rect 14515 7032 14530 7052
rect 14486 7026 14530 7032
rect 14580 7056 14629 7068
rect 16469 7119 16480 7139
rect 16500 7119 16518 7139
rect 16469 7107 16518 7119
rect 16568 7143 16612 7149
rect 16568 7123 16583 7143
rect 16603 7123 16612 7143
rect 16568 7107 16612 7123
rect 16682 7139 16731 7149
rect 16682 7119 16693 7139
rect 16713 7119 16731 7139
rect 16682 7107 16731 7119
rect 16781 7143 16825 7149
rect 16781 7123 16796 7143
rect 16816 7123 16825 7143
rect 16781 7107 16825 7123
rect 16890 7139 16939 7149
rect 16890 7119 16901 7139
rect 16921 7119 16939 7139
rect 16890 7107 16939 7119
rect 16989 7143 17033 7149
rect 16989 7123 17004 7143
rect 17024 7123 17033 7143
rect 16989 7107 17033 7123
rect 17103 7143 17147 7149
rect 17103 7123 17112 7143
rect 17132 7123 17147 7143
rect 17103 7107 17147 7123
rect 17197 7139 17246 7149
rect 17197 7119 17215 7139
rect 17235 7119 17246 7139
rect 17197 7107 17246 7119
rect 18908 7097 18957 7109
rect 18908 7077 18919 7097
rect 18939 7077 18957 7097
rect 18908 7067 18957 7077
rect 19007 7093 19051 7109
rect 19007 7073 19022 7093
rect 19042 7073 19051 7093
rect 19007 7067 19051 7073
rect 19121 7093 19165 7109
rect 19121 7073 19130 7093
rect 19150 7073 19165 7093
rect 19121 7067 19165 7073
rect 19215 7097 19264 7109
rect 19215 7077 19233 7097
rect 19253 7077 19264 7097
rect 19215 7067 19264 7077
rect 19329 7093 19373 7109
rect 19329 7073 19338 7093
rect 19358 7073 19373 7093
rect 19329 7067 19373 7073
rect 19423 7097 19472 7109
rect 19423 7077 19441 7097
rect 19461 7077 19472 7097
rect 19423 7067 19472 7077
rect 19542 7093 19586 7109
rect 19542 7073 19551 7093
rect 19571 7073 19586 7093
rect 19542 7067 19586 7073
rect 19636 7097 19685 7109
rect 19636 7077 19654 7097
rect 19674 7077 19685 7097
rect 19636 7067 19685 7077
rect 14580 7036 14598 7056
rect 14618 7036 14629 7056
rect 14580 7026 14629 7036
rect 5390 6854 5439 6864
rect 5390 6834 5401 6854
rect 5421 6834 5439 6854
rect 5390 6822 5439 6834
rect 5489 6858 5533 6864
rect 5489 6838 5504 6858
rect 5524 6838 5533 6858
rect 5489 6822 5533 6838
rect 5603 6854 5652 6864
rect 5603 6834 5614 6854
rect 5634 6834 5652 6854
rect 5603 6822 5652 6834
rect 5702 6858 5746 6864
rect 5702 6838 5717 6858
rect 5737 6838 5746 6858
rect 5702 6822 5746 6838
rect 5811 6854 5860 6864
rect 5811 6834 5822 6854
rect 5842 6834 5860 6854
rect 5811 6822 5860 6834
rect 5910 6858 5954 6864
rect 5910 6838 5925 6858
rect 5945 6838 5954 6858
rect 5910 6822 5954 6838
rect 6024 6858 6068 6864
rect 6024 6838 6033 6858
rect 6053 6838 6068 6858
rect 6024 6822 6068 6838
rect 6118 6854 6167 6864
rect 6118 6834 6136 6854
rect 6156 6834 6167 6854
rect 6118 6822 6167 6834
rect 2882 6741 2931 6753
rect 2882 6721 2893 6741
rect 2913 6721 2931 6741
rect 2882 6711 2931 6721
rect 2981 6737 3025 6753
rect 2981 6717 2996 6737
rect 3016 6717 3025 6737
rect 2981 6711 3025 6717
rect 3095 6737 3139 6753
rect 3095 6717 3104 6737
rect 3124 6717 3139 6737
rect 3095 6711 3139 6717
rect 3189 6741 3238 6753
rect 3189 6721 3207 6741
rect 3227 6721 3238 6741
rect 3189 6711 3238 6721
rect 3303 6737 3347 6753
rect 3303 6717 3312 6737
rect 3332 6717 3347 6737
rect 3303 6711 3347 6717
rect 3397 6741 3446 6753
rect 3397 6721 3415 6741
rect 3435 6721 3446 6741
rect 3397 6711 3446 6721
rect 3516 6737 3560 6753
rect 3516 6717 3525 6737
rect 3545 6717 3560 6737
rect 3516 6711 3560 6717
rect 3610 6741 3659 6753
rect 3610 6721 3628 6741
rect 3648 6721 3659 6741
rect 3610 6711 3659 6721
rect 1272 6569 1321 6579
rect 1272 6549 1283 6569
rect 1303 6549 1321 6569
rect 1272 6537 1321 6549
rect 1371 6573 1415 6579
rect 1371 6553 1386 6573
rect 1406 6553 1415 6573
rect 1371 6537 1415 6553
rect 1485 6569 1534 6579
rect 1485 6549 1496 6569
rect 1516 6549 1534 6569
rect 1485 6537 1534 6549
rect 1584 6573 1628 6579
rect 1584 6553 1599 6573
rect 1619 6553 1628 6573
rect 1584 6537 1628 6553
rect 1693 6569 1742 6579
rect 1693 6549 1704 6569
rect 1724 6549 1742 6569
rect 1693 6537 1742 6549
rect 1792 6573 1836 6579
rect 1792 6553 1807 6573
rect 1827 6553 1836 6573
rect 1792 6537 1836 6553
rect 1906 6573 1950 6579
rect 1906 6553 1915 6573
rect 1935 6553 1950 6573
rect 1906 6537 1950 6553
rect 2000 6569 2049 6579
rect 2000 6549 2018 6569
rect 2038 6549 2049 6569
rect 2000 6537 2049 6549
rect 7938 6782 7987 6794
rect 7938 6762 7949 6782
rect 7969 6762 7987 6782
rect 7938 6752 7987 6762
rect 8037 6778 8081 6794
rect 8037 6758 8052 6778
rect 8072 6758 8081 6778
rect 8037 6752 8081 6758
rect 8151 6778 8195 6794
rect 8151 6758 8160 6778
rect 8180 6758 8195 6778
rect 8151 6752 8195 6758
rect 8245 6782 8294 6794
rect 8245 6762 8263 6782
rect 8283 6762 8294 6782
rect 8245 6752 8294 6762
rect 8359 6778 8403 6794
rect 8359 6758 8368 6778
rect 8388 6758 8403 6778
rect 8359 6752 8403 6758
rect 8453 6782 8502 6794
rect 8453 6762 8471 6782
rect 8491 6762 8502 6782
rect 8453 6752 8502 6762
rect 8572 6778 8616 6794
rect 8572 6758 8581 6778
rect 8601 6758 8616 6778
rect 8572 6752 8616 6758
rect 8666 6782 8715 6794
rect 8666 6762 8684 6782
rect 8704 6762 8715 6782
rect 8666 6752 8715 6762
rect 10365 6818 10414 6828
rect 10365 6798 10376 6818
rect 10396 6798 10414 6818
rect 10365 6786 10414 6798
rect 10464 6822 10508 6828
rect 10464 6802 10479 6822
rect 10499 6802 10508 6822
rect 10464 6786 10508 6802
rect 10578 6818 10627 6828
rect 10578 6798 10589 6818
rect 10609 6798 10627 6818
rect 10578 6786 10627 6798
rect 10677 6822 10721 6828
rect 10677 6802 10692 6822
rect 10712 6802 10721 6822
rect 10677 6786 10721 6802
rect 10786 6818 10835 6828
rect 10786 6798 10797 6818
rect 10817 6798 10835 6818
rect 10786 6786 10835 6798
rect 10885 6822 10929 6828
rect 10885 6802 10900 6822
rect 10920 6802 10929 6822
rect 10885 6786 10929 6802
rect 10999 6822 11043 6828
rect 10999 6802 11008 6822
rect 11028 6802 11043 6822
rect 10999 6786 11043 6802
rect 11093 6818 11142 6828
rect 11093 6798 11111 6818
rect 11131 6798 11142 6818
rect 11093 6786 11142 6798
rect 15421 6859 15470 6869
rect 15421 6839 15432 6859
rect 15452 6839 15470 6859
rect 15421 6827 15470 6839
rect 15520 6863 15564 6869
rect 15520 6843 15535 6863
rect 15555 6843 15564 6863
rect 15520 6827 15564 6843
rect 15634 6859 15683 6869
rect 15634 6839 15645 6859
rect 15665 6839 15683 6859
rect 15634 6827 15683 6839
rect 15733 6863 15777 6869
rect 15733 6843 15748 6863
rect 15768 6843 15777 6863
rect 15733 6827 15777 6843
rect 15842 6859 15891 6869
rect 15842 6839 15853 6859
rect 15873 6839 15891 6859
rect 15842 6827 15891 6839
rect 15941 6863 15985 6869
rect 15941 6843 15956 6863
rect 15976 6843 15985 6863
rect 15941 6827 15985 6843
rect 16055 6863 16099 6869
rect 16055 6843 16064 6863
rect 16084 6843 16099 6863
rect 16055 6827 16099 6843
rect 16149 6859 16198 6869
rect 16149 6839 16167 6859
rect 16187 6839 16198 6859
rect 16149 6827 16198 6839
rect 6328 6610 6377 6620
rect 6328 6590 6339 6610
rect 6359 6590 6377 6610
rect 6328 6578 6377 6590
rect 6427 6614 6471 6620
rect 6427 6594 6442 6614
rect 6462 6594 6471 6614
rect 6427 6578 6471 6594
rect 6541 6610 6590 6620
rect 6541 6590 6552 6610
rect 6572 6590 6590 6610
rect 6541 6578 6590 6590
rect 6640 6614 6684 6620
rect 6640 6594 6655 6614
rect 6675 6594 6684 6614
rect 6640 6578 6684 6594
rect 6749 6610 6798 6620
rect 6749 6590 6760 6610
rect 6780 6590 6798 6610
rect 6749 6578 6798 6590
rect 6848 6614 6892 6620
rect 6848 6594 6863 6614
rect 6883 6594 6892 6614
rect 6848 6578 6892 6594
rect 6962 6614 7006 6620
rect 6962 6594 6971 6614
rect 6991 6594 7006 6614
rect 6962 6578 7006 6594
rect 7056 6610 7105 6620
rect 7056 6590 7074 6610
rect 7094 6590 7105 6610
rect 7056 6578 7105 6590
rect 12913 6746 12962 6758
rect 12913 6726 12924 6746
rect 12944 6726 12962 6746
rect 12913 6716 12962 6726
rect 13012 6742 13056 6758
rect 13012 6722 13027 6742
rect 13047 6722 13056 6742
rect 13012 6716 13056 6722
rect 13126 6742 13170 6758
rect 13126 6722 13135 6742
rect 13155 6722 13170 6742
rect 13126 6716 13170 6722
rect 13220 6746 13269 6758
rect 13220 6726 13238 6746
rect 13258 6726 13269 6746
rect 13220 6716 13269 6726
rect 13334 6742 13378 6758
rect 13334 6722 13343 6742
rect 13363 6722 13378 6742
rect 13334 6716 13378 6722
rect 13428 6746 13477 6758
rect 13428 6726 13446 6746
rect 13466 6726 13477 6746
rect 13428 6716 13477 6726
rect 13547 6742 13591 6758
rect 13547 6722 13556 6742
rect 13576 6722 13591 6742
rect 13547 6716 13591 6722
rect 13641 6746 13690 6758
rect 13641 6726 13659 6746
rect 13679 6726 13690 6746
rect 13641 6716 13690 6726
rect 3820 6497 3869 6509
rect 3820 6477 3831 6497
rect 3851 6477 3869 6497
rect 3820 6467 3869 6477
rect 3919 6493 3963 6509
rect 3919 6473 3934 6493
rect 3954 6473 3963 6493
rect 3919 6467 3963 6473
rect 4033 6493 4077 6509
rect 4033 6473 4042 6493
rect 4062 6473 4077 6493
rect 4033 6467 4077 6473
rect 4127 6497 4176 6509
rect 4127 6477 4145 6497
rect 4165 6477 4176 6497
rect 4127 6467 4176 6477
rect 4241 6493 4285 6509
rect 4241 6473 4250 6493
rect 4270 6473 4285 6493
rect 4241 6467 4285 6473
rect 4335 6497 4384 6509
rect 4335 6477 4353 6497
rect 4373 6477 4384 6497
rect 4335 6467 4384 6477
rect 4454 6493 4498 6509
rect 4454 6473 4463 6493
rect 4483 6473 4498 6493
rect 4454 6467 4498 6473
rect 4548 6497 4597 6509
rect 4548 6477 4566 6497
rect 4586 6477 4597 6497
rect 4548 6467 4597 6477
rect 8876 6538 8925 6550
rect 8876 6518 8887 6538
rect 8907 6518 8925 6538
rect 8876 6508 8925 6518
rect 8975 6534 9019 6550
rect 8975 6514 8990 6534
rect 9010 6514 9019 6534
rect 8975 6508 9019 6514
rect 9089 6534 9133 6550
rect 9089 6514 9098 6534
rect 9118 6514 9133 6534
rect 9089 6508 9133 6514
rect 9183 6538 9232 6550
rect 9183 6518 9201 6538
rect 9221 6518 9232 6538
rect 9183 6508 9232 6518
rect 9297 6534 9341 6550
rect 9297 6514 9306 6534
rect 9326 6514 9341 6534
rect 9297 6508 9341 6514
rect 9391 6538 9440 6550
rect 9391 6518 9409 6538
rect 9429 6518 9440 6538
rect 9391 6508 9440 6518
rect 9510 6534 9554 6550
rect 9510 6514 9519 6534
rect 9539 6514 9554 6534
rect 9510 6508 9554 6514
rect 9604 6538 9653 6550
rect 9604 6518 9622 6538
rect 9642 6518 9653 6538
rect 9604 6508 9653 6518
rect 11303 6574 11352 6584
rect 11303 6554 11314 6574
rect 11334 6554 11352 6574
rect 11303 6542 11352 6554
rect 11402 6578 11446 6584
rect 11402 6558 11417 6578
rect 11437 6558 11446 6578
rect 11402 6542 11446 6558
rect 11516 6574 11565 6584
rect 11516 6554 11527 6574
rect 11547 6554 11565 6574
rect 11516 6542 11565 6554
rect 11615 6578 11659 6584
rect 11615 6558 11630 6578
rect 11650 6558 11659 6578
rect 11615 6542 11659 6558
rect 11724 6574 11773 6584
rect 11724 6554 11735 6574
rect 11755 6554 11773 6574
rect 11724 6542 11773 6554
rect 11823 6578 11867 6584
rect 11823 6558 11838 6578
rect 11858 6558 11867 6578
rect 11823 6542 11867 6558
rect 11937 6578 11981 6584
rect 11937 6558 11946 6578
rect 11966 6558 11981 6578
rect 11937 6542 11981 6558
rect 12031 6574 12080 6584
rect 12031 6554 12049 6574
rect 12069 6554 12080 6574
rect 12031 6542 12080 6554
rect 17969 6787 18018 6799
rect 17969 6767 17980 6787
rect 18000 6767 18018 6787
rect 17969 6757 18018 6767
rect 18068 6783 18112 6799
rect 18068 6763 18083 6783
rect 18103 6763 18112 6783
rect 18068 6757 18112 6763
rect 18182 6783 18226 6799
rect 18182 6763 18191 6783
rect 18211 6763 18226 6783
rect 18182 6757 18226 6763
rect 18276 6787 18325 6799
rect 18276 6767 18294 6787
rect 18314 6767 18325 6787
rect 18276 6757 18325 6767
rect 18390 6783 18434 6799
rect 18390 6763 18399 6783
rect 18419 6763 18434 6783
rect 18390 6757 18434 6763
rect 18484 6787 18533 6799
rect 18484 6767 18502 6787
rect 18522 6767 18533 6787
rect 18484 6757 18533 6767
rect 18603 6783 18647 6799
rect 18603 6763 18612 6783
rect 18632 6763 18647 6783
rect 18603 6757 18647 6763
rect 18697 6787 18746 6799
rect 18697 6767 18715 6787
rect 18735 6767 18746 6787
rect 18697 6757 18746 6767
rect 16359 6615 16408 6625
rect 16359 6595 16370 6615
rect 16390 6595 16408 6615
rect 16359 6583 16408 6595
rect 16458 6619 16502 6625
rect 16458 6599 16473 6619
rect 16493 6599 16502 6619
rect 16458 6583 16502 6599
rect 16572 6615 16621 6625
rect 16572 6595 16583 6615
rect 16603 6595 16621 6615
rect 16572 6583 16621 6595
rect 16671 6619 16715 6625
rect 16671 6599 16686 6619
rect 16706 6599 16715 6619
rect 16671 6583 16715 6599
rect 16780 6615 16829 6625
rect 16780 6595 16791 6615
rect 16811 6595 16829 6615
rect 16780 6583 16829 6595
rect 16879 6619 16923 6625
rect 16879 6599 16894 6619
rect 16914 6599 16923 6619
rect 16879 6583 16923 6599
rect 16993 6619 17037 6625
rect 16993 6599 17002 6619
rect 17022 6599 17037 6619
rect 16993 6583 17037 6599
rect 17087 6615 17136 6625
rect 17087 6595 17105 6615
rect 17125 6595 17136 6615
rect 17087 6583 17136 6595
rect 13851 6502 13900 6514
rect 13851 6482 13862 6502
rect 13882 6482 13900 6502
rect 13851 6472 13900 6482
rect 13950 6498 13994 6514
rect 13950 6478 13965 6498
rect 13985 6478 13994 6498
rect 13950 6472 13994 6478
rect 14064 6498 14108 6514
rect 14064 6478 14073 6498
rect 14093 6478 14108 6498
rect 14064 6472 14108 6478
rect 14158 6502 14207 6514
rect 14158 6482 14176 6502
rect 14196 6482 14207 6502
rect 14158 6472 14207 6482
rect 14272 6498 14316 6514
rect 14272 6478 14281 6498
rect 14301 6478 14316 6498
rect 14272 6472 14316 6478
rect 14366 6502 14415 6514
rect 14366 6482 14384 6502
rect 14404 6482 14415 6502
rect 14366 6472 14415 6482
rect 14485 6498 14529 6514
rect 14485 6478 14494 6498
rect 14514 6478 14529 6498
rect 14485 6472 14529 6478
rect 14579 6502 14628 6514
rect 14579 6482 14597 6502
rect 14617 6482 14628 6502
rect 14579 6472 14628 6482
rect 5389 6300 5438 6310
rect 5389 6280 5400 6300
rect 5420 6280 5438 6300
rect 333 6259 382 6269
rect 333 6239 344 6259
rect 364 6239 382 6259
rect 333 6227 382 6239
rect 432 6263 476 6269
rect 432 6243 447 6263
rect 467 6243 476 6263
rect 432 6227 476 6243
rect 546 6259 595 6269
rect 546 6239 557 6259
rect 577 6239 595 6259
rect 546 6227 595 6239
rect 645 6263 689 6269
rect 645 6243 660 6263
rect 680 6243 689 6263
rect 645 6227 689 6243
rect 754 6259 803 6269
rect 754 6239 765 6259
rect 785 6239 803 6259
rect 754 6227 803 6239
rect 853 6263 897 6269
rect 853 6243 868 6263
rect 888 6243 897 6263
rect 853 6227 897 6243
rect 967 6263 1011 6269
rect 967 6243 976 6263
rect 996 6243 1011 6263
rect 967 6227 1011 6243
rect 1061 6259 1110 6269
rect 1061 6239 1079 6259
rect 1099 6239 1110 6259
rect 1061 6227 1110 6239
rect 2742 6230 2791 6242
rect 2742 6210 2753 6230
rect 2773 6210 2791 6230
rect 2742 6200 2791 6210
rect 2841 6226 2885 6242
rect 2841 6206 2856 6226
rect 2876 6206 2885 6226
rect 2841 6200 2885 6206
rect 2955 6226 2999 6242
rect 2955 6206 2964 6226
rect 2984 6206 2999 6226
rect 2955 6200 2999 6206
rect 3049 6230 3098 6242
rect 3049 6210 3067 6230
rect 3087 6210 3098 6230
rect 3049 6200 3098 6210
rect 3163 6226 3207 6242
rect 3163 6206 3172 6226
rect 3192 6206 3207 6226
rect 3163 6200 3207 6206
rect 3257 6230 3306 6242
rect 3257 6210 3275 6230
rect 3295 6210 3306 6230
rect 3257 6200 3306 6210
rect 3376 6226 3420 6242
rect 3376 6206 3385 6226
rect 3405 6206 3420 6226
rect 3376 6200 3420 6206
rect 3470 6230 3519 6242
rect 3470 6210 3488 6230
rect 3508 6210 3519 6230
rect 3470 6200 3519 6210
rect 5389 6268 5438 6280
rect 5488 6304 5532 6310
rect 5488 6284 5503 6304
rect 5523 6284 5532 6304
rect 5488 6268 5532 6284
rect 5602 6300 5651 6310
rect 5602 6280 5613 6300
rect 5633 6280 5651 6300
rect 5602 6268 5651 6280
rect 5701 6304 5745 6310
rect 5701 6284 5716 6304
rect 5736 6284 5745 6304
rect 5701 6268 5745 6284
rect 5810 6300 5859 6310
rect 5810 6280 5821 6300
rect 5841 6280 5859 6300
rect 5810 6268 5859 6280
rect 5909 6304 5953 6310
rect 5909 6284 5924 6304
rect 5944 6284 5953 6304
rect 5909 6268 5953 6284
rect 6023 6304 6067 6310
rect 6023 6284 6032 6304
rect 6052 6284 6067 6304
rect 6023 6268 6067 6284
rect 6117 6300 6166 6310
rect 6117 6280 6135 6300
rect 6155 6280 6166 6300
rect 6117 6268 6166 6280
rect 7798 6271 7847 6283
rect 7798 6251 7809 6271
rect 7829 6251 7847 6271
rect 7798 6241 7847 6251
rect 7897 6267 7941 6283
rect 7897 6247 7912 6267
rect 7932 6247 7941 6267
rect 7897 6241 7941 6247
rect 8011 6267 8055 6283
rect 8011 6247 8020 6267
rect 8040 6247 8055 6267
rect 8011 6241 8055 6247
rect 8105 6271 8154 6283
rect 8105 6251 8123 6271
rect 8143 6251 8154 6271
rect 8105 6241 8154 6251
rect 8219 6267 8263 6283
rect 8219 6247 8228 6267
rect 8248 6247 8263 6267
rect 8219 6241 8263 6247
rect 8313 6271 8362 6283
rect 8313 6251 8331 6271
rect 8351 6251 8362 6271
rect 8313 6241 8362 6251
rect 8432 6267 8476 6283
rect 8432 6247 8441 6267
rect 8461 6247 8476 6267
rect 8432 6241 8476 6247
rect 8526 6271 8575 6283
rect 8526 6251 8544 6271
rect 8564 6251 8575 6271
rect 8526 6241 8575 6251
rect 18907 6543 18956 6555
rect 18907 6523 18918 6543
rect 18938 6523 18956 6543
rect 18907 6513 18956 6523
rect 19006 6539 19050 6555
rect 19006 6519 19021 6539
rect 19041 6519 19050 6539
rect 19006 6513 19050 6519
rect 19120 6539 19164 6555
rect 19120 6519 19129 6539
rect 19149 6519 19164 6539
rect 19120 6513 19164 6519
rect 19214 6543 19263 6555
rect 19214 6523 19232 6543
rect 19252 6523 19263 6543
rect 19214 6513 19263 6523
rect 19328 6539 19372 6555
rect 19328 6519 19337 6539
rect 19357 6519 19372 6539
rect 19328 6513 19372 6519
rect 19422 6543 19471 6555
rect 19422 6523 19440 6543
rect 19460 6523 19471 6543
rect 19422 6513 19471 6523
rect 19541 6539 19585 6555
rect 19541 6519 19550 6539
rect 19570 6519 19585 6539
rect 19541 6513 19585 6519
rect 19635 6543 19684 6555
rect 19635 6523 19653 6543
rect 19673 6523 19684 6543
rect 19635 6513 19684 6523
rect 15420 6305 15469 6315
rect 15420 6285 15431 6305
rect 15451 6285 15469 6305
rect 10364 6264 10413 6274
rect 10364 6244 10375 6264
rect 10395 6244 10413 6264
rect 10364 6232 10413 6244
rect 10463 6268 10507 6274
rect 10463 6248 10478 6268
rect 10498 6248 10507 6268
rect 10463 6232 10507 6248
rect 10577 6264 10626 6274
rect 10577 6244 10588 6264
rect 10608 6244 10626 6264
rect 10577 6232 10626 6244
rect 10676 6268 10720 6274
rect 10676 6248 10691 6268
rect 10711 6248 10720 6268
rect 10676 6232 10720 6248
rect 10785 6264 10834 6274
rect 10785 6244 10796 6264
rect 10816 6244 10834 6264
rect 10785 6232 10834 6244
rect 10884 6268 10928 6274
rect 10884 6248 10899 6268
rect 10919 6248 10928 6268
rect 10884 6232 10928 6248
rect 10998 6268 11042 6274
rect 10998 6248 11007 6268
rect 11027 6248 11042 6268
rect 10998 6232 11042 6248
rect 11092 6264 11141 6274
rect 11092 6244 11110 6264
rect 11130 6244 11141 6264
rect 11092 6232 11141 6244
rect 12773 6235 12822 6247
rect 12773 6215 12784 6235
rect 12804 6215 12822 6235
rect 12773 6205 12822 6215
rect 12872 6231 12916 6247
rect 12872 6211 12887 6231
rect 12907 6211 12916 6231
rect 12872 6205 12916 6211
rect 12986 6231 13030 6247
rect 12986 6211 12995 6231
rect 13015 6211 13030 6231
rect 12986 6205 13030 6211
rect 13080 6235 13129 6247
rect 13080 6215 13098 6235
rect 13118 6215 13129 6235
rect 13080 6205 13129 6215
rect 13194 6231 13238 6247
rect 13194 6211 13203 6231
rect 13223 6211 13238 6231
rect 13194 6205 13238 6211
rect 13288 6235 13337 6247
rect 13288 6215 13306 6235
rect 13326 6215 13337 6235
rect 13288 6205 13337 6215
rect 13407 6231 13451 6247
rect 13407 6211 13416 6231
rect 13436 6211 13451 6231
rect 13407 6205 13451 6211
rect 13501 6235 13550 6247
rect 13501 6215 13519 6235
rect 13539 6215 13550 6235
rect 13501 6205 13550 6215
rect 15420 6273 15469 6285
rect 15519 6309 15563 6315
rect 15519 6289 15534 6309
rect 15554 6289 15563 6309
rect 15519 6273 15563 6289
rect 15633 6305 15682 6315
rect 15633 6285 15644 6305
rect 15664 6285 15682 6305
rect 15633 6273 15682 6285
rect 15732 6309 15776 6315
rect 15732 6289 15747 6309
rect 15767 6289 15776 6309
rect 15732 6273 15776 6289
rect 15841 6305 15890 6315
rect 15841 6285 15852 6305
rect 15872 6285 15890 6305
rect 15841 6273 15890 6285
rect 15940 6309 15984 6315
rect 15940 6289 15955 6309
rect 15975 6289 15984 6309
rect 15940 6273 15984 6289
rect 16054 6309 16098 6315
rect 16054 6289 16063 6309
rect 16083 6289 16098 6309
rect 16054 6273 16098 6289
rect 16148 6305 16197 6315
rect 16148 6285 16166 6305
rect 16186 6285 16197 6305
rect 16148 6273 16197 6285
rect 17829 6276 17878 6288
rect 17829 6256 17840 6276
rect 17860 6256 17878 6276
rect 17829 6246 17878 6256
rect 17928 6272 17972 6288
rect 17928 6252 17943 6272
rect 17963 6252 17972 6272
rect 17928 6246 17972 6252
rect 18042 6272 18086 6288
rect 18042 6252 18051 6272
rect 18071 6252 18086 6272
rect 18042 6246 18086 6252
rect 18136 6276 18185 6288
rect 18136 6256 18154 6276
rect 18174 6256 18185 6276
rect 18136 6246 18185 6256
rect 18250 6272 18294 6288
rect 18250 6252 18259 6272
rect 18279 6252 18294 6272
rect 18250 6246 18294 6252
rect 18344 6276 18393 6288
rect 18344 6256 18362 6276
rect 18382 6256 18393 6276
rect 18344 6246 18393 6256
rect 18463 6272 18507 6288
rect 18463 6252 18472 6272
rect 18492 6252 18507 6272
rect 18463 6246 18507 6252
rect 18557 6276 18606 6288
rect 18557 6256 18575 6276
rect 18595 6256 18606 6276
rect 18557 6246 18606 6256
rect 1413 5977 1462 5987
rect 1413 5957 1424 5977
rect 1444 5957 1462 5977
rect 1413 5945 1462 5957
rect 1512 5981 1556 5987
rect 1512 5961 1527 5981
rect 1547 5961 1556 5981
rect 1512 5945 1556 5961
rect 1626 5977 1675 5987
rect 1626 5957 1637 5977
rect 1657 5957 1675 5977
rect 1626 5945 1675 5957
rect 1725 5981 1769 5987
rect 1725 5961 1740 5981
rect 1760 5961 1769 5981
rect 1725 5945 1769 5961
rect 1834 5977 1883 5987
rect 1834 5957 1845 5977
rect 1865 5957 1883 5977
rect 1834 5945 1883 5957
rect 1933 5981 1977 5987
rect 1933 5961 1948 5981
rect 1968 5961 1977 5981
rect 1933 5945 1977 5961
rect 2047 5981 2091 5987
rect 2047 5961 2056 5981
rect 2076 5961 2091 5981
rect 2047 5945 2091 5961
rect 2141 5977 2190 5987
rect 2141 5957 2159 5977
rect 2179 5957 2190 5977
rect 2141 5945 2190 5957
rect 3822 5948 3871 5960
rect 3822 5928 3833 5948
rect 3853 5928 3871 5948
rect 3822 5918 3871 5928
rect 3921 5944 3965 5960
rect 3921 5924 3936 5944
rect 3956 5924 3965 5944
rect 3921 5918 3965 5924
rect 4035 5944 4079 5960
rect 4035 5924 4044 5944
rect 4064 5924 4079 5944
rect 4035 5918 4079 5924
rect 4129 5948 4178 5960
rect 4129 5928 4147 5948
rect 4167 5928 4178 5948
rect 4129 5918 4178 5928
rect 4243 5944 4287 5960
rect 4243 5924 4252 5944
rect 4272 5924 4287 5944
rect 4243 5918 4287 5924
rect 4337 5948 4386 5960
rect 4337 5928 4355 5948
rect 4375 5928 4386 5948
rect 4337 5918 4386 5928
rect 4456 5944 4500 5960
rect 4456 5924 4465 5944
rect 4485 5924 4500 5944
rect 4456 5918 4500 5924
rect 4550 5948 4599 5960
rect 6469 6018 6518 6028
rect 6469 5998 6480 6018
rect 6500 5998 6518 6018
rect 6469 5986 6518 5998
rect 6568 6022 6612 6028
rect 6568 6002 6583 6022
rect 6603 6002 6612 6022
rect 6568 5986 6612 6002
rect 6682 6018 6731 6028
rect 6682 5998 6693 6018
rect 6713 5998 6731 6018
rect 6682 5986 6731 5998
rect 6781 6022 6825 6028
rect 6781 6002 6796 6022
rect 6816 6002 6825 6022
rect 6781 5986 6825 6002
rect 6890 6018 6939 6028
rect 6890 5998 6901 6018
rect 6921 5998 6939 6018
rect 6890 5986 6939 5998
rect 6989 6022 7033 6028
rect 6989 6002 7004 6022
rect 7024 6002 7033 6022
rect 6989 5986 7033 6002
rect 7103 6022 7147 6028
rect 7103 6002 7112 6022
rect 7132 6002 7147 6022
rect 7103 5986 7147 6002
rect 7197 6018 7246 6028
rect 7197 5998 7215 6018
rect 7235 5998 7246 6018
rect 7197 5986 7246 5998
rect 8878 5989 8927 6001
rect 8878 5969 8889 5989
rect 8909 5969 8927 5989
rect 8878 5959 8927 5969
rect 8977 5985 9021 6001
rect 8977 5965 8992 5985
rect 9012 5965 9021 5985
rect 8977 5959 9021 5965
rect 9091 5985 9135 6001
rect 9091 5965 9100 5985
rect 9120 5965 9135 5985
rect 9091 5959 9135 5965
rect 9185 5989 9234 6001
rect 9185 5969 9203 5989
rect 9223 5969 9234 5989
rect 9185 5959 9234 5969
rect 9299 5985 9343 6001
rect 9299 5965 9308 5985
rect 9328 5965 9343 5985
rect 9299 5959 9343 5965
rect 9393 5989 9442 6001
rect 9393 5969 9411 5989
rect 9431 5969 9442 5989
rect 9393 5959 9442 5969
rect 9512 5985 9556 6001
rect 9512 5965 9521 5985
rect 9541 5965 9556 5985
rect 9512 5959 9556 5965
rect 9606 5989 9655 6001
rect 9606 5969 9624 5989
rect 9644 5969 9655 5989
rect 9606 5959 9655 5969
rect 4550 5928 4568 5948
rect 4588 5928 4599 5948
rect 4550 5918 4599 5928
rect 335 5710 384 5720
rect 335 5690 346 5710
rect 366 5690 384 5710
rect 335 5678 384 5690
rect 434 5714 478 5720
rect 434 5694 449 5714
rect 469 5694 478 5714
rect 434 5678 478 5694
rect 548 5710 597 5720
rect 548 5690 559 5710
rect 579 5690 597 5710
rect 548 5678 597 5690
rect 647 5714 691 5720
rect 647 5694 662 5714
rect 682 5694 691 5714
rect 647 5678 691 5694
rect 756 5710 805 5720
rect 756 5690 767 5710
rect 787 5690 805 5710
rect 756 5678 805 5690
rect 855 5714 899 5720
rect 855 5694 870 5714
rect 890 5694 899 5714
rect 855 5678 899 5694
rect 969 5714 1013 5720
rect 969 5694 978 5714
rect 998 5694 1013 5714
rect 969 5678 1013 5694
rect 1063 5710 1112 5720
rect 1063 5690 1081 5710
rect 1101 5690 1112 5710
rect 1063 5678 1112 5690
rect 11444 5982 11493 5992
rect 11444 5962 11455 5982
rect 11475 5962 11493 5982
rect 11444 5950 11493 5962
rect 11543 5986 11587 5992
rect 11543 5966 11558 5986
rect 11578 5966 11587 5986
rect 11543 5950 11587 5966
rect 11657 5982 11706 5992
rect 11657 5962 11668 5982
rect 11688 5962 11706 5982
rect 11657 5950 11706 5962
rect 11756 5986 11800 5992
rect 11756 5966 11771 5986
rect 11791 5966 11800 5986
rect 11756 5950 11800 5966
rect 11865 5982 11914 5992
rect 11865 5962 11876 5982
rect 11896 5962 11914 5982
rect 11865 5950 11914 5962
rect 11964 5986 12008 5992
rect 11964 5966 11979 5986
rect 11999 5966 12008 5986
rect 11964 5950 12008 5966
rect 12078 5986 12122 5992
rect 12078 5966 12087 5986
rect 12107 5966 12122 5986
rect 12078 5950 12122 5966
rect 12172 5982 12221 5992
rect 12172 5962 12190 5982
rect 12210 5962 12221 5982
rect 12172 5950 12221 5962
rect 13853 5953 13902 5965
rect 13853 5933 13864 5953
rect 13884 5933 13902 5953
rect 13853 5923 13902 5933
rect 13952 5949 13996 5965
rect 13952 5929 13967 5949
rect 13987 5929 13996 5949
rect 13952 5923 13996 5929
rect 14066 5949 14110 5965
rect 14066 5929 14075 5949
rect 14095 5929 14110 5949
rect 14066 5923 14110 5929
rect 14160 5953 14209 5965
rect 14160 5933 14178 5953
rect 14198 5933 14209 5953
rect 14160 5923 14209 5933
rect 14274 5949 14318 5965
rect 14274 5929 14283 5949
rect 14303 5929 14318 5949
rect 14274 5923 14318 5929
rect 14368 5953 14417 5965
rect 14368 5933 14386 5953
rect 14406 5933 14417 5953
rect 14368 5923 14417 5933
rect 14487 5949 14531 5965
rect 14487 5929 14496 5949
rect 14516 5929 14531 5949
rect 14487 5923 14531 5929
rect 14581 5953 14630 5965
rect 16500 6023 16549 6033
rect 16500 6003 16511 6023
rect 16531 6003 16549 6023
rect 16500 5991 16549 6003
rect 16599 6027 16643 6033
rect 16599 6007 16614 6027
rect 16634 6007 16643 6027
rect 16599 5991 16643 6007
rect 16713 6023 16762 6033
rect 16713 6003 16724 6023
rect 16744 6003 16762 6023
rect 16713 5991 16762 6003
rect 16812 6027 16856 6033
rect 16812 6007 16827 6027
rect 16847 6007 16856 6027
rect 16812 5991 16856 6007
rect 16921 6023 16970 6033
rect 16921 6003 16932 6023
rect 16952 6003 16970 6023
rect 16921 5991 16970 6003
rect 17020 6027 17064 6033
rect 17020 6007 17035 6027
rect 17055 6007 17064 6027
rect 17020 5991 17064 6007
rect 17134 6027 17178 6033
rect 17134 6007 17143 6027
rect 17163 6007 17178 6027
rect 17134 5991 17178 6007
rect 17228 6023 17277 6033
rect 17228 6003 17246 6023
rect 17266 6003 17277 6023
rect 17228 5991 17277 6003
rect 18909 5994 18958 6006
rect 18909 5974 18920 5994
rect 18940 5974 18958 5994
rect 18909 5964 18958 5974
rect 19008 5990 19052 6006
rect 19008 5970 19023 5990
rect 19043 5970 19052 5990
rect 19008 5964 19052 5970
rect 19122 5990 19166 6006
rect 19122 5970 19131 5990
rect 19151 5970 19166 5990
rect 19122 5964 19166 5970
rect 19216 5994 19265 6006
rect 19216 5974 19234 5994
rect 19254 5974 19265 5994
rect 19216 5964 19265 5974
rect 19330 5990 19374 6006
rect 19330 5970 19339 5990
rect 19359 5970 19374 5990
rect 19330 5964 19374 5970
rect 19424 5994 19473 6006
rect 19424 5974 19442 5994
rect 19462 5974 19473 5994
rect 19424 5964 19473 5974
rect 19543 5990 19587 6006
rect 19543 5970 19552 5990
rect 19572 5970 19587 5990
rect 19543 5964 19587 5970
rect 19637 5994 19686 6006
rect 19637 5974 19655 5994
rect 19675 5974 19686 5994
rect 19637 5964 19686 5974
rect 14581 5933 14599 5953
rect 14619 5933 14630 5953
rect 14581 5923 14630 5933
rect 5391 5751 5440 5761
rect 5391 5731 5402 5751
rect 5422 5731 5440 5751
rect 5391 5719 5440 5731
rect 5490 5755 5534 5761
rect 5490 5735 5505 5755
rect 5525 5735 5534 5755
rect 5490 5719 5534 5735
rect 5604 5751 5653 5761
rect 5604 5731 5615 5751
rect 5635 5731 5653 5751
rect 5604 5719 5653 5731
rect 5703 5755 5747 5761
rect 5703 5735 5718 5755
rect 5738 5735 5747 5755
rect 5703 5719 5747 5735
rect 5812 5751 5861 5761
rect 5812 5731 5823 5751
rect 5843 5731 5861 5751
rect 5812 5719 5861 5731
rect 5911 5755 5955 5761
rect 5911 5735 5926 5755
rect 5946 5735 5955 5755
rect 5911 5719 5955 5735
rect 6025 5755 6069 5761
rect 6025 5735 6034 5755
rect 6054 5735 6069 5755
rect 6025 5719 6069 5735
rect 6119 5751 6168 5761
rect 6119 5731 6137 5751
rect 6157 5731 6168 5751
rect 6119 5719 6168 5731
rect 2883 5638 2932 5650
rect 2883 5618 2894 5638
rect 2914 5618 2932 5638
rect 2883 5608 2932 5618
rect 2982 5634 3026 5650
rect 2982 5614 2997 5634
rect 3017 5614 3026 5634
rect 2982 5608 3026 5614
rect 3096 5634 3140 5650
rect 3096 5614 3105 5634
rect 3125 5614 3140 5634
rect 3096 5608 3140 5614
rect 3190 5638 3239 5650
rect 3190 5618 3208 5638
rect 3228 5618 3239 5638
rect 3190 5608 3239 5618
rect 3304 5634 3348 5650
rect 3304 5614 3313 5634
rect 3333 5614 3348 5634
rect 3304 5608 3348 5614
rect 3398 5638 3447 5650
rect 3398 5618 3416 5638
rect 3436 5618 3447 5638
rect 3398 5608 3447 5618
rect 3517 5634 3561 5650
rect 3517 5614 3526 5634
rect 3546 5614 3561 5634
rect 3517 5608 3561 5614
rect 3611 5638 3660 5650
rect 3611 5618 3629 5638
rect 3649 5618 3660 5638
rect 3611 5608 3660 5618
rect 1273 5466 1322 5476
rect 1273 5446 1284 5466
rect 1304 5446 1322 5466
rect 1273 5434 1322 5446
rect 1372 5470 1416 5476
rect 1372 5450 1387 5470
rect 1407 5450 1416 5470
rect 1372 5434 1416 5450
rect 1486 5466 1535 5476
rect 1486 5446 1497 5466
rect 1517 5446 1535 5466
rect 1486 5434 1535 5446
rect 1585 5470 1629 5476
rect 1585 5450 1600 5470
rect 1620 5450 1629 5470
rect 1585 5434 1629 5450
rect 1694 5466 1743 5476
rect 1694 5446 1705 5466
rect 1725 5446 1743 5466
rect 1694 5434 1743 5446
rect 1793 5470 1837 5476
rect 1793 5450 1808 5470
rect 1828 5450 1837 5470
rect 1793 5434 1837 5450
rect 1907 5470 1951 5476
rect 1907 5450 1916 5470
rect 1936 5450 1951 5470
rect 1907 5434 1951 5450
rect 2001 5466 2050 5476
rect 2001 5446 2019 5466
rect 2039 5446 2050 5466
rect 2001 5434 2050 5446
rect 7939 5679 7988 5691
rect 7939 5659 7950 5679
rect 7970 5659 7988 5679
rect 7939 5649 7988 5659
rect 8038 5675 8082 5691
rect 8038 5655 8053 5675
rect 8073 5655 8082 5675
rect 8038 5649 8082 5655
rect 8152 5675 8196 5691
rect 8152 5655 8161 5675
rect 8181 5655 8196 5675
rect 8152 5649 8196 5655
rect 8246 5679 8295 5691
rect 8246 5659 8264 5679
rect 8284 5659 8295 5679
rect 8246 5649 8295 5659
rect 8360 5675 8404 5691
rect 8360 5655 8369 5675
rect 8389 5655 8404 5675
rect 8360 5649 8404 5655
rect 8454 5679 8503 5691
rect 8454 5659 8472 5679
rect 8492 5659 8503 5679
rect 8454 5649 8503 5659
rect 8573 5675 8617 5691
rect 8573 5655 8582 5675
rect 8602 5655 8617 5675
rect 8573 5649 8617 5655
rect 8667 5679 8716 5691
rect 8667 5659 8685 5679
rect 8705 5659 8716 5679
rect 8667 5649 8716 5659
rect 10366 5715 10415 5725
rect 10366 5695 10377 5715
rect 10397 5695 10415 5715
rect 10366 5683 10415 5695
rect 10465 5719 10509 5725
rect 10465 5699 10480 5719
rect 10500 5699 10509 5719
rect 10465 5683 10509 5699
rect 10579 5715 10628 5725
rect 10579 5695 10590 5715
rect 10610 5695 10628 5715
rect 10579 5683 10628 5695
rect 10678 5719 10722 5725
rect 10678 5699 10693 5719
rect 10713 5699 10722 5719
rect 10678 5683 10722 5699
rect 10787 5715 10836 5725
rect 10787 5695 10798 5715
rect 10818 5695 10836 5715
rect 10787 5683 10836 5695
rect 10886 5719 10930 5725
rect 10886 5699 10901 5719
rect 10921 5699 10930 5719
rect 10886 5683 10930 5699
rect 11000 5719 11044 5725
rect 11000 5699 11009 5719
rect 11029 5699 11044 5719
rect 11000 5683 11044 5699
rect 11094 5715 11143 5725
rect 11094 5695 11112 5715
rect 11132 5695 11143 5715
rect 11094 5683 11143 5695
rect 15422 5756 15471 5766
rect 15422 5736 15433 5756
rect 15453 5736 15471 5756
rect 15422 5724 15471 5736
rect 15521 5760 15565 5766
rect 15521 5740 15536 5760
rect 15556 5740 15565 5760
rect 15521 5724 15565 5740
rect 15635 5756 15684 5766
rect 15635 5736 15646 5756
rect 15666 5736 15684 5756
rect 15635 5724 15684 5736
rect 15734 5760 15778 5766
rect 15734 5740 15749 5760
rect 15769 5740 15778 5760
rect 15734 5724 15778 5740
rect 15843 5756 15892 5766
rect 15843 5736 15854 5756
rect 15874 5736 15892 5756
rect 15843 5724 15892 5736
rect 15942 5760 15986 5766
rect 15942 5740 15957 5760
rect 15977 5740 15986 5760
rect 15942 5724 15986 5740
rect 16056 5760 16100 5766
rect 16056 5740 16065 5760
rect 16085 5740 16100 5760
rect 16056 5724 16100 5740
rect 16150 5756 16199 5766
rect 16150 5736 16168 5756
rect 16188 5736 16199 5756
rect 16150 5724 16199 5736
rect 6329 5507 6378 5517
rect 6329 5487 6340 5507
rect 6360 5487 6378 5507
rect 6329 5475 6378 5487
rect 6428 5511 6472 5517
rect 6428 5491 6443 5511
rect 6463 5491 6472 5511
rect 6428 5475 6472 5491
rect 6542 5507 6591 5517
rect 6542 5487 6553 5507
rect 6573 5487 6591 5507
rect 6542 5475 6591 5487
rect 6641 5511 6685 5517
rect 6641 5491 6656 5511
rect 6676 5491 6685 5511
rect 6641 5475 6685 5491
rect 6750 5507 6799 5517
rect 6750 5487 6761 5507
rect 6781 5487 6799 5507
rect 6750 5475 6799 5487
rect 6849 5511 6893 5517
rect 6849 5491 6864 5511
rect 6884 5491 6893 5511
rect 6849 5475 6893 5491
rect 6963 5511 7007 5517
rect 6963 5491 6972 5511
rect 6992 5491 7007 5511
rect 6963 5475 7007 5491
rect 7057 5507 7106 5517
rect 7057 5487 7075 5507
rect 7095 5487 7106 5507
rect 7057 5475 7106 5487
rect 12914 5643 12963 5655
rect 12914 5623 12925 5643
rect 12945 5623 12963 5643
rect 12914 5613 12963 5623
rect 13013 5639 13057 5655
rect 13013 5619 13028 5639
rect 13048 5619 13057 5639
rect 13013 5613 13057 5619
rect 13127 5639 13171 5655
rect 13127 5619 13136 5639
rect 13156 5619 13171 5639
rect 13127 5613 13171 5619
rect 13221 5643 13270 5655
rect 13221 5623 13239 5643
rect 13259 5623 13270 5643
rect 13221 5613 13270 5623
rect 13335 5639 13379 5655
rect 13335 5619 13344 5639
rect 13364 5619 13379 5639
rect 13335 5613 13379 5619
rect 13429 5643 13478 5655
rect 13429 5623 13447 5643
rect 13467 5623 13478 5643
rect 13429 5613 13478 5623
rect 13548 5639 13592 5655
rect 13548 5619 13557 5639
rect 13577 5619 13592 5639
rect 13548 5613 13592 5619
rect 13642 5643 13691 5655
rect 13642 5623 13660 5643
rect 13680 5623 13691 5643
rect 13642 5613 13691 5623
rect 3821 5394 3870 5406
rect 3821 5374 3832 5394
rect 3852 5374 3870 5394
rect 3821 5364 3870 5374
rect 3920 5390 3964 5406
rect 3920 5370 3935 5390
rect 3955 5370 3964 5390
rect 3920 5364 3964 5370
rect 4034 5390 4078 5406
rect 4034 5370 4043 5390
rect 4063 5370 4078 5390
rect 4034 5364 4078 5370
rect 4128 5394 4177 5406
rect 4128 5374 4146 5394
rect 4166 5374 4177 5394
rect 4128 5364 4177 5374
rect 4242 5390 4286 5406
rect 4242 5370 4251 5390
rect 4271 5370 4286 5390
rect 4242 5364 4286 5370
rect 4336 5394 4385 5406
rect 4336 5374 4354 5394
rect 4374 5374 4385 5394
rect 4336 5364 4385 5374
rect 4455 5390 4499 5406
rect 4455 5370 4464 5390
rect 4484 5370 4499 5390
rect 4455 5364 4499 5370
rect 4549 5394 4598 5406
rect 4549 5374 4567 5394
rect 4587 5374 4598 5394
rect 4549 5364 4598 5374
rect 8877 5435 8926 5447
rect 8877 5415 8888 5435
rect 8908 5415 8926 5435
rect 8877 5405 8926 5415
rect 8976 5431 9020 5447
rect 8976 5411 8991 5431
rect 9011 5411 9020 5431
rect 8976 5405 9020 5411
rect 9090 5431 9134 5447
rect 9090 5411 9099 5431
rect 9119 5411 9134 5431
rect 9090 5405 9134 5411
rect 9184 5435 9233 5447
rect 9184 5415 9202 5435
rect 9222 5415 9233 5435
rect 9184 5405 9233 5415
rect 9298 5431 9342 5447
rect 9298 5411 9307 5431
rect 9327 5411 9342 5431
rect 9298 5405 9342 5411
rect 9392 5435 9441 5447
rect 9392 5415 9410 5435
rect 9430 5415 9441 5435
rect 9392 5405 9441 5415
rect 9511 5431 9555 5447
rect 9511 5411 9520 5431
rect 9540 5411 9555 5431
rect 9511 5405 9555 5411
rect 9605 5435 9654 5447
rect 9605 5415 9623 5435
rect 9643 5415 9654 5435
rect 9605 5405 9654 5415
rect 11304 5471 11353 5481
rect 11304 5451 11315 5471
rect 11335 5451 11353 5471
rect 11304 5439 11353 5451
rect 11403 5475 11447 5481
rect 11403 5455 11418 5475
rect 11438 5455 11447 5475
rect 11403 5439 11447 5455
rect 11517 5471 11566 5481
rect 11517 5451 11528 5471
rect 11548 5451 11566 5471
rect 11517 5439 11566 5451
rect 11616 5475 11660 5481
rect 11616 5455 11631 5475
rect 11651 5455 11660 5475
rect 11616 5439 11660 5455
rect 11725 5471 11774 5481
rect 11725 5451 11736 5471
rect 11756 5451 11774 5471
rect 11725 5439 11774 5451
rect 11824 5475 11868 5481
rect 11824 5455 11839 5475
rect 11859 5455 11868 5475
rect 11824 5439 11868 5455
rect 11938 5475 11982 5481
rect 11938 5455 11947 5475
rect 11967 5455 11982 5475
rect 11938 5439 11982 5455
rect 12032 5471 12081 5481
rect 12032 5451 12050 5471
rect 12070 5451 12081 5471
rect 12032 5439 12081 5451
rect 17970 5684 18019 5696
rect 17970 5664 17981 5684
rect 18001 5664 18019 5684
rect 17970 5654 18019 5664
rect 18069 5680 18113 5696
rect 18069 5660 18084 5680
rect 18104 5660 18113 5680
rect 18069 5654 18113 5660
rect 18183 5680 18227 5696
rect 18183 5660 18192 5680
rect 18212 5660 18227 5680
rect 18183 5654 18227 5660
rect 18277 5684 18326 5696
rect 18277 5664 18295 5684
rect 18315 5664 18326 5684
rect 18277 5654 18326 5664
rect 18391 5680 18435 5696
rect 18391 5660 18400 5680
rect 18420 5660 18435 5680
rect 18391 5654 18435 5660
rect 18485 5684 18534 5696
rect 18485 5664 18503 5684
rect 18523 5664 18534 5684
rect 18485 5654 18534 5664
rect 18604 5680 18648 5696
rect 18604 5660 18613 5680
rect 18633 5660 18648 5680
rect 18604 5654 18648 5660
rect 18698 5684 18747 5696
rect 18698 5664 18716 5684
rect 18736 5664 18747 5684
rect 18698 5654 18747 5664
rect 16360 5512 16409 5522
rect 16360 5492 16371 5512
rect 16391 5492 16409 5512
rect 16360 5480 16409 5492
rect 16459 5516 16503 5522
rect 16459 5496 16474 5516
rect 16494 5496 16503 5516
rect 16459 5480 16503 5496
rect 16573 5512 16622 5522
rect 16573 5492 16584 5512
rect 16604 5492 16622 5512
rect 16573 5480 16622 5492
rect 16672 5516 16716 5522
rect 16672 5496 16687 5516
rect 16707 5496 16716 5516
rect 16672 5480 16716 5496
rect 16781 5512 16830 5522
rect 16781 5492 16792 5512
rect 16812 5492 16830 5512
rect 16781 5480 16830 5492
rect 16880 5516 16924 5522
rect 16880 5496 16895 5516
rect 16915 5496 16924 5516
rect 16880 5480 16924 5496
rect 16994 5516 17038 5522
rect 16994 5496 17003 5516
rect 17023 5496 17038 5516
rect 16994 5480 17038 5496
rect 17088 5512 17137 5522
rect 17088 5492 17106 5512
rect 17126 5492 17137 5512
rect 17088 5480 17137 5492
rect 13852 5399 13901 5411
rect 13852 5379 13863 5399
rect 13883 5379 13901 5399
rect 13852 5369 13901 5379
rect 13951 5395 13995 5411
rect 13951 5375 13966 5395
rect 13986 5375 13995 5395
rect 13951 5369 13995 5375
rect 14065 5395 14109 5411
rect 14065 5375 14074 5395
rect 14094 5375 14109 5395
rect 14065 5369 14109 5375
rect 14159 5399 14208 5411
rect 14159 5379 14177 5399
rect 14197 5379 14208 5399
rect 14159 5369 14208 5379
rect 14273 5395 14317 5411
rect 14273 5375 14282 5395
rect 14302 5375 14317 5395
rect 14273 5369 14317 5375
rect 14367 5399 14416 5411
rect 14367 5379 14385 5399
rect 14405 5379 14416 5399
rect 14367 5369 14416 5379
rect 14486 5395 14530 5411
rect 14486 5375 14495 5395
rect 14515 5375 14530 5395
rect 14486 5369 14530 5375
rect 14580 5399 14629 5411
rect 14580 5379 14598 5399
rect 14618 5379 14629 5399
rect 14580 5369 14629 5379
rect 334 5156 383 5166
rect 334 5136 345 5156
rect 365 5136 383 5156
rect 334 5124 383 5136
rect 433 5160 477 5166
rect 433 5140 448 5160
rect 468 5140 477 5160
rect 433 5124 477 5140
rect 547 5156 596 5166
rect 547 5136 558 5156
rect 578 5136 596 5156
rect 547 5124 596 5136
rect 646 5160 690 5166
rect 646 5140 661 5160
rect 681 5140 690 5160
rect 646 5124 690 5140
rect 755 5156 804 5166
rect 755 5136 766 5156
rect 786 5136 804 5156
rect 755 5124 804 5136
rect 854 5160 898 5166
rect 854 5140 869 5160
rect 889 5140 898 5160
rect 854 5124 898 5140
rect 968 5160 1012 5166
rect 968 5140 977 5160
rect 997 5140 1012 5160
rect 968 5124 1012 5140
rect 1062 5156 1111 5166
rect 1062 5136 1080 5156
rect 1100 5136 1111 5156
rect 1062 5124 1111 5136
rect 5390 5197 5439 5207
rect 5390 5177 5401 5197
rect 5421 5177 5439 5197
rect 2774 5108 2823 5120
rect 2774 5088 2785 5108
rect 2805 5088 2823 5108
rect 2774 5078 2823 5088
rect 2873 5104 2917 5120
rect 2873 5084 2888 5104
rect 2908 5084 2917 5104
rect 2873 5078 2917 5084
rect 2987 5104 3031 5120
rect 2987 5084 2996 5104
rect 3016 5084 3031 5104
rect 2987 5078 3031 5084
rect 3081 5108 3130 5120
rect 3081 5088 3099 5108
rect 3119 5088 3130 5108
rect 3081 5078 3130 5088
rect 3195 5104 3239 5120
rect 3195 5084 3204 5104
rect 3224 5084 3239 5104
rect 3195 5078 3239 5084
rect 3289 5108 3338 5120
rect 3289 5088 3307 5108
rect 3327 5088 3338 5108
rect 3289 5078 3338 5088
rect 3408 5104 3452 5120
rect 3408 5084 3417 5104
rect 3437 5084 3452 5104
rect 3408 5078 3452 5084
rect 3502 5108 3551 5120
rect 3502 5088 3520 5108
rect 3540 5088 3551 5108
rect 5390 5165 5439 5177
rect 5489 5201 5533 5207
rect 5489 5181 5504 5201
rect 5524 5181 5533 5201
rect 5489 5165 5533 5181
rect 5603 5197 5652 5207
rect 5603 5177 5614 5197
rect 5634 5177 5652 5197
rect 5603 5165 5652 5177
rect 5702 5201 5746 5207
rect 5702 5181 5717 5201
rect 5737 5181 5746 5201
rect 5702 5165 5746 5181
rect 5811 5197 5860 5207
rect 5811 5177 5822 5197
rect 5842 5177 5860 5197
rect 5811 5165 5860 5177
rect 5910 5201 5954 5207
rect 5910 5181 5925 5201
rect 5945 5181 5954 5201
rect 5910 5165 5954 5181
rect 6024 5201 6068 5207
rect 6024 5181 6033 5201
rect 6053 5181 6068 5201
rect 6024 5165 6068 5181
rect 6118 5197 6167 5207
rect 6118 5177 6136 5197
rect 6156 5177 6167 5197
rect 6118 5165 6167 5177
rect 7830 5149 7879 5161
rect 3502 5078 3551 5088
rect 7830 5129 7841 5149
rect 7861 5129 7879 5149
rect 7830 5119 7879 5129
rect 7929 5145 7973 5161
rect 7929 5125 7944 5145
rect 7964 5125 7973 5145
rect 7929 5119 7973 5125
rect 8043 5145 8087 5161
rect 8043 5125 8052 5145
rect 8072 5125 8087 5145
rect 8043 5119 8087 5125
rect 8137 5149 8186 5161
rect 8137 5129 8155 5149
rect 8175 5129 8186 5149
rect 8137 5119 8186 5129
rect 8251 5145 8295 5161
rect 8251 5125 8260 5145
rect 8280 5125 8295 5145
rect 8251 5119 8295 5125
rect 8345 5149 8394 5161
rect 8345 5129 8363 5149
rect 8383 5129 8394 5149
rect 8345 5119 8394 5129
rect 8464 5145 8508 5161
rect 8464 5125 8473 5145
rect 8493 5125 8508 5145
rect 8464 5119 8508 5125
rect 8558 5149 8607 5161
rect 8558 5129 8576 5149
rect 8596 5129 8607 5149
rect 18908 5440 18957 5452
rect 18908 5420 18919 5440
rect 18939 5420 18957 5440
rect 18908 5410 18957 5420
rect 19007 5436 19051 5452
rect 19007 5416 19022 5436
rect 19042 5416 19051 5436
rect 19007 5410 19051 5416
rect 19121 5436 19165 5452
rect 19121 5416 19130 5436
rect 19150 5416 19165 5436
rect 19121 5410 19165 5416
rect 19215 5440 19264 5452
rect 19215 5420 19233 5440
rect 19253 5420 19264 5440
rect 19215 5410 19264 5420
rect 19329 5436 19373 5452
rect 19329 5416 19338 5436
rect 19358 5416 19373 5436
rect 19329 5410 19373 5416
rect 19423 5440 19472 5452
rect 19423 5420 19441 5440
rect 19461 5420 19472 5440
rect 19423 5410 19472 5420
rect 19542 5436 19586 5452
rect 19542 5416 19551 5436
rect 19571 5416 19586 5436
rect 19542 5410 19586 5416
rect 19636 5440 19685 5452
rect 19636 5420 19654 5440
rect 19674 5420 19685 5440
rect 19636 5410 19685 5420
rect 8558 5119 8607 5129
rect 10365 5161 10414 5171
rect 10365 5141 10376 5161
rect 10396 5141 10414 5161
rect 10365 5129 10414 5141
rect 10464 5165 10508 5171
rect 10464 5145 10479 5165
rect 10499 5145 10508 5165
rect 10464 5129 10508 5145
rect 10578 5161 10627 5171
rect 10578 5141 10589 5161
rect 10609 5141 10627 5161
rect 10578 5129 10627 5141
rect 10677 5165 10721 5171
rect 10677 5145 10692 5165
rect 10712 5145 10721 5165
rect 10677 5129 10721 5145
rect 10786 5161 10835 5171
rect 10786 5141 10797 5161
rect 10817 5141 10835 5161
rect 10786 5129 10835 5141
rect 10885 5165 10929 5171
rect 10885 5145 10900 5165
rect 10920 5145 10929 5165
rect 10885 5129 10929 5145
rect 10999 5165 11043 5171
rect 10999 5145 11008 5165
rect 11028 5145 11043 5165
rect 10999 5129 11043 5145
rect 11093 5161 11142 5171
rect 11093 5141 11111 5161
rect 11131 5141 11142 5161
rect 11093 5129 11142 5141
rect 15421 5202 15470 5212
rect 15421 5182 15432 5202
rect 15452 5182 15470 5202
rect 12805 5113 12854 5125
rect 12805 5093 12816 5113
rect 12836 5093 12854 5113
rect 1382 4893 1431 4903
rect 1382 4873 1393 4893
rect 1413 4873 1431 4893
rect 1382 4861 1431 4873
rect 1481 4897 1525 4903
rect 1481 4877 1496 4897
rect 1516 4877 1525 4897
rect 1481 4861 1525 4877
rect 1595 4893 1644 4903
rect 1595 4873 1606 4893
rect 1626 4873 1644 4893
rect 1595 4861 1644 4873
rect 1694 4897 1738 4903
rect 1694 4877 1709 4897
rect 1729 4877 1738 4897
rect 1694 4861 1738 4877
rect 1803 4893 1852 4903
rect 1803 4873 1814 4893
rect 1834 4873 1852 4893
rect 1803 4861 1852 4873
rect 1902 4897 1946 4903
rect 1902 4877 1917 4897
rect 1937 4877 1946 4897
rect 1902 4861 1946 4877
rect 2016 4897 2060 4903
rect 2016 4877 2025 4897
rect 2045 4877 2060 4897
rect 2016 4861 2060 4877
rect 2110 4893 2159 4903
rect 2110 4873 2128 4893
rect 2148 4873 2159 4893
rect 6438 4934 6487 4944
rect 2110 4861 2159 4873
rect 3822 4845 3871 4857
rect 3822 4825 3833 4845
rect 3853 4825 3871 4845
rect 3822 4815 3871 4825
rect 3921 4841 3965 4857
rect 3921 4821 3936 4841
rect 3956 4821 3965 4841
rect 3921 4815 3965 4821
rect 4035 4841 4079 4857
rect 4035 4821 4044 4841
rect 4064 4821 4079 4841
rect 4035 4815 4079 4821
rect 4129 4845 4178 4857
rect 4129 4825 4147 4845
rect 4167 4825 4178 4845
rect 4129 4815 4178 4825
rect 4243 4841 4287 4857
rect 4243 4821 4252 4841
rect 4272 4821 4287 4841
rect 4243 4815 4287 4821
rect 4337 4845 4386 4857
rect 4337 4825 4355 4845
rect 4375 4825 4386 4845
rect 4337 4815 4386 4825
rect 4456 4841 4500 4857
rect 4456 4821 4465 4841
rect 4485 4821 4500 4841
rect 4456 4815 4500 4821
rect 4550 4845 4599 4857
rect 6438 4914 6449 4934
rect 6469 4914 6487 4934
rect 6438 4902 6487 4914
rect 6537 4938 6581 4944
rect 6537 4918 6552 4938
rect 6572 4918 6581 4938
rect 6537 4902 6581 4918
rect 6651 4934 6700 4944
rect 6651 4914 6662 4934
rect 6682 4914 6700 4934
rect 6651 4902 6700 4914
rect 6750 4938 6794 4944
rect 6750 4918 6765 4938
rect 6785 4918 6794 4938
rect 6750 4902 6794 4918
rect 6859 4934 6908 4944
rect 6859 4914 6870 4934
rect 6890 4914 6908 4934
rect 6859 4902 6908 4914
rect 6958 4938 7002 4944
rect 6958 4918 6973 4938
rect 6993 4918 7002 4938
rect 6958 4902 7002 4918
rect 7072 4938 7116 4944
rect 7072 4918 7081 4938
rect 7101 4918 7116 4938
rect 7072 4902 7116 4918
rect 7166 4934 7215 4944
rect 12805 5083 12854 5093
rect 12904 5109 12948 5125
rect 12904 5089 12919 5109
rect 12939 5089 12948 5109
rect 12904 5083 12948 5089
rect 13018 5109 13062 5125
rect 13018 5089 13027 5109
rect 13047 5089 13062 5109
rect 13018 5083 13062 5089
rect 13112 5113 13161 5125
rect 13112 5093 13130 5113
rect 13150 5093 13161 5113
rect 13112 5083 13161 5093
rect 13226 5109 13270 5125
rect 13226 5089 13235 5109
rect 13255 5089 13270 5109
rect 13226 5083 13270 5089
rect 13320 5113 13369 5125
rect 13320 5093 13338 5113
rect 13358 5093 13369 5113
rect 13320 5083 13369 5093
rect 13439 5109 13483 5125
rect 13439 5089 13448 5109
rect 13468 5089 13483 5109
rect 13439 5083 13483 5089
rect 13533 5113 13582 5125
rect 13533 5093 13551 5113
rect 13571 5093 13582 5113
rect 15421 5170 15470 5182
rect 15520 5206 15564 5212
rect 15520 5186 15535 5206
rect 15555 5186 15564 5206
rect 15520 5170 15564 5186
rect 15634 5202 15683 5212
rect 15634 5182 15645 5202
rect 15665 5182 15683 5202
rect 15634 5170 15683 5182
rect 15733 5206 15777 5212
rect 15733 5186 15748 5206
rect 15768 5186 15777 5206
rect 15733 5170 15777 5186
rect 15842 5202 15891 5212
rect 15842 5182 15853 5202
rect 15873 5182 15891 5202
rect 15842 5170 15891 5182
rect 15941 5206 15985 5212
rect 15941 5186 15956 5206
rect 15976 5186 15985 5206
rect 15941 5170 15985 5186
rect 16055 5206 16099 5212
rect 16055 5186 16064 5206
rect 16084 5186 16099 5206
rect 16055 5170 16099 5186
rect 16149 5202 16198 5212
rect 16149 5182 16167 5202
rect 16187 5182 16198 5202
rect 16149 5170 16198 5182
rect 17861 5154 17910 5166
rect 13533 5083 13582 5093
rect 17861 5134 17872 5154
rect 17892 5134 17910 5154
rect 17861 5124 17910 5134
rect 17960 5150 18004 5166
rect 17960 5130 17975 5150
rect 17995 5130 18004 5150
rect 17960 5124 18004 5130
rect 18074 5150 18118 5166
rect 18074 5130 18083 5150
rect 18103 5130 18118 5150
rect 18074 5124 18118 5130
rect 18168 5154 18217 5166
rect 18168 5134 18186 5154
rect 18206 5134 18217 5154
rect 18168 5124 18217 5134
rect 18282 5150 18326 5166
rect 18282 5130 18291 5150
rect 18311 5130 18326 5150
rect 18282 5124 18326 5130
rect 18376 5154 18425 5166
rect 18376 5134 18394 5154
rect 18414 5134 18425 5154
rect 18376 5124 18425 5134
rect 18495 5150 18539 5166
rect 18495 5130 18504 5150
rect 18524 5130 18539 5150
rect 18495 5124 18539 5130
rect 18589 5154 18638 5166
rect 18589 5134 18607 5154
rect 18627 5134 18638 5154
rect 18589 5124 18638 5134
rect 7166 4914 7184 4934
rect 7204 4914 7215 4934
rect 7166 4902 7215 4914
rect 4550 4825 4568 4845
rect 4588 4825 4599 4845
rect 4550 4815 4599 4825
rect 8878 4886 8927 4898
rect 8878 4866 8889 4886
rect 8909 4866 8927 4886
rect 8878 4856 8927 4866
rect 8977 4882 9021 4898
rect 8977 4862 8992 4882
rect 9012 4862 9021 4882
rect 8977 4856 9021 4862
rect 9091 4882 9135 4898
rect 9091 4862 9100 4882
rect 9120 4862 9135 4882
rect 9091 4856 9135 4862
rect 9185 4886 9234 4898
rect 9185 4866 9203 4886
rect 9223 4866 9234 4886
rect 9185 4856 9234 4866
rect 9299 4882 9343 4898
rect 9299 4862 9308 4882
rect 9328 4862 9343 4882
rect 9299 4856 9343 4862
rect 9393 4886 9442 4898
rect 9393 4866 9411 4886
rect 9431 4866 9442 4886
rect 9393 4856 9442 4866
rect 9512 4882 9556 4898
rect 9512 4862 9521 4882
rect 9541 4862 9556 4882
rect 9512 4856 9556 4862
rect 9606 4886 9655 4898
rect 9606 4866 9624 4886
rect 9644 4866 9655 4886
rect 9606 4856 9655 4866
rect 11413 4898 11462 4908
rect 335 4607 384 4617
rect 335 4587 346 4607
rect 366 4587 384 4607
rect 335 4575 384 4587
rect 434 4611 478 4617
rect 434 4591 449 4611
rect 469 4591 478 4611
rect 434 4575 478 4591
rect 548 4607 597 4617
rect 548 4587 559 4607
rect 579 4587 597 4607
rect 548 4575 597 4587
rect 647 4611 691 4617
rect 647 4591 662 4611
rect 682 4591 691 4611
rect 647 4575 691 4591
rect 756 4607 805 4617
rect 756 4587 767 4607
rect 787 4587 805 4607
rect 756 4575 805 4587
rect 855 4611 899 4617
rect 855 4591 870 4611
rect 890 4591 899 4611
rect 855 4575 899 4591
rect 969 4611 1013 4617
rect 969 4591 978 4611
rect 998 4591 1013 4611
rect 969 4575 1013 4591
rect 1063 4607 1112 4617
rect 1063 4587 1081 4607
rect 1101 4587 1112 4607
rect 1063 4575 1112 4587
rect 11413 4878 11424 4898
rect 11444 4878 11462 4898
rect 11413 4866 11462 4878
rect 11512 4902 11556 4908
rect 11512 4882 11527 4902
rect 11547 4882 11556 4902
rect 11512 4866 11556 4882
rect 11626 4898 11675 4908
rect 11626 4878 11637 4898
rect 11657 4878 11675 4898
rect 11626 4866 11675 4878
rect 11725 4902 11769 4908
rect 11725 4882 11740 4902
rect 11760 4882 11769 4902
rect 11725 4866 11769 4882
rect 11834 4898 11883 4908
rect 11834 4878 11845 4898
rect 11865 4878 11883 4898
rect 11834 4866 11883 4878
rect 11933 4902 11977 4908
rect 11933 4882 11948 4902
rect 11968 4882 11977 4902
rect 11933 4866 11977 4882
rect 12047 4902 12091 4908
rect 12047 4882 12056 4902
rect 12076 4882 12091 4902
rect 12047 4866 12091 4882
rect 12141 4898 12190 4908
rect 12141 4878 12159 4898
rect 12179 4878 12190 4898
rect 16469 4939 16518 4949
rect 12141 4866 12190 4878
rect 13853 4850 13902 4862
rect 13853 4830 13864 4850
rect 13884 4830 13902 4850
rect 13853 4820 13902 4830
rect 13952 4846 13996 4862
rect 13952 4826 13967 4846
rect 13987 4826 13996 4846
rect 13952 4820 13996 4826
rect 14066 4846 14110 4862
rect 14066 4826 14075 4846
rect 14095 4826 14110 4846
rect 14066 4820 14110 4826
rect 14160 4850 14209 4862
rect 14160 4830 14178 4850
rect 14198 4830 14209 4850
rect 14160 4820 14209 4830
rect 14274 4846 14318 4862
rect 14274 4826 14283 4846
rect 14303 4826 14318 4846
rect 14274 4820 14318 4826
rect 14368 4850 14417 4862
rect 14368 4830 14386 4850
rect 14406 4830 14417 4850
rect 14368 4820 14417 4830
rect 14487 4846 14531 4862
rect 14487 4826 14496 4846
rect 14516 4826 14531 4846
rect 14487 4820 14531 4826
rect 14581 4850 14630 4862
rect 16469 4919 16480 4939
rect 16500 4919 16518 4939
rect 16469 4907 16518 4919
rect 16568 4943 16612 4949
rect 16568 4923 16583 4943
rect 16603 4923 16612 4943
rect 16568 4907 16612 4923
rect 16682 4939 16731 4949
rect 16682 4919 16693 4939
rect 16713 4919 16731 4939
rect 16682 4907 16731 4919
rect 16781 4943 16825 4949
rect 16781 4923 16796 4943
rect 16816 4923 16825 4943
rect 16781 4907 16825 4923
rect 16890 4939 16939 4949
rect 16890 4919 16901 4939
rect 16921 4919 16939 4939
rect 16890 4907 16939 4919
rect 16989 4943 17033 4949
rect 16989 4923 17004 4943
rect 17024 4923 17033 4943
rect 16989 4907 17033 4923
rect 17103 4943 17147 4949
rect 17103 4923 17112 4943
rect 17132 4923 17147 4943
rect 17103 4907 17147 4923
rect 17197 4939 17246 4949
rect 17197 4919 17215 4939
rect 17235 4919 17246 4939
rect 17197 4907 17246 4919
rect 14581 4830 14599 4850
rect 14619 4830 14630 4850
rect 14581 4820 14630 4830
rect 18909 4891 18958 4903
rect 18909 4871 18920 4891
rect 18940 4871 18958 4891
rect 18909 4861 18958 4871
rect 19008 4887 19052 4903
rect 19008 4867 19023 4887
rect 19043 4867 19052 4887
rect 19008 4861 19052 4867
rect 19122 4887 19166 4903
rect 19122 4867 19131 4887
rect 19151 4867 19166 4887
rect 19122 4861 19166 4867
rect 19216 4891 19265 4903
rect 19216 4871 19234 4891
rect 19254 4871 19265 4891
rect 19216 4861 19265 4871
rect 19330 4887 19374 4903
rect 19330 4867 19339 4887
rect 19359 4867 19374 4887
rect 19330 4861 19374 4867
rect 19424 4891 19473 4903
rect 19424 4871 19442 4891
rect 19462 4871 19473 4891
rect 19424 4861 19473 4871
rect 19543 4887 19587 4903
rect 19543 4867 19552 4887
rect 19572 4867 19587 4887
rect 19543 4861 19587 4867
rect 19637 4891 19686 4903
rect 19637 4871 19655 4891
rect 19675 4871 19686 4891
rect 19637 4861 19686 4871
rect 5391 4648 5440 4658
rect 5391 4628 5402 4648
rect 5422 4628 5440 4648
rect 5391 4616 5440 4628
rect 5490 4652 5534 4658
rect 5490 4632 5505 4652
rect 5525 4632 5534 4652
rect 5490 4616 5534 4632
rect 5604 4648 5653 4658
rect 5604 4628 5615 4648
rect 5635 4628 5653 4648
rect 5604 4616 5653 4628
rect 5703 4652 5747 4658
rect 5703 4632 5718 4652
rect 5738 4632 5747 4652
rect 5703 4616 5747 4632
rect 5812 4648 5861 4658
rect 5812 4628 5823 4648
rect 5843 4628 5861 4648
rect 5812 4616 5861 4628
rect 5911 4652 5955 4658
rect 5911 4632 5926 4652
rect 5946 4632 5955 4652
rect 5911 4616 5955 4632
rect 6025 4652 6069 4658
rect 6025 4632 6034 4652
rect 6054 4632 6069 4652
rect 6025 4616 6069 4632
rect 6119 4648 6168 4658
rect 6119 4628 6137 4648
rect 6157 4628 6168 4648
rect 6119 4616 6168 4628
rect 2883 4535 2932 4547
rect 2883 4515 2894 4535
rect 2914 4515 2932 4535
rect 2883 4505 2932 4515
rect 2982 4531 3026 4547
rect 2982 4511 2997 4531
rect 3017 4511 3026 4531
rect 2982 4505 3026 4511
rect 3096 4531 3140 4547
rect 3096 4511 3105 4531
rect 3125 4511 3140 4531
rect 3096 4505 3140 4511
rect 3190 4535 3239 4547
rect 3190 4515 3208 4535
rect 3228 4515 3239 4535
rect 3190 4505 3239 4515
rect 3304 4531 3348 4547
rect 3304 4511 3313 4531
rect 3333 4511 3348 4531
rect 3304 4505 3348 4511
rect 3398 4535 3447 4547
rect 3398 4515 3416 4535
rect 3436 4515 3447 4535
rect 3398 4505 3447 4515
rect 3517 4531 3561 4547
rect 3517 4511 3526 4531
rect 3546 4511 3561 4531
rect 3517 4505 3561 4511
rect 3611 4535 3660 4547
rect 3611 4515 3629 4535
rect 3649 4515 3660 4535
rect 3611 4505 3660 4515
rect 1273 4363 1322 4373
rect 1273 4343 1284 4363
rect 1304 4343 1322 4363
rect 1273 4331 1322 4343
rect 1372 4367 1416 4373
rect 1372 4347 1387 4367
rect 1407 4347 1416 4367
rect 1372 4331 1416 4347
rect 1486 4363 1535 4373
rect 1486 4343 1497 4363
rect 1517 4343 1535 4363
rect 1486 4331 1535 4343
rect 1585 4367 1629 4373
rect 1585 4347 1600 4367
rect 1620 4347 1629 4367
rect 1585 4331 1629 4347
rect 1694 4363 1743 4373
rect 1694 4343 1705 4363
rect 1725 4343 1743 4363
rect 1694 4331 1743 4343
rect 1793 4367 1837 4373
rect 1793 4347 1808 4367
rect 1828 4347 1837 4367
rect 1793 4331 1837 4347
rect 1907 4367 1951 4373
rect 1907 4347 1916 4367
rect 1936 4347 1951 4367
rect 1907 4331 1951 4347
rect 2001 4363 2050 4373
rect 2001 4343 2019 4363
rect 2039 4343 2050 4363
rect 2001 4331 2050 4343
rect 7939 4576 7988 4588
rect 7939 4556 7950 4576
rect 7970 4556 7988 4576
rect 7939 4546 7988 4556
rect 8038 4572 8082 4588
rect 8038 4552 8053 4572
rect 8073 4552 8082 4572
rect 8038 4546 8082 4552
rect 8152 4572 8196 4588
rect 8152 4552 8161 4572
rect 8181 4552 8196 4572
rect 8152 4546 8196 4552
rect 8246 4576 8295 4588
rect 8246 4556 8264 4576
rect 8284 4556 8295 4576
rect 8246 4546 8295 4556
rect 8360 4572 8404 4588
rect 8360 4552 8369 4572
rect 8389 4552 8404 4572
rect 8360 4546 8404 4552
rect 8454 4576 8503 4588
rect 8454 4556 8472 4576
rect 8492 4556 8503 4576
rect 8454 4546 8503 4556
rect 8573 4572 8617 4588
rect 8573 4552 8582 4572
rect 8602 4552 8617 4572
rect 8573 4546 8617 4552
rect 8667 4576 8716 4588
rect 8667 4556 8685 4576
rect 8705 4556 8716 4576
rect 8667 4546 8716 4556
rect 10366 4612 10415 4622
rect 10366 4592 10377 4612
rect 10397 4592 10415 4612
rect 10366 4580 10415 4592
rect 10465 4616 10509 4622
rect 10465 4596 10480 4616
rect 10500 4596 10509 4616
rect 10465 4580 10509 4596
rect 10579 4612 10628 4622
rect 10579 4592 10590 4612
rect 10610 4592 10628 4612
rect 10579 4580 10628 4592
rect 10678 4616 10722 4622
rect 10678 4596 10693 4616
rect 10713 4596 10722 4616
rect 10678 4580 10722 4596
rect 10787 4612 10836 4622
rect 10787 4592 10798 4612
rect 10818 4592 10836 4612
rect 10787 4580 10836 4592
rect 10886 4616 10930 4622
rect 10886 4596 10901 4616
rect 10921 4596 10930 4616
rect 10886 4580 10930 4596
rect 11000 4616 11044 4622
rect 11000 4596 11009 4616
rect 11029 4596 11044 4616
rect 11000 4580 11044 4596
rect 11094 4612 11143 4622
rect 11094 4592 11112 4612
rect 11132 4592 11143 4612
rect 11094 4580 11143 4592
rect 15422 4653 15471 4663
rect 15422 4633 15433 4653
rect 15453 4633 15471 4653
rect 15422 4621 15471 4633
rect 15521 4657 15565 4663
rect 15521 4637 15536 4657
rect 15556 4637 15565 4657
rect 15521 4621 15565 4637
rect 15635 4653 15684 4663
rect 15635 4633 15646 4653
rect 15666 4633 15684 4653
rect 15635 4621 15684 4633
rect 15734 4657 15778 4663
rect 15734 4637 15749 4657
rect 15769 4637 15778 4657
rect 15734 4621 15778 4637
rect 15843 4653 15892 4663
rect 15843 4633 15854 4653
rect 15874 4633 15892 4653
rect 15843 4621 15892 4633
rect 15942 4657 15986 4663
rect 15942 4637 15957 4657
rect 15977 4637 15986 4657
rect 15942 4621 15986 4637
rect 16056 4657 16100 4663
rect 16056 4637 16065 4657
rect 16085 4637 16100 4657
rect 16056 4621 16100 4637
rect 16150 4653 16199 4663
rect 16150 4633 16168 4653
rect 16188 4633 16199 4653
rect 16150 4621 16199 4633
rect 6329 4404 6378 4414
rect 6329 4384 6340 4404
rect 6360 4384 6378 4404
rect 6329 4372 6378 4384
rect 6428 4408 6472 4414
rect 6428 4388 6443 4408
rect 6463 4388 6472 4408
rect 6428 4372 6472 4388
rect 6542 4404 6591 4414
rect 6542 4384 6553 4404
rect 6573 4384 6591 4404
rect 6542 4372 6591 4384
rect 6641 4408 6685 4414
rect 6641 4388 6656 4408
rect 6676 4388 6685 4408
rect 6641 4372 6685 4388
rect 6750 4404 6799 4414
rect 6750 4384 6761 4404
rect 6781 4384 6799 4404
rect 6750 4372 6799 4384
rect 6849 4408 6893 4414
rect 6849 4388 6864 4408
rect 6884 4388 6893 4408
rect 6849 4372 6893 4388
rect 6963 4408 7007 4414
rect 6963 4388 6972 4408
rect 6992 4388 7007 4408
rect 6963 4372 7007 4388
rect 7057 4404 7106 4414
rect 7057 4384 7075 4404
rect 7095 4384 7106 4404
rect 7057 4372 7106 4384
rect 12914 4540 12963 4552
rect 12914 4520 12925 4540
rect 12945 4520 12963 4540
rect 12914 4510 12963 4520
rect 13013 4536 13057 4552
rect 13013 4516 13028 4536
rect 13048 4516 13057 4536
rect 13013 4510 13057 4516
rect 13127 4536 13171 4552
rect 13127 4516 13136 4536
rect 13156 4516 13171 4536
rect 13127 4510 13171 4516
rect 13221 4540 13270 4552
rect 13221 4520 13239 4540
rect 13259 4520 13270 4540
rect 13221 4510 13270 4520
rect 13335 4536 13379 4552
rect 13335 4516 13344 4536
rect 13364 4516 13379 4536
rect 13335 4510 13379 4516
rect 13429 4540 13478 4552
rect 13429 4520 13447 4540
rect 13467 4520 13478 4540
rect 13429 4510 13478 4520
rect 13548 4536 13592 4552
rect 13548 4516 13557 4536
rect 13577 4516 13592 4536
rect 13548 4510 13592 4516
rect 13642 4540 13691 4552
rect 13642 4520 13660 4540
rect 13680 4520 13691 4540
rect 13642 4510 13691 4520
rect 3821 4291 3870 4303
rect 3821 4271 3832 4291
rect 3852 4271 3870 4291
rect 3821 4261 3870 4271
rect 3920 4287 3964 4303
rect 3920 4267 3935 4287
rect 3955 4267 3964 4287
rect 3920 4261 3964 4267
rect 4034 4287 4078 4303
rect 4034 4267 4043 4287
rect 4063 4267 4078 4287
rect 4034 4261 4078 4267
rect 4128 4291 4177 4303
rect 4128 4271 4146 4291
rect 4166 4271 4177 4291
rect 4128 4261 4177 4271
rect 4242 4287 4286 4303
rect 4242 4267 4251 4287
rect 4271 4267 4286 4287
rect 4242 4261 4286 4267
rect 4336 4291 4385 4303
rect 4336 4271 4354 4291
rect 4374 4271 4385 4291
rect 4336 4261 4385 4271
rect 4455 4287 4499 4303
rect 4455 4267 4464 4287
rect 4484 4267 4499 4287
rect 4455 4261 4499 4267
rect 4549 4291 4598 4303
rect 4549 4271 4567 4291
rect 4587 4271 4598 4291
rect 4549 4261 4598 4271
rect 8877 4332 8926 4344
rect 8877 4312 8888 4332
rect 8908 4312 8926 4332
rect 8877 4302 8926 4312
rect 8976 4328 9020 4344
rect 8976 4308 8991 4328
rect 9011 4308 9020 4328
rect 8976 4302 9020 4308
rect 9090 4328 9134 4344
rect 9090 4308 9099 4328
rect 9119 4308 9134 4328
rect 9090 4302 9134 4308
rect 9184 4332 9233 4344
rect 9184 4312 9202 4332
rect 9222 4312 9233 4332
rect 9184 4302 9233 4312
rect 9298 4328 9342 4344
rect 9298 4308 9307 4328
rect 9327 4308 9342 4328
rect 9298 4302 9342 4308
rect 9392 4332 9441 4344
rect 9392 4312 9410 4332
rect 9430 4312 9441 4332
rect 9392 4302 9441 4312
rect 9511 4328 9555 4344
rect 9511 4308 9520 4328
rect 9540 4308 9555 4328
rect 9511 4302 9555 4308
rect 9605 4332 9654 4344
rect 9605 4312 9623 4332
rect 9643 4312 9654 4332
rect 9605 4302 9654 4312
rect 11304 4368 11353 4378
rect 11304 4348 11315 4368
rect 11335 4348 11353 4368
rect 11304 4336 11353 4348
rect 11403 4372 11447 4378
rect 11403 4352 11418 4372
rect 11438 4352 11447 4372
rect 11403 4336 11447 4352
rect 11517 4368 11566 4378
rect 11517 4348 11528 4368
rect 11548 4348 11566 4368
rect 11517 4336 11566 4348
rect 11616 4372 11660 4378
rect 11616 4352 11631 4372
rect 11651 4352 11660 4372
rect 11616 4336 11660 4352
rect 11725 4368 11774 4378
rect 11725 4348 11736 4368
rect 11756 4348 11774 4368
rect 11725 4336 11774 4348
rect 11824 4372 11868 4378
rect 11824 4352 11839 4372
rect 11859 4352 11868 4372
rect 11824 4336 11868 4352
rect 11938 4372 11982 4378
rect 11938 4352 11947 4372
rect 11967 4352 11982 4372
rect 11938 4336 11982 4352
rect 12032 4368 12081 4378
rect 12032 4348 12050 4368
rect 12070 4348 12081 4368
rect 12032 4336 12081 4348
rect 17970 4581 18019 4593
rect 17970 4561 17981 4581
rect 18001 4561 18019 4581
rect 17970 4551 18019 4561
rect 18069 4577 18113 4593
rect 18069 4557 18084 4577
rect 18104 4557 18113 4577
rect 18069 4551 18113 4557
rect 18183 4577 18227 4593
rect 18183 4557 18192 4577
rect 18212 4557 18227 4577
rect 18183 4551 18227 4557
rect 18277 4581 18326 4593
rect 18277 4561 18295 4581
rect 18315 4561 18326 4581
rect 18277 4551 18326 4561
rect 18391 4577 18435 4593
rect 18391 4557 18400 4577
rect 18420 4557 18435 4577
rect 18391 4551 18435 4557
rect 18485 4581 18534 4593
rect 18485 4561 18503 4581
rect 18523 4561 18534 4581
rect 18485 4551 18534 4561
rect 18604 4577 18648 4593
rect 18604 4557 18613 4577
rect 18633 4557 18648 4577
rect 18604 4551 18648 4557
rect 18698 4581 18747 4593
rect 18698 4561 18716 4581
rect 18736 4561 18747 4581
rect 18698 4551 18747 4561
rect 16360 4409 16409 4419
rect 16360 4389 16371 4409
rect 16391 4389 16409 4409
rect 16360 4377 16409 4389
rect 16459 4413 16503 4419
rect 16459 4393 16474 4413
rect 16494 4393 16503 4413
rect 16459 4377 16503 4393
rect 16573 4409 16622 4419
rect 16573 4389 16584 4409
rect 16604 4389 16622 4409
rect 16573 4377 16622 4389
rect 16672 4413 16716 4419
rect 16672 4393 16687 4413
rect 16707 4393 16716 4413
rect 16672 4377 16716 4393
rect 16781 4409 16830 4419
rect 16781 4389 16792 4409
rect 16812 4389 16830 4409
rect 16781 4377 16830 4389
rect 16880 4413 16924 4419
rect 16880 4393 16895 4413
rect 16915 4393 16924 4413
rect 16880 4377 16924 4393
rect 16994 4413 17038 4419
rect 16994 4393 17003 4413
rect 17023 4393 17038 4413
rect 16994 4377 17038 4393
rect 17088 4409 17137 4419
rect 17088 4389 17106 4409
rect 17126 4389 17137 4409
rect 17088 4377 17137 4389
rect 13852 4296 13901 4308
rect 13852 4276 13863 4296
rect 13883 4276 13901 4296
rect 13852 4266 13901 4276
rect 13951 4292 13995 4308
rect 13951 4272 13966 4292
rect 13986 4272 13995 4292
rect 13951 4266 13995 4272
rect 14065 4292 14109 4308
rect 14065 4272 14074 4292
rect 14094 4272 14109 4292
rect 14065 4266 14109 4272
rect 14159 4296 14208 4308
rect 14159 4276 14177 4296
rect 14197 4276 14208 4296
rect 14159 4266 14208 4276
rect 14273 4292 14317 4308
rect 14273 4272 14282 4292
rect 14302 4272 14317 4292
rect 14273 4266 14317 4272
rect 14367 4296 14416 4308
rect 14367 4276 14385 4296
rect 14405 4276 14416 4296
rect 14367 4266 14416 4276
rect 14486 4292 14530 4308
rect 14486 4272 14495 4292
rect 14515 4272 14530 4292
rect 14486 4266 14530 4272
rect 14580 4296 14629 4308
rect 14580 4276 14598 4296
rect 14618 4276 14629 4296
rect 14580 4266 14629 4276
rect 5390 4094 5439 4104
rect 5390 4074 5401 4094
rect 5421 4074 5439 4094
rect 334 4053 383 4063
rect 334 4033 345 4053
rect 365 4033 383 4053
rect 334 4021 383 4033
rect 433 4057 477 4063
rect 433 4037 448 4057
rect 468 4037 477 4057
rect 433 4021 477 4037
rect 547 4053 596 4063
rect 547 4033 558 4053
rect 578 4033 596 4053
rect 547 4021 596 4033
rect 646 4057 690 4063
rect 646 4037 661 4057
rect 681 4037 690 4057
rect 646 4021 690 4037
rect 755 4053 804 4063
rect 755 4033 766 4053
rect 786 4033 804 4053
rect 755 4021 804 4033
rect 854 4057 898 4063
rect 854 4037 869 4057
rect 889 4037 898 4057
rect 854 4021 898 4037
rect 968 4057 1012 4063
rect 968 4037 977 4057
rect 997 4037 1012 4057
rect 968 4021 1012 4037
rect 1062 4053 1111 4063
rect 1062 4033 1080 4053
rect 1100 4033 1111 4053
rect 1062 4021 1111 4033
rect 2743 4024 2792 4036
rect 2743 4004 2754 4024
rect 2774 4004 2792 4024
rect 2743 3994 2792 4004
rect 2842 4020 2886 4036
rect 2842 4000 2857 4020
rect 2877 4000 2886 4020
rect 2842 3994 2886 4000
rect 2956 4020 3000 4036
rect 2956 4000 2965 4020
rect 2985 4000 3000 4020
rect 2956 3994 3000 4000
rect 3050 4024 3099 4036
rect 3050 4004 3068 4024
rect 3088 4004 3099 4024
rect 3050 3994 3099 4004
rect 3164 4020 3208 4036
rect 3164 4000 3173 4020
rect 3193 4000 3208 4020
rect 3164 3994 3208 4000
rect 3258 4024 3307 4036
rect 3258 4004 3276 4024
rect 3296 4004 3307 4024
rect 3258 3994 3307 4004
rect 3377 4020 3421 4036
rect 3377 4000 3386 4020
rect 3406 4000 3421 4020
rect 3377 3994 3421 4000
rect 3471 4024 3520 4036
rect 3471 4004 3489 4024
rect 3509 4004 3520 4024
rect 3471 3994 3520 4004
rect 5390 4062 5439 4074
rect 5489 4098 5533 4104
rect 5489 4078 5504 4098
rect 5524 4078 5533 4098
rect 5489 4062 5533 4078
rect 5603 4094 5652 4104
rect 5603 4074 5614 4094
rect 5634 4074 5652 4094
rect 5603 4062 5652 4074
rect 5702 4098 5746 4104
rect 5702 4078 5717 4098
rect 5737 4078 5746 4098
rect 5702 4062 5746 4078
rect 5811 4094 5860 4104
rect 5811 4074 5822 4094
rect 5842 4074 5860 4094
rect 5811 4062 5860 4074
rect 5910 4098 5954 4104
rect 5910 4078 5925 4098
rect 5945 4078 5954 4098
rect 5910 4062 5954 4078
rect 6024 4098 6068 4104
rect 6024 4078 6033 4098
rect 6053 4078 6068 4098
rect 6024 4062 6068 4078
rect 6118 4094 6167 4104
rect 6118 4074 6136 4094
rect 6156 4074 6167 4094
rect 6118 4062 6167 4074
rect 7799 4065 7848 4077
rect 7799 4045 7810 4065
rect 7830 4045 7848 4065
rect 7799 4035 7848 4045
rect 7898 4061 7942 4077
rect 7898 4041 7913 4061
rect 7933 4041 7942 4061
rect 7898 4035 7942 4041
rect 8012 4061 8056 4077
rect 8012 4041 8021 4061
rect 8041 4041 8056 4061
rect 8012 4035 8056 4041
rect 8106 4065 8155 4077
rect 8106 4045 8124 4065
rect 8144 4045 8155 4065
rect 8106 4035 8155 4045
rect 8220 4061 8264 4077
rect 8220 4041 8229 4061
rect 8249 4041 8264 4061
rect 8220 4035 8264 4041
rect 8314 4065 8363 4077
rect 8314 4045 8332 4065
rect 8352 4045 8363 4065
rect 8314 4035 8363 4045
rect 8433 4061 8477 4077
rect 8433 4041 8442 4061
rect 8462 4041 8477 4061
rect 8433 4035 8477 4041
rect 8527 4065 8576 4077
rect 8527 4045 8545 4065
rect 8565 4045 8576 4065
rect 8527 4035 8576 4045
rect 18908 4337 18957 4349
rect 18908 4317 18919 4337
rect 18939 4317 18957 4337
rect 18908 4307 18957 4317
rect 19007 4333 19051 4349
rect 19007 4313 19022 4333
rect 19042 4313 19051 4333
rect 19007 4307 19051 4313
rect 19121 4333 19165 4349
rect 19121 4313 19130 4333
rect 19150 4313 19165 4333
rect 19121 4307 19165 4313
rect 19215 4337 19264 4349
rect 19215 4317 19233 4337
rect 19253 4317 19264 4337
rect 19215 4307 19264 4317
rect 19329 4333 19373 4349
rect 19329 4313 19338 4333
rect 19358 4313 19373 4333
rect 19329 4307 19373 4313
rect 19423 4337 19472 4349
rect 19423 4317 19441 4337
rect 19461 4317 19472 4337
rect 19423 4307 19472 4317
rect 19542 4333 19586 4349
rect 19542 4313 19551 4333
rect 19571 4313 19586 4333
rect 19542 4307 19586 4313
rect 19636 4337 19685 4349
rect 19636 4317 19654 4337
rect 19674 4317 19685 4337
rect 19636 4307 19685 4317
rect 15421 4099 15470 4109
rect 15421 4079 15432 4099
rect 15452 4079 15470 4099
rect 10365 4058 10414 4068
rect 10365 4038 10376 4058
rect 10396 4038 10414 4058
rect 10365 4026 10414 4038
rect 10464 4062 10508 4068
rect 10464 4042 10479 4062
rect 10499 4042 10508 4062
rect 10464 4026 10508 4042
rect 10578 4058 10627 4068
rect 10578 4038 10589 4058
rect 10609 4038 10627 4058
rect 10578 4026 10627 4038
rect 10677 4062 10721 4068
rect 10677 4042 10692 4062
rect 10712 4042 10721 4062
rect 10677 4026 10721 4042
rect 10786 4058 10835 4068
rect 10786 4038 10797 4058
rect 10817 4038 10835 4058
rect 10786 4026 10835 4038
rect 10885 4062 10929 4068
rect 10885 4042 10900 4062
rect 10920 4042 10929 4062
rect 10885 4026 10929 4042
rect 10999 4062 11043 4068
rect 10999 4042 11008 4062
rect 11028 4042 11043 4062
rect 10999 4026 11043 4042
rect 11093 4058 11142 4068
rect 11093 4038 11111 4058
rect 11131 4038 11142 4058
rect 11093 4026 11142 4038
rect 12774 4029 12823 4041
rect 12774 4009 12785 4029
rect 12805 4009 12823 4029
rect 12774 3999 12823 4009
rect 12873 4025 12917 4041
rect 12873 4005 12888 4025
rect 12908 4005 12917 4025
rect 12873 3999 12917 4005
rect 12987 4025 13031 4041
rect 12987 4005 12996 4025
rect 13016 4005 13031 4025
rect 12987 3999 13031 4005
rect 13081 4029 13130 4041
rect 13081 4009 13099 4029
rect 13119 4009 13130 4029
rect 13081 3999 13130 4009
rect 13195 4025 13239 4041
rect 13195 4005 13204 4025
rect 13224 4005 13239 4025
rect 13195 3999 13239 4005
rect 13289 4029 13338 4041
rect 13289 4009 13307 4029
rect 13327 4009 13338 4029
rect 13289 3999 13338 4009
rect 13408 4025 13452 4041
rect 13408 4005 13417 4025
rect 13437 4005 13452 4025
rect 13408 3999 13452 4005
rect 13502 4029 13551 4041
rect 13502 4009 13520 4029
rect 13540 4009 13551 4029
rect 13502 3999 13551 4009
rect 15421 4067 15470 4079
rect 15520 4103 15564 4109
rect 15520 4083 15535 4103
rect 15555 4083 15564 4103
rect 15520 4067 15564 4083
rect 15634 4099 15683 4109
rect 15634 4079 15645 4099
rect 15665 4079 15683 4099
rect 15634 4067 15683 4079
rect 15733 4103 15777 4109
rect 15733 4083 15748 4103
rect 15768 4083 15777 4103
rect 15733 4067 15777 4083
rect 15842 4099 15891 4109
rect 15842 4079 15853 4099
rect 15873 4079 15891 4099
rect 15842 4067 15891 4079
rect 15941 4103 15985 4109
rect 15941 4083 15956 4103
rect 15976 4083 15985 4103
rect 15941 4067 15985 4083
rect 16055 4103 16099 4109
rect 16055 4083 16064 4103
rect 16084 4083 16099 4103
rect 16055 4067 16099 4083
rect 16149 4099 16198 4109
rect 16149 4079 16167 4099
rect 16187 4079 16198 4099
rect 16149 4067 16198 4079
rect 17830 4070 17879 4082
rect 17830 4050 17841 4070
rect 17861 4050 17879 4070
rect 17830 4040 17879 4050
rect 17929 4066 17973 4082
rect 17929 4046 17944 4066
rect 17964 4046 17973 4066
rect 17929 4040 17973 4046
rect 18043 4066 18087 4082
rect 18043 4046 18052 4066
rect 18072 4046 18087 4066
rect 18043 4040 18087 4046
rect 18137 4070 18186 4082
rect 18137 4050 18155 4070
rect 18175 4050 18186 4070
rect 18137 4040 18186 4050
rect 18251 4066 18295 4082
rect 18251 4046 18260 4066
rect 18280 4046 18295 4066
rect 18251 4040 18295 4046
rect 18345 4070 18394 4082
rect 18345 4050 18363 4070
rect 18383 4050 18394 4070
rect 18345 4040 18394 4050
rect 18464 4066 18508 4082
rect 18464 4046 18473 4066
rect 18493 4046 18508 4066
rect 18464 4040 18508 4046
rect 18558 4070 18607 4082
rect 18558 4050 18576 4070
rect 18596 4050 18607 4070
rect 18558 4040 18607 4050
rect 1414 3771 1463 3781
rect 1414 3751 1425 3771
rect 1445 3751 1463 3771
rect 1414 3739 1463 3751
rect 1513 3775 1557 3781
rect 1513 3755 1528 3775
rect 1548 3755 1557 3775
rect 1513 3739 1557 3755
rect 1627 3771 1676 3781
rect 1627 3751 1638 3771
rect 1658 3751 1676 3771
rect 1627 3739 1676 3751
rect 1726 3775 1770 3781
rect 1726 3755 1741 3775
rect 1761 3755 1770 3775
rect 1726 3739 1770 3755
rect 1835 3771 1884 3781
rect 1835 3751 1846 3771
rect 1866 3751 1884 3771
rect 1835 3739 1884 3751
rect 1934 3775 1978 3781
rect 1934 3755 1949 3775
rect 1969 3755 1978 3775
rect 1934 3739 1978 3755
rect 2048 3775 2092 3781
rect 2048 3755 2057 3775
rect 2077 3755 2092 3775
rect 2048 3739 2092 3755
rect 2142 3771 2191 3781
rect 2142 3751 2160 3771
rect 2180 3751 2191 3771
rect 2142 3739 2191 3751
rect 3823 3742 3872 3754
rect 3823 3722 3834 3742
rect 3854 3722 3872 3742
rect 3823 3712 3872 3722
rect 3922 3738 3966 3754
rect 3922 3718 3937 3738
rect 3957 3718 3966 3738
rect 3922 3712 3966 3718
rect 4036 3738 4080 3754
rect 4036 3718 4045 3738
rect 4065 3718 4080 3738
rect 4036 3712 4080 3718
rect 4130 3742 4179 3754
rect 4130 3722 4148 3742
rect 4168 3722 4179 3742
rect 4130 3712 4179 3722
rect 4244 3738 4288 3754
rect 4244 3718 4253 3738
rect 4273 3718 4288 3738
rect 4244 3712 4288 3718
rect 4338 3742 4387 3754
rect 4338 3722 4356 3742
rect 4376 3722 4387 3742
rect 4338 3712 4387 3722
rect 4457 3738 4501 3754
rect 4457 3718 4466 3738
rect 4486 3718 4501 3738
rect 4457 3712 4501 3718
rect 4551 3742 4600 3754
rect 6470 3812 6519 3822
rect 6470 3792 6481 3812
rect 6501 3792 6519 3812
rect 6470 3780 6519 3792
rect 6569 3816 6613 3822
rect 6569 3796 6584 3816
rect 6604 3796 6613 3816
rect 6569 3780 6613 3796
rect 6683 3812 6732 3822
rect 6683 3792 6694 3812
rect 6714 3792 6732 3812
rect 6683 3780 6732 3792
rect 6782 3816 6826 3822
rect 6782 3796 6797 3816
rect 6817 3796 6826 3816
rect 6782 3780 6826 3796
rect 6891 3812 6940 3822
rect 6891 3792 6902 3812
rect 6922 3792 6940 3812
rect 6891 3780 6940 3792
rect 6990 3816 7034 3822
rect 6990 3796 7005 3816
rect 7025 3796 7034 3816
rect 6990 3780 7034 3796
rect 7104 3816 7148 3822
rect 7104 3796 7113 3816
rect 7133 3796 7148 3816
rect 7104 3780 7148 3796
rect 7198 3812 7247 3822
rect 7198 3792 7216 3812
rect 7236 3792 7247 3812
rect 7198 3780 7247 3792
rect 8879 3783 8928 3795
rect 8879 3763 8890 3783
rect 8910 3763 8928 3783
rect 8879 3753 8928 3763
rect 8978 3779 9022 3795
rect 8978 3759 8993 3779
rect 9013 3759 9022 3779
rect 8978 3753 9022 3759
rect 9092 3779 9136 3795
rect 9092 3759 9101 3779
rect 9121 3759 9136 3779
rect 9092 3753 9136 3759
rect 9186 3783 9235 3795
rect 9186 3763 9204 3783
rect 9224 3763 9235 3783
rect 9186 3753 9235 3763
rect 9300 3779 9344 3795
rect 9300 3759 9309 3779
rect 9329 3759 9344 3779
rect 9300 3753 9344 3759
rect 9394 3783 9443 3795
rect 9394 3763 9412 3783
rect 9432 3763 9443 3783
rect 9394 3753 9443 3763
rect 9513 3779 9557 3795
rect 9513 3759 9522 3779
rect 9542 3759 9557 3779
rect 9513 3753 9557 3759
rect 9607 3783 9656 3795
rect 9607 3763 9625 3783
rect 9645 3763 9656 3783
rect 9607 3753 9656 3763
rect 4551 3722 4569 3742
rect 4589 3722 4600 3742
rect 4551 3712 4600 3722
rect 336 3504 385 3514
rect 336 3484 347 3504
rect 367 3484 385 3504
rect 336 3472 385 3484
rect 435 3508 479 3514
rect 435 3488 450 3508
rect 470 3488 479 3508
rect 435 3472 479 3488
rect 549 3504 598 3514
rect 549 3484 560 3504
rect 580 3484 598 3504
rect 549 3472 598 3484
rect 648 3508 692 3514
rect 648 3488 663 3508
rect 683 3488 692 3508
rect 648 3472 692 3488
rect 757 3504 806 3514
rect 757 3484 768 3504
rect 788 3484 806 3504
rect 757 3472 806 3484
rect 856 3508 900 3514
rect 856 3488 871 3508
rect 891 3488 900 3508
rect 856 3472 900 3488
rect 970 3508 1014 3514
rect 970 3488 979 3508
rect 999 3488 1014 3508
rect 970 3472 1014 3488
rect 1064 3504 1113 3514
rect 1064 3484 1082 3504
rect 1102 3484 1113 3504
rect 1064 3472 1113 3484
rect 11445 3776 11494 3786
rect 11445 3756 11456 3776
rect 11476 3756 11494 3776
rect 11445 3744 11494 3756
rect 11544 3780 11588 3786
rect 11544 3760 11559 3780
rect 11579 3760 11588 3780
rect 11544 3744 11588 3760
rect 11658 3776 11707 3786
rect 11658 3756 11669 3776
rect 11689 3756 11707 3776
rect 11658 3744 11707 3756
rect 11757 3780 11801 3786
rect 11757 3760 11772 3780
rect 11792 3760 11801 3780
rect 11757 3744 11801 3760
rect 11866 3776 11915 3786
rect 11866 3756 11877 3776
rect 11897 3756 11915 3776
rect 11866 3744 11915 3756
rect 11965 3780 12009 3786
rect 11965 3760 11980 3780
rect 12000 3760 12009 3780
rect 11965 3744 12009 3760
rect 12079 3780 12123 3786
rect 12079 3760 12088 3780
rect 12108 3760 12123 3780
rect 12079 3744 12123 3760
rect 12173 3776 12222 3786
rect 12173 3756 12191 3776
rect 12211 3756 12222 3776
rect 12173 3744 12222 3756
rect 13854 3747 13903 3759
rect 13854 3727 13865 3747
rect 13885 3727 13903 3747
rect 13854 3717 13903 3727
rect 13953 3743 13997 3759
rect 13953 3723 13968 3743
rect 13988 3723 13997 3743
rect 13953 3717 13997 3723
rect 14067 3743 14111 3759
rect 14067 3723 14076 3743
rect 14096 3723 14111 3743
rect 14067 3717 14111 3723
rect 14161 3747 14210 3759
rect 14161 3727 14179 3747
rect 14199 3727 14210 3747
rect 14161 3717 14210 3727
rect 14275 3743 14319 3759
rect 14275 3723 14284 3743
rect 14304 3723 14319 3743
rect 14275 3717 14319 3723
rect 14369 3747 14418 3759
rect 14369 3727 14387 3747
rect 14407 3727 14418 3747
rect 14369 3717 14418 3727
rect 14488 3743 14532 3759
rect 14488 3723 14497 3743
rect 14517 3723 14532 3743
rect 14488 3717 14532 3723
rect 14582 3747 14631 3759
rect 16501 3817 16550 3827
rect 16501 3797 16512 3817
rect 16532 3797 16550 3817
rect 16501 3785 16550 3797
rect 16600 3821 16644 3827
rect 16600 3801 16615 3821
rect 16635 3801 16644 3821
rect 16600 3785 16644 3801
rect 16714 3817 16763 3827
rect 16714 3797 16725 3817
rect 16745 3797 16763 3817
rect 16714 3785 16763 3797
rect 16813 3821 16857 3827
rect 16813 3801 16828 3821
rect 16848 3801 16857 3821
rect 16813 3785 16857 3801
rect 16922 3817 16971 3827
rect 16922 3797 16933 3817
rect 16953 3797 16971 3817
rect 16922 3785 16971 3797
rect 17021 3821 17065 3827
rect 17021 3801 17036 3821
rect 17056 3801 17065 3821
rect 17021 3785 17065 3801
rect 17135 3821 17179 3827
rect 17135 3801 17144 3821
rect 17164 3801 17179 3821
rect 17135 3785 17179 3801
rect 17229 3817 17278 3827
rect 17229 3797 17247 3817
rect 17267 3797 17278 3817
rect 17229 3785 17278 3797
rect 18910 3788 18959 3800
rect 18910 3768 18921 3788
rect 18941 3768 18959 3788
rect 18910 3758 18959 3768
rect 19009 3784 19053 3800
rect 19009 3764 19024 3784
rect 19044 3764 19053 3784
rect 19009 3758 19053 3764
rect 19123 3784 19167 3800
rect 19123 3764 19132 3784
rect 19152 3764 19167 3784
rect 19123 3758 19167 3764
rect 19217 3788 19266 3800
rect 19217 3768 19235 3788
rect 19255 3768 19266 3788
rect 19217 3758 19266 3768
rect 19331 3784 19375 3800
rect 19331 3764 19340 3784
rect 19360 3764 19375 3784
rect 19331 3758 19375 3764
rect 19425 3788 19474 3800
rect 19425 3768 19443 3788
rect 19463 3768 19474 3788
rect 19425 3758 19474 3768
rect 19544 3784 19588 3800
rect 19544 3764 19553 3784
rect 19573 3764 19588 3784
rect 19544 3758 19588 3764
rect 19638 3788 19687 3800
rect 19638 3768 19656 3788
rect 19676 3768 19687 3788
rect 19638 3758 19687 3768
rect 14582 3727 14600 3747
rect 14620 3727 14631 3747
rect 14582 3717 14631 3727
rect 5392 3545 5441 3555
rect 5392 3525 5403 3545
rect 5423 3525 5441 3545
rect 5392 3513 5441 3525
rect 5491 3549 5535 3555
rect 5491 3529 5506 3549
rect 5526 3529 5535 3549
rect 5491 3513 5535 3529
rect 5605 3545 5654 3555
rect 5605 3525 5616 3545
rect 5636 3525 5654 3545
rect 5605 3513 5654 3525
rect 5704 3549 5748 3555
rect 5704 3529 5719 3549
rect 5739 3529 5748 3549
rect 5704 3513 5748 3529
rect 5813 3545 5862 3555
rect 5813 3525 5824 3545
rect 5844 3525 5862 3545
rect 5813 3513 5862 3525
rect 5912 3549 5956 3555
rect 5912 3529 5927 3549
rect 5947 3529 5956 3549
rect 5912 3513 5956 3529
rect 6026 3549 6070 3555
rect 6026 3529 6035 3549
rect 6055 3529 6070 3549
rect 6026 3513 6070 3529
rect 6120 3545 6169 3555
rect 6120 3525 6138 3545
rect 6158 3525 6169 3545
rect 6120 3513 6169 3525
rect 2884 3432 2933 3444
rect 2884 3412 2895 3432
rect 2915 3412 2933 3432
rect 2884 3402 2933 3412
rect 2983 3428 3027 3444
rect 2983 3408 2998 3428
rect 3018 3408 3027 3428
rect 2983 3402 3027 3408
rect 3097 3428 3141 3444
rect 3097 3408 3106 3428
rect 3126 3408 3141 3428
rect 3097 3402 3141 3408
rect 3191 3432 3240 3444
rect 3191 3412 3209 3432
rect 3229 3412 3240 3432
rect 3191 3402 3240 3412
rect 3305 3428 3349 3444
rect 3305 3408 3314 3428
rect 3334 3408 3349 3428
rect 3305 3402 3349 3408
rect 3399 3432 3448 3444
rect 3399 3412 3417 3432
rect 3437 3412 3448 3432
rect 3399 3402 3448 3412
rect 3518 3428 3562 3444
rect 3518 3408 3527 3428
rect 3547 3408 3562 3428
rect 3518 3402 3562 3408
rect 3612 3432 3661 3444
rect 3612 3412 3630 3432
rect 3650 3412 3661 3432
rect 3612 3402 3661 3412
rect 1274 3260 1323 3270
rect 1274 3240 1285 3260
rect 1305 3240 1323 3260
rect 1274 3228 1323 3240
rect 1373 3264 1417 3270
rect 1373 3244 1388 3264
rect 1408 3244 1417 3264
rect 1373 3228 1417 3244
rect 1487 3260 1536 3270
rect 1487 3240 1498 3260
rect 1518 3240 1536 3260
rect 1487 3228 1536 3240
rect 1586 3264 1630 3270
rect 1586 3244 1601 3264
rect 1621 3244 1630 3264
rect 1586 3228 1630 3244
rect 1695 3260 1744 3270
rect 1695 3240 1706 3260
rect 1726 3240 1744 3260
rect 1695 3228 1744 3240
rect 1794 3264 1838 3270
rect 1794 3244 1809 3264
rect 1829 3244 1838 3264
rect 1794 3228 1838 3244
rect 1908 3264 1952 3270
rect 1908 3244 1917 3264
rect 1937 3244 1952 3264
rect 1908 3228 1952 3244
rect 2002 3260 2051 3270
rect 2002 3240 2020 3260
rect 2040 3240 2051 3260
rect 2002 3228 2051 3240
rect 7940 3473 7989 3485
rect 7940 3453 7951 3473
rect 7971 3453 7989 3473
rect 7940 3443 7989 3453
rect 8039 3469 8083 3485
rect 8039 3449 8054 3469
rect 8074 3449 8083 3469
rect 8039 3443 8083 3449
rect 8153 3469 8197 3485
rect 8153 3449 8162 3469
rect 8182 3449 8197 3469
rect 8153 3443 8197 3449
rect 8247 3473 8296 3485
rect 8247 3453 8265 3473
rect 8285 3453 8296 3473
rect 8247 3443 8296 3453
rect 8361 3469 8405 3485
rect 8361 3449 8370 3469
rect 8390 3449 8405 3469
rect 8361 3443 8405 3449
rect 8455 3473 8504 3485
rect 8455 3453 8473 3473
rect 8493 3453 8504 3473
rect 8455 3443 8504 3453
rect 8574 3469 8618 3485
rect 8574 3449 8583 3469
rect 8603 3449 8618 3469
rect 8574 3443 8618 3449
rect 8668 3473 8717 3485
rect 8668 3453 8686 3473
rect 8706 3453 8717 3473
rect 8668 3443 8717 3453
rect 10367 3509 10416 3519
rect 10367 3489 10378 3509
rect 10398 3489 10416 3509
rect 10367 3477 10416 3489
rect 10466 3513 10510 3519
rect 10466 3493 10481 3513
rect 10501 3493 10510 3513
rect 10466 3477 10510 3493
rect 10580 3509 10629 3519
rect 10580 3489 10591 3509
rect 10611 3489 10629 3509
rect 10580 3477 10629 3489
rect 10679 3513 10723 3519
rect 10679 3493 10694 3513
rect 10714 3493 10723 3513
rect 10679 3477 10723 3493
rect 10788 3509 10837 3519
rect 10788 3489 10799 3509
rect 10819 3489 10837 3509
rect 10788 3477 10837 3489
rect 10887 3513 10931 3519
rect 10887 3493 10902 3513
rect 10922 3493 10931 3513
rect 10887 3477 10931 3493
rect 11001 3513 11045 3519
rect 11001 3493 11010 3513
rect 11030 3493 11045 3513
rect 11001 3477 11045 3493
rect 11095 3509 11144 3519
rect 11095 3489 11113 3509
rect 11133 3489 11144 3509
rect 11095 3477 11144 3489
rect 15423 3550 15472 3560
rect 15423 3530 15434 3550
rect 15454 3530 15472 3550
rect 15423 3518 15472 3530
rect 15522 3554 15566 3560
rect 15522 3534 15537 3554
rect 15557 3534 15566 3554
rect 15522 3518 15566 3534
rect 15636 3550 15685 3560
rect 15636 3530 15647 3550
rect 15667 3530 15685 3550
rect 15636 3518 15685 3530
rect 15735 3554 15779 3560
rect 15735 3534 15750 3554
rect 15770 3534 15779 3554
rect 15735 3518 15779 3534
rect 15844 3550 15893 3560
rect 15844 3530 15855 3550
rect 15875 3530 15893 3550
rect 15844 3518 15893 3530
rect 15943 3554 15987 3560
rect 15943 3534 15958 3554
rect 15978 3534 15987 3554
rect 15943 3518 15987 3534
rect 16057 3554 16101 3560
rect 16057 3534 16066 3554
rect 16086 3534 16101 3554
rect 16057 3518 16101 3534
rect 16151 3550 16200 3560
rect 16151 3530 16169 3550
rect 16189 3530 16200 3550
rect 16151 3518 16200 3530
rect 6330 3301 6379 3311
rect 6330 3281 6341 3301
rect 6361 3281 6379 3301
rect 6330 3269 6379 3281
rect 6429 3305 6473 3311
rect 6429 3285 6444 3305
rect 6464 3285 6473 3305
rect 6429 3269 6473 3285
rect 6543 3301 6592 3311
rect 6543 3281 6554 3301
rect 6574 3281 6592 3301
rect 6543 3269 6592 3281
rect 6642 3305 6686 3311
rect 6642 3285 6657 3305
rect 6677 3285 6686 3305
rect 6642 3269 6686 3285
rect 6751 3301 6800 3311
rect 6751 3281 6762 3301
rect 6782 3281 6800 3301
rect 6751 3269 6800 3281
rect 6850 3305 6894 3311
rect 6850 3285 6865 3305
rect 6885 3285 6894 3305
rect 6850 3269 6894 3285
rect 6964 3305 7008 3311
rect 6964 3285 6973 3305
rect 6993 3285 7008 3305
rect 6964 3269 7008 3285
rect 7058 3301 7107 3311
rect 7058 3281 7076 3301
rect 7096 3281 7107 3301
rect 7058 3269 7107 3281
rect 12915 3437 12964 3449
rect 12915 3417 12926 3437
rect 12946 3417 12964 3437
rect 12915 3407 12964 3417
rect 13014 3433 13058 3449
rect 13014 3413 13029 3433
rect 13049 3413 13058 3433
rect 13014 3407 13058 3413
rect 13128 3433 13172 3449
rect 13128 3413 13137 3433
rect 13157 3413 13172 3433
rect 13128 3407 13172 3413
rect 13222 3437 13271 3449
rect 13222 3417 13240 3437
rect 13260 3417 13271 3437
rect 13222 3407 13271 3417
rect 13336 3433 13380 3449
rect 13336 3413 13345 3433
rect 13365 3413 13380 3433
rect 13336 3407 13380 3413
rect 13430 3437 13479 3449
rect 13430 3417 13448 3437
rect 13468 3417 13479 3437
rect 13430 3407 13479 3417
rect 13549 3433 13593 3449
rect 13549 3413 13558 3433
rect 13578 3413 13593 3433
rect 13549 3407 13593 3413
rect 13643 3437 13692 3449
rect 13643 3417 13661 3437
rect 13681 3417 13692 3437
rect 13643 3407 13692 3417
rect 3822 3188 3871 3200
rect 3822 3168 3833 3188
rect 3853 3168 3871 3188
rect 3822 3158 3871 3168
rect 3921 3184 3965 3200
rect 3921 3164 3936 3184
rect 3956 3164 3965 3184
rect 3921 3158 3965 3164
rect 4035 3184 4079 3200
rect 4035 3164 4044 3184
rect 4064 3164 4079 3184
rect 4035 3158 4079 3164
rect 4129 3188 4178 3200
rect 4129 3168 4147 3188
rect 4167 3168 4178 3188
rect 4129 3158 4178 3168
rect 4243 3184 4287 3200
rect 4243 3164 4252 3184
rect 4272 3164 4287 3184
rect 4243 3158 4287 3164
rect 4337 3188 4386 3200
rect 4337 3168 4355 3188
rect 4375 3168 4386 3188
rect 4337 3158 4386 3168
rect 4456 3184 4500 3200
rect 4456 3164 4465 3184
rect 4485 3164 4500 3184
rect 4456 3158 4500 3164
rect 4550 3188 4599 3200
rect 4550 3168 4568 3188
rect 4588 3168 4599 3188
rect 4550 3158 4599 3168
rect 8878 3229 8927 3241
rect 8878 3209 8889 3229
rect 8909 3209 8927 3229
rect 8878 3199 8927 3209
rect 8977 3225 9021 3241
rect 8977 3205 8992 3225
rect 9012 3205 9021 3225
rect 8977 3199 9021 3205
rect 9091 3225 9135 3241
rect 9091 3205 9100 3225
rect 9120 3205 9135 3225
rect 9091 3199 9135 3205
rect 9185 3229 9234 3241
rect 9185 3209 9203 3229
rect 9223 3209 9234 3229
rect 9185 3199 9234 3209
rect 9299 3225 9343 3241
rect 9299 3205 9308 3225
rect 9328 3205 9343 3225
rect 9299 3199 9343 3205
rect 9393 3229 9442 3241
rect 9393 3209 9411 3229
rect 9431 3209 9442 3229
rect 9393 3199 9442 3209
rect 9512 3225 9556 3241
rect 9512 3205 9521 3225
rect 9541 3205 9556 3225
rect 9512 3199 9556 3205
rect 9606 3229 9655 3241
rect 9606 3209 9624 3229
rect 9644 3209 9655 3229
rect 9606 3199 9655 3209
rect 11305 3265 11354 3275
rect 11305 3245 11316 3265
rect 11336 3245 11354 3265
rect 11305 3233 11354 3245
rect 11404 3269 11448 3275
rect 11404 3249 11419 3269
rect 11439 3249 11448 3269
rect 11404 3233 11448 3249
rect 11518 3265 11567 3275
rect 11518 3245 11529 3265
rect 11549 3245 11567 3265
rect 11518 3233 11567 3245
rect 11617 3269 11661 3275
rect 11617 3249 11632 3269
rect 11652 3249 11661 3269
rect 11617 3233 11661 3249
rect 11726 3265 11775 3275
rect 11726 3245 11737 3265
rect 11757 3245 11775 3265
rect 11726 3233 11775 3245
rect 11825 3269 11869 3275
rect 11825 3249 11840 3269
rect 11860 3249 11869 3269
rect 11825 3233 11869 3249
rect 11939 3269 11983 3275
rect 11939 3249 11948 3269
rect 11968 3249 11983 3269
rect 11939 3233 11983 3249
rect 12033 3265 12082 3275
rect 12033 3245 12051 3265
rect 12071 3245 12082 3265
rect 12033 3233 12082 3245
rect 17971 3478 18020 3490
rect 17971 3458 17982 3478
rect 18002 3458 18020 3478
rect 17971 3448 18020 3458
rect 18070 3474 18114 3490
rect 18070 3454 18085 3474
rect 18105 3454 18114 3474
rect 18070 3448 18114 3454
rect 18184 3474 18228 3490
rect 18184 3454 18193 3474
rect 18213 3454 18228 3474
rect 18184 3448 18228 3454
rect 18278 3478 18327 3490
rect 18278 3458 18296 3478
rect 18316 3458 18327 3478
rect 18278 3448 18327 3458
rect 18392 3474 18436 3490
rect 18392 3454 18401 3474
rect 18421 3454 18436 3474
rect 18392 3448 18436 3454
rect 18486 3478 18535 3490
rect 18486 3458 18504 3478
rect 18524 3458 18535 3478
rect 18486 3448 18535 3458
rect 18605 3474 18649 3490
rect 18605 3454 18614 3474
rect 18634 3454 18649 3474
rect 18605 3448 18649 3454
rect 18699 3478 18748 3490
rect 18699 3458 18717 3478
rect 18737 3458 18748 3478
rect 18699 3448 18748 3458
rect 16361 3306 16410 3316
rect 16361 3286 16372 3306
rect 16392 3286 16410 3306
rect 16361 3274 16410 3286
rect 16460 3310 16504 3316
rect 16460 3290 16475 3310
rect 16495 3290 16504 3310
rect 16460 3274 16504 3290
rect 16574 3306 16623 3316
rect 16574 3286 16585 3306
rect 16605 3286 16623 3306
rect 16574 3274 16623 3286
rect 16673 3310 16717 3316
rect 16673 3290 16688 3310
rect 16708 3290 16717 3310
rect 16673 3274 16717 3290
rect 16782 3306 16831 3316
rect 16782 3286 16793 3306
rect 16813 3286 16831 3306
rect 16782 3274 16831 3286
rect 16881 3310 16925 3316
rect 16881 3290 16896 3310
rect 16916 3290 16925 3310
rect 16881 3274 16925 3290
rect 16995 3310 17039 3316
rect 16995 3290 17004 3310
rect 17024 3290 17039 3310
rect 16995 3274 17039 3290
rect 17089 3306 17138 3316
rect 17089 3286 17107 3306
rect 17127 3286 17138 3306
rect 17089 3274 17138 3286
rect 13853 3193 13902 3205
rect 13853 3173 13864 3193
rect 13884 3173 13902 3193
rect 13853 3163 13902 3173
rect 13952 3189 13996 3205
rect 13952 3169 13967 3189
rect 13987 3169 13996 3189
rect 13952 3163 13996 3169
rect 14066 3189 14110 3205
rect 14066 3169 14075 3189
rect 14095 3169 14110 3189
rect 14066 3163 14110 3169
rect 14160 3193 14209 3205
rect 14160 3173 14178 3193
rect 14198 3173 14209 3193
rect 14160 3163 14209 3173
rect 14274 3189 14318 3205
rect 14274 3169 14283 3189
rect 14303 3169 14318 3189
rect 14274 3163 14318 3169
rect 14368 3193 14417 3205
rect 14368 3173 14386 3193
rect 14406 3173 14417 3193
rect 14368 3163 14417 3173
rect 14487 3189 14531 3205
rect 14487 3169 14496 3189
rect 14516 3169 14531 3189
rect 14487 3163 14531 3169
rect 14581 3193 14630 3205
rect 14581 3173 14599 3193
rect 14619 3173 14630 3193
rect 14581 3163 14630 3173
rect 5391 2991 5440 3001
rect 5391 2971 5402 2991
rect 5422 2971 5440 2991
rect 335 2950 384 2960
rect 335 2930 346 2950
rect 366 2930 384 2950
rect 335 2918 384 2930
rect 434 2954 478 2960
rect 434 2934 449 2954
rect 469 2934 478 2954
rect 434 2918 478 2934
rect 548 2950 597 2960
rect 548 2930 559 2950
rect 579 2930 597 2950
rect 548 2918 597 2930
rect 647 2954 691 2960
rect 647 2934 662 2954
rect 682 2934 691 2954
rect 647 2918 691 2934
rect 756 2950 805 2960
rect 756 2930 767 2950
rect 787 2930 805 2950
rect 756 2918 805 2930
rect 855 2954 899 2960
rect 855 2934 870 2954
rect 890 2934 899 2954
rect 855 2918 899 2934
rect 969 2954 1013 2960
rect 969 2934 978 2954
rect 998 2934 1013 2954
rect 969 2918 1013 2934
rect 1063 2950 1112 2960
rect 1063 2930 1081 2950
rect 1101 2930 1112 2950
rect 1063 2918 1112 2930
rect 2774 2908 2823 2920
rect 2774 2888 2785 2908
rect 2805 2888 2823 2908
rect 2774 2878 2823 2888
rect 2873 2904 2917 2920
rect 2873 2884 2888 2904
rect 2908 2884 2917 2904
rect 2873 2878 2917 2884
rect 2987 2904 3031 2920
rect 2987 2884 2996 2904
rect 3016 2884 3031 2904
rect 2987 2878 3031 2884
rect 3081 2908 3130 2920
rect 3081 2888 3099 2908
rect 3119 2888 3130 2908
rect 3081 2878 3130 2888
rect 3195 2904 3239 2920
rect 3195 2884 3204 2904
rect 3224 2884 3239 2904
rect 3195 2878 3239 2884
rect 3289 2908 3338 2920
rect 3289 2888 3307 2908
rect 3327 2888 3338 2908
rect 3289 2878 3338 2888
rect 3408 2904 3452 2920
rect 3408 2884 3417 2904
rect 3437 2884 3452 2904
rect 3408 2878 3452 2884
rect 3502 2908 3551 2920
rect 3502 2888 3520 2908
rect 3540 2888 3551 2908
rect 5391 2959 5440 2971
rect 5490 2995 5534 3001
rect 5490 2975 5505 2995
rect 5525 2975 5534 2995
rect 5490 2959 5534 2975
rect 5604 2991 5653 3001
rect 5604 2971 5615 2991
rect 5635 2971 5653 2991
rect 5604 2959 5653 2971
rect 5703 2995 5747 3001
rect 5703 2975 5718 2995
rect 5738 2975 5747 2995
rect 5703 2959 5747 2975
rect 5812 2991 5861 3001
rect 5812 2971 5823 2991
rect 5843 2971 5861 2991
rect 5812 2959 5861 2971
rect 5911 2995 5955 3001
rect 5911 2975 5926 2995
rect 5946 2975 5955 2995
rect 5911 2959 5955 2975
rect 6025 2995 6069 3001
rect 6025 2975 6034 2995
rect 6054 2975 6069 2995
rect 6025 2959 6069 2975
rect 6119 2991 6168 3001
rect 6119 2971 6137 2991
rect 6157 2971 6168 2991
rect 6119 2959 6168 2971
rect 7830 2949 7879 2961
rect 7830 2929 7841 2949
rect 7861 2929 7879 2949
rect 3502 2878 3551 2888
rect 7830 2919 7879 2929
rect 7929 2945 7973 2961
rect 7929 2925 7944 2945
rect 7964 2925 7973 2945
rect 7929 2919 7973 2925
rect 8043 2945 8087 2961
rect 8043 2925 8052 2945
rect 8072 2925 8087 2945
rect 8043 2919 8087 2925
rect 8137 2949 8186 2961
rect 8137 2929 8155 2949
rect 8175 2929 8186 2949
rect 8137 2919 8186 2929
rect 8251 2945 8295 2961
rect 8251 2925 8260 2945
rect 8280 2925 8295 2945
rect 8251 2919 8295 2925
rect 8345 2949 8394 2961
rect 8345 2929 8363 2949
rect 8383 2929 8394 2949
rect 8345 2919 8394 2929
rect 8464 2945 8508 2961
rect 8464 2925 8473 2945
rect 8493 2925 8508 2945
rect 8464 2919 8508 2925
rect 8558 2949 8607 2961
rect 8558 2929 8576 2949
rect 8596 2929 8607 2949
rect 18909 3234 18958 3246
rect 18909 3214 18920 3234
rect 18940 3214 18958 3234
rect 18909 3204 18958 3214
rect 19008 3230 19052 3246
rect 19008 3210 19023 3230
rect 19043 3210 19052 3230
rect 19008 3204 19052 3210
rect 19122 3230 19166 3246
rect 19122 3210 19131 3230
rect 19151 3210 19166 3230
rect 19122 3204 19166 3210
rect 19216 3234 19265 3246
rect 19216 3214 19234 3234
rect 19254 3214 19265 3234
rect 19216 3204 19265 3214
rect 19330 3230 19374 3246
rect 19330 3210 19339 3230
rect 19359 3210 19374 3230
rect 19330 3204 19374 3210
rect 19424 3234 19473 3246
rect 19424 3214 19442 3234
rect 19462 3214 19473 3234
rect 19424 3204 19473 3214
rect 19543 3230 19587 3246
rect 19543 3210 19552 3230
rect 19572 3210 19587 3230
rect 19543 3204 19587 3210
rect 19637 3234 19686 3246
rect 19637 3214 19655 3234
rect 19675 3214 19686 3234
rect 19637 3204 19686 3214
rect 15422 2996 15471 3006
rect 15422 2976 15433 2996
rect 15453 2976 15471 2996
rect 8558 2919 8607 2929
rect 10366 2955 10415 2965
rect 10366 2935 10377 2955
rect 10397 2935 10415 2955
rect 10366 2923 10415 2935
rect 10465 2959 10509 2965
rect 10465 2939 10480 2959
rect 10500 2939 10509 2959
rect 10465 2923 10509 2939
rect 10579 2955 10628 2965
rect 10579 2935 10590 2955
rect 10610 2935 10628 2955
rect 10579 2923 10628 2935
rect 10678 2959 10722 2965
rect 10678 2939 10693 2959
rect 10713 2939 10722 2959
rect 10678 2923 10722 2939
rect 10787 2955 10836 2965
rect 10787 2935 10798 2955
rect 10818 2935 10836 2955
rect 10787 2923 10836 2935
rect 10886 2959 10930 2965
rect 10886 2939 10901 2959
rect 10921 2939 10930 2959
rect 10886 2923 10930 2939
rect 11000 2959 11044 2965
rect 11000 2939 11009 2959
rect 11029 2939 11044 2959
rect 11000 2923 11044 2939
rect 11094 2955 11143 2965
rect 11094 2935 11112 2955
rect 11132 2935 11143 2955
rect 11094 2923 11143 2935
rect 12805 2913 12854 2925
rect 12805 2893 12816 2913
rect 12836 2893 12854 2913
rect 12805 2883 12854 2893
rect 12904 2909 12948 2925
rect 12904 2889 12919 2909
rect 12939 2889 12948 2909
rect 12904 2883 12948 2889
rect 13018 2909 13062 2925
rect 13018 2889 13027 2909
rect 13047 2889 13062 2909
rect 13018 2883 13062 2889
rect 13112 2913 13161 2925
rect 13112 2893 13130 2913
rect 13150 2893 13161 2913
rect 13112 2883 13161 2893
rect 13226 2909 13270 2925
rect 13226 2889 13235 2909
rect 13255 2889 13270 2909
rect 13226 2883 13270 2889
rect 13320 2913 13369 2925
rect 13320 2893 13338 2913
rect 13358 2893 13369 2913
rect 13320 2883 13369 2893
rect 13439 2909 13483 2925
rect 13439 2889 13448 2909
rect 13468 2889 13483 2909
rect 13439 2883 13483 2889
rect 13533 2913 13582 2925
rect 13533 2893 13551 2913
rect 13571 2893 13582 2913
rect 15422 2964 15471 2976
rect 15521 3000 15565 3006
rect 15521 2980 15536 3000
rect 15556 2980 15565 3000
rect 15521 2964 15565 2980
rect 15635 2996 15684 3006
rect 15635 2976 15646 2996
rect 15666 2976 15684 2996
rect 15635 2964 15684 2976
rect 15734 3000 15778 3006
rect 15734 2980 15749 3000
rect 15769 2980 15778 3000
rect 15734 2964 15778 2980
rect 15843 2996 15892 3006
rect 15843 2976 15854 2996
rect 15874 2976 15892 2996
rect 15843 2964 15892 2976
rect 15942 3000 15986 3006
rect 15942 2980 15957 3000
rect 15977 2980 15986 3000
rect 15942 2964 15986 2980
rect 16056 3000 16100 3006
rect 16056 2980 16065 3000
rect 16085 2980 16100 3000
rect 16056 2964 16100 2980
rect 16150 2996 16199 3006
rect 16150 2976 16168 2996
rect 16188 2976 16199 2996
rect 16150 2964 16199 2976
rect 17861 2954 17910 2966
rect 17861 2934 17872 2954
rect 17892 2934 17910 2954
rect 13533 2883 13582 2893
rect 17861 2924 17910 2934
rect 17960 2950 18004 2966
rect 17960 2930 17975 2950
rect 17995 2930 18004 2950
rect 17960 2924 18004 2930
rect 18074 2950 18118 2966
rect 18074 2930 18083 2950
rect 18103 2930 18118 2950
rect 18074 2924 18118 2930
rect 18168 2954 18217 2966
rect 18168 2934 18186 2954
rect 18206 2934 18217 2954
rect 18168 2924 18217 2934
rect 18282 2950 18326 2966
rect 18282 2930 18291 2950
rect 18311 2930 18326 2950
rect 18282 2924 18326 2930
rect 18376 2954 18425 2966
rect 18376 2934 18394 2954
rect 18414 2934 18425 2954
rect 18376 2924 18425 2934
rect 18495 2950 18539 2966
rect 18495 2930 18504 2950
rect 18524 2930 18539 2950
rect 18495 2924 18539 2930
rect 18589 2954 18638 2966
rect 18589 2934 18607 2954
rect 18627 2934 18638 2954
rect 18589 2924 18638 2934
rect 1384 2681 1433 2691
rect 1384 2661 1395 2681
rect 1415 2661 1433 2681
rect 1384 2649 1433 2661
rect 1483 2685 1527 2691
rect 1483 2665 1498 2685
rect 1518 2665 1527 2685
rect 1483 2649 1527 2665
rect 1597 2681 1646 2691
rect 1597 2661 1608 2681
rect 1628 2661 1646 2681
rect 1597 2649 1646 2661
rect 1696 2685 1740 2691
rect 1696 2665 1711 2685
rect 1731 2665 1740 2685
rect 1696 2649 1740 2665
rect 1805 2681 1854 2691
rect 1805 2661 1816 2681
rect 1836 2661 1854 2681
rect 1805 2649 1854 2661
rect 1904 2685 1948 2691
rect 1904 2665 1919 2685
rect 1939 2665 1948 2685
rect 1904 2649 1948 2665
rect 2018 2685 2062 2691
rect 2018 2665 2027 2685
rect 2047 2665 2062 2685
rect 2018 2649 2062 2665
rect 2112 2681 2161 2691
rect 6440 2722 6489 2732
rect 2112 2661 2130 2681
rect 2150 2661 2161 2681
rect 2112 2649 2161 2661
rect 3823 2639 3872 2651
rect 3823 2619 3834 2639
rect 3854 2619 3872 2639
rect 3823 2609 3872 2619
rect 3922 2635 3966 2651
rect 3922 2615 3937 2635
rect 3957 2615 3966 2635
rect 3922 2609 3966 2615
rect 4036 2635 4080 2651
rect 4036 2615 4045 2635
rect 4065 2615 4080 2635
rect 4036 2609 4080 2615
rect 4130 2639 4179 2651
rect 4130 2619 4148 2639
rect 4168 2619 4179 2639
rect 4130 2609 4179 2619
rect 4244 2635 4288 2651
rect 4244 2615 4253 2635
rect 4273 2615 4288 2635
rect 4244 2609 4288 2615
rect 4338 2639 4387 2651
rect 4338 2619 4356 2639
rect 4376 2619 4387 2639
rect 4338 2609 4387 2619
rect 4457 2635 4501 2651
rect 4457 2615 4466 2635
rect 4486 2615 4501 2635
rect 4457 2609 4501 2615
rect 4551 2639 4600 2651
rect 6440 2702 6451 2722
rect 6471 2702 6489 2722
rect 6440 2690 6489 2702
rect 6539 2726 6583 2732
rect 6539 2706 6554 2726
rect 6574 2706 6583 2726
rect 6539 2690 6583 2706
rect 6653 2722 6702 2732
rect 6653 2702 6664 2722
rect 6684 2702 6702 2722
rect 6653 2690 6702 2702
rect 6752 2726 6796 2732
rect 6752 2706 6767 2726
rect 6787 2706 6796 2726
rect 6752 2690 6796 2706
rect 6861 2722 6910 2732
rect 6861 2702 6872 2722
rect 6892 2702 6910 2722
rect 6861 2690 6910 2702
rect 6960 2726 7004 2732
rect 6960 2706 6975 2726
rect 6995 2706 7004 2726
rect 6960 2690 7004 2706
rect 7074 2726 7118 2732
rect 7074 2706 7083 2726
rect 7103 2706 7118 2726
rect 7074 2690 7118 2706
rect 7168 2722 7217 2732
rect 7168 2702 7186 2722
rect 7206 2702 7217 2722
rect 7168 2690 7217 2702
rect 8879 2680 8928 2692
rect 8879 2660 8890 2680
rect 8910 2660 8928 2680
rect 8879 2650 8928 2660
rect 8978 2676 9022 2692
rect 8978 2656 8993 2676
rect 9013 2656 9022 2676
rect 8978 2650 9022 2656
rect 9092 2676 9136 2692
rect 9092 2656 9101 2676
rect 9121 2656 9136 2676
rect 9092 2650 9136 2656
rect 9186 2680 9235 2692
rect 9186 2660 9204 2680
rect 9224 2660 9235 2680
rect 9186 2650 9235 2660
rect 9300 2676 9344 2692
rect 9300 2656 9309 2676
rect 9329 2656 9344 2676
rect 9300 2650 9344 2656
rect 9394 2680 9443 2692
rect 9394 2660 9412 2680
rect 9432 2660 9443 2680
rect 9394 2650 9443 2660
rect 9513 2676 9557 2692
rect 9513 2656 9522 2676
rect 9542 2656 9557 2676
rect 9513 2650 9557 2656
rect 9607 2680 9656 2692
rect 9607 2660 9625 2680
rect 9645 2660 9656 2680
rect 9607 2650 9656 2660
rect 11415 2686 11464 2696
rect 4551 2619 4569 2639
rect 4589 2619 4600 2639
rect 4551 2609 4600 2619
rect 336 2401 385 2411
rect 336 2381 347 2401
rect 367 2381 385 2401
rect 336 2369 385 2381
rect 435 2405 479 2411
rect 435 2385 450 2405
rect 470 2385 479 2405
rect 435 2369 479 2385
rect 549 2401 598 2411
rect 549 2381 560 2401
rect 580 2381 598 2401
rect 549 2369 598 2381
rect 648 2405 692 2411
rect 648 2385 663 2405
rect 683 2385 692 2405
rect 648 2369 692 2385
rect 757 2401 806 2411
rect 757 2381 768 2401
rect 788 2381 806 2401
rect 757 2369 806 2381
rect 856 2405 900 2411
rect 856 2385 871 2405
rect 891 2385 900 2405
rect 856 2369 900 2385
rect 970 2405 1014 2411
rect 970 2385 979 2405
rect 999 2385 1014 2405
rect 970 2369 1014 2385
rect 1064 2401 1113 2411
rect 1064 2381 1082 2401
rect 1102 2381 1113 2401
rect 1064 2369 1113 2381
rect 11415 2666 11426 2686
rect 11446 2666 11464 2686
rect 11415 2654 11464 2666
rect 11514 2690 11558 2696
rect 11514 2670 11529 2690
rect 11549 2670 11558 2690
rect 11514 2654 11558 2670
rect 11628 2686 11677 2696
rect 11628 2666 11639 2686
rect 11659 2666 11677 2686
rect 11628 2654 11677 2666
rect 11727 2690 11771 2696
rect 11727 2670 11742 2690
rect 11762 2670 11771 2690
rect 11727 2654 11771 2670
rect 11836 2686 11885 2696
rect 11836 2666 11847 2686
rect 11867 2666 11885 2686
rect 11836 2654 11885 2666
rect 11935 2690 11979 2696
rect 11935 2670 11950 2690
rect 11970 2670 11979 2690
rect 11935 2654 11979 2670
rect 12049 2690 12093 2696
rect 12049 2670 12058 2690
rect 12078 2670 12093 2690
rect 12049 2654 12093 2670
rect 12143 2686 12192 2696
rect 16471 2727 16520 2737
rect 12143 2666 12161 2686
rect 12181 2666 12192 2686
rect 12143 2654 12192 2666
rect 13854 2644 13903 2656
rect 13854 2624 13865 2644
rect 13885 2624 13903 2644
rect 13854 2614 13903 2624
rect 13953 2640 13997 2656
rect 13953 2620 13968 2640
rect 13988 2620 13997 2640
rect 13953 2614 13997 2620
rect 14067 2640 14111 2656
rect 14067 2620 14076 2640
rect 14096 2620 14111 2640
rect 14067 2614 14111 2620
rect 14161 2644 14210 2656
rect 14161 2624 14179 2644
rect 14199 2624 14210 2644
rect 14161 2614 14210 2624
rect 14275 2640 14319 2656
rect 14275 2620 14284 2640
rect 14304 2620 14319 2640
rect 14275 2614 14319 2620
rect 14369 2644 14418 2656
rect 14369 2624 14387 2644
rect 14407 2624 14418 2644
rect 14369 2614 14418 2624
rect 14488 2640 14532 2656
rect 14488 2620 14497 2640
rect 14517 2620 14532 2640
rect 14488 2614 14532 2620
rect 14582 2644 14631 2656
rect 16471 2707 16482 2727
rect 16502 2707 16520 2727
rect 16471 2695 16520 2707
rect 16570 2731 16614 2737
rect 16570 2711 16585 2731
rect 16605 2711 16614 2731
rect 16570 2695 16614 2711
rect 16684 2727 16733 2737
rect 16684 2707 16695 2727
rect 16715 2707 16733 2727
rect 16684 2695 16733 2707
rect 16783 2731 16827 2737
rect 16783 2711 16798 2731
rect 16818 2711 16827 2731
rect 16783 2695 16827 2711
rect 16892 2727 16941 2737
rect 16892 2707 16903 2727
rect 16923 2707 16941 2727
rect 16892 2695 16941 2707
rect 16991 2731 17035 2737
rect 16991 2711 17006 2731
rect 17026 2711 17035 2731
rect 16991 2695 17035 2711
rect 17105 2731 17149 2737
rect 17105 2711 17114 2731
rect 17134 2711 17149 2731
rect 17105 2695 17149 2711
rect 17199 2727 17248 2737
rect 17199 2707 17217 2727
rect 17237 2707 17248 2727
rect 17199 2695 17248 2707
rect 18910 2685 18959 2697
rect 18910 2665 18921 2685
rect 18941 2665 18959 2685
rect 18910 2655 18959 2665
rect 19009 2681 19053 2697
rect 19009 2661 19024 2681
rect 19044 2661 19053 2681
rect 19009 2655 19053 2661
rect 19123 2681 19167 2697
rect 19123 2661 19132 2681
rect 19152 2661 19167 2681
rect 19123 2655 19167 2661
rect 19217 2685 19266 2697
rect 19217 2665 19235 2685
rect 19255 2665 19266 2685
rect 19217 2655 19266 2665
rect 19331 2681 19375 2697
rect 19331 2661 19340 2681
rect 19360 2661 19375 2681
rect 19331 2655 19375 2661
rect 19425 2685 19474 2697
rect 19425 2665 19443 2685
rect 19463 2665 19474 2685
rect 19425 2655 19474 2665
rect 19544 2681 19588 2697
rect 19544 2661 19553 2681
rect 19573 2661 19588 2681
rect 19544 2655 19588 2661
rect 19638 2685 19687 2697
rect 19638 2665 19656 2685
rect 19676 2665 19687 2685
rect 19638 2655 19687 2665
rect 14582 2624 14600 2644
rect 14620 2624 14631 2644
rect 14582 2614 14631 2624
rect 5392 2442 5441 2452
rect 5392 2422 5403 2442
rect 5423 2422 5441 2442
rect 5392 2410 5441 2422
rect 5491 2446 5535 2452
rect 5491 2426 5506 2446
rect 5526 2426 5535 2446
rect 5491 2410 5535 2426
rect 5605 2442 5654 2452
rect 5605 2422 5616 2442
rect 5636 2422 5654 2442
rect 5605 2410 5654 2422
rect 5704 2446 5748 2452
rect 5704 2426 5719 2446
rect 5739 2426 5748 2446
rect 5704 2410 5748 2426
rect 5813 2442 5862 2452
rect 5813 2422 5824 2442
rect 5844 2422 5862 2442
rect 5813 2410 5862 2422
rect 5912 2446 5956 2452
rect 5912 2426 5927 2446
rect 5947 2426 5956 2446
rect 5912 2410 5956 2426
rect 6026 2446 6070 2452
rect 6026 2426 6035 2446
rect 6055 2426 6070 2446
rect 6026 2410 6070 2426
rect 6120 2442 6169 2452
rect 6120 2422 6138 2442
rect 6158 2422 6169 2442
rect 6120 2410 6169 2422
rect 2884 2329 2933 2341
rect 2884 2309 2895 2329
rect 2915 2309 2933 2329
rect 2884 2299 2933 2309
rect 2983 2325 3027 2341
rect 2983 2305 2998 2325
rect 3018 2305 3027 2325
rect 2983 2299 3027 2305
rect 3097 2325 3141 2341
rect 3097 2305 3106 2325
rect 3126 2305 3141 2325
rect 3097 2299 3141 2305
rect 3191 2329 3240 2341
rect 3191 2309 3209 2329
rect 3229 2309 3240 2329
rect 3191 2299 3240 2309
rect 3305 2325 3349 2341
rect 3305 2305 3314 2325
rect 3334 2305 3349 2325
rect 3305 2299 3349 2305
rect 3399 2329 3448 2341
rect 3399 2309 3417 2329
rect 3437 2309 3448 2329
rect 3399 2299 3448 2309
rect 3518 2325 3562 2341
rect 3518 2305 3527 2325
rect 3547 2305 3562 2325
rect 3518 2299 3562 2305
rect 3612 2329 3661 2341
rect 3612 2309 3630 2329
rect 3650 2309 3661 2329
rect 3612 2299 3661 2309
rect 1274 2157 1323 2167
rect 1274 2137 1285 2157
rect 1305 2137 1323 2157
rect 1274 2125 1323 2137
rect 1373 2161 1417 2167
rect 1373 2141 1388 2161
rect 1408 2141 1417 2161
rect 1373 2125 1417 2141
rect 1487 2157 1536 2167
rect 1487 2137 1498 2157
rect 1518 2137 1536 2157
rect 1487 2125 1536 2137
rect 1586 2161 1630 2167
rect 1586 2141 1601 2161
rect 1621 2141 1630 2161
rect 1586 2125 1630 2141
rect 1695 2157 1744 2167
rect 1695 2137 1706 2157
rect 1726 2137 1744 2157
rect 1695 2125 1744 2137
rect 1794 2161 1838 2167
rect 1794 2141 1809 2161
rect 1829 2141 1838 2161
rect 1794 2125 1838 2141
rect 1908 2161 1952 2167
rect 1908 2141 1917 2161
rect 1937 2141 1952 2161
rect 1908 2125 1952 2141
rect 2002 2157 2051 2167
rect 2002 2137 2020 2157
rect 2040 2137 2051 2157
rect 2002 2125 2051 2137
rect 7940 2370 7989 2382
rect 7940 2350 7951 2370
rect 7971 2350 7989 2370
rect 7940 2340 7989 2350
rect 8039 2366 8083 2382
rect 8039 2346 8054 2366
rect 8074 2346 8083 2366
rect 8039 2340 8083 2346
rect 8153 2366 8197 2382
rect 8153 2346 8162 2366
rect 8182 2346 8197 2366
rect 8153 2340 8197 2346
rect 8247 2370 8296 2382
rect 8247 2350 8265 2370
rect 8285 2350 8296 2370
rect 8247 2340 8296 2350
rect 8361 2366 8405 2382
rect 8361 2346 8370 2366
rect 8390 2346 8405 2366
rect 8361 2340 8405 2346
rect 8455 2370 8504 2382
rect 8455 2350 8473 2370
rect 8493 2350 8504 2370
rect 8455 2340 8504 2350
rect 8574 2366 8618 2382
rect 8574 2346 8583 2366
rect 8603 2346 8618 2366
rect 8574 2340 8618 2346
rect 8668 2370 8717 2382
rect 8668 2350 8686 2370
rect 8706 2350 8717 2370
rect 8668 2340 8717 2350
rect 10367 2406 10416 2416
rect 10367 2386 10378 2406
rect 10398 2386 10416 2406
rect 10367 2374 10416 2386
rect 10466 2410 10510 2416
rect 10466 2390 10481 2410
rect 10501 2390 10510 2410
rect 10466 2374 10510 2390
rect 10580 2406 10629 2416
rect 10580 2386 10591 2406
rect 10611 2386 10629 2406
rect 10580 2374 10629 2386
rect 10679 2410 10723 2416
rect 10679 2390 10694 2410
rect 10714 2390 10723 2410
rect 10679 2374 10723 2390
rect 10788 2406 10837 2416
rect 10788 2386 10799 2406
rect 10819 2386 10837 2406
rect 10788 2374 10837 2386
rect 10887 2410 10931 2416
rect 10887 2390 10902 2410
rect 10922 2390 10931 2410
rect 10887 2374 10931 2390
rect 11001 2410 11045 2416
rect 11001 2390 11010 2410
rect 11030 2390 11045 2410
rect 11001 2374 11045 2390
rect 11095 2406 11144 2416
rect 11095 2386 11113 2406
rect 11133 2386 11144 2406
rect 11095 2374 11144 2386
rect 15423 2447 15472 2457
rect 15423 2427 15434 2447
rect 15454 2427 15472 2447
rect 15423 2415 15472 2427
rect 15522 2451 15566 2457
rect 15522 2431 15537 2451
rect 15557 2431 15566 2451
rect 15522 2415 15566 2431
rect 15636 2447 15685 2457
rect 15636 2427 15647 2447
rect 15667 2427 15685 2447
rect 15636 2415 15685 2427
rect 15735 2451 15779 2457
rect 15735 2431 15750 2451
rect 15770 2431 15779 2451
rect 15735 2415 15779 2431
rect 15844 2447 15893 2457
rect 15844 2427 15855 2447
rect 15875 2427 15893 2447
rect 15844 2415 15893 2427
rect 15943 2451 15987 2457
rect 15943 2431 15958 2451
rect 15978 2431 15987 2451
rect 15943 2415 15987 2431
rect 16057 2451 16101 2457
rect 16057 2431 16066 2451
rect 16086 2431 16101 2451
rect 16057 2415 16101 2431
rect 16151 2447 16200 2457
rect 16151 2427 16169 2447
rect 16189 2427 16200 2447
rect 16151 2415 16200 2427
rect 6330 2198 6379 2208
rect 6330 2178 6341 2198
rect 6361 2178 6379 2198
rect 6330 2166 6379 2178
rect 6429 2202 6473 2208
rect 6429 2182 6444 2202
rect 6464 2182 6473 2202
rect 6429 2166 6473 2182
rect 6543 2198 6592 2208
rect 6543 2178 6554 2198
rect 6574 2178 6592 2198
rect 6543 2166 6592 2178
rect 6642 2202 6686 2208
rect 6642 2182 6657 2202
rect 6677 2182 6686 2202
rect 6642 2166 6686 2182
rect 6751 2198 6800 2208
rect 6751 2178 6762 2198
rect 6782 2178 6800 2198
rect 6751 2166 6800 2178
rect 6850 2202 6894 2208
rect 6850 2182 6865 2202
rect 6885 2182 6894 2202
rect 6850 2166 6894 2182
rect 6964 2202 7008 2208
rect 6964 2182 6973 2202
rect 6993 2182 7008 2202
rect 6964 2166 7008 2182
rect 7058 2198 7107 2208
rect 7058 2178 7076 2198
rect 7096 2178 7107 2198
rect 7058 2166 7107 2178
rect 12915 2334 12964 2346
rect 12915 2314 12926 2334
rect 12946 2314 12964 2334
rect 12915 2304 12964 2314
rect 13014 2330 13058 2346
rect 13014 2310 13029 2330
rect 13049 2310 13058 2330
rect 13014 2304 13058 2310
rect 13128 2330 13172 2346
rect 13128 2310 13137 2330
rect 13157 2310 13172 2330
rect 13128 2304 13172 2310
rect 13222 2334 13271 2346
rect 13222 2314 13240 2334
rect 13260 2314 13271 2334
rect 13222 2304 13271 2314
rect 13336 2330 13380 2346
rect 13336 2310 13345 2330
rect 13365 2310 13380 2330
rect 13336 2304 13380 2310
rect 13430 2334 13479 2346
rect 13430 2314 13448 2334
rect 13468 2314 13479 2334
rect 13430 2304 13479 2314
rect 13549 2330 13593 2346
rect 13549 2310 13558 2330
rect 13578 2310 13593 2330
rect 13549 2304 13593 2310
rect 13643 2334 13692 2346
rect 13643 2314 13661 2334
rect 13681 2314 13692 2334
rect 13643 2304 13692 2314
rect 3822 2085 3871 2097
rect 3822 2065 3833 2085
rect 3853 2065 3871 2085
rect 3822 2055 3871 2065
rect 3921 2081 3965 2097
rect 3921 2061 3936 2081
rect 3956 2061 3965 2081
rect 3921 2055 3965 2061
rect 4035 2081 4079 2097
rect 4035 2061 4044 2081
rect 4064 2061 4079 2081
rect 4035 2055 4079 2061
rect 4129 2085 4178 2097
rect 4129 2065 4147 2085
rect 4167 2065 4178 2085
rect 4129 2055 4178 2065
rect 4243 2081 4287 2097
rect 4243 2061 4252 2081
rect 4272 2061 4287 2081
rect 4243 2055 4287 2061
rect 4337 2085 4386 2097
rect 4337 2065 4355 2085
rect 4375 2065 4386 2085
rect 4337 2055 4386 2065
rect 4456 2081 4500 2097
rect 4456 2061 4465 2081
rect 4485 2061 4500 2081
rect 4456 2055 4500 2061
rect 4550 2085 4599 2097
rect 4550 2065 4568 2085
rect 4588 2065 4599 2085
rect 4550 2055 4599 2065
rect 8878 2126 8927 2138
rect 8878 2106 8889 2126
rect 8909 2106 8927 2126
rect 8878 2096 8927 2106
rect 8977 2122 9021 2138
rect 8977 2102 8992 2122
rect 9012 2102 9021 2122
rect 8977 2096 9021 2102
rect 9091 2122 9135 2138
rect 9091 2102 9100 2122
rect 9120 2102 9135 2122
rect 9091 2096 9135 2102
rect 9185 2126 9234 2138
rect 9185 2106 9203 2126
rect 9223 2106 9234 2126
rect 9185 2096 9234 2106
rect 9299 2122 9343 2138
rect 9299 2102 9308 2122
rect 9328 2102 9343 2122
rect 9299 2096 9343 2102
rect 9393 2126 9442 2138
rect 9393 2106 9411 2126
rect 9431 2106 9442 2126
rect 9393 2096 9442 2106
rect 9512 2122 9556 2138
rect 9512 2102 9521 2122
rect 9541 2102 9556 2122
rect 9512 2096 9556 2102
rect 9606 2126 9655 2138
rect 9606 2106 9624 2126
rect 9644 2106 9655 2126
rect 9606 2096 9655 2106
rect 11305 2162 11354 2172
rect 11305 2142 11316 2162
rect 11336 2142 11354 2162
rect 11305 2130 11354 2142
rect 11404 2166 11448 2172
rect 11404 2146 11419 2166
rect 11439 2146 11448 2166
rect 11404 2130 11448 2146
rect 11518 2162 11567 2172
rect 11518 2142 11529 2162
rect 11549 2142 11567 2162
rect 11518 2130 11567 2142
rect 11617 2166 11661 2172
rect 11617 2146 11632 2166
rect 11652 2146 11661 2166
rect 11617 2130 11661 2146
rect 11726 2162 11775 2172
rect 11726 2142 11737 2162
rect 11757 2142 11775 2162
rect 11726 2130 11775 2142
rect 11825 2166 11869 2172
rect 11825 2146 11840 2166
rect 11860 2146 11869 2166
rect 11825 2130 11869 2146
rect 11939 2166 11983 2172
rect 11939 2146 11948 2166
rect 11968 2146 11983 2166
rect 11939 2130 11983 2146
rect 12033 2162 12082 2172
rect 12033 2142 12051 2162
rect 12071 2142 12082 2162
rect 12033 2130 12082 2142
rect 17971 2375 18020 2387
rect 17971 2355 17982 2375
rect 18002 2355 18020 2375
rect 17971 2345 18020 2355
rect 18070 2371 18114 2387
rect 18070 2351 18085 2371
rect 18105 2351 18114 2371
rect 18070 2345 18114 2351
rect 18184 2371 18228 2387
rect 18184 2351 18193 2371
rect 18213 2351 18228 2371
rect 18184 2345 18228 2351
rect 18278 2375 18327 2387
rect 18278 2355 18296 2375
rect 18316 2355 18327 2375
rect 18278 2345 18327 2355
rect 18392 2371 18436 2387
rect 18392 2351 18401 2371
rect 18421 2351 18436 2371
rect 18392 2345 18436 2351
rect 18486 2375 18535 2387
rect 18486 2355 18504 2375
rect 18524 2355 18535 2375
rect 18486 2345 18535 2355
rect 18605 2371 18649 2387
rect 18605 2351 18614 2371
rect 18634 2351 18649 2371
rect 18605 2345 18649 2351
rect 18699 2375 18748 2387
rect 18699 2355 18717 2375
rect 18737 2355 18748 2375
rect 18699 2345 18748 2355
rect 16361 2203 16410 2213
rect 16361 2183 16372 2203
rect 16392 2183 16410 2203
rect 16361 2171 16410 2183
rect 16460 2207 16504 2213
rect 16460 2187 16475 2207
rect 16495 2187 16504 2207
rect 16460 2171 16504 2187
rect 16574 2203 16623 2213
rect 16574 2183 16585 2203
rect 16605 2183 16623 2203
rect 16574 2171 16623 2183
rect 16673 2207 16717 2213
rect 16673 2187 16688 2207
rect 16708 2187 16717 2207
rect 16673 2171 16717 2187
rect 16782 2203 16831 2213
rect 16782 2183 16793 2203
rect 16813 2183 16831 2203
rect 16782 2171 16831 2183
rect 16881 2207 16925 2213
rect 16881 2187 16896 2207
rect 16916 2187 16925 2207
rect 16881 2171 16925 2187
rect 16995 2207 17039 2213
rect 16995 2187 17004 2207
rect 17024 2187 17039 2207
rect 16995 2171 17039 2187
rect 17089 2203 17138 2213
rect 17089 2183 17107 2203
rect 17127 2183 17138 2203
rect 17089 2171 17138 2183
rect 13853 2090 13902 2102
rect 13853 2070 13864 2090
rect 13884 2070 13902 2090
rect 13853 2060 13902 2070
rect 13952 2086 13996 2102
rect 13952 2066 13967 2086
rect 13987 2066 13996 2086
rect 13952 2060 13996 2066
rect 14066 2086 14110 2102
rect 14066 2066 14075 2086
rect 14095 2066 14110 2086
rect 14066 2060 14110 2066
rect 14160 2090 14209 2102
rect 14160 2070 14178 2090
rect 14198 2070 14209 2090
rect 14160 2060 14209 2070
rect 14274 2086 14318 2102
rect 14274 2066 14283 2086
rect 14303 2066 14318 2086
rect 14274 2060 14318 2066
rect 14368 2090 14417 2102
rect 14368 2070 14386 2090
rect 14406 2070 14417 2090
rect 14368 2060 14417 2070
rect 14487 2086 14531 2102
rect 14487 2066 14496 2086
rect 14516 2066 14531 2086
rect 14487 2060 14531 2066
rect 14581 2090 14630 2102
rect 14581 2070 14599 2090
rect 14619 2070 14630 2090
rect 14581 2060 14630 2070
rect 5391 1888 5440 1898
rect 5391 1868 5402 1888
rect 5422 1868 5440 1888
rect 335 1847 384 1857
rect 335 1827 346 1847
rect 366 1827 384 1847
rect 335 1815 384 1827
rect 434 1851 478 1857
rect 434 1831 449 1851
rect 469 1831 478 1851
rect 434 1815 478 1831
rect 548 1847 597 1857
rect 548 1827 559 1847
rect 579 1827 597 1847
rect 548 1815 597 1827
rect 647 1851 691 1857
rect 647 1831 662 1851
rect 682 1831 691 1851
rect 647 1815 691 1831
rect 756 1847 805 1857
rect 756 1827 767 1847
rect 787 1827 805 1847
rect 756 1815 805 1827
rect 855 1851 899 1857
rect 855 1831 870 1851
rect 890 1831 899 1851
rect 855 1815 899 1831
rect 969 1851 1013 1857
rect 969 1831 978 1851
rect 998 1831 1013 1851
rect 969 1815 1013 1831
rect 1063 1847 1112 1857
rect 1063 1827 1081 1847
rect 1101 1827 1112 1847
rect 1063 1815 1112 1827
rect 2744 1818 2793 1830
rect 2744 1798 2755 1818
rect 2775 1798 2793 1818
rect 2744 1788 2793 1798
rect 2843 1814 2887 1830
rect 2843 1794 2858 1814
rect 2878 1794 2887 1814
rect 2843 1788 2887 1794
rect 2957 1814 3001 1830
rect 2957 1794 2966 1814
rect 2986 1794 3001 1814
rect 2957 1788 3001 1794
rect 3051 1818 3100 1830
rect 3051 1798 3069 1818
rect 3089 1798 3100 1818
rect 3051 1788 3100 1798
rect 3165 1814 3209 1830
rect 3165 1794 3174 1814
rect 3194 1794 3209 1814
rect 3165 1788 3209 1794
rect 3259 1818 3308 1830
rect 3259 1798 3277 1818
rect 3297 1798 3308 1818
rect 3259 1788 3308 1798
rect 3378 1814 3422 1830
rect 3378 1794 3387 1814
rect 3407 1794 3422 1814
rect 3378 1788 3422 1794
rect 3472 1818 3521 1830
rect 3472 1798 3490 1818
rect 3510 1798 3521 1818
rect 3472 1788 3521 1798
rect 5391 1856 5440 1868
rect 5490 1892 5534 1898
rect 5490 1872 5505 1892
rect 5525 1872 5534 1892
rect 5490 1856 5534 1872
rect 5604 1888 5653 1898
rect 5604 1868 5615 1888
rect 5635 1868 5653 1888
rect 5604 1856 5653 1868
rect 5703 1892 5747 1898
rect 5703 1872 5718 1892
rect 5738 1872 5747 1892
rect 5703 1856 5747 1872
rect 5812 1888 5861 1898
rect 5812 1868 5823 1888
rect 5843 1868 5861 1888
rect 5812 1856 5861 1868
rect 5911 1892 5955 1898
rect 5911 1872 5926 1892
rect 5946 1872 5955 1892
rect 5911 1856 5955 1872
rect 6025 1892 6069 1898
rect 6025 1872 6034 1892
rect 6054 1872 6069 1892
rect 6025 1856 6069 1872
rect 6119 1888 6168 1898
rect 6119 1868 6137 1888
rect 6157 1868 6168 1888
rect 6119 1856 6168 1868
rect 7800 1859 7849 1871
rect 7800 1839 7811 1859
rect 7831 1839 7849 1859
rect 7800 1829 7849 1839
rect 7899 1855 7943 1871
rect 7899 1835 7914 1855
rect 7934 1835 7943 1855
rect 7899 1829 7943 1835
rect 8013 1855 8057 1871
rect 8013 1835 8022 1855
rect 8042 1835 8057 1855
rect 8013 1829 8057 1835
rect 8107 1859 8156 1871
rect 8107 1839 8125 1859
rect 8145 1839 8156 1859
rect 8107 1829 8156 1839
rect 8221 1855 8265 1871
rect 8221 1835 8230 1855
rect 8250 1835 8265 1855
rect 8221 1829 8265 1835
rect 8315 1859 8364 1871
rect 8315 1839 8333 1859
rect 8353 1839 8364 1859
rect 8315 1829 8364 1839
rect 8434 1855 8478 1871
rect 8434 1835 8443 1855
rect 8463 1835 8478 1855
rect 8434 1829 8478 1835
rect 8528 1859 8577 1871
rect 8528 1839 8546 1859
rect 8566 1839 8577 1859
rect 8528 1829 8577 1839
rect 18909 2131 18958 2143
rect 18909 2111 18920 2131
rect 18940 2111 18958 2131
rect 18909 2101 18958 2111
rect 19008 2127 19052 2143
rect 19008 2107 19023 2127
rect 19043 2107 19052 2127
rect 19008 2101 19052 2107
rect 19122 2127 19166 2143
rect 19122 2107 19131 2127
rect 19151 2107 19166 2127
rect 19122 2101 19166 2107
rect 19216 2131 19265 2143
rect 19216 2111 19234 2131
rect 19254 2111 19265 2131
rect 19216 2101 19265 2111
rect 19330 2127 19374 2143
rect 19330 2107 19339 2127
rect 19359 2107 19374 2127
rect 19330 2101 19374 2107
rect 19424 2131 19473 2143
rect 19424 2111 19442 2131
rect 19462 2111 19473 2131
rect 19424 2101 19473 2111
rect 19543 2127 19587 2143
rect 19543 2107 19552 2127
rect 19572 2107 19587 2127
rect 19543 2101 19587 2107
rect 19637 2131 19686 2143
rect 19637 2111 19655 2131
rect 19675 2111 19686 2131
rect 19637 2101 19686 2111
rect 15422 1893 15471 1903
rect 15422 1873 15433 1893
rect 15453 1873 15471 1893
rect 10366 1852 10415 1862
rect 10366 1832 10377 1852
rect 10397 1832 10415 1852
rect 10366 1820 10415 1832
rect 10465 1856 10509 1862
rect 10465 1836 10480 1856
rect 10500 1836 10509 1856
rect 10465 1820 10509 1836
rect 10579 1852 10628 1862
rect 10579 1832 10590 1852
rect 10610 1832 10628 1852
rect 10579 1820 10628 1832
rect 10678 1856 10722 1862
rect 10678 1836 10693 1856
rect 10713 1836 10722 1856
rect 10678 1820 10722 1836
rect 10787 1852 10836 1862
rect 10787 1832 10798 1852
rect 10818 1832 10836 1852
rect 10787 1820 10836 1832
rect 10886 1856 10930 1862
rect 10886 1836 10901 1856
rect 10921 1836 10930 1856
rect 10886 1820 10930 1836
rect 11000 1856 11044 1862
rect 11000 1836 11009 1856
rect 11029 1836 11044 1856
rect 11000 1820 11044 1836
rect 11094 1852 11143 1862
rect 11094 1832 11112 1852
rect 11132 1832 11143 1852
rect 11094 1820 11143 1832
rect 12775 1823 12824 1835
rect 12775 1803 12786 1823
rect 12806 1803 12824 1823
rect 12775 1793 12824 1803
rect 12874 1819 12918 1835
rect 12874 1799 12889 1819
rect 12909 1799 12918 1819
rect 12874 1793 12918 1799
rect 12988 1819 13032 1835
rect 12988 1799 12997 1819
rect 13017 1799 13032 1819
rect 12988 1793 13032 1799
rect 13082 1823 13131 1835
rect 13082 1803 13100 1823
rect 13120 1803 13131 1823
rect 13082 1793 13131 1803
rect 13196 1819 13240 1835
rect 13196 1799 13205 1819
rect 13225 1799 13240 1819
rect 13196 1793 13240 1799
rect 13290 1823 13339 1835
rect 13290 1803 13308 1823
rect 13328 1803 13339 1823
rect 13290 1793 13339 1803
rect 13409 1819 13453 1835
rect 13409 1799 13418 1819
rect 13438 1799 13453 1819
rect 13409 1793 13453 1799
rect 13503 1823 13552 1835
rect 13503 1803 13521 1823
rect 13541 1803 13552 1823
rect 13503 1793 13552 1803
rect 15422 1861 15471 1873
rect 15521 1897 15565 1903
rect 15521 1877 15536 1897
rect 15556 1877 15565 1897
rect 15521 1861 15565 1877
rect 15635 1893 15684 1903
rect 15635 1873 15646 1893
rect 15666 1873 15684 1893
rect 15635 1861 15684 1873
rect 15734 1897 15778 1903
rect 15734 1877 15749 1897
rect 15769 1877 15778 1897
rect 15734 1861 15778 1877
rect 15843 1893 15892 1903
rect 15843 1873 15854 1893
rect 15874 1873 15892 1893
rect 15843 1861 15892 1873
rect 15942 1897 15986 1903
rect 15942 1877 15957 1897
rect 15977 1877 15986 1897
rect 15942 1861 15986 1877
rect 16056 1897 16100 1903
rect 16056 1877 16065 1897
rect 16085 1877 16100 1897
rect 16056 1861 16100 1877
rect 16150 1893 16199 1903
rect 16150 1873 16168 1893
rect 16188 1873 16199 1893
rect 16150 1861 16199 1873
rect 17831 1864 17880 1876
rect 17831 1844 17842 1864
rect 17862 1844 17880 1864
rect 17831 1834 17880 1844
rect 17930 1860 17974 1876
rect 17930 1840 17945 1860
rect 17965 1840 17974 1860
rect 17930 1834 17974 1840
rect 18044 1860 18088 1876
rect 18044 1840 18053 1860
rect 18073 1840 18088 1860
rect 18044 1834 18088 1840
rect 18138 1864 18187 1876
rect 18138 1844 18156 1864
rect 18176 1844 18187 1864
rect 18138 1834 18187 1844
rect 18252 1860 18296 1876
rect 18252 1840 18261 1860
rect 18281 1840 18296 1860
rect 18252 1834 18296 1840
rect 18346 1864 18395 1876
rect 18346 1844 18364 1864
rect 18384 1844 18395 1864
rect 18346 1834 18395 1844
rect 18465 1860 18509 1876
rect 18465 1840 18474 1860
rect 18494 1840 18509 1860
rect 18465 1834 18509 1840
rect 18559 1864 18608 1876
rect 18559 1844 18577 1864
rect 18597 1844 18608 1864
rect 18559 1834 18608 1844
rect 1415 1565 1464 1575
rect 1415 1545 1426 1565
rect 1446 1545 1464 1565
rect 1415 1533 1464 1545
rect 1514 1569 1558 1575
rect 1514 1549 1529 1569
rect 1549 1549 1558 1569
rect 1514 1533 1558 1549
rect 1628 1565 1677 1575
rect 1628 1545 1639 1565
rect 1659 1545 1677 1565
rect 1628 1533 1677 1545
rect 1727 1569 1771 1575
rect 1727 1549 1742 1569
rect 1762 1549 1771 1569
rect 1727 1533 1771 1549
rect 1836 1565 1885 1575
rect 1836 1545 1847 1565
rect 1867 1545 1885 1565
rect 1836 1533 1885 1545
rect 1935 1569 1979 1575
rect 1935 1549 1950 1569
rect 1970 1549 1979 1569
rect 1935 1533 1979 1549
rect 2049 1569 2093 1575
rect 2049 1549 2058 1569
rect 2078 1549 2093 1569
rect 2049 1533 2093 1549
rect 2143 1565 2192 1575
rect 2143 1545 2161 1565
rect 2181 1545 2192 1565
rect 2143 1533 2192 1545
rect 3824 1536 3873 1548
rect 3824 1516 3835 1536
rect 3855 1516 3873 1536
rect 3824 1506 3873 1516
rect 3923 1532 3967 1548
rect 3923 1512 3938 1532
rect 3958 1512 3967 1532
rect 3923 1506 3967 1512
rect 4037 1532 4081 1548
rect 4037 1512 4046 1532
rect 4066 1512 4081 1532
rect 4037 1506 4081 1512
rect 4131 1536 4180 1548
rect 4131 1516 4149 1536
rect 4169 1516 4180 1536
rect 4131 1506 4180 1516
rect 4245 1532 4289 1548
rect 4245 1512 4254 1532
rect 4274 1512 4289 1532
rect 4245 1506 4289 1512
rect 4339 1536 4388 1548
rect 4339 1516 4357 1536
rect 4377 1516 4388 1536
rect 4339 1506 4388 1516
rect 4458 1532 4502 1548
rect 4458 1512 4467 1532
rect 4487 1512 4502 1532
rect 4458 1506 4502 1512
rect 4552 1536 4601 1548
rect 6471 1606 6520 1616
rect 6471 1586 6482 1606
rect 6502 1586 6520 1606
rect 6471 1574 6520 1586
rect 6570 1610 6614 1616
rect 6570 1590 6585 1610
rect 6605 1590 6614 1610
rect 6570 1574 6614 1590
rect 6684 1606 6733 1616
rect 6684 1586 6695 1606
rect 6715 1586 6733 1606
rect 6684 1574 6733 1586
rect 6783 1610 6827 1616
rect 6783 1590 6798 1610
rect 6818 1590 6827 1610
rect 6783 1574 6827 1590
rect 6892 1606 6941 1616
rect 6892 1586 6903 1606
rect 6923 1586 6941 1606
rect 6892 1574 6941 1586
rect 6991 1610 7035 1616
rect 6991 1590 7006 1610
rect 7026 1590 7035 1610
rect 6991 1574 7035 1590
rect 7105 1610 7149 1616
rect 7105 1590 7114 1610
rect 7134 1590 7149 1610
rect 7105 1574 7149 1590
rect 7199 1606 7248 1616
rect 7199 1586 7217 1606
rect 7237 1586 7248 1606
rect 7199 1574 7248 1586
rect 8880 1577 8929 1589
rect 8880 1557 8891 1577
rect 8911 1557 8929 1577
rect 8880 1547 8929 1557
rect 8979 1573 9023 1589
rect 8979 1553 8994 1573
rect 9014 1553 9023 1573
rect 8979 1547 9023 1553
rect 9093 1573 9137 1589
rect 9093 1553 9102 1573
rect 9122 1553 9137 1573
rect 9093 1547 9137 1553
rect 9187 1577 9236 1589
rect 9187 1557 9205 1577
rect 9225 1557 9236 1577
rect 9187 1547 9236 1557
rect 9301 1573 9345 1589
rect 9301 1553 9310 1573
rect 9330 1553 9345 1573
rect 9301 1547 9345 1553
rect 9395 1577 9444 1589
rect 9395 1557 9413 1577
rect 9433 1557 9444 1577
rect 9395 1547 9444 1557
rect 9514 1573 9558 1589
rect 9514 1553 9523 1573
rect 9543 1553 9558 1573
rect 9514 1547 9558 1553
rect 9608 1577 9657 1589
rect 9608 1557 9626 1577
rect 9646 1557 9657 1577
rect 9608 1547 9657 1557
rect 4552 1516 4570 1536
rect 4590 1516 4601 1536
rect 4552 1506 4601 1516
rect 337 1298 386 1308
rect 337 1278 348 1298
rect 368 1278 386 1298
rect 337 1266 386 1278
rect 436 1302 480 1308
rect 436 1282 451 1302
rect 471 1282 480 1302
rect 436 1266 480 1282
rect 550 1298 599 1308
rect 550 1278 561 1298
rect 581 1278 599 1298
rect 550 1266 599 1278
rect 649 1302 693 1308
rect 649 1282 664 1302
rect 684 1282 693 1302
rect 649 1266 693 1282
rect 758 1298 807 1308
rect 758 1278 769 1298
rect 789 1278 807 1298
rect 758 1266 807 1278
rect 857 1302 901 1308
rect 857 1282 872 1302
rect 892 1282 901 1302
rect 857 1266 901 1282
rect 971 1302 1015 1308
rect 971 1282 980 1302
rect 1000 1282 1015 1302
rect 971 1266 1015 1282
rect 1065 1298 1114 1308
rect 1065 1278 1083 1298
rect 1103 1278 1114 1298
rect 1065 1266 1114 1278
rect 11446 1570 11495 1580
rect 11446 1550 11457 1570
rect 11477 1550 11495 1570
rect 11446 1538 11495 1550
rect 11545 1574 11589 1580
rect 11545 1554 11560 1574
rect 11580 1554 11589 1574
rect 11545 1538 11589 1554
rect 11659 1570 11708 1580
rect 11659 1550 11670 1570
rect 11690 1550 11708 1570
rect 11659 1538 11708 1550
rect 11758 1574 11802 1580
rect 11758 1554 11773 1574
rect 11793 1554 11802 1574
rect 11758 1538 11802 1554
rect 11867 1570 11916 1580
rect 11867 1550 11878 1570
rect 11898 1550 11916 1570
rect 11867 1538 11916 1550
rect 11966 1574 12010 1580
rect 11966 1554 11981 1574
rect 12001 1554 12010 1574
rect 11966 1538 12010 1554
rect 12080 1574 12124 1580
rect 12080 1554 12089 1574
rect 12109 1554 12124 1574
rect 12080 1538 12124 1554
rect 12174 1570 12223 1580
rect 12174 1550 12192 1570
rect 12212 1550 12223 1570
rect 12174 1538 12223 1550
rect 13855 1541 13904 1553
rect 13855 1521 13866 1541
rect 13886 1521 13904 1541
rect 13855 1511 13904 1521
rect 13954 1537 13998 1553
rect 13954 1517 13969 1537
rect 13989 1517 13998 1537
rect 13954 1511 13998 1517
rect 14068 1537 14112 1553
rect 14068 1517 14077 1537
rect 14097 1517 14112 1537
rect 14068 1511 14112 1517
rect 14162 1541 14211 1553
rect 14162 1521 14180 1541
rect 14200 1521 14211 1541
rect 14162 1511 14211 1521
rect 14276 1537 14320 1553
rect 14276 1517 14285 1537
rect 14305 1517 14320 1537
rect 14276 1511 14320 1517
rect 14370 1541 14419 1553
rect 14370 1521 14388 1541
rect 14408 1521 14419 1541
rect 14370 1511 14419 1521
rect 14489 1537 14533 1553
rect 14489 1517 14498 1537
rect 14518 1517 14533 1537
rect 14489 1511 14533 1517
rect 14583 1541 14632 1553
rect 16502 1611 16551 1621
rect 16502 1591 16513 1611
rect 16533 1591 16551 1611
rect 16502 1579 16551 1591
rect 16601 1615 16645 1621
rect 16601 1595 16616 1615
rect 16636 1595 16645 1615
rect 16601 1579 16645 1595
rect 16715 1611 16764 1621
rect 16715 1591 16726 1611
rect 16746 1591 16764 1611
rect 16715 1579 16764 1591
rect 16814 1615 16858 1621
rect 16814 1595 16829 1615
rect 16849 1595 16858 1615
rect 16814 1579 16858 1595
rect 16923 1611 16972 1621
rect 16923 1591 16934 1611
rect 16954 1591 16972 1611
rect 16923 1579 16972 1591
rect 17022 1615 17066 1621
rect 17022 1595 17037 1615
rect 17057 1595 17066 1615
rect 17022 1579 17066 1595
rect 17136 1615 17180 1621
rect 17136 1595 17145 1615
rect 17165 1595 17180 1615
rect 17136 1579 17180 1595
rect 17230 1611 17279 1621
rect 17230 1591 17248 1611
rect 17268 1591 17279 1611
rect 17230 1579 17279 1591
rect 18911 1582 18960 1594
rect 18911 1562 18922 1582
rect 18942 1562 18960 1582
rect 18911 1552 18960 1562
rect 19010 1578 19054 1594
rect 19010 1558 19025 1578
rect 19045 1558 19054 1578
rect 19010 1552 19054 1558
rect 19124 1578 19168 1594
rect 19124 1558 19133 1578
rect 19153 1558 19168 1578
rect 19124 1552 19168 1558
rect 19218 1582 19267 1594
rect 19218 1562 19236 1582
rect 19256 1562 19267 1582
rect 19218 1552 19267 1562
rect 19332 1578 19376 1594
rect 19332 1558 19341 1578
rect 19361 1558 19376 1578
rect 19332 1552 19376 1558
rect 19426 1582 19475 1594
rect 19426 1562 19444 1582
rect 19464 1562 19475 1582
rect 19426 1552 19475 1562
rect 19545 1578 19589 1594
rect 19545 1558 19554 1578
rect 19574 1558 19589 1578
rect 19545 1552 19589 1558
rect 19639 1582 19688 1594
rect 19639 1562 19657 1582
rect 19677 1562 19688 1582
rect 19639 1552 19688 1562
rect 14583 1521 14601 1541
rect 14621 1521 14632 1541
rect 14583 1511 14632 1521
rect 5393 1339 5442 1349
rect 5393 1319 5404 1339
rect 5424 1319 5442 1339
rect 5393 1307 5442 1319
rect 5492 1343 5536 1349
rect 5492 1323 5507 1343
rect 5527 1323 5536 1343
rect 5492 1307 5536 1323
rect 5606 1339 5655 1349
rect 5606 1319 5617 1339
rect 5637 1319 5655 1339
rect 5606 1307 5655 1319
rect 5705 1343 5749 1349
rect 5705 1323 5720 1343
rect 5740 1323 5749 1343
rect 5705 1307 5749 1323
rect 5814 1339 5863 1349
rect 5814 1319 5825 1339
rect 5845 1319 5863 1339
rect 5814 1307 5863 1319
rect 5913 1343 5957 1349
rect 5913 1323 5928 1343
rect 5948 1323 5957 1343
rect 5913 1307 5957 1323
rect 6027 1343 6071 1349
rect 6027 1323 6036 1343
rect 6056 1323 6071 1343
rect 6027 1307 6071 1323
rect 6121 1339 6170 1349
rect 6121 1319 6139 1339
rect 6159 1319 6170 1339
rect 6121 1307 6170 1319
rect 2885 1226 2934 1238
rect 2885 1206 2896 1226
rect 2916 1206 2934 1226
rect 2885 1196 2934 1206
rect 2984 1222 3028 1238
rect 2984 1202 2999 1222
rect 3019 1202 3028 1222
rect 2984 1196 3028 1202
rect 3098 1222 3142 1238
rect 3098 1202 3107 1222
rect 3127 1202 3142 1222
rect 3098 1196 3142 1202
rect 3192 1226 3241 1238
rect 3192 1206 3210 1226
rect 3230 1206 3241 1226
rect 3192 1196 3241 1206
rect 3306 1222 3350 1238
rect 3306 1202 3315 1222
rect 3335 1202 3350 1222
rect 3306 1196 3350 1202
rect 3400 1226 3449 1238
rect 3400 1206 3418 1226
rect 3438 1206 3449 1226
rect 3400 1196 3449 1206
rect 3519 1222 3563 1238
rect 3519 1202 3528 1222
rect 3548 1202 3563 1222
rect 3519 1196 3563 1202
rect 3613 1226 3662 1238
rect 3613 1206 3631 1226
rect 3651 1206 3662 1226
rect 3613 1196 3662 1206
rect 1275 1054 1324 1064
rect 1275 1034 1286 1054
rect 1306 1034 1324 1054
rect 1275 1022 1324 1034
rect 1374 1058 1418 1064
rect 1374 1038 1389 1058
rect 1409 1038 1418 1058
rect 1374 1022 1418 1038
rect 1488 1054 1537 1064
rect 1488 1034 1499 1054
rect 1519 1034 1537 1054
rect 1488 1022 1537 1034
rect 1587 1058 1631 1064
rect 1587 1038 1602 1058
rect 1622 1038 1631 1058
rect 1587 1022 1631 1038
rect 1696 1054 1745 1064
rect 1696 1034 1707 1054
rect 1727 1034 1745 1054
rect 1696 1022 1745 1034
rect 1795 1058 1839 1064
rect 1795 1038 1810 1058
rect 1830 1038 1839 1058
rect 1795 1022 1839 1038
rect 1909 1058 1953 1064
rect 1909 1038 1918 1058
rect 1938 1038 1953 1058
rect 1909 1022 1953 1038
rect 2003 1054 2052 1064
rect 2003 1034 2021 1054
rect 2041 1034 2052 1054
rect 2003 1022 2052 1034
rect 7941 1267 7990 1279
rect 7941 1247 7952 1267
rect 7972 1247 7990 1267
rect 7941 1237 7990 1247
rect 8040 1263 8084 1279
rect 8040 1243 8055 1263
rect 8075 1243 8084 1263
rect 8040 1237 8084 1243
rect 8154 1263 8198 1279
rect 8154 1243 8163 1263
rect 8183 1243 8198 1263
rect 8154 1237 8198 1243
rect 8248 1267 8297 1279
rect 8248 1247 8266 1267
rect 8286 1247 8297 1267
rect 8248 1237 8297 1247
rect 8362 1263 8406 1279
rect 8362 1243 8371 1263
rect 8391 1243 8406 1263
rect 8362 1237 8406 1243
rect 8456 1267 8505 1279
rect 8456 1247 8474 1267
rect 8494 1247 8505 1267
rect 8456 1237 8505 1247
rect 8575 1263 8619 1279
rect 8575 1243 8584 1263
rect 8604 1243 8619 1263
rect 8575 1237 8619 1243
rect 8669 1267 8718 1279
rect 8669 1247 8687 1267
rect 8707 1247 8718 1267
rect 8669 1237 8718 1247
rect 10368 1303 10417 1313
rect 10368 1283 10379 1303
rect 10399 1283 10417 1303
rect 10368 1271 10417 1283
rect 10467 1307 10511 1313
rect 10467 1287 10482 1307
rect 10502 1287 10511 1307
rect 10467 1271 10511 1287
rect 10581 1303 10630 1313
rect 10581 1283 10592 1303
rect 10612 1283 10630 1303
rect 10581 1271 10630 1283
rect 10680 1307 10724 1313
rect 10680 1287 10695 1307
rect 10715 1287 10724 1307
rect 10680 1271 10724 1287
rect 10789 1303 10838 1313
rect 10789 1283 10800 1303
rect 10820 1283 10838 1303
rect 10789 1271 10838 1283
rect 10888 1307 10932 1313
rect 10888 1287 10903 1307
rect 10923 1287 10932 1307
rect 10888 1271 10932 1287
rect 11002 1307 11046 1313
rect 11002 1287 11011 1307
rect 11031 1287 11046 1307
rect 11002 1271 11046 1287
rect 11096 1303 11145 1313
rect 11096 1283 11114 1303
rect 11134 1283 11145 1303
rect 11096 1271 11145 1283
rect 15424 1344 15473 1354
rect 15424 1324 15435 1344
rect 15455 1324 15473 1344
rect 15424 1312 15473 1324
rect 15523 1348 15567 1354
rect 15523 1328 15538 1348
rect 15558 1328 15567 1348
rect 15523 1312 15567 1328
rect 15637 1344 15686 1354
rect 15637 1324 15648 1344
rect 15668 1324 15686 1344
rect 15637 1312 15686 1324
rect 15736 1348 15780 1354
rect 15736 1328 15751 1348
rect 15771 1328 15780 1348
rect 15736 1312 15780 1328
rect 15845 1344 15894 1354
rect 15845 1324 15856 1344
rect 15876 1324 15894 1344
rect 15845 1312 15894 1324
rect 15944 1348 15988 1354
rect 15944 1328 15959 1348
rect 15979 1328 15988 1348
rect 15944 1312 15988 1328
rect 16058 1348 16102 1354
rect 16058 1328 16067 1348
rect 16087 1328 16102 1348
rect 16058 1312 16102 1328
rect 16152 1344 16201 1354
rect 16152 1324 16170 1344
rect 16190 1324 16201 1344
rect 16152 1312 16201 1324
rect 6331 1095 6380 1105
rect 6331 1075 6342 1095
rect 6362 1075 6380 1095
rect 6331 1063 6380 1075
rect 6430 1099 6474 1105
rect 6430 1079 6445 1099
rect 6465 1079 6474 1099
rect 6430 1063 6474 1079
rect 6544 1095 6593 1105
rect 6544 1075 6555 1095
rect 6575 1075 6593 1095
rect 6544 1063 6593 1075
rect 6643 1099 6687 1105
rect 6643 1079 6658 1099
rect 6678 1079 6687 1099
rect 6643 1063 6687 1079
rect 6752 1095 6801 1105
rect 6752 1075 6763 1095
rect 6783 1075 6801 1095
rect 6752 1063 6801 1075
rect 6851 1099 6895 1105
rect 6851 1079 6866 1099
rect 6886 1079 6895 1099
rect 6851 1063 6895 1079
rect 6965 1099 7009 1105
rect 6965 1079 6974 1099
rect 6994 1079 7009 1099
rect 6965 1063 7009 1079
rect 7059 1095 7108 1105
rect 7059 1075 7077 1095
rect 7097 1075 7108 1095
rect 7059 1063 7108 1075
rect 12916 1231 12965 1243
rect 12916 1211 12927 1231
rect 12947 1211 12965 1231
rect 12916 1201 12965 1211
rect 13015 1227 13059 1243
rect 13015 1207 13030 1227
rect 13050 1207 13059 1227
rect 13015 1201 13059 1207
rect 13129 1227 13173 1243
rect 13129 1207 13138 1227
rect 13158 1207 13173 1227
rect 13129 1201 13173 1207
rect 13223 1231 13272 1243
rect 13223 1211 13241 1231
rect 13261 1211 13272 1231
rect 13223 1201 13272 1211
rect 13337 1227 13381 1243
rect 13337 1207 13346 1227
rect 13366 1207 13381 1227
rect 13337 1201 13381 1207
rect 13431 1231 13480 1243
rect 13431 1211 13449 1231
rect 13469 1211 13480 1231
rect 13431 1201 13480 1211
rect 13550 1227 13594 1243
rect 13550 1207 13559 1227
rect 13579 1207 13594 1227
rect 13550 1201 13594 1207
rect 13644 1231 13693 1243
rect 13644 1211 13662 1231
rect 13682 1211 13693 1231
rect 13644 1201 13693 1211
rect 3823 982 3872 994
rect 3823 962 3834 982
rect 3854 962 3872 982
rect 3823 952 3872 962
rect 3922 978 3966 994
rect 3922 958 3937 978
rect 3957 958 3966 978
rect 3922 952 3966 958
rect 4036 978 4080 994
rect 4036 958 4045 978
rect 4065 958 4080 978
rect 4036 952 4080 958
rect 4130 982 4179 994
rect 4130 962 4148 982
rect 4168 962 4179 982
rect 4130 952 4179 962
rect 4244 978 4288 994
rect 4244 958 4253 978
rect 4273 958 4288 978
rect 4244 952 4288 958
rect 4338 982 4387 994
rect 4338 962 4356 982
rect 4376 962 4387 982
rect 4338 952 4387 962
rect 4457 978 4501 994
rect 4457 958 4466 978
rect 4486 958 4501 978
rect 4457 952 4501 958
rect 4551 982 4600 994
rect 4551 962 4569 982
rect 4589 962 4600 982
rect 4551 952 4600 962
rect 8879 1023 8928 1035
rect 8879 1003 8890 1023
rect 8910 1003 8928 1023
rect 8879 993 8928 1003
rect 8978 1019 9022 1035
rect 8978 999 8993 1019
rect 9013 999 9022 1019
rect 8978 993 9022 999
rect 9092 1019 9136 1035
rect 9092 999 9101 1019
rect 9121 999 9136 1019
rect 9092 993 9136 999
rect 9186 1023 9235 1035
rect 9186 1003 9204 1023
rect 9224 1003 9235 1023
rect 9186 993 9235 1003
rect 9300 1019 9344 1035
rect 9300 999 9309 1019
rect 9329 999 9344 1019
rect 9300 993 9344 999
rect 9394 1023 9443 1035
rect 9394 1003 9412 1023
rect 9432 1003 9443 1023
rect 9394 993 9443 1003
rect 9513 1019 9557 1035
rect 9513 999 9522 1019
rect 9542 999 9557 1019
rect 9513 993 9557 999
rect 9607 1023 9656 1035
rect 9607 1003 9625 1023
rect 9645 1003 9656 1023
rect 9607 993 9656 1003
rect 11306 1059 11355 1069
rect 11306 1039 11317 1059
rect 11337 1039 11355 1059
rect 11306 1027 11355 1039
rect 11405 1063 11449 1069
rect 11405 1043 11420 1063
rect 11440 1043 11449 1063
rect 11405 1027 11449 1043
rect 11519 1059 11568 1069
rect 11519 1039 11530 1059
rect 11550 1039 11568 1059
rect 11519 1027 11568 1039
rect 11618 1063 11662 1069
rect 11618 1043 11633 1063
rect 11653 1043 11662 1063
rect 11618 1027 11662 1043
rect 11727 1059 11776 1069
rect 11727 1039 11738 1059
rect 11758 1039 11776 1059
rect 11727 1027 11776 1039
rect 11826 1063 11870 1069
rect 11826 1043 11841 1063
rect 11861 1043 11870 1063
rect 11826 1027 11870 1043
rect 11940 1063 11984 1069
rect 11940 1043 11949 1063
rect 11969 1043 11984 1063
rect 11940 1027 11984 1043
rect 12034 1059 12083 1069
rect 12034 1039 12052 1059
rect 12072 1039 12083 1059
rect 12034 1027 12083 1039
rect 17972 1272 18021 1284
rect 17972 1252 17983 1272
rect 18003 1252 18021 1272
rect 17972 1242 18021 1252
rect 18071 1268 18115 1284
rect 18071 1248 18086 1268
rect 18106 1248 18115 1268
rect 18071 1242 18115 1248
rect 18185 1268 18229 1284
rect 18185 1248 18194 1268
rect 18214 1248 18229 1268
rect 18185 1242 18229 1248
rect 18279 1272 18328 1284
rect 18279 1252 18297 1272
rect 18317 1252 18328 1272
rect 18279 1242 18328 1252
rect 18393 1268 18437 1284
rect 18393 1248 18402 1268
rect 18422 1248 18437 1268
rect 18393 1242 18437 1248
rect 18487 1272 18536 1284
rect 18487 1252 18505 1272
rect 18525 1252 18536 1272
rect 18487 1242 18536 1252
rect 18606 1268 18650 1284
rect 18606 1248 18615 1268
rect 18635 1248 18650 1268
rect 18606 1242 18650 1248
rect 18700 1272 18749 1284
rect 18700 1252 18718 1272
rect 18738 1252 18749 1272
rect 18700 1242 18749 1252
rect 16362 1100 16411 1110
rect 16362 1080 16373 1100
rect 16393 1080 16411 1100
rect 16362 1068 16411 1080
rect 16461 1104 16505 1110
rect 16461 1084 16476 1104
rect 16496 1084 16505 1104
rect 16461 1068 16505 1084
rect 16575 1100 16624 1110
rect 16575 1080 16586 1100
rect 16606 1080 16624 1100
rect 16575 1068 16624 1080
rect 16674 1104 16718 1110
rect 16674 1084 16689 1104
rect 16709 1084 16718 1104
rect 16674 1068 16718 1084
rect 16783 1100 16832 1110
rect 16783 1080 16794 1100
rect 16814 1080 16832 1100
rect 16783 1068 16832 1080
rect 16882 1104 16926 1110
rect 16882 1084 16897 1104
rect 16917 1084 16926 1104
rect 16882 1068 16926 1084
rect 16996 1104 17040 1110
rect 16996 1084 17005 1104
rect 17025 1084 17040 1104
rect 16996 1068 17040 1084
rect 17090 1100 17139 1110
rect 17090 1080 17108 1100
rect 17128 1080 17139 1100
rect 17090 1068 17139 1080
rect 13854 987 13903 999
rect 13854 967 13865 987
rect 13885 967 13903 987
rect 13854 957 13903 967
rect 13953 983 13997 999
rect 13953 963 13968 983
rect 13988 963 13997 983
rect 13953 957 13997 963
rect 14067 983 14111 999
rect 14067 963 14076 983
rect 14096 963 14111 983
rect 14067 957 14111 963
rect 14161 987 14210 999
rect 14161 967 14179 987
rect 14199 967 14210 987
rect 14161 957 14210 967
rect 14275 983 14319 999
rect 14275 963 14284 983
rect 14304 963 14319 983
rect 14275 957 14319 963
rect 14369 987 14418 999
rect 14369 967 14387 987
rect 14407 967 14418 987
rect 14369 957 14418 967
rect 14488 983 14532 999
rect 14488 963 14497 983
rect 14517 963 14532 983
rect 14488 957 14532 963
rect 14582 987 14631 999
rect 14582 967 14600 987
rect 14620 967 14631 987
rect 14582 957 14631 967
rect 5392 785 5441 795
rect 5392 765 5403 785
rect 5423 765 5441 785
rect 336 744 385 754
rect 336 724 347 744
rect 367 724 385 744
rect 336 712 385 724
rect 435 748 479 754
rect 435 728 450 748
rect 470 728 479 748
rect 435 712 479 728
rect 549 744 598 754
rect 549 724 560 744
rect 580 724 598 744
rect 549 712 598 724
rect 648 748 692 754
rect 648 728 663 748
rect 683 728 692 748
rect 648 712 692 728
rect 757 744 806 754
rect 757 724 768 744
rect 788 724 806 744
rect 757 712 806 724
rect 856 748 900 754
rect 856 728 871 748
rect 891 728 900 748
rect 856 712 900 728
rect 970 748 1014 754
rect 970 728 979 748
rect 999 728 1014 748
rect 970 712 1014 728
rect 1064 744 1113 754
rect 1064 724 1082 744
rect 1102 724 1113 744
rect 1064 712 1113 724
rect 5392 753 5441 765
rect 5491 789 5535 795
rect 5491 769 5506 789
rect 5526 769 5535 789
rect 5491 753 5535 769
rect 5605 785 5654 795
rect 5605 765 5616 785
rect 5636 765 5654 785
rect 5605 753 5654 765
rect 5704 789 5748 795
rect 5704 769 5719 789
rect 5739 769 5748 789
rect 5704 753 5748 769
rect 5813 785 5862 795
rect 5813 765 5824 785
rect 5844 765 5862 785
rect 5813 753 5862 765
rect 5912 789 5956 795
rect 5912 769 5927 789
rect 5947 769 5956 789
rect 5912 753 5956 769
rect 6026 789 6070 795
rect 6026 769 6035 789
rect 6055 769 6070 789
rect 6026 753 6070 769
rect 6120 785 6169 795
rect 6120 765 6138 785
rect 6158 765 6169 785
rect 6120 753 6169 765
rect 18910 1028 18959 1040
rect 18910 1008 18921 1028
rect 18941 1008 18959 1028
rect 18910 998 18959 1008
rect 19009 1024 19053 1040
rect 19009 1004 19024 1024
rect 19044 1004 19053 1024
rect 19009 998 19053 1004
rect 19123 1024 19167 1040
rect 19123 1004 19132 1024
rect 19152 1004 19167 1024
rect 19123 998 19167 1004
rect 19217 1028 19266 1040
rect 19217 1008 19235 1028
rect 19255 1008 19266 1028
rect 19217 998 19266 1008
rect 19331 1024 19375 1040
rect 19331 1004 19340 1024
rect 19360 1004 19375 1024
rect 19331 998 19375 1004
rect 19425 1028 19474 1040
rect 19425 1008 19443 1028
rect 19463 1008 19474 1028
rect 19425 998 19474 1008
rect 19544 1024 19588 1040
rect 19544 1004 19553 1024
rect 19573 1004 19588 1024
rect 19544 998 19588 1004
rect 19638 1028 19687 1040
rect 19638 1008 19656 1028
rect 19676 1008 19687 1028
rect 19638 998 19687 1008
rect 15423 790 15472 800
rect 15423 770 15434 790
rect 15454 770 15472 790
rect 10367 749 10416 759
rect 10367 729 10378 749
rect 10398 729 10416 749
rect 10367 717 10416 729
rect 10466 753 10510 759
rect 10466 733 10481 753
rect 10501 733 10510 753
rect 10466 717 10510 733
rect 10580 749 10629 759
rect 10580 729 10591 749
rect 10611 729 10629 749
rect 10580 717 10629 729
rect 10679 753 10723 759
rect 10679 733 10694 753
rect 10714 733 10723 753
rect 10679 717 10723 733
rect 10788 749 10837 759
rect 10788 729 10799 749
rect 10819 729 10837 749
rect 10788 717 10837 729
rect 10887 753 10931 759
rect 10887 733 10902 753
rect 10922 733 10931 753
rect 10887 717 10931 733
rect 11001 753 11045 759
rect 11001 733 11010 753
rect 11030 733 11045 753
rect 11001 717 11045 733
rect 11095 749 11144 759
rect 11095 729 11113 749
rect 11133 729 11144 749
rect 11095 717 11144 729
rect 15423 758 15472 770
rect 15522 794 15566 800
rect 15522 774 15537 794
rect 15557 774 15566 794
rect 15522 758 15566 774
rect 15636 790 15685 800
rect 15636 770 15647 790
rect 15667 770 15685 790
rect 15636 758 15685 770
rect 15735 794 15779 800
rect 15735 774 15750 794
rect 15770 774 15779 794
rect 15735 758 15779 774
rect 15844 790 15893 800
rect 15844 770 15855 790
rect 15875 770 15893 790
rect 15844 758 15893 770
rect 15943 794 15987 800
rect 15943 774 15958 794
rect 15978 774 15987 794
rect 15943 758 15987 774
rect 16057 794 16101 800
rect 16057 774 16066 794
rect 16086 774 16101 794
rect 16057 758 16101 774
rect 16151 790 16200 800
rect 16151 770 16169 790
rect 16189 770 16200 790
rect 16151 758 16200 770
rect 1583 185 1632 195
rect 1583 165 1594 185
rect 1614 165 1632 185
rect 1583 153 1632 165
rect 1682 189 1726 195
rect 1682 169 1697 189
rect 1717 169 1726 189
rect 1682 153 1726 169
rect 1796 185 1845 195
rect 1796 165 1807 185
rect 1827 165 1845 185
rect 1796 153 1845 165
rect 1895 189 1939 195
rect 1895 169 1910 189
rect 1930 169 1939 189
rect 1895 153 1939 169
rect 2004 185 2053 195
rect 2004 165 2015 185
rect 2035 165 2053 185
rect 2004 153 2053 165
rect 2103 189 2147 195
rect 2103 169 2118 189
rect 2138 169 2147 189
rect 2103 153 2147 169
rect 2217 189 2261 195
rect 2217 169 2226 189
rect 2246 169 2261 189
rect 2217 153 2261 169
rect 2311 185 2360 195
rect 2311 165 2329 185
rect 2349 165 2360 185
rect 6639 226 6688 236
rect 6639 206 6650 226
rect 6670 206 6688 226
rect 6639 194 6688 206
rect 6738 230 6782 236
rect 6738 210 6753 230
rect 6773 210 6782 230
rect 6738 194 6782 210
rect 6852 226 6901 236
rect 6852 206 6863 226
rect 6883 206 6901 226
rect 6852 194 6901 206
rect 6951 230 6995 236
rect 6951 210 6966 230
rect 6986 210 6995 230
rect 6951 194 6995 210
rect 7060 226 7109 236
rect 7060 206 7071 226
rect 7091 206 7109 226
rect 7060 194 7109 206
rect 7159 230 7203 236
rect 7159 210 7174 230
rect 7194 210 7203 230
rect 7159 194 7203 210
rect 7273 230 7317 236
rect 7273 210 7282 230
rect 7302 210 7317 230
rect 7273 194 7317 210
rect 7367 226 7416 236
rect 7367 206 7385 226
rect 7405 206 7416 226
rect 7367 194 7416 206
rect 2311 153 2360 165
rect 4533 165 4582 175
rect 4533 145 4544 165
rect 4564 145 4582 165
rect 4533 133 4582 145
rect 4632 169 4676 175
rect 4632 149 4647 169
rect 4667 149 4676 169
rect 4632 133 4676 149
rect 4746 165 4795 175
rect 4746 145 4757 165
rect 4777 145 4795 165
rect 4746 133 4795 145
rect 4845 169 4889 175
rect 4845 149 4860 169
rect 4880 149 4889 169
rect 4845 133 4889 149
rect 4954 165 5003 175
rect 4954 145 4965 165
rect 4985 145 5003 165
rect 4954 133 5003 145
rect 5053 169 5097 175
rect 5053 149 5068 169
rect 5088 149 5097 169
rect 5053 133 5097 149
rect 5167 169 5211 175
rect 5167 149 5176 169
rect 5196 149 5211 169
rect 5167 133 5211 149
rect 5261 165 5310 175
rect 5261 145 5279 165
rect 5299 145 5310 165
rect 5261 133 5310 145
rect 11614 190 11663 200
rect 11614 170 11625 190
rect 11645 170 11663 190
rect 11614 158 11663 170
rect 11713 194 11757 200
rect 11713 174 11728 194
rect 11748 174 11757 194
rect 11713 158 11757 174
rect 11827 190 11876 200
rect 11827 170 11838 190
rect 11858 170 11876 190
rect 11827 158 11876 170
rect 11926 194 11970 200
rect 11926 174 11941 194
rect 11961 174 11970 194
rect 11926 158 11970 174
rect 12035 190 12084 200
rect 12035 170 12046 190
rect 12066 170 12084 190
rect 12035 158 12084 170
rect 12134 194 12178 200
rect 12134 174 12149 194
rect 12169 174 12178 194
rect 12134 158 12178 174
rect 12248 194 12292 200
rect 12248 174 12257 194
rect 12277 174 12292 194
rect 12248 158 12292 174
rect 12342 190 12391 200
rect 12342 170 12360 190
rect 12380 170 12391 190
rect 16670 231 16719 241
rect 16670 211 16681 231
rect 16701 211 16719 231
rect 16670 199 16719 211
rect 16769 235 16813 241
rect 16769 215 16784 235
rect 16804 215 16813 235
rect 16769 199 16813 215
rect 16883 231 16932 241
rect 16883 211 16894 231
rect 16914 211 16932 231
rect 16883 199 16932 211
rect 16982 235 17026 241
rect 16982 215 16997 235
rect 17017 215 17026 235
rect 16982 199 17026 215
rect 17091 231 17140 241
rect 17091 211 17102 231
rect 17122 211 17140 231
rect 17091 199 17140 211
rect 17190 235 17234 241
rect 17190 215 17205 235
rect 17225 215 17234 235
rect 17190 199 17234 215
rect 17304 235 17348 241
rect 17304 215 17313 235
rect 17333 215 17348 235
rect 17304 199 17348 215
rect 17398 231 17447 241
rect 17398 211 17416 231
rect 17436 211 17447 231
rect 17398 199 17447 211
rect 12342 158 12391 170
rect 14564 170 14613 180
rect 14564 150 14575 170
rect 14595 150 14613 170
rect 14564 138 14613 150
rect 14663 174 14707 180
rect 14663 154 14678 174
rect 14698 154 14707 174
rect 14663 138 14707 154
rect 14777 170 14826 180
rect 14777 150 14788 170
rect 14808 150 14826 170
rect 14777 138 14826 150
rect 14876 174 14920 180
rect 14876 154 14891 174
rect 14911 154 14920 174
rect 14876 138 14920 154
rect 14985 170 15034 180
rect 14985 150 14996 170
rect 15016 150 15034 170
rect 14985 138 15034 150
rect 15084 174 15128 180
rect 15084 154 15099 174
rect 15119 154 15128 174
rect 15084 138 15128 154
rect 15198 174 15242 180
rect 15198 154 15207 174
rect 15227 154 15242 174
rect 15198 138 15242 154
rect 15292 170 15341 180
rect 15292 150 15310 170
rect 15330 150 15341 170
rect 15292 138 15341 150
rect 9467 49 9516 59
rect 9467 29 9478 49
rect 9498 29 9516 49
rect 9467 17 9516 29
rect 9566 53 9610 59
rect 9566 33 9581 53
rect 9601 33 9610 53
rect 9566 17 9610 33
rect 9680 49 9729 59
rect 9680 29 9691 49
rect 9711 29 9729 49
rect 9680 17 9729 29
rect 9779 53 9823 59
rect 9779 33 9794 53
rect 9814 33 9823 53
rect 9779 17 9823 33
rect 9888 49 9937 59
rect 9888 29 9899 49
rect 9919 29 9937 49
rect 9888 17 9937 29
rect 9987 53 10031 59
rect 9987 33 10002 53
rect 10022 33 10031 53
rect 9987 17 10031 33
rect 10101 53 10145 59
rect 10101 33 10110 53
rect 10130 33 10145 53
rect 10101 17 10145 33
rect 10195 49 10244 59
rect 10195 29 10213 49
rect 10233 29 10244 49
rect 10195 17 10244 29
<< pdiff >>
rect 338 9168 382 9206
rect 338 9148 350 9168
rect 370 9148 382 9168
rect 338 9106 382 9148
rect 432 9168 474 9206
rect 432 9148 446 9168
rect 466 9148 474 9168
rect 432 9106 474 9148
rect 551 9168 595 9206
rect 551 9148 563 9168
rect 583 9148 595 9168
rect 551 9106 595 9148
rect 645 9168 687 9206
rect 645 9148 659 9168
rect 679 9148 687 9168
rect 645 9106 687 9148
rect 759 9168 803 9206
rect 759 9148 771 9168
rect 791 9148 803 9168
rect 759 9106 803 9148
rect 853 9168 895 9206
rect 853 9148 867 9168
rect 887 9148 895 9168
rect 853 9106 895 9148
rect 969 9168 1011 9206
rect 969 9148 977 9168
rect 997 9148 1011 9168
rect 969 9106 1011 9148
rect 1061 9175 1106 9206
rect 1061 9168 1105 9175
rect 1061 9148 1073 9168
rect 1093 9148 1105 9168
rect 5394 9209 5438 9247
rect 5394 9189 5406 9209
rect 5426 9189 5438 9209
rect 1061 9106 1105 9148
rect 3825 9108 3869 9150
rect 3825 9088 3837 9108
rect 3857 9088 3869 9108
rect 3825 9081 3869 9088
rect 3824 9050 3869 9081
rect 3919 9108 3961 9150
rect 3919 9088 3933 9108
rect 3953 9088 3961 9108
rect 3919 9050 3961 9088
rect 4035 9108 4077 9150
rect 4035 9088 4043 9108
rect 4063 9088 4077 9108
rect 4035 9050 4077 9088
rect 4127 9108 4171 9150
rect 4127 9088 4139 9108
rect 4159 9088 4171 9108
rect 4127 9050 4171 9088
rect 4243 9108 4285 9150
rect 4243 9088 4251 9108
rect 4271 9088 4285 9108
rect 4243 9050 4285 9088
rect 4335 9108 4379 9150
rect 4335 9088 4347 9108
rect 4367 9088 4379 9108
rect 4335 9050 4379 9088
rect 4456 9108 4498 9150
rect 4456 9088 4464 9108
rect 4484 9088 4498 9108
rect 4456 9050 4498 9088
rect 4548 9108 4592 9150
rect 5394 9147 5438 9189
rect 5488 9209 5530 9247
rect 5488 9189 5502 9209
rect 5522 9189 5530 9209
rect 5488 9147 5530 9189
rect 5607 9209 5651 9247
rect 5607 9189 5619 9209
rect 5639 9189 5651 9209
rect 5607 9147 5651 9189
rect 5701 9209 5743 9247
rect 5701 9189 5715 9209
rect 5735 9189 5743 9209
rect 5701 9147 5743 9189
rect 5815 9209 5859 9247
rect 5815 9189 5827 9209
rect 5847 9189 5859 9209
rect 5815 9147 5859 9189
rect 5909 9209 5951 9247
rect 5909 9189 5923 9209
rect 5943 9189 5951 9209
rect 5909 9147 5951 9189
rect 6025 9209 6067 9247
rect 6025 9189 6033 9209
rect 6053 9189 6067 9209
rect 6025 9147 6067 9189
rect 6117 9216 6162 9247
rect 6117 9209 6161 9216
rect 6117 9189 6129 9209
rect 6149 9189 6161 9209
rect 6117 9147 6161 9189
rect 8881 9149 8925 9191
rect 4548 9088 4560 9108
rect 4580 9088 4592 9108
rect 4548 9050 4592 9088
rect 8881 9129 8893 9149
rect 8913 9129 8925 9149
rect 8881 9122 8925 9129
rect 8880 9091 8925 9122
rect 8975 9149 9017 9191
rect 8975 9129 8989 9149
rect 9009 9129 9017 9149
rect 8975 9091 9017 9129
rect 9091 9149 9133 9191
rect 9091 9129 9099 9149
rect 9119 9129 9133 9149
rect 9091 9091 9133 9129
rect 9183 9149 9227 9191
rect 9183 9129 9195 9149
rect 9215 9129 9227 9149
rect 9183 9091 9227 9129
rect 9299 9149 9341 9191
rect 9299 9129 9307 9149
rect 9327 9129 9341 9149
rect 9299 9091 9341 9129
rect 9391 9149 9435 9191
rect 9391 9129 9403 9149
rect 9423 9129 9435 9149
rect 9391 9091 9435 9129
rect 9512 9149 9554 9191
rect 9512 9129 9520 9149
rect 9540 9129 9554 9149
rect 9512 9091 9554 9129
rect 9604 9149 9648 9191
rect 10369 9173 10413 9211
rect 9604 9129 9616 9149
rect 9636 9129 9648 9149
rect 9604 9091 9648 9129
rect 10369 9153 10381 9173
rect 10401 9153 10413 9173
rect 10369 9111 10413 9153
rect 10463 9173 10505 9211
rect 10463 9153 10477 9173
rect 10497 9153 10505 9173
rect 10463 9111 10505 9153
rect 10582 9173 10626 9211
rect 10582 9153 10594 9173
rect 10614 9153 10626 9173
rect 10582 9111 10626 9153
rect 10676 9173 10718 9211
rect 10676 9153 10690 9173
rect 10710 9153 10718 9173
rect 10676 9111 10718 9153
rect 10790 9173 10834 9211
rect 10790 9153 10802 9173
rect 10822 9153 10834 9173
rect 10790 9111 10834 9153
rect 10884 9173 10926 9211
rect 10884 9153 10898 9173
rect 10918 9153 10926 9173
rect 10884 9111 10926 9153
rect 11000 9173 11042 9211
rect 11000 9153 11008 9173
rect 11028 9153 11042 9173
rect 11000 9111 11042 9153
rect 11092 9180 11137 9211
rect 11092 9173 11136 9180
rect 11092 9153 11104 9173
rect 11124 9153 11136 9173
rect 15425 9214 15469 9252
rect 15425 9194 15437 9214
rect 15457 9194 15469 9214
rect 11092 9111 11136 9153
rect 13856 9113 13900 9155
rect 1276 8924 1320 8962
rect 1276 8904 1288 8924
rect 1308 8904 1320 8924
rect 1276 8862 1320 8904
rect 1370 8924 1412 8962
rect 1370 8904 1384 8924
rect 1404 8904 1412 8924
rect 1370 8862 1412 8904
rect 1489 8924 1533 8962
rect 1489 8904 1501 8924
rect 1521 8904 1533 8924
rect 1489 8862 1533 8904
rect 1583 8924 1625 8962
rect 1583 8904 1597 8924
rect 1617 8904 1625 8924
rect 1583 8862 1625 8904
rect 1697 8924 1741 8962
rect 1697 8904 1709 8924
rect 1729 8904 1741 8924
rect 1697 8862 1741 8904
rect 1791 8924 1833 8962
rect 1791 8904 1805 8924
rect 1825 8904 1833 8924
rect 1791 8862 1833 8904
rect 1907 8924 1949 8962
rect 1907 8904 1915 8924
rect 1935 8904 1949 8924
rect 1907 8862 1949 8904
rect 1999 8931 2044 8962
rect 1999 8924 2043 8931
rect 1999 8904 2011 8924
rect 2031 8904 2043 8924
rect 1999 8862 2043 8904
rect 6332 8965 6376 9003
rect 6332 8945 6344 8965
rect 6364 8945 6376 8965
rect 2886 8798 2930 8840
rect 2886 8778 2898 8798
rect 2918 8778 2930 8798
rect 2886 8771 2930 8778
rect 2885 8740 2930 8771
rect 2980 8798 3022 8840
rect 2980 8778 2994 8798
rect 3014 8778 3022 8798
rect 2980 8740 3022 8778
rect 3096 8798 3138 8840
rect 3096 8778 3104 8798
rect 3124 8778 3138 8798
rect 3096 8740 3138 8778
rect 3188 8798 3232 8840
rect 3188 8778 3200 8798
rect 3220 8778 3232 8798
rect 3188 8740 3232 8778
rect 3304 8798 3346 8840
rect 3304 8778 3312 8798
rect 3332 8778 3346 8798
rect 3304 8740 3346 8778
rect 3396 8798 3440 8840
rect 3396 8778 3408 8798
rect 3428 8778 3440 8798
rect 3396 8740 3440 8778
rect 3517 8798 3559 8840
rect 3517 8778 3525 8798
rect 3545 8778 3559 8798
rect 3517 8740 3559 8778
rect 3609 8798 3653 8840
rect 6332 8903 6376 8945
rect 6426 8965 6468 9003
rect 6426 8945 6440 8965
rect 6460 8945 6468 8965
rect 6426 8903 6468 8945
rect 6545 8965 6589 9003
rect 6545 8945 6557 8965
rect 6577 8945 6589 8965
rect 6545 8903 6589 8945
rect 6639 8965 6681 9003
rect 6639 8945 6653 8965
rect 6673 8945 6681 8965
rect 6639 8903 6681 8945
rect 6753 8965 6797 9003
rect 6753 8945 6765 8965
rect 6785 8945 6797 8965
rect 6753 8903 6797 8945
rect 6847 8965 6889 9003
rect 6847 8945 6861 8965
rect 6881 8945 6889 8965
rect 6847 8903 6889 8945
rect 6963 8965 7005 9003
rect 6963 8945 6971 8965
rect 6991 8945 7005 8965
rect 6963 8903 7005 8945
rect 7055 8972 7100 9003
rect 13856 9093 13868 9113
rect 13888 9093 13900 9113
rect 13856 9086 13900 9093
rect 7055 8965 7099 8972
rect 7055 8945 7067 8965
rect 7087 8945 7099 8965
rect 13855 9055 13900 9086
rect 13950 9113 13992 9155
rect 13950 9093 13964 9113
rect 13984 9093 13992 9113
rect 13950 9055 13992 9093
rect 14066 9113 14108 9155
rect 14066 9093 14074 9113
rect 14094 9093 14108 9113
rect 14066 9055 14108 9093
rect 14158 9113 14202 9155
rect 14158 9093 14170 9113
rect 14190 9093 14202 9113
rect 14158 9055 14202 9093
rect 14274 9113 14316 9155
rect 14274 9093 14282 9113
rect 14302 9093 14316 9113
rect 14274 9055 14316 9093
rect 14366 9113 14410 9155
rect 14366 9093 14378 9113
rect 14398 9093 14410 9113
rect 14366 9055 14410 9093
rect 14487 9113 14529 9155
rect 14487 9093 14495 9113
rect 14515 9093 14529 9113
rect 14487 9055 14529 9093
rect 14579 9113 14623 9155
rect 15425 9152 15469 9194
rect 15519 9214 15561 9252
rect 15519 9194 15533 9214
rect 15553 9194 15561 9214
rect 15519 9152 15561 9194
rect 15638 9214 15682 9252
rect 15638 9194 15650 9214
rect 15670 9194 15682 9214
rect 15638 9152 15682 9194
rect 15732 9214 15774 9252
rect 15732 9194 15746 9214
rect 15766 9194 15774 9214
rect 15732 9152 15774 9194
rect 15846 9214 15890 9252
rect 15846 9194 15858 9214
rect 15878 9194 15890 9214
rect 15846 9152 15890 9194
rect 15940 9214 15982 9252
rect 15940 9194 15954 9214
rect 15974 9194 15982 9214
rect 15940 9152 15982 9194
rect 16056 9214 16098 9252
rect 16056 9194 16064 9214
rect 16084 9194 16098 9214
rect 16056 9152 16098 9194
rect 16148 9221 16193 9252
rect 16148 9214 16192 9221
rect 16148 9194 16160 9214
rect 16180 9194 16192 9214
rect 16148 9152 16192 9194
rect 18912 9154 18956 9196
rect 14579 9093 14591 9113
rect 14611 9093 14623 9113
rect 14579 9055 14623 9093
rect 18912 9134 18924 9154
rect 18944 9134 18956 9154
rect 18912 9127 18956 9134
rect 18911 9096 18956 9127
rect 19006 9154 19048 9196
rect 19006 9134 19020 9154
rect 19040 9134 19048 9154
rect 19006 9096 19048 9134
rect 19122 9154 19164 9196
rect 19122 9134 19130 9154
rect 19150 9134 19164 9154
rect 19122 9096 19164 9134
rect 19214 9154 19258 9196
rect 19214 9134 19226 9154
rect 19246 9134 19258 9154
rect 19214 9096 19258 9134
rect 19330 9154 19372 9196
rect 19330 9134 19338 9154
rect 19358 9134 19372 9154
rect 19330 9096 19372 9134
rect 19422 9154 19466 9196
rect 19422 9134 19434 9154
rect 19454 9134 19466 9154
rect 19422 9096 19466 9134
rect 19543 9154 19585 9196
rect 19543 9134 19551 9154
rect 19571 9134 19585 9154
rect 19543 9096 19585 9134
rect 19635 9154 19679 9196
rect 19635 9134 19647 9154
rect 19667 9134 19679 9154
rect 19635 9096 19679 9134
rect 7055 8903 7099 8945
rect 3609 8778 3621 8798
rect 3641 8778 3653 8798
rect 3609 8740 3653 8778
rect 7942 8839 7986 8881
rect 7942 8819 7954 8839
rect 7974 8819 7986 8839
rect 7942 8812 7986 8819
rect 7941 8781 7986 8812
rect 8036 8839 8078 8881
rect 8036 8819 8050 8839
rect 8070 8819 8078 8839
rect 8036 8781 8078 8819
rect 8152 8839 8194 8881
rect 8152 8819 8160 8839
rect 8180 8819 8194 8839
rect 8152 8781 8194 8819
rect 8244 8839 8288 8881
rect 8244 8819 8256 8839
rect 8276 8819 8288 8839
rect 8244 8781 8288 8819
rect 8360 8839 8402 8881
rect 8360 8819 8368 8839
rect 8388 8819 8402 8839
rect 8360 8781 8402 8819
rect 8452 8839 8496 8881
rect 8452 8819 8464 8839
rect 8484 8819 8496 8839
rect 8452 8781 8496 8819
rect 8573 8839 8615 8881
rect 8573 8819 8581 8839
rect 8601 8819 8615 8839
rect 8573 8781 8615 8819
rect 8665 8839 8709 8881
rect 11307 8929 11351 8967
rect 11307 8909 11319 8929
rect 11339 8909 11351 8929
rect 8665 8819 8677 8839
rect 8697 8819 8709 8839
rect 8665 8781 8709 8819
rect 11307 8867 11351 8909
rect 11401 8929 11443 8967
rect 11401 8909 11415 8929
rect 11435 8909 11443 8929
rect 11401 8867 11443 8909
rect 11520 8929 11564 8967
rect 11520 8909 11532 8929
rect 11552 8909 11564 8929
rect 11520 8867 11564 8909
rect 11614 8929 11656 8967
rect 11614 8909 11628 8929
rect 11648 8909 11656 8929
rect 11614 8867 11656 8909
rect 11728 8929 11772 8967
rect 11728 8909 11740 8929
rect 11760 8909 11772 8929
rect 11728 8867 11772 8909
rect 11822 8929 11864 8967
rect 11822 8909 11836 8929
rect 11856 8909 11864 8929
rect 11822 8867 11864 8909
rect 11938 8929 11980 8967
rect 11938 8909 11946 8929
rect 11966 8909 11980 8929
rect 11938 8867 11980 8909
rect 12030 8936 12075 8967
rect 12030 8929 12074 8936
rect 12030 8909 12042 8929
rect 12062 8909 12074 8929
rect 12030 8867 12074 8909
rect 16363 8970 16407 9008
rect 16363 8950 16375 8970
rect 16395 8950 16407 8970
rect 12917 8803 12961 8845
rect 337 8614 381 8652
rect 337 8594 349 8614
rect 369 8594 381 8614
rect 337 8552 381 8594
rect 431 8614 473 8652
rect 431 8594 445 8614
rect 465 8594 473 8614
rect 431 8552 473 8594
rect 550 8614 594 8652
rect 550 8594 562 8614
rect 582 8594 594 8614
rect 550 8552 594 8594
rect 644 8614 686 8652
rect 644 8594 658 8614
rect 678 8594 686 8614
rect 644 8552 686 8594
rect 758 8614 802 8652
rect 758 8594 770 8614
rect 790 8594 802 8614
rect 758 8552 802 8594
rect 852 8614 894 8652
rect 852 8594 866 8614
rect 886 8594 894 8614
rect 852 8552 894 8594
rect 968 8614 1010 8652
rect 968 8594 976 8614
rect 996 8594 1010 8614
rect 968 8552 1010 8594
rect 1060 8621 1105 8652
rect 1060 8614 1104 8621
rect 1060 8594 1072 8614
rect 1092 8594 1104 8614
rect 5393 8655 5437 8693
rect 5393 8635 5405 8655
rect 5425 8635 5437 8655
rect 1060 8552 1104 8594
rect 3824 8554 3868 8596
rect 3824 8534 3836 8554
rect 3856 8534 3868 8554
rect 3824 8527 3868 8534
rect 3823 8496 3868 8527
rect 3918 8554 3960 8596
rect 3918 8534 3932 8554
rect 3952 8534 3960 8554
rect 3918 8496 3960 8534
rect 4034 8554 4076 8596
rect 4034 8534 4042 8554
rect 4062 8534 4076 8554
rect 4034 8496 4076 8534
rect 4126 8554 4170 8596
rect 4126 8534 4138 8554
rect 4158 8534 4170 8554
rect 4126 8496 4170 8534
rect 4242 8554 4284 8596
rect 4242 8534 4250 8554
rect 4270 8534 4284 8554
rect 4242 8496 4284 8534
rect 4334 8554 4378 8596
rect 4334 8534 4346 8554
rect 4366 8534 4378 8554
rect 4334 8496 4378 8534
rect 4455 8554 4497 8596
rect 4455 8534 4463 8554
rect 4483 8534 4497 8554
rect 4455 8496 4497 8534
rect 4547 8554 4591 8596
rect 5393 8593 5437 8635
rect 5487 8655 5529 8693
rect 5487 8635 5501 8655
rect 5521 8635 5529 8655
rect 5487 8593 5529 8635
rect 5606 8655 5650 8693
rect 5606 8635 5618 8655
rect 5638 8635 5650 8655
rect 5606 8593 5650 8635
rect 5700 8655 5742 8693
rect 5700 8635 5714 8655
rect 5734 8635 5742 8655
rect 5700 8593 5742 8635
rect 5814 8655 5858 8693
rect 5814 8635 5826 8655
rect 5846 8635 5858 8655
rect 5814 8593 5858 8635
rect 5908 8655 5950 8693
rect 5908 8635 5922 8655
rect 5942 8635 5950 8655
rect 5908 8593 5950 8635
rect 6024 8655 6066 8693
rect 6024 8635 6032 8655
rect 6052 8635 6066 8655
rect 6024 8593 6066 8635
rect 6116 8662 6161 8693
rect 12917 8783 12929 8803
rect 12949 8783 12961 8803
rect 12917 8776 12961 8783
rect 6116 8655 6160 8662
rect 6116 8635 6128 8655
rect 6148 8635 6160 8655
rect 12916 8745 12961 8776
rect 13011 8803 13053 8845
rect 13011 8783 13025 8803
rect 13045 8783 13053 8803
rect 13011 8745 13053 8783
rect 13127 8803 13169 8845
rect 13127 8783 13135 8803
rect 13155 8783 13169 8803
rect 13127 8745 13169 8783
rect 13219 8803 13263 8845
rect 13219 8783 13231 8803
rect 13251 8783 13263 8803
rect 13219 8745 13263 8783
rect 13335 8803 13377 8845
rect 13335 8783 13343 8803
rect 13363 8783 13377 8803
rect 13335 8745 13377 8783
rect 13427 8803 13471 8845
rect 13427 8783 13439 8803
rect 13459 8783 13471 8803
rect 13427 8745 13471 8783
rect 13548 8803 13590 8845
rect 13548 8783 13556 8803
rect 13576 8783 13590 8803
rect 13548 8745 13590 8783
rect 13640 8803 13684 8845
rect 16363 8908 16407 8950
rect 16457 8970 16499 9008
rect 16457 8950 16471 8970
rect 16491 8950 16499 8970
rect 16457 8908 16499 8950
rect 16576 8970 16620 9008
rect 16576 8950 16588 8970
rect 16608 8950 16620 8970
rect 16576 8908 16620 8950
rect 16670 8970 16712 9008
rect 16670 8950 16684 8970
rect 16704 8950 16712 8970
rect 16670 8908 16712 8950
rect 16784 8970 16828 9008
rect 16784 8950 16796 8970
rect 16816 8950 16828 8970
rect 16784 8908 16828 8950
rect 16878 8970 16920 9008
rect 16878 8950 16892 8970
rect 16912 8950 16920 8970
rect 16878 8908 16920 8950
rect 16994 8970 17036 9008
rect 16994 8950 17002 8970
rect 17022 8950 17036 8970
rect 16994 8908 17036 8950
rect 17086 8977 17131 9008
rect 17086 8970 17130 8977
rect 17086 8950 17098 8970
rect 17118 8950 17130 8970
rect 17086 8908 17130 8950
rect 13640 8783 13652 8803
rect 13672 8783 13684 8803
rect 13640 8745 13684 8783
rect 17973 8844 18017 8886
rect 17973 8824 17985 8844
rect 18005 8824 18017 8844
rect 17973 8817 18017 8824
rect 17972 8786 18017 8817
rect 18067 8844 18109 8886
rect 18067 8824 18081 8844
rect 18101 8824 18109 8844
rect 18067 8786 18109 8824
rect 18183 8844 18225 8886
rect 18183 8824 18191 8844
rect 18211 8824 18225 8844
rect 18183 8786 18225 8824
rect 18275 8844 18319 8886
rect 18275 8824 18287 8844
rect 18307 8824 18319 8844
rect 18275 8786 18319 8824
rect 18391 8844 18433 8886
rect 18391 8824 18399 8844
rect 18419 8824 18433 8844
rect 18391 8786 18433 8824
rect 18483 8844 18527 8886
rect 18483 8824 18495 8844
rect 18515 8824 18527 8844
rect 18483 8786 18527 8824
rect 18604 8844 18646 8886
rect 18604 8824 18612 8844
rect 18632 8824 18646 8844
rect 18604 8786 18646 8824
rect 18696 8844 18740 8886
rect 18696 8824 18708 8844
rect 18728 8824 18740 8844
rect 18696 8786 18740 8824
rect 6116 8593 6160 8635
rect 8880 8595 8924 8637
rect 4547 8534 4559 8554
rect 4579 8534 4591 8554
rect 4547 8496 4591 8534
rect 8880 8575 8892 8595
rect 8912 8575 8924 8595
rect 8880 8568 8924 8575
rect 8879 8537 8924 8568
rect 8974 8595 9016 8637
rect 8974 8575 8988 8595
rect 9008 8575 9016 8595
rect 8974 8537 9016 8575
rect 9090 8595 9132 8637
rect 9090 8575 9098 8595
rect 9118 8575 9132 8595
rect 9090 8537 9132 8575
rect 9182 8595 9226 8637
rect 9182 8575 9194 8595
rect 9214 8575 9226 8595
rect 9182 8537 9226 8575
rect 9298 8595 9340 8637
rect 9298 8575 9306 8595
rect 9326 8575 9340 8595
rect 9298 8537 9340 8575
rect 9390 8595 9434 8637
rect 9390 8575 9402 8595
rect 9422 8575 9434 8595
rect 9390 8537 9434 8575
rect 9511 8595 9553 8637
rect 9511 8575 9519 8595
rect 9539 8575 9553 8595
rect 9511 8537 9553 8575
rect 9603 8595 9647 8637
rect 9603 8575 9615 8595
rect 9635 8575 9647 8595
rect 10368 8619 10412 8657
rect 10368 8599 10380 8619
rect 10400 8599 10412 8619
rect 9603 8537 9647 8575
rect 10368 8557 10412 8599
rect 10462 8619 10504 8657
rect 10462 8599 10476 8619
rect 10496 8599 10504 8619
rect 10462 8557 10504 8599
rect 10581 8619 10625 8657
rect 10581 8599 10593 8619
rect 10613 8599 10625 8619
rect 10581 8557 10625 8599
rect 10675 8619 10717 8657
rect 10675 8599 10689 8619
rect 10709 8599 10717 8619
rect 10675 8557 10717 8599
rect 10789 8619 10833 8657
rect 10789 8599 10801 8619
rect 10821 8599 10833 8619
rect 10789 8557 10833 8599
rect 10883 8619 10925 8657
rect 10883 8599 10897 8619
rect 10917 8599 10925 8619
rect 10883 8557 10925 8599
rect 10999 8619 11041 8657
rect 10999 8599 11007 8619
rect 11027 8599 11041 8619
rect 10999 8557 11041 8599
rect 11091 8626 11136 8657
rect 11091 8619 11135 8626
rect 11091 8599 11103 8619
rect 11123 8599 11135 8619
rect 15424 8660 15468 8698
rect 15424 8640 15436 8660
rect 15456 8640 15468 8660
rect 11091 8557 11135 8599
rect 13855 8559 13899 8601
rect 13855 8539 13867 8559
rect 13887 8539 13899 8559
rect 13855 8532 13899 8539
rect 13854 8501 13899 8532
rect 13949 8559 13991 8601
rect 13949 8539 13963 8559
rect 13983 8539 13991 8559
rect 13949 8501 13991 8539
rect 14065 8559 14107 8601
rect 14065 8539 14073 8559
rect 14093 8539 14107 8559
rect 14065 8501 14107 8539
rect 14157 8559 14201 8601
rect 14157 8539 14169 8559
rect 14189 8539 14201 8559
rect 14157 8501 14201 8539
rect 14273 8559 14315 8601
rect 14273 8539 14281 8559
rect 14301 8539 14315 8559
rect 14273 8501 14315 8539
rect 14365 8559 14409 8601
rect 14365 8539 14377 8559
rect 14397 8539 14409 8559
rect 14365 8501 14409 8539
rect 14486 8559 14528 8601
rect 14486 8539 14494 8559
rect 14514 8539 14528 8559
rect 14486 8501 14528 8539
rect 14578 8559 14622 8601
rect 15424 8598 15468 8640
rect 15518 8660 15560 8698
rect 15518 8640 15532 8660
rect 15552 8640 15560 8660
rect 15518 8598 15560 8640
rect 15637 8660 15681 8698
rect 15637 8640 15649 8660
rect 15669 8640 15681 8660
rect 15637 8598 15681 8640
rect 15731 8660 15773 8698
rect 15731 8640 15745 8660
rect 15765 8640 15773 8660
rect 15731 8598 15773 8640
rect 15845 8660 15889 8698
rect 15845 8640 15857 8660
rect 15877 8640 15889 8660
rect 15845 8598 15889 8640
rect 15939 8660 15981 8698
rect 15939 8640 15953 8660
rect 15973 8640 15981 8660
rect 15939 8598 15981 8640
rect 16055 8660 16097 8698
rect 16055 8640 16063 8660
rect 16083 8640 16097 8660
rect 16055 8598 16097 8640
rect 16147 8667 16192 8698
rect 16147 8660 16191 8667
rect 16147 8640 16159 8660
rect 16179 8640 16191 8660
rect 16147 8598 16191 8640
rect 18911 8600 18955 8642
rect 14578 8539 14590 8559
rect 14610 8539 14622 8559
rect 14578 8501 14622 8539
rect 18911 8580 18923 8600
rect 18943 8580 18955 8600
rect 18911 8573 18955 8580
rect 18910 8542 18955 8573
rect 19005 8600 19047 8642
rect 19005 8580 19019 8600
rect 19039 8580 19047 8600
rect 19005 8542 19047 8580
rect 19121 8600 19163 8642
rect 19121 8580 19129 8600
rect 19149 8580 19163 8600
rect 19121 8542 19163 8580
rect 19213 8600 19257 8642
rect 19213 8580 19225 8600
rect 19245 8580 19257 8600
rect 19213 8542 19257 8580
rect 19329 8600 19371 8642
rect 19329 8580 19337 8600
rect 19357 8580 19371 8600
rect 19329 8542 19371 8580
rect 19421 8600 19465 8642
rect 19421 8580 19433 8600
rect 19453 8580 19465 8600
rect 19421 8542 19465 8580
rect 19542 8600 19584 8642
rect 19542 8580 19550 8600
rect 19570 8580 19584 8600
rect 19542 8542 19584 8580
rect 19634 8600 19678 8642
rect 19634 8580 19646 8600
rect 19666 8580 19678 8600
rect 19634 8542 19678 8580
rect 1417 8332 1461 8370
rect 1417 8312 1429 8332
rect 1449 8312 1461 8332
rect 1417 8270 1461 8312
rect 1511 8332 1553 8370
rect 1511 8312 1525 8332
rect 1545 8312 1553 8332
rect 1511 8270 1553 8312
rect 1630 8332 1674 8370
rect 1630 8312 1642 8332
rect 1662 8312 1674 8332
rect 1630 8270 1674 8312
rect 1724 8332 1766 8370
rect 1724 8312 1738 8332
rect 1758 8312 1766 8332
rect 1724 8270 1766 8312
rect 1838 8332 1882 8370
rect 1838 8312 1850 8332
rect 1870 8312 1882 8332
rect 1838 8270 1882 8312
rect 1932 8332 1974 8370
rect 1932 8312 1946 8332
rect 1966 8312 1974 8332
rect 1932 8270 1974 8312
rect 2048 8332 2090 8370
rect 2048 8312 2056 8332
rect 2076 8312 2090 8332
rect 2048 8270 2090 8312
rect 2140 8339 2185 8370
rect 2140 8332 2184 8339
rect 2140 8312 2152 8332
rect 2172 8312 2184 8332
rect 6473 8373 6517 8411
rect 6473 8353 6485 8373
rect 6505 8353 6517 8373
rect 2140 8270 2184 8312
rect 2746 8287 2790 8329
rect 2746 8267 2758 8287
rect 2778 8267 2790 8287
rect 2746 8260 2790 8267
rect 2745 8229 2790 8260
rect 2840 8287 2882 8329
rect 2840 8267 2854 8287
rect 2874 8267 2882 8287
rect 2840 8229 2882 8267
rect 2956 8287 2998 8329
rect 2956 8267 2964 8287
rect 2984 8267 2998 8287
rect 2956 8229 2998 8267
rect 3048 8287 3092 8329
rect 3048 8267 3060 8287
rect 3080 8267 3092 8287
rect 3048 8229 3092 8267
rect 3164 8287 3206 8329
rect 3164 8267 3172 8287
rect 3192 8267 3206 8287
rect 3164 8229 3206 8267
rect 3256 8287 3300 8329
rect 3256 8267 3268 8287
rect 3288 8267 3300 8287
rect 3256 8229 3300 8267
rect 3377 8287 3419 8329
rect 3377 8267 3385 8287
rect 3405 8267 3419 8287
rect 3377 8229 3419 8267
rect 3469 8287 3513 8329
rect 6473 8311 6517 8353
rect 6567 8373 6609 8411
rect 6567 8353 6581 8373
rect 6601 8353 6609 8373
rect 6567 8311 6609 8353
rect 6686 8373 6730 8411
rect 6686 8353 6698 8373
rect 6718 8353 6730 8373
rect 6686 8311 6730 8353
rect 6780 8373 6822 8411
rect 6780 8353 6794 8373
rect 6814 8353 6822 8373
rect 6780 8311 6822 8353
rect 6894 8373 6938 8411
rect 6894 8353 6906 8373
rect 6926 8353 6938 8373
rect 6894 8311 6938 8353
rect 6988 8373 7030 8411
rect 6988 8353 7002 8373
rect 7022 8353 7030 8373
rect 6988 8311 7030 8353
rect 7104 8373 7146 8411
rect 7104 8353 7112 8373
rect 7132 8353 7146 8373
rect 7104 8311 7146 8353
rect 7196 8380 7241 8411
rect 7196 8373 7240 8380
rect 7196 8353 7208 8373
rect 7228 8353 7240 8373
rect 7196 8311 7240 8353
rect 7802 8328 7846 8370
rect 3469 8267 3481 8287
rect 3501 8267 3513 8287
rect 3469 8229 3513 8267
rect 7802 8308 7814 8328
rect 7834 8308 7846 8328
rect 7802 8301 7846 8308
rect 7801 8270 7846 8301
rect 7896 8328 7938 8370
rect 7896 8308 7910 8328
rect 7930 8308 7938 8328
rect 7896 8270 7938 8308
rect 8012 8328 8054 8370
rect 8012 8308 8020 8328
rect 8040 8308 8054 8328
rect 8012 8270 8054 8308
rect 8104 8328 8148 8370
rect 8104 8308 8116 8328
rect 8136 8308 8148 8328
rect 8104 8270 8148 8308
rect 8220 8328 8262 8370
rect 8220 8308 8228 8328
rect 8248 8308 8262 8328
rect 8220 8270 8262 8308
rect 8312 8328 8356 8370
rect 8312 8308 8324 8328
rect 8344 8308 8356 8328
rect 8312 8270 8356 8308
rect 8433 8328 8475 8370
rect 8433 8308 8441 8328
rect 8461 8308 8475 8328
rect 8433 8270 8475 8308
rect 8525 8328 8569 8370
rect 8525 8308 8537 8328
rect 8557 8308 8569 8328
rect 8525 8270 8569 8308
rect 11448 8337 11492 8375
rect 11448 8317 11460 8337
rect 11480 8317 11492 8337
rect 11448 8275 11492 8317
rect 11542 8337 11584 8375
rect 11542 8317 11556 8337
rect 11576 8317 11584 8337
rect 11542 8275 11584 8317
rect 11661 8337 11705 8375
rect 11661 8317 11673 8337
rect 11693 8317 11705 8337
rect 11661 8275 11705 8317
rect 11755 8337 11797 8375
rect 11755 8317 11769 8337
rect 11789 8317 11797 8337
rect 11755 8275 11797 8317
rect 11869 8337 11913 8375
rect 11869 8317 11881 8337
rect 11901 8317 11913 8337
rect 11869 8275 11913 8317
rect 11963 8337 12005 8375
rect 11963 8317 11977 8337
rect 11997 8317 12005 8337
rect 11963 8275 12005 8317
rect 12079 8337 12121 8375
rect 12079 8317 12087 8337
rect 12107 8317 12121 8337
rect 12079 8275 12121 8317
rect 12171 8344 12216 8375
rect 12171 8337 12215 8344
rect 12171 8317 12183 8337
rect 12203 8317 12215 8337
rect 16504 8378 16548 8416
rect 16504 8358 16516 8378
rect 16536 8358 16548 8378
rect 12171 8275 12215 8317
rect 12777 8292 12821 8334
rect 12777 8272 12789 8292
rect 12809 8272 12821 8292
rect 12777 8265 12821 8272
rect 12776 8234 12821 8265
rect 12871 8292 12913 8334
rect 12871 8272 12885 8292
rect 12905 8272 12913 8292
rect 12871 8234 12913 8272
rect 12987 8292 13029 8334
rect 12987 8272 12995 8292
rect 13015 8272 13029 8292
rect 12987 8234 13029 8272
rect 13079 8292 13123 8334
rect 13079 8272 13091 8292
rect 13111 8272 13123 8292
rect 13079 8234 13123 8272
rect 13195 8292 13237 8334
rect 13195 8272 13203 8292
rect 13223 8272 13237 8292
rect 13195 8234 13237 8272
rect 13287 8292 13331 8334
rect 13287 8272 13299 8292
rect 13319 8272 13331 8292
rect 13287 8234 13331 8272
rect 13408 8292 13450 8334
rect 13408 8272 13416 8292
rect 13436 8272 13450 8292
rect 13408 8234 13450 8272
rect 13500 8292 13544 8334
rect 16504 8316 16548 8358
rect 16598 8378 16640 8416
rect 16598 8358 16612 8378
rect 16632 8358 16640 8378
rect 16598 8316 16640 8358
rect 16717 8378 16761 8416
rect 16717 8358 16729 8378
rect 16749 8358 16761 8378
rect 16717 8316 16761 8358
rect 16811 8378 16853 8416
rect 16811 8358 16825 8378
rect 16845 8358 16853 8378
rect 16811 8316 16853 8358
rect 16925 8378 16969 8416
rect 16925 8358 16937 8378
rect 16957 8358 16969 8378
rect 16925 8316 16969 8358
rect 17019 8378 17061 8416
rect 17019 8358 17033 8378
rect 17053 8358 17061 8378
rect 17019 8316 17061 8358
rect 17135 8378 17177 8416
rect 17135 8358 17143 8378
rect 17163 8358 17177 8378
rect 17135 8316 17177 8358
rect 17227 8385 17272 8416
rect 17227 8378 17271 8385
rect 17227 8358 17239 8378
rect 17259 8358 17271 8378
rect 17227 8316 17271 8358
rect 17833 8333 17877 8375
rect 13500 8272 13512 8292
rect 13532 8272 13544 8292
rect 13500 8234 13544 8272
rect 17833 8313 17845 8333
rect 17865 8313 17877 8333
rect 17833 8306 17877 8313
rect 17832 8275 17877 8306
rect 17927 8333 17969 8375
rect 17927 8313 17941 8333
rect 17961 8313 17969 8333
rect 17927 8275 17969 8313
rect 18043 8333 18085 8375
rect 18043 8313 18051 8333
rect 18071 8313 18085 8333
rect 18043 8275 18085 8313
rect 18135 8333 18179 8375
rect 18135 8313 18147 8333
rect 18167 8313 18179 8333
rect 18135 8275 18179 8313
rect 18251 8333 18293 8375
rect 18251 8313 18259 8333
rect 18279 8313 18293 8333
rect 18251 8275 18293 8313
rect 18343 8333 18387 8375
rect 18343 8313 18355 8333
rect 18375 8313 18387 8333
rect 18343 8275 18387 8313
rect 18464 8333 18506 8375
rect 18464 8313 18472 8333
rect 18492 8313 18506 8333
rect 18464 8275 18506 8313
rect 18556 8333 18600 8375
rect 18556 8313 18568 8333
rect 18588 8313 18600 8333
rect 18556 8275 18600 8313
rect 339 8065 383 8103
rect 339 8045 351 8065
rect 371 8045 383 8065
rect 339 8003 383 8045
rect 433 8065 475 8103
rect 433 8045 447 8065
rect 467 8045 475 8065
rect 433 8003 475 8045
rect 552 8065 596 8103
rect 552 8045 564 8065
rect 584 8045 596 8065
rect 552 8003 596 8045
rect 646 8065 688 8103
rect 646 8045 660 8065
rect 680 8045 688 8065
rect 646 8003 688 8045
rect 760 8065 804 8103
rect 760 8045 772 8065
rect 792 8045 804 8065
rect 760 8003 804 8045
rect 854 8065 896 8103
rect 854 8045 868 8065
rect 888 8045 896 8065
rect 854 8003 896 8045
rect 970 8065 1012 8103
rect 970 8045 978 8065
rect 998 8045 1012 8065
rect 970 8003 1012 8045
rect 1062 8072 1107 8103
rect 1062 8065 1106 8072
rect 1062 8045 1074 8065
rect 1094 8045 1106 8065
rect 5395 8106 5439 8144
rect 5395 8086 5407 8106
rect 5427 8086 5439 8106
rect 1062 8003 1106 8045
rect 3826 8005 3870 8047
rect 3826 7985 3838 8005
rect 3858 7985 3870 8005
rect 3826 7978 3870 7985
rect 3825 7947 3870 7978
rect 3920 8005 3962 8047
rect 3920 7985 3934 8005
rect 3954 7985 3962 8005
rect 3920 7947 3962 7985
rect 4036 8005 4078 8047
rect 4036 7985 4044 8005
rect 4064 7985 4078 8005
rect 4036 7947 4078 7985
rect 4128 8005 4172 8047
rect 4128 7985 4140 8005
rect 4160 7985 4172 8005
rect 4128 7947 4172 7985
rect 4244 8005 4286 8047
rect 4244 7985 4252 8005
rect 4272 7985 4286 8005
rect 4244 7947 4286 7985
rect 4336 8005 4380 8047
rect 4336 7985 4348 8005
rect 4368 7985 4380 8005
rect 4336 7947 4380 7985
rect 4457 8005 4499 8047
rect 4457 7985 4465 8005
rect 4485 7985 4499 8005
rect 4457 7947 4499 7985
rect 4549 8005 4593 8047
rect 5395 8044 5439 8086
rect 5489 8106 5531 8144
rect 5489 8086 5503 8106
rect 5523 8086 5531 8106
rect 5489 8044 5531 8086
rect 5608 8106 5652 8144
rect 5608 8086 5620 8106
rect 5640 8086 5652 8106
rect 5608 8044 5652 8086
rect 5702 8106 5744 8144
rect 5702 8086 5716 8106
rect 5736 8086 5744 8106
rect 5702 8044 5744 8086
rect 5816 8106 5860 8144
rect 5816 8086 5828 8106
rect 5848 8086 5860 8106
rect 5816 8044 5860 8086
rect 5910 8106 5952 8144
rect 5910 8086 5924 8106
rect 5944 8086 5952 8106
rect 5910 8044 5952 8086
rect 6026 8106 6068 8144
rect 6026 8086 6034 8106
rect 6054 8086 6068 8106
rect 6026 8044 6068 8086
rect 6118 8113 6163 8144
rect 6118 8106 6162 8113
rect 6118 8086 6130 8106
rect 6150 8086 6162 8106
rect 6118 8044 6162 8086
rect 8882 8046 8926 8088
rect 4549 7985 4561 8005
rect 4581 7985 4593 8005
rect 4549 7947 4593 7985
rect 8882 8026 8894 8046
rect 8914 8026 8926 8046
rect 8882 8019 8926 8026
rect 8881 7988 8926 8019
rect 8976 8046 9018 8088
rect 8976 8026 8990 8046
rect 9010 8026 9018 8046
rect 8976 7988 9018 8026
rect 9092 8046 9134 8088
rect 9092 8026 9100 8046
rect 9120 8026 9134 8046
rect 9092 7988 9134 8026
rect 9184 8046 9228 8088
rect 9184 8026 9196 8046
rect 9216 8026 9228 8046
rect 9184 7988 9228 8026
rect 9300 8046 9342 8088
rect 9300 8026 9308 8046
rect 9328 8026 9342 8046
rect 9300 7988 9342 8026
rect 9392 8046 9436 8088
rect 9392 8026 9404 8046
rect 9424 8026 9436 8046
rect 9392 7988 9436 8026
rect 9513 8046 9555 8088
rect 9513 8026 9521 8046
rect 9541 8026 9555 8046
rect 9513 7988 9555 8026
rect 9605 8046 9649 8088
rect 10370 8070 10414 8108
rect 9605 8026 9617 8046
rect 9637 8026 9649 8046
rect 9605 7988 9649 8026
rect 10370 8050 10382 8070
rect 10402 8050 10414 8070
rect 10370 8008 10414 8050
rect 10464 8070 10506 8108
rect 10464 8050 10478 8070
rect 10498 8050 10506 8070
rect 10464 8008 10506 8050
rect 10583 8070 10627 8108
rect 10583 8050 10595 8070
rect 10615 8050 10627 8070
rect 10583 8008 10627 8050
rect 10677 8070 10719 8108
rect 10677 8050 10691 8070
rect 10711 8050 10719 8070
rect 10677 8008 10719 8050
rect 10791 8070 10835 8108
rect 10791 8050 10803 8070
rect 10823 8050 10835 8070
rect 10791 8008 10835 8050
rect 10885 8070 10927 8108
rect 10885 8050 10899 8070
rect 10919 8050 10927 8070
rect 10885 8008 10927 8050
rect 11001 8070 11043 8108
rect 11001 8050 11009 8070
rect 11029 8050 11043 8070
rect 11001 8008 11043 8050
rect 11093 8077 11138 8108
rect 11093 8070 11137 8077
rect 11093 8050 11105 8070
rect 11125 8050 11137 8070
rect 15426 8111 15470 8149
rect 15426 8091 15438 8111
rect 15458 8091 15470 8111
rect 11093 8008 11137 8050
rect 13857 8010 13901 8052
rect 1277 7821 1321 7859
rect 1277 7801 1289 7821
rect 1309 7801 1321 7821
rect 1277 7759 1321 7801
rect 1371 7821 1413 7859
rect 1371 7801 1385 7821
rect 1405 7801 1413 7821
rect 1371 7759 1413 7801
rect 1490 7821 1534 7859
rect 1490 7801 1502 7821
rect 1522 7801 1534 7821
rect 1490 7759 1534 7801
rect 1584 7821 1626 7859
rect 1584 7801 1598 7821
rect 1618 7801 1626 7821
rect 1584 7759 1626 7801
rect 1698 7821 1742 7859
rect 1698 7801 1710 7821
rect 1730 7801 1742 7821
rect 1698 7759 1742 7801
rect 1792 7821 1834 7859
rect 1792 7801 1806 7821
rect 1826 7801 1834 7821
rect 1792 7759 1834 7801
rect 1908 7821 1950 7859
rect 1908 7801 1916 7821
rect 1936 7801 1950 7821
rect 1908 7759 1950 7801
rect 2000 7828 2045 7859
rect 2000 7821 2044 7828
rect 2000 7801 2012 7821
rect 2032 7801 2044 7821
rect 2000 7759 2044 7801
rect 6333 7862 6377 7900
rect 6333 7842 6345 7862
rect 6365 7842 6377 7862
rect 2887 7695 2931 7737
rect 2887 7675 2899 7695
rect 2919 7675 2931 7695
rect 2887 7668 2931 7675
rect 2886 7637 2931 7668
rect 2981 7695 3023 7737
rect 2981 7675 2995 7695
rect 3015 7675 3023 7695
rect 2981 7637 3023 7675
rect 3097 7695 3139 7737
rect 3097 7675 3105 7695
rect 3125 7675 3139 7695
rect 3097 7637 3139 7675
rect 3189 7695 3233 7737
rect 3189 7675 3201 7695
rect 3221 7675 3233 7695
rect 3189 7637 3233 7675
rect 3305 7695 3347 7737
rect 3305 7675 3313 7695
rect 3333 7675 3347 7695
rect 3305 7637 3347 7675
rect 3397 7695 3441 7737
rect 3397 7675 3409 7695
rect 3429 7675 3441 7695
rect 3397 7637 3441 7675
rect 3518 7695 3560 7737
rect 3518 7675 3526 7695
rect 3546 7675 3560 7695
rect 3518 7637 3560 7675
rect 3610 7695 3654 7737
rect 6333 7800 6377 7842
rect 6427 7862 6469 7900
rect 6427 7842 6441 7862
rect 6461 7842 6469 7862
rect 6427 7800 6469 7842
rect 6546 7862 6590 7900
rect 6546 7842 6558 7862
rect 6578 7842 6590 7862
rect 6546 7800 6590 7842
rect 6640 7862 6682 7900
rect 6640 7842 6654 7862
rect 6674 7842 6682 7862
rect 6640 7800 6682 7842
rect 6754 7862 6798 7900
rect 6754 7842 6766 7862
rect 6786 7842 6798 7862
rect 6754 7800 6798 7842
rect 6848 7862 6890 7900
rect 6848 7842 6862 7862
rect 6882 7842 6890 7862
rect 6848 7800 6890 7842
rect 6964 7862 7006 7900
rect 6964 7842 6972 7862
rect 6992 7842 7006 7862
rect 6964 7800 7006 7842
rect 7056 7869 7101 7900
rect 13857 7990 13869 8010
rect 13889 7990 13901 8010
rect 13857 7983 13901 7990
rect 7056 7862 7100 7869
rect 7056 7842 7068 7862
rect 7088 7842 7100 7862
rect 13856 7952 13901 7983
rect 13951 8010 13993 8052
rect 13951 7990 13965 8010
rect 13985 7990 13993 8010
rect 13951 7952 13993 7990
rect 14067 8010 14109 8052
rect 14067 7990 14075 8010
rect 14095 7990 14109 8010
rect 14067 7952 14109 7990
rect 14159 8010 14203 8052
rect 14159 7990 14171 8010
rect 14191 7990 14203 8010
rect 14159 7952 14203 7990
rect 14275 8010 14317 8052
rect 14275 7990 14283 8010
rect 14303 7990 14317 8010
rect 14275 7952 14317 7990
rect 14367 8010 14411 8052
rect 14367 7990 14379 8010
rect 14399 7990 14411 8010
rect 14367 7952 14411 7990
rect 14488 8010 14530 8052
rect 14488 7990 14496 8010
rect 14516 7990 14530 8010
rect 14488 7952 14530 7990
rect 14580 8010 14624 8052
rect 15426 8049 15470 8091
rect 15520 8111 15562 8149
rect 15520 8091 15534 8111
rect 15554 8091 15562 8111
rect 15520 8049 15562 8091
rect 15639 8111 15683 8149
rect 15639 8091 15651 8111
rect 15671 8091 15683 8111
rect 15639 8049 15683 8091
rect 15733 8111 15775 8149
rect 15733 8091 15747 8111
rect 15767 8091 15775 8111
rect 15733 8049 15775 8091
rect 15847 8111 15891 8149
rect 15847 8091 15859 8111
rect 15879 8091 15891 8111
rect 15847 8049 15891 8091
rect 15941 8111 15983 8149
rect 15941 8091 15955 8111
rect 15975 8091 15983 8111
rect 15941 8049 15983 8091
rect 16057 8111 16099 8149
rect 16057 8091 16065 8111
rect 16085 8091 16099 8111
rect 16057 8049 16099 8091
rect 16149 8118 16194 8149
rect 16149 8111 16193 8118
rect 16149 8091 16161 8111
rect 16181 8091 16193 8111
rect 16149 8049 16193 8091
rect 18913 8051 18957 8093
rect 14580 7990 14592 8010
rect 14612 7990 14624 8010
rect 14580 7952 14624 7990
rect 18913 8031 18925 8051
rect 18945 8031 18957 8051
rect 18913 8024 18957 8031
rect 18912 7993 18957 8024
rect 19007 8051 19049 8093
rect 19007 8031 19021 8051
rect 19041 8031 19049 8051
rect 19007 7993 19049 8031
rect 19123 8051 19165 8093
rect 19123 8031 19131 8051
rect 19151 8031 19165 8051
rect 19123 7993 19165 8031
rect 19215 8051 19259 8093
rect 19215 8031 19227 8051
rect 19247 8031 19259 8051
rect 19215 7993 19259 8031
rect 19331 8051 19373 8093
rect 19331 8031 19339 8051
rect 19359 8031 19373 8051
rect 19331 7993 19373 8031
rect 19423 8051 19467 8093
rect 19423 8031 19435 8051
rect 19455 8031 19467 8051
rect 19423 7993 19467 8031
rect 19544 8051 19586 8093
rect 19544 8031 19552 8051
rect 19572 8031 19586 8051
rect 19544 7993 19586 8031
rect 19636 8051 19680 8093
rect 19636 8031 19648 8051
rect 19668 8031 19680 8051
rect 19636 7993 19680 8031
rect 7056 7800 7100 7842
rect 3610 7675 3622 7695
rect 3642 7675 3654 7695
rect 3610 7637 3654 7675
rect 7943 7736 7987 7778
rect 7943 7716 7955 7736
rect 7975 7716 7987 7736
rect 7943 7709 7987 7716
rect 7942 7678 7987 7709
rect 8037 7736 8079 7778
rect 8037 7716 8051 7736
rect 8071 7716 8079 7736
rect 8037 7678 8079 7716
rect 8153 7736 8195 7778
rect 8153 7716 8161 7736
rect 8181 7716 8195 7736
rect 8153 7678 8195 7716
rect 8245 7736 8289 7778
rect 8245 7716 8257 7736
rect 8277 7716 8289 7736
rect 8245 7678 8289 7716
rect 8361 7736 8403 7778
rect 8361 7716 8369 7736
rect 8389 7716 8403 7736
rect 8361 7678 8403 7716
rect 8453 7736 8497 7778
rect 8453 7716 8465 7736
rect 8485 7716 8497 7736
rect 8453 7678 8497 7716
rect 8574 7736 8616 7778
rect 8574 7716 8582 7736
rect 8602 7716 8616 7736
rect 8574 7678 8616 7716
rect 8666 7736 8710 7778
rect 11308 7826 11352 7864
rect 11308 7806 11320 7826
rect 11340 7806 11352 7826
rect 8666 7716 8678 7736
rect 8698 7716 8710 7736
rect 8666 7678 8710 7716
rect 11308 7764 11352 7806
rect 11402 7826 11444 7864
rect 11402 7806 11416 7826
rect 11436 7806 11444 7826
rect 11402 7764 11444 7806
rect 11521 7826 11565 7864
rect 11521 7806 11533 7826
rect 11553 7806 11565 7826
rect 11521 7764 11565 7806
rect 11615 7826 11657 7864
rect 11615 7806 11629 7826
rect 11649 7806 11657 7826
rect 11615 7764 11657 7806
rect 11729 7826 11773 7864
rect 11729 7806 11741 7826
rect 11761 7806 11773 7826
rect 11729 7764 11773 7806
rect 11823 7826 11865 7864
rect 11823 7806 11837 7826
rect 11857 7806 11865 7826
rect 11823 7764 11865 7806
rect 11939 7826 11981 7864
rect 11939 7806 11947 7826
rect 11967 7806 11981 7826
rect 11939 7764 11981 7806
rect 12031 7833 12076 7864
rect 12031 7826 12075 7833
rect 12031 7806 12043 7826
rect 12063 7806 12075 7826
rect 12031 7764 12075 7806
rect 16364 7867 16408 7905
rect 16364 7847 16376 7867
rect 16396 7847 16408 7867
rect 12918 7700 12962 7742
rect 338 7511 382 7549
rect 338 7491 350 7511
rect 370 7491 382 7511
rect 338 7449 382 7491
rect 432 7511 474 7549
rect 432 7491 446 7511
rect 466 7491 474 7511
rect 432 7449 474 7491
rect 551 7511 595 7549
rect 551 7491 563 7511
rect 583 7491 595 7511
rect 551 7449 595 7491
rect 645 7511 687 7549
rect 645 7491 659 7511
rect 679 7491 687 7511
rect 645 7449 687 7491
rect 759 7511 803 7549
rect 759 7491 771 7511
rect 791 7491 803 7511
rect 759 7449 803 7491
rect 853 7511 895 7549
rect 853 7491 867 7511
rect 887 7491 895 7511
rect 853 7449 895 7491
rect 969 7511 1011 7549
rect 969 7491 977 7511
rect 997 7491 1011 7511
rect 969 7449 1011 7491
rect 1061 7518 1106 7549
rect 1061 7511 1105 7518
rect 1061 7491 1073 7511
rect 1093 7491 1105 7511
rect 5394 7552 5438 7590
rect 5394 7532 5406 7552
rect 5426 7532 5438 7552
rect 1061 7449 1105 7491
rect 3825 7451 3869 7493
rect 3825 7431 3837 7451
rect 3857 7431 3869 7451
rect 3825 7424 3869 7431
rect 3824 7393 3869 7424
rect 3919 7451 3961 7493
rect 3919 7431 3933 7451
rect 3953 7431 3961 7451
rect 3919 7393 3961 7431
rect 4035 7451 4077 7493
rect 4035 7431 4043 7451
rect 4063 7431 4077 7451
rect 4035 7393 4077 7431
rect 4127 7451 4171 7493
rect 4127 7431 4139 7451
rect 4159 7431 4171 7451
rect 4127 7393 4171 7431
rect 4243 7451 4285 7493
rect 4243 7431 4251 7451
rect 4271 7431 4285 7451
rect 4243 7393 4285 7431
rect 4335 7451 4379 7493
rect 4335 7431 4347 7451
rect 4367 7431 4379 7451
rect 4335 7393 4379 7431
rect 4456 7451 4498 7493
rect 4456 7431 4464 7451
rect 4484 7431 4498 7451
rect 4456 7393 4498 7431
rect 4548 7451 4592 7493
rect 5394 7490 5438 7532
rect 5488 7552 5530 7590
rect 5488 7532 5502 7552
rect 5522 7532 5530 7552
rect 5488 7490 5530 7532
rect 5607 7552 5651 7590
rect 5607 7532 5619 7552
rect 5639 7532 5651 7552
rect 5607 7490 5651 7532
rect 5701 7552 5743 7590
rect 5701 7532 5715 7552
rect 5735 7532 5743 7552
rect 5701 7490 5743 7532
rect 5815 7552 5859 7590
rect 5815 7532 5827 7552
rect 5847 7532 5859 7552
rect 5815 7490 5859 7532
rect 5909 7552 5951 7590
rect 5909 7532 5923 7552
rect 5943 7532 5951 7552
rect 5909 7490 5951 7532
rect 6025 7552 6067 7590
rect 6025 7532 6033 7552
rect 6053 7532 6067 7552
rect 6025 7490 6067 7532
rect 6117 7559 6162 7590
rect 12918 7680 12930 7700
rect 12950 7680 12962 7700
rect 12918 7673 12962 7680
rect 6117 7552 6161 7559
rect 6117 7532 6129 7552
rect 6149 7532 6161 7552
rect 12917 7642 12962 7673
rect 13012 7700 13054 7742
rect 13012 7680 13026 7700
rect 13046 7680 13054 7700
rect 13012 7642 13054 7680
rect 13128 7700 13170 7742
rect 13128 7680 13136 7700
rect 13156 7680 13170 7700
rect 13128 7642 13170 7680
rect 13220 7700 13264 7742
rect 13220 7680 13232 7700
rect 13252 7680 13264 7700
rect 13220 7642 13264 7680
rect 13336 7700 13378 7742
rect 13336 7680 13344 7700
rect 13364 7680 13378 7700
rect 13336 7642 13378 7680
rect 13428 7700 13472 7742
rect 13428 7680 13440 7700
rect 13460 7680 13472 7700
rect 13428 7642 13472 7680
rect 13549 7700 13591 7742
rect 13549 7680 13557 7700
rect 13577 7680 13591 7700
rect 13549 7642 13591 7680
rect 13641 7700 13685 7742
rect 16364 7805 16408 7847
rect 16458 7867 16500 7905
rect 16458 7847 16472 7867
rect 16492 7847 16500 7867
rect 16458 7805 16500 7847
rect 16577 7867 16621 7905
rect 16577 7847 16589 7867
rect 16609 7847 16621 7867
rect 16577 7805 16621 7847
rect 16671 7867 16713 7905
rect 16671 7847 16685 7867
rect 16705 7847 16713 7867
rect 16671 7805 16713 7847
rect 16785 7867 16829 7905
rect 16785 7847 16797 7867
rect 16817 7847 16829 7867
rect 16785 7805 16829 7847
rect 16879 7867 16921 7905
rect 16879 7847 16893 7867
rect 16913 7847 16921 7867
rect 16879 7805 16921 7847
rect 16995 7867 17037 7905
rect 16995 7847 17003 7867
rect 17023 7847 17037 7867
rect 16995 7805 17037 7847
rect 17087 7874 17132 7905
rect 17087 7867 17131 7874
rect 17087 7847 17099 7867
rect 17119 7847 17131 7867
rect 17087 7805 17131 7847
rect 13641 7680 13653 7700
rect 13673 7680 13685 7700
rect 13641 7642 13685 7680
rect 17974 7741 18018 7783
rect 17974 7721 17986 7741
rect 18006 7721 18018 7741
rect 17974 7714 18018 7721
rect 17973 7683 18018 7714
rect 18068 7741 18110 7783
rect 18068 7721 18082 7741
rect 18102 7721 18110 7741
rect 18068 7683 18110 7721
rect 18184 7741 18226 7783
rect 18184 7721 18192 7741
rect 18212 7721 18226 7741
rect 18184 7683 18226 7721
rect 18276 7741 18320 7783
rect 18276 7721 18288 7741
rect 18308 7721 18320 7741
rect 18276 7683 18320 7721
rect 18392 7741 18434 7783
rect 18392 7721 18400 7741
rect 18420 7721 18434 7741
rect 18392 7683 18434 7721
rect 18484 7741 18528 7783
rect 18484 7721 18496 7741
rect 18516 7721 18528 7741
rect 18484 7683 18528 7721
rect 18605 7741 18647 7783
rect 18605 7721 18613 7741
rect 18633 7721 18647 7741
rect 18605 7683 18647 7721
rect 18697 7741 18741 7783
rect 18697 7721 18709 7741
rect 18729 7721 18741 7741
rect 18697 7683 18741 7721
rect 6117 7490 6161 7532
rect 8881 7492 8925 7534
rect 4548 7431 4560 7451
rect 4580 7431 4592 7451
rect 4548 7393 4592 7431
rect 8881 7472 8893 7492
rect 8913 7472 8925 7492
rect 8881 7465 8925 7472
rect 8880 7434 8925 7465
rect 8975 7492 9017 7534
rect 8975 7472 8989 7492
rect 9009 7472 9017 7492
rect 8975 7434 9017 7472
rect 9091 7492 9133 7534
rect 9091 7472 9099 7492
rect 9119 7472 9133 7492
rect 9091 7434 9133 7472
rect 9183 7492 9227 7534
rect 9183 7472 9195 7492
rect 9215 7472 9227 7492
rect 9183 7434 9227 7472
rect 9299 7492 9341 7534
rect 9299 7472 9307 7492
rect 9327 7472 9341 7492
rect 9299 7434 9341 7472
rect 9391 7492 9435 7534
rect 9391 7472 9403 7492
rect 9423 7472 9435 7492
rect 9391 7434 9435 7472
rect 9512 7492 9554 7534
rect 9512 7472 9520 7492
rect 9540 7472 9554 7492
rect 9512 7434 9554 7472
rect 9604 7492 9648 7534
rect 9604 7472 9616 7492
rect 9636 7472 9648 7492
rect 10369 7516 10413 7554
rect 10369 7496 10381 7516
rect 10401 7496 10413 7516
rect 9604 7434 9648 7472
rect 10369 7454 10413 7496
rect 10463 7516 10505 7554
rect 10463 7496 10477 7516
rect 10497 7496 10505 7516
rect 10463 7454 10505 7496
rect 10582 7516 10626 7554
rect 10582 7496 10594 7516
rect 10614 7496 10626 7516
rect 10582 7454 10626 7496
rect 10676 7516 10718 7554
rect 10676 7496 10690 7516
rect 10710 7496 10718 7516
rect 10676 7454 10718 7496
rect 10790 7516 10834 7554
rect 10790 7496 10802 7516
rect 10822 7496 10834 7516
rect 10790 7454 10834 7496
rect 10884 7516 10926 7554
rect 10884 7496 10898 7516
rect 10918 7496 10926 7516
rect 10884 7454 10926 7496
rect 11000 7516 11042 7554
rect 11000 7496 11008 7516
rect 11028 7496 11042 7516
rect 11000 7454 11042 7496
rect 11092 7523 11137 7554
rect 11092 7516 11136 7523
rect 11092 7496 11104 7516
rect 11124 7496 11136 7516
rect 15425 7557 15469 7595
rect 15425 7537 15437 7557
rect 15457 7537 15469 7557
rect 11092 7454 11136 7496
rect 13856 7456 13900 7498
rect 13856 7436 13868 7456
rect 13888 7436 13900 7456
rect 13856 7429 13900 7436
rect 13855 7398 13900 7429
rect 13950 7456 13992 7498
rect 13950 7436 13964 7456
rect 13984 7436 13992 7456
rect 13950 7398 13992 7436
rect 14066 7456 14108 7498
rect 14066 7436 14074 7456
rect 14094 7436 14108 7456
rect 14066 7398 14108 7436
rect 14158 7456 14202 7498
rect 14158 7436 14170 7456
rect 14190 7436 14202 7456
rect 14158 7398 14202 7436
rect 14274 7456 14316 7498
rect 14274 7436 14282 7456
rect 14302 7436 14316 7456
rect 14274 7398 14316 7436
rect 14366 7456 14410 7498
rect 14366 7436 14378 7456
rect 14398 7436 14410 7456
rect 14366 7398 14410 7436
rect 14487 7456 14529 7498
rect 14487 7436 14495 7456
rect 14515 7436 14529 7456
rect 14487 7398 14529 7436
rect 14579 7456 14623 7498
rect 15425 7495 15469 7537
rect 15519 7557 15561 7595
rect 15519 7537 15533 7557
rect 15553 7537 15561 7557
rect 15519 7495 15561 7537
rect 15638 7557 15682 7595
rect 15638 7537 15650 7557
rect 15670 7537 15682 7557
rect 15638 7495 15682 7537
rect 15732 7557 15774 7595
rect 15732 7537 15746 7557
rect 15766 7537 15774 7557
rect 15732 7495 15774 7537
rect 15846 7557 15890 7595
rect 15846 7537 15858 7557
rect 15878 7537 15890 7557
rect 15846 7495 15890 7537
rect 15940 7557 15982 7595
rect 15940 7537 15954 7557
rect 15974 7537 15982 7557
rect 15940 7495 15982 7537
rect 16056 7557 16098 7595
rect 16056 7537 16064 7557
rect 16084 7537 16098 7557
rect 16056 7495 16098 7537
rect 16148 7564 16193 7595
rect 16148 7557 16192 7564
rect 16148 7537 16160 7557
rect 16180 7537 16192 7557
rect 16148 7495 16192 7537
rect 18912 7497 18956 7539
rect 14579 7436 14591 7456
rect 14611 7436 14623 7456
rect 14579 7398 14623 7436
rect 18912 7477 18924 7497
rect 18944 7477 18956 7497
rect 18912 7470 18956 7477
rect 18911 7439 18956 7470
rect 19006 7497 19048 7539
rect 19006 7477 19020 7497
rect 19040 7477 19048 7497
rect 19006 7439 19048 7477
rect 19122 7497 19164 7539
rect 19122 7477 19130 7497
rect 19150 7477 19164 7497
rect 19122 7439 19164 7477
rect 19214 7497 19258 7539
rect 19214 7477 19226 7497
rect 19246 7477 19258 7497
rect 19214 7439 19258 7477
rect 19330 7497 19372 7539
rect 19330 7477 19338 7497
rect 19358 7477 19372 7497
rect 19330 7439 19372 7477
rect 19422 7497 19466 7539
rect 19422 7477 19434 7497
rect 19454 7477 19466 7497
rect 19422 7439 19466 7477
rect 19543 7497 19585 7539
rect 19543 7477 19551 7497
rect 19571 7477 19585 7497
rect 19543 7439 19585 7477
rect 19635 7497 19679 7539
rect 19635 7477 19647 7497
rect 19667 7477 19679 7497
rect 19635 7439 19679 7477
rect 1387 7242 1431 7280
rect 1387 7222 1399 7242
rect 1419 7222 1431 7242
rect 1387 7180 1431 7222
rect 1481 7242 1523 7280
rect 1481 7222 1495 7242
rect 1515 7222 1523 7242
rect 1481 7180 1523 7222
rect 1600 7242 1644 7280
rect 1600 7222 1612 7242
rect 1632 7222 1644 7242
rect 1600 7180 1644 7222
rect 1694 7242 1736 7280
rect 1694 7222 1708 7242
rect 1728 7222 1736 7242
rect 1694 7180 1736 7222
rect 1808 7242 1852 7280
rect 1808 7222 1820 7242
rect 1840 7222 1852 7242
rect 1808 7180 1852 7222
rect 1902 7242 1944 7280
rect 1902 7222 1916 7242
rect 1936 7222 1944 7242
rect 1902 7180 1944 7222
rect 2018 7242 2060 7280
rect 2018 7222 2026 7242
rect 2046 7222 2060 7242
rect 2018 7180 2060 7222
rect 2110 7249 2155 7280
rect 2110 7242 2154 7249
rect 2110 7222 2122 7242
rect 2142 7222 2154 7242
rect 2110 7180 2154 7222
rect 6443 7283 6487 7321
rect 6443 7263 6455 7283
rect 6475 7263 6487 7283
rect 6443 7221 6487 7263
rect 6537 7283 6579 7321
rect 6537 7263 6551 7283
rect 6571 7263 6579 7283
rect 6537 7221 6579 7263
rect 6656 7283 6700 7321
rect 6656 7263 6668 7283
rect 6688 7263 6700 7283
rect 6656 7221 6700 7263
rect 6750 7283 6792 7321
rect 6750 7263 6764 7283
rect 6784 7263 6792 7283
rect 6750 7221 6792 7263
rect 6864 7283 6908 7321
rect 6864 7263 6876 7283
rect 6896 7263 6908 7283
rect 6864 7221 6908 7263
rect 6958 7283 7000 7321
rect 6958 7263 6972 7283
rect 6992 7263 7000 7283
rect 6958 7221 7000 7263
rect 7074 7283 7116 7321
rect 7074 7263 7082 7283
rect 7102 7263 7116 7283
rect 7074 7221 7116 7263
rect 7166 7290 7211 7321
rect 7166 7283 7210 7290
rect 7166 7263 7178 7283
rect 7198 7263 7210 7283
rect 7166 7221 7210 7263
rect 2777 7171 2821 7213
rect 2777 7151 2789 7171
rect 2809 7151 2821 7171
rect 2777 7144 2821 7151
rect 2776 7113 2821 7144
rect 2871 7171 2913 7213
rect 2871 7151 2885 7171
rect 2905 7151 2913 7171
rect 2871 7113 2913 7151
rect 2987 7171 3029 7213
rect 2987 7151 2995 7171
rect 3015 7151 3029 7171
rect 2987 7113 3029 7151
rect 3079 7171 3123 7213
rect 3079 7151 3091 7171
rect 3111 7151 3123 7171
rect 3079 7113 3123 7151
rect 3195 7171 3237 7213
rect 3195 7151 3203 7171
rect 3223 7151 3237 7171
rect 3195 7113 3237 7151
rect 3287 7171 3331 7213
rect 3287 7151 3299 7171
rect 3319 7151 3331 7171
rect 3287 7113 3331 7151
rect 3408 7171 3450 7213
rect 3408 7151 3416 7171
rect 3436 7151 3450 7171
rect 3408 7113 3450 7151
rect 3500 7171 3544 7213
rect 3500 7151 3512 7171
rect 3532 7151 3544 7171
rect 3500 7113 3544 7151
rect 7833 7212 7877 7254
rect 7833 7192 7845 7212
rect 7865 7192 7877 7212
rect 7833 7185 7877 7192
rect 7832 7154 7877 7185
rect 7927 7212 7969 7254
rect 7927 7192 7941 7212
rect 7961 7192 7969 7212
rect 7927 7154 7969 7192
rect 8043 7212 8085 7254
rect 8043 7192 8051 7212
rect 8071 7192 8085 7212
rect 8043 7154 8085 7192
rect 8135 7212 8179 7254
rect 8135 7192 8147 7212
rect 8167 7192 8179 7212
rect 8135 7154 8179 7192
rect 8251 7212 8293 7254
rect 8251 7192 8259 7212
rect 8279 7192 8293 7212
rect 8251 7154 8293 7192
rect 8343 7212 8387 7254
rect 8343 7192 8355 7212
rect 8375 7192 8387 7212
rect 8343 7154 8387 7192
rect 8464 7212 8506 7254
rect 8464 7192 8472 7212
rect 8492 7192 8506 7212
rect 8464 7154 8506 7192
rect 8556 7212 8600 7254
rect 11418 7247 11462 7285
rect 8556 7192 8568 7212
rect 8588 7192 8600 7212
rect 11418 7227 11430 7247
rect 11450 7227 11462 7247
rect 8556 7154 8600 7192
rect 11418 7185 11462 7227
rect 11512 7247 11554 7285
rect 11512 7227 11526 7247
rect 11546 7227 11554 7247
rect 11512 7185 11554 7227
rect 11631 7247 11675 7285
rect 11631 7227 11643 7247
rect 11663 7227 11675 7247
rect 11631 7185 11675 7227
rect 11725 7247 11767 7285
rect 11725 7227 11739 7247
rect 11759 7227 11767 7247
rect 11725 7185 11767 7227
rect 11839 7247 11883 7285
rect 11839 7227 11851 7247
rect 11871 7227 11883 7247
rect 11839 7185 11883 7227
rect 11933 7247 11975 7285
rect 11933 7227 11947 7247
rect 11967 7227 11975 7247
rect 11933 7185 11975 7227
rect 12049 7247 12091 7285
rect 12049 7227 12057 7247
rect 12077 7227 12091 7247
rect 12049 7185 12091 7227
rect 12141 7254 12186 7285
rect 12141 7247 12185 7254
rect 12141 7227 12153 7247
rect 12173 7227 12185 7247
rect 12141 7185 12185 7227
rect 16474 7288 16518 7326
rect 16474 7268 16486 7288
rect 16506 7268 16518 7288
rect 16474 7226 16518 7268
rect 16568 7288 16610 7326
rect 16568 7268 16582 7288
rect 16602 7268 16610 7288
rect 16568 7226 16610 7268
rect 16687 7288 16731 7326
rect 16687 7268 16699 7288
rect 16719 7268 16731 7288
rect 16687 7226 16731 7268
rect 16781 7288 16823 7326
rect 16781 7268 16795 7288
rect 16815 7268 16823 7288
rect 16781 7226 16823 7268
rect 16895 7288 16939 7326
rect 16895 7268 16907 7288
rect 16927 7268 16939 7288
rect 16895 7226 16939 7268
rect 16989 7288 17031 7326
rect 16989 7268 17003 7288
rect 17023 7268 17031 7288
rect 16989 7226 17031 7268
rect 17105 7288 17147 7326
rect 17105 7268 17113 7288
rect 17133 7268 17147 7288
rect 17105 7226 17147 7268
rect 17197 7295 17242 7326
rect 17197 7288 17241 7295
rect 17197 7268 17209 7288
rect 17229 7268 17241 7288
rect 17197 7226 17241 7268
rect 12808 7176 12852 7218
rect 12808 7156 12820 7176
rect 12840 7156 12852 7176
rect 12808 7149 12852 7156
rect 12807 7118 12852 7149
rect 12902 7176 12944 7218
rect 12902 7156 12916 7176
rect 12936 7156 12944 7176
rect 12902 7118 12944 7156
rect 13018 7176 13060 7218
rect 13018 7156 13026 7176
rect 13046 7156 13060 7176
rect 13018 7118 13060 7156
rect 13110 7176 13154 7218
rect 13110 7156 13122 7176
rect 13142 7156 13154 7176
rect 13110 7118 13154 7156
rect 13226 7176 13268 7218
rect 13226 7156 13234 7176
rect 13254 7156 13268 7176
rect 13226 7118 13268 7156
rect 13318 7176 13362 7218
rect 13318 7156 13330 7176
rect 13350 7156 13362 7176
rect 13318 7118 13362 7156
rect 13439 7176 13481 7218
rect 13439 7156 13447 7176
rect 13467 7156 13481 7176
rect 13439 7118 13481 7156
rect 13531 7176 13575 7218
rect 13531 7156 13543 7176
rect 13563 7156 13575 7176
rect 13531 7118 13575 7156
rect 17864 7217 17908 7259
rect 17864 7197 17876 7217
rect 17896 7197 17908 7217
rect 17864 7190 17908 7197
rect 17863 7159 17908 7190
rect 17958 7217 18000 7259
rect 17958 7197 17972 7217
rect 17992 7197 18000 7217
rect 17958 7159 18000 7197
rect 18074 7217 18116 7259
rect 18074 7197 18082 7217
rect 18102 7197 18116 7217
rect 18074 7159 18116 7197
rect 18166 7217 18210 7259
rect 18166 7197 18178 7217
rect 18198 7197 18210 7217
rect 18166 7159 18210 7197
rect 18282 7217 18324 7259
rect 18282 7197 18290 7217
rect 18310 7197 18324 7217
rect 18282 7159 18324 7197
rect 18374 7217 18418 7259
rect 18374 7197 18386 7217
rect 18406 7197 18418 7217
rect 18374 7159 18418 7197
rect 18495 7217 18537 7259
rect 18495 7197 18503 7217
rect 18523 7197 18537 7217
rect 18495 7159 18537 7197
rect 18587 7217 18631 7259
rect 18587 7197 18599 7217
rect 18619 7197 18631 7217
rect 18587 7159 18631 7197
rect 339 6962 383 7000
rect 339 6942 351 6962
rect 371 6942 383 6962
rect 339 6900 383 6942
rect 433 6962 475 7000
rect 433 6942 447 6962
rect 467 6942 475 6962
rect 433 6900 475 6942
rect 552 6962 596 7000
rect 552 6942 564 6962
rect 584 6942 596 6962
rect 552 6900 596 6942
rect 646 6962 688 7000
rect 646 6942 660 6962
rect 680 6942 688 6962
rect 646 6900 688 6942
rect 760 6962 804 7000
rect 760 6942 772 6962
rect 792 6942 804 6962
rect 760 6900 804 6942
rect 854 6962 896 7000
rect 854 6942 868 6962
rect 888 6942 896 6962
rect 854 6900 896 6942
rect 970 6962 1012 7000
rect 970 6942 978 6962
rect 998 6942 1012 6962
rect 970 6900 1012 6942
rect 1062 6969 1107 7000
rect 1062 6962 1106 6969
rect 1062 6942 1074 6962
rect 1094 6942 1106 6962
rect 5395 7003 5439 7041
rect 5395 6983 5407 7003
rect 5427 6983 5439 7003
rect 1062 6900 1106 6942
rect 3826 6902 3870 6944
rect 3826 6882 3838 6902
rect 3858 6882 3870 6902
rect 3826 6875 3870 6882
rect 3825 6844 3870 6875
rect 3920 6902 3962 6944
rect 3920 6882 3934 6902
rect 3954 6882 3962 6902
rect 3920 6844 3962 6882
rect 4036 6902 4078 6944
rect 4036 6882 4044 6902
rect 4064 6882 4078 6902
rect 4036 6844 4078 6882
rect 4128 6902 4172 6944
rect 4128 6882 4140 6902
rect 4160 6882 4172 6902
rect 4128 6844 4172 6882
rect 4244 6902 4286 6944
rect 4244 6882 4252 6902
rect 4272 6882 4286 6902
rect 4244 6844 4286 6882
rect 4336 6902 4380 6944
rect 4336 6882 4348 6902
rect 4368 6882 4380 6902
rect 4336 6844 4380 6882
rect 4457 6902 4499 6944
rect 4457 6882 4465 6902
rect 4485 6882 4499 6902
rect 4457 6844 4499 6882
rect 4549 6902 4593 6944
rect 5395 6941 5439 6983
rect 5489 7003 5531 7041
rect 5489 6983 5503 7003
rect 5523 6983 5531 7003
rect 5489 6941 5531 6983
rect 5608 7003 5652 7041
rect 5608 6983 5620 7003
rect 5640 6983 5652 7003
rect 5608 6941 5652 6983
rect 5702 7003 5744 7041
rect 5702 6983 5716 7003
rect 5736 6983 5744 7003
rect 5702 6941 5744 6983
rect 5816 7003 5860 7041
rect 5816 6983 5828 7003
rect 5848 6983 5860 7003
rect 5816 6941 5860 6983
rect 5910 7003 5952 7041
rect 5910 6983 5924 7003
rect 5944 6983 5952 7003
rect 5910 6941 5952 6983
rect 6026 7003 6068 7041
rect 6026 6983 6034 7003
rect 6054 6983 6068 7003
rect 6026 6941 6068 6983
rect 6118 7010 6163 7041
rect 6118 7003 6162 7010
rect 6118 6983 6130 7003
rect 6150 6983 6162 7003
rect 6118 6941 6162 6983
rect 8882 6943 8926 6985
rect 4549 6882 4561 6902
rect 4581 6882 4593 6902
rect 4549 6844 4593 6882
rect 8882 6923 8894 6943
rect 8914 6923 8926 6943
rect 8882 6916 8926 6923
rect 8881 6885 8926 6916
rect 8976 6943 9018 6985
rect 8976 6923 8990 6943
rect 9010 6923 9018 6943
rect 8976 6885 9018 6923
rect 9092 6943 9134 6985
rect 9092 6923 9100 6943
rect 9120 6923 9134 6943
rect 9092 6885 9134 6923
rect 9184 6943 9228 6985
rect 9184 6923 9196 6943
rect 9216 6923 9228 6943
rect 9184 6885 9228 6923
rect 9300 6943 9342 6985
rect 9300 6923 9308 6943
rect 9328 6923 9342 6943
rect 9300 6885 9342 6923
rect 9392 6943 9436 6985
rect 9392 6923 9404 6943
rect 9424 6923 9436 6943
rect 9392 6885 9436 6923
rect 9513 6943 9555 6985
rect 9513 6923 9521 6943
rect 9541 6923 9555 6943
rect 9513 6885 9555 6923
rect 9605 6943 9649 6985
rect 10370 6967 10414 7005
rect 9605 6923 9617 6943
rect 9637 6923 9649 6943
rect 9605 6885 9649 6923
rect 10370 6947 10382 6967
rect 10402 6947 10414 6967
rect 10370 6905 10414 6947
rect 10464 6967 10506 7005
rect 10464 6947 10478 6967
rect 10498 6947 10506 6967
rect 10464 6905 10506 6947
rect 10583 6967 10627 7005
rect 10583 6947 10595 6967
rect 10615 6947 10627 6967
rect 10583 6905 10627 6947
rect 10677 6967 10719 7005
rect 10677 6947 10691 6967
rect 10711 6947 10719 6967
rect 10677 6905 10719 6947
rect 10791 6967 10835 7005
rect 10791 6947 10803 6967
rect 10823 6947 10835 6967
rect 10791 6905 10835 6947
rect 10885 6967 10927 7005
rect 10885 6947 10899 6967
rect 10919 6947 10927 6967
rect 10885 6905 10927 6947
rect 11001 6967 11043 7005
rect 11001 6947 11009 6967
rect 11029 6947 11043 6967
rect 11001 6905 11043 6947
rect 11093 6974 11138 7005
rect 11093 6967 11137 6974
rect 11093 6947 11105 6967
rect 11125 6947 11137 6967
rect 15426 7008 15470 7046
rect 15426 6988 15438 7008
rect 15458 6988 15470 7008
rect 11093 6905 11137 6947
rect 13857 6907 13901 6949
rect 1277 6718 1321 6756
rect 1277 6698 1289 6718
rect 1309 6698 1321 6718
rect 1277 6656 1321 6698
rect 1371 6718 1413 6756
rect 1371 6698 1385 6718
rect 1405 6698 1413 6718
rect 1371 6656 1413 6698
rect 1490 6718 1534 6756
rect 1490 6698 1502 6718
rect 1522 6698 1534 6718
rect 1490 6656 1534 6698
rect 1584 6718 1626 6756
rect 1584 6698 1598 6718
rect 1618 6698 1626 6718
rect 1584 6656 1626 6698
rect 1698 6718 1742 6756
rect 1698 6698 1710 6718
rect 1730 6698 1742 6718
rect 1698 6656 1742 6698
rect 1792 6718 1834 6756
rect 1792 6698 1806 6718
rect 1826 6698 1834 6718
rect 1792 6656 1834 6698
rect 1908 6718 1950 6756
rect 1908 6698 1916 6718
rect 1936 6698 1950 6718
rect 1908 6656 1950 6698
rect 2000 6725 2045 6756
rect 2000 6718 2044 6725
rect 2000 6698 2012 6718
rect 2032 6698 2044 6718
rect 2000 6656 2044 6698
rect 6333 6759 6377 6797
rect 6333 6739 6345 6759
rect 6365 6739 6377 6759
rect 2887 6592 2931 6634
rect 2887 6572 2899 6592
rect 2919 6572 2931 6592
rect 2887 6565 2931 6572
rect 2886 6534 2931 6565
rect 2981 6592 3023 6634
rect 2981 6572 2995 6592
rect 3015 6572 3023 6592
rect 2981 6534 3023 6572
rect 3097 6592 3139 6634
rect 3097 6572 3105 6592
rect 3125 6572 3139 6592
rect 3097 6534 3139 6572
rect 3189 6592 3233 6634
rect 3189 6572 3201 6592
rect 3221 6572 3233 6592
rect 3189 6534 3233 6572
rect 3305 6592 3347 6634
rect 3305 6572 3313 6592
rect 3333 6572 3347 6592
rect 3305 6534 3347 6572
rect 3397 6592 3441 6634
rect 3397 6572 3409 6592
rect 3429 6572 3441 6592
rect 3397 6534 3441 6572
rect 3518 6592 3560 6634
rect 3518 6572 3526 6592
rect 3546 6572 3560 6592
rect 3518 6534 3560 6572
rect 3610 6592 3654 6634
rect 6333 6697 6377 6739
rect 6427 6759 6469 6797
rect 6427 6739 6441 6759
rect 6461 6739 6469 6759
rect 6427 6697 6469 6739
rect 6546 6759 6590 6797
rect 6546 6739 6558 6759
rect 6578 6739 6590 6759
rect 6546 6697 6590 6739
rect 6640 6759 6682 6797
rect 6640 6739 6654 6759
rect 6674 6739 6682 6759
rect 6640 6697 6682 6739
rect 6754 6759 6798 6797
rect 6754 6739 6766 6759
rect 6786 6739 6798 6759
rect 6754 6697 6798 6739
rect 6848 6759 6890 6797
rect 6848 6739 6862 6759
rect 6882 6739 6890 6759
rect 6848 6697 6890 6739
rect 6964 6759 7006 6797
rect 6964 6739 6972 6759
rect 6992 6739 7006 6759
rect 6964 6697 7006 6739
rect 7056 6766 7101 6797
rect 13857 6887 13869 6907
rect 13889 6887 13901 6907
rect 13857 6880 13901 6887
rect 7056 6759 7100 6766
rect 7056 6739 7068 6759
rect 7088 6739 7100 6759
rect 13856 6849 13901 6880
rect 13951 6907 13993 6949
rect 13951 6887 13965 6907
rect 13985 6887 13993 6907
rect 13951 6849 13993 6887
rect 14067 6907 14109 6949
rect 14067 6887 14075 6907
rect 14095 6887 14109 6907
rect 14067 6849 14109 6887
rect 14159 6907 14203 6949
rect 14159 6887 14171 6907
rect 14191 6887 14203 6907
rect 14159 6849 14203 6887
rect 14275 6907 14317 6949
rect 14275 6887 14283 6907
rect 14303 6887 14317 6907
rect 14275 6849 14317 6887
rect 14367 6907 14411 6949
rect 14367 6887 14379 6907
rect 14399 6887 14411 6907
rect 14367 6849 14411 6887
rect 14488 6907 14530 6949
rect 14488 6887 14496 6907
rect 14516 6887 14530 6907
rect 14488 6849 14530 6887
rect 14580 6907 14624 6949
rect 15426 6946 15470 6988
rect 15520 7008 15562 7046
rect 15520 6988 15534 7008
rect 15554 6988 15562 7008
rect 15520 6946 15562 6988
rect 15639 7008 15683 7046
rect 15639 6988 15651 7008
rect 15671 6988 15683 7008
rect 15639 6946 15683 6988
rect 15733 7008 15775 7046
rect 15733 6988 15747 7008
rect 15767 6988 15775 7008
rect 15733 6946 15775 6988
rect 15847 7008 15891 7046
rect 15847 6988 15859 7008
rect 15879 6988 15891 7008
rect 15847 6946 15891 6988
rect 15941 7008 15983 7046
rect 15941 6988 15955 7008
rect 15975 6988 15983 7008
rect 15941 6946 15983 6988
rect 16057 7008 16099 7046
rect 16057 6988 16065 7008
rect 16085 6988 16099 7008
rect 16057 6946 16099 6988
rect 16149 7015 16194 7046
rect 16149 7008 16193 7015
rect 16149 6988 16161 7008
rect 16181 6988 16193 7008
rect 16149 6946 16193 6988
rect 18913 6948 18957 6990
rect 14580 6887 14592 6907
rect 14612 6887 14624 6907
rect 14580 6849 14624 6887
rect 18913 6928 18925 6948
rect 18945 6928 18957 6948
rect 18913 6921 18957 6928
rect 18912 6890 18957 6921
rect 19007 6948 19049 6990
rect 19007 6928 19021 6948
rect 19041 6928 19049 6948
rect 19007 6890 19049 6928
rect 19123 6948 19165 6990
rect 19123 6928 19131 6948
rect 19151 6928 19165 6948
rect 19123 6890 19165 6928
rect 19215 6948 19259 6990
rect 19215 6928 19227 6948
rect 19247 6928 19259 6948
rect 19215 6890 19259 6928
rect 19331 6948 19373 6990
rect 19331 6928 19339 6948
rect 19359 6928 19373 6948
rect 19331 6890 19373 6928
rect 19423 6948 19467 6990
rect 19423 6928 19435 6948
rect 19455 6928 19467 6948
rect 19423 6890 19467 6928
rect 19544 6948 19586 6990
rect 19544 6928 19552 6948
rect 19572 6928 19586 6948
rect 19544 6890 19586 6928
rect 19636 6948 19680 6990
rect 19636 6928 19648 6948
rect 19668 6928 19680 6948
rect 19636 6890 19680 6928
rect 7056 6697 7100 6739
rect 3610 6572 3622 6592
rect 3642 6572 3654 6592
rect 3610 6534 3654 6572
rect 7943 6633 7987 6675
rect 7943 6613 7955 6633
rect 7975 6613 7987 6633
rect 7943 6606 7987 6613
rect 7942 6575 7987 6606
rect 8037 6633 8079 6675
rect 8037 6613 8051 6633
rect 8071 6613 8079 6633
rect 8037 6575 8079 6613
rect 8153 6633 8195 6675
rect 8153 6613 8161 6633
rect 8181 6613 8195 6633
rect 8153 6575 8195 6613
rect 8245 6633 8289 6675
rect 8245 6613 8257 6633
rect 8277 6613 8289 6633
rect 8245 6575 8289 6613
rect 8361 6633 8403 6675
rect 8361 6613 8369 6633
rect 8389 6613 8403 6633
rect 8361 6575 8403 6613
rect 8453 6633 8497 6675
rect 8453 6613 8465 6633
rect 8485 6613 8497 6633
rect 8453 6575 8497 6613
rect 8574 6633 8616 6675
rect 8574 6613 8582 6633
rect 8602 6613 8616 6633
rect 8574 6575 8616 6613
rect 8666 6633 8710 6675
rect 11308 6723 11352 6761
rect 11308 6703 11320 6723
rect 11340 6703 11352 6723
rect 8666 6613 8678 6633
rect 8698 6613 8710 6633
rect 8666 6575 8710 6613
rect 11308 6661 11352 6703
rect 11402 6723 11444 6761
rect 11402 6703 11416 6723
rect 11436 6703 11444 6723
rect 11402 6661 11444 6703
rect 11521 6723 11565 6761
rect 11521 6703 11533 6723
rect 11553 6703 11565 6723
rect 11521 6661 11565 6703
rect 11615 6723 11657 6761
rect 11615 6703 11629 6723
rect 11649 6703 11657 6723
rect 11615 6661 11657 6703
rect 11729 6723 11773 6761
rect 11729 6703 11741 6723
rect 11761 6703 11773 6723
rect 11729 6661 11773 6703
rect 11823 6723 11865 6761
rect 11823 6703 11837 6723
rect 11857 6703 11865 6723
rect 11823 6661 11865 6703
rect 11939 6723 11981 6761
rect 11939 6703 11947 6723
rect 11967 6703 11981 6723
rect 11939 6661 11981 6703
rect 12031 6730 12076 6761
rect 12031 6723 12075 6730
rect 12031 6703 12043 6723
rect 12063 6703 12075 6723
rect 12031 6661 12075 6703
rect 16364 6764 16408 6802
rect 16364 6744 16376 6764
rect 16396 6744 16408 6764
rect 12918 6597 12962 6639
rect 338 6408 382 6446
rect 338 6388 350 6408
rect 370 6388 382 6408
rect 338 6346 382 6388
rect 432 6408 474 6446
rect 432 6388 446 6408
rect 466 6388 474 6408
rect 432 6346 474 6388
rect 551 6408 595 6446
rect 551 6388 563 6408
rect 583 6388 595 6408
rect 551 6346 595 6388
rect 645 6408 687 6446
rect 645 6388 659 6408
rect 679 6388 687 6408
rect 645 6346 687 6388
rect 759 6408 803 6446
rect 759 6388 771 6408
rect 791 6388 803 6408
rect 759 6346 803 6388
rect 853 6408 895 6446
rect 853 6388 867 6408
rect 887 6388 895 6408
rect 853 6346 895 6388
rect 969 6408 1011 6446
rect 969 6388 977 6408
rect 997 6388 1011 6408
rect 969 6346 1011 6388
rect 1061 6415 1106 6446
rect 1061 6408 1105 6415
rect 1061 6388 1073 6408
rect 1093 6388 1105 6408
rect 5394 6449 5438 6487
rect 5394 6429 5406 6449
rect 5426 6429 5438 6449
rect 1061 6346 1105 6388
rect 3825 6348 3869 6390
rect 3825 6328 3837 6348
rect 3857 6328 3869 6348
rect 3825 6321 3869 6328
rect 3824 6290 3869 6321
rect 3919 6348 3961 6390
rect 3919 6328 3933 6348
rect 3953 6328 3961 6348
rect 3919 6290 3961 6328
rect 4035 6348 4077 6390
rect 4035 6328 4043 6348
rect 4063 6328 4077 6348
rect 4035 6290 4077 6328
rect 4127 6348 4171 6390
rect 4127 6328 4139 6348
rect 4159 6328 4171 6348
rect 4127 6290 4171 6328
rect 4243 6348 4285 6390
rect 4243 6328 4251 6348
rect 4271 6328 4285 6348
rect 4243 6290 4285 6328
rect 4335 6348 4379 6390
rect 4335 6328 4347 6348
rect 4367 6328 4379 6348
rect 4335 6290 4379 6328
rect 4456 6348 4498 6390
rect 4456 6328 4464 6348
rect 4484 6328 4498 6348
rect 4456 6290 4498 6328
rect 4548 6348 4592 6390
rect 5394 6387 5438 6429
rect 5488 6449 5530 6487
rect 5488 6429 5502 6449
rect 5522 6429 5530 6449
rect 5488 6387 5530 6429
rect 5607 6449 5651 6487
rect 5607 6429 5619 6449
rect 5639 6429 5651 6449
rect 5607 6387 5651 6429
rect 5701 6449 5743 6487
rect 5701 6429 5715 6449
rect 5735 6429 5743 6449
rect 5701 6387 5743 6429
rect 5815 6449 5859 6487
rect 5815 6429 5827 6449
rect 5847 6429 5859 6449
rect 5815 6387 5859 6429
rect 5909 6449 5951 6487
rect 5909 6429 5923 6449
rect 5943 6429 5951 6449
rect 5909 6387 5951 6429
rect 6025 6449 6067 6487
rect 6025 6429 6033 6449
rect 6053 6429 6067 6449
rect 6025 6387 6067 6429
rect 6117 6456 6162 6487
rect 12918 6577 12930 6597
rect 12950 6577 12962 6597
rect 12918 6570 12962 6577
rect 6117 6449 6161 6456
rect 6117 6429 6129 6449
rect 6149 6429 6161 6449
rect 12917 6539 12962 6570
rect 13012 6597 13054 6639
rect 13012 6577 13026 6597
rect 13046 6577 13054 6597
rect 13012 6539 13054 6577
rect 13128 6597 13170 6639
rect 13128 6577 13136 6597
rect 13156 6577 13170 6597
rect 13128 6539 13170 6577
rect 13220 6597 13264 6639
rect 13220 6577 13232 6597
rect 13252 6577 13264 6597
rect 13220 6539 13264 6577
rect 13336 6597 13378 6639
rect 13336 6577 13344 6597
rect 13364 6577 13378 6597
rect 13336 6539 13378 6577
rect 13428 6597 13472 6639
rect 13428 6577 13440 6597
rect 13460 6577 13472 6597
rect 13428 6539 13472 6577
rect 13549 6597 13591 6639
rect 13549 6577 13557 6597
rect 13577 6577 13591 6597
rect 13549 6539 13591 6577
rect 13641 6597 13685 6639
rect 16364 6702 16408 6744
rect 16458 6764 16500 6802
rect 16458 6744 16472 6764
rect 16492 6744 16500 6764
rect 16458 6702 16500 6744
rect 16577 6764 16621 6802
rect 16577 6744 16589 6764
rect 16609 6744 16621 6764
rect 16577 6702 16621 6744
rect 16671 6764 16713 6802
rect 16671 6744 16685 6764
rect 16705 6744 16713 6764
rect 16671 6702 16713 6744
rect 16785 6764 16829 6802
rect 16785 6744 16797 6764
rect 16817 6744 16829 6764
rect 16785 6702 16829 6744
rect 16879 6764 16921 6802
rect 16879 6744 16893 6764
rect 16913 6744 16921 6764
rect 16879 6702 16921 6744
rect 16995 6764 17037 6802
rect 16995 6744 17003 6764
rect 17023 6744 17037 6764
rect 16995 6702 17037 6744
rect 17087 6771 17132 6802
rect 17087 6764 17131 6771
rect 17087 6744 17099 6764
rect 17119 6744 17131 6764
rect 17087 6702 17131 6744
rect 13641 6577 13653 6597
rect 13673 6577 13685 6597
rect 13641 6539 13685 6577
rect 17974 6638 18018 6680
rect 17974 6618 17986 6638
rect 18006 6618 18018 6638
rect 17974 6611 18018 6618
rect 17973 6580 18018 6611
rect 18068 6638 18110 6680
rect 18068 6618 18082 6638
rect 18102 6618 18110 6638
rect 18068 6580 18110 6618
rect 18184 6638 18226 6680
rect 18184 6618 18192 6638
rect 18212 6618 18226 6638
rect 18184 6580 18226 6618
rect 18276 6638 18320 6680
rect 18276 6618 18288 6638
rect 18308 6618 18320 6638
rect 18276 6580 18320 6618
rect 18392 6638 18434 6680
rect 18392 6618 18400 6638
rect 18420 6618 18434 6638
rect 18392 6580 18434 6618
rect 18484 6638 18528 6680
rect 18484 6618 18496 6638
rect 18516 6618 18528 6638
rect 18484 6580 18528 6618
rect 18605 6638 18647 6680
rect 18605 6618 18613 6638
rect 18633 6618 18647 6638
rect 18605 6580 18647 6618
rect 18697 6638 18741 6680
rect 18697 6618 18709 6638
rect 18729 6618 18741 6638
rect 18697 6580 18741 6618
rect 6117 6387 6161 6429
rect 8881 6389 8925 6431
rect 4548 6328 4560 6348
rect 4580 6328 4592 6348
rect 4548 6290 4592 6328
rect 8881 6369 8893 6389
rect 8913 6369 8925 6389
rect 8881 6362 8925 6369
rect 8880 6331 8925 6362
rect 8975 6389 9017 6431
rect 8975 6369 8989 6389
rect 9009 6369 9017 6389
rect 8975 6331 9017 6369
rect 9091 6389 9133 6431
rect 9091 6369 9099 6389
rect 9119 6369 9133 6389
rect 9091 6331 9133 6369
rect 9183 6389 9227 6431
rect 9183 6369 9195 6389
rect 9215 6369 9227 6389
rect 9183 6331 9227 6369
rect 9299 6389 9341 6431
rect 9299 6369 9307 6389
rect 9327 6369 9341 6389
rect 9299 6331 9341 6369
rect 9391 6389 9435 6431
rect 9391 6369 9403 6389
rect 9423 6369 9435 6389
rect 9391 6331 9435 6369
rect 9512 6389 9554 6431
rect 9512 6369 9520 6389
rect 9540 6369 9554 6389
rect 9512 6331 9554 6369
rect 9604 6389 9648 6431
rect 9604 6369 9616 6389
rect 9636 6369 9648 6389
rect 10369 6413 10413 6451
rect 10369 6393 10381 6413
rect 10401 6393 10413 6413
rect 9604 6331 9648 6369
rect 10369 6351 10413 6393
rect 10463 6413 10505 6451
rect 10463 6393 10477 6413
rect 10497 6393 10505 6413
rect 10463 6351 10505 6393
rect 10582 6413 10626 6451
rect 10582 6393 10594 6413
rect 10614 6393 10626 6413
rect 10582 6351 10626 6393
rect 10676 6413 10718 6451
rect 10676 6393 10690 6413
rect 10710 6393 10718 6413
rect 10676 6351 10718 6393
rect 10790 6413 10834 6451
rect 10790 6393 10802 6413
rect 10822 6393 10834 6413
rect 10790 6351 10834 6393
rect 10884 6413 10926 6451
rect 10884 6393 10898 6413
rect 10918 6393 10926 6413
rect 10884 6351 10926 6393
rect 11000 6413 11042 6451
rect 11000 6393 11008 6413
rect 11028 6393 11042 6413
rect 11000 6351 11042 6393
rect 11092 6420 11137 6451
rect 11092 6413 11136 6420
rect 11092 6393 11104 6413
rect 11124 6393 11136 6413
rect 15425 6454 15469 6492
rect 15425 6434 15437 6454
rect 15457 6434 15469 6454
rect 11092 6351 11136 6393
rect 13856 6353 13900 6395
rect 13856 6333 13868 6353
rect 13888 6333 13900 6353
rect 13856 6326 13900 6333
rect 13855 6295 13900 6326
rect 13950 6353 13992 6395
rect 13950 6333 13964 6353
rect 13984 6333 13992 6353
rect 13950 6295 13992 6333
rect 14066 6353 14108 6395
rect 14066 6333 14074 6353
rect 14094 6333 14108 6353
rect 14066 6295 14108 6333
rect 14158 6353 14202 6395
rect 14158 6333 14170 6353
rect 14190 6333 14202 6353
rect 14158 6295 14202 6333
rect 14274 6353 14316 6395
rect 14274 6333 14282 6353
rect 14302 6333 14316 6353
rect 14274 6295 14316 6333
rect 14366 6353 14410 6395
rect 14366 6333 14378 6353
rect 14398 6333 14410 6353
rect 14366 6295 14410 6333
rect 14487 6353 14529 6395
rect 14487 6333 14495 6353
rect 14515 6333 14529 6353
rect 14487 6295 14529 6333
rect 14579 6353 14623 6395
rect 15425 6392 15469 6434
rect 15519 6454 15561 6492
rect 15519 6434 15533 6454
rect 15553 6434 15561 6454
rect 15519 6392 15561 6434
rect 15638 6454 15682 6492
rect 15638 6434 15650 6454
rect 15670 6434 15682 6454
rect 15638 6392 15682 6434
rect 15732 6454 15774 6492
rect 15732 6434 15746 6454
rect 15766 6434 15774 6454
rect 15732 6392 15774 6434
rect 15846 6454 15890 6492
rect 15846 6434 15858 6454
rect 15878 6434 15890 6454
rect 15846 6392 15890 6434
rect 15940 6454 15982 6492
rect 15940 6434 15954 6454
rect 15974 6434 15982 6454
rect 15940 6392 15982 6434
rect 16056 6454 16098 6492
rect 16056 6434 16064 6454
rect 16084 6434 16098 6454
rect 16056 6392 16098 6434
rect 16148 6461 16193 6492
rect 16148 6454 16192 6461
rect 16148 6434 16160 6454
rect 16180 6434 16192 6454
rect 16148 6392 16192 6434
rect 18912 6394 18956 6436
rect 14579 6333 14591 6353
rect 14611 6333 14623 6353
rect 14579 6295 14623 6333
rect 18912 6374 18924 6394
rect 18944 6374 18956 6394
rect 18912 6367 18956 6374
rect 18911 6336 18956 6367
rect 19006 6394 19048 6436
rect 19006 6374 19020 6394
rect 19040 6374 19048 6394
rect 19006 6336 19048 6374
rect 19122 6394 19164 6436
rect 19122 6374 19130 6394
rect 19150 6374 19164 6394
rect 19122 6336 19164 6374
rect 19214 6394 19258 6436
rect 19214 6374 19226 6394
rect 19246 6374 19258 6394
rect 19214 6336 19258 6374
rect 19330 6394 19372 6436
rect 19330 6374 19338 6394
rect 19358 6374 19372 6394
rect 19330 6336 19372 6374
rect 19422 6394 19466 6436
rect 19422 6374 19434 6394
rect 19454 6374 19466 6394
rect 19422 6336 19466 6374
rect 19543 6394 19585 6436
rect 19543 6374 19551 6394
rect 19571 6374 19585 6394
rect 19543 6336 19585 6374
rect 19635 6394 19679 6436
rect 19635 6374 19647 6394
rect 19667 6374 19679 6394
rect 19635 6336 19679 6374
rect 1418 6126 1462 6164
rect 1418 6106 1430 6126
rect 1450 6106 1462 6126
rect 1418 6064 1462 6106
rect 1512 6126 1554 6164
rect 1512 6106 1526 6126
rect 1546 6106 1554 6126
rect 1512 6064 1554 6106
rect 1631 6126 1675 6164
rect 1631 6106 1643 6126
rect 1663 6106 1675 6126
rect 1631 6064 1675 6106
rect 1725 6126 1767 6164
rect 1725 6106 1739 6126
rect 1759 6106 1767 6126
rect 1725 6064 1767 6106
rect 1839 6126 1883 6164
rect 1839 6106 1851 6126
rect 1871 6106 1883 6126
rect 1839 6064 1883 6106
rect 1933 6126 1975 6164
rect 1933 6106 1947 6126
rect 1967 6106 1975 6126
rect 1933 6064 1975 6106
rect 2049 6126 2091 6164
rect 2049 6106 2057 6126
rect 2077 6106 2091 6126
rect 2049 6064 2091 6106
rect 2141 6133 2186 6164
rect 2141 6126 2185 6133
rect 2141 6106 2153 6126
rect 2173 6106 2185 6126
rect 6474 6167 6518 6205
rect 6474 6147 6486 6167
rect 6506 6147 6518 6167
rect 2141 6064 2185 6106
rect 2747 6081 2791 6123
rect 2747 6061 2759 6081
rect 2779 6061 2791 6081
rect 2747 6054 2791 6061
rect 2746 6023 2791 6054
rect 2841 6081 2883 6123
rect 2841 6061 2855 6081
rect 2875 6061 2883 6081
rect 2841 6023 2883 6061
rect 2957 6081 2999 6123
rect 2957 6061 2965 6081
rect 2985 6061 2999 6081
rect 2957 6023 2999 6061
rect 3049 6081 3093 6123
rect 3049 6061 3061 6081
rect 3081 6061 3093 6081
rect 3049 6023 3093 6061
rect 3165 6081 3207 6123
rect 3165 6061 3173 6081
rect 3193 6061 3207 6081
rect 3165 6023 3207 6061
rect 3257 6081 3301 6123
rect 3257 6061 3269 6081
rect 3289 6061 3301 6081
rect 3257 6023 3301 6061
rect 3378 6081 3420 6123
rect 3378 6061 3386 6081
rect 3406 6061 3420 6081
rect 3378 6023 3420 6061
rect 3470 6081 3514 6123
rect 6474 6105 6518 6147
rect 6568 6167 6610 6205
rect 6568 6147 6582 6167
rect 6602 6147 6610 6167
rect 6568 6105 6610 6147
rect 6687 6167 6731 6205
rect 6687 6147 6699 6167
rect 6719 6147 6731 6167
rect 6687 6105 6731 6147
rect 6781 6167 6823 6205
rect 6781 6147 6795 6167
rect 6815 6147 6823 6167
rect 6781 6105 6823 6147
rect 6895 6167 6939 6205
rect 6895 6147 6907 6167
rect 6927 6147 6939 6167
rect 6895 6105 6939 6147
rect 6989 6167 7031 6205
rect 6989 6147 7003 6167
rect 7023 6147 7031 6167
rect 6989 6105 7031 6147
rect 7105 6167 7147 6205
rect 7105 6147 7113 6167
rect 7133 6147 7147 6167
rect 7105 6105 7147 6147
rect 7197 6174 7242 6205
rect 7197 6167 7241 6174
rect 7197 6147 7209 6167
rect 7229 6147 7241 6167
rect 7197 6105 7241 6147
rect 7803 6122 7847 6164
rect 3470 6061 3482 6081
rect 3502 6061 3514 6081
rect 3470 6023 3514 6061
rect 7803 6102 7815 6122
rect 7835 6102 7847 6122
rect 7803 6095 7847 6102
rect 7802 6064 7847 6095
rect 7897 6122 7939 6164
rect 7897 6102 7911 6122
rect 7931 6102 7939 6122
rect 7897 6064 7939 6102
rect 8013 6122 8055 6164
rect 8013 6102 8021 6122
rect 8041 6102 8055 6122
rect 8013 6064 8055 6102
rect 8105 6122 8149 6164
rect 8105 6102 8117 6122
rect 8137 6102 8149 6122
rect 8105 6064 8149 6102
rect 8221 6122 8263 6164
rect 8221 6102 8229 6122
rect 8249 6102 8263 6122
rect 8221 6064 8263 6102
rect 8313 6122 8357 6164
rect 8313 6102 8325 6122
rect 8345 6102 8357 6122
rect 8313 6064 8357 6102
rect 8434 6122 8476 6164
rect 8434 6102 8442 6122
rect 8462 6102 8476 6122
rect 8434 6064 8476 6102
rect 8526 6122 8570 6164
rect 8526 6102 8538 6122
rect 8558 6102 8570 6122
rect 8526 6064 8570 6102
rect 11449 6131 11493 6169
rect 11449 6111 11461 6131
rect 11481 6111 11493 6131
rect 11449 6069 11493 6111
rect 11543 6131 11585 6169
rect 11543 6111 11557 6131
rect 11577 6111 11585 6131
rect 11543 6069 11585 6111
rect 11662 6131 11706 6169
rect 11662 6111 11674 6131
rect 11694 6111 11706 6131
rect 11662 6069 11706 6111
rect 11756 6131 11798 6169
rect 11756 6111 11770 6131
rect 11790 6111 11798 6131
rect 11756 6069 11798 6111
rect 11870 6131 11914 6169
rect 11870 6111 11882 6131
rect 11902 6111 11914 6131
rect 11870 6069 11914 6111
rect 11964 6131 12006 6169
rect 11964 6111 11978 6131
rect 11998 6111 12006 6131
rect 11964 6069 12006 6111
rect 12080 6131 12122 6169
rect 12080 6111 12088 6131
rect 12108 6111 12122 6131
rect 12080 6069 12122 6111
rect 12172 6138 12217 6169
rect 12172 6131 12216 6138
rect 12172 6111 12184 6131
rect 12204 6111 12216 6131
rect 16505 6172 16549 6210
rect 16505 6152 16517 6172
rect 16537 6152 16549 6172
rect 12172 6069 12216 6111
rect 12778 6086 12822 6128
rect 12778 6066 12790 6086
rect 12810 6066 12822 6086
rect 12778 6059 12822 6066
rect 12777 6028 12822 6059
rect 12872 6086 12914 6128
rect 12872 6066 12886 6086
rect 12906 6066 12914 6086
rect 12872 6028 12914 6066
rect 12988 6086 13030 6128
rect 12988 6066 12996 6086
rect 13016 6066 13030 6086
rect 12988 6028 13030 6066
rect 13080 6086 13124 6128
rect 13080 6066 13092 6086
rect 13112 6066 13124 6086
rect 13080 6028 13124 6066
rect 13196 6086 13238 6128
rect 13196 6066 13204 6086
rect 13224 6066 13238 6086
rect 13196 6028 13238 6066
rect 13288 6086 13332 6128
rect 13288 6066 13300 6086
rect 13320 6066 13332 6086
rect 13288 6028 13332 6066
rect 13409 6086 13451 6128
rect 13409 6066 13417 6086
rect 13437 6066 13451 6086
rect 13409 6028 13451 6066
rect 13501 6086 13545 6128
rect 16505 6110 16549 6152
rect 16599 6172 16641 6210
rect 16599 6152 16613 6172
rect 16633 6152 16641 6172
rect 16599 6110 16641 6152
rect 16718 6172 16762 6210
rect 16718 6152 16730 6172
rect 16750 6152 16762 6172
rect 16718 6110 16762 6152
rect 16812 6172 16854 6210
rect 16812 6152 16826 6172
rect 16846 6152 16854 6172
rect 16812 6110 16854 6152
rect 16926 6172 16970 6210
rect 16926 6152 16938 6172
rect 16958 6152 16970 6172
rect 16926 6110 16970 6152
rect 17020 6172 17062 6210
rect 17020 6152 17034 6172
rect 17054 6152 17062 6172
rect 17020 6110 17062 6152
rect 17136 6172 17178 6210
rect 17136 6152 17144 6172
rect 17164 6152 17178 6172
rect 17136 6110 17178 6152
rect 17228 6179 17273 6210
rect 17228 6172 17272 6179
rect 17228 6152 17240 6172
rect 17260 6152 17272 6172
rect 17228 6110 17272 6152
rect 17834 6127 17878 6169
rect 13501 6066 13513 6086
rect 13533 6066 13545 6086
rect 13501 6028 13545 6066
rect 17834 6107 17846 6127
rect 17866 6107 17878 6127
rect 17834 6100 17878 6107
rect 17833 6069 17878 6100
rect 17928 6127 17970 6169
rect 17928 6107 17942 6127
rect 17962 6107 17970 6127
rect 17928 6069 17970 6107
rect 18044 6127 18086 6169
rect 18044 6107 18052 6127
rect 18072 6107 18086 6127
rect 18044 6069 18086 6107
rect 18136 6127 18180 6169
rect 18136 6107 18148 6127
rect 18168 6107 18180 6127
rect 18136 6069 18180 6107
rect 18252 6127 18294 6169
rect 18252 6107 18260 6127
rect 18280 6107 18294 6127
rect 18252 6069 18294 6107
rect 18344 6127 18388 6169
rect 18344 6107 18356 6127
rect 18376 6107 18388 6127
rect 18344 6069 18388 6107
rect 18465 6127 18507 6169
rect 18465 6107 18473 6127
rect 18493 6107 18507 6127
rect 18465 6069 18507 6107
rect 18557 6127 18601 6169
rect 18557 6107 18569 6127
rect 18589 6107 18601 6127
rect 18557 6069 18601 6107
rect 340 5859 384 5897
rect 340 5839 352 5859
rect 372 5839 384 5859
rect 340 5797 384 5839
rect 434 5859 476 5897
rect 434 5839 448 5859
rect 468 5839 476 5859
rect 434 5797 476 5839
rect 553 5859 597 5897
rect 553 5839 565 5859
rect 585 5839 597 5859
rect 553 5797 597 5839
rect 647 5859 689 5897
rect 647 5839 661 5859
rect 681 5839 689 5859
rect 647 5797 689 5839
rect 761 5859 805 5897
rect 761 5839 773 5859
rect 793 5839 805 5859
rect 761 5797 805 5839
rect 855 5859 897 5897
rect 855 5839 869 5859
rect 889 5839 897 5859
rect 855 5797 897 5839
rect 971 5859 1013 5897
rect 971 5839 979 5859
rect 999 5839 1013 5859
rect 971 5797 1013 5839
rect 1063 5866 1108 5897
rect 1063 5859 1107 5866
rect 1063 5839 1075 5859
rect 1095 5839 1107 5859
rect 5396 5900 5440 5938
rect 5396 5880 5408 5900
rect 5428 5880 5440 5900
rect 1063 5797 1107 5839
rect 3827 5799 3871 5841
rect 3827 5779 3839 5799
rect 3859 5779 3871 5799
rect 3827 5772 3871 5779
rect 3826 5741 3871 5772
rect 3921 5799 3963 5841
rect 3921 5779 3935 5799
rect 3955 5779 3963 5799
rect 3921 5741 3963 5779
rect 4037 5799 4079 5841
rect 4037 5779 4045 5799
rect 4065 5779 4079 5799
rect 4037 5741 4079 5779
rect 4129 5799 4173 5841
rect 4129 5779 4141 5799
rect 4161 5779 4173 5799
rect 4129 5741 4173 5779
rect 4245 5799 4287 5841
rect 4245 5779 4253 5799
rect 4273 5779 4287 5799
rect 4245 5741 4287 5779
rect 4337 5799 4381 5841
rect 4337 5779 4349 5799
rect 4369 5779 4381 5799
rect 4337 5741 4381 5779
rect 4458 5799 4500 5841
rect 4458 5779 4466 5799
rect 4486 5779 4500 5799
rect 4458 5741 4500 5779
rect 4550 5799 4594 5841
rect 5396 5838 5440 5880
rect 5490 5900 5532 5938
rect 5490 5880 5504 5900
rect 5524 5880 5532 5900
rect 5490 5838 5532 5880
rect 5609 5900 5653 5938
rect 5609 5880 5621 5900
rect 5641 5880 5653 5900
rect 5609 5838 5653 5880
rect 5703 5900 5745 5938
rect 5703 5880 5717 5900
rect 5737 5880 5745 5900
rect 5703 5838 5745 5880
rect 5817 5900 5861 5938
rect 5817 5880 5829 5900
rect 5849 5880 5861 5900
rect 5817 5838 5861 5880
rect 5911 5900 5953 5938
rect 5911 5880 5925 5900
rect 5945 5880 5953 5900
rect 5911 5838 5953 5880
rect 6027 5900 6069 5938
rect 6027 5880 6035 5900
rect 6055 5880 6069 5900
rect 6027 5838 6069 5880
rect 6119 5907 6164 5938
rect 6119 5900 6163 5907
rect 6119 5880 6131 5900
rect 6151 5880 6163 5900
rect 6119 5838 6163 5880
rect 8883 5840 8927 5882
rect 4550 5779 4562 5799
rect 4582 5779 4594 5799
rect 4550 5741 4594 5779
rect 8883 5820 8895 5840
rect 8915 5820 8927 5840
rect 8883 5813 8927 5820
rect 8882 5782 8927 5813
rect 8977 5840 9019 5882
rect 8977 5820 8991 5840
rect 9011 5820 9019 5840
rect 8977 5782 9019 5820
rect 9093 5840 9135 5882
rect 9093 5820 9101 5840
rect 9121 5820 9135 5840
rect 9093 5782 9135 5820
rect 9185 5840 9229 5882
rect 9185 5820 9197 5840
rect 9217 5820 9229 5840
rect 9185 5782 9229 5820
rect 9301 5840 9343 5882
rect 9301 5820 9309 5840
rect 9329 5820 9343 5840
rect 9301 5782 9343 5820
rect 9393 5840 9437 5882
rect 9393 5820 9405 5840
rect 9425 5820 9437 5840
rect 9393 5782 9437 5820
rect 9514 5840 9556 5882
rect 9514 5820 9522 5840
rect 9542 5820 9556 5840
rect 9514 5782 9556 5820
rect 9606 5840 9650 5882
rect 10371 5864 10415 5902
rect 9606 5820 9618 5840
rect 9638 5820 9650 5840
rect 9606 5782 9650 5820
rect 10371 5844 10383 5864
rect 10403 5844 10415 5864
rect 10371 5802 10415 5844
rect 10465 5864 10507 5902
rect 10465 5844 10479 5864
rect 10499 5844 10507 5864
rect 10465 5802 10507 5844
rect 10584 5864 10628 5902
rect 10584 5844 10596 5864
rect 10616 5844 10628 5864
rect 10584 5802 10628 5844
rect 10678 5864 10720 5902
rect 10678 5844 10692 5864
rect 10712 5844 10720 5864
rect 10678 5802 10720 5844
rect 10792 5864 10836 5902
rect 10792 5844 10804 5864
rect 10824 5844 10836 5864
rect 10792 5802 10836 5844
rect 10886 5864 10928 5902
rect 10886 5844 10900 5864
rect 10920 5844 10928 5864
rect 10886 5802 10928 5844
rect 11002 5864 11044 5902
rect 11002 5844 11010 5864
rect 11030 5844 11044 5864
rect 11002 5802 11044 5844
rect 11094 5871 11139 5902
rect 11094 5864 11138 5871
rect 11094 5844 11106 5864
rect 11126 5844 11138 5864
rect 15427 5905 15471 5943
rect 15427 5885 15439 5905
rect 15459 5885 15471 5905
rect 11094 5802 11138 5844
rect 13858 5804 13902 5846
rect 1278 5615 1322 5653
rect 1278 5595 1290 5615
rect 1310 5595 1322 5615
rect 1278 5553 1322 5595
rect 1372 5615 1414 5653
rect 1372 5595 1386 5615
rect 1406 5595 1414 5615
rect 1372 5553 1414 5595
rect 1491 5615 1535 5653
rect 1491 5595 1503 5615
rect 1523 5595 1535 5615
rect 1491 5553 1535 5595
rect 1585 5615 1627 5653
rect 1585 5595 1599 5615
rect 1619 5595 1627 5615
rect 1585 5553 1627 5595
rect 1699 5615 1743 5653
rect 1699 5595 1711 5615
rect 1731 5595 1743 5615
rect 1699 5553 1743 5595
rect 1793 5615 1835 5653
rect 1793 5595 1807 5615
rect 1827 5595 1835 5615
rect 1793 5553 1835 5595
rect 1909 5615 1951 5653
rect 1909 5595 1917 5615
rect 1937 5595 1951 5615
rect 1909 5553 1951 5595
rect 2001 5622 2046 5653
rect 2001 5615 2045 5622
rect 2001 5595 2013 5615
rect 2033 5595 2045 5615
rect 2001 5553 2045 5595
rect 6334 5656 6378 5694
rect 6334 5636 6346 5656
rect 6366 5636 6378 5656
rect 2888 5489 2932 5531
rect 2888 5469 2900 5489
rect 2920 5469 2932 5489
rect 2888 5462 2932 5469
rect 2887 5431 2932 5462
rect 2982 5489 3024 5531
rect 2982 5469 2996 5489
rect 3016 5469 3024 5489
rect 2982 5431 3024 5469
rect 3098 5489 3140 5531
rect 3098 5469 3106 5489
rect 3126 5469 3140 5489
rect 3098 5431 3140 5469
rect 3190 5489 3234 5531
rect 3190 5469 3202 5489
rect 3222 5469 3234 5489
rect 3190 5431 3234 5469
rect 3306 5489 3348 5531
rect 3306 5469 3314 5489
rect 3334 5469 3348 5489
rect 3306 5431 3348 5469
rect 3398 5489 3442 5531
rect 3398 5469 3410 5489
rect 3430 5469 3442 5489
rect 3398 5431 3442 5469
rect 3519 5489 3561 5531
rect 3519 5469 3527 5489
rect 3547 5469 3561 5489
rect 3519 5431 3561 5469
rect 3611 5489 3655 5531
rect 6334 5594 6378 5636
rect 6428 5656 6470 5694
rect 6428 5636 6442 5656
rect 6462 5636 6470 5656
rect 6428 5594 6470 5636
rect 6547 5656 6591 5694
rect 6547 5636 6559 5656
rect 6579 5636 6591 5656
rect 6547 5594 6591 5636
rect 6641 5656 6683 5694
rect 6641 5636 6655 5656
rect 6675 5636 6683 5656
rect 6641 5594 6683 5636
rect 6755 5656 6799 5694
rect 6755 5636 6767 5656
rect 6787 5636 6799 5656
rect 6755 5594 6799 5636
rect 6849 5656 6891 5694
rect 6849 5636 6863 5656
rect 6883 5636 6891 5656
rect 6849 5594 6891 5636
rect 6965 5656 7007 5694
rect 6965 5636 6973 5656
rect 6993 5636 7007 5656
rect 6965 5594 7007 5636
rect 7057 5663 7102 5694
rect 13858 5784 13870 5804
rect 13890 5784 13902 5804
rect 13858 5777 13902 5784
rect 7057 5656 7101 5663
rect 7057 5636 7069 5656
rect 7089 5636 7101 5656
rect 13857 5746 13902 5777
rect 13952 5804 13994 5846
rect 13952 5784 13966 5804
rect 13986 5784 13994 5804
rect 13952 5746 13994 5784
rect 14068 5804 14110 5846
rect 14068 5784 14076 5804
rect 14096 5784 14110 5804
rect 14068 5746 14110 5784
rect 14160 5804 14204 5846
rect 14160 5784 14172 5804
rect 14192 5784 14204 5804
rect 14160 5746 14204 5784
rect 14276 5804 14318 5846
rect 14276 5784 14284 5804
rect 14304 5784 14318 5804
rect 14276 5746 14318 5784
rect 14368 5804 14412 5846
rect 14368 5784 14380 5804
rect 14400 5784 14412 5804
rect 14368 5746 14412 5784
rect 14489 5804 14531 5846
rect 14489 5784 14497 5804
rect 14517 5784 14531 5804
rect 14489 5746 14531 5784
rect 14581 5804 14625 5846
rect 15427 5843 15471 5885
rect 15521 5905 15563 5943
rect 15521 5885 15535 5905
rect 15555 5885 15563 5905
rect 15521 5843 15563 5885
rect 15640 5905 15684 5943
rect 15640 5885 15652 5905
rect 15672 5885 15684 5905
rect 15640 5843 15684 5885
rect 15734 5905 15776 5943
rect 15734 5885 15748 5905
rect 15768 5885 15776 5905
rect 15734 5843 15776 5885
rect 15848 5905 15892 5943
rect 15848 5885 15860 5905
rect 15880 5885 15892 5905
rect 15848 5843 15892 5885
rect 15942 5905 15984 5943
rect 15942 5885 15956 5905
rect 15976 5885 15984 5905
rect 15942 5843 15984 5885
rect 16058 5905 16100 5943
rect 16058 5885 16066 5905
rect 16086 5885 16100 5905
rect 16058 5843 16100 5885
rect 16150 5912 16195 5943
rect 16150 5905 16194 5912
rect 16150 5885 16162 5905
rect 16182 5885 16194 5905
rect 16150 5843 16194 5885
rect 18914 5845 18958 5887
rect 14581 5784 14593 5804
rect 14613 5784 14625 5804
rect 14581 5746 14625 5784
rect 18914 5825 18926 5845
rect 18946 5825 18958 5845
rect 18914 5818 18958 5825
rect 18913 5787 18958 5818
rect 19008 5845 19050 5887
rect 19008 5825 19022 5845
rect 19042 5825 19050 5845
rect 19008 5787 19050 5825
rect 19124 5845 19166 5887
rect 19124 5825 19132 5845
rect 19152 5825 19166 5845
rect 19124 5787 19166 5825
rect 19216 5845 19260 5887
rect 19216 5825 19228 5845
rect 19248 5825 19260 5845
rect 19216 5787 19260 5825
rect 19332 5845 19374 5887
rect 19332 5825 19340 5845
rect 19360 5825 19374 5845
rect 19332 5787 19374 5825
rect 19424 5845 19468 5887
rect 19424 5825 19436 5845
rect 19456 5825 19468 5845
rect 19424 5787 19468 5825
rect 19545 5845 19587 5887
rect 19545 5825 19553 5845
rect 19573 5825 19587 5845
rect 19545 5787 19587 5825
rect 19637 5845 19681 5887
rect 19637 5825 19649 5845
rect 19669 5825 19681 5845
rect 19637 5787 19681 5825
rect 7057 5594 7101 5636
rect 3611 5469 3623 5489
rect 3643 5469 3655 5489
rect 3611 5431 3655 5469
rect 7944 5530 7988 5572
rect 7944 5510 7956 5530
rect 7976 5510 7988 5530
rect 7944 5503 7988 5510
rect 7943 5472 7988 5503
rect 8038 5530 8080 5572
rect 8038 5510 8052 5530
rect 8072 5510 8080 5530
rect 8038 5472 8080 5510
rect 8154 5530 8196 5572
rect 8154 5510 8162 5530
rect 8182 5510 8196 5530
rect 8154 5472 8196 5510
rect 8246 5530 8290 5572
rect 8246 5510 8258 5530
rect 8278 5510 8290 5530
rect 8246 5472 8290 5510
rect 8362 5530 8404 5572
rect 8362 5510 8370 5530
rect 8390 5510 8404 5530
rect 8362 5472 8404 5510
rect 8454 5530 8498 5572
rect 8454 5510 8466 5530
rect 8486 5510 8498 5530
rect 8454 5472 8498 5510
rect 8575 5530 8617 5572
rect 8575 5510 8583 5530
rect 8603 5510 8617 5530
rect 8575 5472 8617 5510
rect 8667 5530 8711 5572
rect 11309 5620 11353 5658
rect 11309 5600 11321 5620
rect 11341 5600 11353 5620
rect 8667 5510 8679 5530
rect 8699 5510 8711 5530
rect 8667 5472 8711 5510
rect 11309 5558 11353 5600
rect 11403 5620 11445 5658
rect 11403 5600 11417 5620
rect 11437 5600 11445 5620
rect 11403 5558 11445 5600
rect 11522 5620 11566 5658
rect 11522 5600 11534 5620
rect 11554 5600 11566 5620
rect 11522 5558 11566 5600
rect 11616 5620 11658 5658
rect 11616 5600 11630 5620
rect 11650 5600 11658 5620
rect 11616 5558 11658 5600
rect 11730 5620 11774 5658
rect 11730 5600 11742 5620
rect 11762 5600 11774 5620
rect 11730 5558 11774 5600
rect 11824 5620 11866 5658
rect 11824 5600 11838 5620
rect 11858 5600 11866 5620
rect 11824 5558 11866 5600
rect 11940 5620 11982 5658
rect 11940 5600 11948 5620
rect 11968 5600 11982 5620
rect 11940 5558 11982 5600
rect 12032 5627 12077 5658
rect 12032 5620 12076 5627
rect 12032 5600 12044 5620
rect 12064 5600 12076 5620
rect 12032 5558 12076 5600
rect 16365 5661 16409 5699
rect 16365 5641 16377 5661
rect 16397 5641 16409 5661
rect 12919 5494 12963 5536
rect 339 5305 383 5343
rect 339 5285 351 5305
rect 371 5285 383 5305
rect 339 5243 383 5285
rect 433 5305 475 5343
rect 433 5285 447 5305
rect 467 5285 475 5305
rect 433 5243 475 5285
rect 552 5305 596 5343
rect 552 5285 564 5305
rect 584 5285 596 5305
rect 552 5243 596 5285
rect 646 5305 688 5343
rect 646 5285 660 5305
rect 680 5285 688 5305
rect 646 5243 688 5285
rect 760 5305 804 5343
rect 760 5285 772 5305
rect 792 5285 804 5305
rect 760 5243 804 5285
rect 854 5305 896 5343
rect 854 5285 868 5305
rect 888 5285 896 5305
rect 854 5243 896 5285
rect 970 5305 1012 5343
rect 970 5285 978 5305
rect 998 5285 1012 5305
rect 970 5243 1012 5285
rect 1062 5312 1107 5343
rect 1062 5305 1106 5312
rect 1062 5285 1074 5305
rect 1094 5285 1106 5305
rect 5395 5346 5439 5384
rect 5395 5326 5407 5346
rect 5427 5326 5439 5346
rect 1062 5243 1106 5285
rect 3826 5245 3870 5287
rect 3826 5225 3838 5245
rect 3858 5225 3870 5245
rect 3826 5218 3870 5225
rect 3825 5187 3870 5218
rect 3920 5245 3962 5287
rect 3920 5225 3934 5245
rect 3954 5225 3962 5245
rect 3920 5187 3962 5225
rect 4036 5245 4078 5287
rect 4036 5225 4044 5245
rect 4064 5225 4078 5245
rect 4036 5187 4078 5225
rect 4128 5245 4172 5287
rect 4128 5225 4140 5245
rect 4160 5225 4172 5245
rect 4128 5187 4172 5225
rect 4244 5245 4286 5287
rect 4244 5225 4252 5245
rect 4272 5225 4286 5245
rect 4244 5187 4286 5225
rect 4336 5245 4380 5287
rect 4336 5225 4348 5245
rect 4368 5225 4380 5245
rect 4336 5187 4380 5225
rect 4457 5245 4499 5287
rect 4457 5225 4465 5245
rect 4485 5225 4499 5245
rect 4457 5187 4499 5225
rect 4549 5245 4593 5287
rect 5395 5284 5439 5326
rect 5489 5346 5531 5384
rect 5489 5326 5503 5346
rect 5523 5326 5531 5346
rect 5489 5284 5531 5326
rect 5608 5346 5652 5384
rect 5608 5326 5620 5346
rect 5640 5326 5652 5346
rect 5608 5284 5652 5326
rect 5702 5346 5744 5384
rect 5702 5326 5716 5346
rect 5736 5326 5744 5346
rect 5702 5284 5744 5326
rect 5816 5346 5860 5384
rect 5816 5326 5828 5346
rect 5848 5326 5860 5346
rect 5816 5284 5860 5326
rect 5910 5346 5952 5384
rect 5910 5326 5924 5346
rect 5944 5326 5952 5346
rect 5910 5284 5952 5326
rect 6026 5346 6068 5384
rect 6026 5326 6034 5346
rect 6054 5326 6068 5346
rect 6026 5284 6068 5326
rect 6118 5353 6163 5384
rect 12919 5474 12931 5494
rect 12951 5474 12963 5494
rect 12919 5467 12963 5474
rect 6118 5346 6162 5353
rect 6118 5326 6130 5346
rect 6150 5326 6162 5346
rect 12918 5436 12963 5467
rect 13013 5494 13055 5536
rect 13013 5474 13027 5494
rect 13047 5474 13055 5494
rect 13013 5436 13055 5474
rect 13129 5494 13171 5536
rect 13129 5474 13137 5494
rect 13157 5474 13171 5494
rect 13129 5436 13171 5474
rect 13221 5494 13265 5536
rect 13221 5474 13233 5494
rect 13253 5474 13265 5494
rect 13221 5436 13265 5474
rect 13337 5494 13379 5536
rect 13337 5474 13345 5494
rect 13365 5474 13379 5494
rect 13337 5436 13379 5474
rect 13429 5494 13473 5536
rect 13429 5474 13441 5494
rect 13461 5474 13473 5494
rect 13429 5436 13473 5474
rect 13550 5494 13592 5536
rect 13550 5474 13558 5494
rect 13578 5474 13592 5494
rect 13550 5436 13592 5474
rect 13642 5494 13686 5536
rect 16365 5599 16409 5641
rect 16459 5661 16501 5699
rect 16459 5641 16473 5661
rect 16493 5641 16501 5661
rect 16459 5599 16501 5641
rect 16578 5661 16622 5699
rect 16578 5641 16590 5661
rect 16610 5641 16622 5661
rect 16578 5599 16622 5641
rect 16672 5661 16714 5699
rect 16672 5641 16686 5661
rect 16706 5641 16714 5661
rect 16672 5599 16714 5641
rect 16786 5661 16830 5699
rect 16786 5641 16798 5661
rect 16818 5641 16830 5661
rect 16786 5599 16830 5641
rect 16880 5661 16922 5699
rect 16880 5641 16894 5661
rect 16914 5641 16922 5661
rect 16880 5599 16922 5641
rect 16996 5661 17038 5699
rect 16996 5641 17004 5661
rect 17024 5641 17038 5661
rect 16996 5599 17038 5641
rect 17088 5668 17133 5699
rect 17088 5661 17132 5668
rect 17088 5641 17100 5661
rect 17120 5641 17132 5661
rect 17088 5599 17132 5641
rect 13642 5474 13654 5494
rect 13674 5474 13686 5494
rect 13642 5436 13686 5474
rect 17975 5535 18019 5577
rect 17975 5515 17987 5535
rect 18007 5515 18019 5535
rect 17975 5508 18019 5515
rect 17974 5477 18019 5508
rect 18069 5535 18111 5577
rect 18069 5515 18083 5535
rect 18103 5515 18111 5535
rect 18069 5477 18111 5515
rect 18185 5535 18227 5577
rect 18185 5515 18193 5535
rect 18213 5515 18227 5535
rect 18185 5477 18227 5515
rect 18277 5535 18321 5577
rect 18277 5515 18289 5535
rect 18309 5515 18321 5535
rect 18277 5477 18321 5515
rect 18393 5535 18435 5577
rect 18393 5515 18401 5535
rect 18421 5515 18435 5535
rect 18393 5477 18435 5515
rect 18485 5535 18529 5577
rect 18485 5515 18497 5535
rect 18517 5515 18529 5535
rect 18485 5477 18529 5515
rect 18606 5535 18648 5577
rect 18606 5515 18614 5535
rect 18634 5515 18648 5535
rect 18606 5477 18648 5515
rect 18698 5535 18742 5577
rect 18698 5515 18710 5535
rect 18730 5515 18742 5535
rect 18698 5477 18742 5515
rect 6118 5284 6162 5326
rect 8882 5286 8926 5328
rect 4549 5225 4561 5245
rect 4581 5225 4593 5245
rect 4549 5187 4593 5225
rect 8882 5266 8894 5286
rect 8914 5266 8926 5286
rect 8882 5259 8926 5266
rect 8881 5228 8926 5259
rect 8976 5286 9018 5328
rect 8976 5266 8990 5286
rect 9010 5266 9018 5286
rect 8976 5228 9018 5266
rect 9092 5286 9134 5328
rect 9092 5266 9100 5286
rect 9120 5266 9134 5286
rect 9092 5228 9134 5266
rect 9184 5286 9228 5328
rect 9184 5266 9196 5286
rect 9216 5266 9228 5286
rect 9184 5228 9228 5266
rect 9300 5286 9342 5328
rect 9300 5266 9308 5286
rect 9328 5266 9342 5286
rect 9300 5228 9342 5266
rect 9392 5286 9436 5328
rect 9392 5266 9404 5286
rect 9424 5266 9436 5286
rect 9392 5228 9436 5266
rect 9513 5286 9555 5328
rect 9513 5266 9521 5286
rect 9541 5266 9555 5286
rect 9513 5228 9555 5266
rect 9605 5286 9649 5328
rect 9605 5266 9617 5286
rect 9637 5266 9649 5286
rect 10370 5310 10414 5348
rect 10370 5290 10382 5310
rect 10402 5290 10414 5310
rect 9605 5228 9649 5266
rect 10370 5248 10414 5290
rect 10464 5310 10506 5348
rect 10464 5290 10478 5310
rect 10498 5290 10506 5310
rect 10464 5248 10506 5290
rect 10583 5310 10627 5348
rect 10583 5290 10595 5310
rect 10615 5290 10627 5310
rect 10583 5248 10627 5290
rect 10677 5310 10719 5348
rect 10677 5290 10691 5310
rect 10711 5290 10719 5310
rect 10677 5248 10719 5290
rect 10791 5310 10835 5348
rect 10791 5290 10803 5310
rect 10823 5290 10835 5310
rect 10791 5248 10835 5290
rect 10885 5310 10927 5348
rect 10885 5290 10899 5310
rect 10919 5290 10927 5310
rect 10885 5248 10927 5290
rect 11001 5310 11043 5348
rect 11001 5290 11009 5310
rect 11029 5290 11043 5310
rect 11001 5248 11043 5290
rect 11093 5317 11138 5348
rect 11093 5310 11137 5317
rect 11093 5290 11105 5310
rect 11125 5290 11137 5310
rect 15426 5351 15470 5389
rect 15426 5331 15438 5351
rect 15458 5331 15470 5351
rect 11093 5248 11137 5290
rect 13857 5250 13901 5292
rect 1387 5042 1431 5080
rect 1387 5022 1399 5042
rect 1419 5022 1431 5042
rect 1387 4980 1431 5022
rect 1481 5042 1523 5080
rect 1481 5022 1495 5042
rect 1515 5022 1523 5042
rect 1481 4980 1523 5022
rect 1600 5042 1644 5080
rect 1600 5022 1612 5042
rect 1632 5022 1644 5042
rect 1600 4980 1644 5022
rect 1694 5042 1736 5080
rect 1694 5022 1708 5042
rect 1728 5022 1736 5042
rect 1694 4980 1736 5022
rect 1808 5042 1852 5080
rect 1808 5022 1820 5042
rect 1840 5022 1852 5042
rect 1808 4980 1852 5022
rect 1902 5042 1944 5080
rect 1902 5022 1916 5042
rect 1936 5022 1944 5042
rect 1902 4980 1944 5022
rect 2018 5042 2060 5080
rect 2018 5022 2026 5042
rect 2046 5022 2060 5042
rect 2018 4980 2060 5022
rect 2110 5049 2155 5080
rect 2110 5042 2154 5049
rect 2110 5022 2122 5042
rect 2142 5022 2154 5042
rect 2110 4980 2154 5022
rect 6443 5083 6487 5121
rect 6443 5063 6455 5083
rect 6475 5063 6487 5083
rect 6443 5021 6487 5063
rect 6537 5083 6579 5121
rect 6537 5063 6551 5083
rect 6571 5063 6579 5083
rect 6537 5021 6579 5063
rect 6656 5083 6700 5121
rect 6656 5063 6668 5083
rect 6688 5063 6700 5083
rect 6656 5021 6700 5063
rect 6750 5083 6792 5121
rect 6750 5063 6764 5083
rect 6784 5063 6792 5083
rect 6750 5021 6792 5063
rect 6864 5083 6908 5121
rect 6864 5063 6876 5083
rect 6896 5063 6908 5083
rect 6864 5021 6908 5063
rect 6958 5083 7000 5121
rect 6958 5063 6972 5083
rect 6992 5063 7000 5083
rect 6958 5021 7000 5063
rect 7074 5083 7116 5121
rect 7074 5063 7082 5083
rect 7102 5063 7116 5083
rect 7074 5021 7116 5063
rect 7166 5090 7211 5121
rect 13857 5230 13869 5250
rect 13889 5230 13901 5250
rect 13857 5223 13901 5230
rect 13856 5192 13901 5223
rect 13951 5250 13993 5292
rect 13951 5230 13965 5250
rect 13985 5230 13993 5250
rect 13951 5192 13993 5230
rect 14067 5250 14109 5292
rect 14067 5230 14075 5250
rect 14095 5230 14109 5250
rect 14067 5192 14109 5230
rect 14159 5250 14203 5292
rect 14159 5230 14171 5250
rect 14191 5230 14203 5250
rect 14159 5192 14203 5230
rect 14275 5250 14317 5292
rect 14275 5230 14283 5250
rect 14303 5230 14317 5250
rect 14275 5192 14317 5230
rect 14367 5250 14411 5292
rect 14367 5230 14379 5250
rect 14399 5230 14411 5250
rect 14367 5192 14411 5230
rect 14488 5250 14530 5292
rect 14488 5230 14496 5250
rect 14516 5230 14530 5250
rect 14488 5192 14530 5230
rect 14580 5250 14624 5292
rect 15426 5289 15470 5331
rect 15520 5351 15562 5389
rect 15520 5331 15534 5351
rect 15554 5331 15562 5351
rect 15520 5289 15562 5331
rect 15639 5351 15683 5389
rect 15639 5331 15651 5351
rect 15671 5331 15683 5351
rect 15639 5289 15683 5331
rect 15733 5351 15775 5389
rect 15733 5331 15747 5351
rect 15767 5331 15775 5351
rect 15733 5289 15775 5331
rect 15847 5351 15891 5389
rect 15847 5331 15859 5351
rect 15879 5331 15891 5351
rect 15847 5289 15891 5331
rect 15941 5351 15983 5389
rect 15941 5331 15955 5351
rect 15975 5331 15983 5351
rect 15941 5289 15983 5331
rect 16057 5351 16099 5389
rect 16057 5331 16065 5351
rect 16085 5331 16099 5351
rect 16057 5289 16099 5331
rect 16149 5358 16194 5389
rect 16149 5351 16193 5358
rect 16149 5331 16161 5351
rect 16181 5331 16193 5351
rect 16149 5289 16193 5331
rect 18913 5291 18957 5333
rect 14580 5230 14592 5250
rect 14612 5230 14624 5250
rect 14580 5192 14624 5230
rect 18913 5271 18925 5291
rect 18945 5271 18957 5291
rect 18913 5264 18957 5271
rect 18912 5233 18957 5264
rect 19007 5291 19049 5333
rect 19007 5271 19021 5291
rect 19041 5271 19049 5291
rect 19007 5233 19049 5271
rect 19123 5291 19165 5333
rect 19123 5271 19131 5291
rect 19151 5271 19165 5291
rect 19123 5233 19165 5271
rect 19215 5291 19259 5333
rect 19215 5271 19227 5291
rect 19247 5271 19259 5291
rect 19215 5233 19259 5271
rect 19331 5291 19373 5333
rect 19331 5271 19339 5291
rect 19359 5271 19373 5291
rect 19331 5233 19373 5271
rect 19423 5291 19467 5333
rect 19423 5271 19435 5291
rect 19455 5271 19467 5291
rect 19423 5233 19467 5271
rect 19544 5291 19586 5333
rect 19544 5271 19552 5291
rect 19572 5271 19586 5291
rect 19544 5233 19586 5271
rect 19636 5291 19680 5333
rect 19636 5271 19648 5291
rect 19668 5271 19680 5291
rect 19636 5233 19680 5271
rect 7166 5083 7210 5090
rect 7166 5063 7178 5083
rect 7198 5063 7210 5083
rect 7166 5021 7210 5063
rect 2779 4959 2823 5001
rect 2779 4939 2791 4959
rect 2811 4939 2823 4959
rect 2779 4932 2823 4939
rect 2778 4901 2823 4932
rect 2873 4959 2915 5001
rect 2873 4939 2887 4959
rect 2907 4939 2915 4959
rect 2873 4901 2915 4939
rect 2989 4959 3031 5001
rect 2989 4939 2997 4959
rect 3017 4939 3031 4959
rect 2989 4901 3031 4939
rect 3081 4959 3125 5001
rect 3081 4939 3093 4959
rect 3113 4939 3125 4959
rect 3081 4901 3125 4939
rect 3197 4959 3239 5001
rect 3197 4939 3205 4959
rect 3225 4939 3239 4959
rect 3197 4901 3239 4939
rect 3289 4959 3333 5001
rect 3289 4939 3301 4959
rect 3321 4939 3333 4959
rect 3289 4901 3333 4939
rect 3410 4959 3452 5001
rect 3410 4939 3418 4959
rect 3438 4939 3452 4959
rect 3410 4901 3452 4939
rect 3502 4959 3546 5001
rect 3502 4939 3514 4959
rect 3534 4939 3546 4959
rect 3502 4901 3546 4939
rect 7835 5000 7879 5042
rect 7835 4980 7847 5000
rect 7867 4980 7879 5000
rect 7835 4973 7879 4980
rect 7834 4942 7879 4973
rect 7929 5000 7971 5042
rect 7929 4980 7943 5000
rect 7963 4980 7971 5000
rect 7929 4942 7971 4980
rect 8045 5000 8087 5042
rect 8045 4980 8053 5000
rect 8073 4980 8087 5000
rect 8045 4942 8087 4980
rect 8137 5000 8181 5042
rect 8137 4980 8149 5000
rect 8169 4980 8181 5000
rect 8137 4942 8181 4980
rect 8253 5000 8295 5042
rect 8253 4980 8261 5000
rect 8281 4980 8295 5000
rect 8253 4942 8295 4980
rect 8345 5000 8389 5042
rect 8345 4980 8357 5000
rect 8377 4980 8389 5000
rect 8345 4942 8389 4980
rect 8466 5000 8508 5042
rect 8466 4980 8474 5000
rect 8494 4980 8508 5000
rect 8466 4942 8508 4980
rect 8558 5000 8602 5042
rect 11418 5047 11462 5085
rect 8558 4980 8570 5000
rect 8590 4980 8602 5000
rect 11418 5027 11430 5047
rect 11450 5027 11462 5047
rect 8558 4942 8602 4980
rect 11418 4985 11462 5027
rect 11512 5047 11554 5085
rect 11512 5027 11526 5047
rect 11546 5027 11554 5047
rect 11512 4985 11554 5027
rect 11631 5047 11675 5085
rect 11631 5027 11643 5047
rect 11663 5027 11675 5047
rect 11631 4985 11675 5027
rect 11725 5047 11767 5085
rect 11725 5027 11739 5047
rect 11759 5027 11767 5047
rect 11725 4985 11767 5027
rect 11839 5047 11883 5085
rect 11839 5027 11851 5047
rect 11871 5027 11883 5047
rect 11839 4985 11883 5027
rect 11933 5047 11975 5085
rect 11933 5027 11947 5047
rect 11967 5027 11975 5047
rect 11933 4985 11975 5027
rect 12049 5047 12091 5085
rect 12049 5027 12057 5047
rect 12077 5027 12091 5047
rect 12049 4985 12091 5027
rect 12141 5054 12186 5085
rect 12141 5047 12185 5054
rect 12141 5027 12153 5047
rect 12173 5027 12185 5047
rect 12141 4985 12185 5027
rect 16474 5088 16518 5126
rect 16474 5068 16486 5088
rect 16506 5068 16518 5088
rect 16474 5026 16518 5068
rect 16568 5088 16610 5126
rect 16568 5068 16582 5088
rect 16602 5068 16610 5088
rect 16568 5026 16610 5068
rect 16687 5088 16731 5126
rect 16687 5068 16699 5088
rect 16719 5068 16731 5088
rect 16687 5026 16731 5068
rect 16781 5088 16823 5126
rect 16781 5068 16795 5088
rect 16815 5068 16823 5088
rect 16781 5026 16823 5068
rect 16895 5088 16939 5126
rect 16895 5068 16907 5088
rect 16927 5068 16939 5088
rect 16895 5026 16939 5068
rect 16989 5088 17031 5126
rect 16989 5068 17003 5088
rect 17023 5068 17031 5088
rect 16989 5026 17031 5068
rect 17105 5088 17147 5126
rect 17105 5068 17113 5088
rect 17133 5068 17147 5088
rect 17105 5026 17147 5068
rect 17197 5095 17242 5126
rect 17197 5088 17241 5095
rect 17197 5068 17209 5088
rect 17229 5068 17241 5088
rect 17197 5026 17241 5068
rect 12810 4964 12854 5006
rect 12810 4944 12822 4964
rect 12842 4944 12854 4964
rect 12810 4937 12854 4944
rect 340 4756 384 4794
rect 340 4736 352 4756
rect 372 4736 384 4756
rect 340 4694 384 4736
rect 434 4756 476 4794
rect 434 4736 448 4756
rect 468 4736 476 4756
rect 434 4694 476 4736
rect 553 4756 597 4794
rect 553 4736 565 4756
rect 585 4736 597 4756
rect 553 4694 597 4736
rect 647 4756 689 4794
rect 647 4736 661 4756
rect 681 4736 689 4756
rect 647 4694 689 4736
rect 761 4756 805 4794
rect 761 4736 773 4756
rect 793 4736 805 4756
rect 761 4694 805 4736
rect 855 4756 897 4794
rect 855 4736 869 4756
rect 889 4736 897 4756
rect 855 4694 897 4736
rect 971 4756 1013 4794
rect 971 4736 979 4756
rect 999 4736 1013 4756
rect 971 4694 1013 4736
rect 1063 4763 1108 4794
rect 1063 4756 1107 4763
rect 1063 4736 1075 4756
rect 1095 4736 1107 4756
rect 5396 4797 5440 4835
rect 5396 4777 5408 4797
rect 5428 4777 5440 4797
rect 1063 4694 1107 4736
rect 3827 4696 3871 4738
rect 3827 4676 3839 4696
rect 3859 4676 3871 4696
rect 3827 4669 3871 4676
rect 3826 4638 3871 4669
rect 3921 4696 3963 4738
rect 3921 4676 3935 4696
rect 3955 4676 3963 4696
rect 3921 4638 3963 4676
rect 4037 4696 4079 4738
rect 4037 4676 4045 4696
rect 4065 4676 4079 4696
rect 4037 4638 4079 4676
rect 4129 4696 4173 4738
rect 4129 4676 4141 4696
rect 4161 4676 4173 4696
rect 4129 4638 4173 4676
rect 4245 4696 4287 4738
rect 4245 4676 4253 4696
rect 4273 4676 4287 4696
rect 4245 4638 4287 4676
rect 4337 4696 4381 4738
rect 4337 4676 4349 4696
rect 4369 4676 4381 4696
rect 4337 4638 4381 4676
rect 4458 4696 4500 4738
rect 4458 4676 4466 4696
rect 4486 4676 4500 4696
rect 4458 4638 4500 4676
rect 4550 4696 4594 4738
rect 5396 4735 5440 4777
rect 5490 4797 5532 4835
rect 5490 4777 5504 4797
rect 5524 4777 5532 4797
rect 5490 4735 5532 4777
rect 5609 4797 5653 4835
rect 5609 4777 5621 4797
rect 5641 4777 5653 4797
rect 5609 4735 5653 4777
rect 5703 4797 5745 4835
rect 5703 4777 5717 4797
rect 5737 4777 5745 4797
rect 5703 4735 5745 4777
rect 5817 4797 5861 4835
rect 5817 4777 5829 4797
rect 5849 4777 5861 4797
rect 5817 4735 5861 4777
rect 5911 4797 5953 4835
rect 5911 4777 5925 4797
rect 5945 4777 5953 4797
rect 5911 4735 5953 4777
rect 6027 4797 6069 4835
rect 6027 4777 6035 4797
rect 6055 4777 6069 4797
rect 6027 4735 6069 4777
rect 6119 4804 6164 4835
rect 6119 4797 6163 4804
rect 6119 4777 6131 4797
rect 6151 4777 6163 4797
rect 12809 4906 12854 4937
rect 12904 4964 12946 5006
rect 12904 4944 12918 4964
rect 12938 4944 12946 4964
rect 12904 4906 12946 4944
rect 13020 4964 13062 5006
rect 13020 4944 13028 4964
rect 13048 4944 13062 4964
rect 13020 4906 13062 4944
rect 13112 4964 13156 5006
rect 13112 4944 13124 4964
rect 13144 4944 13156 4964
rect 13112 4906 13156 4944
rect 13228 4964 13270 5006
rect 13228 4944 13236 4964
rect 13256 4944 13270 4964
rect 13228 4906 13270 4944
rect 13320 4964 13364 5006
rect 13320 4944 13332 4964
rect 13352 4944 13364 4964
rect 13320 4906 13364 4944
rect 13441 4964 13483 5006
rect 13441 4944 13449 4964
rect 13469 4944 13483 4964
rect 13441 4906 13483 4944
rect 13533 4964 13577 5006
rect 13533 4944 13545 4964
rect 13565 4944 13577 4964
rect 13533 4906 13577 4944
rect 17866 5005 17910 5047
rect 17866 4985 17878 5005
rect 17898 4985 17910 5005
rect 17866 4978 17910 4985
rect 17865 4947 17910 4978
rect 17960 5005 18002 5047
rect 17960 4985 17974 5005
rect 17994 4985 18002 5005
rect 17960 4947 18002 4985
rect 18076 5005 18118 5047
rect 18076 4985 18084 5005
rect 18104 4985 18118 5005
rect 18076 4947 18118 4985
rect 18168 5005 18212 5047
rect 18168 4985 18180 5005
rect 18200 4985 18212 5005
rect 18168 4947 18212 4985
rect 18284 5005 18326 5047
rect 18284 4985 18292 5005
rect 18312 4985 18326 5005
rect 18284 4947 18326 4985
rect 18376 5005 18420 5047
rect 18376 4985 18388 5005
rect 18408 4985 18420 5005
rect 18376 4947 18420 4985
rect 18497 5005 18539 5047
rect 18497 4985 18505 5005
rect 18525 4985 18539 5005
rect 18497 4947 18539 4985
rect 18589 5005 18633 5047
rect 18589 4985 18601 5005
rect 18621 4985 18633 5005
rect 18589 4947 18633 4985
rect 6119 4735 6163 4777
rect 8883 4737 8927 4779
rect 4550 4676 4562 4696
rect 4582 4676 4594 4696
rect 4550 4638 4594 4676
rect 8883 4717 8895 4737
rect 8915 4717 8927 4737
rect 8883 4710 8927 4717
rect 8882 4679 8927 4710
rect 8977 4737 9019 4779
rect 8977 4717 8991 4737
rect 9011 4717 9019 4737
rect 8977 4679 9019 4717
rect 9093 4737 9135 4779
rect 9093 4717 9101 4737
rect 9121 4717 9135 4737
rect 9093 4679 9135 4717
rect 9185 4737 9229 4779
rect 9185 4717 9197 4737
rect 9217 4717 9229 4737
rect 9185 4679 9229 4717
rect 9301 4737 9343 4779
rect 9301 4717 9309 4737
rect 9329 4717 9343 4737
rect 9301 4679 9343 4717
rect 9393 4737 9437 4779
rect 9393 4717 9405 4737
rect 9425 4717 9437 4737
rect 9393 4679 9437 4717
rect 9514 4737 9556 4779
rect 9514 4717 9522 4737
rect 9542 4717 9556 4737
rect 9514 4679 9556 4717
rect 9606 4737 9650 4779
rect 10371 4761 10415 4799
rect 9606 4717 9618 4737
rect 9638 4717 9650 4737
rect 9606 4679 9650 4717
rect 10371 4741 10383 4761
rect 10403 4741 10415 4761
rect 10371 4699 10415 4741
rect 10465 4761 10507 4799
rect 10465 4741 10479 4761
rect 10499 4741 10507 4761
rect 10465 4699 10507 4741
rect 10584 4761 10628 4799
rect 10584 4741 10596 4761
rect 10616 4741 10628 4761
rect 10584 4699 10628 4741
rect 10678 4761 10720 4799
rect 10678 4741 10692 4761
rect 10712 4741 10720 4761
rect 10678 4699 10720 4741
rect 10792 4761 10836 4799
rect 10792 4741 10804 4761
rect 10824 4741 10836 4761
rect 10792 4699 10836 4741
rect 10886 4761 10928 4799
rect 10886 4741 10900 4761
rect 10920 4741 10928 4761
rect 10886 4699 10928 4741
rect 11002 4761 11044 4799
rect 11002 4741 11010 4761
rect 11030 4741 11044 4761
rect 11002 4699 11044 4741
rect 11094 4768 11139 4799
rect 11094 4761 11138 4768
rect 11094 4741 11106 4761
rect 11126 4741 11138 4761
rect 15427 4802 15471 4840
rect 15427 4782 15439 4802
rect 15459 4782 15471 4802
rect 11094 4699 11138 4741
rect 13858 4701 13902 4743
rect 1278 4512 1322 4550
rect 1278 4492 1290 4512
rect 1310 4492 1322 4512
rect 1278 4450 1322 4492
rect 1372 4512 1414 4550
rect 1372 4492 1386 4512
rect 1406 4492 1414 4512
rect 1372 4450 1414 4492
rect 1491 4512 1535 4550
rect 1491 4492 1503 4512
rect 1523 4492 1535 4512
rect 1491 4450 1535 4492
rect 1585 4512 1627 4550
rect 1585 4492 1599 4512
rect 1619 4492 1627 4512
rect 1585 4450 1627 4492
rect 1699 4512 1743 4550
rect 1699 4492 1711 4512
rect 1731 4492 1743 4512
rect 1699 4450 1743 4492
rect 1793 4512 1835 4550
rect 1793 4492 1807 4512
rect 1827 4492 1835 4512
rect 1793 4450 1835 4492
rect 1909 4512 1951 4550
rect 1909 4492 1917 4512
rect 1937 4492 1951 4512
rect 1909 4450 1951 4492
rect 2001 4519 2046 4550
rect 2001 4512 2045 4519
rect 2001 4492 2013 4512
rect 2033 4492 2045 4512
rect 2001 4450 2045 4492
rect 6334 4553 6378 4591
rect 6334 4533 6346 4553
rect 6366 4533 6378 4553
rect 2888 4386 2932 4428
rect 2888 4366 2900 4386
rect 2920 4366 2932 4386
rect 2888 4359 2932 4366
rect 2887 4328 2932 4359
rect 2982 4386 3024 4428
rect 2982 4366 2996 4386
rect 3016 4366 3024 4386
rect 2982 4328 3024 4366
rect 3098 4386 3140 4428
rect 3098 4366 3106 4386
rect 3126 4366 3140 4386
rect 3098 4328 3140 4366
rect 3190 4386 3234 4428
rect 3190 4366 3202 4386
rect 3222 4366 3234 4386
rect 3190 4328 3234 4366
rect 3306 4386 3348 4428
rect 3306 4366 3314 4386
rect 3334 4366 3348 4386
rect 3306 4328 3348 4366
rect 3398 4386 3442 4428
rect 3398 4366 3410 4386
rect 3430 4366 3442 4386
rect 3398 4328 3442 4366
rect 3519 4386 3561 4428
rect 3519 4366 3527 4386
rect 3547 4366 3561 4386
rect 3519 4328 3561 4366
rect 3611 4386 3655 4428
rect 6334 4491 6378 4533
rect 6428 4553 6470 4591
rect 6428 4533 6442 4553
rect 6462 4533 6470 4553
rect 6428 4491 6470 4533
rect 6547 4553 6591 4591
rect 6547 4533 6559 4553
rect 6579 4533 6591 4553
rect 6547 4491 6591 4533
rect 6641 4553 6683 4591
rect 6641 4533 6655 4553
rect 6675 4533 6683 4553
rect 6641 4491 6683 4533
rect 6755 4553 6799 4591
rect 6755 4533 6767 4553
rect 6787 4533 6799 4553
rect 6755 4491 6799 4533
rect 6849 4553 6891 4591
rect 6849 4533 6863 4553
rect 6883 4533 6891 4553
rect 6849 4491 6891 4533
rect 6965 4553 7007 4591
rect 6965 4533 6973 4553
rect 6993 4533 7007 4553
rect 6965 4491 7007 4533
rect 7057 4560 7102 4591
rect 13858 4681 13870 4701
rect 13890 4681 13902 4701
rect 13858 4674 13902 4681
rect 7057 4553 7101 4560
rect 7057 4533 7069 4553
rect 7089 4533 7101 4553
rect 13857 4643 13902 4674
rect 13952 4701 13994 4743
rect 13952 4681 13966 4701
rect 13986 4681 13994 4701
rect 13952 4643 13994 4681
rect 14068 4701 14110 4743
rect 14068 4681 14076 4701
rect 14096 4681 14110 4701
rect 14068 4643 14110 4681
rect 14160 4701 14204 4743
rect 14160 4681 14172 4701
rect 14192 4681 14204 4701
rect 14160 4643 14204 4681
rect 14276 4701 14318 4743
rect 14276 4681 14284 4701
rect 14304 4681 14318 4701
rect 14276 4643 14318 4681
rect 14368 4701 14412 4743
rect 14368 4681 14380 4701
rect 14400 4681 14412 4701
rect 14368 4643 14412 4681
rect 14489 4701 14531 4743
rect 14489 4681 14497 4701
rect 14517 4681 14531 4701
rect 14489 4643 14531 4681
rect 14581 4701 14625 4743
rect 15427 4740 15471 4782
rect 15521 4802 15563 4840
rect 15521 4782 15535 4802
rect 15555 4782 15563 4802
rect 15521 4740 15563 4782
rect 15640 4802 15684 4840
rect 15640 4782 15652 4802
rect 15672 4782 15684 4802
rect 15640 4740 15684 4782
rect 15734 4802 15776 4840
rect 15734 4782 15748 4802
rect 15768 4782 15776 4802
rect 15734 4740 15776 4782
rect 15848 4802 15892 4840
rect 15848 4782 15860 4802
rect 15880 4782 15892 4802
rect 15848 4740 15892 4782
rect 15942 4802 15984 4840
rect 15942 4782 15956 4802
rect 15976 4782 15984 4802
rect 15942 4740 15984 4782
rect 16058 4802 16100 4840
rect 16058 4782 16066 4802
rect 16086 4782 16100 4802
rect 16058 4740 16100 4782
rect 16150 4809 16195 4840
rect 16150 4802 16194 4809
rect 16150 4782 16162 4802
rect 16182 4782 16194 4802
rect 16150 4740 16194 4782
rect 18914 4742 18958 4784
rect 14581 4681 14593 4701
rect 14613 4681 14625 4701
rect 14581 4643 14625 4681
rect 18914 4722 18926 4742
rect 18946 4722 18958 4742
rect 18914 4715 18958 4722
rect 18913 4684 18958 4715
rect 19008 4742 19050 4784
rect 19008 4722 19022 4742
rect 19042 4722 19050 4742
rect 19008 4684 19050 4722
rect 19124 4742 19166 4784
rect 19124 4722 19132 4742
rect 19152 4722 19166 4742
rect 19124 4684 19166 4722
rect 19216 4742 19260 4784
rect 19216 4722 19228 4742
rect 19248 4722 19260 4742
rect 19216 4684 19260 4722
rect 19332 4742 19374 4784
rect 19332 4722 19340 4742
rect 19360 4722 19374 4742
rect 19332 4684 19374 4722
rect 19424 4742 19468 4784
rect 19424 4722 19436 4742
rect 19456 4722 19468 4742
rect 19424 4684 19468 4722
rect 19545 4742 19587 4784
rect 19545 4722 19553 4742
rect 19573 4722 19587 4742
rect 19545 4684 19587 4722
rect 19637 4742 19681 4784
rect 19637 4722 19649 4742
rect 19669 4722 19681 4742
rect 19637 4684 19681 4722
rect 7057 4491 7101 4533
rect 3611 4366 3623 4386
rect 3643 4366 3655 4386
rect 3611 4328 3655 4366
rect 7944 4427 7988 4469
rect 7944 4407 7956 4427
rect 7976 4407 7988 4427
rect 7944 4400 7988 4407
rect 7943 4369 7988 4400
rect 8038 4427 8080 4469
rect 8038 4407 8052 4427
rect 8072 4407 8080 4427
rect 8038 4369 8080 4407
rect 8154 4427 8196 4469
rect 8154 4407 8162 4427
rect 8182 4407 8196 4427
rect 8154 4369 8196 4407
rect 8246 4427 8290 4469
rect 8246 4407 8258 4427
rect 8278 4407 8290 4427
rect 8246 4369 8290 4407
rect 8362 4427 8404 4469
rect 8362 4407 8370 4427
rect 8390 4407 8404 4427
rect 8362 4369 8404 4407
rect 8454 4427 8498 4469
rect 8454 4407 8466 4427
rect 8486 4407 8498 4427
rect 8454 4369 8498 4407
rect 8575 4427 8617 4469
rect 8575 4407 8583 4427
rect 8603 4407 8617 4427
rect 8575 4369 8617 4407
rect 8667 4427 8711 4469
rect 11309 4517 11353 4555
rect 11309 4497 11321 4517
rect 11341 4497 11353 4517
rect 8667 4407 8679 4427
rect 8699 4407 8711 4427
rect 8667 4369 8711 4407
rect 11309 4455 11353 4497
rect 11403 4517 11445 4555
rect 11403 4497 11417 4517
rect 11437 4497 11445 4517
rect 11403 4455 11445 4497
rect 11522 4517 11566 4555
rect 11522 4497 11534 4517
rect 11554 4497 11566 4517
rect 11522 4455 11566 4497
rect 11616 4517 11658 4555
rect 11616 4497 11630 4517
rect 11650 4497 11658 4517
rect 11616 4455 11658 4497
rect 11730 4517 11774 4555
rect 11730 4497 11742 4517
rect 11762 4497 11774 4517
rect 11730 4455 11774 4497
rect 11824 4517 11866 4555
rect 11824 4497 11838 4517
rect 11858 4497 11866 4517
rect 11824 4455 11866 4497
rect 11940 4517 11982 4555
rect 11940 4497 11948 4517
rect 11968 4497 11982 4517
rect 11940 4455 11982 4497
rect 12032 4524 12077 4555
rect 12032 4517 12076 4524
rect 12032 4497 12044 4517
rect 12064 4497 12076 4517
rect 12032 4455 12076 4497
rect 16365 4558 16409 4596
rect 16365 4538 16377 4558
rect 16397 4538 16409 4558
rect 12919 4391 12963 4433
rect 339 4202 383 4240
rect 339 4182 351 4202
rect 371 4182 383 4202
rect 339 4140 383 4182
rect 433 4202 475 4240
rect 433 4182 447 4202
rect 467 4182 475 4202
rect 433 4140 475 4182
rect 552 4202 596 4240
rect 552 4182 564 4202
rect 584 4182 596 4202
rect 552 4140 596 4182
rect 646 4202 688 4240
rect 646 4182 660 4202
rect 680 4182 688 4202
rect 646 4140 688 4182
rect 760 4202 804 4240
rect 760 4182 772 4202
rect 792 4182 804 4202
rect 760 4140 804 4182
rect 854 4202 896 4240
rect 854 4182 868 4202
rect 888 4182 896 4202
rect 854 4140 896 4182
rect 970 4202 1012 4240
rect 970 4182 978 4202
rect 998 4182 1012 4202
rect 970 4140 1012 4182
rect 1062 4209 1107 4240
rect 1062 4202 1106 4209
rect 1062 4182 1074 4202
rect 1094 4182 1106 4202
rect 5395 4243 5439 4281
rect 5395 4223 5407 4243
rect 5427 4223 5439 4243
rect 1062 4140 1106 4182
rect 3826 4142 3870 4184
rect 3826 4122 3838 4142
rect 3858 4122 3870 4142
rect 3826 4115 3870 4122
rect 3825 4084 3870 4115
rect 3920 4142 3962 4184
rect 3920 4122 3934 4142
rect 3954 4122 3962 4142
rect 3920 4084 3962 4122
rect 4036 4142 4078 4184
rect 4036 4122 4044 4142
rect 4064 4122 4078 4142
rect 4036 4084 4078 4122
rect 4128 4142 4172 4184
rect 4128 4122 4140 4142
rect 4160 4122 4172 4142
rect 4128 4084 4172 4122
rect 4244 4142 4286 4184
rect 4244 4122 4252 4142
rect 4272 4122 4286 4142
rect 4244 4084 4286 4122
rect 4336 4142 4380 4184
rect 4336 4122 4348 4142
rect 4368 4122 4380 4142
rect 4336 4084 4380 4122
rect 4457 4142 4499 4184
rect 4457 4122 4465 4142
rect 4485 4122 4499 4142
rect 4457 4084 4499 4122
rect 4549 4142 4593 4184
rect 5395 4181 5439 4223
rect 5489 4243 5531 4281
rect 5489 4223 5503 4243
rect 5523 4223 5531 4243
rect 5489 4181 5531 4223
rect 5608 4243 5652 4281
rect 5608 4223 5620 4243
rect 5640 4223 5652 4243
rect 5608 4181 5652 4223
rect 5702 4243 5744 4281
rect 5702 4223 5716 4243
rect 5736 4223 5744 4243
rect 5702 4181 5744 4223
rect 5816 4243 5860 4281
rect 5816 4223 5828 4243
rect 5848 4223 5860 4243
rect 5816 4181 5860 4223
rect 5910 4243 5952 4281
rect 5910 4223 5924 4243
rect 5944 4223 5952 4243
rect 5910 4181 5952 4223
rect 6026 4243 6068 4281
rect 6026 4223 6034 4243
rect 6054 4223 6068 4243
rect 6026 4181 6068 4223
rect 6118 4250 6163 4281
rect 12919 4371 12931 4391
rect 12951 4371 12963 4391
rect 12919 4364 12963 4371
rect 6118 4243 6162 4250
rect 6118 4223 6130 4243
rect 6150 4223 6162 4243
rect 12918 4333 12963 4364
rect 13013 4391 13055 4433
rect 13013 4371 13027 4391
rect 13047 4371 13055 4391
rect 13013 4333 13055 4371
rect 13129 4391 13171 4433
rect 13129 4371 13137 4391
rect 13157 4371 13171 4391
rect 13129 4333 13171 4371
rect 13221 4391 13265 4433
rect 13221 4371 13233 4391
rect 13253 4371 13265 4391
rect 13221 4333 13265 4371
rect 13337 4391 13379 4433
rect 13337 4371 13345 4391
rect 13365 4371 13379 4391
rect 13337 4333 13379 4371
rect 13429 4391 13473 4433
rect 13429 4371 13441 4391
rect 13461 4371 13473 4391
rect 13429 4333 13473 4371
rect 13550 4391 13592 4433
rect 13550 4371 13558 4391
rect 13578 4371 13592 4391
rect 13550 4333 13592 4371
rect 13642 4391 13686 4433
rect 16365 4496 16409 4538
rect 16459 4558 16501 4596
rect 16459 4538 16473 4558
rect 16493 4538 16501 4558
rect 16459 4496 16501 4538
rect 16578 4558 16622 4596
rect 16578 4538 16590 4558
rect 16610 4538 16622 4558
rect 16578 4496 16622 4538
rect 16672 4558 16714 4596
rect 16672 4538 16686 4558
rect 16706 4538 16714 4558
rect 16672 4496 16714 4538
rect 16786 4558 16830 4596
rect 16786 4538 16798 4558
rect 16818 4538 16830 4558
rect 16786 4496 16830 4538
rect 16880 4558 16922 4596
rect 16880 4538 16894 4558
rect 16914 4538 16922 4558
rect 16880 4496 16922 4538
rect 16996 4558 17038 4596
rect 16996 4538 17004 4558
rect 17024 4538 17038 4558
rect 16996 4496 17038 4538
rect 17088 4565 17133 4596
rect 17088 4558 17132 4565
rect 17088 4538 17100 4558
rect 17120 4538 17132 4558
rect 17088 4496 17132 4538
rect 13642 4371 13654 4391
rect 13674 4371 13686 4391
rect 13642 4333 13686 4371
rect 17975 4432 18019 4474
rect 17975 4412 17987 4432
rect 18007 4412 18019 4432
rect 17975 4405 18019 4412
rect 17974 4374 18019 4405
rect 18069 4432 18111 4474
rect 18069 4412 18083 4432
rect 18103 4412 18111 4432
rect 18069 4374 18111 4412
rect 18185 4432 18227 4474
rect 18185 4412 18193 4432
rect 18213 4412 18227 4432
rect 18185 4374 18227 4412
rect 18277 4432 18321 4474
rect 18277 4412 18289 4432
rect 18309 4412 18321 4432
rect 18277 4374 18321 4412
rect 18393 4432 18435 4474
rect 18393 4412 18401 4432
rect 18421 4412 18435 4432
rect 18393 4374 18435 4412
rect 18485 4432 18529 4474
rect 18485 4412 18497 4432
rect 18517 4412 18529 4432
rect 18485 4374 18529 4412
rect 18606 4432 18648 4474
rect 18606 4412 18614 4432
rect 18634 4412 18648 4432
rect 18606 4374 18648 4412
rect 18698 4432 18742 4474
rect 18698 4412 18710 4432
rect 18730 4412 18742 4432
rect 18698 4374 18742 4412
rect 6118 4181 6162 4223
rect 8882 4183 8926 4225
rect 4549 4122 4561 4142
rect 4581 4122 4593 4142
rect 4549 4084 4593 4122
rect 8882 4163 8894 4183
rect 8914 4163 8926 4183
rect 8882 4156 8926 4163
rect 8881 4125 8926 4156
rect 8976 4183 9018 4225
rect 8976 4163 8990 4183
rect 9010 4163 9018 4183
rect 8976 4125 9018 4163
rect 9092 4183 9134 4225
rect 9092 4163 9100 4183
rect 9120 4163 9134 4183
rect 9092 4125 9134 4163
rect 9184 4183 9228 4225
rect 9184 4163 9196 4183
rect 9216 4163 9228 4183
rect 9184 4125 9228 4163
rect 9300 4183 9342 4225
rect 9300 4163 9308 4183
rect 9328 4163 9342 4183
rect 9300 4125 9342 4163
rect 9392 4183 9436 4225
rect 9392 4163 9404 4183
rect 9424 4163 9436 4183
rect 9392 4125 9436 4163
rect 9513 4183 9555 4225
rect 9513 4163 9521 4183
rect 9541 4163 9555 4183
rect 9513 4125 9555 4163
rect 9605 4183 9649 4225
rect 9605 4163 9617 4183
rect 9637 4163 9649 4183
rect 10370 4207 10414 4245
rect 10370 4187 10382 4207
rect 10402 4187 10414 4207
rect 9605 4125 9649 4163
rect 10370 4145 10414 4187
rect 10464 4207 10506 4245
rect 10464 4187 10478 4207
rect 10498 4187 10506 4207
rect 10464 4145 10506 4187
rect 10583 4207 10627 4245
rect 10583 4187 10595 4207
rect 10615 4187 10627 4207
rect 10583 4145 10627 4187
rect 10677 4207 10719 4245
rect 10677 4187 10691 4207
rect 10711 4187 10719 4207
rect 10677 4145 10719 4187
rect 10791 4207 10835 4245
rect 10791 4187 10803 4207
rect 10823 4187 10835 4207
rect 10791 4145 10835 4187
rect 10885 4207 10927 4245
rect 10885 4187 10899 4207
rect 10919 4187 10927 4207
rect 10885 4145 10927 4187
rect 11001 4207 11043 4245
rect 11001 4187 11009 4207
rect 11029 4187 11043 4207
rect 11001 4145 11043 4187
rect 11093 4214 11138 4245
rect 11093 4207 11137 4214
rect 11093 4187 11105 4207
rect 11125 4187 11137 4207
rect 15426 4248 15470 4286
rect 15426 4228 15438 4248
rect 15458 4228 15470 4248
rect 11093 4145 11137 4187
rect 13857 4147 13901 4189
rect 13857 4127 13869 4147
rect 13889 4127 13901 4147
rect 13857 4120 13901 4127
rect 13856 4089 13901 4120
rect 13951 4147 13993 4189
rect 13951 4127 13965 4147
rect 13985 4127 13993 4147
rect 13951 4089 13993 4127
rect 14067 4147 14109 4189
rect 14067 4127 14075 4147
rect 14095 4127 14109 4147
rect 14067 4089 14109 4127
rect 14159 4147 14203 4189
rect 14159 4127 14171 4147
rect 14191 4127 14203 4147
rect 14159 4089 14203 4127
rect 14275 4147 14317 4189
rect 14275 4127 14283 4147
rect 14303 4127 14317 4147
rect 14275 4089 14317 4127
rect 14367 4147 14411 4189
rect 14367 4127 14379 4147
rect 14399 4127 14411 4147
rect 14367 4089 14411 4127
rect 14488 4147 14530 4189
rect 14488 4127 14496 4147
rect 14516 4127 14530 4147
rect 14488 4089 14530 4127
rect 14580 4147 14624 4189
rect 15426 4186 15470 4228
rect 15520 4248 15562 4286
rect 15520 4228 15534 4248
rect 15554 4228 15562 4248
rect 15520 4186 15562 4228
rect 15639 4248 15683 4286
rect 15639 4228 15651 4248
rect 15671 4228 15683 4248
rect 15639 4186 15683 4228
rect 15733 4248 15775 4286
rect 15733 4228 15747 4248
rect 15767 4228 15775 4248
rect 15733 4186 15775 4228
rect 15847 4248 15891 4286
rect 15847 4228 15859 4248
rect 15879 4228 15891 4248
rect 15847 4186 15891 4228
rect 15941 4248 15983 4286
rect 15941 4228 15955 4248
rect 15975 4228 15983 4248
rect 15941 4186 15983 4228
rect 16057 4248 16099 4286
rect 16057 4228 16065 4248
rect 16085 4228 16099 4248
rect 16057 4186 16099 4228
rect 16149 4255 16194 4286
rect 16149 4248 16193 4255
rect 16149 4228 16161 4248
rect 16181 4228 16193 4248
rect 16149 4186 16193 4228
rect 18913 4188 18957 4230
rect 14580 4127 14592 4147
rect 14612 4127 14624 4147
rect 14580 4089 14624 4127
rect 18913 4168 18925 4188
rect 18945 4168 18957 4188
rect 18913 4161 18957 4168
rect 18912 4130 18957 4161
rect 19007 4188 19049 4230
rect 19007 4168 19021 4188
rect 19041 4168 19049 4188
rect 19007 4130 19049 4168
rect 19123 4188 19165 4230
rect 19123 4168 19131 4188
rect 19151 4168 19165 4188
rect 19123 4130 19165 4168
rect 19215 4188 19259 4230
rect 19215 4168 19227 4188
rect 19247 4168 19259 4188
rect 19215 4130 19259 4168
rect 19331 4188 19373 4230
rect 19331 4168 19339 4188
rect 19359 4168 19373 4188
rect 19331 4130 19373 4168
rect 19423 4188 19467 4230
rect 19423 4168 19435 4188
rect 19455 4168 19467 4188
rect 19423 4130 19467 4168
rect 19544 4188 19586 4230
rect 19544 4168 19552 4188
rect 19572 4168 19586 4188
rect 19544 4130 19586 4168
rect 19636 4188 19680 4230
rect 19636 4168 19648 4188
rect 19668 4168 19680 4188
rect 19636 4130 19680 4168
rect 1419 3920 1463 3958
rect 1419 3900 1431 3920
rect 1451 3900 1463 3920
rect 1419 3858 1463 3900
rect 1513 3920 1555 3958
rect 1513 3900 1527 3920
rect 1547 3900 1555 3920
rect 1513 3858 1555 3900
rect 1632 3920 1676 3958
rect 1632 3900 1644 3920
rect 1664 3900 1676 3920
rect 1632 3858 1676 3900
rect 1726 3920 1768 3958
rect 1726 3900 1740 3920
rect 1760 3900 1768 3920
rect 1726 3858 1768 3900
rect 1840 3920 1884 3958
rect 1840 3900 1852 3920
rect 1872 3900 1884 3920
rect 1840 3858 1884 3900
rect 1934 3920 1976 3958
rect 1934 3900 1948 3920
rect 1968 3900 1976 3920
rect 1934 3858 1976 3900
rect 2050 3920 2092 3958
rect 2050 3900 2058 3920
rect 2078 3900 2092 3920
rect 2050 3858 2092 3900
rect 2142 3927 2187 3958
rect 2142 3920 2186 3927
rect 2142 3900 2154 3920
rect 2174 3900 2186 3920
rect 6475 3961 6519 3999
rect 6475 3941 6487 3961
rect 6507 3941 6519 3961
rect 2142 3858 2186 3900
rect 2748 3875 2792 3917
rect 2748 3855 2760 3875
rect 2780 3855 2792 3875
rect 2748 3848 2792 3855
rect 2747 3817 2792 3848
rect 2842 3875 2884 3917
rect 2842 3855 2856 3875
rect 2876 3855 2884 3875
rect 2842 3817 2884 3855
rect 2958 3875 3000 3917
rect 2958 3855 2966 3875
rect 2986 3855 3000 3875
rect 2958 3817 3000 3855
rect 3050 3875 3094 3917
rect 3050 3855 3062 3875
rect 3082 3855 3094 3875
rect 3050 3817 3094 3855
rect 3166 3875 3208 3917
rect 3166 3855 3174 3875
rect 3194 3855 3208 3875
rect 3166 3817 3208 3855
rect 3258 3875 3302 3917
rect 3258 3855 3270 3875
rect 3290 3855 3302 3875
rect 3258 3817 3302 3855
rect 3379 3875 3421 3917
rect 3379 3855 3387 3875
rect 3407 3855 3421 3875
rect 3379 3817 3421 3855
rect 3471 3875 3515 3917
rect 6475 3899 6519 3941
rect 6569 3961 6611 3999
rect 6569 3941 6583 3961
rect 6603 3941 6611 3961
rect 6569 3899 6611 3941
rect 6688 3961 6732 3999
rect 6688 3941 6700 3961
rect 6720 3941 6732 3961
rect 6688 3899 6732 3941
rect 6782 3961 6824 3999
rect 6782 3941 6796 3961
rect 6816 3941 6824 3961
rect 6782 3899 6824 3941
rect 6896 3961 6940 3999
rect 6896 3941 6908 3961
rect 6928 3941 6940 3961
rect 6896 3899 6940 3941
rect 6990 3961 7032 3999
rect 6990 3941 7004 3961
rect 7024 3941 7032 3961
rect 6990 3899 7032 3941
rect 7106 3961 7148 3999
rect 7106 3941 7114 3961
rect 7134 3941 7148 3961
rect 7106 3899 7148 3941
rect 7198 3968 7243 3999
rect 7198 3961 7242 3968
rect 7198 3941 7210 3961
rect 7230 3941 7242 3961
rect 7198 3899 7242 3941
rect 7804 3916 7848 3958
rect 3471 3855 3483 3875
rect 3503 3855 3515 3875
rect 3471 3817 3515 3855
rect 7804 3896 7816 3916
rect 7836 3896 7848 3916
rect 7804 3889 7848 3896
rect 7803 3858 7848 3889
rect 7898 3916 7940 3958
rect 7898 3896 7912 3916
rect 7932 3896 7940 3916
rect 7898 3858 7940 3896
rect 8014 3916 8056 3958
rect 8014 3896 8022 3916
rect 8042 3896 8056 3916
rect 8014 3858 8056 3896
rect 8106 3916 8150 3958
rect 8106 3896 8118 3916
rect 8138 3896 8150 3916
rect 8106 3858 8150 3896
rect 8222 3916 8264 3958
rect 8222 3896 8230 3916
rect 8250 3896 8264 3916
rect 8222 3858 8264 3896
rect 8314 3916 8358 3958
rect 8314 3896 8326 3916
rect 8346 3896 8358 3916
rect 8314 3858 8358 3896
rect 8435 3916 8477 3958
rect 8435 3896 8443 3916
rect 8463 3896 8477 3916
rect 8435 3858 8477 3896
rect 8527 3916 8571 3958
rect 8527 3896 8539 3916
rect 8559 3896 8571 3916
rect 8527 3858 8571 3896
rect 11450 3925 11494 3963
rect 11450 3905 11462 3925
rect 11482 3905 11494 3925
rect 11450 3863 11494 3905
rect 11544 3925 11586 3963
rect 11544 3905 11558 3925
rect 11578 3905 11586 3925
rect 11544 3863 11586 3905
rect 11663 3925 11707 3963
rect 11663 3905 11675 3925
rect 11695 3905 11707 3925
rect 11663 3863 11707 3905
rect 11757 3925 11799 3963
rect 11757 3905 11771 3925
rect 11791 3905 11799 3925
rect 11757 3863 11799 3905
rect 11871 3925 11915 3963
rect 11871 3905 11883 3925
rect 11903 3905 11915 3925
rect 11871 3863 11915 3905
rect 11965 3925 12007 3963
rect 11965 3905 11979 3925
rect 11999 3905 12007 3925
rect 11965 3863 12007 3905
rect 12081 3925 12123 3963
rect 12081 3905 12089 3925
rect 12109 3905 12123 3925
rect 12081 3863 12123 3905
rect 12173 3932 12218 3963
rect 12173 3925 12217 3932
rect 12173 3905 12185 3925
rect 12205 3905 12217 3925
rect 16506 3966 16550 4004
rect 16506 3946 16518 3966
rect 16538 3946 16550 3966
rect 12173 3863 12217 3905
rect 12779 3880 12823 3922
rect 12779 3860 12791 3880
rect 12811 3860 12823 3880
rect 12779 3853 12823 3860
rect 12778 3822 12823 3853
rect 12873 3880 12915 3922
rect 12873 3860 12887 3880
rect 12907 3860 12915 3880
rect 12873 3822 12915 3860
rect 12989 3880 13031 3922
rect 12989 3860 12997 3880
rect 13017 3860 13031 3880
rect 12989 3822 13031 3860
rect 13081 3880 13125 3922
rect 13081 3860 13093 3880
rect 13113 3860 13125 3880
rect 13081 3822 13125 3860
rect 13197 3880 13239 3922
rect 13197 3860 13205 3880
rect 13225 3860 13239 3880
rect 13197 3822 13239 3860
rect 13289 3880 13333 3922
rect 13289 3860 13301 3880
rect 13321 3860 13333 3880
rect 13289 3822 13333 3860
rect 13410 3880 13452 3922
rect 13410 3860 13418 3880
rect 13438 3860 13452 3880
rect 13410 3822 13452 3860
rect 13502 3880 13546 3922
rect 16506 3904 16550 3946
rect 16600 3966 16642 4004
rect 16600 3946 16614 3966
rect 16634 3946 16642 3966
rect 16600 3904 16642 3946
rect 16719 3966 16763 4004
rect 16719 3946 16731 3966
rect 16751 3946 16763 3966
rect 16719 3904 16763 3946
rect 16813 3966 16855 4004
rect 16813 3946 16827 3966
rect 16847 3946 16855 3966
rect 16813 3904 16855 3946
rect 16927 3966 16971 4004
rect 16927 3946 16939 3966
rect 16959 3946 16971 3966
rect 16927 3904 16971 3946
rect 17021 3966 17063 4004
rect 17021 3946 17035 3966
rect 17055 3946 17063 3966
rect 17021 3904 17063 3946
rect 17137 3966 17179 4004
rect 17137 3946 17145 3966
rect 17165 3946 17179 3966
rect 17137 3904 17179 3946
rect 17229 3973 17274 4004
rect 17229 3966 17273 3973
rect 17229 3946 17241 3966
rect 17261 3946 17273 3966
rect 17229 3904 17273 3946
rect 17835 3921 17879 3963
rect 13502 3860 13514 3880
rect 13534 3860 13546 3880
rect 13502 3822 13546 3860
rect 17835 3901 17847 3921
rect 17867 3901 17879 3921
rect 17835 3894 17879 3901
rect 17834 3863 17879 3894
rect 17929 3921 17971 3963
rect 17929 3901 17943 3921
rect 17963 3901 17971 3921
rect 17929 3863 17971 3901
rect 18045 3921 18087 3963
rect 18045 3901 18053 3921
rect 18073 3901 18087 3921
rect 18045 3863 18087 3901
rect 18137 3921 18181 3963
rect 18137 3901 18149 3921
rect 18169 3901 18181 3921
rect 18137 3863 18181 3901
rect 18253 3921 18295 3963
rect 18253 3901 18261 3921
rect 18281 3901 18295 3921
rect 18253 3863 18295 3901
rect 18345 3921 18389 3963
rect 18345 3901 18357 3921
rect 18377 3901 18389 3921
rect 18345 3863 18389 3901
rect 18466 3921 18508 3963
rect 18466 3901 18474 3921
rect 18494 3901 18508 3921
rect 18466 3863 18508 3901
rect 18558 3921 18602 3963
rect 18558 3901 18570 3921
rect 18590 3901 18602 3921
rect 18558 3863 18602 3901
rect 341 3653 385 3691
rect 341 3633 353 3653
rect 373 3633 385 3653
rect 341 3591 385 3633
rect 435 3653 477 3691
rect 435 3633 449 3653
rect 469 3633 477 3653
rect 435 3591 477 3633
rect 554 3653 598 3691
rect 554 3633 566 3653
rect 586 3633 598 3653
rect 554 3591 598 3633
rect 648 3653 690 3691
rect 648 3633 662 3653
rect 682 3633 690 3653
rect 648 3591 690 3633
rect 762 3653 806 3691
rect 762 3633 774 3653
rect 794 3633 806 3653
rect 762 3591 806 3633
rect 856 3653 898 3691
rect 856 3633 870 3653
rect 890 3633 898 3653
rect 856 3591 898 3633
rect 972 3653 1014 3691
rect 972 3633 980 3653
rect 1000 3633 1014 3653
rect 972 3591 1014 3633
rect 1064 3660 1109 3691
rect 1064 3653 1108 3660
rect 1064 3633 1076 3653
rect 1096 3633 1108 3653
rect 5397 3694 5441 3732
rect 5397 3674 5409 3694
rect 5429 3674 5441 3694
rect 1064 3591 1108 3633
rect 3828 3593 3872 3635
rect 3828 3573 3840 3593
rect 3860 3573 3872 3593
rect 3828 3566 3872 3573
rect 3827 3535 3872 3566
rect 3922 3593 3964 3635
rect 3922 3573 3936 3593
rect 3956 3573 3964 3593
rect 3922 3535 3964 3573
rect 4038 3593 4080 3635
rect 4038 3573 4046 3593
rect 4066 3573 4080 3593
rect 4038 3535 4080 3573
rect 4130 3593 4174 3635
rect 4130 3573 4142 3593
rect 4162 3573 4174 3593
rect 4130 3535 4174 3573
rect 4246 3593 4288 3635
rect 4246 3573 4254 3593
rect 4274 3573 4288 3593
rect 4246 3535 4288 3573
rect 4338 3593 4382 3635
rect 4338 3573 4350 3593
rect 4370 3573 4382 3593
rect 4338 3535 4382 3573
rect 4459 3593 4501 3635
rect 4459 3573 4467 3593
rect 4487 3573 4501 3593
rect 4459 3535 4501 3573
rect 4551 3593 4595 3635
rect 5397 3632 5441 3674
rect 5491 3694 5533 3732
rect 5491 3674 5505 3694
rect 5525 3674 5533 3694
rect 5491 3632 5533 3674
rect 5610 3694 5654 3732
rect 5610 3674 5622 3694
rect 5642 3674 5654 3694
rect 5610 3632 5654 3674
rect 5704 3694 5746 3732
rect 5704 3674 5718 3694
rect 5738 3674 5746 3694
rect 5704 3632 5746 3674
rect 5818 3694 5862 3732
rect 5818 3674 5830 3694
rect 5850 3674 5862 3694
rect 5818 3632 5862 3674
rect 5912 3694 5954 3732
rect 5912 3674 5926 3694
rect 5946 3674 5954 3694
rect 5912 3632 5954 3674
rect 6028 3694 6070 3732
rect 6028 3674 6036 3694
rect 6056 3674 6070 3694
rect 6028 3632 6070 3674
rect 6120 3701 6165 3732
rect 6120 3694 6164 3701
rect 6120 3674 6132 3694
rect 6152 3674 6164 3694
rect 6120 3632 6164 3674
rect 8884 3634 8928 3676
rect 4551 3573 4563 3593
rect 4583 3573 4595 3593
rect 4551 3535 4595 3573
rect 8884 3614 8896 3634
rect 8916 3614 8928 3634
rect 8884 3607 8928 3614
rect 8883 3576 8928 3607
rect 8978 3634 9020 3676
rect 8978 3614 8992 3634
rect 9012 3614 9020 3634
rect 8978 3576 9020 3614
rect 9094 3634 9136 3676
rect 9094 3614 9102 3634
rect 9122 3614 9136 3634
rect 9094 3576 9136 3614
rect 9186 3634 9230 3676
rect 9186 3614 9198 3634
rect 9218 3614 9230 3634
rect 9186 3576 9230 3614
rect 9302 3634 9344 3676
rect 9302 3614 9310 3634
rect 9330 3614 9344 3634
rect 9302 3576 9344 3614
rect 9394 3634 9438 3676
rect 9394 3614 9406 3634
rect 9426 3614 9438 3634
rect 9394 3576 9438 3614
rect 9515 3634 9557 3676
rect 9515 3614 9523 3634
rect 9543 3614 9557 3634
rect 9515 3576 9557 3614
rect 9607 3634 9651 3676
rect 10372 3658 10416 3696
rect 9607 3614 9619 3634
rect 9639 3614 9651 3634
rect 9607 3576 9651 3614
rect 10372 3638 10384 3658
rect 10404 3638 10416 3658
rect 10372 3596 10416 3638
rect 10466 3658 10508 3696
rect 10466 3638 10480 3658
rect 10500 3638 10508 3658
rect 10466 3596 10508 3638
rect 10585 3658 10629 3696
rect 10585 3638 10597 3658
rect 10617 3638 10629 3658
rect 10585 3596 10629 3638
rect 10679 3658 10721 3696
rect 10679 3638 10693 3658
rect 10713 3638 10721 3658
rect 10679 3596 10721 3638
rect 10793 3658 10837 3696
rect 10793 3638 10805 3658
rect 10825 3638 10837 3658
rect 10793 3596 10837 3638
rect 10887 3658 10929 3696
rect 10887 3638 10901 3658
rect 10921 3638 10929 3658
rect 10887 3596 10929 3638
rect 11003 3658 11045 3696
rect 11003 3638 11011 3658
rect 11031 3638 11045 3658
rect 11003 3596 11045 3638
rect 11095 3665 11140 3696
rect 11095 3658 11139 3665
rect 11095 3638 11107 3658
rect 11127 3638 11139 3658
rect 15428 3699 15472 3737
rect 15428 3679 15440 3699
rect 15460 3679 15472 3699
rect 11095 3596 11139 3638
rect 13859 3598 13903 3640
rect 1279 3409 1323 3447
rect 1279 3389 1291 3409
rect 1311 3389 1323 3409
rect 1279 3347 1323 3389
rect 1373 3409 1415 3447
rect 1373 3389 1387 3409
rect 1407 3389 1415 3409
rect 1373 3347 1415 3389
rect 1492 3409 1536 3447
rect 1492 3389 1504 3409
rect 1524 3389 1536 3409
rect 1492 3347 1536 3389
rect 1586 3409 1628 3447
rect 1586 3389 1600 3409
rect 1620 3389 1628 3409
rect 1586 3347 1628 3389
rect 1700 3409 1744 3447
rect 1700 3389 1712 3409
rect 1732 3389 1744 3409
rect 1700 3347 1744 3389
rect 1794 3409 1836 3447
rect 1794 3389 1808 3409
rect 1828 3389 1836 3409
rect 1794 3347 1836 3389
rect 1910 3409 1952 3447
rect 1910 3389 1918 3409
rect 1938 3389 1952 3409
rect 1910 3347 1952 3389
rect 2002 3416 2047 3447
rect 2002 3409 2046 3416
rect 2002 3389 2014 3409
rect 2034 3389 2046 3409
rect 2002 3347 2046 3389
rect 6335 3450 6379 3488
rect 6335 3430 6347 3450
rect 6367 3430 6379 3450
rect 2889 3283 2933 3325
rect 2889 3263 2901 3283
rect 2921 3263 2933 3283
rect 2889 3256 2933 3263
rect 2888 3225 2933 3256
rect 2983 3283 3025 3325
rect 2983 3263 2997 3283
rect 3017 3263 3025 3283
rect 2983 3225 3025 3263
rect 3099 3283 3141 3325
rect 3099 3263 3107 3283
rect 3127 3263 3141 3283
rect 3099 3225 3141 3263
rect 3191 3283 3235 3325
rect 3191 3263 3203 3283
rect 3223 3263 3235 3283
rect 3191 3225 3235 3263
rect 3307 3283 3349 3325
rect 3307 3263 3315 3283
rect 3335 3263 3349 3283
rect 3307 3225 3349 3263
rect 3399 3283 3443 3325
rect 3399 3263 3411 3283
rect 3431 3263 3443 3283
rect 3399 3225 3443 3263
rect 3520 3283 3562 3325
rect 3520 3263 3528 3283
rect 3548 3263 3562 3283
rect 3520 3225 3562 3263
rect 3612 3283 3656 3325
rect 6335 3388 6379 3430
rect 6429 3450 6471 3488
rect 6429 3430 6443 3450
rect 6463 3430 6471 3450
rect 6429 3388 6471 3430
rect 6548 3450 6592 3488
rect 6548 3430 6560 3450
rect 6580 3430 6592 3450
rect 6548 3388 6592 3430
rect 6642 3450 6684 3488
rect 6642 3430 6656 3450
rect 6676 3430 6684 3450
rect 6642 3388 6684 3430
rect 6756 3450 6800 3488
rect 6756 3430 6768 3450
rect 6788 3430 6800 3450
rect 6756 3388 6800 3430
rect 6850 3450 6892 3488
rect 6850 3430 6864 3450
rect 6884 3430 6892 3450
rect 6850 3388 6892 3430
rect 6966 3450 7008 3488
rect 6966 3430 6974 3450
rect 6994 3430 7008 3450
rect 6966 3388 7008 3430
rect 7058 3457 7103 3488
rect 13859 3578 13871 3598
rect 13891 3578 13903 3598
rect 13859 3571 13903 3578
rect 7058 3450 7102 3457
rect 7058 3430 7070 3450
rect 7090 3430 7102 3450
rect 13858 3540 13903 3571
rect 13953 3598 13995 3640
rect 13953 3578 13967 3598
rect 13987 3578 13995 3598
rect 13953 3540 13995 3578
rect 14069 3598 14111 3640
rect 14069 3578 14077 3598
rect 14097 3578 14111 3598
rect 14069 3540 14111 3578
rect 14161 3598 14205 3640
rect 14161 3578 14173 3598
rect 14193 3578 14205 3598
rect 14161 3540 14205 3578
rect 14277 3598 14319 3640
rect 14277 3578 14285 3598
rect 14305 3578 14319 3598
rect 14277 3540 14319 3578
rect 14369 3598 14413 3640
rect 14369 3578 14381 3598
rect 14401 3578 14413 3598
rect 14369 3540 14413 3578
rect 14490 3598 14532 3640
rect 14490 3578 14498 3598
rect 14518 3578 14532 3598
rect 14490 3540 14532 3578
rect 14582 3598 14626 3640
rect 15428 3637 15472 3679
rect 15522 3699 15564 3737
rect 15522 3679 15536 3699
rect 15556 3679 15564 3699
rect 15522 3637 15564 3679
rect 15641 3699 15685 3737
rect 15641 3679 15653 3699
rect 15673 3679 15685 3699
rect 15641 3637 15685 3679
rect 15735 3699 15777 3737
rect 15735 3679 15749 3699
rect 15769 3679 15777 3699
rect 15735 3637 15777 3679
rect 15849 3699 15893 3737
rect 15849 3679 15861 3699
rect 15881 3679 15893 3699
rect 15849 3637 15893 3679
rect 15943 3699 15985 3737
rect 15943 3679 15957 3699
rect 15977 3679 15985 3699
rect 15943 3637 15985 3679
rect 16059 3699 16101 3737
rect 16059 3679 16067 3699
rect 16087 3679 16101 3699
rect 16059 3637 16101 3679
rect 16151 3706 16196 3737
rect 16151 3699 16195 3706
rect 16151 3679 16163 3699
rect 16183 3679 16195 3699
rect 16151 3637 16195 3679
rect 18915 3639 18959 3681
rect 14582 3578 14594 3598
rect 14614 3578 14626 3598
rect 14582 3540 14626 3578
rect 18915 3619 18927 3639
rect 18947 3619 18959 3639
rect 18915 3612 18959 3619
rect 18914 3581 18959 3612
rect 19009 3639 19051 3681
rect 19009 3619 19023 3639
rect 19043 3619 19051 3639
rect 19009 3581 19051 3619
rect 19125 3639 19167 3681
rect 19125 3619 19133 3639
rect 19153 3619 19167 3639
rect 19125 3581 19167 3619
rect 19217 3639 19261 3681
rect 19217 3619 19229 3639
rect 19249 3619 19261 3639
rect 19217 3581 19261 3619
rect 19333 3639 19375 3681
rect 19333 3619 19341 3639
rect 19361 3619 19375 3639
rect 19333 3581 19375 3619
rect 19425 3639 19469 3681
rect 19425 3619 19437 3639
rect 19457 3619 19469 3639
rect 19425 3581 19469 3619
rect 19546 3639 19588 3681
rect 19546 3619 19554 3639
rect 19574 3619 19588 3639
rect 19546 3581 19588 3619
rect 19638 3639 19682 3681
rect 19638 3619 19650 3639
rect 19670 3619 19682 3639
rect 19638 3581 19682 3619
rect 7058 3388 7102 3430
rect 3612 3263 3624 3283
rect 3644 3263 3656 3283
rect 3612 3225 3656 3263
rect 7945 3324 7989 3366
rect 7945 3304 7957 3324
rect 7977 3304 7989 3324
rect 7945 3297 7989 3304
rect 7944 3266 7989 3297
rect 8039 3324 8081 3366
rect 8039 3304 8053 3324
rect 8073 3304 8081 3324
rect 8039 3266 8081 3304
rect 8155 3324 8197 3366
rect 8155 3304 8163 3324
rect 8183 3304 8197 3324
rect 8155 3266 8197 3304
rect 8247 3324 8291 3366
rect 8247 3304 8259 3324
rect 8279 3304 8291 3324
rect 8247 3266 8291 3304
rect 8363 3324 8405 3366
rect 8363 3304 8371 3324
rect 8391 3304 8405 3324
rect 8363 3266 8405 3304
rect 8455 3324 8499 3366
rect 8455 3304 8467 3324
rect 8487 3304 8499 3324
rect 8455 3266 8499 3304
rect 8576 3324 8618 3366
rect 8576 3304 8584 3324
rect 8604 3304 8618 3324
rect 8576 3266 8618 3304
rect 8668 3324 8712 3366
rect 11310 3414 11354 3452
rect 11310 3394 11322 3414
rect 11342 3394 11354 3414
rect 8668 3304 8680 3324
rect 8700 3304 8712 3324
rect 8668 3266 8712 3304
rect 11310 3352 11354 3394
rect 11404 3414 11446 3452
rect 11404 3394 11418 3414
rect 11438 3394 11446 3414
rect 11404 3352 11446 3394
rect 11523 3414 11567 3452
rect 11523 3394 11535 3414
rect 11555 3394 11567 3414
rect 11523 3352 11567 3394
rect 11617 3414 11659 3452
rect 11617 3394 11631 3414
rect 11651 3394 11659 3414
rect 11617 3352 11659 3394
rect 11731 3414 11775 3452
rect 11731 3394 11743 3414
rect 11763 3394 11775 3414
rect 11731 3352 11775 3394
rect 11825 3414 11867 3452
rect 11825 3394 11839 3414
rect 11859 3394 11867 3414
rect 11825 3352 11867 3394
rect 11941 3414 11983 3452
rect 11941 3394 11949 3414
rect 11969 3394 11983 3414
rect 11941 3352 11983 3394
rect 12033 3421 12078 3452
rect 12033 3414 12077 3421
rect 12033 3394 12045 3414
rect 12065 3394 12077 3414
rect 12033 3352 12077 3394
rect 16366 3455 16410 3493
rect 16366 3435 16378 3455
rect 16398 3435 16410 3455
rect 12920 3288 12964 3330
rect 340 3099 384 3137
rect 340 3079 352 3099
rect 372 3079 384 3099
rect 340 3037 384 3079
rect 434 3099 476 3137
rect 434 3079 448 3099
rect 468 3079 476 3099
rect 434 3037 476 3079
rect 553 3099 597 3137
rect 553 3079 565 3099
rect 585 3079 597 3099
rect 553 3037 597 3079
rect 647 3099 689 3137
rect 647 3079 661 3099
rect 681 3079 689 3099
rect 647 3037 689 3079
rect 761 3099 805 3137
rect 761 3079 773 3099
rect 793 3079 805 3099
rect 761 3037 805 3079
rect 855 3099 897 3137
rect 855 3079 869 3099
rect 889 3079 897 3099
rect 855 3037 897 3079
rect 971 3099 1013 3137
rect 971 3079 979 3099
rect 999 3079 1013 3099
rect 971 3037 1013 3079
rect 1063 3106 1108 3137
rect 1063 3099 1107 3106
rect 1063 3079 1075 3099
rect 1095 3079 1107 3099
rect 5396 3140 5440 3178
rect 5396 3120 5408 3140
rect 5428 3120 5440 3140
rect 1063 3037 1107 3079
rect 3827 3039 3871 3081
rect 3827 3019 3839 3039
rect 3859 3019 3871 3039
rect 3827 3012 3871 3019
rect 3826 2981 3871 3012
rect 3921 3039 3963 3081
rect 3921 3019 3935 3039
rect 3955 3019 3963 3039
rect 3921 2981 3963 3019
rect 4037 3039 4079 3081
rect 4037 3019 4045 3039
rect 4065 3019 4079 3039
rect 4037 2981 4079 3019
rect 4129 3039 4173 3081
rect 4129 3019 4141 3039
rect 4161 3019 4173 3039
rect 4129 2981 4173 3019
rect 4245 3039 4287 3081
rect 4245 3019 4253 3039
rect 4273 3019 4287 3039
rect 4245 2981 4287 3019
rect 4337 3039 4381 3081
rect 4337 3019 4349 3039
rect 4369 3019 4381 3039
rect 4337 2981 4381 3019
rect 4458 3039 4500 3081
rect 4458 3019 4466 3039
rect 4486 3019 4500 3039
rect 4458 2981 4500 3019
rect 4550 3039 4594 3081
rect 5396 3078 5440 3120
rect 5490 3140 5532 3178
rect 5490 3120 5504 3140
rect 5524 3120 5532 3140
rect 5490 3078 5532 3120
rect 5609 3140 5653 3178
rect 5609 3120 5621 3140
rect 5641 3120 5653 3140
rect 5609 3078 5653 3120
rect 5703 3140 5745 3178
rect 5703 3120 5717 3140
rect 5737 3120 5745 3140
rect 5703 3078 5745 3120
rect 5817 3140 5861 3178
rect 5817 3120 5829 3140
rect 5849 3120 5861 3140
rect 5817 3078 5861 3120
rect 5911 3140 5953 3178
rect 5911 3120 5925 3140
rect 5945 3120 5953 3140
rect 5911 3078 5953 3120
rect 6027 3140 6069 3178
rect 6027 3120 6035 3140
rect 6055 3120 6069 3140
rect 6027 3078 6069 3120
rect 6119 3147 6164 3178
rect 12920 3268 12932 3288
rect 12952 3268 12964 3288
rect 12920 3261 12964 3268
rect 6119 3140 6163 3147
rect 6119 3120 6131 3140
rect 6151 3120 6163 3140
rect 12919 3230 12964 3261
rect 13014 3288 13056 3330
rect 13014 3268 13028 3288
rect 13048 3268 13056 3288
rect 13014 3230 13056 3268
rect 13130 3288 13172 3330
rect 13130 3268 13138 3288
rect 13158 3268 13172 3288
rect 13130 3230 13172 3268
rect 13222 3288 13266 3330
rect 13222 3268 13234 3288
rect 13254 3268 13266 3288
rect 13222 3230 13266 3268
rect 13338 3288 13380 3330
rect 13338 3268 13346 3288
rect 13366 3268 13380 3288
rect 13338 3230 13380 3268
rect 13430 3288 13474 3330
rect 13430 3268 13442 3288
rect 13462 3268 13474 3288
rect 13430 3230 13474 3268
rect 13551 3288 13593 3330
rect 13551 3268 13559 3288
rect 13579 3268 13593 3288
rect 13551 3230 13593 3268
rect 13643 3288 13687 3330
rect 16366 3393 16410 3435
rect 16460 3455 16502 3493
rect 16460 3435 16474 3455
rect 16494 3435 16502 3455
rect 16460 3393 16502 3435
rect 16579 3455 16623 3493
rect 16579 3435 16591 3455
rect 16611 3435 16623 3455
rect 16579 3393 16623 3435
rect 16673 3455 16715 3493
rect 16673 3435 16687 3455
rect 16707 3435 16715 3455
rect 16673 3393 16715 3435
rect 16787 3455 16831 3493
rect 16787 3435 16799 3455
rect 16819 3435 16831 3455
rect 16787 3393 16831 3435
rect 16881 3455 16923 3493
rect 16881 3435 16895 3455
rect 16915 3435 16923 3455
rect 16881 3393 16923 3435
rect 16997 3455 17039 3493
rect 16997 3435 17005 3455
rect 17025 3435 17039 3455
rect 16997 3393 17039 3435
rect 17089 3462 17134 3493
rect 17089 3455 17133 3462
rect 17089 3435 17101 3455
rect 17121 3435 17133 3455
rect 17089 3393 17133 3435
rect 13643 3268 13655 3288
rect 13675 3268 13687 3288
rect 13643 3230 13687 3268
rect 17976 3329 18020 3371
rect 17976 3309 17988 3329
rect 18008 3309 18020 3329
rect 17976 3302 18020 3309
rect 17975 3271 18020 3302
rect 18070 3329 18112 3371
rect 18070 3309 18084 3329
rect 18104 3309 18112 3329
rect 18070 3271 18112 3309
rect 18186 3329 18228 3371
rect 18186 3309 18194 3329
rect 18214 3309 18228 3329
rect 18186 3271 18228 3309
rect 18278 3329 18322 3371
rect 18278 3309 18290 3329
rect 18310 3309 18322 3329
rect 18278 3271 18322 3309
rect 18394 3329 18436 3371
rect 18394 3309 18402 3329
rect 18422 3309 18436 3329
rect 18394 3271 18436 3309
rect 18486 3329 18530 3371
rect 18486 3309 18498 3329
rect 18518 3309 18530 3329
rect 18486 3271 18530 3309
rect 18607 3329 18649 3371
rect 18607 3309 18615 3329
rect 18635 3309 18649 3329
rect 18607 3271 18649 3309
rect 18699 3329 18743 3371
rect 18699 3309 18711 3329
rect 18731 3309 18743 3329
rect 18699 3271 18743 3309
rect 6119 3078 6163 3120
rect 8883 3080 8927 3122
rect 4550 3019 4562 3039
rect 4582 3019 4594 3039
rect 4550 2981 4594 3019
rect 8883 3060 8895 3080
rect 8915 3060 8927 3080
rect 8883 3053 8927 3060
rect 8882 3022 8927 3053
rect 8977 3080 9019 3122
rect 8977 3060 8991 3080
rect 9011 3060 9019 3080
rect 8977 3022 9019 3060
rect 9093 3080 9135 3122
rect 9093 3060 9101 3080
rect 9121 3060 9135 3080
rect 9093 3022 9135 3060
rect 9185 3080 9229 3122
rect 9185 3060 9197 3080
rect 9217 3060 9229 3080
rect 9185 3022 9229 3060
rect 9301 3080 9343 3122
rect 9301 3060 9309 3080
rect 9329 3060 9343 3080
rect 9301 3022 9343 3060
rect 9393 3080 9437 3122
rect 9393 3060 9405 3080
rect 9425 3060 9437 3080
rect 9393 3022 9437 3060
rect 9514 3080 9556 3122
rect 9514 3060 9522 3080
rect 9542 3060 9556 3080
rect 9514 3022 9556 3060
rect 9606 3080 9650 3122
rect 9606 3060 9618 3080
rect 9638 3060 9650 3080
rect 10371 3104 10415 3142
rect 10371 3084 10383 3104
rect 10403 3084 10415 3104
rect 9606 3022 9650 3060
rect 10371 3042 10415 3084
rect 10465 3104 10507 3142
rect 10465 3084 10479 3104
rect 10499 3084 10507 3104
rect 10465 3042 10507 3084
rect 10584 3104 10628 3142
rect 10584 3084 10596 3104
rect 10616 3084 10628 3104
rect 10584 3042 10628 3084
rect 10678 3104 10720 3142
rect 10678 3084 10692 3104
rect 10712 3084 10720 3104
rect 10678 3042 10720 3084
rect 10792 3104 10836 3142
rect 10792 3084 10804 3104
rect 10824 3084 10836 3104
rect 10792 3042 10836 3084
rect 10886 3104 10928 3142
rect 10886 3084 10900 3104
rect 10920 3084 10928 3104
rect 10886 3042 10928 3084
rect 11002 3104 11044 3142
rect 11002 3084 11010 3104
rect 11030 3084 11044 3104
rect 11002 3042 11044 3084
rect 11094 3111 11139 3142
rect 11094 3104 11138 3111
rect 11094 3084 11106 3104
rect 11126 3084 11138 3104
rect 15427 3145 15471 3183
rect 15427 3125 15439 3145
rect 15459 3125 15471 3145
rect 11094 3042 11138 3084
rect 13858 3044 13902 3086
rect 13858 3024 13870 3044
rect 13890 3024 13902 3044
rect 13858 3017 13902 3024
rect 13857 2986 13902 3017
rect 13952 3044 13994 3086
rect 13952 3024 13966 3044
rect 13986 3024 13994 3044
rect 13952 2986 13994 3024
rect 14068 3044 14110 3086
rect 14068 3024 14076 3044
rect 14096 3024 14110 3044
rect 14068 2986 14110 3024
rect 14160 3044 14204 3086
rect 14160 3024 14172 3044
rect 14192 3024 14204 3044
rect 14160 2986 14204 3024
rect 14276 3044 14318 3086
rect 14276 3024 14284 3044
rect 14304 3024 14318 3044
rect 14276 2986 14318 3024
rect 14368 3044 14412 3086
rect 14368 3024 14380 3044
rect 14400 3024 14412 3044
rect 14368 2986 14412 3024
rect 14489 3044 14531 3086
rect 14489 3024 14497 3044
rect 14517 3024 14531 3044
rect 14489 2986 14531 3024
rect 14581 3044 14625 3086
rect 15427 3083 15471 3125
rect 15521 3145 15563 3183
rect 15521 3125 15535 3145
rect 15555 3125 15563 3145
rect 15521 3083 15563 3125
rect 15640 3145 15684 3183
rect 15640 3125 15652 3145
rect 15672 3125 15684 3145
rect 15640 3083 15684 3125
rect 15734 3145 15776 3183
rect 15734 3125 15748 3145
rect 15768 3125 15776 3145
rect 15734 3083 15776 3125
rect 15848 3145 15892 3183
rect 15848 3125 15860 3145
rect 15880 3125 15892 3145
rect 15848 3083 15892 3125
rect 15942 3145 15984 3183
rect 15942 3125 15956 3145
rect 15976 3125 15984 3145
rect 15942 3083 15984 3125
rect 16058 3145 16100 3183
rect 16058 3125 16066 3145
rect 16086 3125 16100 3145
rect 16058 3083 16100 3125
rect 16150 3152 16195 3183
rect 16150 3145 16194 3152
rect 16150 3125 16162 3145
rect 16182 3125 16194 3145
rect 16150 3083 16194 3125
rect 18914 3085 18958 3127
rect 14581 3024 14593 3044
rect 14613 3024 14625 3044
rect 14581 2986 14625 3024
rect 18914 3065 18926 3085
rect 18946 3065 18958 3085
rect 18914 3058 18958 3065
rect 18913 3027 18958 3058
rect 19008 3085 19050 3127
rect 19008 3065 19022 3085
rect 19042 3065 19050 3085
rect 19008 3027 19050 3065
rect 19124 3085 19166 3127
rect 19124 3065 19132 3085
rect 19152 3065 19166 3085
rect 19124 3027 19166 3065
rect 19216 3085 19260 3127
rect 19216 3065 19228 3085
rect 19248 3065 19260 3085
rect 19216 3027 19260 3065
rect 19332 3085 19374 3127
rect 19332 3065 19340 3085
rect 19360 3065 19374 3085
rect 19332 3027 19374 3065
rect 19424 3085 19468 3127
rect 19424 3065 19436 3085
rect 19456 3065 19468 3085
rect 19424 3027 19468 3065
rect 19545 3085 19587 3127
rect 19545 3065 19553 3085
rect 19573 3065 19587 3085
rect 19545 3027 19587 3065
rect 19637 3085 19681 3127
rect 19637 3065 19649 3085
rect 19669 3065 19681 3085
rect 19637 3027 19681 3065
rect 1389 2830 1433 2868
rect 1389 2810 1401 2830
rect 1421 2810 1433 2830
rect 1389 2768 1433 2810
rect 1483 2830 1525 2868
rect 1483 2810 1497 2830
rect 1517 2810 1525 2830
rect 1483 2768 1525 2810
rect 1602 2830 1646 2868
rect 1602 2810 1614 2830
rect 1634 2810 1646 2830
rect 1602 2768 1646 2810
rect 1696 2830 1738 2868
rect 1696 2810 1710 2830
rect 1730 2810 1738 2830
rect 1696 2768 1738 2810
rect 1810 2830 1854 2868
rect 1810 2810 1822 2830
rect 1842 2810 1854 2830
rect 1810 2768 1854 2810
rect 1904 2830 1946 2868
rect 1904 2810 1918 2830
rect 1938 2810 1946 2830
rect 1904 2768 1946 2810
rect 2020 2830 2062 2868
rect 2020 2810 2028 2830
rect 2048 2810 2062 2830
rect 2020 2768 2062 2810
rect 2112 2837 2157 2868
rect 2112 2830 2156 2837
rect 2112 2810 2124 2830
rect 2144 2810 2156 2830
rect 2112 2768 2156 2810
rect 6445 2871 6489 2909
rect 6445 2851 6457 2871
rect 6477 2851 6489 2871
rect 6445 2809 6489 2851
rect 6539 2871 6581 2909
rect 6539 2851 6553 2871
rect 6573 2851 6581 2871
rect 6539 2809 6581 2851
rect 6658 2871 6702 2909
rect 6658 2851 6670 2871
rect 6690 2851 6702 2871
rect 6658 2809 6702 2851
rect 6752 2871 6794 2909
rect 6752 2851 6766 2871
rect 6786 2851 6794 2871
rect 6752 2809 6794 2851
rect 6866 2871 6910 2909
rect 6866 2851 6878 2871
rect 6898 2851 6910 2871
rect 6866 2809 6910 2851
rect 6960 2871 7002 2909
rect 6960 2851 6974 2871
rect 6994 2851 7002 2871
rect 6960 2809 7002 2851
rect 7076 2871 7118 2909
rect 7076 2851 7084 2871
rect 7104 2851 7118 2871
rect 7076 2809 7118 2851
rect 7168 2878 7213 2909
rect 7168 2871 7212 2878
rect 7168 2851 7180 2871
rect 7200 2851 7212 2871
rect 7168 2809 7212 2851
rect 2779 2759 2823 2801
rect 2779 2739 2791 2759
rect 2811 2739 2823 2759
rect 2779 2732 2823 2739
rect 2778 2701 2823 2732
rect 2873 2759 2915 2801
rect 2873 2739 2887 2759
rect 2907 2739 2915 2759
rect 2873 2701 2915 2739
rect 2989 2759 3031 2801
rect 2989 2739 2997 2759
rect 3017 2739 3031 2759
rect 2989 2701 3031 2739
rect 3081 2759 3125 2801
rect 3081 2739 3093 2759
rect 3113 2739 3125 2759
rect 3081 2701 3125 2739
rect 3197 2759 3239 2801
rect 3197 2739 3205 2759
rect 3225 2739 3239 2759
rect 3197 2701 3239 2739
rect 3289 2759 3333 2801
rect 3289 2739 3301 2759
rect 3321 2739 3333 2759
rect 3289 2701 3333 2739
rect 3410 2759 3452 2801
rect 3410 2739 3418 2759
rect 3438 2739 3452 2759
rect 3410 2701 3452 2739
rect 3502 2759 3546 2801
rect 3502 2739 3514 2759
rect 3534 2739 3546 2759
rect 3502 2701 3546 2739
rect 7835 2800 7879 2842
rect 7835 2780 7847 2800
rect 7867 2780 7879 2800
rect 7835 2773 7879 2780
rect 7834 2742 7879 2773
rect 7929 2800 7971 2842
rect 7929 2780 7943 2800
rect 7963 2780 7971 2800
rect 7929 2742 7971 2780
rect 8045 2800 8087 2842
rect 8045 2780 8053 2800
rect 8073 2780 8087 2800
rect 8045 2742 8087 2780
rect 8137 2800 8181 2842
rect 8137 2780 8149 2800
rect 8169 2780 8181 2800
rect 8137 2742 8181 2780
rect 8253 2800 8295 2842
rect 8253 2780 8261 2800
rect 8281 2780 8295 2800
rect 8253 2742 8295 2780
rect 8345 2800 8389 2842
rect 8345 2780 8357 2800
rect 8377 2780 8389 2800
rect 8345 2742 8389 2780
rect 8466 2800 8508 2842
rect 8466 2780 8474 2800
rect 8494 2780 8508 2800
rect 8466 2742 8508 2780
rect 8558 2800 8602 2842
rect 11420 2835 11464 2873
rect 8558 2780 8570 2800
rect 8590 2780 8602 2800
rect 11420 2815 11432 2835
rect 11452 2815 11464 2835
rect 8558 2742 8602 2780
rect 11420 2773 11464 2815
rect 11514 2835 11556 2873
rect 11514 2815 11528 2835
rect 11548 2815 11556 2835
rect 11514 2773 11556 2815
rect 11633 2835 11677 2873
rect 11633 2815 11645 2835
rect 11665 2815 11677 2835
rect 11633 2773 11677 2815
rect 11727 2835 11769 2873
rect 11727 2815 11741 2835
rect 11761 2815 11769 2835
rect 11727 2773 11769 2815
rect 11841 2835 11885 2873
rect 11841 2815 11853 2835
rect 11873 2815 11885 2835
rect 11841 2773 11885 2815
rect 11935 2835 11977 2873
rect 11935 2815 11949 2835
rect 11969 2815 11977 2835
rect 11935 2773 11977 2815
rect 12051 2835 12093 2873
rect 12051 2815 12059 2835
rect 12079 2815 12093 2835
rect 12051 2773 12093 2815
rect 12143 2842 12188 2873
rect 12143 2835 12187 2842
rect 12143 2815 12155 2835
rect 12175 2815 12187 2835
rect 12143 2773 12187 2815
rect 16476 2876 16520 2914
rect 16476 2856 16488 2876
rect 16508 2856 16520 2876
rect 16476 2814 16520 2856
rect 16570 2876 16612 2914
rect 16570 2856 16584 2876
rect 16604 2856 16612 2876
rect 16570 2814 16612 2856
rect 16689 2876 16733 2914
rect 16689 2856 16701 2876
rect 16721 2856 16733 2876
rect 16689 2814 16733 2856
rect 16783 2876 16825 2914
rect 16783 2856 16797 2876
rect 16817 2856 16825 2876
rect 16783 2814 16825 2856
rect 16897 2876 16941 2914
rect 16897 2856 16909 2876
rect 16929 2856 16941 2876
rect 16897 2814 16941 2856
rect 16991 2876 17033 2914
rect 16991 2856 17005 2876
rect 17025 2856 17033 2876
rect 16991 2814 17033 2856
rect 17107 2876 17149 2914
rect 17107 2856 17115 2876
rect 17135 2856 17149 2876
rect 17107 2814 17149 2856
rect 17199 2883 17244 2914
rect 17199 2876 17243 2883
rect 17199 2856 17211 2876
rect 17231 2856 17243 2876
rect 17199 2814 17243 2856
rect 12810 2764 12854 2806
rect 12810 2744 12822 2764
rect 12842 2744 12854 2764
rect 12810 2737 12854 2744
rect 12809 2706 12854 2737
rect 12904 2764 12946 2806
rect 12904 2744 12918 2764
rect 12938 2744 12946 2764
rect 12904 2706 12946 2744
rect 13020 2764 13062 2806
rect 13020 2744 13028 2764
rect 13048 2744 13062 2764
rect 13020 2706 13062 2744
rect 13112 2764 13156 2806
rect 13112 2744 13124 2764
rect 13144 2744 13156 2764
rect 13112 2706 13156 2744
rect 13228 2764 13270 2806
rect 13228 2744 13236 2764
rect 13256 2744 13270 2764
rect 13228 2706 13270 2744
rect 13320 2764 13364 2806
rect 13320 2744 13332 2764
rect 13352 2744 13364 2764
rect 13320 2706 13364 2744
rect 13441 2764 13483 2806
rect 13441 2744 13449 2764
rect 13469 2744 13483 2764
rect 13441 2706 13483 2744
rect 13533 2764 13577 2806
rect 13533 2744 13545 2764
rect 13565 2744 13577 2764
rect 13533 2706 13577 2744
rect 17866 2805 17910 2847
rect 17866 2785 17878 2805
rect 17898 2785 17910 2805
rect 17866 2778 17910 2785
rect 17865 2747 17910 2778
rect 17960 2805 18002 2847
rect 17960 2785 17974 2805
rect 17994 2785 18002 2805
rect 17960 2747 18002 2785
rect 18076 2805 18118 2847
rect 18076 2785 18084 2805
rect 18104 2785 18118 2805
rect 18076 2747 18118 2785
rect 18168 2805 18212 2847
rect 18168 2785 18180 2805
rect 18200 2785 18212 2805
rect 18168 2747 18212 2785
rect 18284 2805 18326 2847
rect 18284 2785 18292 2805
rect 18312 2785 18326 2805
rect 18284 2747 18326 2785
rect 18376 2805 18420 2847
rect 18376 2785 18388 2805
rect 18408 2785 18420 2805
rect 18376 2747 18420 2785
rect 18497 2805 18539 2847
rect 18497 2785 18505 2805
rect 18525 2785 18539 2805
rect 18497 2747 18539 2785
rect 18589 2805 18633 2847
rect 18589 2785 18601 2805
rect 18621 2785 18633 2805
rect 18589 2747 18633 2785
rect 341 2550 385 2588
rect 341 2530 353 2550
rect 373 2530 385 2550
rect 341 2488 385 2530
rect 435 2550 477 2588
rect 435 2530 449 2550
rect 469 2530 477 2550
rect 435 2488 477 2530
rect 554 2550 598 2588
rect 554 2530 566 2550
rect 586 2530 598 2550
rect 554 2488 598 2530
rect 648 2550 690 2588
rect 648 2530 662 2550
rect 682 2530 690 2550
rect 648 2488 690 2530
rect 762 2550 806 2588
rect 762 2530 774 2550
rect 794 2530 806 2550
rect 762 2488 806 2530
rect 856 2550 898 2588
rect 856 2530 870 2550
rect 890 2530 898 2550
rect 856 2488 898 2530
rect 972 2550 1014 2588
rect 972 2530 980 2550
rect 1000 2530 1014 2550
rect 972 2488 1014 2530
rect 1064 2557 1109 2588
rect 1064 2550 1108 2557
rect 1064 2530 1076 2550
rect 1096 2530 1108 2550
rect 5397 2591 5441 2629
rect 5397 2571 5409 2591
rect 5429 2571 5441 2591
rect 1064 2488 1108 2530
rect 3828 2490 3872 2532
rect 3828 2470 3840 2490
rect 3860 2470 3872 2490
rect 3828 2463 3872 2470
rect 3827 2432 3872 2463
rect 3922 2490 3964 2532
rect 3922 2470 3936 2490
rect 3956 2470 3964 2490
rect 3922 2432 3964 2470
rect 4038 2490 4080 2532
rect 4038 2470 4046 2490
rect 4066 2470 4080 2490
rect 4038 2432 4080 2470
rect 4130 2490 4174 2532
rect 4130 2470 4142 2490
rect 4162 2470 4174 2490
rect 4130 2432 4174 2470
rect 4246 2490 4288 2532
rect 4246 2470 4254 2490
rect 4274 2470 4288 2490
rect 4246 2432 4288 2470
rect 4338 2490 4382 2532
rect 4338 2470 4350 2490
rect 4370 2470 4382 2490
rect 4338 2432 4382 2470
rect 4459 2490 4501 2532
rect 4459 2470 4467 2490
rect 4487 2470 4501 2490
rect 4459 2432 4501 2470
rect 4551 2490 4595 2532
rect 5397 2529 5441 2571
rect 5491 2591 5533 2629
rect 5491 2571 5505 2591
rect 5525 2571 5533 2591
rect 5491 2529 5533 2571
rect 5610 2591 5654 2629
rect 5610 2571 5622 2591
rect 5642 2571 5654 2591
rect 5610 2529 5654 2571
rect 5704 2591 5746 2629
rect 5704 2571 5718 2591
rect 5738 2571 5746 2591
rect 5704 2529 5746 2571
rect 5818 2591 5862 2629
rect 5818 2571 5830 2591
rect 5850 2571 5862 2591
rect 5818 2529 5862 2571
rect 5912 2591 5954 2629
rect 5912 2571 5926 2591
rect 5946 2571 5954 2591
rect 5912 2529 5954 2571
rect 6028 2591 6070 2629
rect 6028 2571 6036 2591
rect 6056 2571 6070 2591
rect 6028 2529 6070 2571
rect 6120 2598 6165 2629
rect 6120 2591 6164 2598
rect 6120 2571 6132 2591
rect 6152 2571 6164 2591
rect 6120 2529 6164 2571
rect 8884 2531 8928 2573
rect 4551 2470 4563 2490
rect 4583 2470 4595 2490
rect 4551 2432 4595 2470
rect 8884 2511 8896 2531
rect 8916 2511 8928 2531
rect 8884 2504 8928 2511
rect 8883 2473 8928 2504
rect 8978 2531 9020 2573
rect 8978 2511 8992 2531
rect 9012 2511 9020 2531
rect 8978 2473 9020 2511
rect 9094 2531 9136 2573
rect 9094 2511 9102 2531
rect 9122 2511 9136 2531
rect 9094 2473 9136 2511
rect 9186 2531 9230 2573
rect 9186 2511 9198 2531
rect 9218 2511 9230 2531
rect 9186 2473 9230 2511
rect 9302 2531 9344 2573
rect 9302 2511 9310 2531
rect 9330 2511 9344 2531
rect 9302 2473 9344 2511
rect 9394 2531 9438 2573
rect 9394 2511 9406 2531
rect 9426 2511 9438 2531
rect 9394 2473 9438 2511
rect 9515 2531 9557 2573
rect 9515 2511 9523 2531
rect 9543 2511 9557 2531
rect 9515 2473 9557 2511
rect 9607 2531 9651 2573
rect 10372 2555 10416 2593
rect 9607 2511 9619 2531
rect 9639 2511 9651 2531
rect 9607 2473 9651 2511
rect 10372 2535 10384 2555
rect 10404 2535 10416 2555
rect 10372 2493 10416 2535
rect 10466 2555 10508 2593
rect 10466 2535 10480 2555
rect 10500 2535 10508 2555
rect 10466 2493 10508 2535
rect 10585 2555 10629 2593
rect 10585 2535 10597 2555
rect 10617 2535 10629 2555
rect 10585 2493 10629 2535
rect 10679 2555 10721 2593
rect 10679 2535 10693 2555
rect 10713 2535 10721 2555
rect 10679 2493 10721 2535
rect 10793 2555 10837 2593
rect 10793 2535 10805 2555
rect 10825 2535 10837 2555
rect 10793 2493 10837 2535
rect 10887 2555 10929 2593
rect 10887 2535 10901 2555
rect 10921 2535 10929 2555
rect 10887 2493 10929 2535
rect 11003 2555 11045 2593
rect 11003 2535 11011 2555
rect 11031 2535 11045 2555
rect 11003 2493 11045 2535
rect 11095 2562 11140 2593
rect 11095 2555 11139 2562
rect 11095 2535 11107 2555
rect 11127 2535 11139 2555
rect 15428 2596 15472 2634
rect 15428 2576 15440 2596
rect 15460 2576 15472 2596
rect 11095 2493 11139 2535
rect 13859 2495 13903 2537
rect 1279 2306 1323 2344
rect 1279 2286 1291 2306
rect 1311 2286 1323 2306
rect 1279 2244 1323 2286
rect 1373 2306 1415 2344
rect 1373 2286 1387 2306
rect 1407 2286 1415 2306
rect 1373 2244 1415 2286
rect 1492 2306 1536 2344
rect 1492 2286 1504 2306
rect 1524 2286 1536 2306
rect 1492 2244 1536 2286
rect 1586 2306 1628 2344
rect 1586 2286 1600 2306
rect 1620 2286 1628 2306
rect 1586 2244 1628 2286
rect 1700 2306 1744 2344
rect 1700 2286 1712 2306
rect 1732 2286 1744 2306
rect 1700 2244 1744 2286
rect 1794 2306 1836 2344
rect 1794 2286 1808 2306
rect 1828 2286 1836 2306
rect 1794 2244 1836 2286
rect 1910 2306 1952 2344
rect 1910 2286 1918 2306
rect 1938 2286 1952 2306
rect 1910 2244 1952 2286
rect 2002 2313 2047 2344
rect 2002 2306 2046 2313
rect 2002 2286 2014 2306
rect 2034 2286 2046 2306
rect 2002 2244 2046 2286
rect 6335 2347 6379 2385
rect 6335 2327 6347 2347
rect 6367 2327 6379 2347
rect 2889 2180 2933 2222
rect 2889 2160 2901 2180
rect 2921 2160 2933 2180
rect 2889 2153 2933 2160
rect 2888 2122 2933 2153
rect 2983 2180 3025 2222
rect 2983 2160 2997 2180
rect 3017 2160 3025 2180
rect 2983 2122 3025 2160
rect 3099 2180 3141 2222
rect 3099 2160 3107 2180
rect 3127 2160 3141 2180
rect 3099 2122 3141 2160
rect 3191 2180 3235 2222
rect 3191 2160 3203 2180
rect 3223 2160 3235 2180
rect 3191 2122 3235 2160
rect 3307 2180 3349 2222
rect 3307 2160 3315 2180
rect 3335 2160 3349 2180
rect 3307 2122 3349 2160
rect 3399 2180 3443 2222
rect 3399 2160 3411 2180
rect 3431 2160 3443 2180
rect 3399 2122 3443 2160
rect 3520 2180 3562 2222
rect 3520 2160 3528 2180
rect 3548 2160 3562 2180
rect 3520 2122 3562 2160
rect 3612 2180 3656 2222
rect 6335 2285 6379 2327
rect 6429 2347 6471 2385
rect 6429 2327 6443 2347
rect 6463 2327 6471 2347
rect 6429 2285 6471 2327
rect 6548 2347 6592 2385
rect 6548 2327 6560 2347
rect 6580 2327 6592 2347
rect 6548 2285 6592 2327
rect 6642 2347 6684 2385
rect 6642 2327 6656 2347
rect 6676 2327 6684 2347
rect 6642 2285 6684 2327
rect 6756 2347 6800 2385
rect 6756 2327 6768 2347
rect 6788 2327 6800 2347
rect 6756 2285 6800 2327
rect 6850 2347 6892 2385
rect 6850 2327 6864 2347
rect 6884 2327 6892 2347
rect 6850 2285 6892 2327
rect 6966 2347 7008 2385
rect 6966 2327 6974 2347
rect 6994 2327 7008 2347
rect 6966 2285 7008 2327
rect 7058 2354 7103 2385
rect 13859 2475 13871 2495
rect 13891 2475 13903 2495
rect 13859 2468 13903 2475
rect 7058 2347 7102 2354
rect 7058 2327 7070 2347
rect 7090 2327 7102 2347
rect 13858 2437 13903 2468
rect 13953 2495 13995 2537
rect 13953 2475 13967 2495
rect 13987 2475 13995 2495
rect 13953 2437 13995 2475
rect 14069 2495 14111 2537
rect 14069 2475 14077 2495
rect 14097 2475 14111 2495
rect 14069 2437 14111 2475
rect 14161 2495 14205 2537
rect 14161 2475 14173 2495
rect 14193 2475 14205 2495
rect 14161 2437 14205 2475
rect 14277 2495 14319 2537
rect 14277 2475 14285 2495
rect 14305 2475 14319 2495
rect 14277 2437 14319 2475
rect 14369 2495 14413 2537
rect 14369 2475 14381 2495
rect 14401 2475 14413 2495
rect 14369 2437 14413 2475
rect 14490 2495 14532 2537
rect 14490 2475 14498 2495
rect 14518 2475 14532 2495
rect 14490 2437 14532 2475
rect 14582 2495 14626 2537
rect 15428 2534 15472 2576
rect 15522 2596 15564 2634
rect 15522 2576 15536 2596
rect 15556 2576 15564 2596
rect 15522 2534 15564 2576
rect 15641 2596 15685 2634
rect 15641 2576 15653 2596
rect 15673 2576 15685 2596
rect 15641 2534 15685 2576
rect 15735 2596 15777 2634
rect 15735 2576 15749 2596
rect 15769 2576 15777 2596
rect 15735 2534 15777 2576
rect 15849 2596 15893 2634
rect 15849 2576 15861 2596
rect 15881 2576 15893 2596
rect 15849 2534 15893 2576
rect 15943 2596 15985 2634
rect 15943 2576 15957 2596
rect 15977 2576 15985 2596
rect 15943 2534 15985 2576
rect 16059 2596 16101 2634
rect 16059 2576 16067 2596
rect 16087 2576 16101 2596
rect 16059 2534 16101 2576
rect 16151 2603 16196 2634
rect 16151 2596 16195 2603
rect 16151 2576 16163 2596
rect 16183 2576 16195 2596
rect 16151 2534 16195 2576
rect 18915 2536 18959 2578
rect 14582 2475 14594 2495
rect 14614 2475 14626 2495
rect 14582 2437 14626 2475
rect 18915 2516 18927 2536
rect 18947 2516 18959 2536
rect 18915 2509 18959 2516
rect 18914 2478 18959 2509
rect 19009 2536 19051 2578
rect 19009 2516 19023 2536
rect 19043 2516 19051 2536
rect 19009 2478 19051 2516
rect 19125 2536 19167 2578
rect 19125 2516 19133 2536
rect 19153 2516 19167 2536
rect 19125 2478 19167 2516
rect 19217 2536 19261 2578
rect 19217 2516 19229 2536
rect 19249 2516 19261 2536
rect 19217 2478 19261 2516
rect 19333 2536 19375 2578
rect 19333 2516 19341 2536
rect 19361 2516 19375 2536
rect 19333 2478 19375 2516
rect 19425 2536 19469 2578
rect 19425 2516 19437 2536
rect 19457 2516 19469 2536
rect 19425 2478 19469 2516
rect 19546 2536 19588 2578
rect 19546 2516 19554 2536
rect 19574 2516 19588 2536
rect 19546 2478 19588 2516
rect 19638 2536 19682 2578
rect 19638 2516 19650 2536
rect 19670 2516 19682 2536
rect 19638 2478 19682 2516
rect 7058 2285 7102 2327
rect 3612 2160 3624 2180
rect 3644 2160 3656 2180
rect 3612 2122 3656 2160
rect 7945 2221 7989 2263
rect 7945 2201 7957 2221
rect 7977 2201 7989 2221
rect 7945 2194 7989 2201
rect 7944 2163 7989 2194
rect 8039 2221 8081 2263
rect 8039 2201 8053 2221
rect 8073 2201 8081 2221
rect 8039 2163 8081 2201
rect 8155 2221 8197 2263
rect 8155 2201 8163 2221
rect 8183 2201 8197 2221
rect 8155 2163 8197 2201
rect 8247 2221 8291 2263
rect 8247 2201 8259 2221
rect 8279 2201 8291 2221
rect 8247 2163 8291 2201
rect 8363 2221 8405 2263
rect 8363 2201 8371 2221
rect 8391 2201 8405 2221
rect 8363 2163 8405 2201
rect 8455 2221 8499 2263
rect 8455 2201 8467 2221
rect 8487 2201 8499 2221
rect 8455 2163 8499 2201
rect 8576 2221 8618 2263
rect 8576 2201 8584 2221
rect 8604 2201 8618 2221
rect 8576 2163 8618 2201
rect 8668 2221 8712 2263
rect 11310 2311 11354 2349
rect 11310 2291 11322 2311
rect 11342 2291 11354 2311
rect 8668 2201 8680 2221
rect 8700 2201 8712 2221
rect 8668 2163 8712 2201
rect 11310 2249 11354 2291
rect 11404 2311 11446 2349
rect 11404 2291 11418 2311
rect 11438 2291 11446 2311
rect 11404 2249 11446 2291
rect 11523 2311 11567 2349
rect 11523 2291 11535 2311
rect 11555 2291 11567 2311
rect 11523 2249 11567 2291
rect 11617 2311 11659 2349
rect 11617 2291 11631 2311
rect 11651 2291 11659 2311
rect 11617 2249 11659 2291
rect 11731 2311 11775 2349
rect 11731 2291 11743 2311
rect 11763 2291 11775 2311
rect 11731 2249 11775 2291
rect 11825 2311 11867 2349
rect 11825 2291 11839 2311
rect 11859 2291 11867 2311
rect 11825 2249 11867 2291
rect 11941 2311 11983 2349
rect 11941 2291 11949 2311
rect 11969 2291 11983 2311
rect 11941 2249 11983 2291
rect 12033 2318 12078 2349
rect 12033 2311 12077 2318
rect 12033 2291 12045 2311
rect 12065 2291 12077 2311
rect 12033 2249 12077 2291
rect 16366 2352 16410 2390
rect 16366 2332 16378 2352
rect 16398 2332 16410 2352
rect 12920 2185 12964 2227
rect 340 1996 384 2034
rect 340 1976 352 1996
rect 372 1976 384 1996
rect 340 1934 384 1976
rect 434 1996 476 2034
rect 434 1976 448 1996
rect 468 1976 476 1996
rect 434 1934 476 1976
rect 553 1996 597 2034
rect 553 1976 565 1996
rect 585 1976 597 1996
rect 553 1934 597 1976
rect 647 1996 689 2034
rect 647 1976 661 1996
rect 681 1976 689 1996
rect 647 1934 689 1976
rect 761 1996 805 2034
rect 761 1976 773 1996
rect 793 1976 805 1996
rect 761 1934 805 1976
rect 855 1996 897 2034
rect 855 1976 869 1996
rect 889 1976 897 1996
rect 855 1934 897 1976
rect 971 1996 1013 2034
rect 971 1976 979 1996
rect 999 1976 1013 1996
rect 971 1934 1013 1976
rect 1063 2003 1108 2034
rect 1063 1996 1107 2003
rect 1063 1976 1075 1996
rect 1095 1976 1107 1996
rect 5396 2037 5440 2075
rect 5396 2017 5408 2037
rect 5428 2017 5440 2037
rect 1063 1934 1107 1976
rect 3827 1936 3871 1978
rect 3827 1916 3839 1936
rect 3859 1916 3871 1936
rect 3827 1909 3871 1916
rect 3826 1878 3871 1909
rect 3921 1936 3963 1978
rect 3921 1916 3935 1936
rect 3955 1916 3963 1936
rect 3921 1878 3963 1916
rect 4037 1936 4079 1978
rect 4037 1916 4045 1936
rect 4065 1916 4079 1936
rect 4037 1878 4079 1916
rect 4129 1936 4173 1978
rect 4129 1916 4141 1936
rect 4161 1916 4173 1936
rect 4129 1878 4173 1916
rect 4245 1936 4287 1978
rect 4245 1916 4253 1936
rect 4273 1916 4287 1936
rect 4245 1878 4287 1916
rect 4337 1936 4381 1978
rect 4337 1916 4349 1936
rect 4369 1916 4381 1936
rect 4337 1878 4381 1916
rect 4458 1936 4500 1978
rect 4458 1916 4466 1936
rect 4486 1916 4500 1936
rect 4458 1878 4500 1916
rect 4550 1936 4594 1978
rect 5396 1975 5440 2017
rect 5490 2037 5532 2075
rect 5490 2017 5504 2037
rect 5524 2017 5532 2037
rect 5490 1975 5532 2017
rect 5609 2037 5653 2075
rect 5609 2017 5621 2037
rect 5641 2017 5653 2037
rect 5609 1975 5653 2017
rect 5703 2037 5745 2075
rect 5703 2017 5717 2037
rect 5737 2017 5745 2037
rect 5703 1975 5745 2017
rect 5817 2037 5861 2075
rect 5817 2017 5829 2037
rect 5849 2017 5861 2037
rect 5817 1975 5861 2017
rect 5911 2037 5953 2075
rect 5911 2017 5925 2037
rect 5945 2017 5953 2037
rect 5911 1975 5953 2017
rect 6027 2037 6069 2075
rect 6027 2017 6035 2037
rect 6055 2017 6069 2037
rect 6027 1975 6069 2017
rect 6119 2044 6164 2075
rect 12920 2165 12932 2185
rect 12952 2165 12964 2185
rect 12920 2158 12964 2165
rect 6119 2037 6163 2044
rect 6119 2017 6131 2037
rect 6151 2017 6163 2037
rect 12919 2127 12964 2158
rect 13014 2185 13056 2227
rect 13014 2165 13028 2185
rect 13048 2165 13056 2185
rect 13014 2127 13056 2165
rect 13130 2185 13172 2227
rect 13130 2165 13138 2185
rect 13158 2165 13172 2185
rect 13130 2127 13172 2165
rect 13222 2185 13266 2227
rect 13222 2165 13234 2185
rect 13254 2165 13266 2185
rect 13222 2127 13266 2165
rect 13338 2185 13380 2227
rect 13338 2165 13346 2185
rect 13366 2165 13380 2185
rect 13338 2127 13380 2165
rect 13430 2185 13474 2227
rect 13430 2165 13442 2185
rect 13462 2165 13474 2185
rect 13430 2127 13474 2165
rect 13551 2185 13593 2227
rect 13551 2165 13559 2185
rect 13579 2165 13593 2185
rect 13551 2127 13593 2165
rect 13643 2185 13687 2227
rect 16366 2290 16410 2332
rect 16460 2352 16502 2390
rect 16460 2332 16474 2352
rect 16494 2332 16502 2352
rect 16460 2290 16502 2332
rect 16579 2352 16623 2390
rect 16579 2332 16591 2352
rect 16611 2332 16623 2352
rect 16579 2290 16623 2332
rect 16673 2352 16715 2390
rect 16673 2332 16687 2352
rect 16707 2332 16715 2352
rect 16673 2290 16715 2332
rect 16787 2352 16831 2390
rect 16787 2332 16799 2352
rect 16819 2332 16831 2352
rect 16787 2290 16831 2332
rect 16881 2352 16923 2390
rect 16881 2332 16895 2352
rect 16915 2332 16923 2352
rect 16881 2290 16923 2332
rect 16997 2352 17039 2390
rect 16997 2332 17005 2352
rect 17025 2332 17039 2352
rect 16997 2290 17039 2332
rect 17089 2359 17134 2390
rect 17089 2352 17133 2359
rect 17089 2332 17101 2352
rect 17121 2332 17133 2352
rect 17089 2290 17133 2332
rect 13643 2165 13655 2185
rect 13675 2165 13687 2185
rect 13643 2127 13687 2165
rect 17976 2226 18020 2268
rect 17976 2206 17988 2226
rect 18008 2206 18020 2226
rect 17976 2199 18020 2206
rect 17975 2168 18020 2199
rect 18070 2226 18112 2268
rect 18070 2206 18084 2226
rect 18104 2206 18112 2226
rect 18070 2168 18112 2206
rect 18186 2226 18228 2268
rect 18186 2206 18194 2226
rect 18214 2206 18228 2226
rect 18186 2168 18228 2206
rect 18278 2226 18322 2268
rect 18278 2206 18290 2226
rect 18310 2206 18322 2226
rect 18278 2168 18322 2206
rect 18394 2226 18436 2268
rect 18394 2206 18402 2226
rect 18422 2206 18436 2226
rect 18394 2168 18436 2206
rect 18486 2226 18530 2268
rect 18486 2206 18498 2226
rect 18518 2206 18530 2226
rect 18486 2168 18530 2206
rect 18607 2226 18649 2268
rect 18607 2206 18615 2226
rect 18635 2206 18649 2226
rect 18607 2168 18649 2206
rect 18699 2226 18743 2268
rect 18699 2206 18711 2226
rect 18731 2206 18743 2226
rect 18699 2168 18743 2206
rect 6119 1975 6163 2017
rect 8883 1977 8927 2019
rect 4550 1916 4562 1936
rect 4582 1916 4594 1936
rect 4550 1878 4594 1916
rect 8883 1957 8895 1977
rect 8915 1957 8927 1977
rect 8883 1950 8927 1957
rect 8882 1919 8927 1950
rect 8977 1977 9019 2019
rect 8977 1957 8991 1977
rect 9011 1957 9019 1977
rect 8977 1919 9019 1957
rect 9093 1977 9135 2019
rect 9093 1957 9101 1977
rect 9121 1957 9135 1977
rect 9093 1919 9135 1957
rect 9185 1977 9229 2019
rect 9185 1957 9197 1977
rect 9217 1957 9229 1977
rect 9185 1919 9229 1957
rect 9301 1977 9343 2019
rect 9301 1957 9309 1977
rect 9329 1957 9343 1977
rect 9301 1919 9343 1957
rect 9393 1977 9437 2019
rect 9393 1957 9405 1977
rect 9425 1957 9437 1977
rect 9393 1919 9437 1957
rect 9514 1977 9556 2019
rect 9514 1957 9522 1977
rect 9542 1957 9556 1977
rect 9514 1919 9556 1957
rect 9606 1977 9650 2019
rect 9606 1957 9618 1977
rect 9638 1957 9650 1977
rect 10371 2001 10415 2039
rect 10371 1981 10383 2001
rect 10403 1981 10415 2001
rect 9606 1919 9650 1957
rect 10371 1939 10415 1981
rect 10465 2001 10507 2039
rect 10465 1981 10479 2001
rect 10499 1981 10507 2001
rect 10465 1939 10507 1981
rect 10584 2001 10628 2039
rect 10584 1981 10596 2001
rect 10616 1981 10628 2001
rect 10584 1939 10628 1981
rect 10678 2001 10720 2039
rect 10678 1981 10692 2001
rect 10712 1981 10720 2001
rect 10678 1939 10720 1981
rect 10792 2001 10836 2039
rect 10792 1981 10804 2001
rect 10824 1981 10836 2001
rect 10792 1939 10836 1981
rect 10886 2001 10928 2039
rect 10886 1981 10900 2001
rect 10920 1981 10928 2001
rect 10886 1939 10928 1981
rect 11002 2001 11044 2039
rect 11002 1981 11010 2001
rect 11030 1981 11044 2001
rect 11002 1939 11044 1981
rect 11094 2008 11139 2039
rect 11094 2001 11138 2008
rect 11094 1981 11106 2001
rect 11126 1981 11138 2001
rect 15427 2042 15471 2080
rect 15427 2022 15439 2042
rect 15459 2022 15471 2042
rect 11094 1939 11138 1981
rect 13858 1941 13902 1983
rect 13858 1921 13870 1941
rect 13890 1921 13902 1941
rect 13858 1914 13902 1921
rect 13857 1883 13902 1914
rect 13952 1941 13994 1983
rect 13952 1921 13966 1941
rect 13986 1921 13994 1941
rect 13952 1883 13994 1921
rect 14068 1941 14110 1983
rect 14068 1921 14076 1941
rect 14096 1921 14110 1941
rect 14068 1883 14110 1921
rect 14160 1941 14204 1983
rect 14160 1921 14172 1941
rect 14192 1921 14204 1941
rect 14160 1883 14204 1921
rect 14276 1941 14318 1983
rect 14276 1921 14284 1941
rect 14304 1921 14318 1941
rect 14276 1883 14318 1921
rect 14368 1941 14412 1983
rect 14368 1921 14380 1941
rect 14400 1921 14412 1941
rect 14368 1883 14412 1921
rect 14489 1941 14531 1983
rect 14489 1921 14497 1941
rect 14517 1921 14531 1941
rect 14489 1883 14531 1921
rect 14581 1941 14625 1983
rect 15427 1980 15471 2022
rect 15521 2042 15563 2080
rect 15521 2022 15535 2042
rect 15555 2022 15563 2042
rect 15521 1980 15563 2022
rect 15640 2042 15684 2080
rect 15640 2022 15652 2042
rect 15672 2022 15684 2042
rect 15640 1980 15684 2022
rect 15734 2042 15776 2080
rect 15734 2022 15748 2042
rect 15768 2022 15776 2042
rect 15734 1980 15776 2022
rect 15848 2042 15892 2080
rect 15848 2022 15860 2042
rect 15880 2022 15892 2042
rect 15848 1980 15892 2022
rect 15942 2042 15984 2080
rect 15942 2022 15956 2042
rect 15976 2022 15984 2042
rect 15942 1980 15984 2022
rect 16058 2042 16100 2080
rect 16058 2022 16066 2042
rect 16086 2022 16100 2042
rect 16058 1980 16100 2022
rect 16150 2049 16195 2080
rect 16150 2042 16194 2049
rect 16150 2022 16162 2042
rect 16182 2022 16194 2042
rect 16150 1980 16194 2022
rect 18914 1982 18958 2024
rect 14581 1921 14593 1941
rect 14613 1921 14625 1941
rect 14581 1883 14625 1921
rect 18914 1962 18926 1982
rect 18946 1962 18958 1982
rect 18914 1955 18958 1962
rect 18913 1924 18958 1955
rect 19008 1982 19050 2024
rect 19008 1962 19022 1982
rect 19042 1962 19050 1982
rect 19008 1924 19050 1962
rect 19124 1982 19166 2024
rect 19124 1962 19132 1982
rect 19152 1962 19166 1982
rect 19124 1924 19166 1962
rect 19216 1982 19260 2024
rect 19216 1962 19228 1982
rect 19248 1962 19260 1982
rect 19216 1924 19260 1962
rect 19332 1982 19374 2024
rect 19332 1962 19340 1982
rect 19360 1962 19374 1982
rect 19332 1924 19374 1962
rect 19424 1982 19468 2024
rect 19424 1962 19436 1982
rect 19456 1962 19468 1982
rect 19424 1924 19468 1962
rect 19545 1982 19587 2024
rect 19545 1962 19553 1982
rect 19573 1962 19587 1982
rect 19545 1924 19587 1962
rect 19637 1982 19681 2024
rect 19637 1962 19649 1982
rect 19669 1962 19681 1982
rect 19637 1924 19681 1962
rect 1420 1714 1464 1752
rect 1420 1694 1432 1714
rect 1452 1694 1464 1714
rect 1420 1652 1464 1694
rect 1514 1714 1556 1752
rect 1514 1694 1528 1714
rect 1548 1694 1556 1714
rect 1514 1652 1556 1694
rect 1633 1714 1677 1752
rect 1633 1694 1645 1714
rect 1665 1694 1677 1714
rect 1633 1652 1677 1694
rect 1727 1714 1769 1752
rect 1727 1694 1741 1714
rect 1761 1694 1769 1714
rect 1727 1652 1769 1694
rect 1841 1714 1885 1752
rect 1841 1694 1853 1714
rect 1873 1694 1885 1714
rect 1841 1652 1885 1694
rect 1935 1714 1977 1752
rect 1935 1694 1949 1714
rect 1969 1694 1977 1714
rect 1935 1652 1977 1694
rect 2051 1714 2093 1752
rect 2051 1694 2059 1714
rect 2079 1694 2093 1714
rect 2051 1652 2093 1694
rect 2143 1721 2188 1752
rect 2143 1714 2187 1721
rect 2143 1694 2155 1714
rect 2175 1694 2187 1714
rect 6476 1755 6520 1793
rect 6476 1735 6488 1755
rect 6508 1735 6520 1755
rect 2143 1652 2187 1694
rect 2749 1669 2793 1711
rect 2749 1649 2761 1669
rect 2781 1649 2793 1669
rect 2749 1642 2793 1649
rect 2748 1611 2793 1642
rect 2843 1669 2885 1711
rect 2843 1649 2857 1669
rect 2877 1649 2885 1669
rect 2843 1611 2885 1649
rect 2959 1669 3001 1711
rect 2959 1649 2967 1669
rect 2987 1649 3001 1669
rect 2959 1611 3001 1649
rect 3051 1669 3095 1711
rect 3051 1649 3063 1669
rect 3083 1649 3095 1669
rect 3051 1611 3095 1649
rect 3167 1669 3209 1711
rect 3167 1649 3175 1669
rect 3195 1649 3209 1669
rect 3167 1611 3209 1649
rect 3259 1669 3303 1711
rect 3259 1649 3271 1669
rect 3291 1649 3303 1669
rect 3259 1611 3303 1649
rect 3380 1669 3422 1711
rect 3380 1649 3388 1669
rect 3408 1649 3422 1669
rect 3380 1611 3422 1649
rect 3472 1669 3516 1711
rect 6476 1693 6520 1735
rect 6570 1755 6612 1793
rect 6570 1735 6584 1755
rect 6604 1735 6612 1755
rect 6570 1693 6612 1735
rect 6689 1755 6733 1793
rect 6689 1735 6701 1755
rect 6721 1735 6733 1755
rect 6689 1693 6733 1735
rect 6783 1755 6825 1793
rect 6783 1735 6797 1755
rect 6817 1735 6825 1755
rect 6783 1693 6825 1735
rect 6897 1755 6941 1793
rect 6897 1735 6909 1755
rect 6929 1735 6941 1755
rect 6897 1693 6941 1735
rect 6991 1755 7033 1793
rect 6991 1735 7005 1755
rect 7025 1735 7033 1755
rect 6991 1693 7033 1735
rect 7107 1755 7149 1793
rect 7107 1735 7115 1755
rect 7135 1735 7149 1755
rect 7107 1693 7149 1735
rect 7199 1762 7244 1793
rect 7199 1755 7243 1762
rect 7199 1735 7211 1755
rect 7231 1735 7243 1755
rect 7199 1693 7243 1735
rect 7805 1710 7849 1752
rect 3472 1649 3484 1669
rect 3504 1649 3516 1669
rect 3472 1611 3516 1649
rect 7805 1690 7817 1710
rect 7837 1690 7849 1710
rect 7805 1683 7849 1690
rect 7804 1652 7849 1683
rect 7899 1710 7941 1752
rect 7899 1690 7913 1710
rect 7933 1690 7941 1710
rect 7899 1652 7941 1690
rect 8015 1710 8057 1752
rect 8015 1690 8023 1710
rect 8043 1690 8057 1710
rect 8015 1652 8057 1690
rect 8107 1710 8151 1752
rect 8107 1690 8119 1710
rect 8139 1690 8151 1710
rect 8107 1652 8151 1690
rect 8223 1710 8265 1752
rect 8223 1690 8231 1710
rect 8251 1690 8265 1710
rect 8223 1652 8265 1690
rect 8315 1710 8359 1752
rect 8315 1690 8327 1710
rect 8347 1690 8359 1710
rect 8315 1652 8359 1690
rect 8436 1710 8478 1752
rect 8436 1690 8444 1710
rect 8464 1690 8478 1710
rect 8436 1652 8478 1690
rect 8528 1710 8572 1752
rect 8528 1690 8540 1710
rect 8560 1690 8572 1710
rect 8528 1652 8572 1690
rect 11451 1719 11495 1757
rect 11451 1699 11463 1719
rect 11483 1699 11495 1719
rect 11451 1657 11495 1699
rect 11545 1719 11587 1757
rect 11545 1699 11559 1719
rect 11579 1699 11587 1719
rect 11545 1657 11587 1699
rect 11664 1719 11708 1757
rect 11664 1699 11676 1719
rect 11696 1699 11708 1719
rect 11664 1657 11708 1699
rect 11758 1719 11800 1757
rect 11758 1699 11772 1719
rect 11792 1699 11800 1719
rect 11758 1657 11800 1699
rect 11872 1719 11916 1757
rect 11872 1699 11884 1719
rect 11904 1699 11916 1719
rect 11872 1657 11916 1699
rect 11966 1719 12008 1757
rect 11966 1699 11980 1719
rect 12000 1699 12008 1719
rect 11966 1657 12008 1699
rect 12082 1719 12124 1757
rect 12082 1699 12090 1719
rect 12110 1699 12124 1719
rect 12082 1657 12124 1699
rect 12174 1726 12219 1757
rect 12174 1719 12218 1726
rect 12174 1699 12186 1719
rect 12206 1699 12218 1719
rect 16507 1760 16551 1798
rect 16507 1740 16519 1760
rect 16539 1740 16551 1760
rect 12174 1657 12218 1699
rect 12780 1674 12824 1716
rect 12780 1654 12792 1674
rect 12812 1654 12824 1674
rect 12780 1647 12824 1654
rect 12779 1616 12824 1647
rect 12874 1674 12916 1716
rect 12874 1654 12888 1674
rect 12908 1654 12916 1674
rect 12874 1616 12916 1654
rect 12990 1674 13032 1716
rect 12990 1654 12998 1674
rect 13018 1654 13032 1674
rect 12990 1616 13032 1654
rect 13082 1674 13126 1716
rect 13082 1654 13094 1674
rect 13114 1654 13126 1674
rect 13082 1616 13126 1654
rect 13198 1674 13240 1716
rect 13198 1654 13206 1674
rect 13226 1654 13240 1674
rect 13198 1616 13240 1654
rect 13290 1674 13334 1716
rect 13290 1654 13302 1674
rect 13322 1654 13334 1674
rect 13290 1616 13334 1654
rect 13411 1674 13453 1716
rect 13411 1654 13419 1674
rect 13439 1654 13453 1674
rect 13411 1616 13453 1654
rect 13503 1674 13547 1716
rect 16507 1698 16551 1740
rect 16601 1760 16643 1798
rect 16601 1740 16615 1760
rect 16635 1740 16643 1760
rect 16601 1698 16643 1740
rect 16720 1760 16764 1798
rect 16720 1740 16732 1760
rect 16752 1740 16764 1760
rect 16720 1698 16764 1740
rect 16814 1760 16856 1798
rect 16814 1740 16828 1760
rect 16848 1740 16856 1760
rect 16814 1698 16856 1740
rect 16928 1760 16972 1798
rect 16928 1740 16940 1760
rect 16960 1740 16972 1760
rect 16928 1698 16972 1740
rect 17022 1760 17064 1798
rect 17022 1740 17036 1760
rect 17056 1740 17064 1760
rect 17022 1698 17064 1740
rect 17138 1760 17180 1798
rect 17138 1740 17146 1760
rect 17166 1740 17180 1760
rect 17138 1698 17180 1740
rect 17230 1767 17275 1798
rect 17230 1760 17274 1767
rect 17230 1740 17242 1760
rect 17262 1740 17274 1760
rect 17230 1698 17274 1740
rect 17836 1715 17880 1757
rect 13503 1654 13515 1674
rect 13535 1654 13547 1674
rect 13503 1616 13547 1654
rect 17836 1695 17848 1715
rect 17868 1695 17880 1715
rect 17836 1688 17880 1695
rect 17835 1657 17880 1688
rect 17930 1715 17972 1757
rect 17930 1695 17944 1715
rect 17964 1695 17972 1715
rect 17930 1657 17972 1695
rect 18046 1715 18088 1757
rect 18046 1695 18054 1715
rect 18074 1695 18088 1715
rect 18046 1657 18088 1695
rect 18138 1715 18182 1757
rect 18138 1695 18150 1715
rect 18170 1695 18182 1715
rect 18138 1657 18182 1695
rect 18254 1715 18296 1757
rect 18254 1695 18262 1715
rect 18282 1695 18296 1715
rect 18254 1657 18296 1695
rect 18346 1715 18390 1757
rect 18346 1695 18358 1715
rect 18378 1695 18390 1715
rect 18346 1657 18390 1695
rect 18467 1715 18509 1757
rect 18467 1695 18475 1715
rect 18495 1695 18509 1715
rect 18467 1657 18509 1695
rect 18559 1715 18603 1757
rect 18559 1695 18571 1715
rect 18591 1695 18603 1715
rect 18559 1657 18603 1695
rect 342 1447 386 1485
rect 342 1427 354 1447
rect 374 1427 386 1447
rect 342 1385 386 1427
rect 436 1447 478 1485
rect 436 1427 450 1447
rect 470 1427 478 1447
rect 436 1385 478 1427
rect 555 1447 599 1485
rect 555 1427 567 1447
rect 587 1427 599 1447
rect 555 1385 599 1427
rect 649 1447 691 1485
rect 649 1427 663 1447
rect 683 1427 691 1447
rect 649 1385 691 1427
rect 763 1447 807 1485
rect 763 1427 775 1447
rect 795 1427 807 1447
rect 763 1385 807 1427
rect 857 1447 899 1485
rect 857 1427 871 1447
rect 891 1427 899 1447
rect 857 1385 899 1427
rect 973 1447 1015 1485
rect 973 1427 981 1447
rect 1001 1427 1015 1447
rect 973 1385 1015 1427
rect 1065 1454 1110 1485
rect 1065 1447 1109 1454
rect 1065 1427 1077 1447
rect 1097 1427 1109 1447
rect 5398 1488 5442 1526
rect 5398 1468 5410 1488
rect 5430 1468 5442 1488
rect 1065 1385 1109 1427
rect 3829 1387 3873 1429
rect 3829 1367 3841 1387
rect 3861 1367 3873 1387
rect 3829 1360 3873 1367
rect 3828 1329 3873 1360
rect 3923 1387 3965 1429
rect 3923 1367 3937 1387
rect 3957 1367 3965 1387
rect 3923 1329 3965 1367
rect 4039 1387 4081 1429
rect 4039 1367 4047 1387
rect 4067 1367 4081 1387
rect 4039 1329 4081 1367
rect 4131 1387 4175 1429
rect 4131 1367 4143 1387
rect 4163 1367 4175 1387
rect 4131 1329 4175 1367
rect 4247 1387 4289 1429
rect 4247 1367 4255 1387
rect 4275 1367 4289 1387
rect 4247 1329 4289 1367
rect 4339 1387 4383 1429
rect 4339 1367 4351 1387
rect 4371 1367 4383 1387
rect 4339 1329 4383 1367
rect 4460 1387 4502 1429
rect 4460 1367 4468 1387
rect 4488 1367 4502 1387
rect 4460 1329 4502 1367
rect 4552 1387 4596 1429
rect 5398 1426 5442 1468
rect 5492 1488 5534 1526
rect 5492 1468 5506 1488
rect 5526 1468 5534 1488
rect 5492 1426 5534 1468
rect 5611 1488 5655 1526
rect 5611 1468 5623 1488
rect 5643 1468 5655 1488
rect 5611 1426 5655 1468
rect 5705 1488 5747 1526
rect 5705 1468 5719 1488
rect 5739 1468 5747 1488
rect 5705 1426 5747 1468
rect 5819 1488 5863 1526
rect 5819 1468 5831 1488
rect 5851 1468 5863 1488
rect 5819 1426 5863 1468
rect 5913 1488 5955 1526
rect 5913 1468 5927 1488
rect 5947 1468 5955 1488
rect 5913 1426 5955 1468
rect 6029 1488 6071 1526
rect 6029 1468 6037 1488
rect 6057 1468 6071 1488
rect 6029 1426 6071 1468
rect 6121 1495 6166 1526
rect 6121 1488 6165 1495
rect 6121 1468 6133 1488
rect 6153 1468 6165 1488
rect 6121 1426 6165 1468
rect 8885 1428 8929 1470
rect 4552 1367 4564 1387
rect 4584 1367 4596 1387
rect 4552 1329 4596 1367
rect 8885 1408 8897 1428
rect 8917 1408 8929 1428
rect 8885 1401 8929 1408
rect 8884 1370 8929 1401
rect 8979 1428 9021 1470
rect 8979 1408 8993 1428
rect 9013 1408 9021 1428
rect 8979 1370 9021 1408
rect 9095 1428 9137 1470
rect 9095 1408 9103 1428
rect 9123 1408 9137 1428
rect 9095 1370 9137 1408
rect 9187 1428 9231 1470
rect 9187 1408 9199 1428
rect 9219 1408 9231 1428
rect 9187 1370 9231 1408
rect 9303 1428 9345 1470
rect 9303 1408 9311 1428
rect 9331 1408 9345 1428
rect 9303 1370 9345 1408
rect 9395 1428 9439 1470
rect 9395 1408 9407 1428
rect 9427 1408 9439 1428
rect 9395 1370 9439 1408
rect 9516 1428 9558 1470
rect 9516 1408 9524 1428
rect 9544 1408 9558 1428
rect 9516 1370 9558 1408
rect 9608 1428 9652 1470
rect 10373 1452 10417 1490
rect 9608 1408 9620 1428
rect 9640 1408 9652 1428
rect 9608 1370 9652 1408
rect 10373 1432 10385 1452
rect 10405 1432 10417 1452
rect 10373 1390 10417 1432
rect 10467 1452 10509 1490
rect 10467 1432 10481 1452
rect 10501 1432 10509 1452
rect 10467 1390 10509 1432
rect 10586 1452 10630 1490
rect 10586 1432 10598 1452
rect 10618 1432 10630 1452
rect 10586 1390 10630 1432
rect 10680 1452 10722 1490
rect 10680 1432 10694 1452
rect 10714 1432 10722 1452
rect 10680 1390 10722 1432
rect 10794 1452 10838 1490
rect 10794 1432 10806 1452
rect 10826 1432 10838 1452
rect 10794 1390 10838 1432
rect 10888 1452 10930 1490
rect 10888 1432 10902 1452
rect 10922 1432 10930 1452
rect 10888 1390 10930 1432
rect 11004 1452 11046 1490
rect 11004 1432 11012 1452
rect 11032 1432 11046 1452
rect 11004 1390 11046 1432
rect 11096 1459 11141 1490
rect 11096 1452 11140 1459
rect 11096 1432 11108 1452
rect 11128 1432 11140 1452
rect 15429 1493 15473 1531
rect 15429 1473 15441 1493
rect 15461 1473 15473 1493
rect 11096 1390 11140 1432
rect 13860 1392 13904 1434
rect 1280 1203 1324 1241
rect 1280 1183 1292 1203
rect 1312 1183 1324 1203
rect 1280 1141 1324 1183
rect 1374 1203 1416 1241
rect 1374 1183 1388 1203
rect 1408 1183 1416 1203
rect 1374 1141 1416 1183
rect 1493 1203 1537 1241
rect 1493 1183 1505 1203
rect 1525 1183 1537 1203
rect 1493 1141 1537 1183
rect 1587 1203 1629 1241
rect 1587 1183 1601 1203
rect 1621 1183 1629 1203
rect 1587 1141 1629 1183
rect 1701 1203 1745 1241
rect 1701 1183 1713 1203
rect 1733 1183 1745 1203
rect 1701 1141 1745 1183
rect 1795 1203 1837 1241
rect 1795 1183 1809 1203
rect 1829 1183 1837 1203
rect 1795 1141 1837 1183
rect 1911 1203 1953 1241
rect 1911 1183 1919 1203
rect 1939 1183 1953 1203
rect 1911 1141 1953 1183
rect 2003 1210 2048 1241
rect 2003 1203 2047 1210
rect 2003 1183 2015 1203
rect 2035 1183 2047 1203
rect 2003 1141 2047 1183
rect 6336 1244 6380 1282
rect 6336 1224 6348 1244
rect 6368 1224 6380 1244
rect 2890 1077 2934 1119
rect 2890 1057 2902 1077
rect 2922 1057 2934 1077
rect 2890 1050 2934 1057
rect 2889 1019 2934 1050
rect 2984 1077 3026 1119
rect 2984 1057 2998 1077
rect 3018 1057 3026 1077
rect 2984 1019 3026 1057
rect 3100 1077 3142 1119
rect 3100 1057 3108 1077
rect 3128 1057 3142 1077
rect 3100 1019 3142 1057
rect 3192 1077 3236 1119
rect 3192 1057 3204 1077
rect 3224 1057 3236 1077
rect 3192 1019 3236 1057
rect 3308 1077 3350 1119
rect 3308 1057 3316 1077
rect 3336 1057 3350 1077
rect 3308 1019 3350 1057
rect 3400 1077 3444 1119
rect 3400 1057 3412 1077
rect 3432 1057 3444 1077
rect 3400 1019 3444 1057
rect 3521 1077 3563 1119
rect 3521 1057 3529 1077
rect 3549 1057 3563 1077
rect 3521 1019 3563 1057
rect 3613 1077 3657 1119
rect 6336 1182 6380 1224
rect 6430 1244 6472 1282
rect 6430 1224 6444 1244
rect 6464 1224 6472 1244
rect 6430 1182 6472 1224
rect 6549 1244 6593 1282
rect 6549 1224 6561 1244
rect 6581 1224 6593 1244
rect 6549 1182 6593 1224
rect 6643 1244 6685 1282
rect 6643 1224 6657 1244
rect 6677 1224 6685 1244
rect 6643 1182 6685 1224
rect 6757 1244 6801 1282
rect 6757 1224 6769 1244
rect 6789 1224 6801 1244
rect 6757 1182 6801 1224
rect 6851 1244 6893 1282
rect 6851 1224 6865 1244
rect 6885 1224 6893 1244
rect 6851 1182 6893 1224
rect 6967 1244 7009 1282
rect 6967 1224 6975 1244
rect 6995 1224 7009 1244
rect 6967 1182 7009 1224
rect 7059 1251 7104 1282
rect 13860 1372 13872 1392
rect 13892 1372 13904 1392
rect 13860 1365 13904 1372
rect 7059 1244 7103 1251
rect 7059 1224 7071 1244
rect 7091 1224 7103 1244
rect 13859 1334 13904 1365
rect 13954 1392 13996 1434
rect 13954 1372 13968 1392
rect 13988 1372 13996 1392
rect 13954 1334 13996 1372
rect 14070 1392 14112 1434
rect 14070 1372 14078 1392
rect 14098 1372 14112 1392
rect 14070 1334 14112 1372
rect 14162 1392 14206 1434
rect 14162 1372 14174 1392
rect 14194 1372 14206 1392
rect 14162 1334 14206 1372
rect 14278 1392 14320 1434
rect 14278 1372 14286 1392
rect 14306 1372 14320 1392
rect 14278 1334 14320 1372
rect 14370 1392 14414 1434
rect 14370 1372 14382 1392
rect 14402 1372 14414 1392
rect 14370 1334 14414 1372
rect 14491 1392 14533 1434
rect 14491 1372 14499 1392
rect 14519 1372 14533 1392
rect 14491 1334 14533 1372
rect 14583 1392 14627 1434
rect 15429 1431 15473 1473
rect 15523 1493 15565 1531
rect 15523 1473 15537 1493
rect 15557 1473 15565 1493
rect 15523 1431 15565 1473
rect 15642 1493 15686 1531
rect 15642 1473 15654 1493
rect 15674 1473 15686 1493
rect 15642 1431 15686 1473
rect 15736 1493 15778 1531
rect 15736 1473 15750 1493
rect 15770 1473 15778 1493
rect 15736 1431 15778 1473
rect 15850 1493 15894 1531
rect 15850 1473 15862 1493
rect 15882 1473 15894 1493
rect 15850 1431 15894 1473
rect 15944 1493 15986 1531
rect 15944 1473 15958 1493
rect 15978 1473 15986 1493
rect 15944 1431 15986 1473
rect 16060 1493 16102 1531
rect 16060 1473 16068 1493
rect 16088 1473 16102 1493
rect 16060 1431 16102 1473
rect 16152 1500 16197 1531
rect 16152 1493 16196 1500
rect 16152 1473 16164 1493
rect 16184 1473 16196 1493
rect 16152 1431 16196 1473
rect 18916 1433 18960 1475
rect 14583 1372 14595 1392
rect 14615 1372 14627 1392
rect 14583 1334 14627 1372
rect 18916 1413 18928 1433
rect 18948 1413 18960 1433
rect 18916 1406 18960 1413
rect 18915 1375 18960 1406
rect 19010 1433 19052 1475
rect 19010 1413 19024 1433
rect 19044 1413 19052 1433
rect 19010 1375 19052 1413
rect 19126 1433 19168 1475
rect 19126 1413 19134 1433
rect 19154 1413 19168 1433
rect 19126 1375 19168 1413
rect 19218 1433 19262 1475
rect 19218 1413 19230 1433
rect 19250 1413 19262 1433
rect 19218 1375 19262 1413
rect 19334 1433 19376 1475
rect 19334 1413 19342 1433
rect 19362 1413 19376 1433
rect 19334 1375 19376 1413
rect 19426 1433 19470 1475
rect 19426 1413 19438 1433
rect 19458 1413 19470 1433
rect 19426 1375 19470 1413
rect 19547 1433 19589 1475
rect 19547 1413 19555 1433
rect 19575 1413 19589 1433
rect 19547 1375 19589 1413
rect 19639 1433 19683 1475
rect 19639 1413 19651 1433
rect 19671 1413 19683 1433
rect 19639 1375 19683 1413
rect 7059 1182 7103 1224
rect 3613 1057 3625 1077
rect 3645 1057 3657 1077
rect 3613 1019 3657 1057
rect 7946 1118 7990 1160
rect 7946 1098 7958 1118
rect 7978 1098 7990 1118
rect 7946 1091 7990 1098
rect 7945 1060 7990 1091
rect 8040 1118 8082 1160
rect 8040 1098 8054 1118
rect 8074 1098 8082 1118
rect 8040 1060 8082 1098
rect 8156 1118 8198 1160
rect 8156 1098 8164 1118
rect 8184 1098 8198 1118
rect 8156 1060 8198 1098
rect 8248 1118 8292 1160
rect 8248 1098 8260 1118
rect 8280 1098 8292 1118
rect 8248 1060 8292 1098
rect 8364 1118 8406 1160
rect 8364 1098 8372 1118
rect 8392 1098 8406 1118
rect 8364 1060 8406 1098
rect 8456 1118 8500 1160
rect 8456 1098 8468 1118
rect 8488 1098 8500 1118
rect 8456 1060 8500 1098
rect 8577 1118 8619 1160
rect 8577 1098 8585 1118
rect 8605 1098 8619 1118
rect 8577 1060 8619 1098
rect 8669 1118 8713 1160
rect 11311 1208 11355 1246
rect 11311 1188 11323 1208
rect 11343 1188 11355 1208
rect 8669 1098 8681 1118
rect 8701 1098 8713 1118
rect 8669 1060 8713 1098
rect 11311 1146 11355 1188
rect 11405 1208 11447 1246
rect 11405 1188 11419 1208
rect 11439 1188 11447 1208
rect 11405 1146 11447 1188
rect 11524 1208 11568 1246
rect 11524 1188 11536 1208
rect 11556 1188 11568 1208
rect 11524 1146 11568 1188
rect 11618 1208 11660 1246
rect 11618 1188 11632 1208
rect 11652 1188 11660 1208
rect 11618 1146 11660 1188
rect 11732 1208 11776 1246
rect 11732 1188 11744 1208
rect 11764 1188 11776 1208
rect 11732 1146 11776 1188
rect 11826 1208 11868 1246
rect 11826 1188 11840 1208
rect 11860 1188 11868 1208
rect 11826 1146 11868 1188
rect 11942 1208 11984 1246
rect 11942 1188 11950 1208
rect 11970 1188 11984 1208
rect 11942 1146 11984 1188
rect 12034 1215 12079 1246
rect 12034 1208 12078 1215
rect 12034 1188 12046 1208
rect 12066 1188 12078 1208
rect 12034 1146 12078 1188
rect 16367 1249 16411 1287
rect 16367 1229 16379 1249
rect 16399 1229 16411 1249
rect 12921 1082 12965 1124
rect 341 893 385 931
rect 341 873 353 893
rect 373 873 385 893
rect 341 831 385 873
rect 435 893 477 931
rect 435 873 449 893
rect 469 873 477 893
rect 435 831 477 873
rect 554 893 598 931
rect 554 873 566 893
rect 586 873 598 893
rect 554 831 598 873
rect 648 893 690 931
rect 648 873 662 893
rect 682 873 690 893
rect 648 831 690 873
rect 762 893 806 931
rect 762 873 774 893
rect 794 873 806 893
rect 762 831 806 873
rect 856 893 898 931
rect 856 873 870 893
rect 890 873 898 893
rect 856 831 898 873
rect 972 893 1014 931
rect 972 873 980 893
rect 1000 873 1014 893
rect 972 831 1014 873
rect 1064 900 1109 931
rect 1064 893 1108 900
rect 1064 873 1076 893
rect 1096 873 1108 893
rect 5397 934 5441 972
rect 5397 914 5409 934
rect 5429 914 5441 934
rect 1064 831 1108 873
rect 3828 833 3872 875
rect 3828 813 3840 833
rect 3860 813 3872 833
rect 3828 806 3872 813
rect 3827 775 3872 806
rect 3922 833 3964 875
rect 3922 813 3936 833
rect 3956 813 3964 833
rect 3922 775 3964 813
rect 4038 833 4080 875
rect 4038 813 4046 833
rect 4066 813 4080 833
rect 4038 775 4080 813
rect 4130 833 4174 875
rect 4130 813 4142 833
rect 4162 813 4174 833
rect 4130 775 4174 813
rect 4246 833 4288 875
rect 4246 813 4254 833
rect 4274 813 4288 833
rect 4246 775 4288 813
rect 4338 833 4382 875
rect 4338 813 4350 833
rect 4370 813 4382 833
rect 4338 775 4382 813
rect 4459 833 4501 875
rect 4459 813 4467 833
rect 4487 813 4501 833
rect 4459 775 4501 813
rect 4551 833 4595 875
rect 5397 872 5441 914
rect 5491 934 5533 972
rect 5491 914 5505 934
rect 5525 914 5533 934
rect 5491 872 5533 914
rect 5610 934 5654 972
rect 5610 914 5622 934
rect 5642 914 5654 934
rect 5610 872 5654 914
rect 5704 934 5746 972
rect 5704 914 5718 934
rect 5738 914 5746 934
rect 5704 872 5746 914
rect 5818 934 5862 972
rect 5818 914 5830 934
rect 5850 914 5862 934
rect 5818 872 5862 914
rect 5912 934 5954 972
rect 5912 914 5926 934
rect 5946 914 5954 934
rect 5912 872 5954 914
rect 6028 934 6070 972
rect 6028 914 6036 934
rect 6056 914 6070 934
rect 6028 872 6070 914
rect 6120 941 6165 972
rect 12921 1062 12933 1082
rect 12953 1062 12965 1082
rect 12921 1055 12965 1062
rect 6120 934 6164 941
rect 6120 914 6132 934
rect 6152 914 6164 934
rect 12920 1024 12965 1055
rect 13015 1082 13057 1124
rect 13015 1062 13029 1082
rect 13049 1062 13057 1082
rect 13015 1024 13057 1062
rect 13131 1082 13173 1124
rect 13131 1062 13139 1082
rect 13159 1062 13173 1082
rect 13131 1024 13173 1062
rect 13223 1082 13267 1124
rect 13223 1062 13235 1082
rect 13255 1062 13267 1082
rect 13223 1024 13267 1062
rect 13339 1082 13381 1124
rect 13339 1062 13347 1082
rect 13367 1062 13381 1082
rect 13339 1024 13381 1062
rect 13431 1082 13475 1124
rect 13431 1062 13443 1082
rect 13463 1062 13475 1082
rect 13431 1024 13475 1062
rect 13552 1082 13594 1124
rect 13552 1062 13560 1082
rect 13580 1062 13594 1082
rect 13552 1024 13594 1062
rect 13644 1082 13688 1124
rect 16367 1187 16411 1229
rect 16461 1249 16503 1287
rect 16461 1229 16475 1249
rect 16495 1229 16503 1249
rect 16461 1187 16503 1229
rect 16580 1249 16624 1287
rect 16580 1229 16592 1249
rect 16612 1229 16624 1249
rect 16580 1187 16624 1229
rect 16674 1249 16716 1287
rect 16674 1229 16688 1249
rect 16708 1229 16716 1249
rect 16674 1187 16716 1229
rect 16788 1249 16832 1287
rect 16788 1229 16800 1249
rect 16820 1229 16832 1249
rect 16788 1187 16832 1229
rect 16882 1249 16924 1287
rect 16882 1229 16896 1249
rect 16916 1229 16924 1249
rect 16882 1187 16924 1229
rect 16998 1249 17040 1287
rect 16998 1229 17006 1249
rect 17026 1229 17040 1249
rect 16998 1187 17040 1229
rect 17090 1256 17135 1287
rect 17090 1249 17134 1256
rect 17090 1229 17102 1249
rect 17122 1229 17134 1249
rect 17090 1187 17134 1229
rect 13644 1062 13656 1082
rect 13676 1062 13688 1082
rect 13644 1024 13688 1062
rect 17977 1123 18021 1165
rect 17977 1103 17989 1123
rect 18009 1103 18021 1123
rect 17977 1096 18021 1103
rect 17976 1065 18021 1096
rect 18071 1123 18113 1165
rect 18071 1103 18085 1123
rect 18105 1103 18113 1123
rect 18071 1065 18113 1103
rect 18187 1123 18229 1165
rect 18187 1103 18195 1123
rect 18215 1103 18229 1123
rect 18187 1065 18229 1103
rect 18279 1123 18323 1165
rect 18279 1103 18291 1123
rect 18311 1103 18323 1123
rect 18279 1065 18323 1103
rect 18395 1123 18437 1165
rect 18395 1103 18403 1123
rect 18423 1103 18437 1123
rect 18395 1065 18437 1103
rect 18487 1123 18531 1165
rect 18487 1103 18499 1123
rect 18519 1103 18531 1123
rect 18487 1065 18531 1103
rect 18608 1123 18650 1165
rect 18608 1103 18616 1123
rect 18636 1103 18650 1123
rect 18608 1065 18650 1103
rect 18700 1123 18744 1165
rect 18700 1103 18712 1123
rect 18732 1103 18744 1123
rect 18700 1065 18744 1103
rect 6120 872 6164 914
rect 8884 874 8928 916
rect 4551 813 4563 833
rect 4583 813 4595 833
rect 4551 775 4595 813
rect 8884 854 8896 874
rect 8916 854 8928 874
rect 8884 847 8928 854
rect 8883 816 8928 847
rect 8978 874 9020 916
rect 8978 854 8992 874
rect 9012 854 9020 874
rect 8978 816 9020 854
rect 9094 874 9136 916
rect 9094 854 9102 874
rect 9122 854 9136 874
rect 9094 816 9136 854
rect 9186 874 9230 916
rect 9186 854 9198 874
rect 9218 854 9230 874
rect 9186 816 9230 854
rect 9302 874 9344 916
rect 9302 854 9310 874
rect 9330 854 9344 874
rect 9302 816 9344 854
rect 9394 874 9438 916
rect 9394 854 9406 874
rect 9426 854 9438 874
rect 9394 816 9438 854
rect 9515 874 9557 916
rect 9515 854 9523 874
rect 9543 854 9557 874
rect 9515 816 9557 854
rect 9607 874 9651 916
rect 9607 854 9619 874
rect 9639 854 9651 874
rect 10372 898 10416 936
rect 10372 878 10384 898
rect 10404 878 10416 898
rect 9607 816 9651 854
rect 10372 836 10416 878
rect 10466 898 10508 936
rect 10466 878 10480 898
rect 10500 878 10508 898
rect 10466 836 10508 878
rect 10585 898 10629 936
rect 10585 878 10597 898
rect 10617 878 10629 898
rect 10585 836 10629 878
rect 10679 898 10721 936
rect 10679 878 10693 898
rect 10713 878 10721 898
rect 10679 836 10721 878
rect 10793 898 10837 936
rect 10793 878 10805 898
rect 10825 878 10837 898
rect 10793 836 10837 878
rect 10887 898 10929 936
rect 10887 878 10901 898
rect 10921 878 10929 898
rect 10887 836 10929 878
rect 11003 898 11045 936
rect 11003 878 11011 898
rect 11031 878 11045 898
rect 11003 836 11045 878
rect 11095 905 11140 936
rect 11095 898 11139 905
rect 11095 878 11107 898
rect 11127 878 11139 898
rect 15428 939 15472 977
rect 15428 919 15440 939
rect 15460 919 15472 939
rect 11095 836 11139 878
rect 13859 838 13903 880
rect 13859 818 13871 838
rect 13891 818 13903 838
rect 13859 811 13903 818
rect 13858 780 13903 811
rect 13953 838 13995 880
rect 13953 818 13967 838
rect 13987 818 13995 838
rect 13953 780 13995 818
rect 14069 838 14111 880
rect 14069 818 14077 838
rect 14097 818 14111 838
rect 14069 780 14111 818
rect 14161 838 14205 880
rect 14161 818 14173 838
rect 14193 818 14205 838
rect 14161 780 14205 818
rect 14277 838 14319 880
rect 14277 818 14285 838
rect 14305 818 14319 838
rect 14277 780 14319 818
rect 14369 838 14413 880
rect 14369 818 14381 838
rect 14401 818 14413 838
rect 14369 780 14413 818
rect 14490 838 14532 880
rect 14490 818 14498 838
rect 14518 818 14532 838
rect 14490 780 14532 818
rect 14582 838 14626 880
rect 15428 877 15472 919
rect 15522 939 15564 977
rect 15522 919 15536 939
rect 15556 919 15564 939
rect 15522 877 15564 919
rect 15641 939 15685 977
rect 15641 919 15653 939
rect 15673 919 15685 939
rect 15641 877 15685 919
rect 15735 939 15777 977
rect 15735 919 15749 939
rect 15769 919 15777 939
rect 15735 877 15777 919
rect 15849 939 15893 977
rect 15849 919 15861 939
rect 15881 919 15893 939
rect 15849 877 15893 919
rect 15943 939 15985 977
rect 15943 919 15957 939
rect 15977 919 15985 939
rect 15943 877 15985 919
rect 16059 939 16101 977
rect 16059 919 16067 939
rect 16087 919 16101 939
rect 16059 877 16101 919
rect 16151 946 16196 977
rect 16151 939 16195 946
rect 16151 919 16163 939
rect 16183 919 16195 939
rect 16151 877 16195 919
rect 18915 879 18959 921
rect 14582 818 14594 838
rect 14614 818 14626 838
rect 14582 780 14626 818
rect 18915 859 18927 879
rect 18947 859 18959 879
rect 18915 852 18959 859
rect 18914 821 18959 852
rect 19009 879 19051 921
rect 19009 859 19023 879
rect 19043 859 19051 879
rect 19009 821 19051 859
rect 19125 879 19167 921
rect 19125 859 19133 879
rect 19153 859 19167 879
rect 19125 821 19167 859
rect 19217 879 19261 921
rect 19217 859 19229 879
rect 19249 859 19261 879
rect 19217 821 19261 859
rect 19333 879 19375 921
rect 19333 859 19341 879
rect 19361 859 19375 879
rect 19333 821 19375 859
rect 19425 879 19469 921
rect 19425 859 19437 879
rect 19457 859 19469 879
rect 19425 821 19469 859
rect 19546 879 19588 921
rect 19546 859 19554 879
rect 19574 859 19588 879
rect 19546 821 19588 859
rect 19638 879 19682 921
rect 19638 859 19650 879
rect 19670 859 19682 879
rect 19638 821 19682 859
rect 6644 375 6688 413
rect 1588 334 1632 372
rect 1588 314 1600 334
rect 1620 314 1632 334
rect 1588 272 1632 314
rect 1682 334 1724 372
rect 1682 314 1696 334
rect 1716 314 1724 334
rect 1682 272 1724 314
rect 1801 334 1845 372
rect 1801 314 1813 334
rect 1833 314 1845 334
rect 1801 272 1845 314
rect 1895 334 1937 372
rect 1895 314 1909 334
rect 1929 314 1937 334
rect 1895 272 1937 314
rect 2009 334 2053 372
rect 2009 314 2021 334
rect 2041 314 2053 334
rect 2009 272 2053 314
rect 2103 334 2145 372
rect 2103 314 2117 334
rect 2137 314 2145 334
rect 2103 272 2145 314
rect 2219 334 2261 372
rect 2219 314 2227 334
rect 2247 314 2261 334
rect 2219 272 2261 314
rect 2311 341 2356 372
rect 6644 355 6656 375
rect 6676 355 6688 375
rect 2311 334 2355 341
rect 2311 314 2323 334
rect 2343 314 2355 334
rect 2311 272 2355 314
rect 4538 314 4582 352
rect 4538 294 4550 314
rect 4570 294 4582 314
rect 4538 252 4582 294
rect 4632 314 4674 352
rect 4632 294 4646 314
rect 4666 294 4674 314
rect 4632 252 4674 294
rect 4751 314 4795 352
rect 4751 294 4763 314
rect 4783 294 4795 314
rect 4751 252 4795 294
rect 4845 314 4887 352
rect 4845 294 4859 314
rect 4879 294 4887 314
rect 4845 252 4887 294
rect 4959 314 5003 352
rect 4959 294 4971 314
rect 4991 294 5003 314
rect 4959 252 5003 294
rect 5053 314 5095 352
rect 5053 294 5067 314
rect 5087 294 5095 314
rect 5053 252 5095 294
rect 5169 314 5211 352
rect 5169 294 5177 314
rect 5197 294 5211 314
rect 5169 252 5211 294
rect 5261 321 5306 352
rect 5261 314 5305 321
rect 5261 294 5273 314
rect 5293 294 5305 314
rect 6644 313 6688 355
rect 6738 375 6780 413
rect 6738 355 6752 375
rect 6772 355 6780 375
rect 6738 313 6780 355
rect 6857 375 6901 413
rect 6857 355 6869 375
rect 6889 355 6901 375
rect 6857 313 6901 355
rect 6951 375 6993 413
rect 6951 355 6965 375
rect 6985 355 6993 375
rect 6951 313 6993 355
rect 7065 375 7109 413
rect 7065 355 7077 375
rect 7097 355 7109 375
rect 7065 313 7109 355
rect 7159 375 7201 413
rect 7159 355 7173 375
rect 7193 355 7201 375
rect 7159 313 7201 355
rect 7275 375 7317 413
rect 7275 355 7283 375
rect 7303 355 7317 375
rect 7275 313 7317 355
rect 7367 382 7412 413
rect 7367 375 7411 382
rect 16675 380 16719 418
rect 7367 355 7379 375
rect 7399 355 7411 375
rect 7367 313 7411 355
rect 11619 339 11663 377
rect 5261 252 5305 294
rect 11619 319 11631 339
rect 11651 319 11663 339
rect 11619 277 11663 319
rect 11713 339 11755 377
rect 11713 319 11727 339
rect 11747 319 11755 339
rect 11713 277 11755 319
rect 11832 339 11876 377
rect 11832 319 11844 339
rect 11864 319 11876 339
rect 11832 277 11876 319
rect 11926 339 11968 377
rect 11926 319 11940 339
rect 11960 319 11968 339
rect 11926 277 11968 319
rect 12040 339 12084 377
rect 12040 319 12052 339
rect 12072 319 12084 339
rect 12040 277 12084 319
rect 12134 339 12176 377
rect 12134 319 12148 339
rect 12168 319 12176 339
rect 12134 277 12176 319
rect 12250 339 12292 377
rect 12250 319 12258 339
rect 12278 319 12292 339
rect 12250 277 12292 319
rect 12342 346 12387 377
rect 16675 360 16687 380
rect 16707 360 16719 380
rect 12342 339 12386 346
rect 12342 319 12354 339
rect 12374 319 12386 339
rect 12342 277 12386 319
rect 14569 319 14613 357
rect 14569 299 14581 319
rect 14601 299 14613 319
rect 9472 198 9516 236
rect 9472 178 9484 198
rect 9504 178 9516 198
rect 9472 136 9516 178
rect 9566 198 9608 236
rect 9566 178 9580 198
rect 9600 178 9608 198
rect 9566 136 9608 178
rect 9685 198 9729 236
rect 9685 178 9697 198
rect 9717 178 9729 198
rect 9685 136 9729 178
rect 9779 198 9821 236
rect 9779 178 9793 198
rect 9813 178 9821 198
rect 9779 136 9821 178
rect 9893 198 9937 236
rect 9893 178 9905 198
rect 9925 178 9937 198
rect 9893 136 9937 178
rect 9987 198 10029 236
rect 9987 178 10001 198
rect 10021 178 10029 198
rect 9987 136 10029 178
rect 10103 198 10145 236
rect 10103 178 10111 198
rect 10131 178 10145 198
rect 10103 136 10145 178
rect 10195 205 10240 236
rect 10195 198 10239 205
rect 14569 257 14613 299
rect 14663 319 14705 357
rect 14663 299 14677 319
rect 14697 299 14705 319
rect 14663 257 14705 299
rect 14782 319 14826 357
rect 14782 299 14794 319
rect 14814 299 14826 319
rect 14782 257 14826 299
rect 14876 319 14918 357
rect 14876 299 14890 319
rect 14910 299 14918 319
rect 14876 257 14918 299
rect 14990 319 15034 357
rect 14990 299 15002 319
rect 15022 299 15034 319
rect 14990 257 15034 299
rect 15084 319 15126 357
rect 15084 299 15098 319
rect 15118 299 15126 319
rect 15084 257 15126 299
rect 15200 319 15242 357
rect 15200 299 15208 319
rect 15228 299 15242 319
rect 15200 257 15242 299
rect 15292 326 15337 357
rect 15292 319 15336 326
rect 15292 299 15304 319
rect 15324 299 15336 319
rect 16675 318 16719 360
rect 16769 380 16811 418
rect 16769 360 16783 380
rect 16803 360 16811 380
rect 16769 318 16811 360
rect 16888 380 16932 418
rect 16888 360 16900 380
rect 16920 360 16932 380
rect 16888 318 16932 360
rect 16982 380 17024 418
rect 16982 360 16996 380
rect 17016 360 17024 380
rect 16982 318 17024 360
rect 17096 380 17140 418
rect 17096 360 17108 380
rect 17128 360 17140 380
rect 17096 318 17140 360
rect 17190 380 17232 418
rect 17190 360 17204 380
rect 17224 360 17232 380
rect 17190 318 17232 360
rect 17306 380 17348 418
rect 17306 360 17314 380
rect 17334 360 17348 380
rect 17306 318 17348 360
rect 17398 387 17443 418
rect 17398 380 17442 387
rect 17398 360 17410 380
rect 17430 360 17442 380
rect 17398 318 17442 360
rect 15292 257 15336 299
rect 10195 178 10207 198
rect 10227 178 10239 198
rect 10195 136 10239 178
<< ndiffc >>
rect 5172 9325 5190 9343
rect 116 9284 134 9302
rect 3831 9237 3851 9257
rect 3934 9233 3954 9253
rect 4042 9233 4062 9253
rect 4145 9237 4165 9257
rect 4250 9233 4270 9253
rect 4353 9237 4373 9257
rect 4463 9233 4483 9253
rect 8887 9278 8907 9298
rect 8990 9274 9010 9294
rect 9098 9274 9118 9294
rect 9201 9278 9221 9298
rect 9306 9274 9326 9294
rect 9409 9278 9429 9298
rect 9519 9274 9539 9294
rect 15203 9330 15221 9348
rect 9622 9278 9642 9298
rect 10147 9289 10165 9307
rect 4566 9237 4586 9257
rect 118 9185 136 9203
rect 116 9097 134 9115
rect 5174 9226 5192 9244
rect 118 8998 136 9016
rect 344 8999 364 9019
rect 447 9003 467 9023
rect 557 8999 577 9019
rect 660 9003 680 9023
rect 765 8999 785 9019
rect 868 9003 888 9023
rect 976 9003 996 9023
rect 1079 8999 1099 9019
rect 4793 9145 4811 9163
rect 5172 9138 5190 9156
rect 13862 9242 13882 9262
rect 13965 9238 13985 9258
rect 14073 9238 14093 9258
rect 14176 9242 14196 9262
rect 14281 9238 14301 9258
rect 14384 9242 14404 9262
rect 14494 9238 14514 9258
rect 18918 9283 18938 9303
rect 19021 9279 19041 9299
rect 19129 9279 19149 9299
rect 19232 9283 19252 9303
rect 19337 9279 19357 9299
rect 19440 9283 19460 9303
rect 19550 9279 19570 9299
rect 19653 9283 19673 9303
rect 14597 9242 14617 9262
rect 4795 9046 4813 9064
rect 5174 9039 5192 9057
rect 5400 9040 5420 9060
rect 5503 9044 5523 9064
rect 5613 9040 5633 9060
rect 5716 9044 5736 9064
rect 5821 9040 5841 9060
rect 5924 9044 5944 9064
rect 6032 9044 6052 9064
rect 6135 9040 6155 9060
rect 9849 9186 9867 9204
rect 10149 9190 10167 9208
rect 9851 9087 9869 9105
rect 10147 9102 10165 9120
rect 15205 9231 15223 9249
rect 116 8868 134 8886
rect 2892 8927 2912 8947
rect 2995 8923 3015 8943
rect 3103 8923 3123 8943
rect 3206 8927 3226 8947
rect 3311 8923 3331 8943
rect 3414 8927 3434 8947
rect 3524 8923 3544 8943
rect 3627 8927 3647 8947
rect 118 8769 136 8787
rect 4793 8915 4811 8933
rect 5172 8909 5190 8927
rect 1282 8755 1302 8775
rect 1385 8759 1405 8779
rect 1495 8755 1515 8775
rect 1598 8759 1618 8779
rect 1703 8755 1723 8775
rect 1806 8759 1826 8779
rect 1914 8759 1934 8779
rect 2017 8755 2037 8775
rect 10149 9003 10167 9021
rect 7948 8968 7968 8988
rect 8051 8964 8071 8984
rect 8159 8964 8179 8984
rect 8262 8968 8282 8988
rect 8367 8964 8387 8984
rect 8470 8968 8490 8988
rect 8580 8964 8600 8984
rect 8683 8968 8703 8988
rect 10375 9004 10395 9024
rect 10478 9008 10498 9028
rect 10588 9004 10608 9024
rect 10691 9008 10711 9028
rect 10796 9004 10816 9024
rect 10899 9008 10919 9028
rect 11007 9008 11027 9028
rect 11110 9004 11130 9024
rect 14824 9150 14842 9168
rect 15203 9143 15221 9161
rect 14826 9051 14844 9069
rect 15205 9044 15223 9062
rect 15431 9045 15451 9065
rect 15534 9049 15554 9069
rect 15644 9045 15664 9065
rect 15747 9049 15767 9069
rect 15852 9045 15872 9065
rect 15955 9049 15975 9069
rect 16063 9049 16083 9069
rect 16166 9045 16186 9065
rect 19880 9191 19898 9209
rect 19882 9092 19900 9110
rect 4795 8816 4813 8834
rect 5174 8810 5192 8828
rect 9849 8956 9867 8974
rect 6338 8796 6358 8816
rect 6441 8800 6461 8820
rect 6551 8796 6571 8816
rect 6654 8800 6674 8820
rect 6759 8796 6779 8816
rect 6862 8800 6882 8820
rect 6970 8800 6990 8820
rect 7073 8796 7093 8816
rect 9851 8857 9869 8875
rect 10147 8873 10165 8891
rect 12923 8932 12943 8952
rect 13026 8928 13046 8948
rect 13134 8928 13154 8948
rect 13237 8932 13257 8952
rect 13342 8928 13362 8948
rect 13445 8932 13465 8952
rect 13555 8928 13575 8948
rect 13658 8932 13678 8952
rect 10149 8774 10167 8792
rect 14824 8920 14842 8938
rect 15203 8914 15221 8932
rect 116 8638 134 8656
rect 118 8539 136 8557
rect 3830 8683 3850 8703
rect 3933 8679 3953 8699
rect 4041 8679 4061 8699
rect 4144 8683 4164 8703
rect 4249 8679 4269 8699
rect 4352 8683 4372 8703
rect 4462 8679 4482 8699
rect 4565 8683 4585 8703
rect 4793 8686 4811 8704
rect 5172 8679 5190 8697
rect 4795 8587 4813 8605
rect 5174 8580 5192 8598
rect 8886 8724 8906 8744
rect 8989 8720 9009 8740
rect 9097 8720 9117 8740
rect 9200 8724 9220 8744
rect 9305 8720 9325 8740
rect 9408 8724 9428 8744
rect 9518 8720 9538 8740
rect 9621 8724 9641 8744
rect 11313 8760 11333 8780
rect 11416 8764 11436 8784
rect 11526 8760 11546 8780
rect 11629 8764 11649 8784
rect 11734 8760 11754 8780
rect 11837 8764 11857 8784
rect 11945 8764 11965 8784
rect 12048 8760 12068 8780
rect 9849 8727 9867 8745
rect 17979 8973 17999 8993
rect 18082 8969 18102 8989
rect 18190 8969 18210 8989
rect 18293 8973 18313 8993
rect 18398 8969 18418 8989
rect 18501 8973 18521 8993
rect 18611 8969 18631 8989
rect 18714 8973 18734 8993
rect 14826 8821 14844 8839
rect 15205 8815 15223 8833
rect 19880 8961 19898 8979
rect 16369 8801 16389 8821
rect 16472 8805 16492 8825
rect 16582 8801 16602 8821
rect 16685 8805 16705 8825
rect 16790 8801 16810 8821
rect 16893 8805 16913 8825
rect 17001 8805 17021 8825
rect 17104 8801 17124 8821
rect 19882 8862 19900 8880
rect 4793 8499 4811 8517
rect 9851 8628 9869 8646
rect 10147 8643 10165 8661
rect 9849 8540 9867 8558
rect 10149 8544 10167 8562
rect 13861 8688 13881 8708
rect 13964 8684 13984 8704
rect 14072 8684 14092 8704
rect 14175 8688 14195 8708
rect 14280 8684 14300 8704
rect 14383 8688 14403 8708
rect 14493 8684 14513 8704
rect 14596 8688 14616 8708
rect 14824 8691 14842 8709
rect 15203 8684 15221 8702
rect 5399 8486 5419 8506
rect 343 8445 363 8465
rect 446 8449 466 8469
rect 556 8445 576 8465
rect 659 8449 679 8469
rect 764 8445 784 8465
rect 867 8449 887 8469
rect 975 8449 995 8469
rect 1078 8445 1098 8465
rect 2752 8416 2772 8436
rect 2855 8412 2875 8432
rect 2963 8412 2983 8432
rect 3066 8416 3086 8436
rect 3171 8412 3191 8432
rect 3274 8416 3294 8436
rect 3384 8412 3404 8432
rect 3487 8416 3507 8436
rect 5502 8490 5522 8510
rect 5612 8486 5632 8506
rect 5715 8490 5735 8510
rect 5820 8486 5840 8506
rect 5923 8490 5943 8510
rect 6031 8490 6051 8510
rect 6134 8486 6154 8506
rect 7808 8457 7828 8477
rect 7911 8453 7931 8473
rect 8019 8453 8039 8473
rect 8122 8457 8142 8477
rect 8227 8453 8247 8473
rect 8330 8457 8350 8477
rect 8440 8453 8460 8473
rect 8543 8457 8563 8477
rect 14826 8592 14844 8610
rect 15205 8585 15223 8603
rect 18917 8729 18937 8749
rect 19020 8725 19040 8745
rect 19128 8725 19148 8745
rect 19231 8729 19251 8749
rect 19336 8725 19356 8745
rect 19439 8729 19459 8749
rect 19549 8725 19569 8745
rect 19652 8729 19672 8749
rect 19880 8732 19898 8750
rect 14824 8504 14842 8522
rect 19882 8633 19900 8651
rect 19880 8545 19898 8563
rect 15430 8491 15450 8511
rect 4795 8400 4813 8418
rect 117 8181 135 8199
rect 9851 8441 9869 8459
rect 10374 8450 10394 8470
rect 10477 8454 10497 8474
rect 10587 8450 10607 8470
rect 10690 8454 10710 8474
rect 10795 8450 10815 8470
rect 10898 8454 10918 8474
rect 11006 8454 11026 8474
rect 11109 8450 11129 8470
rect 12783 8421 12803 8441
rect 12886 8417 12906 8437
rect 12994 8417 13014 8437
rect 13097 8421 13117 8441
rect 13202 8417 13222 8437
rect 13305 8421 13325 8441
rect 13415 8417 13435 8437
rect 13518 8421 13538 8441
rect 15533 8495 15553 8515
rect 15643 8491 15663 8511
rect 15746 8495 15766 8515
rect 15851 8491 15871 8511
rect 15954 8495 15974 8515
rect 16062 8495 16082 8515
rect 16165 8491 16185 8511
rect 17839 8462 17859 8482
rect 17942 8458 17962 8478
rect 18050 8458 18070 8478
rect 18153 8462 18173 8482
rect 18258 8458 18278 8478
rect 18361 8462 18381 8482
rect 18471 8458 18491 8478
rect 18574 8462 18594 8482
rect 5173 8222 5191 8240
rect 14826 8405 14844 8423
rect 1423 8163 1443 8183
rect 1526 8167 1546 8187
rect 1636 8163 1656 8183
rect 1739 8167 1759 8187
rect 1844 8163 1864 8183
rect 1947 8167 1967 8187
rect 2055 8167 2075 8187
rect 2158 8163 2178 8183
rect 3832 8134 3852 8154
rect 3935 8130 3955 8150
rect 4043 8130 4063 8150
rect 4146 8134 4166 8154
rect 4251 8130 4271 8150
rect 4354 8134 4374 8154
rect 4464 8130 4484 8150
rect 6479 8204 6499 8224
rect 6582 8208 6602 8228
rect 6692 8204 6712 8224
rect 6795 8208 6815 8228
rect 6900 8204 6920 8224
rect 7003 8208 7023 8228
rect 7111 8208 7131 8228
rect 7214 8204 7234 8224
rect 8888 8175 8908 8195
rect 8991 8171 9011 8191
rect 9099 8171 9119 8191
rect 9202 8175 9222 8195
rect 9307 8171 9327 8191
rect 9410 8175 9430 8195
rect 9520 8171 9540 8191
rect 9623 8175 9643 8195
rect 10148 8186 10166 8204
rect 19882 8446 19900 8464
rect 15204 8227 15222 8245
rect 4567 8134 4587 8154
rect 119 8082 137 8100
rect 117 7994 135 8012
rect 5175 8123 5193 8141
rect 119 7895 137 7913
rect 345 7896 365 7916
rect 448 7900 468 7920
rect 558 7896 578 7916
rect 661 7900 681 7920
rect 766 7896 786 7916
rect 869 7900 889 7920
rect 977 7900 997 7920
rect 1080 7896 1100 7916
rect 4794 8042 4812 8060
rect 5173 8035 5191 8053
rect 11454 8168 11474 8188
rect 11557 8172 11577 8192
rect 11667 8168 11687 8188
rect 11770 8172 11790 8192
rect 11875 8168 11895 8188
rect 11978 8172 11998 8192
rect 12086 8172 12106 8192
rect 12189 8168 12209 8188
rect 13863 8139 13883 8159
rect 13966 8135 13986 8155
rect 14074 8135 14094 8155
rect 14177 8139 14197 8159
rect 14282 8135 14302 8155
rect 14385 8139 14405 8159
rect 14495 8135 14515 8155
rect 16510 8209 16530 8229
rect 16613 8213 16633 8233
rect 16723 8209 16743 8229
rect 16826 8213 16846 8233
rect 16931 8209 16951 8229
rect 17034 8213 17054 8233
rect 17142 8213 17162 8233
rect 17245 8209 17265 8229
rect 18919 8180 18939 8200
rect 19022 8176 19042 8196
rect 19130 8176 19150 8196
rect 19233 8180 19253 8200
rect 19338 8176 19358 8196
rect 19441 8180 19461 8200
rect 19551 8176 19571 8196
rect 19654 8180 19674 8200
rect 14598 8139 14618 8159
rect 4796 7943 4814 7961
rect 5175 7936 5193 7954
rect 5401 7937 5421 7957
rect 5504 7941 5524 7961
rect 5614 7937 5634 7957
rect 5717 7941 5737 7961
rect 5822 7937 5842 7957
rect 5925 7941 5945 7961
rect 6033 7941 6053 7961
rect 6136 7937 6156 7957
rect 9850 8083 9868 8101
rect 10150 8087 10168 8105
rect 9852 7984 9870 8002
rect 10148 7999 10166 8017
rect 15206 8128 15224 8146
rect 117 7765 135 7783
rect 2893 7824 2913 7844
rect 2996 7820 3016 7840
rect 3104 7820 3124 7840
rect 3207 7824 3227 7844
rect 3312 7820 3332 7840
rect 3415 7824 3435 7844
rect 3525 7820 3545 7840
rect 3628 7824 3648 7844
rect 119 7666 137 7684
rect 4794 7812 4812 7830
rect 5173 7806 5191 7824
rect 1283 7652 1303 7672
rect 1386 7656 1406 7676
rect 1496 7652 1516 7672
rect 1599 7656 1619 7676
rect 1704 7652 1724 7672
rect 1807 7656 1827 7676
rect 1915 7656 1935 7676
rect 2018 7652 2038 7672
rect 10150 7900 10168 7918
rect 7949 7865 7969 7885
rect 8052 7861 8072 7881
rect 8160 7861 8180 7881
rect 8263 7865 8283 7885
rect 8368 7861 8388 7881
rect 8471 7865 8491 7885
rect 8581 7861 8601 7881
rect 8684 7865 8704 7885
rect 10376 7901 10396 7921
rect 10479 7905 10499 7925
rect 10589 7901 10609 7921
rect 10692 7905 10712 7925
rect 10797 7901 10817 7921
rect 10900 7905 10920 7925
rect 11008 7905 11028 7925
rect 11111 7901 11131 7921
rect 14825 8047 14843 8065
rect 15204 8040 15222 8058
rect 14827 7948 14845 7966
rect 15206 7941 15224 7959
rect 15432 7942 15452 7962
rect 15535 7946 15555 7966
rect 15645 7942 15665 7962
rect 15748 7946 15768 7966
rect 15853 7942 15873 7962
rect 15956 7946 15976 7966
rect 16064 7946 16084 7966
rect 16167 7942 16187 7962
rect 19881 8088 19899 8106
rect 19883 7989 19901 8007
rect 4796 7713 4814 7731
rect 5175 7707 5193 7725
rect 9850 7853 9868 7871
rect 6339 7693 6359 7713
rect 6442 7697 6462 7717
rect 6552 7693 6572 7713
rect 6655 7697 6675 7717
rect 6760 7693 6780 7713
rect 6863 7697 6883 7717
rect 6971 7697 6991 7717
rect 7074 7693 7094 7713
rect 9852 7754 9870 7772
rect 10148 7770 10166 7788
rect 12924 7829 12944 7849
rect 13027 7825 13047 7845
rect 13135 7825 13155 7845
rect 13238 7829 13258 7849
rect 13343 7825 13363 7845
rect 13446 7829 13466 7849
rect 13556 7825 13576 7845
rect 13659 7829 13679 7849
rect 10150 7671 10168 7689
rect 14825 7817 14843 7835
rect 15204 7811 15222 7829
rect 117 7535 135 7553
rect 119 7436 137 7454
rect 3831 7580 3851 7600
rect 3934 7576 3954 7596
rect 4042 7576 4062 7596
rect 4145 7580 4165 7600
rect 4250 7576 4270 7596
rect 4353 7580 4373 7600
rect 4463 7576 4483 7596
rect 4566 7580 4586 7600
rect 4794 7583 4812 7601
rect 5173 7576 5191 7594
rect 4796 7484 4814 7502
rect 5175 7477 5193 7495
rect 8887 7621 8907 7641
rect 8990 7617 9010 7637
rect 9098 7617 9118 7637
rect 9201 7621 9221 7641
rect 9306 7617 9326 7637
rect 9409 7621 9429 7641
rect 9519 7617 9539 7637
rect 9622 7621 9642 7641
rect 11314 7657 11334 7677
rect 11417 7661 11437 7681
rect 11527 7657 11547 7677
rect 11630 7661 11650 7681
rect 11735 7657 11755 7677
rect 11838 7661 11858 7681
rect 11946 7661 11966 7681
rect 12049 7657 12069 7677
rect 9850 7624 9868 7642
rect 17980 7870 18000 7890
rect 18083 7866 18103 7886
rect 18191 7866 18211 7886
rect 18294 7870 18314 7890
rect 18399 7866 18419 7886
rect 18502 7870 18522 7890
rect 18612 7866 18632 7886
rect 18715 7870 18735 7890
rect 14827 7718 14845 7736
rect 15206 7712 15224 7730
rect 19881 7858 19899 7876
rect 16370 7698 16390 7718
rect 16473 7702 16493 7722
rect 16583 7698 16603 7718
rect 16686 7702 16706 7722
rect 16791 7698 16811 7718
rect 16894 7702 16914 7722
rect 17002 7702 17022 7722
rect 17105 7698 17125 7718
rect 19883 7759 19901 7777
rect 4794 7396 4812 7414
rect 9852 7525 9870 7543
rect 10148 7540 10166 7558
rect 9850 7437 9868 7455
rect 10150 7441 10168 7459
rect 13862 7585 13882 7605
rect 13965 7581 13985 7601
rect 14073 7581 14093 7601
rect 14176 7585 14196 7605
rect 14281 7581 14301 7601
rect 14384 7585 14404 7605
rect 14494 7581 14514 7601
rect 14597 7585 14617 7605
rect 14825 7588 14843 7606
rect 15204 7581 15222 7599
rect 5400 7383 5420 7403
rect 344 7342 364 7362
rect 447 7346 467 7366
rect 557 7342 577 7362
rect 660 7346 680 7366
rect 765 7342 785 7362
rect 868 7346 888 7366
rect 976 7346 996 7366
rect 1079 7342 1099 7362
rect 2783 7300 2803 7320
rect 2886 7296 2906 7316
rect 2994 7296 3014 7316
rect 3097 7300 3117 7320
rect 3202 7296 3222 7316
rect 3305 7300 3325 7320
rect 3415 7296 3435 7316
rect 3518 7300 3538 7320
rect 5503 7387 5523 7407
rect 5613 7383 5633 7403
rect 5716 7387 5736 7407
rect 5821 7383 5841 7403
rect 5924 7387 5944 7407
rect 6032 7387 6052 7407
rect 6135 7383 6155 7403
rect 7839 7341 7859 7361
rect 4796 7297 4814 7315
rect 7942 7337 7962 7357
rect 8050 7337 8070 7357
rect 8153 7341 8173 7361
rect 8258 7337 8278 7357
rect 8361 7341 8381 7361
rect 8471 7337 8491 7357
rect 8574 7341 8594 7361
rect 14827 7489 14845 7507
rect 15206 7482 15224 7500
rect 18918 7626 18938 7646
rect 19021 7622 19041 7642
rect 19129 7622 19149 7642
rect 19232 7626 19252 7646
rect 19337 7622 19357 7642
rect 19440 7626 19460 7646
rect 19550 7622 19570 7642
rect 19653 7626 19673 7646
rect 19881 7629 19899 7647
rect 14825 7401 14843 7419
rect 19883 7530 19901 7548
rect 19881 7442 19899 7460
rect 15431 7388 15451 7408
rect 9852 7338 9870 7356
rect 10375 7347 10395 7367
rect 10478 7351 10498 7371
rect 10588 7347 10608 7367
rect 10691 7351 10711 7371
rect 10796 7347 10816 7367
rect 10899 7351 10919 7371
rect 11007 7351 11027 7371
rect 11110 7347 11130 7367
rect 12814 7305 12834 7325
rect 12917 7301 12937 7321
rect 13025 7301 13045 7321
rect 13128 7305 13148 7325
rect 13233 7301 13253 7321
rect 13336 7305 13356 7325
rect 13446 7301 13466 7321
rect 13549 7305 13569 7325
rect 15534 7392 15554 7412
rect 15644 7388 15664 7408
rect 15747 7392 15767 7412
rect 15852 7388 15872 7408
rect 15955 7392 15975 7412
rect 16063 7392 16083 7412
rect 16166 7388 16186 7408
rect 17870 7346 17890 7366
rect 14827 7302 14845 7320
rect 17973 7342 17993 7362
rect 18081 7342 18101 7362
rect 18184 7346 18204 7366
rect 18289 7342 18309 7362
rect 18392 7346 18412 7366
rect 18502 7342 18522 7362
rect 18605 7346 18625 7366
rect 19883 7343 19901 7361
rect 117 7078 135 7096
rect 1393 7073 1413 7093
rect 1496 7077 1516 7097
rect 1606 7073 1626 7093
rect 1709 7077 1729 7097
rect 1814 7073 1834 7093
rect 1917 7077 1937 7097
rect 2025 7077 2045 7097
rect 5173 7119 5191 7137
rect 2128 7073 2148 7093
rect 3832 7031 3852 7051
rect 3935 7027 3955 7047
rect 4043 7027 4063 7047
rect 4146 7031 4166 7051
rect 4251 7027 4271 7047
rect 4354 7031 4374 7051
rect 4464 7027 4484 7047
rect 6449 7114 6469 7134
rect 6552 7118 6572 7138
rect 6662 7114 6682 7134
rect 6765 7118 6785 7138
rect 6870 7114 6890 7134
rect 6973 7118 6993 7138
rect 7081 7118 7101 7138
rect 7184 7114 7204 7134
rect 8888 7072 8908 7092
rect 8991 7068 9011 7088
rect 9099 7068 9119 7088
rect 9202 7072 9222 7092
rect 9307 7068 9327 7088
rect 9410 7072 9430 7092
rect 9520 7068 9540 7088
rect 9623 7072 9643 7092
rect 10148 7083 10166 7101
rect 4567 7031 4587 7051
rect 119 6979 137 6997
rect 117 6891 135 6909
rect 5175 7020 5193 7038
rect 119 6792 137 6810
rect 345 6793 365 6813
rect 448 6797 468 6817
rect 558 6793 578 6813
rect 661 6797 681 6817
rect 766 6793 786 6813
rect 869 6797 889 6817
rect 977 6797 997 6817
rect 1080 6793 1100 6813
rect 4794 6939 4812 6957
rect 5173 6932 5191 6950
rect 11424 7078 11444 7098
rect 11527 7082 11547 7102
rect 11637 7078 11657 7098
rect 11740 7082 11760 7102
rect 11845 7078 11865 7098
rect 11948 7082 11968 7102
rect 12056 7082 12076 7102
rect 15204 7124 15222 7142
rect 12159 7078 12179 7098
rect 13863 7036 13883 7056
rect 13966 7032 13986 7052
rect 14074 7032 14094 7052
rect 14177 7036 14197 7056
rect 14282 7032 14302 7052
rect 14385 7036 14405 7056
rect 14495 7032 14515 7052
rect 16480 7119 16500 7139
rect 16583 7123 16603 7143
rect 16693 7119 16713 7139
rect 16796 7123 16816 7143
rect 16901 7119 16921 7139
rect 17004 7123 17024 7143
rect 17112 7123 17132 7143
rect 17215 7119 17235 7139
rect 18919 7077 18939 7097
rect 19022 7073 19042 7093
rect 19130 7073 19150 7093
rect 19233 7077 19253 7097
rect 19338 7073 19358 7093
rect 19441 7077 19461 7097
rect 19551 7073 19571 7093
rect 19654 7077 19674 7097
rect 14598 7036 14618 7056
rect 4796 6840 4814 6858
rect 5175 6833 5193 6851
rect 5401 6834 5421 6854
rect 5504 6838 5524 6858
rect 5614 6834 5634 6854
rect 5717 6838 5737 6858
rect 5822 6834 5842 6854
rect 5925 6838 5945 6858
rect 6033 6838 6053 6858
rect 6136 6834 6156 6854
rect 9850 6980 9868 6998
rect 10150 6984 10168 7002
rect 9852 6881 9870 6899
rect 10148 6896 10166 6914
rect 15206 7025 15224 7043
rect 117 6662 135 6680
rect 2893 6721 2913 6741
rect 2996 6717 3016 6737
rect 3104 6717 3124 6737
rect 3207 6721 3227 6741
rect 3312 6717 3332 6737
rect 3415 6721 3435 6741
rect 3525 6717 3545 6737
rect 3628 6721 3648 6741
rect 119 6563 137 6581
rect 4794 6709 4812 6727
rect 5173 6703 5191 6721
rect 1283 6549 1303 6569
rect 1386 6553 1406 6573
rect 1496 6549 1516 6569
rect 1599 6553 1619 6573
rect 1704 6549 1724 6569
rect 1807 6553 1827 6573
rect 1915 6553 1935 6573
rect 2018 6549 2038 6569
rect 10150 6797 10168 6815
rect 7949 6762 7969 6782
rect 8052 6758 8072 6778
rect 8160 6758 8180 6778
rect 8263 6762 8283 6782
rect 8368 6758 8388 6778
rect 8471 6762 8491 6782
rect 8581 6758 8601 6778
rect 8684 6762 8704 6782
rect 10376 6798 10396 6818
rect 10479 6802 10499 6822
rect 10589 6798 10609 6818
rect 10692 6802 10712 6822
rect 10797 6798 10817 6818
rect 10900 6802 10920 6822
rect 11008 6802 11028 6822
rect 11111 6798 11131 6818
rect 14825 6944 14843 6962
rect 15204 6937 15222 6955
rect 14827 6845 14845 6863
rect 15206 6838 15224 6856
rect 15432 6839 15452 6859
rect 15535 6843 15555 6863
rect 15645 6839 15665 6859
rect 15748 6843 15768 6863
rect 15853 6839 15873 6859
rect 15956 6843 15976 6863
rect 16064 6843 16084 6863
rect 16167 6839 16187 6859
rect 19881 6985 19899 7003
rect 19883 6886 19901 6904
rect 4796 6610 4814 6628
rect 5175 6604 5193 6622
rect 9850 6750 9868 6768
rect 6339 6590 6359 6610
rect 6442 6594 6462 6614
rect 6552 6590 6572 6610
rect 6655 6594 6675 6614
rect 6760 6590 6780 6610
rect 6863 6594 6883 6614
rect 6971 6594 6991 6614
rect 7074 6590 7094 6610
rect 9852 6651 9870 6669
rect 10148 6667 10166 6685
rect 12924 6726 12944 6746
rect 13027 6722 13047 6742
rect 13135 6722 13155 6742
rect 13238 6726 13258 6746
rect 13343 6722 13363 6742
rect 13446 6726 13466 6746
rect 13556 6722 13576 6742
rect 13659 6726 13679 6746
rect 10150 6568 10168 6586
rect 14825 6714 14843 6732
rect 15204 6708 15222 6726
rect 117 6432 135 6450
rect 119 6333 137 6351
rect 3831 6477 3851 6497
rect 3934 6473 3954 6493
rect 4042 6473 4062 6493
rect 4145 6477 4165 6497
rect 4250 6473 4270 6493
rect 4353 6477 4373 6497
rect 4463 6473 4483 6493
rect 4566 6477 4586 6497
rect 4794 6480 4812 6498
rect 5173 6473 5191 6491
rect 4796 6381 4814 6399
rect 5175 6374 5193 6392
rect 8887 6518 8907 6538
rect 8990 6514 9010 6534
rect 9098 6514 9118 6534
rect 9201 6518 9221 6538
rect 9306 6514 9326 6534
rect 9409 6518 9429 6538
rect 9519 6514 9539 6534
rect 9622 6518 9642 6538
rect 11314 6554 11334 6574
rect 11417 6558 11437 6578
rect 11527 6554 11547 6574
rect 11630 6558 11650 6578
rect 11735 6554 11755 6574
rect 11838 6558 11858 6578
rect 11946 6558 11966 6578
rect 12049 6554 12069 6574
rect 9850 6521 9868 6539
rect 17980 6767 18000 6787
rect 18083 6763 18103 6783
rect 18191 6763 18211 6783
rect 18294 6767 18314 6787
rect 18399 6763 18419 6783
rect 18502 6767 18522 6787
rect 18612 6763 18632 6783
rect 18715 6767 18735 6787
rect 14827 6615 14845 6633
rect 15206 6609 15224 6627
rect 19881 6755 19899 6773
rect 16370 6595 16390 6615
rect 16473 6599 16493 6619
rect 16583 6595 16603 6615
rect 16686 6599 16706 6619
rect 16791 6595 16811 6615
rect 16894 6599 16914 6619
rect 17002 6599 17022 6619
rect 17105 6595 17125 6615
rect 19883 6656 19901 6674
rect 4794 6293 4812 6311
rect 9852 6422 9870 6440
rect 10148 6437 10166 6455
rect 9850 6334 9868 6352
rect 10150 6338 10168 6356
rect 13862 6482 13882 6502
rect 13965 6478 13985 6498
rect 14073 6478 14093 6498
rect 14176 6482 14196 6502
rect 14281 6478 14301 6498
rect 14384 6482 14404 6502
rect 14494 6478 14514 6498
rect 14597 6482 14617 6502
rect 14825 6485 14843 6503
rect 15204 6478 15222 6496
rect 5400 6280 5420 6300
rect 344 6239 364 6259
rect 447 6243 467 6263
rect 557 6239 577 6259
rect 660 6243 680 6263
rect 765 6239 785 6259
rect 868 6243 888 6263
rect 976 6243 996 6263
rect 1079 6239 1099 6259
rect 2753 6210 2773 6230
rect 2856 6206 2876 6226
rect 2964 6206 2984 6226
rect 3067 6210 3087 6230
rect 3172 6206 3192 6226
rect 3275 6210 3295 6230
rect 3385 6206 3405 6226
rect 3488 6210 3508 6230
rect 5503 6284 5523 6304
rect 5613 6280 5633 6300
rect 5716 6284 5736 6304
rect 5821 6280 5841 6300
rect 5924 6284 5944 6304
rect 6032 6284 6052 6304
rect 6135 6280 6155 6300
rect 7809 6251 7829 6271
rect 7912 6247 7932 6267
rect 8020 6247 8040 6267
rect 8123 6251 8143 6271
rect 8228 6247 8248 6267
rect 8331 6251 8351 6271
rect 8441 6247 8461 6267
rect 8544 6251 8564 6271
rect 14827 6386 14845 6404
rect 15206 6379 15224 6397
rect 18918 6523 18938 6543
rect 19021 6519 19041 6539
rect 19129 6519 19149 6539
rect 19232 6523 19252 6543
rect 19337 6519 19357 6539
rect 19440 6523 19460 6543
rect 19550 6519 19570 6539
rect 19653 6523 19673 6543
rect 19881 6526 19899 6544
rect 14825 6298 14843 6316
rect 19883 6427 19901 6445
rect 19881 6339 19899 6357
rect 15431 6285 15451 6305
rect 4796 6194 4814 6212
rect 118 5975 136 5993
rect 9852 6235 9870 6253
rect 10375 6244 10395 6264
rect 10478 6248 10498 6268
rect 10588 6244 10608 6264
rect 10691 6248 10711 6268
rect 10796 6244 10816 6264
rect 10899 6248 10919 6268
rect 11007 6248 11027 6268
rect 11110 6244 11130 6264
rect 12784 6215 12804 6235
rect 12887 6211 12907 6231
rect 12995 6211 13015 6231
rect 13098 6215 13118 6235
rect 13203 6211 13223 6231
rect 13306 6215 13326 6235
rect 13416 6211 13436 6231
rect 13519 6215 13539 6235
rect 15534 6289 15554 6309
rect 15644 6285 15664 6305
rect 15747 6289 15767 6309
rect 15852 6285 15872 6305
rect 15955 6289 15975 6309
rect 16063 6289 16083 6309
rect 16166 6285 16186 6305
rect 17840 6256 17860 6276
rect 17943 6252 17963 6272
rect 18051 6252 18071 6272
rect 18154 6256 18174 6276
rect 18259 6252 18279 6272
rect 18362 6256 18382 6276
rect 18472 6252 18492 6272
rect 18575 6256 18595 6276
rect 5174 6016 5192 6034
rect 14827 6199 14845 6217
rect 1424 5957 1444 5977
rect 1527 5961 1547 5981
rect 1637 5957 1657 5977
rect 1740 5961 1760 5981
rect 1845 5957 1865 5977
rect 1948 5961 1968 5981
rect 2056 5961 2076 5981
rect 2159 5957 2179 5977
rect 3833 5928 3853 5948
rect 3936 5924 3956 5944
rect 4044 5924 4064 5944
rect 4147 5928 4167 5948
rect 4252 5924 4272 5944
rect 4355 5928 4375 5948
rect 4465 5924 4485 5944
rect 6480 5998 6500 6018
rect 6583 6002 6603 6022
rect 6693 5998 6713 6018
rect 6796 6002 6816 6022
rect 6901 5998 6921 6018
rect 7004 6002 7024 6022
rect 7112 6002 7132 6022
rect 7215 5998 7235 6018
rect 8889 5969 8909 5989
rect 8992 5965 9012 5985
rect 9100 5965 9120 5985
rect 9203 5969 9223 5989
rect 9308 5965 9328 5985
rect 9411 5969 9431 5989
rect 9521 5965 9541 5985
rect 9624 5969 9644 5989
rect 10149 5980 10167 5998
rect 19883 6240 19901 6258
rect 15205 6021 15223 6039
rect 4568 5928 4588 5948
rect 120 5876 138 5894
rect 118 5788 136 5806
rect 5176 5917 5194 5935
rect 120 5689 138 5707
rect 346 5690 366 5710
rect 449 5694 469 5714
rect 559 5690 579 5710
rect 662 5694 682 5714
rect 767 5690 787 5710
rect 870 5694 890 5714
rect 978 5694 998 5714
rect 1081 5690 1101 5710
rect 4795 5836 4813 5854
rect 5174 5829 5192 5847
rect 11455 5962 11475 5982
rect 11558 5966 11578 5986
rect 11668 5962 11688 5982
rect 11771 5966 11791 5986
rect 11876 5962 11896 5982
rect 11979 5966 11999 5986
rect 12087 5966 12107 5986
rect 12190 5962 12210 5982
rect 13864 5933 13884 5953
rect 13967 5929 13987 5949
rect 14075 5929 14095 5949
rect 14178 5933 14198 5953
rect 14283 5929 14303 5949
rect 14386 5933 14406 5953
rect 14496 5929 14516 5949
rect 16511 6003 16531 6023
rect 16614 6007 16634 6027
rect 16724 6003 16744 6023
rect 16827 6007 16847 6027
rect 16932 6003 16952 6023
rect 17035 6007 17055 6027
rect 17143 6007 17163 6027
rect 17246 6003 17266 6023
rect 18920 5974 18940 5994
rect 19023 5970 19043 5990
rect 19131 5970 19151 5990
rect 19234 5974 19254 5994
rect 19339 5970 19359 5990
rect 19442 5974 19462 5994
rect 19552 5970 19572 5990
rect 19655 5974 19675 5994
rect 14599 5933 14619 5953
rect 4797 5737 4815 5755
rect 5176 5730 5194 5748
rect 5402 5731 5422 5751
rect 5505 5735 5525 5755
rect 5615 5731 5635 5751
rect 5718 5735 5738 5755
rect 5823 5731 5843 5751
rect 5926 5735 5946 5755
rect 6034 5735 6054 5755
rect 6137 5731 6157 5751
rect 9851 5877 9869 5895
rect 10151 5881 10169 5899
rect 9853 5778 9871 5796
rect 10149 5793 10167 5811
rect 15207 5922 15225 5940
rect 118 5559 136 5577
rect 2894 5618 2914 5638
rect 2997 5614 3017 5634
rect 3105 5614 3125 5634
rect 3208 5618 3228 5638
rect 3313 5614 3333 5634
rect 3416 5618 3436 5638
rect 3526 5614 3546 5634
rect 3629 5618 3649 5638
rect 120 5460 138 5478
rect 4795 5606 4813 5624
rect 5174 5600 5192 5618
rect 1284 5446 1304 5466
rect 1387 5450 1407 5470
rect 1497 5446 1517 5466
rect 1600 5450 1620 5470
rect 1705 5446 1725 5466
rect 1808 5450 1828 5470
rect 1916 5450 1936 5470
rect 2019 5446 2039 5466
rect 10151 5694 10169 5712
rect 7950 5659 7970 5679
rect 8053 5655 8073 5675
rect 8161 5655 8181 5675
rect 8264 5659 8284 5679
rect 8369 5655 8389 5675
rect 8472 5659 8492 5679
rect 8582 5655 8602 5675
rect 8685 5659 8705 5679
rect 10377 5695 10397 5715
rect 10480 5699 10500 5719
rect 10590 5695 10610 5715
rect 10693 5699 10713 5719
rect 10798 5695 10818 5715
rect 10901 5699 10921 5719
rect 11009 5699 11029 5719
rect 11112 5695 11132 5715
rect 14826 5841 14844 5859
rect 15205 5834 15223 5852
rect 14828 5742 14846 5760
rect 15207 5735 15225 5753
rect 15433 5736 15453 5756
rect 15536 5740 15556 5760
rect 15646 5736 15666 5756
rect 15749 5740 15769 5760
rect 15854 5736 15874 5756
rect 15957 5740 15977 5760
rect 16065 5740 16085 5760
rect 16168 5736 16188 5756
rect 19882 5882 19900 5900
rect 19884 5783 19902 5801
rect 4797 5507 4815 5525
rect 5176 5501 5194 5519
rect 9851 5647 9869 5665
rect 6340 5487 6360 5507
rect 6443 5491 6463 5511
rect 6553 5487 6573 5507
rect 6656 5491 6676 5511
rect 6761 5487 6781 5507
rect 6864 5491 6884 5511
rect 6972 5491 6992 5511
rect 7075 5487 7095 5507
rect 9853 5548 9871 5566
rect 10149 5564 10167 5582
rect 12925 5623 12945 5643
rect 13028 5619 13048 5639
rect 13136 5619 13156 5639
rect 13239 5623 13259 5643
rect 13344 5619 13364 5639
rect 13447 5623 13467 5643
rect 13557 5619 13577 5639
rect 13660 5623 13680 5643
rect 10151 5465 10169 5483
rect 14826 5611 14844 5629
rect 15205 5605 15223 5623
rect 118 5329 136 5347
rect 120 5230 138 5248
rect 3832 5374 3852 5394
rect 3935 5370 3955 5390
rect 4043 5370 4063 5390
rect 4146 5374 4166 5394
rect 4251 5370 4271 5390
rect 4354 5374 4374 5394
rect 4464 5370 4484 5390
rect 4567 5374 4587 5394
rect 4795 5377 4813 5395
rect 5174 5370 5192 5388
rect 4797 5278 4815 5296
rect 5176 5271 5194 5289
rect 8888 5415 8908 5435
rect 8991 5411 9011 5431
rect 9099 5411 9119 5431
rect 9202 5415 9222 5435
rect 9307 5411 9327 5431
rect 9410 5415 9430 5435
rect 9520 5411 9540 5431
rect 9623 5415 9643 5435
rect 11315 5451 11335 5471
rect 11418 5455 11438 5475
rect 11528 5451 11548 5471
rect 11631 5455 11651 5475
rect 11736 5451 11756 5471
rect 11839 5455 11859 5475
rect 11947 5455 11967 5475
rect 12050 5451 12070 5471
rect 9851 5418 9869 5436
rect 17981 5664 18001 5684
rect 18084 5660 18104 5680
rect 18192 5660 18212 5680
rect 18295 5664 18315 5684
rect 18400 5660 18420 5680
rect 18503 5664 18523 5684
rect 18613 5660 18633 5680
rect 18716 5664 18736 5684
rect 14828 5512 14846 5530
rect 15207 5506 15225 5524
rect 19882 5652 19900 5670
rect 16371 5492 16391 5512
rect 16474 5496 16494 5516
rect 16584 5492 16604 5512
rect 16687 5496 16707 5516
rect 16792 5492 16812 5512
rect 16895 5496 16915 5516
rect 17003 5496 17023 5516
rect 17106 5492 17126 5512
rect 19884 5553 19902 5571
rect 4795 5190 4813 5208
rect 9853 5319 9871 5337
rect 10149 5334 10167 5352
rect 9851 5231 9869 5249
rect 10151 5235 10169 5253
rect 13863 5379 13883 5399
rect 13966 5375 13986 5395
rect 14074 5375 14094 5395
rect 14177 5379 14197 5399
rect 14282 5375 14302 5395
rect 14385 5379 14405 5399
rect 14495 5375 14515 5395
rect 14598 5379 14618 5399
rect 14826 5382 14844 5400
rect 15205 5375 15223 5393
rect 345 5136 365 5156
rect 448 5140 468 5160
rect 558 5136 578 5156
rect 661 5140 681 5160
rect 766 5136 786 5156
rect 869 5140 889 5160
rect 977 5140 997 5160
rect 1080 5136 1100 5156
rect 5401 5177 5421 5197
rect 2785 5088 2805 5108
rect 2888 5084 2908 5104
rect 2996 5084 3016 5104
rect 3099 5088 3119 5108
rect 3204 5084 3224 5104
rect 3307 5088 3327 5108
rect 3417 5084 3437 5104
rect 3520 5088 3540 5108
rect 5504 5181 5524 5201
rect 5614 5177 5634 5197
rect 5717 5181 5737 5201
rect 5822 5177 5842 5197
rect 5925 5181 5945 5201
rect 6033 5181 6053 5201
rect 6136 5177 6156 5197
rect 4797 5091 4815 5109
rect 7841 5129 7861 5149
rect 7944 5125 7964 5145
rect 8052 5125 8072 5145
rect 8155 5129 8175 5149
rect 8260 5125 8280 5145
rect 8363 5129 8383 5149
rect 8473 5125 8493 5145
rect 8576 5129 8596 5149
rect 14828 5283 14846 5301
rect 15207 5276 15225 5294
rect 18919 5420 18939 5440
rect 19022 5416 19042 5436
rect 19130 5416 19150 5436
rect 19233 5420 19253 5440
rect 19338 5416 19358 5436
rect 19441 5420 19461 5440
rect 19551 5416 19571 5436
rect 19654 5420 19674 5440
rect 19882 5423 19900 5441
rect 14826 5195 14844 5213
rect 19884 5324 19902 5342
rect 19882 5236 19900 5254
rect 9853 5132 9871 5150
rect 10376 5141 10396 5161
rect 10479 5145 10499 5165
rect 10589 5141 10609 5161
rect 10692 5145 10712 5165
rect 10797 5141 10817 5161
rect 10900 5145 10920 5165
rect 11008 5145 11028 5165
rect 11111 5141 11131 5161
rect 15432 5182 15452 5202
rect 12816 5093 12836 5113
rect 118 4872 136 4890
rect 1393 4873 1413 4893
rect 1496 4877 1516 4897
rect 1606 4873 1626 4893
rect 1709 4877 1729 4897
rect 1814 4873 1834 4893
rect 1917 4877 1937 4897
rect 2025 4877 2045 4897
rect 2128 4873 2148 4893
rect 5174 4913 5192 4931
rect 3833 4825 3853 4845
rect 3936 4821 3956 4841
rect 4044 4821 4064 4841
rect 4147 4825 4167 4845
rect 4252 4821 4272 4841
rect 4355 4825 4375 4845
rect 4465 4821 4485 4841
rect 6449 4914 6469 4934
rect 6552 4918 6572 4938
rect 6662 4914 6682 4934
rect 6765 4918 6785 4938
rect 6870 4914 6890 4934
rect 6973 4918 6993 4938
rect 7081 4918 7101 4938
rect 12919 5089 12939 5109
rect 13027 5089 13047 5109
rect 13130 5093 13150 5113
rect 13235 5089 13255 5109
rect 13338 5093 13358 5113
rect 13448 5089 13468 5109
rect 13551 5093 13571 5113
rect 15535 5186 15555 5206
rect 15645 5182 15665 5202
rect 15748 5186 15768 5206
rect 15853 5182 15873 5202
rect 15956 5186 15976 5206
rect 16064 5186 16084 5206
rect 16167 5182 16187 5202
rect 14828 5096 14846 5114
rect 17872 5134 17892 5154
rect 17975 5130 17995 5150
rect 18083 5130 18103 5150
rect 18186 5134 18206 5154
rect 18291 5130 18311 5150
rect 18394 5134 18414 5154
rect 18504 5130 18524 5150
rect 18607 5134 18627 5154
rect 19884 5137 19902 5155
rect 7184 4914 7204 4934
rect 4568 4825 4588 4845
rect 8889 4866 8909 4886
rect 8992 4862 9012 4882
rect 9100 4862 9120 4882
rect 9203 4866 9223 4886
rect 9308 4862 9328 4882
rect 9411 4866 9431 4886
rect 9521 4862 9541 4882
rect 9624 4866 9644 4886
rect 10149 4877 10167 4895
rect 120 4773 138 4791
rect 118 4685 136 4703
rect 5176 4814 5194 4832
rect 120 4586 138 4604
rect 346 4587 366 4607
rect 449 4591 469 4611
rect 559 4587 579 4607
rect 662 4591 682 4611
rect 767 4587 787 4607
rect 870 4591 890 4611
rect 978 4591 998 4611
rect 1081 4587 1101 4607
rect 4795 4733 4813 4751
rect 5174 4726 5192 4744
rect 11424 4878 11444 4898
rect 11527 4882 11547 4902
rect 11637 4878 11657 4898
rect 11740 4882 11760 4902
rect 11845 4878 11865 4898
rect 11948 4882 11968 4902
rect 12056 4882 12076 4902
rect 12159 4878 12179 4898
rect 15205 4918 15223 4936
rect 13864 4830 13884 4850
rect 13967 4826 13987 4846
rect 14075 4826 14095 4846
rect 14178 4830 14198 4850
rect 14283 4826 14303 4846
rect 14386 4830 14406 4850
rect 14496 4826 14516 4846
rect 16480 4919 16500 4939
rect 16583 4923 16603 4943
rect 16693 4919 16713 4939
rect 16796 4923 16816 4943
rect 16901 4919 16921 4939
rect 17004 4923 17024 4943
rect 17112 4923 17132 4943
rect 17215 4919 17235 4939
rect 14599 4830 14619 4850
rect 18920 4871 18940 4891
rect 19023 4867 19043 4887
rect 19131 4867 19151 4887
rect 19234 4871 19254 4891
rect 19339 4867 19359 4887
rect 19442 4871 19462 4891
rect 19552 4867 19572 4887
rect 19655 4871 19675 4891
rect 4797 4634 4815 4652
rect 5176 4627 5194 4645
rect 5402 4628 5422 4648
rect 5505 4632 5525 4652
rect 5615 4628 5635 4648
rect 5718 4632 5738 4652
rect 5823 4628 5843 4648
rect 5926 4632 5946 4652
rect 6034 4632 6054 4652
rect 6137 4628 6157 4648
rect 9851 4774 9869 4792
rect 10151 4778 10169 4796
rect 9853 4675 9871 4693
rect 10149 4690 10167 4708
rect 15207 4819 15225 4837
rect 118 4456 136 4474
rect 2894 4515 2914 4535
rect 2997 4511 3017 4531
rect 3105 4511 3125 4531
rect 3208 4515 3228 4535
rect 3313 4511 3333 4531
rect 3416 4515 3436 4535
rect 3526 4511 3546 4531
rect 3629 4515 3649 4535
rect 120 4357 138 4375
rect 4795 4503 4813 4521
rect 5174 4497 5192 4515
rect 1284 4343 1304 4363
rect 1387 4347 1407 4367
rect 1497 4343 1517 4363
rect 1600 4347 1620 4367
rect 1705 4343 1725 4363
rect 1808 4347 1828 4367
rect 1916 4347 1936 4367
rect 2019 4343 2039 4363
rect 10151 4591 10169 4609
rect 7950 4556 7970 4576
rect 8053 4552 8073 4572
rect 8161 4552 8181 4572
rect 8264 4556 8284 4576
rect 8369 4552 8389 4572
rect 8472 4556 8492 4576
rect 8582 4552 8602 4572
rect 8685 4556 8705 4576
rect 10377 4592 10397 4612
rect 10480 4596 10500 4616
rect 10590 4592 10610 4612
rect 10693 4596 10713 4616
rect 10798 4592 10818 4612
rect 10901 4596 10921 4616
rect 11009 4596 11029 4616
rect 11112 4592 11132 4612
rect 14826 4738 14844 4756
rect 15205 4731 15223 4749
rect 14828 4639 14846 4657
rect 15207 4632 15225 4650
rect 15433 4633 15453 4653
rect 15536 4637 15556 4657
rect 15646 4633 15666 4653
rect 15749 4637 15769 4657
rect 15854 4633 15874 4653
rect 15957 4637 15977 4657
rect 16065 4637 16085 4657
rect 16168 4633 16188 4653
rect 19882 4779 19900 4797
rect 19884 4680 19902 4698
rect 4797 4404 4815 4422
rect 5176 4398 5194 4416
rect 9851 4544 9869 4562
rect 6340 4384 6360 4404
rect 6443 4388 6463 4408
rect 6553 4384 6573 4404
rect 6656 4388 6676 4408
rect 6761 4384 6781 4404
rect 6864 4388 6884 4408
rect 6972 4388 6992 4408
rect 7075 4384 7095 4404
rect 9853 4445 9871 4463
rect 10149 4461 10167 4479
rect 12925 4520 12945 4540
rect 13028 4516 13048 4536
rect 13136 4516 13156 4536
rect 13239 4520 13259 4540
rect 13344 4516 13364 4536
rect 13447 4520 13467 4540
rect 13557 4516 13577 4536
rect 13660 4520 13680 4540
rect 10151 4362 10169 4380
rect 14826 4508 14844 4526
rect 15205 4502 15223 4520
rect 118 4226 136 4244
rect 120 4127 138 4145
rect 3832 4271 3852 4291
rect 3935 4267 3955 4287
rect 4043 4267 4063 4287
rect 4146 4271 4166 4291
rect 4251 4267 4271 4287
rect 4354 4271 4374 4291
rect 4464 4267 4484 4287
rect 4567 4271 4587 4291
rect 4795 4274 4813 4292
rect 5174 4267 5192 4285
rect 4797 4175 4815 4193
rect 5176 4168 5194 4186
rect 8888 4312 8908 4332
rect 8991 4308 9011 4328
rect 9099 4308 9119 4328
rect 9202 4312 9222 4332
rect 9307 4308 9327 4328
rect 9410 4312 9430 4332
rect 9520 4308 9540 4328
rect 9623 4312 9643 4332
rect 11315 4348 11335 4368
rect 11418 4352 11438 4372
rect 11528 4348 11548 4368
rect 11631 4352 11651 4372
rect 11736 4348 11756 4368
rect 11839 4352 11859 4372
rect 11947 4352 11967 4372
rect 12050 4348 12070 4368
rect 9851 4315 9869 4333
rect 17981 4561 18001 4581
rect 18084 4557 18104 4577
rect 18192 4557 18212 4577
rect 18295 4561 18315 4581
rect 18400 4557 18420 4577
rect 18503 4561 18523 4581
rect 18613 4557 18633 4577
rect 18716 4561 18736 4581
rect 14828 4409 14846 4427
rect 15207 4403 15225 4421
rect 19882 4549 19900 4567
rect 16371 4389 16391 4409
rect 16474 4393 16494 4413
rect 16584 4389 16604 4409
rect 16687 4393 16707 4413
rect 16792 4389 16812 4409
rect 16895 4393 16915 4413
rect 17003 4393 17023 4413
rect 17106 4389 17126 4409
rect 19884 4450 19902 4468
rect 4795 4087 4813 4105
rect 9853 4216 9871 4234
rect 10149 4231 10167 4249
rect 9851 4128 9869 4146
rect 10151 4132 10169 4150
rect 13863 4276 13883 4296
rect 13966 4272 13986 4292
rect 14074 4272 14094 4292
rect 14177 4276 14197 4296
rect 14282 4272 14302 4292
rect 14385 4276 14405 4296
rect 14495 4272 14515 4292
rect 14598 4276 14618 4296
rect 14826 4279 14844 4297
rect 15205 4272 15223 4290
rect 5401 4074 5421 4094
rect 345 4033 365 4053
rect 448 4037 468 4057
rect 558 4033 578 4053
rect 661 4037 681 4057
rect 766 4033 786 4053
rect 869 4037 889 4057
rect 977 4037 997 4057
rect 1080 4033 1100 4053
rect 2754 4004 2774 4024
rect 2857 4000 2877 4020
rect 2965 4000 2985 4020
rect 3068 4004 3088 4024
rect 3173 4000 3193 4020
rect 3276 4004 3296 4024
rect 3386 4000 3406 4020
rect 3489 4004 3509 4024
rect 5504 4078 5524 4098
rect 5614 4074 5634 4094
rect 5717 4078 5737 4098
rect 5822 4074 5842 4094
rect 5925 4078 5945 4098
rect 6033 4078 6053 4098
rect 6136 4074 6156 4094
rect 7810 4045 7830 4065
rect 7913 4041 7933 4061
rect 8021 4041 8041 4061
rect 8124 4045 8144 4065
rect 8229 4041 8249 4061
rect 8332 4045 8352 4065
rect 8442 4041 8462 4061
rect 8545 4045 8565 4065
rect 14828 4180 14846 4198
rect 15207 4173 15225 4191
rect 18919 4317 18939 4337
rect 19022 4313 19042 4333
rect 19130 4313 19150 4333
rect 19233 4317 19253 4337
rect 19338 4313 19358 4333
rect 19441 4317 19461 4337
rect 19551 4313 19571 4333
rect 19654 4317 19674 4337
rect 19882 4320 19900 4338
rect 14826 4092 14844 4110
rect 19884 4221 19902 4239
rect 19882 4133 19900 4151
rect 15432 4079 15452 4099
rect 4797 3988 4815 4006
rect 119 3769 137 3787
rect 9853 4029 9871 4047
rect 10376 4038 10396 4058
rect 10479 4042 10499 4062
rect 10589 4038 10609 4058
rect 10692 4042 10712 4062
rect 10797 4038 10817 4058
rect 10900 4042 10920 4062
rect 11008 4042 11028 4062
rect 11111 4038 11131 4058
rect 12785 4009 12805 4029
rect 12888 4005 12908 4025
rect 12996 4005 13016 4025
rect 13099 4009 13119 4029
rect 13204 4005 13224 4025
rect 13307 4009 13327 4029
rect 13417 4005 13437 4025
rect 13520 4009 13540 4029
rect 15535 4083 15555 4103
rect 15645 4079 15665 4099
rect 15748 4083 15768 4103
rect 15853 4079 15873 4099
rect 15956 4083 15976 4103
rect 16064 4083 16084 4103
rect 16167 4079 16187 4099
rect 17841 4050 17861 4070
rect 17944 4046 17964 4066
rect 18052 4046 18072 4066
rect 18155 4050 18175 4070
rect 18260 4046 18280 4066
rect 18363 4050 18383 4070
rect 18473 4046 18493 4066
rect 18576 4050 18596 4070
rect 5175 3810 5193 3828
rect 14828 3993 14846 4011
rect 1425 3751 1445 3771
rect 1528 3755 1548 3775
rect 1638 3751 1658 3771
rect 1741 3755 1761 3775
rect 1846 3751 1866 3771
rect 1949 3755 1969 3775
rect 2057 3755 2077 3775
rect 2160 3751 2180 3771
rect 3834 3722 3854 3742
rect 3937 3718 3957 3738
rect 4045 3718 4065 3738
rect 4148 3722 4168 3742
rect 4253 3718 4273 3738
rect 4356 3722 4376 3742
rect 4466 3718 4486 3738
rect 6481 3792 6501 3812
rect 6584 3796 6604 3816
rect 6694 3792 6714 3812
rect 6797 3796 6817 3816
rect 6902 3792 6922 3812
rect 7005 3796 7025 3816
rect 7113 3796 7133 3816
rect 7216 3792 7236 3812
rect 8890 3763 8910 3783
rect 8993 3759 9013 3779
rect 9101 3759 9121 3779
rect 9204 3763 9224 3783
rect 9309 3759 9329 3779
rect 9412 3763 9432 3783
rect 9522 3759 9542 3779
rect 9625 3763 9645 3783
rect 10150 3774 10168 3792
rect 19884 4034 19902 4052
rect 15206 3815 15224 3833
rect 4569 3722 4589 3742
rect 121 3670 139 3688
rect 119 3582 137 3600
rect 5177 3711 5195 3729
rect 121 3483 139 3501
rect 347 3484 367 3504
rect 450 3488 470 3508
rect 560 3484 580 3504
rect 663 3488 683 3508
rect 768 3484 788 3504
rect 871 3488 891 3508
rect 979 3488 999 3508
rect 1082 3484 1102 3504
rect 4796 3630 4814 3648
rect 5175 3623 5193 3641
rect 11456 3756 11476 3776
rect 11559 3760 11579 3780
rect 11669 3756 11689 3776
rect 11772 3760 11792 3780
rect 11877 3756 11897 3776
rect 11980 3760 12000 3780
rect 12088 3760 12108 3780
rect 12191 3756 12211 3776
rect 13865 3727 13885 3747
rect 13968 3723 13988 3743
rect 14076 3723 14096 3743
rect 14179 3727 14199 3747
rect 14284 3723 14304 3743
rect 14387 3727 14407 3747
rect 14497 3723 14517 3743
rect 16512 3797 16532 3817
rect 16615 3801 16635 3821
rect 16725 3797 16745 3817
rect 16828 3801 16848 3821
rect 16933 3797 16953 3817
rect 17036 3801 17056 3821
rect 17144 3801 17164 3821
rect 17247 3797 17267 3817
rect 18921 3768 18941 3788
rect 19024 3764 19044 3784
rect 19132 3764 19152 3784
rect 19235 3768 19255 3788
rect 19340 3764 19360 3784
rect 19443 3768 19463 3788
rect 19553 3764 19573 3784
rect 19656 3768 19676 3788
rect 14600 3727 14620 3747
rect 4798 3531 4816 3549
rect 5177 3524 5195 3542
rect 5403 3525 5423 3545
rect 5506 3529 5526 3549
rect 5616 3525 5636 3545
rect 5719 3529 5739 3549
rect 5824 3525 5844 3545
rect 5927 3529 5947 3549
rect 6035 3529 6055 3549
rect 6138 3525 6158 3545
rect 9852 3671 9870 3689
rect 10152 3675 10170 3693
rect 9854 3572 9872 3590
rect 10150 3587 10168 3605
rect 15208 3716 15226 3734
rect 119 3353 137 3371
rect 2895 3412 2915 3432
rect 2998 3408 3018 3428
rect 3106 3408 3126 3428
rect 3209 3412 3229 3432
rect 3314 3408 3334 3428
rect 3417 3412 3437 3432
rect 3527 3408 3547 3428
rect 3630 3412 3650 3432
rect 121 3254 139 3272
rect 4796 3400 4814 3418
rect 5175 3394 5193 3412
rect 1285 3240 1305 3260
rect 1388 3244 1408 3264
rect 1498 3240 1518 3260
rect 1601 3244 1621 3264
rect 1706 3240 1726 3260
rect 1809 3244 1829 3264
rect 1917 3244 1937 3264
rect 2020 3240 2040 3260
rect 10152 3488 10170 3506
rect 7951 3453 7971 3473
rect 8054 3449 8074 3469
rect 8162 3449 8182 3469
rect 8265 3453 8285 3473
rect 8370 3449 8390 3469
rect 8473 3453 8493 3473
rect 8583 3449 8603 3469
rect 8686 3453 8706 3473
rect 10378 3489 10398 3509
rect 10481 3493 10501 3513
rect 10591 3489 10611 3509
rect 10694 3493 10714 3513
rect 10799 3489 10819 3509
rect 10902 3493 10922 3513
rect 11010 3493 11030 3513
rect 11113 3489 11133 3509
rect 14827 3635 14845 3653
rect 15206 3628 15224 3646
rect 14829 3536 14847 3554
rect 15208 3529 15226 3547
rect 15434 3530 15454 3550
rect 15537 3534 15557 3554
rect 15647 3530 15667 3550
rect 15750 3534 15770 3554
rect 15855 3530 15875 3550
rect 15958 3534 15978 3554
rect 16066 3534 16086 3554
rect 16169 3530 16189 3550
rect 19883 3676 19901 3694
rect 19885 3577 19903 3595
rect 4798 3301 4816 3319
rect 5177 3295 5195 3313
rect 9852 3441 9870 3459
rect 6341 3281 6361 3301
rect 6444 3285 6464 3305
rect 6554 3281 6574 3301
rect 6657 3285 6677 3305
rect 6762 3281 6782 3301
rect 6865 3285 6885 3305
rect 6973 3285 6993 3305
rect 7076 3281 7096 3301
rect 9854 3342 9872 3360
rect 10150 3358 10168 3376
rect 12926 3417 12946 3437
rect 13029 3413 13049 3433
rect 13137 3413 13157 3433
rect 13240 3417 13260 3437
rect 13345 3413 13365 3433
rect 13448 3417 13468 3437
rect 13558 3413 13578 3433
rect 13661 3417 13681 3437
rect 10152 3259 10170 3277
rect 14827 3405 14845 3423
rect 15206 3399 15224 3417
rect 119 3123 137 3141
rect 121 3024 139 3042
rect 3833 3168 3853 3188
rect 3936 3164 3956 3184
rect 4044 3164 4064 3184
rect 4147 3168 4167 3188
rect 4252 3164 4272 3184
rect 4355 3168 4375 3188
rect 4465 3164 4485 3184
rect 4568 3168 4588 3188
rect 4796 3171 4814 3189
rect 5175 3164 5193 3182
rect 4798 3072 4816 3090
rect 5177 3065 5195 3083
rect 8889 3209 8909 3229
rect 8992 3205 9012 3225
rect 9100 3205 9120 3225
rect 9203 3209 9223 3229
rect 9308 3205 9328 3225
rect 9411 3209 9431 3229
rect 9521 3205 9541 3225
rect 9624 3209 9644 3229
rect 11316 3245 11336 3265
rect 11419 3249 11439 3269
rect 11529 3245 11549 3265
rect 11632 3249 11652 3269
rect 11737 3245 11757 3265
rect 11840 3249 11860 3269
rect 11948 3249 11968 3269
rect 12051 3245 12071 3265
rect 9852 3212 9870 3230
rect 17982 3458 18002 3478
rect 18085 3454 18105 3474
rect 18193 3454 18213 3474
rect 18296 3458 18316 3478
rect 18401 3454 18421 3474
rect 18504 3458 18524 3478
rect 18614 3454 18634 3474
rect 18717 3458 18737 3478
rect 14829 3306 14847 3324
rect 15208 3300 15226 3318
rect 19883 3446 19901 3464
rect 16372 3286 16392 3306
rect 16475 3290 16495 3310
rect 16585 3286 16605 3306
rect 16688 3290 16708 3310
rect 16793 3286 16813 3306
rect 16896 3290 16916 3310
rect 17004 3290 17024 3310
rect 17107 3286 17127 3306
rect 19885 3347 19903 3365
rect 4796 2984 4814 3002
rect 9854 3113 9872 3131
rect 10150 3128 10168 3146
rect 9852 3025 9870 3043
rect 10152 3029 10170 3047
rect 13864 3173 13884 3193
rect 13967 3169 13987 3189
rect 14075 3169 14095 3189
rect 14178 3173 14198 3193
rect 14283 3169 14303 3189
rect 14386 3173 14406 3193
rect 14496 3169 14516 3189
rect 14599 3173 14619 3193
rect 14827 3176 14845 3194
rect 15206 3169 15224 3187
rect 5402 2971 5422 2991
rect 346 2930 366 2950
rect 449 2934 469 2954
rect 559 2930 579 2950
rect 662 2934 682 2954
rect 767 2930 787 2950
rect 870 2934 890 2954
rect 978 2934 998 2954
rect 1081 2930 1101 2950
rect 2785 2888 2805 2908
rect 2888 2884 2908 2904
rect 2996 2884 3016 2904
rect 3099 2888 3119 2908
rect 3204 2884 3224 2904
rect 3307 2888 3327 2908
rect 3417 2884 3437 2904
rect 3520 2888 3540 2908
rect 5505 2975 5525 2995
rect 5615 2971 5635 2991
rect 5718 2975 5738 2995
rect 5823 2971 5843 2991
rect 5926 2975 5946 2995
rect 6034 2975 6054 2995
rect 6137 2971 6157 2991
rect 7841 2929 7861 2949
rect 4798 2885 4816 2903
rect 7944 2925 7964 2945
rect 8052 2925 8072 2945
rect 8155 2929 8175 2949
rect 8260 2925 8280 2945
rect 8363 2929 8383 2949
rect 8473 2925 8493 2945
rect 8576 2929 8596 2949
rect 14829 3077 14847 3095
rect 15208 3070 15226 3088
rect 18920 3214 18940 3234
rect 19023 3210 19043 3230
rect 19131 3210 19151 3230
rect 19234 3214 19254 3234
rect 19339 3210 19359 3230
rect 19442 3214 19462 3234
rect 19552 3210 19572 3230
rect 19655 3214 19675 3234
rect 19883 3217 19901 3235
rect 14827 2989 14845 3007
rect 19885 3118 19903 3136
rect 19883 3030 19901 3048
rect 15433 2976 15453 2996
rect 9854 2926 9872 2944
rect 10377 2935 10397 2955
rect 10480 2939 10500 2959
rect 10590 2935 10610 2955
rect 10693 2939 10713 2959
rect 10798 2935 10818 2955
rect 10901 2939 10921 2959
rect 11009 2939 11029 2959
rect 11112 2935 11132 2955
rect 12816 2893 12836 2913
rect 12919 2889 12939 2909
rect 13027 2889 13047 2909
rect 13130 2893 13150 2913
rect 13235 2889 13255 2909
rect 13338 2893 13358 2913
rect 13448 2889 13468 2909
rect 13551 2893 13571 2913
rect 15536 2980 15556 3000
rect 15646 2976 15666 2996
rect 15749 2980 15769 3000
rect 15854 2976 15874 2996
rect 15957 2980 15977 3000
rect 16065 2980 16085 3000
rect 16168 2976 16188 2996
rect 17872 2934 17892 2954
rect 14829 2890 14847 2908
rect 17975 2930 17995 2950
rect 18083 2930 18103 2950
rect 18186 2934 18206 2954
rect 18291 2930 18311 2950
rect 18394 2934 18414 2954
rect 18504 2930 18524 2950
rect 18607 2934 18627 2954
rect 19885 2931 19903 2949
rect 119 2666 137 2684
rect 1395 2661 1415 2681
rect 1498 2665 1518 2685
rect 1608 2661 1628 2681
rect 1711 2665 1731 2685
rect 1816 2661 1836 2681
rect 1919 2665 1939 2685
rect 2027 2665 2047 2685
rect 5175 2707 5193 2725
rect 2130 2661 2150 2681
rect 3834 2619 3854 2639
rect 3937 2615 3957 2635
rect 4045 2615 4065 2635
rect 4148 2619 4168 2639
rect 4253 2615 4273 2635
rect 4356 2619 4376 2639
rect 4466 2615 4486 2635
rect 6451 2702 6471 2722
rect 6554 2706 6574 2726
rect 6664 2702 6684 2722
rect 6767 2706 6787 2726
rect 6872 2702 6892 2722
rect 6975 2706 6995 2726
rect 7083 2706 7103 2726
rect 7186 2702 7206 2722
rect 8890 2660 8910 2680
rect 8993 2656 9013 2676
rect 9101 2656 9121 2676
rect 9204 2660 9224 2680
rect 9309 2656 9329 2676
rect 9412 2660 9432 2680
rect 9522 2656 9542 2676
rect 9625 2660 9645 2680
rect 10150 2671 10168 2689
rect 4569 2619 4589 2639
rect 121 2567 139 2585
rect 119 2479 137 2497
rect 5177 2608 5195 2626
rect 121 2380 139 2398
rect 347 2381 367 2401
rect 450 2385 470 2405
rect 560 2381 580 2401
rect 663 2385 683 2405
rect 768 2381 788 2401
rect 871 2385 891 2405
rect 979 2385 999 2405
rect 1082 2381 1102 2401
rect 4796 2527 4814 2545
rect 5175 2520 5193 2538
rect 11426 2666 11446 2686
rect 11529 2670 11549 2690
rect 11639 2666 11659 2686
rect 11742 2670 11762 2690
rect 11847 2666 11867 2686
rect 11950 2670 11970 2690
rect 12058 2670 12078 2690
rect 15206 2712 15224 2730
rect 12161 2666 12181 2686
rect 13865 2624 13885 2644
rect 13968 2620 13988 2640
rect 14076 2620 14096 2640
rect 14179 2624 14199 2644
rect 14284 2620 14304 2640
rect 14387 2624 14407 2644
rect 14497 2620 14517 2640
rect 16482 2707 16502 2727
rect 16585 2711 16605 2731
rect 16695 2707 16715 2727
rect 16798 2711 16818 2731
rect 16903 2707 16923 2727
rect 17006 2711 17026 2731
rect 17114 2711 17134 2731
rect 17217 2707 17237 2727
rect 18921 2665 18941 2685
rect 19024 2661 19044 2681
rect 19132 2661 19152 2681
rect 19235 2665 19255 2685
rect 19340 2661 19360 2681
rect 19443 2665 19463 2685
rect 19553 2661 19573 2681
rect 19656 2665 19676 2685
rect 14600 2624 14620 2644
rect 4798 2428 4816 2446
rect 5177 2421 5195 2439
rect 5403 2422 5423 2442
rect 5506 2426 5526 2446
rect 5616 2422 5636 2442
rect 5719 2426 5739 2446
rect 5824 2422 5844 2442
rect 5927 2426 5947 2446
rect 6035 2426 6055 2446
rect 6138 2422 6158 2442
rect 9852 2568 9870 2586
rect 10152 2572 10170 2590
rect 9854 2469 9872 2487
rect 10150 2484 10168 2502
rect 15208 2613 15226 2631
rect 119 2250 137 2268
rect 2895 2309 2915 2329
rect 2998 2305 3018 2325
rect 3106 2305 3126 2325
rect 3209 2309 3229 2329
rect 3314 2305 3334 2325
rect 3417 2309 3437 2329
rect 3527 2305 3547 2325
rect 3630 2309 3650 2329
rect 121 2151 139 2169
rect 4796 2297 4814 2315
rect 5175 2291 5193 2309
rect 1285 2137 1305 2157
rect 1388 2141 1408 2161
rect 1498 2137 1518 2157
rect 1601 2141 1621 2161
rect 1706 2137 1726 2157
rect 1809 2141 1829 2161
rect 1917 2141 1937 2161
rect 2020 2137 2040 2157
rect 10152 2385 10170 2403
rect 7951 2350 7971 2370
rect 8054 2346 8074 2366
rect 8162 2346 8182 2366
rect 8265 2350 8285 2370
rect 8370 2346 8390 2366
rect 8473 2350 8493 2370
rect 8583 2346 8603 2366
rect 8686 2350 8706 2370
rect 10378 2386 10398 2406
rect 10481 2390 10501 2410
rect 10591 2386 10611 2406
rect 10694 2390 10714 2410
rect 10799 2386 10819 2406
rect 10902 2390 10922 2410
rect 11010 2390 11030 2410
rect 11113 2386 11133 2406
rect 14827 2532 14845 2550
rect 15206 2525 15224 2543
rect 14829 2433 14847 2451
rect 15208 2426 15226 2444
rect 15434 2427 15454 2447
rect 15537 2431 15557 2451
rect 15647 2427 15667 2447
rect 15750 2431 15770 2451
rect 15855 2427 15875 2447
rect 15958 2431 15978 2451
rect 16066 2431 16086 2451
rect 16169 2427 16189 2447
rect 19883 2573 19901 2591
rect 19885 2474 19903 2492
rect 4798 2198 4816 2216
rect 5177 2192 5195 2210
rect 9852 2338 9870 2356
rect 6341 2178 6361 2198
rect 6444 2182 6464 2202
rect 6554 2178 6574 2198
rect 6657 2182 6677 2202
rect 6762 2178 6782 2198
rect 6865 2182 6885 2202
rect 6973 2182 6993 2202
rect 7076 2178 7096 2198
rect 9854 2239 9872 2257
rect 10150 2255 10168 2273
rect 12926 2314 12946 2334
rect 13029 2310 13049 2330
rect 13137 2310 13157 2330
rect 13240 2314 13260 2334
rect 13345 2310 13365 2330
rect 13448 2314 13468 2334
rect 13558 2310 13578 2330
rect 13661 2314 13681 2334
rect 10152 2156 10170 2174
rect 14827 2302 14845 2320
rect 15206 2296 15224 2314
rect 119 2020 137 2038
rect 121 1921 139 1939
rect 3833 2065 3853 2085
rect 3936 2061 3956 2081
rect 4044 2061 4064 2081
rect 4147 2065 4167 2085
rect 4252 2061 4272 2081
rect 4355 2065 4375 2085
rect 4465 2061 4485 2081
rect 4568 2065 4588 2085
rect 4796 2068 4814 2086
rect 5175 2061 5193 2079
rect 4798 1969 4816 1987
rect 5177 1962 5195 1980
rect 8889 2106 8909 2126
rect 8992 2102 9012 2122
rect 9100 2102 9120 2122
rect 9203 2106 9223 2126
rect 9308 2102 9328 2122
rect 9411 2106 9431 2126
rect 9521 2102 9541 2122
rect 9624 2106 9644 2126
rect 11316 2142 11336 2162
rect 11419 2146 11439 2166
rect 11529 2142 11549 2162
rect 11632 2146 11652 2166
rect 11737 2142 11757 2162
rect 11840 2146 11860 2166
rect 11948 2146 11968 2166
rect 12051 2142 12071 2162
rect 9852 2109 9870 2127
rect 17982 2355 18002 2375
rect 18085 2351 18105 2371
rect 18193 2351 18213 2371
rect 18296 2355 18316 2375
rect 18401 2351 18421 2371
rect 18504 2355 18524 2375
rect 18614 2351 18634 2371
rect 18717 2355 18737 2375
rect 14829 2203 14847 2221
rect 15208 2197 15226 2215
rect 19883 2343 19901 2361
rect 16372 2183 16392 2203
rect 16475 2187 16495 2207
rect 16585 2183 16605 2203
rect 16688 2187 16708 2207
rect 16793 2183 16813 2203
rect 16896 2187 16916 2207
rect 17004 2187 17024 2207
rect 17107 2183 17127 2203
rect 19885 2244 19903 2262
rect 4796 1881 4814 1899
rect 9854 2010 9872 2028
rect 10150 2025 10168 2043
rect 9852 1922 9870 1940
rect 10152 1926 10170 1944
rect 13864 2070 13884 2090
rect 13967 2066 13987 2086
rect 14075 2066 14095 2086
rect 14178 2070 14198 2090
rect 14283 2066 14303 2086
rect 14386 2070 14406 2090
rect 14496 2066 14516 2086
rect 14599 2070 14619 2090
rect 14827 2073 14845 2091
rect 15206 2066 15224 2084
rect 5402 1868 5422 1888
rect 346 1827 366 1847
rect 449 1831 469 1851
rect 559 1827 579 1847
rect 662 1831 682 1851
rect 767 1827 787 1847
rect 870 1831 890 1851
rect 978 1831 998 1851
rect 1081 1827 1101 1847
rect 2755 1798 2775 1818
rect 2858 1794 2878 1814
rect 2966 1794 2986 1814
rect 3069 1798 3089 1818
rect 3174 1794 3194 1814
rect 3277 1798 3297 1818
rect 3387 1794 3407 1814
rect 3490 1798 3510 1818
rect 5505 1872 5525 1892
rect 5615 1868 5635 1888
rect 5718 1872 5738 1892
rect 5823 1868 5843 1888
rect 5926 1872 5946 1892
rect 6034 1872 6054 1892
rect 6137 1868 6157 1888
rect 7811 1839 7831 1859
rect 7914 1835 7934 1855
rect 8022 1835 8042 1855
rect 8125 1839 8145 1859
rect 8230 1835 8250 1855
rect 8333 1839 8353 1859
rect 8443 1835 8463 1855
rect 8546 1839 8566 1859
rect 14829 1974 14847 1992
rect 15208 1967 15226 1985
rect 18920 2111 18940 2131
rect 19023 2107 19043 2127
rect 19131 2107 19151 2127
rect 19234 2111 19254 2131
rect 19339 2107 19359 2127
rect 19442 2111 19462 2131
rect 19552 2107 19572 2127
rect 19655 2111 19675 2131
rect 19883 2114 19901 2132
rect 14827 1886 14845 1904
rect 19885 2015 19903 2033
rect 19883 1927 19901 1945
rect 15433 1873 15453 1893
rect 4798 1782 4816 1800
rect 120 1563 138 1581
rect 9854 1823 9872 1841
rect 10377 1832 10397 1852
rect 10480 1836 10500 1856
rect 10590 1832 10610 1852
rect 10693 1836 10713 1856
rect 10798 1832 10818 1852
rect 10901 1836 10921 1856
rect 11009 1836 11029 1856
rect 11112 1832 11132 1852
rect 12786 1803 12806 1823
rect 12889 1799 12909 1819
rect 12997 1799 13017 1819
rect 13100 1803 13120 1823
rect 13205 1799 13225 1819
rect 13308 1803 13328 1823
rect 13418 1799 13438 1819
rect 13521 1803 13541 1823
rect 15536 1877 15556 1897
rect 15646 1873 15666 1893
rect 15749 1877 15769 1897
rect 15854 1873 15874 1893
rect 15957 1877 15977 1897
rect 16065 1877 16085 1897
rect 16168 1873 16188 1893
rect 17842 1844 17862 1864
rect 17945 1840 17965 1860
rect 18053 1840 18073 1860
rect 18156 1844 18176 1864
rect 18261 1840 18281 1860
rect 18364 1844 18384 1864
rect 18474 1840 18494 1860
rect 18577 1844 18597 1864
rect 5176 1604 5194 1622
rect 14829 1787 14847 1805
rect 1426 1545 1446 1565
rect 1529 1549 1549 1569
rect 1639 1545 1659 1565
rect 1742 1549 1762 1569
rect 1847 1545 1867 1565
rect 1950 1549 1970 1569
rect 2058 1549 2078 1569
rect 2161 1545 2181 1565
rect 3835 1516 3855 1536
rect 3938 1512 3958 1532
rect 4046 1512 4066 1532
rect 4149 1516 4169 1536
rect 4254 1512 4274 1532
rect 4357 1516 4377 1536
rect 4467 1512 4487 1532
rect 6482 1586 6502 1606
rect 6585 1590 6605 1610
rect 6695 1586 6715 1606
rect 6798 1590 6818 1610
rect 6903 1586 6923 1606
rect 7006 1590 7026 1610
rect 7114 1590 7134 1610
rect 7217 1586 7237 1606
rect 8891 1557 8911 1577
rect 8994 1553 9014 1573
rect 9102 1553 9122 1573
rect 9205 1557 9225 1577
rect 9310 1553 9330 1573
rect 9413 1557 9433 1577
rect 9523 1553 9543 1573
rect 9626 1557 9646 1577
rect 10151 1568 10169 1586
rect 19885 1828 19903 1846
rect 15207 1609 15225 1627
rect 4570 1516 4590 1536
rect 122 1464 140 1482
rect 120 1376 138 1394
rect 5178 1505 5196 1523
rect 122 1277 140 1295
rect 348 1278 368 1298
rect 451 1282 471 1302
rect 561 1278 581 1298
rect 664 1282 684 1302
rect 769 1278 789 1298
rect 872 1282 892 1302
rect 980 1282 1000 1302
rect 1083 1278 1103 1298
rect 4797 1424 4815 1442
rect 5176 1417 5194 1435
rect 11457 1550 11477 1570
rect 11560 1554 11580 1574
rect 11670 1550 11690 1570
rect 11773 1554 11793 1574
rect 11878 1550 11898 1570
rect 11981 1554 12001 1574
rect 12089 1554 12109 1574
rect 12192 1550 12212 1570
rect 13866 1521 13886 1541
rect 13969 1517 13989 1537
rect 14077 1517 14097 1537
rect 14180 1521 14200 1541
rect 14285 1517 14305 1537
rect 14388 1521 14408 1541
rect 14498 1517 14518 1537
rect 16513 1591 16533 1611
rect 16616 1595 16636 1615
rect 16726 1591 16746 1611
rect 16829 1595 16849 1615
rect 16934 1591 16954 1611
rect 17037 1595 17057 1615
rect 17145 1595 17165 1615
rect 17248 1591 17268 1611
rect 18922 1562 18942 1582
rect 19025 1558 19045 1578
rect 19133 1558 19153 1578
rect 19236 1562 19256 1582
rect 19341 1558 19361 1578
rect 19444 1562 19464 1582
rect 19554 1558 19574 1578
rect 19657 1562 19677 1582
rect 14601 1521 14621 1541
rect 4799 1325 4817 1343
rect 5178 1318 5196 1336
rect 5404 1319 5424 1339
rect 5507 1323 5527 1343
rect 5617 1319 5637 1339
rect 5720 1323 5740 1343
rect 5825 1319 5845 1339
rect 5928 1323 5948 1343
rect 6036 1323 6056 1343
rect 6139 1319 6159 1339
rect 9853 1465 9871 1483
rect 10153 1469 10171 1487
rect 9855 1366 9873 1384
rect 10151 1381 10169 1399
rect 15209 1510 15227 1528
rect 120 1147 138 1165
rect 2896 1206 2916 1226
rect 2999 1202 3019 1222
rect 3107 1202 3127 1222
rect 3210 1206 3230 1226
rect 3315 1202 3335 1222
rect 3418 1206 3438 1226
rect 3528 1202 3548 1222
rect 3631 1206 3651 1226
rect 122 1048 140 1066
rect 4797 1194 4815 1212
rect 5176 1188 5194 1206
rect 1286 1034 1306 1054
rect 1389 1038 1409 1058
rect 1499 1034 1519 1054
rect 1602 1038 1622 1058
rect 1707 1034 1727 1054
rect 1810 1038 1830 1058
rect 1918 1038 1938 1058
rect 2021 1034 2041 1054
rect 10153 1282 10171 1300
rect 7952 1247 7972 1267
rect 8055 1243 8075 1263
rect 8163 1243 8183 1263
rect 8266 1247 8286 1267
rect 8371 1243 8391 1263
rect 8474 1247 8494 1267
rect 8584 1243 8604 1263
rect 8687 1247 8707 1267
rect 10379 1283 10399 1303
rect 10482 1287 10502 1307
rect 10592 1283 10612 1303
rect 10695 1287 10715 1307
rect 10800 1283 10820 1303
rect 10903 1287 10923 1307
rect 11011 1287 11031 1307
rect 11114 1283 11134 1303
rect 14828 1429 14846 1447
rect 15207 1422 15225 1440
rect 14830 1330 14848 1348
rect 15209 1323 15227 1341
rect 15435 1324 15455 1344
rect 15538 1328 15558 1348
rect 15648 1324 15668 1344
rect 15751 1328 15771 1348
rect 15856 1324 15876 1344
rect 15959 1328 15979 1348
rect 16067 1328 16087 1348
rect 16170 1324 16190 1344
rect 19884 1470 19902 1488
rect 19886 1371 19904 1389
rect 4799 1095 4817 1113
rect 5178 1089 5196 1107
rect 9853 1235 9871 1253
rect 6342 1075 6362 1095
rect 6445 1079 6465 1099
rect 6555 1075 6575 1095
rect 6658 1079 6678 1099
rect 6763 1075 6783 1095
rect 6866 1079 6886 1099
rect 6974 1079 6994 1099
rect 7077 1075 7097 1095
rect 9855 1136 9873 1154
rect 10151 1152 10169 1170
rect 12927 1211 12947 1231
rect 13030 1207 13050 1227
rect 13138 1207 13158 1227
rect 13241 1211 13261 1231
rect 13346 1207 13366 1227
rect 13449 1211 13469 1231
rect 13559 1207 13579 1227
rect 13662 1211 13682 1231
rect 10153 1053 10171 1071
rect 14828 1199 14846 1217
rect 15207 1193 15225 1211
rect 120 917 138 935
rect 122 818 140 836
rect 3834 962 3854 982
rect 3937 958 3957 978
rect 4045 958 4065 978
rect 4148 962 4168 982
rect 4253 958 4273 978
rect 4356 962 4376 982
rect 4466 958 4486 978
rect 4569 962 4589 982
rect 4797 965 4815 983
rect 5176 958 5194 976
rect 4799 866 4817 884
rect 5178 859 5196 877
rect 8890 1003 8910 1023
rect 8993 999 9013 1019
rect 9101 999 9121 1019
rect 9204 1003 9224 1023
rect 9309 999 9329 1019
rect 9412 1003 9432 1023
rect 9522 999 9542 1019
rect 9625 1003 9645 1023
rect 11317 1039 11337 1059
rect 11420 1043 11440 1063
rect 11530 1039 11550 1059
rect 11633 1043 11653 1063
rect 11738 1039 11758 1059
rect 11841 1043 11861 1063
rect 11949 1043 11969 1063
rect 12052 1039 12072 1059
rect 9853 1006 9871 1024
rect 17983 1252 18003 1272
rect 18086 1248 18106 1268
rect 18194 1248 18214 1268
rect 18297 1252 18317 1272
rect 18402 1248 18422 1268
rect 18505 1252 18525 1272
rect 18615 1248 18635 1268
rect 18718 1252 18738 1272
rect 14830 1100 14848 1118
rect 15209 1094 15227 1112
rect 19884 1240 19902 1258
rect 16373 1080 16393 1100
rect 16476 1084 16496 1104
rect 16586 1080 16606 1100
rect 16689 1084 16709 1104
rect 16794 1080 16814 1100
rect 16897 1084 16917 1104
rect 17005 1084 17025 1104
rect 17108 1080 17128 1100
rect 19886 1141 19904 1159
rect 4797 778 4815 796
rect 9855 907 9873 925
rect 10151 922 10169 940
rect 9853 819 9871 837
rect 10153 823 10171 841
rect 13865 967 13885 987
rect 13968 963 13988 983
rect 14076 963 14096 983
rect 14179 967 14199 987
rect 14284 963 14304 983
rect 14387 967 14407 987
rect 14497 963 14517 983
rect 14600 967 14620 987
rect 14828 970 14846 988
rect 15207 963 15225 981
rect 5403 765 5423 785
rect 347 724 367 744
rect 450 728 470 748
rect 560 724 580 744
rect 663 728 683 748
rect 768 724 788 744
rect 871 728 891 748
rect 979 728 999 748
rect 1082 724 1102 744
rect 5506 769 5526 789
rect 5616 765 5636 785
rect 5719 769 5739 789
rect 5824 765 5844 785
rect 5927 769 5947 789
rect 6035 769 6055 789
rect 6138 765 6158 785
rect 14830 871 14848 889
rect 15209 864 15227 882
rect 18921 1008 18941 1028
rect 19024 1004 19044 1024
rect 19132 1004 19152 1024
rect 19235 1008 19255 1028
rect 19340 1004 19360 1024
rect 19443 1008 19463 1028
rect 19553 1004 19573 1024
rect 19656 1008 19676 1028
rect 19884 1011 19902 1029
rect 14828 783 14846 801
rect 19886 912 19904 930
rect 19884 824 19902 842
rect 15434 770 15454 790
rect 9855 720 9873 738
rect 10378 729 10398 749
rect 4799 679 4817 697
rect 10481 733 10501 753
rect 10591 729 10611 749
rect 10694 733 10714 753
rect 10799 729 10819 749
rect 10902 733 10922 753
rect 11010 733 11030 753
rect 11113 729 11133 749
rect 15537 774 15557 794
rect 15647 770 15667 790
rect 15750 774 15770 794
rect 15855 770 15875 790
rect 15958 774 15978 794
rect 16066 774 16086 794
rect 16169 770 16189 790
rect 19886 725 19904 743
rect 14830 684 14848 702
rect 1594 165 1614 185
rect 1697 169 1717 189
rect 1807 165 1827 185
rect 1910 169 1930 189
rect 2015 165 2035 185
rect 2118 169 2138 189
rect 2226 169 2246 189
rect 2329 165 2349 185
rect 6650 206 6670 226
rect 6753 210 6773 230
rect 6863 206 6883 226
rect 6966 210 6986 230
rect 7071 206 7091 226
rect 7174 210 7194 230
rect 7282 210 7302 230
rect 7385 206 7405 226
rect 4544 145 4564 165
rect 4647 149 4667 169
rect 4757 145 4777 165
rect 4860 149 4880 169
rect 4965 145 4985 165
rect 5068 149 5088 169
rect 5176 149 5196 169
rect 5279 145 5299 165
rect 11625 170 11645 190
rect 11728 174 11748 194
rect 11838 170 11858 190
rect 11941 174 11961 194
rect 12046 170 12066 190
rect 12149 174 12169 194
rect 12257 174 12277 194
rect 12360 170 12380 190
rect 16681 211 16701 231
rect 16784 215 16804 235
rect 16894 211 16914 231
rect 16997 215 17017 235
rect 17102 211 17122 231
rect 17205 215 17225 235
rect 17313 215 17333 235
rect 17416 211 17436 231
rect 14575 150 14595 170
rect 14678 154 14698 174
rect 14788 150 14808 170
rect 14891 154 14911 174
rect 14996 150 15016 170
rect 15099 154 15119 174
rect 15207 154 15227 174
rect 15310 150 15330 170
rect 9478 29 9498 49
rect 9581 33 9601 53
rect 9691 29 9711 49
rect 9794 33 9814 53
rect 9899 29 9919 49
rect 10002 33 10022 53
rect 10110 33 10130 53
rect 10213 29 10233 49
<< pdiffc >>
rect 350 9148 370 9168
rect 446 9148 466 9168
rect 563 9148 583 9168
rect 659 9148 679 9168
rect 771 9148 791 9168
rect 867 9148 887 9168
rect 977 9148 997 9168
rect 1073 9148 1093 9168
rect 5406 9189 5426 9209
rect 3837 9088 3857 9108
rect 3933 9088 3953 9108
rect 4043 9088 4063 9108
rect 4139 9088 4159 9108
rect 4251 9088 4271 9108
rect 4347 9088 4367 9108
rect 4464 9088 4484 9108
rect 5502 9189 5522 9209
rect 5619 9189 5639 9209
rect 5715 9189 5735 9209
rect 5827 9189 5847 9209
rect 5923 9189 5943 9209
rect 6033 9189 6053 9209
rect 6129 9189 6149 9209
rect 4560 9088 4580 9108
rect 8893 9129 8913 9149
rect 8989 9129 9009 9149
rect 9099 9129 9119 9149
rect 9195 9129 9215 9149
rect 9307 9129 9327 9149
rect 9403 9129 9423 9149
rect 9520 9129 9540 9149
rect 9616 9129 9636 9149
rect 10381 9153 10401 9173
rect 10477 9153 10497 9173
rect 10594 9153 10614 9173
rect 10690 9153 10710 9173
rect 10802 9153 10822 9173
rect 10898 9153 10918 9173
rect 11008 9153 11028 9173
rect 11104 9153 11124 9173
rect 15437 9194 15457 9214
rect 1288 8904 1308 8924
rect 1384 8904 1404 8924
rect 1501 8904 1521 8924
rect 1597 8904 1617 8924
rect 1709 8904 1729 8924
rect 1805 8904 1825 8924
rect 1915 8904 1935 8924
rect 2011 8904 2031 8924
rect 6344 8945 6364 8965
rect 2898 8778 2918 8798
rect 2994 8778 3014 8798
rect 3104 8778 3124 8798
rect 3200 8778 3220 8798
rect 3312 8778 3332 8798
rect 3408 8778 3428 8798
rect 3525 8778 3545 8798
rect 6440 8945 6460 8965
rect 6557 8945 6577 8965
rect 6653 8945 6673 8965
rect 6765 8945 6785 8965
rect 6861 8945 6881 8965
rect 6971 8945 6991 8965
rect 13868 9093 13888 9113
rect 7067 8945 7087 8965
rect 13964 9093 13984 9113
rect 14074 9093 14094 9113
rect 14170 9093 14190 9113
rect 14282 9093 14302 9113
rect 14378 9093 14398 9113
rect 14495 9093 14515 9113
rect 15533 9194 15553 9214
rect 15650 9194 15670 9214
rect 15746 9194 15766 9214
rect 15858 9194 15878 9214
rect 15954 9194 15974 9214
rect 16064 9194 16084 9214
rect 16160 9194 16180 9214
rect 14591 9093 14611 9113
rect 18924 9134 18944 9154
rect 19020 9134 19040 9154
rect 19130 9134 19150 9154
rect 19226 9134 19246 9154
rect 19338 9134 19358 9154
rect 19434 9134 19454 9154
rect 19551 9134 19571 9154
rect 19647 9134 19667 9154
rect 3621 8778 3641 8798
rect 7954 8819 7974 8839
rect 8050 8819 8070 8839
rect 8160 8819 8180 8839
rect 8256 8819 8276 8839
rect 8368 8819 8388 8839
rect 8464 8819 8484 8839
rect 8581 8819 8601 8839
rect 11319 8909 11339 8929
rect 8677 8819 8697 8839
rect 11415 8909 11435 8929
rect 11532 8909 11552 8929
rect 11628 8909 11648 8929
rect 11740 8909 11760 8929
rect 11836 8909 11856 8929
rect 11946 8909 11966 8929
rect 12042 8909 12062 8929
rect 16375 8950 16395 8970
rect 349 8594 369 8614
rect 445 8594 465 8614
rect 562 8594 582 8614
rect 658 8594 678 8614
rect 770 8594 790 8614
rect 866 8594 886 8614
rect 976 8594 996 8614
rect 1072 8594 1092 8614
rect 5405 8635 5425 8655
rect 3836 8534 3856 8554
rect 3932 8534 3952 8554
rect 4042 8534 4062 8554
rect 4138 8534 4158 8554
rect 4250 8534 4270 8554
rect 4346 8534 4366 8554
rect 4463 8534 4483 8554
rect 5501 8635 5521 8655
rect 5618 8635 5638 8655
rect 5714 8635 5734 8655
rect 5826 8635 5846 8655
rect 5922 8635 5942 8655
rect 6032 8635 6052 8655
rect 12929 8783 12949 8803
rect 6128 8635 6148 8655
rect 13025 8783 13045 8803
rect 13135 8783 13155 8803
rect 13231 8783 13251 8803
rect 13343 8783 13363 8803
rect 13439 8783 13459 8803
rect 13556 8783 13576 8803
rect 16471 8950 16491 8970
rect 16588 8950 16608 8970
rect 16684 8950 16704 8970
rect 16796 8950 16816 8970
rect 16892 8950 16912 8970
rect 17002 8950 17022 8970
rect 17098 8950 17118 8970
rect 13652 8783 13672 8803
rect 17985 8824 18005 8844
rect 18081 8824 18101 8844
rect 18191 8824 18211 8844
rect 18287 8824 18307 8844
rect 18399 8824 18419 8844
rect 18495 8824 18515 8844
rect 18612 8824 18632 8844
rect 18708 8824 18728 8844
rect 4559 8534 4579 8554
rect 8892 8575 8912 8595
rect 8988 8575 9008 8595
rect 9098 8575 9118 8595
rect 9194 8575 9214 8595
rect 9306 8575 9326 8595
rect 9402 8575 9422 8595
rect 9519 8575 9539 8595
rect 9615 8575 9635 8595
rect 10380 8599 10400 8619
rect 10476 8599 10496 8619
rect 10593 8599 10613 8619
rect 10689 8599 10709 8619
rect 10801 8599 10821 8619
rect 10897 8599 10917 8619
rect 11007 8599 11027 8619
rect 11103 8599 11123 8619
rect 15436 8640 15456 8660
rect 13867 8539 13887 8559
rect 13963 8539 13983 8559
rect 14073 8539 14093 8559
rect 14169 8539 14189 8559
rect 14281 8539 14301 8559
rect 14377 8539 14397 8559
rect 14494 8539 14514 8559
rect 15532 8640 15552 8660
rect 15649 8640 15669 8660
rect 15745 8640 15765 8660
rect 15857 8640 15877 8660
rect 15953 8640 15973 8660
rect 16063 8640 16083 8660
rect 16159 8640 16179 8660
rect 14590 8539 14610 8559
rect 18923 8580 18943 8600
rect 19019 8580 19039 8600
rect 19129 8580 19149 8600
rect 19225 8580 19245 8600
rect 19337 8580 19357 8600
rect 19433 8580 19453 8600
rect 19550 8580 19570 8600
rect 19646 8580 19666 8600
rect 1429 8312 1449 8332
rect 1525 8312 1545 8332
rect 1642 8312 1662 8332
rect 1738 8312 1758 8332
rect 1850 8312 1870 8332
rect 1946 8312 1966 8332
rect 2056 8312 2076 8332
rect 2152 8312 2172 8332
rect 6485 8353 6505 8373
rect 2758 8267 2778 8287
rect 2854 8267 2874 8287
rect 2964 8267 2984 8287
rect 3060 8267 3080 8287
rect 3172 8267 3192 8287
rect 3268 8267 3288 8287
rect 3385 8267 3405 8287
rect 6581 8353 6601 8373
rect 6698 8353 6718 8373
rect 6794 8353 6814 8373
rect 6906 8353 6926 8373
rect 7002 8353 7022 8373
rect 7112 8353 7132 8373
rect 7208 8353 7228 8373
rect 3481 8267 3501 8287
rect 7814 8308 7834 8328
rect 7910 8308 7930 8328
rect 8020 8308 8040 8328
rect 8116 8308 8136 8328
rect 8228 8308 8248 8328
rect 8324 8308 8344 8328
rect 8441 8308 8461 8328
rect 8537 8308 8557 8328
rect 11460 8317 11480 8337
rect 11556 8317 11576 8337
rect 11673 8317 11693 8337
rect 11769 8317 11789 8337
rect 11881 8317 11901 8337
rect 11977 8317 11997 8337
rect 12087 8317 12107 8337
rect 12183 8317 12203 8337
rect 16516 8358 16536 8378
rect 12789 8272 12809 8292
rect 12885 8272 12905 8292
rect 12995 8272 13015 8292
rect 13091 8272 13111 8292
rect 13203 8272 13223 8292
rect 13299 8272 13319 8292
rect 13416 8272 13436 8292
rect 16612 8358 16632 8378
rect 16729 8358 16749 8378
rect 16825 8358 16845 8378
rect 16937 8358 16957 8378
rect 17033 8358 17053 8378
rect 17143 8358 17163 8378
rect 17239 8358 17259 8378
rect 13512 8272 13532 8292
rect 17845 8313 17865 8333
rect 17941 8313 17961 8333
rect 18051 8313 18071 8333
rect 18147 8313 18167 8333
rect 18259 8313 18279 8333
rect 18355 8313 18375 8333
rect 18472 8313 18492 8333
rect 18568 8313 18588 8333
rect 351 8045 371 8065
rect 447 8045 467 8065
rect 564 8045 584 8065
rect 660 8045 680 8065
rect 772 8045 792 8065
rect 868 8045 888 8065
rect 978 8045 998 8065
rect 1074 8045 1094 8065
rect 5407 8086 5427 8106
rect 3838 7985 3858 8005
rect 3934 7985 3954 8005
rect 4044 7985 4064 8005
rect 4140 7985 4160 8005
rect 4252 7985 4272 8005
rect 4348 7985 4368 8005
rect 4465 7985 4485 8005
rect 5503 8086 5523 8106
rect 5620 8086 5640 8106
rect 5716 8086 5736 8106
rect 5828 8086 5848 8106
rect 5924 8086 5944 8106
rect 6034 8086 6054 8106
rect 6130 8086 6150 8106
rect 4561 7985 4581 8005
rect 8894 8026 8914 8046
rect 8990 8026 9010 8046
rect 9100 8026 9120 8046
rect 9196 8026 9216 8046
rect 9308 8026 9328 8046
rect 9404 8026 9424 8046
rect 9521 8026 9541 8046
rect 9617 8026 9637 8046
rect 10382 8050 10402 8070
rect 10478 8050 10498 8070
rect 10595 8050 10615 8070
rect 10691 8050 10711 8070
rect 10803 8050 10823 8070
rect 10899 8050 10919 8070
rect 11009 8050 11029 8070
rect 11105 8050 11125 8070
rect 15438 8091 15458 8111
rect 1289 7801 1309 7821
rect 1385 7801 1405 7821
rect 1502 7801 1522 7821
rect 1598 7801 1618 7821
rect 1710 7801 1730 7821
rect 1806 7801 1826 7821
rect 1916 7801 1936 7821
rect 2012 7801 2032 7821
rect 6345 7842 6365 7862
rect 2899 7675 2919 7695
rect 2995 7675 3015 7695
rect 3105 7675 3125 7695
rect 3201 7675 3221 7695
rect 3313 7675 3333 7695
rect 3409 7675 3429 7695
rect 3526 7675 3546 7695
rect 6441 7842 6461 7862
rect 6558 7842 6578 7862
rect 6654 7842 6674 7862
rect 6766 7842 6786 7862
rect 6862 7842 6882 7862
rect 6972 7842 6992 7862
rect 13869 7990 13889 8010
rect 7068 7842 7088 7862
rect 13965 7990 13985 8010
rect 14075 7990 14095 8010
rect 14171 7990 14191 8010
rect 14283 7990 14303 8010
rect 14379 7990 14399 8010
rect 14496 7990 14516 8010
rect 15534 8091 15554 8111
rect 15651 8091 15671 8111
rect 15747 8091 15767 8111
rect 15859 8091 15879 8111
rect 15955 8091 15975 8111
rect 16065 8091 16085 8111
rect 16161 8091 16181 8111
rect 14592 7990 14612 8010
rect 18925 8031 18945 8051
rect 19021 8031 19041 8051
rect 19131 8031 19151 8051
rect 19227 8031 19247 8051
rect 19339 8031 19359 8051
rect 19435 8031 19455 8051
rect 19552 8031 19572 8051
rect 19648 8031 19668 8051
rect 3622 7675 3642 7695
rect 7955 7716 7975 7736
rect 8051 7716 8071 7736
rect 8161 7716 8181 7736
rect 8257 7716 8277 7736
rect 8369 7716 8389 7736
rect 8465 7716 8485 7736
rect 8582 7716 8602 7736
rect 11320 7806 11340 7826
rect 8678 7716 8698 7736
rect 11416 7806 11436 7826
rect 11533 7806 11553 7826
rect 11629 7806 11649 7826
rect 11741 7806 11761 7826
rect 11837 7806 11857 7826
rect 11947 7806 11967 7826
rect 12043 7806 12063 7826
rect 16376 7847 16396 7867
rect 350 7491 370 7511
rect 446 7491 466 7511
rect 563 7491 583 7511
rect 659 7491 679 7511
rect 771 7491 791 7511
rect 867 7491 887 7511
rect 977 7491 997 7511
rect 1073 7491 1093 7511
rect 5406 7532 5426 7552
rect 3837 7431 3857 7451
rect 3933 7431 3953 7451
rect 4043 7431 4063 7451
rect 4139 7431 4159 7451
rect 4251 7431 4271 7451
rect 4347 7431 4367 7451
rect 4464 7431 4484 7451
rect 5502 7532 5522 7552
rect 5619 7532 5639 7552
rect 5715 7532 5735 7552
rect 5827 7532 5847 7552
rect 5923 7532 5943 7552
rect 6033 7532 6053 7552
rect 12930 7680 12950 7700
rect 6129 7532 6149 7552
rect 13026 7680 13046 7700
rect 13136 7680 13156 7700
rect 13232 7680 13252 7700
rect 13344 7680 13364 7700
rect 13440 7680 13460 7700
rect 13557 7680 13577 7700
rect 16472 7847 16492 7867
rect 16589 7847 16609 7867
rect 16685 7847 16705 7867
rect 16797 7847 16817 7867
rect 16893 7847 16913 7867
rect 17003 7847 17023 7867
rect 17099 7847 17119 7867
rect 13653 7680 13673 7700
rect 17986 7721 18006 7741
rect 18082 7721 18102 7741
rect 18192 7721 18212 7741
rect 18288 7721 18308 7741
rect 18400 7721 18420 7741
rect 18496 7721 18516 7741
rect 18613 7721 18633 7741
rect 18709 7721 18729 7741
rect 4560 7431 4580 7451
rect 8893 7472 8913 7492
rect 8989 7472 9009 7492
rect 9099 7472 9119 7492
rect 9195 7472 9215 7492
rect 9307 7472 9327 7492
rect 9403 7472 9423 7492
rect 9520 7472 9540 7492
rect 9616 7472 9636 7492
rect 10381 7496 10401 7516
rect 10477 7496 10497 7516
rect 10594 7496 10614 7516
rect 10690 7496 10710 7516
rect 10802 7496 10822 7516
rect 10898 7496 10918 7516
rect 11008 7496 11028 7516
rect 11104 7496 11124 7516
rect 15437 7537 15457 7557
rect 13868 7436 13888 7456
rect 13964 7436 13984 7456
rect 14074 7436 14094 7456
rect 14170 7436 14190 7456
rect 14282 7436 14302 7456
rect 14378 7436 14398 7456
rect 14495 7436 14515 7456
rect 15533 7537 15553 7557
rect 15650 7537 15670 7557
rect 15746 7537 15766 7557
rect 15858 7537 15878 7557
rect 15954 7537 15974 7557
rect 16064 7537 16084 7557
rect 16160 7537 16180 7557
rect 14591 7436 14611 7456
rect 18924 7477 18944 7497
rect 19020 7477 19040 7497
rect 19130 7477 19150 7497
rect 19226 7477 19246 7497
rect 19338 7477 19358 7497
rect 19434 7477 19454 7497
rect 19551 7477 19571 7497
rect 19647 7477 19667 7497
rect 1399 7222 1419 7242
rect 1495 7222 1515 7242
rect 1612 7222 1632 7242
rect 1708 7222 1728 7242
rect 1820 7222 1840 7242
rect 1916 7222 1936 7242
rect 2026 7222 2046 7242
rect 2122 7222 2142 7242
rect 6455 7263 6475 7283
rect 6551 7263 6571 7283
rect 6668 7263 6688 7283
rect 6764 7263 6784 7283
rect 6876 7263 6896 7283
rect 6972 7263 6992 7283
rect 7082 7263 7102 7283
rect 7178 7263 7198 7283
rect 2789 7151 2809 7171
rect 2885 7151 2905 7171
rect 2995 7151 3015 7171
rect 3091 7151 3111 7171
rect 3203 7151 3223 7171
rect 3299 7151 3319 7171
rect 3416 7151 3436 7171
rect 3512 7151 3532 7171
rect 7845 7192 7865 7212
rect 7941 7192 7961 7212
rect 8051 7192 8071 7212
rect 8147 7192 8167 7212
rect 8259 7192 8279 7212
rect 8355 7192 8375 7212
rect 8472 7192 8492 7212
rect 8568 7192 8588 7212
rect 11430 7227 11450 7247
rect 11526 7227 11546 7247
rect 11643 7227 11663 7247
rect 11739 7227 11759 7247
rect 11851 7227 11871 7247
rect 11947 7227 11967 7247
rect 12057 7227 12077 7247
rect 12153 7227 12173 7247
rect 16486 7268 16506 7288
rect 16582 7268 16602 7288
rect 16699 7268 16719 7288
rect 16795 7268 16815 7288
rect 16907 7268 16927 7288
rect 17003 7268 17023 7288
rect 17113 7268 17133 7288
rect 17209 7268 17229 7288
rect 12820 7156 12840 7176
rect 12916 7156 12936 7176
rect 13026 7156 13046 7176
rect 13122 7156 13142 7176
rect 13234 7156 13254 7176
rect 13330 7156 13350 7176
rect 13447 7156 13467 7176
rect 13543 7156 13563 7176
rect 17876 7197 17896 7217
rect 17972 7197 17992 7217
rect 18082 7197 18102 7217
rect 18178 7197 18198 7217
rect 18290 7197 18310 7217
rect 18386 7197 18406 7217
rect 18503 7197 18523 7217
rect 18599 7197 18619 7217
rect 351 6942 371 6962
rect 447 6942 467 6962
rect 564 6942 584 6962
rect 660 6942 680 6962
rect 772 6942 792 6962
rect 868 6942 888 6962
rect 978 6942 998 6962
rect 1074 6942 1094 6962
rect 5407 6983 5427 7003
rect 3838 6882 3858 6902
rect 3934 6882 3954 6902
rect 4044 6882 4064 6902
rect 4140 6882 4160 6902
rect 4252 6882 4272 6902
rect 4348 6882 4368 6902
rect 4465 6882 4485 6902
rect 5503 6983 5523 7003
rect 5620 6983 5640 7003
rect 5716 6983 5736 7003
rect 5828 6983 5848 7003
rect 5924 6983 5944 7003
rect 6034 6983 6054 7003
rect 6130 6983 6150 7003
rect 4561 6882 4581 6902
rect 8894 6923 8914 6943
rect 8990 6923 9010 6943
rect 9100 6923 9120 6943
rect 9196 6923 9216 6943
rect 9308 6923 9328 6943
rect 9404 6923 9424 6943
rect 9521 6923 9541 6943
rect 9617 6923 9637 6943
rect 10382 6947 10402 6967
rect 10478 6947 10498 6967
rect 10595 6947 10615 6967
rect 10691 6947 10711 6967
rect 10803 6947 10823 6967
rect 10899 6947 10919 6967
rect 11009 6947 11029 6967
rect 11105 6947 11125 6967
rect 15438 6988 15458 7008
rect 1289 6698 1309 6718
rect 1385 6698 1405 6718
rect 1502 6698 1522 6718
rect 1598 6698 1618 6718
rect 1710 6698 1730 6718
rect 1806 6698 1826 6718
rect 1916 6698 1936 6718
rect 2012 6698 2032 6718
rect 6345 6739 6365 6759
rect 2899 6572 2919 6592
rect 2995 6572 3015 6592
rect 3105 6572 3125 6592
rect 3201 6572 3221 6592
rect 3313 6572 3333 6592
rect 3409 6572 3429 6592
rect 3526 6572 3546 6592
rect 6441 6739 6461 6759
rect 6558 6739 6578 6759
rect 6654 6739 6674 6759
rect 6766 6739 6786 6759
rect 6862 6739 6882 6759
rect 6972 6739 6992 6759
rect 13869 6887 13889 6907
rect 7068 6739 7088 6759
rect 13965 6887 13985 6907
rect 14075 6887 14095 6907
rect 14171 6887 14191 6907
rect 14283 6887 14303 6907
rect 14379 6887 14399 6907
rect 14496 6887 14516 6907
rect 15534 6988 15554 7008
rect 15651 6988 15671 7008
rect 15747 6988 15767 7008
rect 15859 6988 15879 7008
rect 15955 6988 15975 7008
rect 16065 6988 16085 7008
rect 16161 6988 16181 7008
rect 14592 6887 14612 6907
rect 18925 6928 18945 6948
rect 19021 6928 19041 6948
rect 19131 6928 19151 6948
rect 19227 6928 19247 6948
rect 19339 6928 19359 6948
rect 19435 6928 19455 6948
rect 19552 6928 19572 6948
rect 19648 6928 19668 6948
rect 3622 6572 3642 6592
rect 7955 6613 7975 6633
rect 8051 6613 8071 6633
rect 8161 6613 8181 6633
rect 8257 6613 8277 6633
rect 8369 6613 8389 6633
rect 8465 6613 8485 6633
rect 8582 6613 8602 6633
rect 11320 6703 11340 6723
rect 8678 6613 8698 6633
rect 11416 6703 11436 6723
rect 11533 6703 11553 6723
rect 11629 6703 11649 6723
rect 11741 6703 11761 6723
rect 11837 6703 11857 6723
rect 11947 6703 11967 6723
rect 12043 6703 12063 6723
rect 16376 6744 16396 6764
rect 350 6388 370 6408
rect 446 6388 466 6408
rect 563 6388 583 6408
rect 659 6388 679 6408
rect 771 6388 791 6408
rect 867 6388 887 6408
rect 977 6388 997 6408
rect 1073 6388 1093 6408
rect 5406 6429 5426 6449
rect 3837 6328 3857 6348
rect 3933 6328 3953 6348
rect 4043 6328 4063 6348
rect 4139 6328 4159 6348
rect 4251 6328 4271 6348
rect 4347 6328 4367 6348
rect 4464 6328 4484 6348
rect 5502 6429 5522 6449
rect 5619 6429 5639 6449
rect 5715 6429 5735 6449
rect 5827 6429 5847 6449
rect 5923 6429 5943 6449
rect 6033 6429 6053 6449
rect 12930 6577 12950 6597
rect 6129 6429 6149 6449
rect 13026 6577 13046 6597
rect 13136 6577 13156 6597
rect 13232 6577 13252 6597
rect 13344 6577 13364 6597
rect 13440 6577 13460 6597
rect 13557 6577 13577 6597
rect 16472 6744 16492 6764
rect 16589 6744 16609 6764
rect 16685 6744 16705 6764
rect 16797 6744 16817 6764
rect 16893 6744 16913 6764
rect 17003 6744 17023 6764
rect 17099 6744 17119 6764
rect 13653 6577 13673 6597
rect 17986 6618 18006 6638
rect 18082 6618 18102 6638
rect 18192 6618 18212 6638
rect 18288 6618 18308 6638
rect 18400 6618 18420 6638
rect 18496 6618 18516 6638
rect 18613 6618 18633 6638
rect 18709 6618 18729 6638
rect 4560 6328 4580 6348
rect 8893 6369 8913 6389
rect 8989 6369 9009 6389
rect 9099 6369 9119 6389
rect 9195 6369 9215 6389
rect 9307 6369 9327 6389
rect 9403 6369 9423 6389
rect 9520 6369 9540 6389
rect 9616 6369 9636 6389
rect 10381 6393 10401 6413
rect 10477 6393 10497 6413
rect 10594 6393 10614 6413
rect 10690 6393 10710 6413
rect 10802 6393 10822 6413
rect 10898 6393 10918 6413
rect 11008 6393 11028 6413
rect 11104 6393 11124 6413
rect 15437 6434 15457 6454
rect 13868 6333 13888 6353
rect 13964 6333 13984 6353
rect 14074 6333 14094 6353
rect 14170 6333 14190 6353
rect 14282 6333 14302 6353
rect 14378 6333 14398 6353
rect 14495 6333 14515 6353
rect 15533 6434 15553 6454
rect 15650 6434 15670 6454
rect 15746 6434 15766 6454
rect 15858 6434 15878 6454
rect 15954 6434 15974 6454
rect 16064 6434 16084 6454
rect 16160 6434 16180 6454
rect 14591 6333 14611 6353
rect 18924 6374 18944 6394
rect 19020 6374 19040 6394
rect 19130 6374 19150 6394
rect 19226 6374 19246 6394
rect 19338 6374 19358 6394
rect 19434 6374 19454 6394
rect 19551 6374 19571 6394
rect 19647 6374 19667 6394
rect 1430 6106 1450 6126
rect 1526 6106 1546 6126
rect 1643 6106 1663 6126
rect 1739 6106 1759 6126
rect 1851 6106 1871 6126
rect 1947 6106 1967 6126
rect 2057 6106 2077 6126
rect 2153 6106 2173 6126
rect 6486 6147 6506 6167
rect 2759 6061 2779 6081
rect 2855 6061 2875 6081
rect 2965 6061 2985 6081
rect 3061 6061 3081 6081
rect 3173 6061 3193 6081
rect 3269 6061 3289 6081
rect 3386 6061 3406 6081
rect 6582 6147 6602 6167
rect 6699 6147 6719 6167
rect 6795 6147 6815 6167
rect 6907 6147 6927 6167
rect 7003 6147 7023 6167
rect 7113 6147 7133 6167
rect 7209 6147 7229 6167
rect 3482 6061 3502 6081
rect 7815 6102 7835 6122
rect 7911 6102 7931 6122
rect 8021 6102 8041 6122
rect 8117 6102 8137 6122
rect 8229 6102 8249 6122
rect 8325 6102 8345 6122
rect 8442 6102 8462 6122
rect 8538 6102 8558 6122
rect 11461 6111 11481 6131
rect 11557 6111 11577 6131
rect 11674 6111 11694 6131
rect 11770 6111 11790 6131
rect 11882 6111 11902 6131
rect 11978 6111 11998 6131
rect 12088 6111 12108 6131
rect 12184 6111 12204 6131
rect 16517 6152 16537 6172
rect 12790 6066 12810 6086
rect 12886 6066 12906 6086
rect 12996 6066 13016 6086
rect 13092 6066 13112 6086
rect 13204 6066 13224 6086
rect 13300 6066 13320 6086
rect 13417 6066 13437 6086
rect 16613 6152 16633 6172
rect 16730 6152 16750 6172
rect 16826 6152 16846 6172
rect 16938 6152 16958 6172
rect 17034 6152 17054 6172
rect 17144 6152 17164 6172
rect 17240 6152 17260 6172
rect 13513 6066 13533 6086
rect 17846 6107 17866 6127
rect 17942 6107 17962 6127
rect 18052 6107 18072 6127
rect 18148 6107 18168 6127
rect 18260 6107 18280 6127
rect 18356 6107 18376 6127
rect 18473 6107 18493 6127
rect 18569 6107 18589 6127
rect 352 5839 372 5859
rect 448 5839 468 5859
rect 565 5839 585 5859
rect 661 5839 681 5859
rect 773 5839 793 5859
rect 869 5839 889 5859
rect 979 5839 999 5859
rect 1075 5839 1095 5859
rect 5408 5880 5428 5900
rect 3839 5779 3859 5799
rect 3935 5779 3955 5799
rect 4045 5779 4065 5799
rect 4141 5779 4161 5799
rect 4253 5779 4273 5799
rect 4349 5779 4369 5799
rect 4466 5779 4486 5799
rect 5504 5880 5524 5900
rect 5621 5880 5641 5900
rect 5717 5880 5737 5900
rect 5829 5880 5849 5900
rect 5925 5880 5945 5900
rect 6035 5880 6055 5900
rect 6131 5880 6151 5900
rect 4562 5779 4582 5799
rect 8895 5820 8915 5840
rect 8991 5820 9011 5840
rect 9101 5820 9121 5840
rect 9197 5820 9217 5840
rect 9309 5820 9329 5840
rect 9405 5820 9425 5840
rect 9522 5820 9542 5840
rect 9618 5820 9638 5840
rect 10383 5844 10403 5864
rect 10479 5844 10499 5864
rect 10596 5844 10616 5864
rect 10692 5844 10712 5864
rect 10804 5844 10824 5864
rect 10900 5844 10920 5864
rect 11010 5844 11030 5864
rect 11106 5844 11126 5864
rect 15439 5885 15459 5905
rect 1290 5595 1310 5615
rect 1386 5595 1406 5615
rect 1503 5595 1523 5615
rect 1599 5595 1619 5615
rect 1711 5595 1731 5615
rect 1807 5595 1827 5615
rect 1917 5595 1937 5615
rect 2013 5595 2033 5615
rect 6346 5636 6366 5656
rect 2900 5469 2920 5489
rect 2996 5469 3016 5489
rect 3106 5469 3126 5489
rect 3202 5469 3222 5489
rect 3314 5469 3334 5489
rect 3410 5469 3430 5489
rect 3527 5469 3547 5489
rect 6442 5636 6462 5656
rect 6559 5636 6579 5656
rect 6655 5636 6675 5656
rect 6767 5636 6787 5656
rect 6863 5636 6883 5656
rect 6973 5636 6993 5656
rect 13870 5784 13890 5804
rect 7069 5636 7089 5656
rect 13966 5784 13986 5804
rect 14076 5784 14096 5804
rect 14172 5784 14192 5804
rect 14284 5784 14304 5804
rect 14380 5784 14400 5804
rect 14497 5784 14517 5804
rect 15535 5885 15555 5905
rect 15652 5885 15672 5905
rect 15748 5885 15768 5905
rect 15860 5885 15880 5905
rect 15956 5885 15976 5905
rect 16066 5885 16086 5905
rect 16162 5885 16182 5905
rect 14593 5784 14613 5804
rect 18926 5825 18946 5845
rect 19022 5825 19042 5845
rect 19132 5825 19152 5845
rect 19228 5825 19248 5845
rect 19340 5825 19360 5845
rect 19436 5825 19456 5845
rect 19553 5825 19573 5845
rect 19649 5825 19669 5845
rect 3623 5469 3643 5489
rect 7956 5510 7976 5530
rect 8052 5510 8072 5530
rect 8162 5510 8182 5530
rect 8258 5510 8278 5530
rect 8370 5510 8390 5530
rect 8466 5510 8486 5530
rect 8583 5510 8603 5530
rect 11321 5600 11341 5620
rect 8679 5510 8699 5530
rect 11417 5600 11437 5620
rect 11534 5600 11554 5620
rect 11630 5600 11650 5620
rect 11742 5600 11762 5620
rect 11838 5600 11858 5620
rect 11948 5600 11968 5620
rect 12044 5600 12064 5620
rect 16377 5641 16397 5661
rect 351 5285 371 5305
rect 447 5285 467 5305
rect 564 5285 584 5305
rect 660 5285 680 5305
rect 772 5285 792 5305
rect 868 5285 888 5305
rect 978 5285 998 5305
rect 1074 5285 1094 5305
rect 5407 5326 5427 5346
rect 3838 5225 3858 5245
rect 3934 5225 3954 5245
rect 4044 5225 4064 5245
rect 4140 5225 4160 5245
rect 4252 5225 4272 5245
rect 4348 5225 4368 5245
rect 4465 5225 4485 5245
rect 5503 5326 5523 5346
rect 5620 5326 5640 5346
rect 5716 5326 5736 5346
rect 5828 5326 5848 5346
rect 5924 5326 5944 5346
rect 6034 5326 6054 5346
rect 12931 5474 12951 5494
rect 6130 5326 6150 5346
rect 13027 5474 13047 5494
rect 13137 5474 13157 5494
rect 13233 5474 13253 5494
rect 13345 5474 13365 5494
rect 13441 5474 13461 5494
rect 13558 5474 13578 5494
rect 16473 5641 16493 5661
rect 16590 5641 16610 5661
rect 16686 5641 16706 5661
rect 16798 5641 16818 5661
rect 16894 5641 16914 5661
rect 17004 5641 17024 5661
rect 17100 5641 17120 5661
rect 13654 5474 13674 5494
rect 17987 5515 18007 5535
rect 18083 5515 18103 5535
rect 18193 5515 18213 5535
rect 18289 5515 18309 5535
rect 18401 5515 18421 5535
rect 18497 5515 18517 5535
rect 18614 5515 18634 5535
rect 18710 5515 18730 5535
rect 4561 5225 4581 5245
rect 8894 5266 8914 5286
rect 8990 5266 9010 5286
rect 9100 5266 9120 5286
rect 9196 5266 9216 5286
rect 9308 5266 9328 5286
rect 9404 5266 9424 5286
rect 9521 5266 9541 5286
rect 9617 5266 9637 5286
rect 10382 5290 10402 5310
rect 10478 5290 10498 5310
rect 10595 5290 10615 5310
rect 10691 5290 10711 5310
rect 10803 5290 10823 5310
rect 10899 5290 10919 5310
rect 11009 5290 11029 5310
rect 11105 5290 11125 5310
rect 15438 5331 15458 5351
rect 1399 5022 1419 5042
rect 1495 5022 1515 5042
rect 1612 5022 1632 5042
rect 1708 5022 1728 5042
rect 1820 5022 1840 5042
rect 1916 5022 1936 5042
rect 2026 5022 2046 5042
rect 2122 5022 2142 5042
rect 6455 5063 6475 5083
rect 6551 5063 6571 5083
rect 6668 5063 6688 5083
rect 6764 5063 6784 5083
rect 6876 5063 6896 5083
rect 6972 5063 6992 5083
rect 7082 5063 7102 5083
rect 13869 5230 13889 5250
rect 13965 5230 13985 5250
rect 14075 5230 14095 5250
rect 14171 5230 14191 5250
rect 14283 5230 14303 5250
rect 14379 5230 14399 5250
rect 14496 5230 14516 5250
rect 15534 5331 15554 5351
rect 15651 5331 15671 5351
rect 15747 5331 15767 5351
rect 15859 5331 15879 5351
rect 15955 5331 15975 5351
rect 16065 5331 16085 5351
rect 16161 5331 16181 5351
rect 14592 5230 14612 5250
rect 18925 5271 18945 5291
rect 19021 5271 19041 5291
rect 19131 5271 19151 5291
rect 19227 5271 19247 5291
rect 19339 5271 19359 5291
rect 19435 5271 19455 5291
rect 19552 5271 19572 5291
rect 19648 5271 19668 5291
rect 7178 5063 7198 5083
rect 2791 4939 2811 4959
rect 2887 4939 2907 4959
rect 2997 4939 3017 4959
rect 3093 4939 3113 4959
rect 3205 4939 3225 4959
rect 3301 4939 3321 4959
rect 3418 4939 3438 4959
rect 3514 4939 3534 4959
rect 7847 4980 7867 5000
rect 7943 4980 7963 5000
rect 8053 4980 8073 5000
rect 8149 4980 8169 5000
rect 8261 4980 8281 5000
rect 8357 4980 8377 5000
rect 8474 4980 8494 5000
rect 8570 4980 8590 5000
rect 11430 5027 11450 5047
rect 11526 5027 11546 5047
rect 11643 5027 11663 5047
rect 11739 5027 11759 5047
rect 11851 5027 11871 5047
rect 11947 5027 11967 5047
rect 12057 5027 12077 5047
rect 12153 5027 12173 5047
rect 16486 5068 16506 5088
rect 16582 5068 16602 5088
rect 16699 5068 16719 5088
rect 16795 5068 16815 5088
rect 16907 5068 16927 5088
rect 17003 5068 17023 5088
rect 17113 5068 17133 5088
rect 17209 5068 17229 5088
rect 12822 4944 12842 4964
rect 352 4736 372 4756
rect 448 4736 468 4756
rect 565 4736 585 4756
rect 661 4736 681 4756
rect 773 4736 793 4756
rect 869 4736 889 4756
rect 979 4736 999 4756
rect 1075 4736 1095 4756
rect 5408 4777 5428 4797
rect 3839 4676 3859 4696
rect 3935 4676 3955 4696
rect 4045 4676 4065 4696
rect 4141 4676 4161 4696
rect 4253 4676 4273 4696
rect 4349 4676 4369 4696
rect 4466 4676 4486 4696
rect 5504 4777 5524 4797
rect 5621 4777 5641 4797
rect 5717 4777 5737 4797
rect 5829 4777 5849 4797
rect 5925 4777 5945 4797
rect 6035 4777 6055 4797
rect 6131 4777 6151 4797
rect 12918 4944 12938 4964
rect 13028 4944 13048 4964
rect 13124 4944 13144 4964
rect 13236 4944 13256 4964
rect 13332 4944 13352 4964
rect 13449 4944 13469 4964
rect 13545 4944 13565 4964
rect 17878 4985 17898 5005
rect 17974 4985 17994 5005
rect 18084 4985 18104 5005
rect 18180 4985 18200 5005
rect 18292 4985 18312 5005
rect 18388 4985 18408 5005
rect 18505 4985 18525 5005
rect 18601 4985 18621 5005
rect 4562 4676 4582 4696
rect 8895 4717 8915 4737
rect 8991 4717 9011 4737
rect 9101 4717 9121 4737
rect 9197 4717 9217 4737
rect 9309 4717 9329 4737
rect 9405 4717 9425 4737
rect 9522 4717 9542 4737
rect 9618 4717 9638 4737
rect 10383 4741 10403 4761
rect 10479 4741 10499 4761
rect 10596 4741 10616 4761
rect 10692 4741 10712 4761
rect 10804 4741 10824 4761
rect 10900 4741 10920 4761
rect 11010 4741 11030 4761
rect 11106 4741 11126 4761
rect 15439 4782 15459 4802
rect 1290 4492 1310 4512
rect 1386 4492 1406 4512
rect 1503 4492 1523 4512
rect 1599 4492 1619 4512
rect 1711 4492 1731 4512
rect 1807 4492 1827 4512
rect 1917 4492 1937 4512
rect 2013 4492 2033 4512
rect 6346 4533 6366 4553
rect 2900 4366 2920 4386
rect 2996 4366 3016 4386
rect 3106 4366 3126 4386
rect 3202 4366 3222 4386
rect 3314 4366 3334 4386
rect 3410 4366 3430 4386
rect 3527 4366 3547 4386
rect 6442 4533 6462 4553
rect 6559 4533 6579 4553
rect 6655 4533 6675 4553
rect 6767 4533 6787 4553
rect 6863 4533 6883 4553
rect 6973 4533 6993 4553
rect 13870 4681 13890 4701
rect 7069 4533 7089 4553
rect 13966 4681 13986 4701
rect 14076 4681 14096 4701
rect 14172 4681 14192 4701
rect 14284 4681 14304 4701
rect 14380 4681 14400 4701
rect 14497 4681 14517 4701
rect 15535 4782 15555 4802
rect 15652 4782 15672 4802
rect 15748 4782 15768 4802
rect 15860 4782 15880 4802
rect 15956 4782 15976 4802
rect 16066 4782 16086 4802
rect 16162 4782 16182 4802
rect 14593 4681 14613 4701
rect 18926 4722 18946 4742
rect 19022 4722 19042 4742
rect 19132 4722 19152 4742
rect 19228 4722 19248 4742
rect 19340 4722 19360 4742
rect 19436 4722 19456 4742
rect 19553 4722 19573 4742
rect 19649 4722 19669 4742
rect 3623 4366 3643 4386
rect 7956 4407 7976 4427
rect 8052 4407 8072 4427
rect 8162 4407 8182 4427
rect 8258 4407 8278 4427
rect 8370 4407 8390 4427
rect 8466 4407 8486 4427
rect 8583 4407 8603 4427
rect 11321 4497 11341 4517
rect 8679 4407 8699 4427
rect 11417 4497 11437 4517
rect 11534 4497 11554 4517
rect 11630 4497 11650 4517
rect 11742 4497 11762 4517
rect 11838 4497 11858 4517
rect 11948 4497 11968 4517
rect 12044 4497 12064 4517
rect 16377 4538 16397 4558
rect 351 4182 371 4202
rect 447 4182 467 4202
rect 564 4182 584 4202
rect 660 4182 680 4202
rect 772 4182 792 4202
rect 868 4182 888 4202
rect 978 4182 998 4202
rect 1074 4182 1094 4202
rect 5407 4223 5427 4243
rect 3838 4122 3858 4142
rect 3934 4122 3954 4142
rect 4044 4122 4064 4142
rect 4140 4122 4160 4142
rect 4252 4122 4272 4142
rect 4348 4122 4368 4142
rect 4465 4122 4485 4142
rect 5503 4223 5523 4243
rect 5620 4223 5640 4243
rect 5716 4223 5736 4243
rect 5828 4223 5848 4243
rect 5924 4223 5944 4243
rect 6034 4223 6054 4243
rect 12931 4371 12951 4391
rect 6130 4223 6150 4243
rect 13027 4371 13047 4391
rect 13137 4371 13157 4391
rect 13233 4371 13253 4391
rect 13345 4371 13365 4391
rect 13441 4371 13461 4391
rect 13558 4371 13578 4391
rect 16473 4538 16493 4558
rect 16590 4538 16610 4558
rect 16686 4538 16706 4558
rect 16798 4538 16818 4558
rect 16894 4538 16914 4558
rect 17004 4538 17024 4558
rect 17100 4538 17120 4558
rect 13654 4371 13674 4391
rect 17987 4412 18007 4432
rect 18083 4412 18103 4432
rect 18193 4412 18213 4432
rect 18289 4412 18309 4432
rect 18401 4412 18421 4432
rect 18497 4412 18517 4432
rect 18614 4412 18634 4432
rect 18710 4412 18730 4432
rect 4561 4122 4581 4142
rect 8894 4163 8914 4183
rect 8990 4163 9010 4183
rect 9100 4163 9120 4183
rect 9196 4163 9216 4183
rect 9308 4163 9328 4183
rect 9404 4163 9424 4183
rect 9521 4163 9541 4183
rect 9617 4163 9637 4183
rect 10382 4187 10402 4207
rect 10478 4187 10498 4207
rect 10595 4187 10615 4207
rect 10691 4187 10711 4207
rect 10803 4187 10823 4207
rect 10899 4187 10919 4207
rect 11009 4187 11029 4207
rect 11105 4187 11125 4207
rect 15438 4228 15458 4248
rect 13869 4127 13889 4147
rect 13965 4127 13985 4147
rect 14075 4127 14095 4147
rect 14171 4127 14191 4147
rect 14283 4127 14303 4147
rect 14379 4127 14399 4147
rect 14496 4127 14516 4147
rect 15534 4228 15554 4248
rect 15651 4228 15671 4248
rect 15747 4228 15767 4248
rect 15859 4228 15879 4248
rect 15955 4228 15975 4248
rect 16065 4228 16085 4248
rect 16161 4228 16181 4248
rect 14592 4127 14612 4147
rect 18925 4168 18945 4188
rect 19021 4168 19041 4188
rect 19131 4168 19151 4188
rect 19227 4168 19247 4188
rect 19339 4168 19359 4188
rect 19435 4168 19455 4188
rect 19552 4168 19572 4188
rect 19648 4168 19668 4188
rect 1431 3900 1451 3920
rect 1527 3900 1547 3920
rect 1644 3900 1664 3920
rect 1740 3900 1760 3920
rect 1852 3900 1872 3920
rect 1948 3900 1968 3920
rect 2058 3900 2078 3920
rect 2154 3900 2174 3920
rect 6487 3941 6507 3961
rect 2760 3855 2780 3875
rect 2856 3855 2876 3875
rect 2966 3855 2986 3875
rect 3062 3855 3082 3875
rect 3174 3855 3194 3875
rect 3270 3855 3290 3875
rect 3387 3855 3407 3875
rect 6583 3941 6603 3961
rect 6700 3941 6720 3961
rect 6796 3941 6816 3961
rect 6908 3941 6928 3961
rect 7004 3941 7024 3961
rect 7114 3941 7134 3961
rect 7210 3941 7230 3961
rect 3483 3855 3503 3875
rect 7816 3896 7836 3916
rect 7912 3896 7932 3916
rect 8022 3896 8042 3916
rect 8118 3896 8138 3916
rect 8230 3896 8250 3916
rect 8326 3896 8346 3916
rect 8443 3896 8463 3916
rect 8539 3896 8559 3916
rect 11462 3905 11482 3925
rect 11558 3905 11578 3925
rect 11675 3905 11695 3925
rect 11771 3905 11791 3925
rect 11883 3905 11903 3925
rect 11979 3905 11999 3925
rect 12089 3905 12109 3925
rect 12185 3905 12205 3925
rect 16518 3946 16538 3966
rect 12791 3860 12811 3880
rect 12887 3860 12907 3880
rect 12997 3860 13017 3880
rect 13093 3860 13113 3880
rect 13205 3860 13225 3880
rect 13301 3860 13321 3880
rect 13418 3860 13438 3880
rect 16614 3946 16634 3966
rect 16731 3946 16751 3966
rect 16827 3946 16847 3966
rect 16939 3946 16959 3966
rect 17035 3946 17055 3966
rect 17145 3946 17165 3966
rect 17241 3946 17261 3966
rect 13514 3860 13534 3880
rect 17847 3901 17867 3921
rect 17943 3901 17963 3921
rect 18053 3901 18073 3921
rect 18149 3901 18169 3921
rect 18261 3901 18281 3921
rect 18357 3901 18377 3921
rect 18474 3901 18494 3921
rect 18570 3901 18590 3921
rect 353 3633 373 3653
rect 449 3633 469 3653
rect 566 3633 586 3653
rect 662 3633 682 3653
rect 774 3633 794 3653
rect 870 3633 890 3653
rect 980 3633 1000 3653
rect 1076 3633 1096 3653
rect 5409 3674 5429 3694
rect 3840 3573 3860 3593
rect 3936 3573 3956 3593
rect 4046 3573 4066 3593
rect 4142 3573 4162 3593
rect 4254 3573 4274 3593
rect 4350 3573 4370 3593
rect 4467 3573 4487 3593
rect 5505 3674 5525 3694
rect 5622 3674 5642 3694
rect 5718 3674 5738 3694
rect 5830 3674 5850 3694
rect 5926 3674 5946 3694
rect 6036 3674 6056 3694
rect 6132 3674 6152 3694
rect 4563 3573 4583 3593
rect 8896 3614 8916 3634
rect 8992 3614 9012 3634
rect 9102 3614 9122 3634
rect 9198 3614 9218 3634
rect 9310 3614 9330 3634
rect 9406 3614 9426 3634
rect 9523 3614 9543 3634
rect 9619 3614 9639 3634
rect 10384 3638 10404 3658
rect 10480 3638 10500 3658
rect 10597 3638 10617 3658
rect 10693 3638 10713 3658
rect 10805 3638 10825 3658
rect 10901 3638 10921 3658
rect 11011 3638 11031 3658
rect 11107 3638 11127 3658
rect 15440 3679 15460 3699
rect 1291 3389 1311 3409
rect 1387 3389 1407 3409
rect 1504 3389 1524 3409
rect 1600 3389 1620 3409
rect 1712 3389 1732 3409
rect 1808 3389 1828 3409
rect 1918 3389 1938 3409
rect 2014 3389 2034 3409
rect 6347 3430 6367 3450
rect 2901 3263 2921 3283
rect 2997 3263 3017 3283
rect 3107 3263 3127 3283
rect 3203 3263 3223 3283
rect 3315 3263 3335 3283
rect 3411 3263 3431 3283
rect 3528 3263 3548 3283
rect 6443 3430 6463 3450
rect 6560 3430 6580 3450
rect 6656 3430 6676 3450
rect 6768 3430 6788 3450
rect 6864 3430 6884 3450
rect 6974 3430 6994 3450
rect 13871 3578 13891 3598
rect 7070 3430 7090 3450
rect 13967 3578 13987 3598
rect 14077 3578 14097 3598
rect 14173 3578 14193 3598
rect 14285 3578 14305 3598
rect 14381 3578 14401 3598
rect 14498 3578 14518 3598
rect 15536 3679 15556 3699
rect 15653 3679 15673 3699
rect 15749 3679 15769 3699
rect 15861 3679 15881 3699
rect 15957 3679 15977 3699
rect 16067 3679 16087 3699
rect 16163 3679 16183 3699
rect 14594 3578 14614 3598
rect 18927 3619 18947 3639
rect 19023 3619 19043 3639
rect 19133 3619 19153 3639
rect 19229 3619 19249 3639
rect 19341 3619 19361 3639
rect 19437 3619 19457 3639
rect 19554 3619 19574 3639
rect 19650 3619 19670 3639
rect 3624 3263 3644 3283
rect 7957 3304 7977 3324
rect 8053 3304 8073 3324
rect 8163 3304 8183 3324
rect 8259 3304 8279 3324
rect 8371 3304 8391 3324
rect 8467 3304 8487 3324
rect 8584 3304 8604 3324
rect 11322 3394 11342 3414
rect 8680 3304 8700 3324
rect 11418 3394 11438 3414
rect 11535 3394 11555 3414
rect 11631 3394 11651 3414
rect 11743 3394 11763 3414
rect 11839 3394 11859 3414
rect 11949 3394 11969 3414
rect 12045 3394 12065 3414
rect 16378 3435 16398 3455
rect 352 3079 372 3099
rect 448 3079 468 3099
rect 565 3079 585 3099
rect 661 3079 681 3099
rect 773 3079 793 3099
rect 869 3079 889 3099
rect 979 3079 999 3099
rect 1075 3079 1095 3099
rect 5408 3120 5428 3140
rect 3839 3019 3859 3039
rect 3935 3019 3955 3039
rect 4045 3019 4065 3039
rect 4141 3019 4161 3039
rect 4253 3019 4273 3039
rect 4349 3019 4369 3039
rect 4466 3019 4486 3039
rect 5504 3120 5524 3140
rect 5621 3120 5641 3140
rect 5717 3120 5737 3140
rect 5829 3120 5849 3140
rect 5925 3120 5945 3140
rect 6035 3120 6055 3140
rect 12932 3268 12952 3288
rect 6131 3120 6151 3140
rect 13028 3268 13048 3288
rect 13138 3268 13158 3288
rect 13234 3268 13254 3288
rect 13346 3268 13366 3288
rect 13442 3268 13462 3288
rect 13559 3268 13579 3288
rect 16474 3435 16494 3455
rect 16591 3435 16611 3455
rect 16687 3435 16707 3455
rect 16799 3435 16819 3455
rect 16895 3435 16915 3455
rect 17005 3435 17025 3455
rect 17101 3435 17121 3455
rect 13655 3268 13675 3288
rect 17988 3309 18008 3329
rect 18084 3309 18104 3329
rect 18194 3309 18214 3329
rect 18290 3309 18310 3329
rect 18402 3309 18422 3329
rect 18498 3309 18518 3329
rect 18615 3309 18635 3329
rect 18711 3309 18731 3329
rect 4562 3019 4582 3039
rect 8895 3060 8915 3080
rect 8991 3060 9011 3080
rect 9101 3060 9121 3080
rect 9197 3060 9217 3080
rect 9309 3060 9329 3080
rect 9405 3060 9425 3080
rect 9522 3060 9542 3080
rect 9618 3060 9638 3080
rect 10383 3084 10403 3104
rect 10479 3084 10499 3104
rect 10596 3084 10616 3104
rect 10692 3084 10712 3104
rect 10804 3084 10824 3104
rect 10900 3084 10920 3104
rect 11010 3084 11030 3104
rect 11106 3084 11126 3104
rect 15439 3125 15459 3145
rect 13870 3024 13890 3044
rect 13966 3024 13986 3044
rect 14076 3024 14096 3044
rect 14172 3024 14192 3044
rect 14284 3024 14304 3044
rect 14380 3024 14400 3044
rect 14497 3024 14517 3044
rect 15535 3125 15555 3145
rect 15652 3125 15672 3145
rect 15748 3125 15768 3145
rect 15860 3125 15880 3145
rect 15956 3125 15976 3145
rect 16066 3125 16086 3145
rect 16162 3125 16182 3145
rect 14593 3024 14613 3044
rect 18926 3065 18946 3085
rect 19022 3065 19042 3085
rect 19132 3065 19152 3085
rect 19228 3065 19248 3085
rect 19340 3065 19360 3085
rect 19436 3065 19456 3085
rect 19553 3065 19573 3085
rect 19649 3065 19669 3085
rect 1401 2810 1421 2830
rect 1497 2810 1517 2830
rect 1614 2810 1634 2830
rect 1710 2810 1730 2830
rect 1822 2810 1842 2830
rect 1918 2810 1938 2830
rect 2028 2810 2048 2830
rect 2124 2810 2144 2830
rect 6457 2851 6477 2871
rect 6553 2851 6573 2871
rect 6670 2851 6690 2871
rect 6766 2851 6786 2871
rect 6878 2851 6898 2871
rect 6974 2851 6994 2871
rect 7084 2851 7104 2871
rect 7180 2851 7200 2871
rect 2791 2739 2811 2759
rect 2887 2739 2907 2759
rect 2997 2739 3017 2759
rect 3093 2739 3113 2759
rect 3205 2739 3225 2759
rect 3301 2739 3321 2759
rect 3418 2739 3438 2759
rect 3514 2739 3534 2759
rect 7847 2780 7867 2800
rect 7943 2780 7963 2800
rect 8053 2780 8073 2800
rect 8149 2780 8169 2800
rect 8261 2780 8281 2800
rect 8357 2780 8377 2800
rect 8474 2780 8494 2800
rect 8570 2780 8590 2800
rect 11432 2815 11452 2835
rect 11528 2815 11548 2835
rect 11645 2815 11665 2835
rect 11741 2815 11761 2835
rect 11853 2815 11873 2835
rect 11949 2815 11969 2835
rect 12059 2815 12079 2835
rect 12155 2815 12175 2835
rect 16488 2856 16508 2876
rect 16584 2856 16604 2876
rect 16701 2856 16721 2876
rect 16797 2856 16817 2876
rect 16909 2856 16929 2876
rect 17005 2856 17025 2876
rect 17115 2856 17135 2876
rect 17211 2856 17231 2876
rect 12822 2744 12842 2764
rect 12918 2744 12938 2764
rect 13028 2744 13048 2764
rect 13124 2744 13144 2764
rect 13236 2744 13256 2764
rect 13332 2744 13352 2764
rect 13449 2744 13469 2764
rect 13545 2744 13565 2764
rect 17878 2785 17898 2805
rect 17974 2785 17994 2805
rect 18084 2785 18104 2805
rect 18180 2785 18200 2805
rect 18292 2785 18312 2805
rect 18388 2785 18408 2805
rect 18505 2785 18525 2805
rect 18601 2785 18621 2805
rect 353 2530 373 2550
rect 449 2530 469 2550
rect 566 2530 586 2550
rect 662 2530 682 2550
rect 774 2530 794 2550
rect 870 2530 890 2550
rect 980 2530 1000 2550
rect 1076 2530 1096 2550
rect 5409 2571 5429 2591
rect 3840 2470 3860 2490
rect 3936 2470 3956 2490
rect 4046 2470 4066 2490
rect 4142 2470 4162 2490
rect 4254 2470 4274 2490
rect 4350 2470 4370 2490
rect 4467 2470 4487 2490
rect 5505 2571 5525 2591
rect 5622 2571 5642 2591
rect 5718 2571 5738 2591
rect 5830 2571 5850 2591
rect 5926 2571 5946 2591
rect 6036 2571 6056 2591
rect 6132 2571 6152 2591
rect 4563 2470 4583 2490
rect 8896 2511 8916 2531
rect 8992 2511 9012 2531
rect 9102 2511 9122 2531
rect 9198 2511 9218 2531
rect 9310 2511 9330 2531
rect 9406 2511 9426 2531
rect 9523 2511 9543 2531
rect 9619 2511 9639 2531
rect 10384 2535 10404 2555
rect 10480 2535 10500 2555
rect 10597 2535 10617 2555
rect 10693 2535 10713 2555
rect 10805 2535 10825 2555
rect 10901 2535 10921 2555
rect 11011 2535 11031 2555
rect 11107 2535 11127 2555
rect 15440 2576 15460 2596
rect 1291 2286 1311 2306
rect 1387 2286 1407 2306
rect 1504 2286 1524 2306
rect 1600 2286 1620 2306
rect 1712 2286 1732 2306
rect 1808 2286 1828 2306
rect 1918 2286 1938 2306
rect 2014 2286 2034 2306
rect 6347 2327 6367 2347
rect 2901 2160 2921 2180
rect 2997 2160 3017 2180
rect 3107 2160 3127 2180
rect 3203 2160 3223 2180
rect 3315 2160 3335 2180
rect 3411 2160 3431 2180
rect 3528 2160 3548 2180
rect 6443 2327 6463 2347
rect 6560 2327 6580 2347
rect 6656 2327 6676 2347
rect 6768 2327 6788 2347
rect 6864 2327 6884 2347
rect 6974 2327 6994 2347
rect 13871 2475 13891 2495
rect 7070 2327 7090 2347
rect 13967 2475 13987 2495
rect 14077 2475 14097 2495
rect 14173 2475 14193 2495
rect 14285 2475 14305 2495
rect 14381 2475 14401 2495
rect 14498 2475 14518 2495
rect 15536 2576 15556 2596
rect 15653 2576 15673 2596
rect 15749 2576 15769 2596
rect 15861 2576 15881 2596
rect 15957 2576 15977 2596
rect 16067 2576 16087 2596
rect 16163 2576 16183 2596
rect 14594 2475 14614 2495
rect 18927 2516 18947 2536
rect 19023 2516 19043 2536
rect 19133 2516 19153 2536
rect 19229 2516 19249 2536
rect 19341 2516 19361 2536
rect 19437 2516 19457 2536
rect 19554 2516 19574 2536
rect 19650 2516 19670 2536
rect 3624 2160 3644 2180
rect 7957 2201 7977 2221
rect 8053 2201 8073 2221
rect 8163 2201 8183 2221
rect 8259 2201 8279 2221
rect 8371 2201 8391 2221
rect 8467 2201 8487 2221
rect 8584 2201 8604 2221
rect 11322 2291 11342 2311
rect 8680 2201 8700 2221
rect 11418 2291 11438 2311
rect 11535 2291 11555 2311
rect 11631 2291 11651 2311
rect 11743 2291 11763 2311
rect 11839 2291 11859 2311
rect 11949 2291 11969 2311
rect 12045 2291 12065 2311
rect 16378 2332 16398 2352
rect 352 1976 372 1996
rect 448 1976 468 1996
rect 565 1976 585 1996
rect 661 1976 681 1996
rect 773 1976 793 1996
rect 869 1976 889 1996
rect 979 1976 999 1996
rect 1075 1976 1095 1996
rect 5408 2017 5428 2037
rect 3839 1916 3859 1936
rect 3935 1916 3955 1936
rect 4045 1916 4065 1936
rect 4141 1916 4161 1936
rect 4253 1916 4273 1936
rect 4349 1916 4369 1936
rect 4466 1916 4486 1936
rect 5504 2017 5524 2037
rect 5621 2017 5641 2037
rect 5717 2017 5737 2037
rect 5829 2017 5849 2037
rect 5925 2017 5945 2037
rect 6035 2017 6055 2037
rect 12932 2165 12952 2185
rect 6131 2017 6151 2037
rect 13028 2165 13048 2185
rect 13138 2165 13158 2185
rect 13234 2165 13254 2185
rect 13346 2165 13366 2185
rect 13442 2165 13462 2185
rect 13559 2165 13579 2185
rect 16474 2332 16494 2352
rect 16591 2332 16611 2352
rect 16687 2332 16707 2352
rect 16799 2332 16819 2352
rect 16895 2332 16915 2352
rect 17005 2332 17025 2352
rect 17101 2332 17121 2352
rect 13655 2165 13675 2185
rect 17988 2206 18008 2226
rect 18084 2206 18104 2226
rect 18194 2206 18214 2226
rect 18290 2206 18310 2226
rect 18402 2206 18422 2226
rect 18498 2206 18518 2226
rect 18615 2206 18635 2226
rect 18711 2206 18731 2226
rect 4562 1916 4582 1936
rect 8895 1957 8915 1977
rect 8991 1957 9011 1977
rect 9101 1957 9121 1977
rect 9197 1957 9217 1977
rect 9309 1957 9329 1977
rect 9405 1957 9425 1977
rect 9522 1957 9542 1977
rect 9618 1957 9638 1977
rect 10383 1981 10403 2001
rect 10479 1981 10499 2001
rect 10596 1981 10616 2001
rect 10692 1981 10712 2001
rect 10804 1981 10824 2001
rect 10900 1981 10920 2001
rect 11010 1981 11030 2001
rect 11106 1981 11126 2001
rect 15439 2022 15459 2042
rect 13870 1921 13890 1941
rect 13966 1921 13986 1941
rect 14076 1921 14096 1941
rect 14172 1921 14192 1941
rect 14284 1921 14304 1941
rect 14380 1921 14400 1941
rect 14497 1921 14517 1941
rect 15535 2022 15555 2042
rect 15652 2022 15672 2042
rect 15748 2022 15768 2042
rect 15860 2022 15880 2042
rect 15956 2022 15976 2042
rect 16066 2022 16086 2042
rect 16162 2022 16182 2042
rect 14593 1921 14613 1941
rect 18926 1962 18946 1982
rect 19022 1962 19042 1982
rect 19132 1962 19152 1982
rect 19228 1962 19248 1982
rect 19340 1962 19360 1982
rect 19436 1962 19456 1982
rect 19553 1962 19573 1982
rect 19649 1962 19669 1982
rect 1432 1694 1452 1714
rect 1528 1694 1548 1714
rect 1645 1694 1665 1714
rect 1741 1694 1761 1714
rect 1853 1694 1873 1714
rect 1949 1694 1969 1714
rect 2059 1694 2079 1714
rect 2155 1694 2175 1714
rect 6488 1735 6508 1755
rect 2761 1649 2781 1669
rect 2857 1649 2877 1669
rect 2967 1649 2987 1669
rect 3063 1649 3083 1669
rect 3175 1649 3195 1669
rect 3271 1649 3291 1669
rect 3388 1649 3408 1669
rect 6584 1735 6604 1755
rect 6701 1735 6721 1755
rect 6797 1735 6817 1755
rect 6909 1735 6929 1755
rect 7005 1735 7025 1755
rect 7115 1735 7135 1755
rect 7211 1735 7231 1755
rect 3484 1649 3504 1669
rect 7817 1690 7837 1710
rect 7913 1690 7933 1710
rect 8023 1690 8043 1710
rect 8119 1690 8139 1710
rect 8231 1690 8251 1710
rect 8327 1690 8347 1710
rect 8444 1690 8464 1710
rect 8540 1690 8560 1710
rect 11463 1699 11483 1719
rect 11559 1699 11579 1719
rect 11676 1699 11696 1719
rect 11772 1699 11792 1719
rect 11884 1699 11904 1719
rect 11980 1699 12000 1719
rect 12090 1699 12110 1719
rect 12186 1699 12206 1719
rect 16519 1740 16539 1760
rect 12792 1654 12812 1674
rect 12888 1654 12908 1674
rect 12998 1654 13018 1674
rect 13094 1654 13114 1674
rect 13206 1654 13226 1674
rect 13302 1654 13322 1674
rect 13419 1654 13439 1674
rect 16615 1740 16635 1760
rect 16732 1740 16752 1760
rect 16828 1740 16848 1760
rect 16940 1740 16960 1760
rect 17036 1740 17056 1760
rect 17146 1740 17166 1760
rect 17242 1740 17262 1760
rect 13515 1654 13535 1674
rect 17848 1695 17868 1715
rect 17944 1695 17964 1715
rect 18054 1695 18074 1715
rect 18150 1695 18170 1715
rect 18262 1695 18282 1715
rect 18358 1695 18378 1715
rect 18475 1695 18495 1715
rect 18571 1695 18591 1715
rect 354 1427 374 1447
rect 450 1427 470 1447
rect 567 1427 587 1447
rect 663 1427 683 1447
rect 775 1427 795 1447
rect 871 1427 891 1447
rect 981 1427 1001 1447
rect 1077 1427 1097 1447
rect 5410 1468 5430 1488
rect 3841 1367 3861 1387
rect 3937 1367 3957 1387
rect 4047 1367 4067 1387
rect 4143 1367 4163 1387
rect 4255 1367 4275 1387
rect 4351 1367 4371 1387
rect 4468 1367 4488 1387
rect 5506 1468 5526 1488
rect 5623 1468 5643 1488
rect 5719 1468 5739 1488
rect 5831 1468 5851 1488
rect 5927 1468 5947 1488
rect 6037 1468 6057 1488
rect 6133 1468 6153 1488
rect 4564 1367 4584 1387
rect 8897 1408 8917 1428
rect 8993 1408 9013 1428
rect 9103 1408 9123 1428
rect 9199 1408 9219 1428
rect 9311 1408 9331 1428
rect 9407 1408 9427 1428
rect 9524 1408 9544 1428
rect 9620 1408 9640 1428
rect 10385 1432 10405 1452
rect 10481 1432 10501 1452
rect 10598 1432 10618 1452
rect 10694 1432 10714 1452
rect 10806 1432 10826 1452
rect 10902 1432 10922 1452
rect 11012 1432 11032 1452
rect 11108 1432 11128 1452
rect 15441 1473 15461 1493
rect 1292 1183 1312 1203
rect 1388 1183 1408 1203
rect 1505 1183 1525 1203
rect 1601 1183 1621 1203
rect 1713 1183 1733 1203
rect 1809 1183 1829 1203
rect 1919 1183 1939 1203
rect 2015 1183 2035 1203
rect 6348 1224 6368 1244
rect 2902 1057 2922 1077
rect 2998 1057 3018 1077
rect 3108 1057 3128 1077
rect 3204 1057 3224 1077
rect 3316 1057 3336 1077
rect 3412 1057 3432 1077
rect 3529 1057 3549 1077
rect 6444 1224 6464 1244
rect 6561 1224 6581 1244
rect 6657 1224 6677 1244
rect 6769 1224 6789 1244
rect 6865 1224 6885 1244
rect 6975 1224 6995 1244
rect 13872 1372 13892 1392
rect 7071 1224 7091 1244
rect 13968 1372 13988 1392
rect 14078 1372 14098 1392
rect 14174 1372 14194 1392
rect 14286 1372 14306 1392
rect 14382 1372 14402 1392
rect 14499 1372 14519 1392
rect 15537 1473 15557 1493
rect 15654 1473 15674 1493
rect 15750 1473 15770 1493
rect 15862 1473 15882 1493
rect 15958 1473 15978 1493
rect 16068 1473 16088 1493
rect 16164 1473 16184 1493
rect 14595 1372 14615 1392
rect 18928 1413 18948 1433
rect 19024 1413 19044 1433
rect 19134 1413 19154 1433
rect 19230 1413 19250 1433
rect 19342 1413 19362 1433
rect 19438 1413 19458 1433
rect 19555 1413 19575 1433
rect 19651 1413 19671 1433
rect 3625 1057 3645 1077
rect 7958 1098 7978 1118
rect 8054 1098 8074 1118
rect 8164 1098 8184 1118
rect 8260 1098 8280 1118
rect 8372 1098 8392 1118
rect 8468 1098 8488 1118
rect 8585 1098 8605 1118
rect 11323 1188 11343 1208
rect 8681 1098 8701 1118
rect 11419 1188 11439 1208
rect 11536 1188 11556 1208
rect 11632 1188 11652 1208
rect 11744 1188 11764 1208
rect 11840 1188 11860 1208
rect 11950 1188 11970 1208
rect 12046 1188 12066 1208
rect 16379 1229 16399 1249
rect 353 873 373 893
rect 449 873 469 893
rect 566 873 586 893
rect 662 873 682 893
rect 774 873 794 893
rect 870 873 890 893
rect 980 873 1000 893
rect 1076 873 1096 893
rect 5409 914 5429 934
rect 3840 813 3860 833
rect 3936 813 3956 833
rect 4046 813 4066 833
rect 4142 813 4162 833
rect 4254 813 4274 833
rect 4350 813 4370 833
rect 4467 813 4487 833
rect 5505 914 5525 934
rect 5622 914 5642 934
rect 5718 914 5738 934
rect 5830 914 5850 934
rect 5926 914 5946 934
rect 6036 914 6056 934
rect 12933 1062 12953 1082
rect 6132 914 6152 934
rect 13029 1062 13049 1082
rect 13139 1062 13159 1082
rect 13235 1062 13255 1082
rect 13347 1062 13367 1082
rect 13443 1062 13463 1082
rect 13560 1062 13580 1082
rect 16475 1229 16495 1249
rect 16592 1229 16612 1249
rect 16688 1229 16708 1249
rect 16800 1229 16820 1249
rect 16896 1229 16916 1249
rect 17006 1229 17026 1249
rect 17102 1229 17122 1249
rect 13656 1062 13676 1082
rect 17989 1103 18009 1123
rect 18085 1103 18105 1123
rect 18195 1103 18215 1123
rect 18291 1103 18311 1123
rect 18403 1103 18423 1123
rect 18499 1103 18519 1123
rect 18616 1103 18636 1123
rect 18712 1103 18732 1123
rect 4563 813 4583 833
rect 8896 854 8916 874
rect 8992 854 9012 874
rect 9102 854 9122 874
rect 9198 854 9218 874
rect 9310 854 9330 874
rect 9406 854 9426 874
rect 9523 854 9543 874
rect 9619 854 9639 874
rect 10384 878 10404 898
rect 10480 878 10500 898
rect 10597 878 10617 898
rect 10693 878 10713 898
rect 10805 878 10825 898
rect 10901 878 10921 898
rect 11011 878 11031 898
rect 11107 878 11127 898
rect 15440 919 15460 939
rect 13871 818 13891 838
rect 13967 818 13987 838
rect 14077 818 14097 838
rect 14173 818 14193 838
rect 14285 818 14305 838
rect 14381 818 14401 838
rect 14498 818 14518 838
rect 15536 919 15556 939
rect 15653 919 15673 939
rect 15749 919 15769 939
rect 15861 919 15881 939
rect 15957 919 15977 939
rect 16067 919 16087 939
rect 16163 919 16183 939
rect 14594 818 14614 838
rect 18927 859 18947 879
rect 19023 859 19043 879
rect 19133 859 19153 879
rect 19229 859 19249 879
rect 19341 859 19361 879
rect 19437 859 19457 879
rect 19554 859 19574 879
rect 19650 859 19670 879
rect 1600 314 1620 334
rect 1696 314 1716 334
rect 1813 314 1833 334
rect 1909 314 1929 334
rect 2021 314 2041 334
rect 2117 314 2137 334
rect 2227 314 2247 334
rect 6656 355 6676 375
rect 2323 314 2343 334
rect 4550 294 4570 314
rect 4646 294 4666 314
rect 4763 294 4783 314
rect 4859 294 4879 314
rect 4971 294 4991 314
rect 5067 294 5087 314
rect 5177 294 5197 314
rect 5273 294 5293 314
rect 6752 355 6772 375
rect 6869 355 6889 375
rect 6965 355 6985 375
rect 7077 355 7097 375
rect 7173 355 7193 375
rect 7283 355 7303 375
rect 7379 355 7399 375
rect 11631 319 11651 339
rect 11727 319 11747 339
rect 11844 319 11864 339
rect 11940 319 11960 339
rect 12052 319 12072 339
rect 12148 319 12168 339
rect 12258 319 12278 339
rect 16687 360 16707 380
rect 12354 319 12374 339
rect 14581 299 14601 319
rect 9484 178 9504 198
rect 9580 178 9600 198
rect 9697 178 9717 198
rect 9793 178 9813 198
rect 9905 178 9925 198
rect 10001 178 10021 198
rect 10111 178 10131 198
rect 14677 299 14697 319
rect 14794 299 14814 319
rect 14890 299 14910 319
rect 15002 299 15022 319
rect 15098 299 15118 319
rect 15208 299 15228 319
rect 15304 299 15324 319
rect 16783 360 16803 380
rect 16900 360 16920 380
rect 16996 360 17016 380
rect 17108 360 17128 380
rect 17204 360 17224 380
rect 17314 360 17334 380
rect 17410 360 17430 380
rect 10207 178 10227 198
<< psubdiff >>
rect 9457 9395 9568 9408
rect 4401 9354 4512 9369
rect 9457 9365 9499 9395
rect 9527 9365 9568 9395
rect 19488 9400 19599 9415
rect 4401 9324 4443 9354
rect 4471 9324 4512 9354
rect 9457 9351 9568 9365
rect 14432 9359 14543 9374
rect 19488 9370 19530 9400
rect 19558 9370 19599 9400
rect 4401 9310 4512 9324
rect 14432 9329 14474 9359
rect 14502 9329 14543 9359
rect 19488 9356 19599 9370
rect 14432 9315 14543 9329
rect 3462 9044 3573 9059
rect 3462 9014 3504 9044
rect 3532 9014 3573 9044
rect 3462 9000 3573 9014
rect 8518 9085 8629 9100
rect 8518 9055 8560 9085
rect 8588 9055 8629 9085
rect 8518 9041 8629 9055
rect 418 8932 529 8946
rect 418 8902 459 8932
rect 487 8902 529 8932
rect 418 8887 529 8902
rect 5474 8973 5585 8987
rect 5474 8943 5515 8973
rect 5543 8943 5585 8973
rect 5474 8928 5585 8943
rect 13493 9049 13604 9064
rect 13493 9019 13535 9049
rect 13563 9019 13604 9049
rect 13493 9005 13604 9019
rect 18549 9090 18660 9105
rect 18549 9060 18591 9090
rect 18619 9060 18660 9090
rect 18549 9046 18660 9060
rect 4400 8800 4511 8815
rect 4400 8770 4442 8800
rect 4470 8770 4511 8800
rect 10449 8937 10560 8951
rect 4400 8756 4511 8770
rect 10449 8907 10490 8937
rect 10518 8907 10560 8937
rect 10449 8892 10560 8907
rect 9456 8841 9567 8856
rect 9456 8811 9498 8841
rect 9526 8811 9567 8841
rect 15505 8978 15616 8992
rect 9456 8797 9567 8811
rect 15505 8948 15546 8978
rect 15574 8948 15616 8978
rect 15505 8933 15616 8948
rect 1356 8688 1467 8702
rect 1356 8658 1397 8688
rect 1425 8658 1467 8688
rect 1356 8643 1467 8658
rect 6412 8729 6523 8743
rect 6412 8699 6453 8729
rect 6481 8699 6523 8729
rect 3322 8533 3433 8548
rect 3322 8503 3364 8533
rect 3392 8503 3433 8533
rect 3322 8489 3433 8503
rect 6412 8684 6523 8699
rect 14431 8805 14542 8820
rect 14431 8775 14473 8805
rect 14501 8775 14542 8805
rect 14431 8761 14542 8775
rect 19487 8846 19598 8861
rect 19487 8816 19529 8846
rect 19557 8816 19598 8846
rect 19487 8802 19598 8816
rect 11387 8693 11498 8707
rect 8378 8574 8489 8589
rect 8378 8544 8420 8574
rect 8448 8544 8489 8574
rect 8378 8530 8489 8544
rect 11387 8663 11428 8693
rect 11456 8663 11498 8693
rect 11387 8648 11498 8663
rect 16443 8734 16554 8748
rect 16443 8704 16484 8734
rect 16512 8704 16554 8734
rect 13353 8538 13464 8553
rect 13353 8508 13395 8538
rect 13423 8508 13464 8538
rect 13353 8494 13464 8508
rect 16443 8689 16554 8704
rect 18409 8579 18520 8594
rect 18409 8549 18451 8579
rect 18479 8549 18520 8579
rect 18409 8535 18520 8549
rect 417 8378 528 8392
rect 417 8348 458 8378
rect 486 8348 528 8378
rect 417 8333 528 8348
rect 5473 8419 5584 8433
rect 5473 8389 5514 8419
rect 5542 8389 5584 8419
rect 5473 8374 5584 8389
rect 10448 8383 10559 8397
rect 4402 8251 4513 8266
rect 4402 8221 4444 8251
rect 4472 8221 4513 8251
rect 4402 8207 4513 8221
rect 10448 8353 10489 8383
rect 10517 8353 10559 8383
rect 10448 8338 10559 8353
rect 9458 8292 9569 8307
rect 9458 8262 9500 8292
rect 9528 8262 9569 8292
rect 15504 8424 15615 8438
rect 15504 8394 15545 8424
rect 15573 8394 15615 8424
rect 15504 8379 15615 8394
rect 9458 8248 9569 8262
rect 14433 8256 14544 8271
rect 14433 8226 14475 8256
rect 14503 8226 14544 8256
rect 14433 8212 14544 8226
rect 19489 8297 19600 8312
rect 19489 8267 19531 8297
rect 19559 8267 19600 8297
rect 19489 8253 19600 8267
rect 1497 8096 1608 8110
rect 1497 8066 1538 8096
rect 1566 8066 1608 8096
rect 1497 8051 1608 8066
rect 3463 7941 3574 7956
rect 6553 8137 6664 8151
rect 6553 8107 6594 8137
rect 6622 8107 6664 8137
rect 6553 8092 6664 8107
rect 3463 7911 3505 7941
rect 3533 7911 3574 7941
rect 3463 7897 3574 7911
rect 8519 7982 8630 7997
rect 8519 7952 8561 7982
rect 8589 7952 8630 7982
rect 11528 8101 11639 8115
rect 11528 8071 11569 8101
rect 11597 8071 11639 8101
rect 11528 8056 11639 8071
rect 8519 7938 8630 7952
rect 419 7829 530 7843
rect 419 7799 460 7829
rect 488 7799 530 7829
rect 419 7784 530 7799
rect 5475 7870 5586 7884
rect 5475 7840 5516 7870
rect 5544 7840 5586 7870
rect 5475 7825 5586 7840
rect 13494 7946 13605 7961
rect 16584 8142 16695 8156
rect 16584 8112 16625 8142
rect 16653 8112 16695 8142
rect 16584 8097 16695 8112
rect 13494 7916 13536 7946
rect 13564 7916 13605 7946
rect 13494 7902 13605 7916
rect 18550 7987 18661 8002
rect 18550 7957 18592 7987
rect 18620 7957 18661 7987
rect 18550 7943 18661 7957
rect 4401 7697 4512 7712
rect 4401 7667 4443 7697
rect 4471 7667 4512 7697
rect 10450 7834 10561 7848
rect 4401 7653 4512 7667
rect 10450 7804 10491 7834
rect 10519 7804 10561 7834
rect 10450 7789 10561 7804
rect 9457 7738 9568 7753
rect 9457 7708 9499 7738
rect 9527 7708 9568 7738
rect 15506 7875 15617 7889
rect 9457 7694 9568 7708
rect 15506 7845 15547 7875
rect 15575 7845 15617 7875
rect 15506 7830 15617 7845
rect 1357 7585 1468 7599
rect 1357 7555 1398 7585
rect 1426 7555 1468 7585
rect 1357 7540 1468 7555
rect 6413 7626 6524 7640
rect 6413 7596 6454 7626
rect 6482 7596 6524 7626
rect 3353 7417 3464 7432
rect 3353 7387 3395 7417
rect 3423 7387 3464 7417
rect 6413 7581 6524 7596
rect 14432 7702 14543 7717
rect 14432 7672 14474 7702
rect 14502 7672 14543 7702
rect 14432 7658 14543 7672
rect 19488 7743 19599 7758
rect 19488 7713 19530 7743
rect 19558 7713 19599 7743
rect 19488 7699 19599 7713
rect 11388 7590 11499 7604
rect 8409 7458 8520 7473
rect 8409 7428 8451 7458
rect 8479 7428 8520 7458
rect 11388 7560 11429 7590
rect 11457 7560 11499 7590
rect 11388 7545 11499 7560
rect 16444 7631 16555 7645
rect 16444 7601 16485 7631
rect 16513 7601 16555 7631
rect 8409 7414 8520 7428
rect 3353 7373 3464 7387
rect 418 7275 529 7289
rect 5474 7316 5585 7330
rect 13384 7422 13495 7437
rect 13384 7392 13426 7422
rect 13454 7392 13495 7422
rect 16444 7586 16555 7601
rect 18440 7463 18551 7478
rect 18440 7433 18482 7463
rect 18510 7433 18551 7463
rect 18440 7419 18551 7433
rect 13384 7378 13495 7392
rect 418 7245 459 7275
rect 487 7245 529 7275
rect 418 7231 529 7245
rect 5474 7286 5515 7316
rect 5543 7286 5585 7316
rect 5474 7272 5585 7286
rect 10449 7280 10560 7294
rect 15505 7321 15616 7335
rect 4402 7148 4513 7162
rect 4402 7118 4444 7148
rect 4472 7118 4513 7148
rect 10449 7250 10490 7280
rect 10518 7250 10560 7280
rect 10449 7236 10560 7250
rect 9458 7189 9569 7203
rect 9458 7159 9500 7189
rect 9528 7159 9569 7189
rect 15505 7291 15546 7321
rect 15574 7291 15616 7321
rect 15505 7277 15616 7291
rect 4402 7104 4513 7118
rect 9458 7145 9569 7159
rect 14433 7153 14544 7167
rect 14433 7123 14475 7153
rect 14503 7123 14544 7153
rect 19489 7194 19600 7208
rect 19489 7164 19531 7194
rect 19559 7164 19600 7194
rect 6523 7047 6634 7061
rect 1467 7006 1578 7020
rect 1467 6976 1508 7006
rect 1536 6976 1578 7006
rect 1467 6961 1578 6976
rect 3463 6838 3574 6853
rect 6523 7017 6564 7047
rect 6592 7017 6634 7047
rect 6523 7002 6634 7017
rect 14433 7109 14544 7123
rect 19489 7150 19600 7164
rect 16554 7052 16665 7066
rect 11498 7011 11609 7025
rect 3463 6808 3505 6838
rect 3533 6808 3574 6838
rect 3463 6794 3574 6808
rect 8519 6879 8630 6894
rect 8519 6849 8561 6879
rect 8589 6849 8630 6879
rect 11498 6981 11539 7011
rect 11567 6981 11609 7011
rect 11498 6966 11609 6981
rect 8519 6835 8630 6849
rect 419 6726 530 6740
rect 419 6696 460 6726
rect 488 6696 530 6726
rect 419 6681 530 6696
rect 5475 6767 5586 6781
rect 5475 6737 5516 6767
rect 5544 6737 5586 6767
rect 5475 6722 5586 6737
rect 13494 6843 13605 6858
rect 16554 7022 16595 7052
rect 16623 7022 16665 7052
rect 16554 7007 16665 7022
rect 13494 6813 13536 6843
rect 13564 6813 13605 6843
rect 13494 6799 13605 6813
rect 18550 6884 18661 6899
rect 18550 6854 18592 6884
rect 18620 6854 18661 6884
rect 18550 6840 18661 6854
rect 4401 6594 4512 6609
rect 4401 6564 4443 6594
rect 4471 6564 4512 6594
rect 10450 6731 10561 6745
rect 4401 6550 4512 6564
rect 10450 6701 10491 6731
rect 10519 6701 10561 6731
rect 10450 6686 10561 6701
rect 9457 6635 9568 6650
rect 9457 6605 9499 6635
rect 9527 6605 9568 6635
rect 15506 6772 15617 6786
rect 9457 6591 9568 6605
rect 15506 6742 15547 6772
rect 15575 6742 15617 6772
rect 15506 6727 15617 6742
rect 1357 6482 1468 6496
rect 1357 6452 1398 6482
rect 1426 6452 1468 6482
rect 1357 6437 1468 6452
rect 6413 6523 6524 6537
rect 6413 6493 6454 6523
rect 6482 6493 6524 6523
rect 3323 6327 3434 6342
rect 3323 6297 3365 6327
rect 3393 6297 3434 6327
rect 3323 6283 3434 6297
rect 6413 6478 6524 6493
rect 14432 6599 14543 6614
rect 14432 6569 14474 6599
rect 14502 6569 14543 6599
rect 14432 6555 14543 6569
rect 19488 6640 19599 6655
rect 19488 6610 19530 6640
rect 19558 6610 19599 6640
rect 19488 6596 19599 6610
rect 11388 6487 11499 6501
rect 8379 6368 8490 6383
rect 8379 6338 8421 6368
rect 8449 6338 8490 6368
rect 8379 6324 8490 6338
rect 11388 6457 11429 6487
rect 11457 6457 11499 6487
rect 11388 6442 11499 6457
rect 16444 6528 16555 6542
rect 16444 6498 16485 6528
rect 16513 6498 16555 6528
rect 13354 6332 13465 6347
rect 13354 6302 13396 6332
rect 13424 6302 13465 6332
rect 13354 6288 13465 6302
rect 16444 6483 16555 6498
rect 18410 6373 18521 6388
rect 18410 6343 18452 6373
rect 18480 6343 18521 6373
rect 18410 6329 18521 6343
rect 418 6172 529 6186
rect 418 6142 459 6172
rect 487 6142 529 6172
rect 418 6127 529 6142
rect 5474 6213 5585 6227
rect 5474 6183 5515 6213
rect 5543 6183 5585 6213
rect 5474 6168 5585 6183
rect 10449 6177 10560 6191
rect 4403 6045 4514 6060
rect 4403 6015 4445 6045
rect 4473 6015 4514 6045
rect 4403 6001 4514 6015
rect 10449 6147 10490 6177
rect 10518 6147 10560 6177
rect 10449 6132 10560 6147
rect 9459 6086 9570 6101
rect 9459 6056 9501 6086
rect 9529 6056 9570 6086
rect 15505 6218 15616 6232
rect 15505 6188 15546 6218
rect 15574 6188 15616 6218
rect 15505 6173 15616 6188
rect 9459 6042 9570 6056
rect 14434 6050 14545 6065
rect 14434 6020 14476 6050
rect 14504 6020 14545 6050
rect 14434 6006 14545 6020
rect 19490 6091 19601 6106
rect 19490 6061 19532 6091
rect 19560 6061 19601 6091
rect 19490 6047 19601 6061
rect 1498 5890 1609 5904
rect 1498 5860 1539 5890
rect 1567 5860 1609 5890
rect 1498 5845 1609 5860
rect 3464 5735 3575 5750
rect 6554 5931 6665 5945
rect 6554 5901 6595 5931
rect 6623 5901 6665 5931
rect 6554 5886 6665 5901
rect 3464 5705 3506 5735
rect 3534 5705 3575 5735
rect 3464 5691 3575 5705
rect 8520 5776 8631 5791
rect 8520 5746 8562 5776
rect 8590 5746 8631 5776
rect 11529 5895 11640 5909
rect 11529 5865 11570 5895
rect 11598 5865 11640 5895
rect 11529 5850 11640 5865
rect 8520 5732 8631 5746
rect 420 5623 531 5637
rect 420 5593 461 5623
rect 489 5593 531 5623
rect 420 5578 531 5593
rect 5476 5664 5587 5678
rect 5476 5634 5517 5664
rect 5545 5634 5587 5664
rect 5476 5619 5587 5634
rect 13495 5740 13606 5755
rect 16585 5936 16696 5950
rect 16585 5906 16626 5936
rect 16654 5906 16696 5936
rect 16585 5891 16696 5906
rect 13495 5710 13537 5740
rect 13565 5710 13606 5740
rect 13495 5696 13606 5710
rect 18551 5781 18662 5796
rect 18551 5751 18593 5781
rect 18621 5751 18662 5781
rect 18551 5737 18662 5751
rect 4402 5491 4513 5506
rect 4402 5461 4444 5491
rect 4472 5461 4513 5491
rect 10451 5628 10562 5642
rect 4402 5447 4513 5461
rect 10451 5598 10492 5628
rect 10520 5598 10562 5628
rect 10451 5583 10562 5598
rect 9458 5532 9569 5547
rect 9458 5502 9500 5532
rect 9528 5502 9569 5532
rect 15507 5669 15618 5683
rect 9458 5488 9569 5502
rect 15507 5639 15548 5669
rect 15576 5639 15618 5669
rect 15507 5624 15618 5639
rect 1358 5379 1469 5393
rect 1358 5349 1399 5379
rect 1427 5349 1469 5379
rect 1358 5334 1469 5349
rect 6414 5420 6525 5434
rect 6414 5390 6455 5420
rect 6483 5390 6525 5420
rect 3355 5205 3466 5220
rect 3355 5175 3397 5205
rect 3425 5175 3466 5205
rect 6414 5375 6525 5390
rect 14433 5496 14544 5511
rect 14433 5466 14475 5496
rect 14503 5466 14544 5496
rect 14433 5452 14544 5466
rect 19489 5537 19600 5552
rect 19489 5507 19531 5537
rect 19559 5507 19600 5537
rect 19489 5493 19600 5507
rect 11389 5384 11500 5398
rect 8411 5246 8522 5261
rect 8411 5216 8453 5246
rect 8481 5216 8522 5246
rect 11389 5354 11430 5384
rect 11458 5354 11500 5384
rect 11389 5339 11500 5354
rect 16445 5425 16556 5439
rect 16445 5395 16486 5425
rect 16514 5395 16556 5425
rect 3355 5161 3466 5175
rect 419 5069 530 5083
rect 419 5039 460 5069
rect 488 5039 530 5069
rect 419 5024 530 5039
rect 8411 5202 8522 5216
rect 5475 5110 5586 5124
rect 5475 5080 5516 5110
rect 5544 5080 5586 5110
rect 5475 5065 5586 5080
rect 13386 5210 13497 5225
rect 13386 5180 13428 5210
rect 13456 5180 13497 5210
rect 16445 5380 16556 5395
rect 18442 5251 18553 5266
rect 18442 5221 18484 5251
rect 18512 5221 18553 5251
rect 13386 5166 13497 5180
rect 10450 5074 10561 5088
rect 10450 5044 10491 5074
rect 10519 5044 10561 5074
rect 4403 4942 4514 4957
rect 4403 4912 4445 4942
rect 4473 4912 4514 4942
rect 4403 4898 4514 4912
rect 1467 4806 1578 4820
rect 10450 5029 10561 5044
rect 9459 4983 9570 4998
rect 18442 5207 18553 5221
rect 15506 5115 15617 5129
rect 15506 5085 15547 5115
rect 15575 5085 15617 5115
rect 15506 5070 15617 5085
rect 9459 4953 9501 4983
rect 9529 4953 9570 4983
rect 9459 4939 9570 4953
rect 6523 4847 6634 4861
rect 1467 4776 1508 4806
rect 1536 4776 1578 4806
rect 1467 4761 1578 4776
rect 3464 4632 3575 4647
rect 6523 4817 6564 4847
rect 6592 4817 6634 4847
rect 6523 4802 6634 4817
rect 14434 4947 14545 4962
rect 14434 4917 14476 4947
rect 14504 4917 14545 4947
rect 14434 4903 14545 4917
rect 11498 4811 11609 4825
rect 19490 4988 19601 5003
rect 19490 4958 19532 4988
rect 19560 4958 19601 4988
rect 19490 4944 19601 4958
rect 16554 4852 16665 4866
rect 3464 4602 3506 4632
rect 3534 4602 3575 4632
rect 3464 4588 3575 4602
rect 8520 4673 8631 4688
rect 8520 4643 8562 4673
rect 8590 4643 8631 4673
rect 11498 4781 11539 4811
rect 11567 4781 11609 4811
rect 11498 4766 11609 4781
rect 8520 4629 8631 4643
rect 420 4520 531 4534
rect 420 4490 461 4520
rect 489 4490 531 4520
rect 420 4475 531 4490
rect 5476 4561 5587 4575
rect 5476 4531 5517 4561
rect 5545 4531 5587 4561
rect 5476 4516 5587 4531
rect 13495 4637 13606 4652
rect 16554 4822 16595 4852
rect 16623 4822 16665 4852
rect 16554 4807 16665 4822
rect 13495 4607 13537 4637
rect 13565 4607 13606 4637
rect 13495 4593 13606 4607
rect 18551 4678 18662 4693
rect 18551 4648 18593 4678
rect 18621 4648 18662 4678
rect 18551 4634 18662 4648
rect 4402 4388 4513 4403
rect 4402 4358 4444 4388
rect 4472 4358 4513 4388
rect 10451 4525 10562 4539
rect 4402 4344 4513 4358
rect 10451 4495 10492 4525
rect 10520 4495 10562 4525
rect 10451 4480 10562 4495
rect 9458 4429 9569 4444
rect 9458 4399 9500 4429
rect 9528 4399 9569 4429
rect 15507 4566 15618 4580
rect 9458 4385 9569 4399
rect 15507 4536 15548 4566
rect 15576 4536 15618 4566
rect 15507 4521 15618 4536
rect 1358 4276 1469 4290
rect 1358 4246 1399 4276
rect 1427 4246 1469 4276
rect 1358 4231 1469 4246
rect 6414 4317 6525 4331
rect 6414 4287 6455 4317
rect 6483 4287 6525 4317
rect 3324 4121 3435 4136
rect 3324 4091 3366 4121
rect 3394 4091 3435 4121
rect 3324 4077 3435 4091
rect 6414 4272 6525 4287
rect 14433 4393 14544 4408
rect 14433 4363 14475 4393
rect 14503 4363 14544 4393
rect 14433 4349 14544 4363
rect 19489 4434 19600 4449
rect 19489 4404 19531 4434
rect 19559 4404 19600 4434
rect 19489 4390 19600 4404
rect 11389 4281 11500 4295
rect 8380 4162 8491 4177
rect 8380 4132 8422 4162
rect 8450 4132 8491 4162
rect 8380 4118 8491 4132
rect 11389 4251 11430 4281
rect 11458 4251 11500 4281
rect 11389 4236 11500 4251
rect 16445 4322 16556 4336
rect 16445 4292 16486 4322
rect 16514 4292 16556 4322
rect 13355 4126 13466 4141
rect 13355 4096 13397 4126
rect 13425 4096 13466 4126
rect 13355 4082 13466 4096
rect 16445 4277 16556 4292
rect 18411 4167 18522 4182
rect 18411 4137 18453 4167
rect 18481 4137 18522 4167
rect 18411 4123 18522 4137
rect 419 3966 530 3980
rect 419 3936 460 3966
rect 488 3936 530 3966
rect 419 3921 530 3936
rect 5475 4007 5586 4021
rect 5475 3977 5516 4007
rect 5544 3977 5586 4007
rect 5475 3962 5586 3977
rect 10450 3971 10561 3985
rect 4404 3839 4515 3854
rect 4404 3809 4446 3839
rect 4474 3809 4515 3839
rect 4404 3795 4515 3809
rect 10450 3941 10491 3971
rect 10519 3941 10561 3971
rect 10450 3926 10561 3941
rect 9460 3880 9571 3895
rect 9460 3850 9502 3880
rect 9530 3850 9571 3880
rect 15506 4012 15617 4026
rect 15506 3982 15547 4012
rect 15575 3982 15617 4012
rect 15506 3967 15617 3982
rect 9460 3836 9571 3850
rect 14435 3844 14546 3859
rect 14435 3814 14477 3844
rect 14505 3814 14546 3844
rect 14435 3800 14546 3814
rect 19491 3885 19602 3900
rect 19491 3855 19533 3885
rect 19561 3855 19602 3885
rect 19491 3841 19602 3855
rect 1499 3684 1610 3698
rect 1499 3654 1540 3684
rect 1568 3654 1610 3684
rect 1499 3639 1610 3654
rect 3465 3529 3576 3544
rect 6555 3725 6666 3739
rect 6555 3695 6596 3725
rect 6624 3695 6666 3725
rect 6555 3680 6666 3695
rect 3465 3499 3507 3529
rect 3535 3499 3576 3529
rect 3465 3485 3576 3499
rect 8521 3570 8632 3585
rect 8521 3540 8563 3570
rect 8591 3540 8632 3570
rect 11530 3689 11641 3703
rect 11530 3659 11571 3689
rect 11599 3659 11641 3689
rect 11530 3644 11641 3659
rect 8521 3526 8632 3540
rect 421 3417 532 3431
rect 421 3387 462 3417
rect 490 3387 532 3417
rect 421 3372 532 3387
rect 5477 3458 5588 3472
rect 5477 3428 5518 3458
rect 5546 3428 5588 3458
rect 5477 3413 5588 3428
rect 13496 3534 13607 3549
rect 16586 3730 16697 3744
rect 16586 3700 16627 3730
rect 16655 3700 16697 3730
rect 16586 3685 16697 3700
rect 13496 3504 13538 3534
rect 13566 3504 13607 3534
rect 13496 3490 13607 3504
rect 18552 3575 18663 3590
rect 18552 3545 18594 3575
rect 18622 3545 18663 3575
rect 18552 3531 18663 3545
rect 4403 3285 4514 3300
rect 4403 3255 4445 3285
rect 4473 3255 4514 3285
rect 10452 3422 10563 3436
rect 4403 3241 4514 3255
rect 10452 3392 10493 3422
rect 10521 3392 10563 3422
rect 10452 3377 10563 3392
rect 9459 3326 9570 3341
rect 9459 3296 9501 3326
rect 9529 3296 9570 3326
rect 15508 3463 15619 3477
rect 9459 3282 9570 3296
rect 15508 3433 15549 3463
rect 15577 3433 15619 3463
rect 15508 3418 15619 3433
rect 1359 3173 1470 3187
rect 1359 3143 1400 3173
rect 1428 3143 1470 3173
rect 1359 3128 1470 3143
rect 6415 3214 6526 3228
rect 6415 3184 6456 3214
rect 6484 3184 6526 3214
rect 3355 3005 3466 3020
rect 3355 2975 3397 3005
rect 3425 2975 3466 3005
rect 6415 3169 6526 3184
rect 14434 3290 14545 3305
rect 14434 3260 14476 3290
rect 14504 3260 14545 3290
rect 14434 3246 14545 3260
rect 19490 3331 19601 3346
rect 19490 3301 19532 3331
rect 19560 3301 19601 3331
rect 19490 3287 19601 3301
rect 11390 3178 11501 3192
rect 8411 3046 8522 3061
rect 8411 3016 8453 3046
rect 8481 3016 8522 3046
rect 11390 3148 11431 3178
rect 11459 3148 11501 3178
rect 11390 3133 11501 3148
rect 16446 3219 16557 3233
rect 16446 3189 16487 3219
rect 16515 3189 16557 3219
rect 8411 3002 8522 3016
rect 3355 2961 3466 2975
rect 420 2863 531 2877
rect 5476 2904 5587 2918
rect 13386 3010 13497 3025
rect 13386 2980 13428 3010
rect 13456 2980 13497 3010
rect 16446 3174 16557 3189
rect 18442 3051 18553 3066
rect 18442 3021 18484 3051
rect 18512 3021 18553 3051
rect 18442 3007 18553 3021
rect 13386 2966 13497 2980
rect 420 2833 461 2863
rect 489 2833 531 2863
rect 420 2819 531 2833
rect 5476 2874 5517 2904
rect 5545 2874 5587 2904
rect 5476 2860 5587 2874
rect 10451 2868 10562 2882
rect 15507 2909 15618 2923
rect 4404 2736 4515 2750
rect 4404 2706 4446 2736
rect 4474 2706 4515 2736
rect 10451 2838 10492 2868
rect 10520 2838 10562 2868
rect 10451 2824 10562 2838
rect 9460 2777 9571 2791
rect 9460 2747 9502 2777
rect 9530 2747 9571 2777
rect 15507 2879 15548 2909
rect 15576 2879 15618 2909
rect 15507 2865 15618 2879
rect 4404 2692 4515 2706
rect 9460 2733 9571 2747
rect 14435 2741 14546 2755
rect 14435 2711 14477 2741
rect 14505 2711 14546 2741
rect 19491 2782 19602 2796
rect 19491 2752 19533 2782
rect 19561 2752 19602 2782
rect 6525 2635 6636 2649
rect 1469 2594 1580 2608
rect 1469 2564 1510 2594
rect 1538 2564 1580 2594
rect 1469 2549 1580 2564
rect 3465 2426 3576 2441
rect 6525 2605 6566 2635
rect 6594 2605 6636 2635
rect 6525 2590 6636 2605
rect 14435 2697 14546 2711
rect 19491 2738 19602 2752
rect 16556 2640 16667 2654
rect 11500 2599 11611 2613
rect 3465 2396 3507 2426
rect 3535 2396 3576 2426
rect 3465 2382 3576 2396
rect 8521 2467 8632 2482
rect 8521 2437 8563 2467
rect 8591 2437 8632 2467
rect 11500 2569 11541 2599
rect 11569 2569 11611 2599
rect 11500 2554 11611 2569
rect 8521 2423 8632 2437
rect 421 2314 532 2328
rect 421 2284 462 2314
rect 490 2284 532 2314
rect 421 2269 532 2284
rect 5477 2355 5588 2369
rect 5477 2325 5518 2355
rect 5546 2325 5588 2355
rect 5477 2310 5588 2325
rect 13496 2431 13607 2446
rect 16556 2610 16597 2640
rect 16625 2610 16667 2640
rect 16556 2595 16667 2610
rect 13496 2401 13538 2431
rect 13566 2401 13607 2431
rect 13496 2387 13607 2401
rect 18552 2472 18663 2487
rect 18552 2442 18594 2472
rect 18622 2442 18663 2472
rect 18552 2428 18663 2442
rect 4403 2182 4514 2197
rect 4403 2152 4445 2182
rect 4473 2152 4514 2182
rect 10452 2319 10563 2333
rect 4403 2138 4514 2152
rect 10452 2289 10493 2319
rect 10521 2289 10563 2319
rect 10452 2274 10563 2289
rect 9459 2223 9570 2238
rect 9459 2193 9501 2223
rect 9529 2193 9570 2223
rect 15508 2360 15619 2374
rect 9459 2179 9570 2193
rect 15508 2330 15549 2360
rect 15577 2330 15619 2360
rect 15508 2315 15619 2330
rect 1359 2070 1470 2084
rect 1359 2040 1400 2070
rect 1428 2040 1470 2070
rect 1359 2025 1470 2040
rect 6415 2111 6526 2125
rect 6415 2081 6456 2111
rect 6484 2081 6526 2111
rect 3325 1915 3436 1930
rect 3325 1885 3367 1915
rect 3395 1885 3436 1915
rect 3325 1871 3436 1885
rect 6415 2066 6526 2081
rect 14434 2187 14545 2202
rect 14434 2157 14476 2187
rect 14504 2157 14545 2187
rect 14434 2143 14545 2157
rect 19490 2228 19601 2243
rect 19490 2198 19532 2228
rect 19560 2198 19601 2228
rect 19490 2184 19601 2198
rect 11390 2075 11501 2089
rect 8381 1956 8492 1971
rect 8381 1926 8423 1956
rect 8451 1926 8492 1956
rect 8381 1912 8492 1926
rect 11390 2045 11431 2075
rect 11459 2045 11501 2075
rect 11390 2030 11501 2045
rect 16446 2116 16557 2130
rect 16446 2086 16487 2116
rect 16515 2086 16557 2116
rect 13356 1920 13467 1935
rect 13356 1890 13398 1920
rect 13426 1890 13467 1920
rect 13356 1876 13467 1890
rect 16446 2071 16557 2086
rect 18412 1961 18523 1976
rect 18412 1931 18454 1961
rect 18482 1931 18523 1961
rect 18412 1917 18523 1931
rect 420 1760 531 1774
rect 420 1730 461 1760
rect 489 1730 531 1760
rect 420 1715 531 1730
rect 5476 1801 5587 1815
rect 5476 1771 5517 1801
rect 5545 1771 5587 1801
rect 5476 1756 5587 1771
rect 10451 1765 10562 1779
rect 4405 1633 4516 1648
rect 4405 1603 4447 1633
rect 4475 1603 4516 1633
rect 4405 1589 4516 1603
rect 10451 1735 10492 1765
rect 10520 1735 10562 1765
rect 10451 1720 10562 1735
rect 9461 1674 9572 1689
rect 9461 1644 9503 1674
rect 9531 1644 9572 1674
rect 15507 1806 15618 1820
rect 15507 1776 15548 1806
rect 15576 1776 15618 1806
rect 15507 1761 15618 1776
rect 9461 1630 9572 1644
rect 14436 1638 14547 1653
rect 14436 1608 14478 1638
rect 14506 1608 14547 1638
rect 14436 1594 14547 1608
rect 19492 1679 19603 1694
rect 19492 1649 19534 1679
rect 19562 1649 19603 1679
rect 19492 1635 19603 1649
rect 1500 1478 1611 1492
rect 1500 1448 1541 1478
rect 1569 1448 1611 1478
rect 1500 1433 1611 1448
rect 3466 1323 3577 1338
rect 6556 1519 6667 1533
rect 6556 1489 6597 1519
rect 6625 1489 6667 1519
rect 6556 1474 6667 1489
rect 3466 1293 3508 1323
rect 3536 1293 3577 1323
rect 3466 1279 3577 1293
rect 8522 1364 8633 1379
rect 8522 1334 8564 1364
rect 8592 1334 8633 1364
rect 11531 1483 11642 1497
rect 11531 1453 11572 1483
rect 11600 1453 11642 1483
rect 11531 1438 11642 1453
rect 8522 1320 8633 1334
rect 422 1211 533 1225
rect 422 1181 463 1211
rect 491 1181 533 1211
rect 422 1166 533 1181
rect 5478 1252 5589 1266
rect 5478 1222 5519 1252
rect 5547 1222 5589 1252
rect 5478 1207 5589 1222
rect 13497 1328 13608 1343
rect 16587 1524 16698 1538
rect 16587 1494 16628 1524
rect 16656 1494 16698 1524
rect 16587 1479 16698 1494
rect 13497 1298 13539 1328
rect 13567 1298 13608 1328
rect 13497 1284 13608 1298
rect 18553 1369 18664 1384
rect 18553 1339 18595 1369
rect 18623 1339 18664 1369
rect 18553 1325 18664 1339
rect 4404 1079 4515 1094
rect 4404 1049 4446 1079
rect 4474 1049 4515 1079
rect 10453 1216 10564 1230
rect 4404 1035 4515 1049
rect 10453 1186 10494 1216
rect 10522 1186 10564 1216
rect 10453 1171 10564 1186
rect 9460 1120 9571 1135
rect 9460 1090 9502 1120
rect 9530 1090 9571 1120
rect 15509 1257 15620 1271
rect 9460 1076 9571 1090
rect 15509 1227 15550 1257
rect 15578 1227 15620 1257
rect 15509 1212 15620 1227
rect 1360 967 1471 981
rect 1360 937 1401 967
rect 1429 937 1471 967
rect 1360 922 1471 937
rect 6416 1008 6527 1022
rect 6416 978 6457 1008
rect 6485 978 6527 1008
rect 6416 963 6527 978
rect 14435 1084 14546 1099
rect 14435 1054 14477 1084
rect 14505 1054 14546 1084
rect 14435 1040 14546 1054
rect 19491 1125 19602 1140
rect 19491 1095 19533 1125
rect 19561 1095 19602 1125
rect 19491 1081 19602 1095
rect 11391 972 11502 986
rect 11391 942 11432 972
rect 11460 942 11502 972
rect 11391 927 11502 942
rect 16447 1013 16558 1027
rect 16447 983 16488 1013
rect 16516 983 16558 1013
rect 16447 968 16558 983
rect 5477 698 5588 712
rect 421 657 532 671
rect 5477 668 5518 698
rect 5546 692 5588 698
rect 5546 668 5587 692
rect 15508 703 15619 717
rect 421 627 462 657
rect 490 651 532 657
rect 5477 653 5587 668
rect 10452 662 10563 676
rect 15508 673 15549 703
rect 15577 697 15619 703
rect 15577 673 15618 697
rect 490 627 531 651
rect 421 612 531 627
rect 10452 632 10493 662
rect 10521 656 10563 662
rect 15508 658 15618 673
rect 10521 632 10562 656
rect 10452 617 10562 632
rect 6724 139 6835 153
rect 1668 98 1779 112
rect 1668 68 1709 98
rect 1737 68 1779 98
rect 6724 109 6765 139
rect 6793 109 6835 139
rect 16755 144 16866 158
rect 6724 94 6835 109
rect 1668 53 1779 68
rect 4618 78 4729 92
rect 4618 48 4659 78
rect 4687 48 4729 78
rect 11699 103 11810 117
rect 11699 73 11740 103
rect 11768 73 11810 103
rect 16755 114 16796 144
rect 16824 114 16866 144
rect 16755 99 16866 114
rect 4618 33 4729 48
rect 11699 58 11810 73
rect 14649 83 14760 97
rect 14649 53 14690 83
rect 14718 53 14760 83
rect 14649 38 14760 53
rect 9552 -38 9663 -24
rect 9552 -68 9593 -38
rect 9621 -68 9663 -38
rect 9552 -83 9663 -68
<< nsubdiff >>
rect 5475 9320 5585 9334
rect 419 9279 529 9293
rect 419 9249 462 9279
rect 490 9249 529 9279
rect 419 9234 529 9249
rect 5475 9290 5518 9320
rect 5546 9290 5585 9320
rect 5475 9275 5585 9290
rect 15506 9325 15616 9339
rect 1357 9035 1467 9049
rect 1357 9005 1400 9035
rect 1428 9005 1467 9035
rect 1357 8990 1467 9005
rect 10450 9284 10560 9298
rect 10450 9254 10493 9284
rect 10521 9254 10560 9284
rect 10450 9239 10560 9254
rect 15506 9295 15549 9325
rect 15577 9295 15616 9325
rect 15506 9280 15616 9295
rect 6413 9076 6523 9090
rect 4401 9007 4511 9022
rect 6413 9046 6456 9076
rect 6484 9046 6523 9076
rect 6413 9031 6523 9046
rect 9457 9048 9567 9063
rect 9457 9018 9496 9048
rect 9524 9018 9567 9048
rect 4401 8977 4440 9007
rect 4468 8977 4511 9007
rect 4401 8963 4511 8977
rect 418 8725 528 8739
rect 9457 9004 9567 9018
rect 11388 9040 11498 9054
rect 11388 9010 11431 9040
rect 11459 9010 11498 9040
rect 11388 8995 11498 9010
rect 16444 9081 16554 9095
rect 14432 9012 14542 9027
rect 16444 9051 16487 9081
rect 16515 9051 16554 9081
rect 16444 9036 16554 9051
rect 19488 9053 19598 9068
rect 19488 9023 19527 9053
rect 19555 9023 19598 9053
rect 14432 8982 14471 9012
rect 14499 8982 14542 9012
rect 5474 8766 5584 8780
rect 14432 8968 14542 8982
rect 5474 8736 5517 8766
rect 5545 8736 5584 8766
rect 418 8695 461 8725
rect 489 8695 528 8725
rect 418 8680 528 8695
rect 3462 8697 3572 8712
rect 3462 8667 3501 8697
rect 3529 8667 3572 8697
rect 5474 8721 5584 8736
rect 3462 8653 3572 8667
rect 8518 8738 8628 8753
rect 8518 8708 8557 8738
rect 8585 8708 8628 8738
rect 8518 8694 8628 8708
rect 10449 8730 10559 8744
rect 19488 9009 19598 9023
rect 15505 8771 15615 8785
rect 15505 8741 15548 8771
rect 15576 8741 15615 8771
rect 10449 8700 10492 8730
rect 10520 8700 10559 8730
rect 10449 8685 10559 8700
rect 13493 8702 13603 8717
rect 13493 8672 13532 8702
rect 13560 8672 13603 8702
rect 15505 8726 15615 8741
rect 13493 8658 13603 8672
rect 1498 8443 1608 8457
rect 4400 8453 4510 8468
rect 1498 8413 1541 8443
rect 1569 8413 1608 8443
rect 1498 8398 1608 8413
rect 4400 8423 4439 8453
rect 4467 8423 4510 8453
rect 6554 8484 6664 8498
rect 9456 8494 9566 8509
rect 4400 8409 4510 8423
rect 6554 8454 6597 8484
rect 6625 8454 6664 8484
rect 6554 8439 6664 8454
rect 9456 8464 9495 8494
rect 9523 8464 9566 8494
rect 9456 8450 9566 8464
rect 18549 8743 18659 8758
rect 18549 8713 18588 8743
rect 18616 8713 18659 8743
rect 18549 8699 18659 8713
rect 11529 8448 11639 8462
rect 14431 8458 14541 8473
rect 11529 8418 11572 8448
rect 11600 8418 11639 8448
rect 11529 8403 11639 8418
rect 14431 8428 14470 8458
rect 14498 8428 14541 8458
rect 16585 8489 16695 8503
rect 19487 8499 19597 8514
rect 14431 8414 14541 8428
rect 16585 8459 16628 8489
rect 16656 8459 16695 8489
rect 16585 8444 16695 8459
rect 19487 8469 19526 8499
rect 19554 8469 19597 8499
rect 19487 8455 19597 8469
rect 420 8176 530 8190
rect 420 8146 463 8176
rect 491 8146 530 8176
rect 3322 8186 3432 8201
rect 3322 8156 3361 8186
rect 3389 8156 3432 8186
rect 5476 8217 5586 8231
rect 420 8131 530 8146
rect 3322 8142 3432 8156
rect 5476 8187 5519 8217
rect 5547 8187 5586 8217
rect 8378 8227 8488 8242
rect 8378 8197 8417 8227
rect 8445 8197 8488 8227
rect 5476 8172 5586 8187
rect 8378 8183 8488 8197
rect 1358 7932 1468 7946
rect 1358 7902 1401 7932
rect 1429 7902 1468 7932
rect 1358 7887 1468 7902
rect 10451 8181 10561 8195
rect 10451 8151 10494 8181
rect 10522 8151 10561 8181
rect 13353 8191 13463 8206
rect 13353 8161 13392 8191
rect 13420 8161 13463 8191
rect 15507 8222 15617 8236
rect 10451 8136 10561 8151
rect 13353 8147 13463 8161
rect 15507 8192 15550 8222
rect 15578 8192 15617 8222
rect 18409 8232 18519 8247
rect 18409 8202 18448 8232
rect 18476 8202 18519 8232
rect 15507 8177 15617 8192
rect 18409 8188 18519 8202
rect 6414 7973 6524 7987
rect 4402 7904 4512 7919
rect 6414 7943 6457 7973
rect 6485 7943 6524 7973
rect 6414 7928 6524 7943
rect 9458 7945 9568 7960
rect 9458 7915 9497 7945
rect 9525 7915 9568 7945
rect 4402 7874 4441 7904
rect 4469 7874 4512 7904
rect 4402 7860 4512 7874
rect 419 7622 529 7636
rect 9458 7901 9568 7915
rect 11389 7937 11499 7951
rect 11389 7907 11432 7937
rect 11460 7907 11499 7937
rect 11389 7892 11499 7907
rect 16445 7978 16555 7992
rect 14433 7909 14543 7924
rect 16445 7948 16488 7978
rect 16516 7948 16555 7978
rect 16445 7933 16555 7948
rect 19489 7950 19599 7965
rect 19489 7920 19528 7950
rect 19556 7920 19599 7950
rect 14433 7879 14472 7909
rect 14500 7879 14543 7909
rect 5475 7663 5585 7677
rect 14433 7865 14543 7879
rect 5475 7633 5518 7663
rect 5546 7633 5585 7663
rect 419 7592 462 7622
rect 490 7592 529 7622
rect 419 7577 529 7592
rect 3463 7594 3573 7609
rect 3463 7564 3502 7594
rect 3530 7564 3573 7594
rect 5475 7618 5585 7633
rect 3463 7550 3573 7564
rect 8519 7635 8629 7650
rect 8519 7605 8558 7635
rect 8586 7605 8629 7635
rect 8519 7591 8629 7605
rect 10450 7627 10560 7641
rect 19489 7906 19599 7920
rect 15506 7668 15616 7682
rect 15506 7638 15549 7668
rect 15577 7638 15616 7668
rect 10450 7597 10493 7627
rect 10521 7597 10560 7627
rect 10450 7582 10560 7597
rect 13494 7599 13604 7614
rect 13494 7569 13533 7599
rect 13561 7569 13604 7599
rect 15506 7623 15616 7638
rect 13494 7555 13604 7569
rect 1468 7353 1578 7367
rect 1468 7323 1511 7353
rect 1539 7323 1578 7353
rect 4401 7350 4511 7365
rect 1468 7308 1578 7323
rect 4401 7320 4440 7350
rect 4468 7320 4511 7350
rect 6524 7394 6634 7408
rect 6524 7364 6567 7394
rect 6595 7364 6634 7394
rect 9457 7391 9567 7406
rect 6524 7349 6634 7364
rect 4401 7306 4511 7320
rect 9457 7361 9496 7391
rect 9524 7361 9567 7391
rect 9457 7347 9567 7361
rect 18550 7640 18660 7655
rect 18550 7610 18589 7640
rect 18617 7610 18660 7640
rect 18550 7596 18660 7610
rect 11499 7358 11609 7372
rect 11499 7328 11542 7358
rect 11570 7328 11609 7358
rect 14432 7355 14542 7370
rect 11499 7313 11609 7328
rect 14432 7325 14471 7355
rect 14499 7325 14542 7355
rect 16555 7399 16665 7413
rect 16555 7369 16598 7399
rect 16626 7369 16665 7399
rect 19488 7396 19598 7411
rect 16555 7354 16665 7369
rect 14432 7311 14542 7325
rect 19488 7366 19527 7396
rect 19555 7366 19598 7396
rect 19488 7352 19598 7366
rect 420 7073 530 7087
rect 420 7043 463 7073
rect 491 7043 530 7073
rect 5476 7114 5586 7128
rect 3353 7070 3463 7085
rect 420 7028 530 7043
rect 3353 7040 3392 7070
rect 3420 7040 3463 7070
rect 3353 7026 3463 7040
rect 5476 7084 5519 7114
rect 5547 7084 5586 7114
rect 8409 7111 8519 7126
rect 5476 7069 5586 7084
rect 8409 7081 8448 7111
rect 8476 7081 8519 7111
rect 8409 7067 8519 7081
rect 1358 6829 1468 6843
rect 1358 6799 1401 6829
rect 1429 6799 1468 6829
rect 1358 6784 1468 6799
rect 10451 7078 10561 7092
rect 10451 7048 10494 7078
rect 10522 7048 10561 7078
rect 15507 7119 15617 7133
rect 13384 7075 13494 7090
rect 10451 7033 10561 7048
rect 13384 7045 13423 7075
rect 13451 7045 13494 7075
rect 13384 7031 13494 7045
rect 15507 7089 15550 7119
rect 15578 7089 15617 7119
rect 18440 7116 18550 7131
rect 15507 7074 15617 7089
rect 18440 7086 18479 7116
rect 18507 7086 18550 7116
rect 18440 7072 18550 7086
rect 6414 6870 6524 6884
rect 4402 6801 4512 6816
rect 6414 6840 6457 6870
rect 6485 6840 6524 6870
rect 6414 6825 6524 6840
rect 9458 6842 9568 6857
rect 9458 6812 9497 6842
rect 9525 6812 9568 6842
rect 4402 6771 4441 6801
rect 4469 6771 4512 6801
rect 4402 6757 4512 6771
rect 419 6519 529 6533
rect 9458 6798 9568 6812
rect 11389 6834 11499 6848
rect 11389 6804 11432 6834
rect 11460 6804 11499 6834
rect 11389 6789 11499 6804
rect 16445 6875 16555 6889
rect 14433 6806 14543 6821
rect 16445 6845 16488 6875
rect 16516 6845 16555 6875
rect 16445 6830 16555 6845
rect 19489 6847 19599 6862
rect 19489 6817 19528 6847
rect 19556 6817 19599 6847
rect 14433 6776 14472 6806
rect 14500 6776 14543 6806
rect 5475 6560 5585 6574
rect 14433 6762 14543 6776
rect 5475 6530 5518 6560
rect 5546 6530 5585 6560
rect 419 6489 462 6519
rect 490 6489 529 6519
rect 419 6474 529 6489
rect 3463 6491 3573 6506
rect 3463 6461 3502 6491
rect 3530 6461 3573 6491
rect 5475 6515 5585 6530
rect 3463 6447 3573 6461
rect 8519 6532 8629 6547
rect 8519 6502 8558 6532
rect 8586 6502 8629 6532
rect 8519 6488 8629 6502
rect 10450 6524 10560 6538
rect 19489 6803 19599 6817
rect 15506 6565 15616 6579
rect 15506 6535 15549 6565
rect 15577 6535 15616 6565
rect 10450 6494 10493 6524
rect 10521 6494 10560 6524
rect 10450 6479 10560 6494
rect 13494 6496 13604 6511
rect 13494 6466 13533 6496
rect 13561 6466 13604 6496
rect 15506 6520 15616 6535
rect 13494 6452 13604 6466
rect 1499 6237 1609 6251
rect 4401 6247 4511 6262
rect 1499 6207 1542 6237
rect 1570 6207 1609 6237
rect 1499 6192 1609 6207
rect 4401 6217 4440 6247
rect 4468 6217 4511 6247
rect 6555 6278 6665 6292
rect 9457 6288 9567 6303
rect 4401 6203 4511 6217
rect 6555 6248 6598 6278
rect 6626 6248 6665 6278
rect 6555 6233 6665 6248
rect 9457 6258 9496 6288
rect 9524 6258 9567 6288
rect 9457 6244 9567 6258
rect 18550 6537 18660 6552
rect 18550 6507 18589 6537
rect 18617 6507 18660 6537
rect 18550 6493 18660 6507
rect 11530 6242 11640 6256
rect 14432 6252 14542 6267
rect 11530 6212 11573 6242
rect 11601 6212 11640 6242
rect 11530 6197 11640 6212
rect 14432 6222 14471 6252
rect 14499 6222 14542 6252
rect 16586 6283 16696 6297
rect 19488 6293 19598 6308
rect 14432 6208 14542 6222
rect 16586 6253 16629 6283
rect 16657 6253 16696 6283
rect 16586 6238 16696 6253
rect 19488 6263 19527 6293
rect 19555 6263 19598 6293
rect 19488 6249 19598 6263
rect 421 5970 531 5984
rect 421 5940 464 5970
rect 492 5940 531 5970
rect 3323 5980 3433 5995
rect 3323 5950 3362 5980
rect 3390 5950 3433 5980
rect 5477 6011 5587 6025
rect 421 5925 531 5940
rect 3323 5936 3433 5950
rect 5477 5981 5520 6011
rect 5548 5981 5587 6011
rect 8379 6021 8489 6036
rect 8379 5991 8418 6021
rect 8446 5991 8489 6021
rect 5477 5966 5587 5981
rect 8379 5977 8489 5991
rect 1359 5726 1469 5740
rect 1359 5696 1402 5726
rect 1430 5696 1469 5726
rect 1359 5681 1469 5696
rect 10452 5975 10562 5989
rect 10452 5945 10495 5975
rect 10523 5945 10562 5975
rect 13354 5985 13464 6000
rect 13354 5955 13393 5985
rect 13421 5955 13464 5985
rect 15508 6016 15618 6030
rect 10452 5930 10562 5945
rect 13354 5941 13464 5955
rect 15508 5986 15551 6016
rect 15579 5986 15618 6016
rect 18410 6026 18520 6041
rect 18410 5996 18449 6026
rect 18477 5996 18520 6026
rect 15508 5971 15618 5986
rect 18410 5982 18520 5996
rect 6415 5767 6525 5781
rect 4403 5698 4513 5713
rect 6415 5737 6458 5767
rect 6486 5737 6525 5767
rect 6415 5722 6525 5737
rect 9459 5739 9569 5754
rect 9459 5709 9498 5739
rect 9526 5709 9569 5739
rect 4403 5668 4442 5698
rect 4470 5668 4513 5698
rect 4403 5654 4513 5668
rect 420 5416 530 5430
rect 9459 5695 9569 5709
rect 11390 5731 11500 5745
rect 11390 5701 11433 5731
rect 11461 5701 11500 5731
rect 11390 5686 11500 5701
rect 16446 5772 16556 5786
rect 14434 5703 14544 5718
rect 16446 5742 16489 5772
rect 16517 5742 16556 5772
rect 16446 5727 16556 5742
rect 19490 5744 19600 5759
rect 19490 5714 19529 5744
rect 19557 5714 19600 5744
rect 14434 5673 14473 5703
rect 14501 5673 14544 5703
rect 5476 5457 5586 5471
rect 14434 5659 14544 5673
rect 5476 5427 5519 5457
rect 5547 5427 5586 5457
rect 420 5386 463 5416
rect 491 5386 530 5416
rect 420 5371 530 5386
rect 3464 5388 3574 5403
rect 3464 5358 3503 5388
rect 3531 5358 3574 5388
rect 5476 5412 5586 5427
rect 3464 5344 3574 5358
rect 8520 5429 8630 5444
rect 8520 5399 8559 5429
rect 8587 5399 8630 5429
rect 8520 5385 8630 5399
rect 10451 5421 10561 5435
rect 19490 5700 19600 5714
rect 15507 5462 15617 5476
rect 15507 5432 15550 5462
rect 15578 5432 15617 5462
rect 10451 5391 10494 5421
rect 10522 5391 10561 5421
rect 10451 5376 10561 5391
rect 13495 5393 13605 5408
rect 13495 5363 13534 5393
rect 13562 5363 13605 5393
rect 15507 5417 15617 5432
rect 13495 5349 13605 5363
rect 1468 5153 1578 5167
rect 1468 5123 1511 5153
rect 1539 5123 1578 5153
rect 4402 5144 4512 5159
rect 1468 5108 1578 5123
rect 4402 5114 4441 5144
rect 4469 5114 4512 5144
rect 6524 5194 6634 5208
rect 6524 5164 6567 5194
rect 6595 5164 6634 5194
rect 9458 5185 9568 5200
rect 6524 5149 6634 5164
rect 4402 5100 4512 5114
rect 9458 5155 9497 5185
rect 9525 5155 9568 5185
rect 9458 5141 9568 5155
rect 18551 5434 18661 5449
rect 18551 5404 18590 5434
rect 18618 5404 18661 5434
rect 18551 5390 18661 5404
rect 11499 5158 11609 5172
rect 11499 5128 11542 5158
rect 11570 5128 11609 5158
rect 14433 5149 14543 5164
rect 11499 5113 11609 5128
rect 421 4867 531 4881
rect 421 4837 464 4867
rect 492 4837 531 4867
rect 5477 4908 5587 4922
rect 3355 4858 3465 4873
rect 421 4822 531 4837
rect 3355 4828 3394 4858
rect 3422 4828 3465 4858
rect 3355 4814 3465 4828
rect 5477 4878 5520 4908
rect 5548 4878 5587 4908
rect 14433 5119 14472 5149
rect 14500 5119 14543 5149
rect 16555 5199 16665 5213
rect 16555 5169 16598 5199
rect 16626 5169 16665 5199
rect 19489 5190 19599 5205
rect 16555 5154 16665 5169
rect 14433 5105 14543 5119
rect 19489 5160 19528 5190
rect 19556 5160 19599 5190
rect 19489 5146 19599 5160
rect 8411 4899 8521 4914
rect 5477 4863 5587 4878
rect 8411 4869 8450 4899
rect 8478 4869 8521 4899
rect 8411 4855 8521 4869
rect 1359 4623 1469 4637
rect 1359 4593 1402 4623
rect 1430 4593 1469 4623
rect 1359 4578 1469 4593
rect 10452 4872 10562 4886
rect 10452 4842 10495 4872
rect 10523 4842 10562 4872
rect 15508 4913 15618 4927
rect 13386 4863 13496 4878
rect 10452 4827 10562 4842
rect 13386 4833 13425 4863
rect 13453 4833 13496 4863
rect 13386 4819 13496 4833
rect 15508 4883 15551 4913
rect 15579 4883 15618 4913
rect 18442 4904 18552 4919
rect 15508 4868 15618 4883
rect 18442 4874 18481 4904
rect 18509 4874 18552 4904
rect 18442 4860 18552 4874
rect 6415 4664 6525 4678
rect 4403 4595 4513 4610
rect 6415 4634 6458 4664
rect 6486 4634 6525 4664
rect 6415 4619 6525 4634
rect 9459 4636 9569 4651
rect 9459 4606 9498 4636
rect 9526 4606 9569 4636
rect 4403 4565 4442 4595
rect 4470 4565 4513 4595
rect 4403 4551 4513 4565
rect 420 4313 530 4327
rect 9459 4592 9569 4606
rect 11390 4628 11500 4642
rect 11390 4598 11433 4628
rect 11461 4598 11500 4628
rect 11390 4583 11500 4598
rect 16446 4669 16556 4683
rect 14434 4600 14544 4615
rect 16446 4639 16489 4669
rect 16517 4639 16556 4669
rect 16446 4624 16556 4639
rect 19490 4641 19600 4656
rect 19490 4611 19529 4641
rect 19557 4611 19600 4641
rect 14434 4570 14473 4600
rect 14501 4570 14544 4600
rect 5476 4354 5586 4368
rect 14434 4556 14544 4570
rect 5476 4324 5519 4354
rect 5547 4324 5586 4354
rect 420 4283 463 4313
rect 491 4283 530 4313
rect 420 4268 530 4283
rect 3464 4285 3574 4300
rect 3464 4255 3503 4285
rect 3531 4255 3574 4285
rect 5476 4309 5586 4324
rect 3464 4241 3574 4255
rect 8520 4326 8630 4341
rect 8520 4296 8559 4326
rect 8587 4296 8630 4326
rect 8520 4282 8630 4296
rect 10451 4318 10561 4332
rect 19490 4597 19600 4611
rect 15507 4359 15617 4373
rect 15507 4329 15550 4359
rect 15578 4329 15617 4359
rect 10451 4288 10494 4318
rect 10522 4288 10561 4318
rect 10451 4273 10561 4288
rect 13495 4290 13605 4305
rect 13495 4260 13534 4290
rect 13562 4260 13605 4290
rect 15507 4314 15617 4329
rect 13495 4246 13605 4260
rect 1500 4031 1610 4045
rect 4402 4041 4512 4056
rect 1500 4001 1543 4031
rect 1571 4001 1610 4031
rect 1500 3986 1610 4001
rect 4402 4011 4441 4041
rect 4469 4011 4512 4041
rect 6556 4072 6666 4086
rect 9458 4082 9568 4097
rect 4402 3997 4512 4011
rect 6556 4042 6599 4072
rect 6627 4042 6666 4072
rect 6556 4027 6666 4042
rect 9458 4052 9497 4082
rect 9525 4052 9568 4082
rect 9458 4038 9568 4052
rect 18551 4331 18661 4346
rect 18551 4301 18590 4331
rect 18618 4301 18661 4331
rect 18551 4287 18661 4301
rect 11531 4036 11641 4050
rect 14433 4046 14543 4061
rect 11531 4006 11574 4036
rect 11602 4006 11641 4036
rect 11531 3991 11641 4006
rect 14433 4016 14472 4046
rect 14500 4016 14543 4046
rect 16587 4077 16697 4091
rect 19489 4087 19599 4102
rect 14433 4002 14543 4016
rect 16587 4047 16630 4077
rect 16658 4047 16697 4077
rect 16587 4032 16697 4047
rect 19489 4057 19528 4087
rect 19556 4057 19599 4087
rect 19489 4043 19599 4057
rect 422 3764 532 3778
rect 422 3734 465 3764
rect 493 3734 532 3764
rect 3324 3774 3434 3789
rect 3324 3744 3363 3774
rect 3391 3744 3434 3774
rect 5478 3805 5588 3819
rect 422 3719 532 3734
rect 3324 3730 3434 3744
rect 5478 3775 5521 3805
rect 5549 3775 5588 3805
rect 8380 3815 8490 3830
rect 8380 3785 8419 3815
rect 8447 3785 8490 3815
rect 5478 3760 5588 3775
rect 8380 3771 8490 3785
rect 1360 3520 1470 3534
rect 1360 3490 1403 3520
rect 1431 3490 1470 3520
rect 1360 3475 1470 3490
rect 10453 3769 10563 3783
rect 10453 3739 10496 3769
rect 10524 3739 10563 3769
rect 13355 3779 13465 3794
rect 13355 3749 13394 3779
rect 13422 3749 13465 3779
rect 15509 3810 15619 3824
rect 10453 3724 10563 3739
rect 13355 3735 13465 3749
rect 15509 3780 15552 3810
rect 15580 3780 15619 3810
rect 18411 3820 18521 3835
rect 18411 3790 18450 3820
rect 18478 3790 18521 3820
rect 15509 3765 15619 3780
rect 18411 3776 18521 3790
rect 6416 3561 6526 3575
rect 4404 3492 4514 3507
rect 6416 3531 6459 3561
rect 6487 3531 6526 3561
rect 6416 3516 6526 3531
rect 9460 3533 9570 3548
rect 9460 3503 9499 3533
rect 9527 3503 9570 3533
rect 4404 3462 4443 3492
rect 4471 3462 4514 3492
rect 4404 3448 4514 3462
rect 421 3210 531 3224
rect 9460 3489 9570 3503
rect 11391 3525 11501 3539
rect 11391 3495 11434 3525
rect 11462 3495 11501 3525
rect 11391 3480 11501 3495
rect 16447 3566 16557 3580
rect 14435 3497 14545 3512
rect 16447 3536 16490 3566
rect 16518 3536 16557 3566
rect 16447 3521 16557 3536
rect 19491 3538 19601 3553
rect 19491 3508 19530 3538
rect 19558 3508 19601 3538
rect 14435 3467 14474 3497
rect 14502 3467 14545 3497
rect 5477 3251 5587 3265
rect 14435 3453 14545 3467
rect 5477 3221 5520 3251
rect 5548 3221 5587 3251
rect 421 3180 464 3210
rect 492 3180 531 3210
rect 421 3165 531 3180
rect 3465 3182 3575 3197
rect 3465 3152 3504 3182
rect 3532 3152 3575 3182
rect 5477 3206 5587 3221
rect 3465 3138 3575 3152
rect 8521 3223 8631 3238
rect 8521 3193 8560 3223
rect 8588 3193 8631 3223
rect 8521 3179 8631 3193
rect 10452 3215 10562 3229
rect 19491 3494 19601 3508
rect 15508 3256 15618 3270
rect 15508 3226 15551 3256
rect 15579 3226 15618 3256
rect 10452 3185 10495 3215
rect 10523 3185 10562 3215
rect 10452 3170 10562 3185
rect 13496 3187 13606 3202
rect 13496 3157 13535 3187
rect 13563 3157 13606 3187
rect 15508 3211 15618 3226
rect 13496 3143 13606 3157
rect 1470 2941 1580 2955
rect 1470 2911 1513 2941
rect 1541 2911 1580 2941
rect 4403 2938 4513 2953
rect 1470 2896 1580 2911
rect 4403 2908 4442 2938
rect 4470 2908 4513 2938
rect 6526 2982 6636 2996
rect 6526 2952 6569 2982
rect 6597 2952 6636 2982
rect 9459 2979 9569 2994
rect 6526 2937 6636 2952
rect 4403 2894 4513 2908
rect 9459 2949 9498 2979
rect 9526 2949 9569 2979
rect 9459 2935 9569 2949
rect 18552 3228 18662 3243
rect 18552 3198 18591 3228
rect 18619 3198 18662 3228
rect 18552 3184 18662 3198
rect 11501 2946 11611 2960
rect 11501 2916 11544 2946
rect 11572 2916 11611 2946
rect 14434 2943 14544 2958
rect 11501 2901 11611 2916
rect 14434 2913 14473 2943
rect 14501 2913 14544 2943
rect 16557 2987 16667 3001
rect 16557 2957 16600 2987
rect 16628 2957 16667 2987
rect 19490 2984 19600 2999
rect 16557 2942 16667 2957
rect 14434 2899 14544 2913
rect 19490 2954 19529 2984
rect 19557 2954 19600 2984
rect 19490 2940 19600 2954
rect 422 2661 532 2675
rect 422 2631 465 2661
rect 493 2631 532 2661
rect 5478 2702 5588 2716
rect 3355 2658 3465 2673
rect 422 2616 532 2631
rect 3355 2628 3394 2658
rect 3422 2628 3465 2658
rect 3355 2614 3465 2628
rect 5478 2672 5521 2702
rect 5549 2672 5588 2702
rect 8411 2699 8521 2714
rect 5478 2657 5588 2672
rect 8411 2669 8450 2699
rect 8478 2669 8521 2699
rect 8411 2655 8521 2669
rect 1360 2417 1470 2431
rect 1360 2387 1403 2417
rect 1431 2387 1470 2417
rect 1360 2372 1470 2387
rect 10453 2666 10563 2680
rect 10453 2636 10496 2666
rect 10524 2636 10563 2666
rect 15509 2707 15619 2721
rect 13386 2663 13496 2678
rect 10453 2621 10563 2636
rect 13386 2633 13425 2663
rect 13453 2633 13496 2663
rect 13386 2619 13496 2633
rect 15509 2677 15552 2707
rect 15580 2677 15619 2707
rect 18442 2704 18552 2719
rect 15509 2662 15619 2677
rect 18442 2674 18481 2704
rect 18509 2674 18552 2704
rect 18442 2660 18552 2674
rect 6416 2458 6526 2472
rect 4404 2389 4514 2404
rect 6416 2428 6459 2458
rect 6487 2428 6526 2458
rect 6416 2413 6526 2428
rect 9460 2430 9570 2445
rect 9460 2400 9499 2430
rect 9527 2400 9570 2430
rect 4404 2359 4443 2389
rect 4471 2359 4514 2389
rect 4404 2345 4514 2359
rect 421 2107 531 2121
rect 9460 2386 9570 2400
rect 11391 2422 11501 2436
rect 11391 2392 11434 2422
rect 11462 2392 11501 2422
rect 11391 2377 11501 2392
rect 16447 2463 16557 2477
rect 14435 2394 14545 2409
rect 16447 2433 16490 2463
rect 16518 2433 16557 2463
rect 16447 2418 16557 2433
rect 19491 2435 19601 2450
rect 19491 2405 19530 2435
rect 19558 2405 19601 2435
rect 14435 2364 14474 2394
rect 14502 2364 14545 2394
rect 5477 2148 5587 2162
rect 14435 2350 14545 2364
rect 5477 2118 5520 2148
rect 5548 2118 5587 2148
rect 421 2077 464 2107
rect 492 2077 531 2107
rect 421 2062 531 2077
rect 3465 2079 3575 2094
rect 3465 2049 3504 2079
rect 3532 2049 3575 2079
rect 5477 2103 5587 2118
rect 3465 2035 3575 2049
rect 8521 2120 8631 2135
rect 8521 2090 8560 2120
rect 8588 2090 8631 2120
rect 8521 2076 8631 2090
rect 10452 2112 10562 2126
rect 19491 2391 19601 2405
rect 15508 2153 15618 2167
rect 15508 2123 15551 2153
rect 15579 2123 15618 2153
rect 10452 2082 10495 2112
rect 10523 2082 10562 2112
rect 10452 2067 10562 2082
rect 13496 2084 13606 2099
rect 13496 2054 13535 2084
rect 13563 2054 13606 2084
rect 15508 2108 15618 2123
rect 13496 2040 13606 2054
rect 1501 1825 1611 1839
rect 4403 1835 4513 1850
rect 1501 1795 1544 1825
rect 1572 1795 1611 1825
rect 1501 1780 1611 1795
rect 4403 1805 4442 1835
rect 4470 1805 4513 1835
rect 6557 1866 6667 1880
rect 9459 1876 9569 1891
rect 4403 1791 4513 1805
rect 6557 1836 6600 1866
rect 6628 1836 6667 1866
rect 6557 1821 6667 1836
rect 9459 1846 9498 1876
rect 9526 1846 9569 1876
rect 9459 1832 9569 1846
rect 18552 2125 18662 2140
rect 18552 2095 18591 2125
rect 18619 2095 18662 2125
rect 18552 2081 18662 2095
rect 11532 1830 11642 1844
rect 14434 1840 14544 1855
rect 11532 1800 11575 1830
rect 11603 1800 11642 1830
rect 11532 1785 11642 1800
rect 14434 1810 14473 1840
rect 14501 1810 14544 1840
rect 16588 1871 16698 1885
rect 19490 1881 19600 1896
rect 14434 1796 14544 1810
rect 16588 1841 16631 1871
rect 16659 1841 16698 1871
rect 16588 1826 16698 1841
rect 19490 1851 19529 1881
rect 19557 1851 19600 1881
rect 19490 1837 19600 1851
rect 423 1558 533 1572
rect 423 1528 466 1558
rect 494 1528 533 1558
rect 3325 1568 3435 1583
rect 3325 1538 3364 1568
rect 3392 1538 3435 1568
rect 5479 1599 5589 1613
rect 423 1513 533 1528
rect 3325 1524 3435 1538
rect 5479 1569 5522 1599
rect 5550 1569 5589 1599
rect 8381 1609 8491 1624
rect 8381 1579 8420 1609
rect 8448 1579 8491 1609
rect 5479 1554 5589 1569
rect 8381 1565 8491 1579
rect 1361 1314 1471 1328
rect 1361 1284 1404 1314
rect 1432 1284 1471 1314
rect 1361 1269 1471 1284
rect 10454 1563 10564 1577
rect 10454 1533 10497 1563
rect 10525 1533 10564 1563
rect 13356 1573 13466 1588
rect 13356 1543 13395 1573
rect 13423 1543 13466 1573
rect 15510 1604 15620 1618
rect 10454 1518 10564 1533
rect 13356 1529 13466 1543
rect 15510 1574 15553 1604
rect 15581 1574 15620 1604
rect 18412 1614 18522 1629
rect 18412 1584 18451 1614
rect 18479 1584 18522 1614
rect 15510 1559 15620 1574
rect 18412 1570 18522 1584
rect 6417 1355 6527 1369
rect 4405 1286 4515 1301
rect 6417 1325 6460 1355
rect 6488 1325 6527 1355
rect 6417 1310 6527 1325
rect 9461 1327 9571 1342
rect 9461 1297 9500 1327
rect 9528 1297 9571 1327
rect 4405 1256 4444 1286
rect 4472 1256 4515 1286
rect 4405 1242 4515 1256
rect 422 1004 532 1018
rect 9461 1283 9571 1297
rect 11392 1319 11502 1333
rect 11392 1289 11435 1319
rect 11463 1289 11502 1319
rect 11392 1274 11502 1289
rect 16448 1360 16558 1374
rect 14436 1291 14546 1306
rect 16448 1330 16491 1360
rect 16519 1330 16558 1360
rect 16448 1315 16558 1330
rect 19492 1332 19602 1347
rect 19492 1302 19531 1332
rect 19559 1302 19602 1332
rect 14436 1261 14475 1291
rect 14503 1261 14546 1291
rect 5478 1045 5588 1059
rect 14436 1247 14546 1261
rect 5478 1015 5521 1045
rect 5549 1015 5588 1045
rect 422 974 465 1004
rect 493 974 532 1004
rect 422 959 532 974
rect 3466 976 3576 991
rect 3466 946 3505 976
rect 3533 946 3576 976
rect 5478 1000 5588 1015
rect 3466 932 3576 946
rect 8522 1017 8632 1032
rect 8522 987 8561 1017
rect 8589 987 8632 1017
rect 8522 973 8632 987
rect 10453 1009 10563 1023
rect 19492 1288 19602 1302
rect 15509 1050 15619 1064
rect 15509 1020 15552 1050
rect 15580 1020 15619 1050
rect 10453 979 10496 1009
rect 10524 979 10563 1009
rect 10453 964 10563 979
rect 13497 981 13607 996
rect 13497 951 13536 981
rect 13564 951 13607 981
rect 15509 1005 15619 1020
rect 13497 937 13607 951
rect 4404 732 4514 747
rect 4404 702 4443 732
rect 4471 702 4514 732
rect 9460 773 9570 788
rect 9460 743 9499 773
rect 9527 743 9570 773
rect 9460 729 9570 743
rect 18553 1022 18663 1037
rect 18553 992 18592 1022
rect 18620 992 18663 1022
rect 18553 978 18663 992
rect 4404 688 4514 702
rect 14435 737 14545 752
rect 14435 707 14474 737
rect 14502 707 14545 737
rect 19491 778 19601 793
rect 19491 748 19530 778
rect 19558 748 19601 778
rect 19491 734 19601 748
rect 14435 693 14545 707
rect 6725 486 6835 500
rect 1669 445 1779 459
rect 1669 415 1712 445
rect 1740 415 1779 445
rect 6725 456 6768 486
rect 6796 456 6835 486
rect 16756 491 16866 505
rect 6725 441 6835 456
rect 11700 450 11810 464
rect 1669 400 1779 415
rect 4619 425 4729 439
rect 4619 395 4662 425
rect 4690 395 4729 425
rect 11700 420 11743 450
rect 11771 420 11810 450
rect 16756 461 16799 491
rect 16827 461 16866 491
rect 16756 446 16866 461
rect 4619 380 4729 395
rect 11700 405 11810 420
rect 14650 430 14760 444
rect 14650 400 14693 430
rect 14721 400 14760 430
rect 14650 385 14760 400
rect 9553 309 9663 323
rect 9553 279 9596 309
rect 9624 279 9663 309
rect 9553 264 9663 279
<< psubdiffcont >>
rect 9499 9365 9527 9395
rect 4443 9324 4471 9354
rect 19530 9370 19558 9400
rect 14474 9329 14502 9359
rect 3504 9014 3532 9044
rect 8560 9055 8588 9085
rect 459 8902 487 8932
rect 5515 8943 5543 8973
rect 13535 9019 13563 9049
rect 18591 9060 18619 9090
rect 4442 8770 4470 8800
rect 10490 8907 10518 8937
rect 9498 8811 9526 8841
rect 15546 8948 15574 8978
rect 1397 8658 1425 8688
rect 6453 8699 6481 8729
rect 3364 8503 3392 8533
rect 14473 8775 14501 8805
rect 19529 8816 19557 8846
rect 8420 8544 8448 8574
rect 11428 8663 11456 8693
rect 16484 8704 16512 8734
rect 13395 8508 13423 8538
rect 18451 8549 18479 8579
rect 458 8348 486 8378
rect 5514 8389 5542 8419
rect 4444 8221 4472 8251
rect 10489 8353 10517 8383
rect 9500 8262 9528 8292
rect 15545 8394 15573 8424
rect 14475 8226 14503 8256
rect 19531 8267 19559 8297
rect 1538 8066 1566 8096
rect 6594 8107 6622 8137
rect 3505 7911 3533 7941
rect 8561 7952 8589 7982
rect 11569 8071 11597 8101
rect 460 7799 488 7829
rect 5516 7840 5544 7870
rect 16625 8112 16653 8142
rect 13536 7916 13564 7946
rect 18592 7957 18620 7987
rect 4443 7667 4471 7697
rect 10491 7804 10519 7834
rect 9499 7708 9527 7738
rect 15547 7845 15575 7875
rect 1398 7555 1426 7585
rect 6454 7596 6482 7626
rect 3395 7387 3423 7417
rect 14474 7672 14502 7702
rect 19530 7713 19558 7743
rect 8451 7428 8479 7458
rect 11429 7560 11457 7590
rect 16485 7601 16513 7631
rect 13426 7392 13454 7422
rect 18482 7433 18510 7463
rect 459 7245 487 7275
rect 5515 7286 5543 7316
rect 4444 7118 4472 7148
rect 10490 7250 10518 7280
rect 9500 7159 9528 7189
rect 15546 7291 15574 7321
rect 14475 7123 14503 7153
rect 19531 7164 19559 7194
rect 1508 6976 1536 7006
rect 6564 7017 6592 7047
rect 3505 6808 3533 6838
rect 8561 6849 8589 6879
rect 11539 6981 11567 7011
rect 460 6696 488 6726
rect 5516 6737 5544 6767
rect 16595 7022 16623 7052
rect 13536 6813 13564 6843
rect 18592 6854 18620 6884
rect 4443 6564 4471 6594
rect 10491 6701 10519 6731
rect 9499 6605 9527 6635
rect 15547 6742 15575 6772
rect 1398 6452 1426 6482
rect 6454 6493 6482 6523
rect 3365 6297 3393 6327
rect 14474 6569 14502 6599
rect 19530 6610 19558 6640
rect 8421 6338 8449 6368
rect 11429 6457 11457 6487
rect 16485 6498 16513 6528
rect 13396 6302 13424 6332
rect 18452 6343 18480 6373
rect 459 6142 487 6172
rect 5515 6183 5543 6213
rect 4445 6015 4473 6045
rect 10490 6147 10518 6177
rect 9501 6056 9529 6086
rect 15546 6188 15574 6218
rect 14476 6020 14504 6050
rect 19532 6061 19560 6091
rect 1539 5860 1567 5890
rect 6595 5901 6623 5931
rect 3506 5705 3534 5735
rect 8562 5746 8590 5776
rect 11570 5865 11598 5895
rect 461 5593 489 5623
rect 5517 5634 5545 5664
rect 16626 5906 16654 5936
rect 13537 5710 13565 5740
rect 18593 5751 18621 5781
rect 4444 5461 4472 5491
rect 10492 5598 10520 5628
rect 9500 5502 9528 5532
rect 15548 5639 15576 5669
rect 1399 5349 1427 5379
rect 6455 5390 6483 5420
rect 3397 5175 3425 5205
rect 14475 5466 14503 5496
rect 19531 5507 19559 5537
rect 8453 5216 8481 5246
rect 11430 5354 11458 5384
rect 16486 5395 16514 5425
rect 460 5039 488 5069
rect 5516 5080 5544 5110
rect 13428 5180 13456 5210
rect 18484 5221 18512 5251
rect 10491 5044 10519 5074
rect 4445 4912 4473 4942
rect 15547 5085 15575 5115
rect 9501 4953 9529 4983
rect 1508 4776 1536 4806
rect 6564 4817 6592 4847
rect 14476 4917 14504 4947
rect 19532 4958 19560 4988
rect 3506 4602 3534 4632
rect 8562 4643 8590 4673
rect 11539 4781 11567 4811
rect 461 4490 489 4520
rect 5517 4531 5545 4561
rect 16595 4822 16623 4852
rect 13537 4607 13565 4637
rect 18593 4648 18621 4678
rect 4444 4358 4472 4388
rect 10492 4495 10520 4525
rect 9500 4399 9528 4429
rect 15548 4536 15576 4566
rect 1399 4246 1427 4276
rect 6455 4287 6483 4317
rect 3366 4091 3394 4121
rect 14475 4363 14503 4393
rect 19531 4404 19559 4434
rect 8422 4132 8450 4162
rect 11430 4251 11458 4281
rect 16486 4292 16514 4322
rect 13397 4096 13425 4126
rect 18453 4137 18481 4167
rect 460 3936 488 3966
rect 5516 3977 5544 4007
rect 4446 3809 4474 3839
rect 10491 3941 10519 3971
rect 9502 3850 9530 3880
rect 15547 3982 15575 4012
rect 14477 3814 14505 3844
rect 19533 3855 19561 3885
rect 1540 3654 1568 3684
rect 6596 3695 6624 3725
rect 3507 3499 3535 3529
rect 8563 3540 8591 3570
rect 11571 3659 11599 3689
rect 462 3387 490 3417
rect 5518 3428 5546 3458
rect 16627 3700 16655 3730
rect 13538 3504 13566 3534
rect 18594 3545 18622 3575
rect 4445 3255 4473 3285
rect 10493 3392 10521 3422
rect 9501 3296 9529 3326
rect 15549 3433 15577 3463
rect 1400 3143 1428 3173
rect 6456 3184 6484 3214
rect 3397 2975 3425 3005
rect 14476 3260 14504 3290
rect 19532 3301 19560 3331
rect 8453 3016 8481 3046
rect 11431 3148 11459 3178
rect 16487 3189 16515 3219
rect 13428 2980 13456 3010
rect 18484 3021 18512 3051
rect 461 2833 489 2863
rect 5517 2874 5545 2904
rect 4446 2706 4474 2736
rect 10492 2838 10520 2868
rect 9502 2747 9530 2777
rect 15548 2879 15576 2909
rect 14477 2711 14505 2741
rect 19533 2752 19561 2782
rect 1510 2564 1538 2594
rect 6566 2605 6594 2635
rect 3507 2396 3535 2426
rect 8563 2437 8591 2467
rect 11541 2569 11569 2599
rect 462 2284 490 2314
rect 5518 2325 5546 2355
rect 16597 2610 16625 2640
rect 13538 2401 13566 2431
rect 18594 2442 18622 2472
rect 4445 2152 4473 2182
rect 10493 2289 10521 2319
rect 9501 2193 9529 2223
rect 15549 2330 15577 2360
rect 1400 2040 1428 2070
rect 6456 2081 6484 2111
rect 3367 1885 3395 1915
rect 14476 2157 14504 2187
rect 19532 2198 19560 2228
rect 8423 1926 8451 1956
rect 11431 2045 11459 2075
rect 16487 2086 16515 2116
rect 13398 1890 13426 1920
rect 18454 1931 18482 1961
rect 461 1730 489 1760
rect 5517 1771 5545 1801
rect 4447 1603 4475 1633
rect 10492 1735 10520 1765
rect 9503 1644 9531 1674
rect 15548 1776 15576 1806
rect 14478 1608 14506 1638
rect 19534 1649 19562 1679
rect 1541 1448 1569 1478
rect 6597 1489 6625 1519
rect 3508 1293 3536 1323
rect 8564 1334 8592 1364
rect 11572 1453 11600 1483
rect 463 1181 491 1211
rect 5519 1222 5547 1252
rect 16628 1494 16656 1524
rect 13539 1298 13567 1328
rect 18595 1339 18623 1369
rect 4446 1049 4474 1079
rect 10494 1186 10522 1216
rect 9502 1090 9530 1120
rect 15550 1227 15578 1257
rect 1401 937 1429 967
rect 6457 978 6485 1008
rect 14477 1054 14505 1084
rect 19533 1095 19561 1125
rect 11432 942 11460 972
rect 16488 983 16516 1013
rect 5518 668 5546 698
rect 462 627 490 657
rect 15549 673 15577 703
rect 10493 632 10521 662
rect 1709 68 1737 98
rect 6765 109 6793 139
rect 4659 48 4687 78
rect 11740 73 11768 103
rect 16796 114 16824 144
rect 14690 53 14718 83
rect 9593 -68 9621 -38
<< nsubdiffcont >>
rect 462 9249 490 9279
rect 5518 9290 5546 9320
rect 1400 9005 1428 9035
rect 10493 9254 10521 9284
rect 15549 9295 15577 9325
rect 6456 9046 6484 9076
rect 9496 9018 9524 9048
rect 4440 8977 4468 9007
rect 11431 9010 11459 9040
rect 16487 9051 16515 9081
rect 19527 9023 19555 9053
rect 14471 8982 14499 9012
rect 5517 8736 5545 8766
rect 461 8695 489 8725
rect 3501 8667 3529 8697
rect 8557 8708 8585 8738
rect 15548 8741 15576 8771
rect 10492 8700 10520 8730
rect 13532 8672 13560 8702
rect 1541 8413 1569 8443
rect 4439 8423 4467 8453
rect 6597 8454 6625 8484
rect 9495 8464 9523 8494
rect 18588 8713 18616 8743
rect 11572 8418 11600 8448
rect 14470 8428 14498 8458
rect 16628 8459 16656 8489
rect 19526 8469 19554 8499
rect 463 8146 491 8176
rect 3361 8156 3389 8186
rect 5519 8187 5547 8217
rect 8417 8197 8445 8227
rect 1401 7902 1429 7932
rect 10494 8151 10522 8181
rect 13392 8161 13420 8191
rect 15550 8192 15578 8222
rect 18448 8202 18476 8232
rect 6457 7943 6485 7973
rect 9497 7915 9525 7945
rect 4441 7874 4469 7904
rect 11432 7907 11460 7937
rect 16488 7948 16516 7978
rect 19528 7920 19556 7950
rect 14472 7879 14500 7909
rect 5518 7633 5546 7663
rect 462 7592 490 7622
rect 3502 7564 3530 7594
rect 8558 7605 8586 7635
rect 15549 7638 15577 7668
rect 10493 7597 10521 7627
rect 13533 7569 13561 7599
rect 1511 7323 1539 7353
rect 4440 7320 4468 7350
rect 6567 7364 6595 7394
rect 9496 7361 9524 7391
rect 18589 7610 18617 7640
rect 11542 7328 11570 7358
rect 14471 7325 14499 7355
rect 16598 7369 16626 7399
rect 19527 7366 19555 7396
rect 463 7043 491 7073
rect 3392 7040 3420 7070
rect 5519 7084 5547 7114
rect 8448 7081 8476 7111
rect 1401 6799 1429 6829
rect 10494 7048 10522 7078
rect 13423 7045 13451 7075
rect 15550 7089 15578 7119
rect 18479 7086 18507 7116
rect 6457 6840 6485 6870
rect 9497 6812 9525 6842
rect 4441 6771 4469 6801
rect 11432 6804 11460 6834
rect 16488 6845 16516 6875
rect 19528 6817 19556 6847
rect 14472 6776 14500 6806
rect 5518 6530 5546 6560
rect 462 6489 490 6519
rect 3502 6461 3530 6491
rect 8558 6502 8586 6532
rect 15549 6535 15577 6565
rect 10493 6494 10521 6524
rect 13533 6466 13561 6496
rect 1542 6207 1570 6237
rect 4440 6217 4468 6247
rect 6598 6248 6626 6278
rect 9496 6258 9524 6288
rect 18589 6507 18617 6537
rect 11573 6212 11601 6242
rect 14471 6222 14499 6252
rect 16629 6253 16657 6283
rect 19527 6263 19555 6293
rect 464 5940 492 5970
rect 3362 5950 3390 5980
rect 5520 5981 5548 6011
rect 8418 5991 8446 6021
rect 1402 5696 1430 5726
rect 10495 5945 10523 5975
rect 13393 5955 13421 5985
rect 15551 5986 15579 6016
rect 18449 5996 18477 6026
rect 6458 5737 6486 5767
rect 9498 5709 9526 5739
rect 4442 5668 4470 5698
rect 11433 5701 11461 5731
rect 16489 5742 16517 5772
rect 19529 5714 19557 5744
rect 14473 5673 14501 5703
rect 5519 5427 5547 5457
rect 463 5386 491 5416
rect 3503 5358 3531 5388
rect 8559 5399 8587 5429
rect 15550 5432 15578 5462
rect 10494 5391 10522 5421
rect 13534 5363 13562 5393
rect 1511 5123 1539 5153
rect 4441 5114 4469 5144
rect 6567 5164 6595 5194
rect 9497 5155 9525 5185
rect 18590 5404 18618 5434
rect 11542 5128 11570 5158
rect 464 4837 492 4867
rect 3394 4828 3422 4858
rect 5520 4878 5548 4908
rect 14472 5119 14500 5149
rect 16598 5169 16626 5199
rect 19528 5160 19556 5190
rect 8450 4869 8478 4899
rect 1402 4593 1430 4623
rect 10495 4842 10523 4872
rect 13425 4833 13453 4863
rect 15551 4883 15579 4913
rect 18481 4874 18509 4904
rect 6458 4634 6486 4664
rect 9498 4606 9526 4636
rect 4442 4565 4470 4595
rect 11433 4598 11461 4628
rect 16489 4639 16517 4669
rect 19529 4611 19557 4641
rect 14473 4570 14501 4600
rect 5519 4324 5547 4354
rect 463 4283 491 4313
rect 3503 4255 3531 4285
rect 8559 4296 8587 4326
rect 15550 4329 15578 4359
rect 10494 4288 10522 4318
rect 13534 4260 13562 4290
rect 1543 4001 1571 4031
rect 4441 4011 4469 4041
rect 6599 4042 6627 4072
rect 9497 4052 9525 4082
rect 18590 4301 18618 4331
rect 11574 4006 11602 4036
rect 14472 4016 14500 4046
rect 16630 4047 16658 4077
rect 19528 4057 19556 4087
rect 465 3734 493 3764
rect 3363 3744 3391 3774
rect 5521 3775 5549 3805
rect 8419 3785 8447 3815
rect 1403 3490 1431 3520
rect 10496 3739 10524 3769
rect 13394 3749 13422 3779
rect 15552 3780 15580 3810
rect 18450 3790 18478 3820
rect 6459 3531 6487 3561
rect 9499 3503 9527 3533
rect 4443 3462 4471 3492
rect 11434 3495 11462 3525
rect 16490 3536 16518 3566
rect 19530 3508 19558 3538
rect 14474 3467 14502 3497
rect 5520 3221 5548 3251
rect 464 3180 492 3210
rect 3504 3152 3532 3182
rect 8560 3193 8588 3223
rect 15551 3226 15579 3256
rect 10495 3185 10523 3215
rect 13535 3157 13563 3187
rect 1513 2911 1541 2941
rect 4442 2908 4470 2938
rect 6569 2952 6597 2982
rect 9498 2949 9526 2979
rect 18591 3198 18619 3228
rect 11544 2916 11572 2946
rect 14473 2913 14501 2943
rect 16600 2957 16628 2987
rect 19529 2954 19557 2984
rect 465 2631 493 2661
rect 3394 2628 3422 2658
rect 5521 2672 5549 2702
rect 8450 2669 8478 2699
rect 1403 2387 1431 2417
rect 10496 2636 10524 2666
rect 13425 2633 13453 2663
rect 15552 2677 15580 2707
rect 18481 2674 18509 2704
rect 6459 2428 6487 2458
rect 9499 2400 9527 2430
rect 4443 2359 4471 2389
rect 11434 2392 11462 2422
rect 16490 2433 16518 2463
rect 19530 2405 19558 2435
rect 14474 2364 14502 2394
rect 5520 2118 5548 2148
rect 464 2077 492 2107
rect 3504 2049 3532 2079
rect 8560 2090 8588 2120
rect 15551 2123 15579 2153
rect 10495 2082 10523 2112
rect 13535 2054 13563 2084
rect 1544 1795 1572 1825
rect 4442 1805 4470 1835
rect 6600 1836 6628 1866
rect 9498 1846 9526 1876
rect 18591 2095 18619 2125
rect 11575 1800 11603 1830
rect 14473 1810 14501 1840
rect 16631 1841 16659 1871
rect 19529 1851 19557 1881
rect 466 1528 494 1558
rect 3364 1538 3392 1568
rect 5522 1569 5550 1599
rect 8420 1579 8448 1609
rect 1404 1284 1432 1314
rect 10497 1533 10525 1563
rect 13395 1543 13423 1573
rect 15553 1574 15581 1604
rect 18451 1584 18479 1614
rect 6460 1325 6488 1355
rect 9500 1297 9528 1327
rect 4444 1256 4472 1286
rect 11435 1289 11463 1319
rect 16491 1330 16519 1360
rect 19531 1302 19559 1332
rect 14475 1261 14503 1291
rect 5521 1015 5549 1045
rect 465 974 493 1004
rect 3505 946 3533 976
rect 8561 987 8589 1017
rect 15552 1020 15580 1050
rect 10496 979 10524 1009
rect 13536 951 13564 981
rect 4443 702 4471 732
rect 9499 743 9527 773
rect 18592 992 18620 1022
rect 14474 707 14502 737
rect 19530 748 19558 778
rect 1712 415 1740 445
rect 6768 456 6796 486
rect 4662 395 4690 425
rect 11743 420 11771 450
rect 16799 461 16827 491
rect 14693 400 14721 430
rect 9596 279 9624 309
<< poly >>
rect 3869 9269 3919 9285
rect 4077 9269 4127 9285
rect 4285 9269 4335 9285
rect 4498 9269 4548 9285
rect 8925 9310 8975 9326
rect 9133 9310 9183 9326
rect 9341 9310 9391 9326
rect 9554 9310 9604 9326
rect 5438 9247 5488 9260
rect 5651 9247 5701 9260
rect 5859 9247 5909 9260
rect 6067 9247 6117 9260
rect 382 9206 432 9219
rect 595 9206 645 9219
rect 803 9206 853 9219
rect 1011 9206 1061 9219
rect 3869 9202 3919 9227
rect 3869 9176 3875 9202
rect 3901 9176 3919 9202
rect 3869 9150 3919 9176
rect 4077 9198 4127 9227
rect 4077 9174 4091 9198
rect 4115 9174 4127 9198
rect 4077 9150 4127 9174
rect 4285 9203 4335 9227
rect 4285 9179 4300 9203
rect 4324 9179 4335 9203
rect 4285 9150 4335 9179
rect 4498 9198 4548 9227
rect 4498 9178 4515 9198
rect 4535 9178 4548 9198
rect 4498 9150 4548 9178
rect 382 9078 432 9106
rect 382 9058 395 9078
rect 415 9058 432 9078
rect 382 9029 432 9058
rect 595 9077 645 9106
rect 595 9053 606 9077
rect 630 9053 645 9077
rect 595 9029 645 9053
rect 803 9082 853 9106
rect 803 9058 815 9082
rect 839 9058 853 9082
rect 803 9029 853 9058
rect 1011 9080 1061 9106
rect 1011 9054 1029 9080
rect 1055 9054 1061 9080
rect 1011 9029 1061 9054
rect 8925 9243 8975 9268
rect 8925 9217 8931 9243
rect 8957 9217 8975 9243
rect 8925 9191 8975 9217
rect 9133 9239 9183 9268
rect 9133 9215 9147 9239
rect 9171 9215 9183 9239
rect 9133 9191 9183 9215
rect 9341 9244 9391 9268
rect 9341 9220 9356 9244
rect 9380 9220 9391 9244
rect 9341 9191 9391 9220
rect 9554 9239 9604 9268
rect 9554 9219 9571 9239
rect 9591 9219 9604 9239
rect 13900 9274 13950 9290
rect 14108 9274 14158 9290
rect 14316 9274 14366 9290
rect 14529 9274 14579 9290
rect 18956 9315 19006 9331
rect 19164 9315 19214 9331
rect 19372 9315 19422 9331
rect 19585 9315 19635 9331
rect 15469 9252 15519 9265
rect 15682 9252 15732 9265
rect 15890 9252 15940 9265
rect 16098 9252 16148 9265
rect 9554 9191 9604 9219
rect 10413 9211 10463 9224
rect 10626 9211 10676 9224
rect 10834 9211 10884 9224
rect 11042 9211 11092 9224
rect 5438 9119 5488 9147
rect 5438 9099 5451 9119
rect 5471 9099 5488 9119
rect 3869 9037 3919 9050
rect 4077 9037 4127 9050
rect 4285 9037 4335 9050
rect 4498 9037 4548 9050
rect 5438 9070 5488 9099
rect 5651 9118 5701 9147
rect 5651 9094 5662 9118
rect 5686 9094 5701 9118
rect 5651 9070 5701 9094
rect 5859 9123 5909 9147
rect 5859 9099 5871 9123
rect 5895 9099 5909 9123
rect 5859 9070 5909 9099
rect 6067 9121 6117 9147
rect 6067 9095 6085 9121
rect 6111 9095 6117 9121
rect 6067 9070 6117 9095
rect 8925 9078 8975 9091
rect 9133 9078 9183 9091
rect 9341 9078 9391 9091
rect 9554 9078 9604 9091
rect 13900 9207 13950 9232
rect 13900 9181 13906 9207
rect 13932 9181 13950 9207
rect 13900 9155 13950 9181
rect 14108 9203 14158 9232
rect 14108 9179 14122 9203
rect 14146 9179 14158 9203
rect 14108 9155 14158 9179
rect 14316 9208 14366 9232
rect 14316 9184 14331 9208
rect 14355 9184 14366 9208
rect 14316 9155 14366 9184
rect 14529 9203 14579 9232
rect 14529 9183 14546 9203
rect 14566 9183 14579 9203
rect 14529 9155 14579 9183
rect 10413 9083 10463 9111
rect 5438 9012 5488 9028
rect 5651 9012 5701 9028
rect 5859 9012 5909 9028
rect 6067 9012 6117 9028
rect 10413 9063 10426 9083
rect 10446 9063 10463 9083
rect 382 8971 432 8987
rect 595 8971 645 8987
rect 803 8971 853 8987
rect 1011 8971 1061 8987
rect 6376 9003 6426 9016
rect 6589 9003 6639 9016
rect 6797 9003 6847 9016
rect 7005 9003 7055 9016
rect 1320 8962 1370 8975
rect 1533 8962 1583 8975
rect 1741 8962 1791 8975
rect 1949 8962 1999 8975
rect 2930 8959 2980 8975
rect 3138 8959 3188 8975
rect 3346 8959 3396 8975
rect 3559 8959 3609 8975
rect 2930 8892 2980 8917
rect 2930 8866 2936 8892
rect 2962 8866 2980 8892
rect 1320 8834 1370 8862
rect 1320 8814 1333 8834
rect 1353 8814 1370 8834
rect 1320 8785 1370 8814
rect 1533 8833 1583 8862
rect 1533 8809 1544 8833
rect 1568 8809 1583 8833
rect 1533 8785 1583 8809
rect 1741 8838 1791 8862
rect 1741 8814 1753 8838
rect 1777 8814 1791 8838
rect 1741 8785 1791 8814
rect 1949 8836 1999 8862
rect 2930 8840 2980 8866
rect 3138 8888 3188 8917
rect 3138 8864 3152 8888
rect 3176 8864 3188 8888
rect 3138 8840 3188 8864
rect 3346 8893 3396 8917
rect 3346 8869 3361 8893
rect 3385 8869 3396 8893
rect 3346 8840 3396 8869
rect 3559 8888 3609 8917
rect 3559 8868 3576 8888
rect 3596 8868 3609 8888
rect 3559 8840 3609 8868
rect 1949 8810 1967 8836
rect 1993 8810 1999 8836
rect 1949 8785 1999 8810
rect 1320 8727 1370 8743
rect 1533 8727 1583 8743
rect 1741 8727 1791 8743
rect 1949 8727 1999 8743
rect 7986 9000 8036 9016
rect 8194 9000 8244 9016
rect 8402 9000 8452 9016
rect 8615 9000 8665 9016
rect 10413 9034 10463 9063
rect 10626 9082 10676 9111
rect 10626 9058 10637 9082
rect 10661 9058 10676 9082
rect 10626 9034 10676 9058
rect 10834 9087 10884 9111
rect 10834 9063 10846 9087
rect 10870 9063 10884 9087
rect 10834 9034 10884 9063
rect 11042 9085 11092 9111
rect 11042 9059 11060 9085
rect 11086 9059 11092 9085
rect 11042 9034 11092 9059
rect 18956 9248 19006 9273
rect 18956 9222 18962 9248
rect 18988 9222 19006 9248
rect 18956 9196 19006 9222
rect 19164 9244 19214 9273
rect 19164 9220 19178 9244
rect 19202 9220 19214 9244
rect 19164 9196 19214 9220
rect 19372 9249 19422 9273
rect 19372 9225 19387 9249
rect 19411 9225 19422 9249
rect 19372 9196 19422 9225
rect 19585 9244 19635 9273
rect 19585 9224 19602 9244
rect 19622 9224 19635 9244
rect 19585 9196 19635 9224
rect 15469 9124 15519 9152
rect 15469 9104 15482 9124
rect 15502 9104 15519 9124
rect 13900 9042 13950 9055
rect 14108 9042 14158 9055
rect 14316 9042 14366 9055
rect 14529 9042 14579 9055
rect 15469 9075 15519 9104
rect 15682 9123 15732 9152
rect 15682 9099 15693 9123
rect 15717 9099 15732 9123
rect 15682 9075 15732 9099
rect 15890 9128 15940 9152
rect 15890 9104 15902 9128
rect 15926 9104 15940 9128
rect 15890 9075 15940 9104
rect 16098 9126 16148 9152
rect 16098 9100 16116 9126
rect 16142 9100 16148 9126
rect 16098 9075 16148 9100
rect 18956 9083 19006 9096
rect 19164 9083 19214 9096
rect 19372 9083 19422 9096
rect 19585 9083 19635 9096
rect 15469 9017 15519 9033
rect 15682 9017 15732 9033
rect 15890 9017 15940 9033
rect 16098 9017 16148 9033
rect 10413 8976 10463 8992
rect 10626 8976 10676 8992
rect 10834 8976 10884 8992
rect 11042 8976 11092 8992
rect 16407 9008 16457 9021
rect 16620 9008 16670 9021
rect 16828 9008 16878 9021
rect 17036 9008 17086 9021
rect 7986 8933 8036 8958
rect 7986 8907 7992 8933
rect 8018 8907 8036 8933
rect 6376 8875 6426 8903
rect 6376 8855 6389 8875
rect 6409 8855 6426 8875
rect 6376 8826 6426 8855
rect 6589 8874 6639 8903
rect 6589 8850 6600 8874
rect 6624 8850 6639 8874
rect 6589 8826 6639 8850
rect 6797 8879 6847 8903
rect 6797 8855 6809 8879
rect 6833 8855 6847 8879
rect 6797 8826 6847 8855
rect 7005 8877 7055 8903
rect 7986 8881 8036 8907
rect 8194 8929 8244 8958
rect 8194 8905 8208 8929
rect 8232 8905 8244 8929
rect 8194 8881 8244 8905
rect 8402 8934 8452 8958
rect 8402 8910 8417 8934
rect 8441 8910 8452 8934
rect 8402 8881 8452 8910
rect 8615 8929 8665 8958
rect 11351 8967 11401 8980
rect 11564 8967 11614 8980
rect 11772 8967 11822 8980
rect 11980 8967 12030 8980
rect 8615 8909 8632 8929
rect 8652 8909 8665 8929
rect 8615 8881 8665 8909
rect 7005 8851 7023 8877
rect 7049 8851 7055 8877
rect 7005 8826 7055 8851
rect 6376 8768 6426 8784
rect 6589 8768 6639 8784
rect 6797 8768 6847 8784
rect 7005 8768 7055 8784
rect 12961 8964 13011 8980
rect 13169 8964 13219 8980
rect 13377 8964 13427 8980
rect 13590 8964 13640 8980
rect 12961 8897 13011 8922
rect 12961 8871 12967 8897
rect 12993 8871 13011 8897
rect 11351 8839 11401 8867
rect 11351 8819 11364 8839
rect 11384 8819 11401 8839
rect 7986 8768 8036 8781
rect 8194 8768 8244 8781
rect 8402 8768 8452 8781
rect 8615 8768 8665 8781
rect 11351 8790 11401 8819
rect 11564 8838 11614 8867
rect 11564 8814 11575 8838
rect 11599 8814 11614 8838
rect 11564 8790 11614 8814
rect 11772 8843 11822 8867
rect 11772 8819 11784 8843
rect 11808 8819 11822 8843
rect 11772 8790 11822 8819
rect 11980 8841 12030 8867
rect 12961 8845 13011 8871
rect 13169 8893 13219 8922
rect 13169 8869 13183 8893
rect 13207 8869 13219 8893
rect 13169 8845 13219 8869
rect 13377 8898 13427 8922
rect 13377 8874 13392 8898
rect 13416 8874 13427 8898
rect 13377 8845 13427 8874
rect 13590 8893 13640 8922
rect 13590 8873 13607 8893
rect 13627 8873 13640 8893
rect 13590 8845 13640 8873
rect 11980 8815 11998 8841
rect 12024 8815 12030 8841
rect 11980 8790 12030 8815
rect 2930 8727 2980 8740
rect 3138 8727 3188 8740
rect 3346 8727 3396 8740
rect 3559 8727 3609 8740
rect 8924 8756 8974 8772
rect 9132 8756 9182 8772
rect 9340 8756 9390 8772
rect 9553 8756 9603 8772
rect 3868 8715 3918 8731
rect 4076 8715 4126 8731
rect 4284 8715 4334 8731
rect 4497 8715 4547 8731
rect 381 8652 431 8665
rect 594 8652 644 8665
rect 802 8652 852 8665
rect 1010 8652 1060 8665
rect 3868 8648 3918 8673
rect 3868 8622 3874 8648
rect 3900 8622 3918 8648
rect 3868 8596 3918 8622
rect 4076 8644 4126 8673
rect 4076 8620 4090 8644
rect 4114 8620 4126 8644
rect 4076 8596 4126 8620
rect 4284 8649 4334 8673
rect 4284 8625 4299 8649
rect 4323 8625 4334 8649
rect 4284 8596 4334 8625
rect 4497 8644 4547 8673
rect 5437 8693 5487 8706
rect 5650 8693 5700 8706
rect 5858 8693 5908 8706
rect 6066 8693 6116 8706
rect 4497 8624 4514 8644
rect 4534 8624 4547 8644
rect 4497 8596 4547 8624
rect 381 8524 431 8552
rect 381 8504 394 8524
rect 414 8504 431 8524
rect 381 8475 431 8504
rect 594 8523 644 8552
rect 594 8499 605 8523
rect 629 8499 644 8523
rect 594 8475 644 8499
rect 802 8528 852 8552
rect 802 8504 814 8528
rect 838 8504 852 8528
rect 802 8475 852 8504
rect 1010 8526 1060 8552
rect 1010 8500 1028 8526
rect 1054 8500 1060 8526
rect 1010 8475 1060 8500
rect 8924 8689 8974 8714
rect 8924 8663 8930 8689
rect 8956 8663 8974 8689
rect 8924 8637 8974 8663
rect 9132 8685 9182 8714
rect 9132 8661 9146 8685
rect 9170 8661 9182 8685
rect 9132 8637 9182 8661
rect 9340 8690 9390 8714
rect 9340 8666 9355 8690
rect 9379 8666 9390 8690
rect 9340 8637 9390 8666
rect 9553 8685 9603 8714
rect 11351 8732 11401 8748
rect 11564 8732 11614 8748
rect 11772 8732 11822 8748
rect 11980 8732 12030 8748
rect 18017 9005 18067 9021
rect 18225 9005 18275 9021
rect 18433 9005 18483 9021
rect 18646 9005 18696 9021
rect 18017 8938 18067 8963
rect 18017 8912 18023 8938
rect 18049 8912 18067 8938
rect 16407 8880 16457 8908
rect 16407 8860 16420 8880
rect 16440 8860 16457 8880
rect 16407 8831 16457 8860
rect 16620 8879 16670 8908
rect 16620 8855 16631 8879
rect 16655 8855 16670 8879
rect 16620 8831 16670 8855
rect 16828 8884 16878 8908
rect 16828 8860 16840 8884
rect 16864 8860 16878 8884
rect 16828 8831 16878 8860
rect 17036 8882 17086 8908
rect 18017 8886 18067 8912
rect 18225 8934 18275 8963
rect 18225 8910 18239 8934
rect 18263 8910 18275 8934
rect 18225 8886 18275 8910
rect 18433 8939 18483 8963
rect 18433 8915 18448 8939
rect 18472 8915 18483 8939
rect 18433 8886 18483 8915
rect 18646 8934 18696 8963
rect 18646 8914 18663 8934
rect 18683 8914 18696 8934
rect 18646 8886 18696 8914
rect 17036 8856 17054 8882
rect 17080 8856 17086 8882
rect 17036 8831 17086 8856
rect 16407 8773 16457 8789
rect 16620 8773 16670 8789
rect 16828 8773 16878 8789
rect 17036 8773 17086 8789
rect 18017 8773 18067 8786
rect 18225 8773 18275 8786
rect 18433 8773 18483 8786
rect 18646 8773 18696 8786
rect 12961 8732 13011 8745
rect 13169 8732 13219 8745
rect 13377 8732 13427 8745
rect 13590 8732 13640 8745
rect 18955 8761 19005 8777
rect 19163 8761 19213 8777
rect 19371 8761 19421 8777
rect 19584 8761 19634 8777
rect 9553 8665 9570 8685
rect 9590 8665 9603 8685
rect 13899 8720 13949 8736
rect 14107 8720 14157 8736
rect 14315 8720 14365 8736
rect 14528 8720 14578 8736
rect 9553 8637 9603 8665
rect 5437 8565 5487 8593
rect 5437 8545 5450 8565
rect 5470 8545 5487 8565
rect 5437 8516 5487 8545
rect 5650 8564 5700 8593
rect 5650 8540 5661 8564
rect 5685 8540 5700 8564
rect 5650 8516 5700 8540
rect 5858 8569 5908 8593
rect 5858 8545 5870 8569
rect 5894 8545 5908 8569
rect 5858 8516 5908 8545
rect 6066 8567 6116 8593
rect 6066 8541 6084 8567
rect 6110 8541 6116 8567
rect 6066 8516 6116 8541
rect 10412 8657 10462 8670
rect 10625 8657 10675 8670
rect 10833 8657 10883 8670
rect 11041 8657 11091 8670
rect 13899 8653 13949 8678
rect 13899 8627 13905 8653
rect 13931 8627 13949 8653
rect 13899 8601 13949 8627
rect 14107 8649 14157 8678
rect 14107 8625 14121 8649
rect 14145 8625 14157 8649
rect 14107 8601 14157 8625
rect 14315 8654 14365 8678
rect 14315 8630 14330 8654
rect 14354 8630 14365 8654
rect 14315 8601 14365 8630
rect 14528 8649 14578 8678
rect 15468 8698 15518 8711
rect 15681 8698 15731 8711
rect 15889 8698 15939 8711
rect 16097 8698 16147 8711
rect 14528 8629 14545 8649
rect 14565 8629 14578 8649
rect 14528 8601 14578 8629
rect 8924 8524 8974 8537
rect 9132 8524 9182 8537
rect 9340 8524 9390 8537
rect 9553 8524 9603 8537
rect 10412 8529 10462 8557
rect 3868 8483 3918 8496
rect 4076 8483 4126 8496
rect 4284 8483 4334 8496
rect 4497 8483 4547 8496
rect 2790 8448 2840 8464
rect 2998 8448 3048 8464
rect 3206 8448 3256 8464
rect 3419 8448 3469 8464
rect 381 8417 431 8433
rect 594 8417 644 8433
rect 802 8417 852 8433
rect 1010 8417 1060 8433
rect 7846 8489 7896 8505
rect 8054 8489 8104 8505
rect 8262 8489 8312 8505
rect 8475 8489 8525 8505
rect 5437 8458 5487 8474
rect 5650 8458 5700 8474
rect 5858 8458 5908 8474
rect 6066 8458 6116 8474
rect 10412 8509 10425 8529
rect 10445 8509 10462 8529
rect 10412 8480 10462 8509
rect 10625 8528 10675 8557
rect 10625 8504 10636 8528
rect 10660 8504 10675 8528
rect 10625 8480 10675 8504
rect 10833 8533 10883 8557
rect 10833 8509 10845 8533
rect 10869 8509 10883 8533
rect 10833 8480 10883 8509
rect 11041 8531 11091 8557
rect 11041 8505 11059 8531
rect 11085 8505 11091 8531
rect 11041 8480 11091 8505
rect 18955 8694 19005 8719
rect 18955 8668 18961 8694
rect 18987 8668 19005 8694
rect 18955 8642 19005 8668
rect 19163 8690 19213 8719
rect 19163 8666 19177 8690
rect 19201 8666 19213 8690
rect 19163 8642 19213 8666
rect 19371 8695 19421 8719
rect 19371 8671 19386 8695
rect 19410 8671 19421 8695
rect 19371 8642 19421 8671
rect 19584 8690 19634 8719
rect 19584 8670 19601 8690
rect 19621 8670 19634 8690
rect 19584 8642 19634 8670
rect 15468 8570 15518 8598
rect 15468 8550 15481 8570
rect 15501 8550 15518 8570
rect 15468 8521 15518 8550
rect 15681 8569 15731 8598
rect 15681 8545 15692 8569
rect 15716 8545 15731 8569
rect 15681 8521 15731 8545
rect 15889 8574 15939 8598
rect 15889 8550 15901 8574
rect 15925 8550 15939 8574
rect 15889 8521 15939 8550
rect 16097 8572 16147 8598
rect 16097 8546 16115 8572
rect 16141 8546 16147 8572
rect 16097 8521 16147 8546
rect 18955 8529 19005 8542
rect 19163 8529 19213 8542
rect 19371 8529 19421 8542
rect 19584 8529 19634 8542
rect 13899 8488 13949 8501
rect 14107 8488 14157 8501
rect 14315 8488 14365 8501
rect 14528 8488 14578 8501
rect 1461 8370 1511 8383
rect 1674 8370 1724 8383
rect 1882 8370 1932 8383
rect 2090 8370 2140 8383
rect 2790 8381 2840 8406
rect 2790 8355 2796 8381
rect 2822 8355 2840 8381
rect 2790 8329 2840 8355
rect 2998 8377 3048 8406
rect 2998 8353 3012 8377
rect 3036 8353 3048 8377
rect 2998 8329 3048 8353
rect 3206 8382 3256 8406
rect 3206 8358 3221 8382
rect 3245 8358 3256 8382
rect 3206 8329 3256 8358
rect 3419 8377 3469 8406
rect 6517 8411 6567 8424
rect 6730 8411 6780 8424
rect 6938 8411 6988 8424
rect 7146 8411 7196 8424
rect 7846 8422 7896 8447
rect 3419 8357 3436 8377
rect 3456 8357 3469 8377
rect 3419 8329 3469 8357
rect 1461 8242 1511 8270
rect 1461 8222 1474 8242
rect 1494 8222 1511 8242
rect 1461 8193 1511 8222
rect 1674 8241 1724 8270
rect 1674 8217 1685 8241
rect 1709 8217 1724 8241
rect 1674 8193 1724 8217
rect 1882 8246 1932 8270
rect 1882 8222 1894 8246
rect 1918 8222 1932 8246
rect 1882 8193 1932 8222
rect 2090 8244 2140 8270
rect 2090 8218 2108 8244
rect 2134 8218 2140 8244
rect 7846 8396 7852 8422
rect 7878 8396 7896 8422
rect 7846 8370 7896 8396
rect 8054 8418 8104 8447
rect 8054 8394 8068 8418
rect 8092 8394 8104 8418
rect 8054 8370 8104 8394
rect 8262 8423 8312 8447
rect 8262 8399 8277 8423
rect 8301 8399 8312 8423
rect 8262 8370 8312 8399
rect 8475 8418 8525 8447
rect 12821 8453 12871 8469
rect 13029 8453 13079 8469
rect 13237 8453 13287 8469
rect 13450 8453 13500 8469
rect 10412 8422 10462 8438
rect 10625 8422 10675 8438
rect 10833 8422 10883 8438
rect 11041 8422 11091 8438
rect 8475 8398 8492 8418
rect 8512 8398 8525 8418
rect 17877 8494 17927 8510
rect 18085 8494 18135 8510
rect 18293 8494 18343 8510
rect 18506 8494 18556 8510
rect 15468 8463 15518 8479
rect 15681 8463 15731 8479
rect 15889 8463 15939 8479
rect 16097 8463 16147 8479
rect 8475 8370 8525 8398
rect 6517 8283 6567 8311
rect 6517 8263 6530 8283
rect 6550 8263 6567 8283
rect 2090 8193 2140 8218
rect 2790 8216 2840 8229
rect 2998 8216 3048 8229
rect 3206 8216 3256 8229
rect 3419 8216 3469 8229
rect 6517 8234 6567 8263
rect 6730 8282 6780 8311
rect 6730 8258 6741 8282
rect 6765 8258 6780 8282
rect 6730 8234 6780 8258
rect 6938 8287 6988 8311
rect 6938 8263 6950 8287
rect 6974 8263 6988 8287
rect 6938 8234 6988 8263
rect 7146 8285 7196 8311
rect 7146 8259 7164 8285
rect 7190 8259 7196 8285
rect 11492 8375 11542 8388
rect 11705 8375 11755 8388
rect 11913 8375 11963 8388
rect 12121 8375 12171 8388
rect 12821 8386 12871 8411
rect 7146 8234 7196 8259
rect 7846 8257 7896 8270
rect 8054 8257 8104 8270
rect 8262 8257 8312 8270
rect 8475 8257 8525 8270
rect 12821 8360 12827 8386
rect 12853 8360 12871 8386
rect 12821 8334 12871 8360
rect 13029 8382 13079 8411
rect 13029 8358 13043 8382
rect 13067 8358 13079 8382
rect 13029 8334 13079 8358
rect 13237 8387 13287 8411
rect 13237 8363 13252 8387
rect 13276 8363 13287 8387
rect 13237 8334 13287 8363
rect 13450 8382 13500 8411
rect 16548 8416 16598 8429
rect 16761 8416 16811 8429
rect 16969 8416 17019 8429
rect 17177 8416 17227 8429
rect 17877 8427 17927 8452
rect 13450 8362 13467 8382
rect 13487 8362 13500 8382
rect 13450 8334 13500 8362
rect 11492 8247 11542 8275
rect 3870 8166 3920 8182
rect 4078 8166 4128 8182
rect 4286 8166 4336 8182
rect 4499 8166 4549 8182
rect 1461 8135 1511 8151
rect 1674 8135 1724 8151
rect 1882 8135 1932 8151
rect 2090 8135 2140 8151
rect 11492 8227 11505 8247
rect 11525 8227 11542 8247
rect 8926 8207 8976 8223
rect 9134 8207 9184 8223
rect 9342 8207 9392 8223
rect 9555 8207 9605 8223
rect 6517 8176 6567 8192
rect 6730 8176 6780 8192
rect 6938 8176 6988 8192
rect 7146 8176 7196 8192
rect 11492 8198 11542 8227
rect 11705 8246 11755 8275
rect 11705 8222 11716 8246
rect 11740 8222 11755 8246
rect 11705 8198 11755 8222
rect 11913 8251 11963 8275
rect 11913 8227 11925 8251
rect 11949 8227 11963 8251
rect 11913 8198 11963 8227
rect 12121 8249 12171 8275
rect 12121 8223 12139 8249
rect 12165 8223 12171 8249
rect 17877 8401 17883 8427
rect 17909 8401 17927 8427
rect 17877 8375 17927 8401
rect 18085 8423 18135 8452
rect 18085 8399 18099 8423
rect 18123 8399 18135 8423
rect 18085 8375 18135 8399
rect 18293 8428 18343 8452
rect 18293 8404 18308 8428
rect 18332 8404 18343 8428
rect 18293 8375 18343 8404
rect 18506 8423 18556 8452
rect 18506 8403 18523 8423
rect 18543 8403 18556 8423
rect 18506 8375 18556 8403
rect 16548 8288 16598 8316
rect 16548 8268 16561 8288
rect 16581 8268 16598 8288
rect 12121 8198 12171 8223
rect 12821 8221 12871 8234
rect 13029 8221 13079 8234
rect 13237 8221 13287 8234
rect 13450 8221 13500 8234
rect 16548 8239 16598 8268
rect 16761 8287 16811 8316
rect 16761 8263 16772 8287
rect 16796 8263 16811 8287
rect 16761 8239 16811 8263
rect 16969 8292 17019 8316
rect 16969 8268 16981 8292
rect 17005 8268 17019 8292
rect 16969 8239 17019 8268
rect 17177 8290 17227 8316
rect 17177 8264 17195 8290
rect 17221 8264 17227 8290
rect 17177 8239 17227 8264
rect 17877 8262 17927 8275
rect 18085 8262 18135 8275
rect 18293 8262 18343 8275
rect 18506 8262 18556 8275
rect 5439 8144 5489 8157
rect 5652 8144 5702 8157
rect 5860 8144 5910 8157
rect 6068 8144 6118 8157
rect 383 8103 433 8116
rect 596 8103 646 8116
rect 804 8103 854 8116
rect 1012 8103 1062 8116
rect 3870 8099 3920 8124
rect 3870 8073 3876 8099
rect 3902 8073 3920 8099
rect 3870 8047 3920 8073
rect 4078 8095 4128 8124
rect 4078 8071 4092 8095
rect 4116 8071 4128 8095
rect 4078 8047 4128 8071
rect 4286 8100 4336 8124
rect 4286 8076 4301 8100
rect 4325 8076 4336 8100
rect 4286 8047 4336 8076
rect 4499 8095 4549 8124
rect 4499 8075 4516 8095
rect 4536 8075 4549 8095
rect 4499 8047 4549 8075
rect 383 7975 433 8003
rect 383 7955 396 7975
rect 416 7955 433 7975
rect 383 7926 433 7955
rect 596 7974 646 8003
rect 596 7950 607 7974
rect 631 7950 646 7974
rect 596 7926 646 7950
rect 804 7979 854 8003
rect 804 7955 816 7979
rect 840 7955 854 7979
rect 804 7926 854 7955
rect 1012 7977 1062 8003
rect 1012 7951 1030 7977
rect 1056 7951 1062 7977
rect 1012 7926 1062 7951
rect 8926 8140 8976 8165
rect 8926 8114 8932 8140
rect 8958 8114 8976 8140
rect 8926 8088 8976 8114
rect 9134 8136 9184 8165
rect 9134 8112 9148 8136
rect 9172 8112 9184 8136
rect 9134 8088 9184 8112
rect 9342 8141 9392 8165
rect 9342 8117 9357 8141
rect 9381 8117 9392 8141
rect 9342 8088 9392 8117
rect 9555 8136 9605 8165
rect 9555 8116 9572 8136
rect 9592 8116 9605 8136
rect 13901 8171 13951 8187
rect 14109 8171 14159 8187
rect 14317 8171 14367 8187
rect 14530 8171 14580 8187
rect 11492 8140 11542 8156
rect 11705 8140 11755 8156
rect 11913 8140 11963 8156
rect 12121 8140 12171 8156
rect 18957 8212 19007 8228
rect 19165 8212 19215 8228
rect 19373 8212 19423 8228
rect 19586 8212 19636 8228
rect 16548 8181 16598 8197
rect 16761 8181 16811 8197
rect 16969 8181 17019 8197
rect 17177 8181 17227 8197
rect 15470 8149 15520 8162
rect 15683 8149 15733 8162
rect 15891 8149 15941 8162
rect 16099 8149 16149 8162
rect 9555 8088 9605 8116
rect 10414 8108 10464 8121
rect 10627 8108 10677 8121
rect 10835 8108 10885 8121
rect 11043 8108 11093 8121
rect 5439 8016 5489 8044
rect 5439 7996 5452 8016
rect 5472 7996 5489 8016
rect 3870 7934 3920 7947
rect 4078 7934 4128 7947
rect 4286 7934 4336 7947
rect 4499 7934 4549 7947
rect 5439 7967 5489 7996
rect 5652 8015 5702 8044
rect 5652 7991 5663 8015
rect 5687 7991 5702 8015
rect 5652 7967 5702 7991
rect 5860 8020 5910 8044
rect 5860 7996 5872 8020
rect 5896 7996 5910 8020
rect 5860 7967 5910 7996
rect 6068 8018 6118 8044
rect 6068 7992 6086 8018
rect 6112 7992 6118 8018
rect 6068 7967 6118 7992
rect 8926 7975 8976 7988
rect 9134 7975 9184 7988
rect 9342 7975 9392 7988
rect 9555 7975 9605 7988
rect 13901 8104 13951 8129
rect 13901 8078 13907 8104
rect 13933 8078 13951 8104
rect 13901 8052 13951 8078
rect 14109 8100 14159 8129
rect 14109 8076 14123 8100
rect 14147 8076 14159 8100
rect 14109 8052 14159 8076
rect 14317 8105 14367 8129
rect 14317 8081 14332 8105
rect 14356 8081 14367 8105
rect 14317 8052 14367 8081
rect 14530 8100 14580 8129
rect 14530 8080 14547 8100
rect 14567 8080 14580 8100
rect 14530 8052 14580 8080
rect 10414 7980 10464 8008
rect 5439 7909 5489 7925
rect 5652 7909 5702 7925
rect 5860 7909 5910 7925
rect 6068 7909 6118 7925
rect 10414 7960 10427 7980
rect 10447 7960 10464 7980
rect 383 7868 433 7884
rect 596 7868 646 7884
rect 804 7868 854 7884
rect 1012 7868 1062 7884
rect 6377 7900 6427 7913
rect 6590 7900 6640 7913
rect 6798 7900 6848 7913
rect 7006 7900 7056 7913
rect 1321 7859 1371 7872
rect 1534 7859 1584 7872
rect 1742 7859 1792 7872
rect 1950 7859 2000 7872
rect 2931 7856 2981 7872
rect 3139 7856 3189 7872
rect 3347 7856 3397 7872
rect 3560 7856 3610 7872
rect 2931 7789 2981 7814
rect 2931 7763 2937 7789
rect 2963 7763 2981 7789
rect 1321 7731 1371 7759
rect 1321 7711 1334 7731
rect 1354 7711 1371 7731
rect 1321 7682 1371 7711
rect 1534 7730 1584 7759
rect 1534 7706 1545 7730
rect 1569 7706 1584 7730
rect 1534 7682 1584 7706
rect 1742 7735 1792 7759
rect 1742 7711 1754 7735
rect 1778 7711 1792 7735
rect 1742 7682 1792 7711
rect 1950 7733 2000 7759
rect 2931 7737 2981 7763
rect 3139 7785 3189 7814
rect 3139 7761 3153 7785
rect 3177 7761 3189 7785
rect 3139 7737 3189 7761
rect 3347 7790 3397 7814
rect 3347 7766 3362 7790
rect 3386 7766 3397 7790
rect 3347 7737 3397 7766
rect 3560 7785 3610 7814
rect 3560 7765 3577 7785
rect 3597 7765 3610 7785
rect 3560 7737 3610 7765
rect 1950 7707 1968 7733
rect 1994 7707 2000 7733
rect 1950 7682 2000 7707
rect 1321 7624 1371 7640
rect 1534 7624 1584 7640
rect 1742 7624 1792 7640
rect 1950 7624 2000 7640
rect 7987 7897 8037 7913
rect 8195 7897 8245 7913
rect 8403 7897 8453 7913
rect 8616 7897 8666 7913
rect 10414 7931 10464 7960
rect 10627 7979 10677 8008
rect 10627 7955 10638 7979
rect 10662 7955 10677 7979
rect 10627 7931 10677 7955
rect 10835 7984 10885 8008
rect 10835 7960 10847 7984
rect 10871 7960 10885 7984
rect 10835 7931 10885 7960
rect 11043 7982 11093 8008
rect 11043 7956 11061 7982
rect 11087 7956 11093 7982
rect 11043 7931 11093 7956
rect 18957 8145 19007 8170
rect 18957 8119 18963 8145
rect 18989 8119 19007 8145
rect 18957 8093 19007 8119
rect 19165 8141 19215 8170
rect 19165 8117 19179 8141
rect 19203 8117 19215 8141
rect 19165 8093 19215 8117
rect 19373 8146 19423 8170
rect 19373 8122 19388 8146
rect 19412 8122 19423 8146
rect 19373 8093 19423 8122
rect 19586 8141 19636 8170
rect 19586 8121 19603 8141
rect 19623 8121 19636 8141
rect 19586 8093 19636 8121
rect 15470 8021 15520 8049
rect 15470 8001 15483 8021
rect 15503 8001 15520 8021
rect 13901 7939 13951 7952
rect 14109 7939 14159 7952
rect 14317 7939 14367 7952
rect 14530 7939 14580 7952
rect 15470 7972 15520 8001
rect 15683 8020 15733 8049
rect 15683 7996 15694 8020
rect 15718 7996 15733 8020
rect 15683 7972 15733 7996
rect 15891 8025 15941 8049
rect 15891 8001 15903 8025
rect 15927 8001 15941 8025
rect 15891 7972 15941 8001
rect 16099 8023 16149 8049
rect 16099 7997 16117 8023
rect 16143 7997 16149 8023
rect 16099 7972 16149 7997
rect 18957 7980 19007 7993
rect 19165 7980 19215 7993
rect 19373 7980 19423 7993
rect 19586 7980 19636 7993
rect 15470 7914 15520 7930
rect 15683 7914 15733 7930
rect 15891 7914 15941 7930
rect 16099 7914 16149 7930
rect 10414 7873 10464 7889
rect 10627 7873 10677 7889
rect 10835 7873 10885 7889
rect 11043 7873 11093 7889
rect 16408 7905 16458 7918
rect 16621 7905 16671 7918
rect 16829 7905 16879 7918
rect 17037 7905 17087 7918
rect 7987 7830 8037 7855
rect 7987 7804 7993 7830
rect 8019 7804 8037 7830
rect 6377 7772 6427 7800
rect 6377 7752 6390 7772
rect 6410 7752 6427 7772
rect 6377 7723 6427 7752
rect 6590 7771 6640 7800
rect 6590 7747 6601 7771
rect 6625 7747 6640 7771
rect 6590 7723 6640 7747
rect 6798 7776 6848 7800
rect 6798 7752 6810 7776
rect 6834 7752 6848 7776
rect 6798 7723 6848 7752
rect 7006 7774 7056 7800
rect 7987 7778 8037 7804
rect 8195 7826 8245 7855
rect 8195 7802 8209 7826
rect 8233 7802 8245 7826
rect 8195 7778 8245 7802
rect 8403 7831 8453 7855
rect 8403 7807 8418 7831
rect 8442 7807 8453 7831
rect 8403 7778 8453 7807
rect 8616 7826 8666 7855
rect 11352 7864 11402 7877
rect 11565 7864 11615 7877
rect 11773 7864 11823 7877
rect 11981 7864 12031 7877
rect 8616 7806 8633 7826
rect 8653 7806 8666 7826
rect 8616 7778 8666 7806
rect 7006 7748 7024 7774
rect 7050 7748 7056 7774
rect 7006 7723 7056 7748
rect 6377 7665 6427 7681
rect 6590 7665 6640 7681
rect 6798 7665 6848 7681
rect 7006 7665 7056 7681
rect 12962 7861 13012 7877
rect 13170 7861 13220 7877
rect 13378 7861 13428 7877
rect 13591 7861 13641 7877
rect 12962 7794 13012 7819
rect 12962 7768 12968 7794
rect 12994 7768 13012 7794
rect 11352 7736 11402 7764
rect 11352 7716 11365 7736
rect 11385 7716 11402 7736
rect 7987 7665 8037 7678
rect 8195 7665 8245 7678
rect 8403 7665 8453 7678
rect 8616 7665 8666 7678
rect 11352 7687 11402 7716
rect 11565 7735 11615 7764
rect 11565 7711 11576 7735
rect 11600 7711 11615 7735
rect 11565 7687 11615 7711
rect 11773 7740 11823 7764
rect 11773 7716 11785 7740
rect 11809 7716 11823 7740
rect 11773 7687 11823 7716
rect 11981 7738 12031 7764
rect 12962 7742 13012 7768
rect 13170 7790 13220 7819
rect 13170 7766 13184 7790
rect 13208 7766 13220 7790
rect 13170 7742 13220 7766
rect 13378 7795 13428 7819
rect 13378 7771 13393 7795
rect 13417 7771 13428 7795
rect 13378 7742 13428 7771
rect 13591 7790 13641 7819
rect 13591 7770 13608 7790
rect 13628 7770 13641 7790
rect 13591 7742 13641 7770
rect 11981 7712 11999 7738
rect 12025 7712 12031 7738
rect 11981 7687 12031 7712
rect 2931 7624 2981 7637
rect 3139 7624 3189 7637
rect 3347 7624 3397 7637
rect 3560 7624 3610 7637
rect 8925 7653 8975 7669
rect 9133 7653 9183 7669
rect 9341 7653 9391 7669
rect 9554 7653 9604 7669
rect 3869 7612 3919 7628
rect 4077 7612 4127 7628
rect 4285 7612 4335 7628
rect 4498 7612 4548 7628
rect 382 7549 432 7562
rect 595 7549 645 7562
rect 803 7549 853 7562
rect 1011 7549 1061 7562
rect 3869 7545 3919 7570
rect 3869 7519 3875 7545
rect 3901 7519 3919 7545
rect 3869 7493 3919 7519
rect 4077 7541 4127 7570
rect 4077 7517 4091 7541
rect 4115 7517 4127 7541
rect 4077 7493 4127 7517
rect 4285 7546 4335 7570
rect 4285 7522 4300 7546
rect 4324 7522 4335 7546
rect 4285 7493 4335 7522
rect 4498 7541 4548 7570
rect 5438 7590 5488 7603
rect 5651 7590 5701 7603
rect 5859 7590 5909 7603
rect 6067 7590 6117 7603
rect 4498 7521 4515 7541
rect 4535 7521 4548 7541
rect 4498 7493 4548 7521
rect 382 7421 432 7449
rect 382 7401 395 7421
rect 415 7401 432 7421
rect 382 7372 432 7401
rect 595 7420 645 7449
rect 595 7396 606 7420
rect 630 7396 645 7420
rect 595 7372 645 7396
rect 803 7425 853 7449
rect 803 7401 815 7425
rect 839 7401 853 7425
rect 803 7372 853 7401
rect 1011 7423 1061 7449
rect 1011 7397 1029 7423
rect 1055 7397 1061 7423
rect 1011 7372 1061 7397
rect 8925 7586 8975 7611
rect 8925 7560 8931 7586
rect 8957 7560 8975 7586
rect 8925 7534 8975 7560
rect 9133 7582 9183 7611
rect 9133 7558 9147 7582
rect 9171 7558 9183 7582
rect 9133 7534 9183 7558
rect 9341 7587 9391 7611
rect 9341 7563 9356 7587
rect 9380 7563 9391 7587
rect 9341 7534 9391 7563
rect 9554 7582 9604 7611
rect 11352 7629 11402 7645
rect 11565 7629 11615 7645
rect 11773 7629 11823 7645
rect 11981 7629 12031 7645
rect 18018 7902 18068 7918
rect 18226 7902 18276 7918
rect 18434 7902 18484 7918
rect 18647 7902 18697 7918
rect 18018 7835 18068 7860
rect 18018 7809 18024 7835
rect 18050 7809 18068 7835
rect 16408 7777 16458 7805
rect 16408 7757 16421 7777
rect 16441 7757 16458 7777
rect 16408 7728 16458 7757
rect 16621 7776 16671 7805
rect 16621 7752 16632 7776
rect 16656 7752 16671 7776
rect 16621 7728 16671 7752
rect 16829 7781 16879 7805
rect 16829 7757 16841 7781
rect 16865 7757 16879 7781
rect 16829 7728 16879 7757
rect 17037 7779 17087 7805
rect 18018 7783 18068 7809
rect 18226 7831 18276 7860
rect 18226 7807 18240 7831
rect 18264 7807 18276 7831
rect 18226 7783 18276 7807
rect 18434 7836 18484 7860
rect 18434 7812 18449 7836
rect 18473 7812 18484 7836
rect 18434 7783 18484 7812
rect 18647 7831 18697 7860
rect 18647 7811 18664 7831
rect 18684 7811 18697 7831
rect 18647 7783 18697 7811
rect 17037 7753 17055 7779
rect 17081 7753 17087 7779
rect 17037 7728 17087 7753
rect 16408 7670 16458 7686
rect 16621 7670 16671 7686
rect 16829 7670 16879 7686
rect 17037 7670 17087 7686
rect 18018 7670 18068 7683
rect 18226 7670 18276 7683
rect 18434 7670 18484 7683
rect 18647 7670 18697 7683
rect 12962 7629 13012 7642
rect 13170 7629 13220 7642
rect 13378 7629 13428 7642
rect 13591 7629 13641 7642
rect 18956 7658 19006 7674
rect 19164 7658 19214 7674
rect 19372 7658 19422 7674
rect 19585 7658 19635 7674
rect 9554 7562 9571 7582
rect 9591 7562 9604 7582
rect 13900 7617 13950 7633
rect 14108 7617 14158 7633
rect 14316 7617 14366 7633
rect 14529 7617 14579 7633
rect 9554 7534 9604 7562
rect 5438 7462 5488 7490
rect 5438 7442 5451 7462
rect 5471 7442 5488 7462
rect 5438 7413 5488 7442
rect 5651 7461 5701 7490
rect 5651 7437 5662 7461
rect 5686 7437 5701 7461
rect 5651 7413 5701 7437
rect 5859 7466 5909 7490
rect 5859 7442 5871 7466
rect 5895 7442 5909 7466
rect 5859 7413 5909 7442
rect 6067 7464 6117 7490
rect 6067 7438 6085 7464
rect 6111 7438 6117 7464
rect 6067 7413 6117 7438
rect 10413 7554 10463 7567
rect 10626 7554 10676 7567
rect 10834 7554 10884 7567
rect 11042 7554 11092 7567
rect 13900 7550 13950 7575
rect 13900 7524 13906 7550
rect 13932 7524 13950 7550
rect 13900 7498 13950 7524
rect 14108 7546 14158 7575
rect 14108 7522 14122 7546
rect 14146 7522 14158 7546
rect 14108 7498 14158 7522
rect 14316 7551 14366 7575
rect 14316 7527 14331 7551
rect 14355 7527 14366 7551
rect 14316 7498 14366 7527
rect 14529 7546 14579 7575
rect 15469 7595 15519 7608
rect 15682 7595 15732 7608
rect 15890 7595 15940 7608
rect 16098 7595 16148 7608
rect 14529 7526 14546 7546
rect 14566 7526 14579 7546
rect 14529 7498 14579 7526
rect 8925 7421 8975 7434
rect 9133 7421 9183 7434
rect 9341 7421 9391 7434
rect 9554 7421 9604 7434
rect 10413 7426 10463 7454
rect 3869 7380 3919 7393
rect 4077 7380 4127 7393
rect 4285 7380 4335 7393
rect 4498 7380 4548 7393
rect 382 7314 432 7330
rect 595 7314 645 7330
rect 803 7314 853 7330
rect 1011 7314 1061 7330
rect 2821 7332 2871 7348
rect 3029 7332 3079 7348
rect 3237 7332 3287 7348
rect 3450 7332 3500 7348
rect 1431 7280 1481 7293
rect 1644 7280 1694 7293
rect 1852 7280 1902 7293
rect 2060 7280 2110 7293
rect 5438 7355 5488 7371
rect 5651 7355 5701 7371
rect 5859 7355 5909 7371
rect 6067 7355 6117 7371
rect 7877 7373 7927 7389
rect 8085 7373 8135 7389
rect 8293 7373 8343 7389
rect 8506 7373 8556 7389
rect 6487 7321 6537 7334
rect 6700 7321 6750 7334
rect 6908 7321 6958 7334
rect 7116 7321 7166 7334
rect 10413 7406 10426 7426
rect 10446 7406 10463 7426
rect 10413 7377 10463 7406
rect 10626 7425 10676 7454
rect 10626 7401 10637 7425
rect 10661 7401 10676 7425
rect 10626 7377 10676 7401
rect 10834 7430 10884 7454
rect 10834 7406 10846 7430
rect 10870 7406 10884 7430
rect 10834 7377 10884 7406
rect 11042 7428 11092 7454
rect 11042 7402 11060 7428
rect 11086 7402 11092 7428
rect 11042 7377 11092 7402
rect 18956 7591 19006 7616
rect 18956 7565 18962 7591
rect 18988 7565 19006 7591
rect 18956 7539 19006 7565
rect 19164 7587 19214 7616
rect 19164 7563 19178 7587
rect 19202 7563 19214 7587
rect 19164 7539 19214 7563
rect 19372 7592 19422 7616
rect 19372 7568 19387 7592
rect 19411 7568 19422 7592
rect 19372 7539 19422 7568
rect 19585 7587 19635 7616
rect 19585 7567 19602 7587
rect 19622 7567 19635 7587
rect 19585 7539 19635 7567
rect 15469 7467 15519 7495
rect 15469 7447 15482 7467
rect 15502 7447 15519 7467
rect 15469 7418 15519 7447
rect 15682 7466 15732 7495
rect 15682 7442 15693 7466
rect 15717 7442 15732 7466
rect 15682 7418 15732 7442
rect 15890 7471 15940 7495
rect 15890 7447 15902 7471
rect 15926 7447 15940 7471
rect 15890 7418 15940 7447
rect 16098 7469 16148 7495
rect 16098 7443 16116 7469
rect 16142 7443 16148 7469
rect 16098 7418 16148 7443
rect 18956 7426 19006 7439
rect 19164 7426 19214 7439
rect 19372 7426 19422 7439
rect 19585 7426 19635 7439
rect 13900 7385 13950 7398
rect 14108 7385 14158 7398
rect 14316 7385 14366 7398
rect 14529 7385 14579 7398
rect 2821 7265 2871 7290
rect 2821 7239 2827 7265
rect 2853 7239 2871 7265
rect 2821 7213 2871 7239
rect 3029 7261 3079 7290
rect 3029 7237 3043 7261
rect 3067 7237 3079 7261
rect 3029 7213 3079 7237
rect 3237 7266 3287 7290
rect 3237 7242 3252 7266
rect 3276 7242 3287 7266
rect 3237 7213 3287 7242
rect 3450 7261 3500 7290
rect 3450 7241 3467 7261
rect 3487 7241 3500 7261
rect 3450 7213 3500 7241
rect 7877 7306 7927 7331
rect 7877 7280 7883 7306
rect 7909 7280 7927 7306
rect 7877 7254 7927 7280
rect 8085 7302 8135 7331
rect 8085 7278 8099 7302
rect 8123 7278 8135 7302
rect 8085 7254 8135 7278
rect 8293 7307 8343 7331
rect 8293 7283 8308 7307
rect 8332 7283 8343 7307
rect 8293 7254 8343 7283
rect 8506 7302 8556 7331
rect 10413 7319 10463 7335
rect 10626 7319 10676 7335
rect 10834 7319 10884 7335
rect 11042 7319 11092 7335
rect 12852 7337 12902 7353
rect 13060 7337 13110 7353
rect 13268 7337 13318 7353
rect 13481 7337 13531 7353
rect 8506 7282 8523 7302
rect 8543 7282 8556 7302
rect 8506 7254 8556 7282
rect 11462 7285 11512 7298
rect 11675 7285 11725 7298
rect 11883 7285 11933 7298
rect 12091 7285 12141 7298
rect 15469 7360 15519 7376
rect 15682 7360 15732 7376
rect 15890 7360 15940 7376
rect 16098 7360 16148 7376
rect 17908 7378 17958 7394
rect 18116 7378 18166 7394
rect 18324 7378 18374 7394
rect 18537 7378 18587 7394
rect 16518 7326 16568 7339
rect 16731 7326 16781 7339
rect 16939 7326 16989 7339
rect 17147 7326 17197 7339
rect 1431 7152 1481 7180
rect 1431 7132 1444 7152
rect 1464 7132 1481 7152
rect 1431 7103 1481 7132
rect 1644 7151 1694 7180
rect 1644 7127 1655 7151
rect 1679 7127 1694 7151
rect 1644 7103 1694 7127
rect 1852 7156 1902 7180
rect 1852 7132 1864 7156
rect 1888 7132 1902 7156
rect 1852 7103 1902 7132
rect 2060 7154 2110 7180
rect 2060 7128 2078 7154
rect 2104 7128 2110 7154
rect 2060 7103 2110 7128
rect 6487 7193 6537 7221
rect 6487 7173 6500 7193
rect 6520 7173 6537 7193
rect 6487 7144 6537 7173
rect 6700 7192 6750 7221
rect 6700 7168 6711 7192
rect 6735 7168 6750 7192
rect 6700 7144 6750 7168
rect 6908 7197 6958 7221
rect 6908 7173 6920 7197
rect 6944 7173 6958 7197
rect 6908 7144 6958 7173
rect 7116 7195 7166 7221
rect 7116 7169 7134 7195
rect 7160 7169 7166 7195
rect 7116 7144 7166 7169
rect 12852 7270 12902 7295
rect 12852 7244 12858 7270
rect 12884 7244 12902 7270
rect 12852 7218 12902 7244
rect 13060 7266 13110 7295
rect 13060 7242 13074 7266
rect 13098 7242 13110 7266
rect 13060 7218 13110 7242
rect 13268 7271 13318 7295
rect 13268 7247 13283 7271
rect 13307 7247 13318 7271
rect 13268 7218 13318 7247
rect 13481 7266 13531 7295
rect 13481 7246 13498 7266
rect 13518 7246 13531 7266
rect 13481 7218 13531 7246
rect 17908 7311 17958 7336
rect 17908 7285 17914 7311
rect 17940 7285 17958 7311
rect 17908 7259 17958 7285
rect 18116 7307 18166 7336
rect 18116 7283 18130 7307
rect 18154 7283 18166 7307
rect 18116 7259 18166 7283
rect 18324 7312 18374 7336
rect 18324 7288 18339 7312
rect 18363 7288 18374 7312
rect 18324 7259 18374 7288
rect 18537 7307 18587 7336
rect 18537 7287 18554 7307
rect 18574 7287 18587 7307
rect 18537 7259 18587 7287
rect 2821 7100 2871 7113
rect 3029 7100 3079 7113
rect 3237 7100 3287 7113
rect 3450 7100 3500 7113
rect 1431 7045 1481 7061
rect 1644 7045 1694 7061
rect 1852 7045 1902 7061
rect 2060 7045 2110 7061
rect 3870 7063 3920 7079
rect 4078 7063 4128 7079
rect 4286 7063 4336 7079
rect 4499 7063 4549 7079
rect 7877 7141 7927 7154
rect 8085 7141 8135 7154
rect 8293 7141 8343 7154
rect 8506 7141 8556 7154
rect 11462 7157 11512 7185
rect 11462 7137 11475 7157
rect 11495 7137 11512 7157
rect 6487 7086 6537 7102
rect 6700 7086 6750 7102
rect 6908 7086 6958 7102
rect 7116 7086 7166 7102
rect 8926 7104 8976 7120
rect 9134 7104 9184 7120
rect 9342 7104 9392 7120
rect 9555 7104 9605 7120
rect 11462 7108 11512 7137
rect 11675 7156 11725 7185
rect 11675 7132 11686 7156
rect 11710 7132 11725 7156
rect 11675 7108 11725 7132
rect 11883 7161 11933 7185
rect 11883 7137 11895 7161
rect 11919 7137 11933 7161
rect 11883 7108 11933 7137
rect 12091 7159 12141 7185
rect 12091 7133 12109 7159
rect 12135 7133 12141 7159
rect 12091 7108 12141 7133
rect 16518 7198 16568 7226
rect 16518 7178 16531 7198
rect 16551 7178 16568 7198
rect 16518 7149 16568 7178
rect 16731 7197 16781 7226
rect 16731 7173 16742 7197
rect 16766 7173 16781 7197
rect 16731 7149 16781 7173
rect 16939 7202 16989 7226
rect 16939 7178 16951 7202
rect 16975 7178 16989 7202
rect 16939 7149 16989 7178
rect 17147 7200 17197 7226
rect 17147 7174 17165 7200
rect 17191 7174 17197 7200
rect 17147 7149 17197 7174
rect 5439 7041 5489 7054
rect 5652 7041 5702 7054
rect 5860 7041 5910 7054
rect 6068 7041 6118 7054
rect 383 7000 433 7013
rect 596 7000 646 7013
rect 804 7000 854 7013
rect 1012 7000 1062 7013
rect 3870 6996 3920 7021
rect 3870 6970 3876 6996
rect 3902 6970 3920 6996
rect 3870 6944 3920 6970
rect 4078 6992 4128 7021
rect 4078 6968 4092 6992
rect 4116 6968 4128 6992
rect 4078 6944 4128 6968
rect 4286 6997 4336 7021
rect 4286 6973 4301 6997
rect 4325 6973 4336 6997
rect 4286 6944 4336 6973
rect 4499 6992 4549 7021
rect 4499 6972 4516 6992
rect 4536 6972 4549 6992
rect 4499 6944 4549 6972
rect 383 6872 433 6900
rect 383 6852 396 6872
rect 416 6852 433 6872
rect 383 6823 433 6852
rect 596 6871 646 6900
rect 596 6847 607 6871
rect 631 6847 646 6871
rect 596 6823 646 6847
rect 804 6876 854 6900
rect 804 6852 816 6876
rect 840 6852 854 6876
rect 804 6823 854 6852
rect 1012 6874 1062 6900
rect 1012 6848 1030 6874
rect 1056 6848 1062 6874
rect 1012 6823 1062 6848
rect 8926 7037 8976 7062
rect 8926 7011 8932 7037
rect 8958 7011 8976 7037
rect 8926 6985 8976 7011
rect 9134 7033 9184 7062
rect 9134 7009 9148 7033
rect 9172 7009 9184 7033
rect 9134 6985 9184 7009
rect 9342 7038 9392 7062
rect 9342 7014 9357 7038
rect 9381 7014 9392 7038
rect 9342 6985 9392 7014
rect 9555 7033 9605 7062
rect 9555 7013 9572 7033
rect 9592 7013 9605 7033
rect 12852 7105 12902 7118
rect 13060 7105 13110 7118
rect 13268 7105 13318 7118
rect 13481 7105 13531 7118
rect 11462 7050 11512 7066
rect 11675 7050 11725 7066
rect 11883 7050 11933 7066
rect 12091 7050 12141 7066
rect 13901 7068 13951 7084
rect 14109 7068 14159 7084
rect 14317 7068 14367 7084
rect 14530 7068 14580 7084
rect 17908 7146 17958 7159
rect 18116 7146 18166 7159
rect 18324 7146 18374 7159
rect 18537 7146 18587 7159
rect 16518 7091 16568 7107
rect 16731 7091 16781 7107
rect 16939 7091 16989 7107
rect 17147 7091 17197 7107
rect 18957 7109 19007 7125
rect 19165 7109 19215 7125
rect 19373 7109 19423 7125
rect 19586 7109 19636 7125
rect 15470 7046 15520 7059
rect 15683 7046 15733 7059
rect 15891 7046 15941 7059
rect 16099 7046 16149 7059
rect 9555 6985 9605 7013
rect 10414 7005 10464 7018
rect 10627 7005 10677 7018
rect 10835 7005 10885 7018
rect 11043 7005 11093 7018
rect 5439 6913 5489 6941
rect 5439 6893 5452 6913
rect 5472 6893 5489 6913
rect 3870 6831 3920 6844
rect 4078 6831 4128 6844
rect 4286 6831 4336 6844
rect 4499 6831 4549 6844
rect 5439 6864 5489 6893
rect 5652 6912 5702 6941
rect 5652 6888 5663 6912
rect 5687 6888 5702 6912
rect 5652 6864 5702 6888
rect 5860 6917 5910 6941
rect 5860 6893 5872 6917
rect 5896 6893 5910 6917
rect 5860 6864 5910 6893
rect 6068 6915 6118 6941
rect 6068 6889 6086 6915
rect 6112 6889 6118 6915
rect 6068 6864 6118 6889
rect 8926 6872 8976 6885
rect 9134 6872 9184 6885
rect 9342 6872 9392 6885
rect 9555 6872 9605 6885
rect 13901 7001 13951 7026
rect 13901 6975 13907 7001
rect 13933 6975 13951 7001
rect 13901 6949 13951 6975
rect 14109 6997 14159 7026
rect 14109 6973 14123 6997
rect 14147 6973 14159 6997
rect 14109 6949 14159 6973
rect 14317 7002 14367 7026
rect 14317 6978 14332 7002
rect 14356 6978 14367 7002
rect 14317 6949 14367 6978
rect 14530 6997 14580 7026
rect 14530 6977 14547 6997
rect 14567 6977 14580 6997
rect 14530 6949 14580 6977
rect 10414 6877 10464 6905
rect 5439 6806 5489 6822
rect 5652 6806 5702 6822
rect 5860 6806 5910 6822
rect 6068 6806 6118 6822
rect 10414 6857 10427 6877
rect 10447 6857 10464 6877
rect 383 6765 433 6781
rect 596 6765 646 6781
rect 804 6765 854 6781
rect 1012 6765 1062 6781
rect 6377 6797 6427 6810
rect 6590 6797 6640 6810
rect 6798 6797 6848 6810
rect 7006 6797 7056 6810
rect 1321 6756 1371 6769
rect 1534 6756 1584 6769
rect 1742 6756 1792 6769
rect 1950 6756 2000 6769
rect 2931 6753 2981 6769
rect 3139 6753 3189 6769
rect 3347 6753 3397 6769
rect 3560 6753 3610 6769
rect 2931 6686 2981 6711
rect 2931 6660 2937 6686
rect 2963 6660 2981 6686
rect 1321 6628 1371 6656
rect 1321 6608 1334 6628
rect 1354 6608 1371 6628
rect 1321 6579 1371 6608
rect 1534 6627 1584 6656
rect 1534 6603 1545 6627
rect 1569 6603 1584 6627
rect 1534 6579 1584 6603
rect 1742 6632 1792 6656
rect 1742 6608 1754 6632
rect 1778 6608 1792 6632
rect 1742 6579 1792 6608
rect 1950 6630 2000 6656
rect 2931 6634 2981 6660
rect 3139 6682 3189 6711
rect 3139 6658 3153 6682
rect 3177 6658 3189 6682
rect 3139 6634 3189 6658
rect 3347 6687 3397 6711
rect 3347 6663 3362 6687
rect 3386 6663 3397 6687
rect 3347 6634 3397 6663
rect 3560 6682 3610 6711
rect 3560 6662 3577 6682
rect 3597 6662 3610 6682
rect 3560 6634 3610 6662
rect 1950 6604 1968 6630
rect 1994 6604 2000 6630
rect 1950 6579 2000 6604
rect 1321 6521 1371 6537
rect 1534 6521 1584 6537
rect 1742 6521 1792 6537
rect 1950 6521 2000 6537
rect 7987 6794 8037 6810
rect 8195 6794 8245 6810
rect 8403 6794 8453 6810
rect 8616 6794 8666 6810
rect 10414 6828 10464 6857
rect 10627 6876 10677 6905
rect 10627 6852 10638 6876
rect 10662 6852 10677 6876
rect 10627 6828 10677 6852
rect 10835 6881 10885 6905
rect 10835 6857 10847 6881
rect 10871 6857 10885 6881
rect 10835 6828 10885 6857
rect 11043 6879 11093 6905
rect 11043 6853 11061 6879
rect 11087 6853 11093 6879
rect 11043 6828 11093 6853
rect 18957 7042 19007 7067
rect 18957 7016 18963 7042
rect 18989 7016 19007 7042
rect 18957 6990 19007 7016
rect 19165 7038 19215 7067
rect 19165 7014 19179 7038
rect 19203 7014 19215 7038
rect 19165 6990 19215 7014
rect 19373 7043 19423 7067
rect 19373 7019 19388 7043
rect 19412 7019 19423 7043
rect 19373 6990 19423 7019
rect 19586 7038 19636 7067
rect 19586 7018 19603 7038
rect 19623 7018 19636 7038
rect 19586 6990 19636 7018
rect 15470 6918 15520 6946
rect 15470 6898 15483 6918
rect 15503 6898 15520 6918
rect 13901 6836 13951 6849
rect 14109 6836 14159 6849
rect 14317 6836 14367 6849
rect 14530 6836 14580 6849
rect 15470 6869 15520 6898
rect 15683 6917 15733 6946
rect 15683 6893 15694 6917
rect 15718 6893 15733 6917
rect 15683 6869 15733 6893
rect 15891 6922 15941 6946
rect 15891 6898 15903 6922
rect 15927 6898 15941 6922
rect 15891 6869 15941 6898
rect 16099 6920 16149 6946
rect 16099 6894 16117 6920
rect 16143 6894 16149 6920
rect 16099 6869 16149 6894
rect 18957 6877 19007 6890
rect 19165 6877 19215 6890
rect 19373 6877 19423 6890
rect 19586 6877 19636 6890
rect 15470 6811 15520 6827
rect 15683 6811 15733 6827
rect 15891 6811 15941 6827
rect 16099 6811 16149 6827
rect 10414 6770 10464 6786
rect 10627 6770 10677 6786
rect 10835 6770 10885 6786
rect 11043 6770 11093 6786
rect 16408 6802 16458 6815
rect 16621 6802 16671 6815
rect 16829 6802 16879 6815
rect 17037 6802 17087 6815
rect 7987 6727 8037 6752
rect 7987 6701 7993 6727
rect 8019 6701 8037 6727
rect 6377 6669 6427 6697
rect 6377 6649 6390 6669
rect 6410 6649 6427 6669
rect 6377 6620 6427 6649
rect 6590 6668 6640 6697
rect 6590 6644 6601 6668
rect 6625 6644 6640 6668
rect 6590 6620 6640 6644
rect 6798 6673 6848 6697
rect 6798 6649 6810 6673
rect 6834 6649 6848 6673
rect 6798 6620 6848 6649
rect 7006 6671 7056 6697
rect 7987 6675 8037 6701
rect 8195 6723 8245 6752
rect 8195 6699 8209 6723
rect 8233 6699 8245 6723
rect 8195 6675 8245 6699
rect 8403 6728 8453 6752
rect 8403 6704 8418 6728
rect 8442 6704 8453 6728
rect 8403 6675 8453 6704
rect 8616 6723 8666 6752
rect 11352 6761 11402 6774
rect 11565 6761 11615 6774
rect 11773 6761 11823 6774
rect 11981 6761 12031 6774
rect 8616 6703 8633 6723
rect 8653 6703 8666 6723
rect 8616 6675 8666 6703
rect 7006 6645 7024 6671
rect 7050 6645 7056 6671
rect 7006 6620 7056 6645
rect 6377 6562 6427 6578
rect 6590 6562 6640 6578
rect 6798 6562 6848 6578
rect 7006 6562 7056 6578
rect 12962 6758 13012 6774
rect 13170 6758 13220 6774
rect 13378 6758 13428 6774
rect 13591 6758 13641 6774
rect 12962 6691 13012 6716
rect 12962 6665 12968 6691
rect 12994 6665 13012 6691
rect 11352 6633 11402 6661
rect 11352 6613 11365 6633
rect 11385 6613 11402 6633
rect 7987 6562 8037 6575
rect 8195 6562 8245 6575
rect 8403 6562 8453 6575
rect 8616 6562 8666 6575
rect 11352 6584 11402 6613
rect 11565 6632 11615 6661
rect 11565 6608 11576 6632
rect 11600 6608 11615 6632
rect 11565 6584 11615 6608
rect 11773 6637 11823 6661
rect 11773 6613 11785 6637
rect 11809 6613 11823 6637
rect 11773 6584 11823 6613
rect 11981 6635 12031 6661
rect 12962 6639 13012 6665
rect 13170 6687 13220 6716
rect 13170 6663 13184 6687
rect 13208 6663 13220 6687
rect 13170 6639 13220 6663
rect 13378 6692 13428 6716
rect 13378 6668 13393 6692
rect 13417 6668 13428 6692
rect 13378 6639 13428 6668
rect 13591 6687 13641 6716
rect 13591 6667 13608 6687
rect 13628 6667 13641 6687
rect 13591 6639 13641 6667
rect 11981 6609 11999 6635
rect 12025 6609 12031 6635
rect 11981 6584 12031 6609
rect 2931 6521 2981 6534
rect 3139 6521 3189 6534
rect 3347 6521 3397 6534
rect 3560 6521 3610 6534
rect 8925 6550 8975 6566
rect 9133 6550 9183 6566
rect 9341 6550 9391 6566
rect 9554 6550 9604 6566
rect 3869 6509 3919 6525
rect 4077 6509 4127 6525
rect 4285 6509 4335 6525
rect 4498 6509 4548 6525
rect 382 6446 432 6459
rect 595 6446 645 6459
rect 803 6446 853 6459
rect 1011 6446 1061 6459
rect 3869 6442 3919 6467
rect 3869 6416 3875 6442
rect 3901 6416 3919 6442
rect 3869 6390 3919 6416
rect 4077 6438 4127 6467
rect 4077 6414 4091 6438
rect 4115 6414 4127 6438
rect 4077 6390 4127 6414
rect 4285 6443 4335 6467
rect 4285 6419 4300 6443
rect 4324 6419 4335 6443
rect 4285 6390 4335 6419
rect 4498 6438 4548 6467
rect 5438 6487 5488 6500
rect 5651 6487 5701 6500
rect 5859 6487 5909 6500
rect 6067 6487 6117 6500
rect 4498 6418 4515 6438
rect 4535 6418 4548 6438
rect 4498 6390 4548 6418
rect 382 6318 432 6346
rect 382 6298 395 6318
rect 415 6298 432 6318
rect 382 6269 432 6298
rect 595 6317 645 6346
rect 595 6293 606 6317
rect 630 6293 645 6317
rect 595 6269 645 6293
rect 803 6322 853 6346
rect 803 6298 815 6322
rect 839 6298 853 6322
rect 803 6269 853 6298
rect 1011 6320 1061 6346
rect 1011 6294 1029 6320
rect 1055 6294 1061 6320
rect 1011 6269 1061 6294
rect 8925 6483 8975 6508
rect 8925 6457 8931 6483
rect 8957 6457 8975 6483
rect 8925 6431 8975 6457
rect 9133 6479 9183 6508
rect 9133 6455 9147 6479
rect 9171 6455 9183 6479
rect 9133 6431 9183 6455
rect 9341 6484 9391 6508
rect 9341 6460 9356 6484
rect 9380 6460 9391 6484
rect 9341 6431 9391 6460
rect 9554 6479 9604 6508
rect 11352 6526 11402 6542
rect 11565 6526 11615 6542
rect 11773 6526 11823 6542
rect 11981 6526 12031 6542
rect 18018 6799 18068 6815
rect 18226 6799 18276 6815
rect 18434 6799 18484 6815
rect 18647 6799 18697 6815
rect 18018 6732 18068 6757
rect 18018 6706 18024 6732
rect 18050 6706 18068 6732
rect 16408 6674 16458 6702
rect 16408 6654 16421 6674
rect 16441 6654 16458 6674
rect 16408 6625 16458 6654
rect 16621 6673 16671 6702
rect 16621 6649 16632 6673
rect 16656 6649 16671 6673
rect 16621 6625 16671 6649
rect 16829 6678 16879 6702
rect 16829 6654 16841 6678
rect 16865 6654 16879 6678
rect 16829 6625 16879 6654
rect 17037 6676 17087 6702
rect 18018 6680 18068 6706
rect 18226 6728 18276 6757
rect 18226 6704 18240 6728
rect 18264 6704 18276 6728
rect 18226 6680 18276 6704
rect 18434 6733 18484 6757
rect 18434 6709 18449 6733
rect 18473 6709 18484 6733
rect 18434 6680 18484 6709
rect 18647 6728 18697 6757
rect 18647 6708 18664 6728
rect 18684 6708 18697 6728
rect 18647 6680 18697 6708
rect 17037 6650 17055 6676
rect 17081 6650 17087 6676
rect 17037 6625 17087 6650
rect 16408 6567 16458 6583
rect 16621 6567 16671 6583
rect 16829 6567 16879 6583
rect 17037 6567 17087 6583
rect 18018 6567 18068 6580
rect 18226 6567 18276 6580
rect 18434 6567 18484 6580
rect 18647 6567 18697 6580
rect 12962 6526 13012 6539
rect 13170 6526 13220 6539
rect 13378 6526 13428 6539
rect 13591 6526 13641 6539
rect 18956 6555 19006 6571
rect 19164 6555 19214 6571
rect 19372 6555 19422 6571
rect 19585 6555 19635 6571
rect 9554 6459 9571 6479
rect 9591 6459 9604 6479
rect 13900 6514 13950 6530
rect 14108 6514 14158 6530
rect 14316 6514 14366 6530
rect 14529 6514 14579 6530
rect 9554 6431 9604 6459
rect 5438 6359 5488 6387
rect 5438 6339 5451 6359
rect 5471 6339 5488 6359
rect 5438 6310 5488 6339
rect 5651 6358 5701 6387
rect 5651 6334 5662 6358
rect 5686 6334 5701 6358
rect 5651 6310 5701 6334
rect 5859 6363 5909 6387
rect 5859 6339 5871 6363
rect 5895 6339 5909 6363
rect 5859 6310 5909 6339
rect 6067 6361 6117 6387
rect 6067 6335 6085 6361
rect 6111 6335 6117 6361
rect 6067 6310 6117 6335
rect 10413 6451 10463 6464
rect 10626 6451 10676 6464
rect 10834 6451 10884 6464
rect 11042 6451 11092 6464
rect 13900 6447 13950 6472
rect 13900 6421 13906 6447
rect 13932 6421 13950 6447
rect 13900 6395 13950 6421
rect 14108 6443 14158 6472
rect 14108 6419 14122 6443
rect 14146 6419 14158 6443
rect 14108 6395 14158 6419
rect 14316 6448 14366 6472
rect 14316 6424 14331 6448
rect 14355 6424 14366 6448
rect 14316 6395 14366 6424
rect 14529 6443 14579 6472
rect 15469 6492 15519 6505
rect 15682 6492 15732 6505
rect 15890 6492 15940 6505
rect 16098 6492 16148 6505
rect 14529 6423 14546 6443
rect 14566 6423 14579 6443
rect 14529 6395 14579 6423
rect 8925 6318 8975 6331
rect 9133 6318 9183 6331
rect 9341 6318 9391 6331
rect 9554 6318 9604 6331
rect 10413 6323 10463 6351
rect 3869 6277 3919 6290
rect 4077 6277 4127 6290
rect 4285 6277 4335 6290
rect 4498 6277 4548 6290
rect 2791 6242 2841 6258
rect 2999 6242 3049 6258
rect 3207 6242 3257 6258
rect 3420 6242 3470 6258
rect 382 6211 432 6227
rect 595 6211 645 6227
rect 803 6211 853 6227
rect 1011 6211 1061 6227
rect 7847 6283 7897 6299
rect 8055 6283 8105 6299
rect 8263 6283 8313 6299
rect 8476 6283 8526 6299
rect 5438 6252 5488 6268
rect 5651 6252 5701 6268
rect 5859 6252 5909 6268
rect 6067 6252 6117 6268
rect 10413 6303 10426 6323
rect 10446 6303 10463 6323
rect 10413 6274 10463 6303
rect 10626 6322 10676 6351
rect 10626 6298 10637 6322
rect 10661 6298 10676 6322
rect 10626 6274 10676 6298
rect 10834 6327 10884 6351
rect 10834 6303 10846 6327
rect 10870 6303 10884 6327
rect 10834 6274 10884 6303
rect 11042 6325 11092 6351
rect 11042 6299 11060 6325
rect 11086 6299 11092 6325
rect 11042 6274 11092 6299
rect 18956 6488 19006 6513
rect 18956 6462 18962 6488
rect 18988 6462 19006 6488
rect 18956 6436 19006 6462
rect 19164 6484 19214 6513
rect 19164 6460 19178 6484
rect 19202 6460 19214 6484
rect 19164 6436 19214 6460
rect 19372 6489 19422 6513
rect 19372 6465 19387 6489
rect 19411 6465 19422 6489
rect 19372 6436 19422 6465
rect 19585 6484 19635 6513
rect 19585 6464 19602 6484
rect 19622 6464 19635 6484
rect 19585 6436 19635 6464
rect 15469 6364 15519 6392
rect 15469 6344 15482 6364
rect 15502 6344 15519 6364
rect 15469 6315 15519 6344
rect 15682 6363 15732 6392
rect 15682 6339 15693 6363
rect 15717 6339 15732 6363
rect 15682 6315 15732 6339
rect 15890 6368 15940 6392
rect 15890 6344 15902 6368
rect 15926 6344 15940 6368
rect 15890 6315 15940 6344
rect 16098 6366 16148 6392
rect 16098 6340 16116 6366
rect 16142 6340 16148 6366
rect 16098 6315 16148 6340
rect 18956 6323 19006 6336
rect 19164 6323 19214 6336
rect 19372 6323 19422 6336
rect 19585 6323 19635 6336
rect 13900 6282 13950 6295
rect 14108 6282 14158 6295
rect 14316 6282 14366 6295
rect 14529 6282 14579 6295
rect 1462 6164 1512 6177
rect 1675 6164 1725 6177
rect 1883 6164 1933 6177
rect 2091 6164 2141 6177
rect 2791 6175 2841 6200
rect 2791 6149 2797 6175
rect 2823 6149 2841 6175
rect 2791 6123 2841 6149
rect 2999 6171 3049 6200
rect 2999 6147 3013 6171
rect 3037 6147 3049 6171
rect 2999 6123 3049 6147
rect 3207 6176 3257 6200
rect 3207 6152 3222 6176
rect 3246 6152 3257 6176
rect 3207 6123 3257 6152
rect 3420 6171 3470 6200
rect 6518 6205 6568 6218
rect 6731 6205 6781 6218
rect 6939 6205 6989 6218
rect 7147 6205 7197 6218
rect 7847 6216 7897 6241
rect 3420 6151 3437 6171
rect 3457 6151 3470 6171
rect 3420 6123 3470 6151
rect 1462 6036 1512 6064
rect 1462 6016 1475 6036
rect 1495 6016 1512 6036
rect 1462 5987 1512 6016
rect 1675 6035 1725 6064
rect 1675 6011 1686 6035
rect 1710 6011 1725 6035
rect 1675 5987 1725 6011
rect 1883 6040 1933 6064
rect 1883 6016 1895 6040
rect 1919 6016 1933 6040
rect 1883 5987 1933 6016
rect 2091 6038 2141 6064
rect 2091 6012 2109 6038
rect 2135 6012 2141 6038
rect 7847 6190 7853 6216
rect 7879 6190 7897 6216
rect 7847 6164 7897 6190
rect 8055 6212 8105 6241
rect 8055 6188 8069 6212
rect 8093 6188 8105 6212
rect 8055 6164 8105 6188
rect 8263 6217 8313 6241
rect 8263 6193 8278 6217
rect 8302 6193 8313 6217
rect 8263 6164 8313 6193
rect 8476 6212 8526 6241
rect 12822 6247 12872 6263
rect 13030 6247 13080 6263
rect 13238 6247 13288 6263
rect 13451 6247 13501 6263
rect 10413 6216 10463 6232
rect 10626 6216 10676 6232
rect 10834 6216 10884 6232
rect 11042 6216 11092 6232
rect 8476 6192 8493 6212
rect 8513 6192 8526 6212
rect 17878 6288 17928 6304
rect 18086 6288 18136 6304
rect 18294 6288 18344 6304
rect 18507 6288 18557 6304
rect 15469 6257 15519 6273
rect 15682 6257 15732 6273
rect 15890 6257 15940 6273
rect 16098 6257 16148 6273
rect 8476 6164 8526 6192
rect 6518 6077 6568 6105
rect 6518 6057 6531 6077
rect 6551 6057 6568 6077
rect 2091 5987 2141 6012
rect 2791 6010 2841 6023
rect 2999 6010 3049 6023
rect 3207 6010 3257 6023
rect 3420 6010 3470 6023
rect 6518 6028 6568 6057
rect 6731 6076 6781 6105
rect 6731 6052 6742 6076
rect 6766 6052 6781 6076
rect 6731 6028 6781 6052
rect 6939 6081 6989 6105
rect 6939 6057 6951 6081
rect 6975 6057 6989 6081
rect 6939 6028 6989 6057
rect 7147 6079 7197 6105
rect 7147 6053 7165 6079
rect 7191 6053 7197 6079
rect 11493 6169 11543 6182
rect 11706 6169 11756 6182
rect 11914 6169 11964 6182
rect 12122 6169 12172 6182
rect 12822 6180 12872 6205
rect 7147 6028 7197 6053
rect 7847 6051 7897 6064
rect 8055 6051 8105 6064
rect 8263 6051 8313 6064
rect 8476 6051 8526 6064
rect 12822 6154 12828 6180
rect 12854 6154 12872 6180
rect 12822 6128 12872 6154
rect 13030 6176 13080 6205
rect 13030 6152 13044 6176
rect 13068 6152 13080 6176
rect 13030 6128 13080 6152
rect 13238 6181 13288 6205
rect 13238 6157 13253 6181
rect 13277 6157 13288 6181
rect 13238 6128 13288 6157
rect 13451 6176 13501 6205
rect 16549 6210 16599 6223
rect 16762 6210 16812 6223
rect 16970 6210 17020 6223
rect 17178 6210 17228 6223
rect 17878 6221 17928 6246
rect 13451 6156 13468 6176
rect 13488 6156 13501 6176
rect 13451 6128 13501 6156
rect 11493 6041 11543 6069
rect 3871 5960 3921 5976
rect 4079 5960 4129 5976
rect 4287 5960 4337 5976
rect 4500 5960 4550 5976
rect 1462 5929 1512 5945
rect 1675 5929 1725 5945
rect 1883 5929 1933 5945
rect 2091 5929 2141 5945
rect 11493 6021 11506 6041
rect 11526 6021 11543 6041
rect 8927 6001 8977 6017
rect 9135 6001 9185 6017
rect 9343 6001 9393 6017
rect 9556 6001 9606 6017
rect 6518 5970 6568 5986
rect 6731 5970 6781 5986
rect 6939 5970 6989 5986
rect 7147 5970 7197 5986
rect 11493 5992 11543 6021
rect 11706 6040 11756 6069
rect 11706 6016 11717 6040
rect 11741 6016 11756 6040
rect 11706 5992 11756 6016
rect 11914 6045 11964 6069
rect 11914 6021 11926 6045
rect 11950 6021 11964 6045
rect 11914 5992 11964 6021
rect 12122 6043 12172 6069
rect 12122 6017 12140 6043
rect 12166 6017 12172 6043
rect 17878 6195 17884 6221
rect 17910 6195 17928 6221
rect 17878 6169 17928 6195
rect 18086 6217 18136 6246
rect 18086 6193 18100 6217
rect 18124 6193 18136 6217
rect 18086 6169 18136 6193
rect 18294 6222 18344 6246
rect 18294 6198 18309 6222
rect 18333 6198 18344 6222
rect 18294 6169 18344 6198
rect 18507 6217 18557 6246
rect 18507 6197 18524 6217
rect 18544 6197 18557 6217
rect 18507 6169 18557 6197
rect 16549 6082 16599 6110
rect 16549 6062 16562 6082
rect 16582 6062 16599 6082
rect 12122 5992 12172 6017
rect 12822 6015 12872 6028
rect 13030 6015 13080 6028
rect 13238 6015 13288 6028
rect 13451 6015 13501 6028
rect 16549 6033 16599 6062
rect 16762 6081 16812 6110
rect 16762 6057 16773 6081
rect 16797 6057 16812 6081
rect 16762 6033 16812 6057
rect 16970 6086 17020 6110
rect 16970 6062 16982 6086
rect 17006 6062 17020 6086
rect 16970 6033 17020 6062
rect 17178 6084 17228 6110
rect 17178 6058 17196 6084
rect 17222 6058 17228 6084
rect 17178 6033 17228 6058
rect 17878 6056 17928 6069
rect 18086 6056 18136 6069
rect 18294 6056 18344 6069
rect 18507 6056 18557 6069
rect 5440 5938 5490 5951
rect 5653 5938 5703 5951
rect 5861 5938 5911 5951
rect 6069 5938 6119 5951
rect 384 5897 434 5910
rect 597 5897 647 5910
rect 805 5897 855 5910
rect 1013 5897 1063 5910
rect 3871 5893 3921 5918
rect 3871 5867 3877 5893
rect 3903 5867 3921 5893
rect 3871 5841 3921 5867
rect 4079 5889 4129 5918
rect 4079 5865 4093 5889
rect 4117 5865 4129 5889
rect 4079 5841 4129 5865
rect 4287 5894 4337 5918
rect 4287 5870 4302 5894
rect 4326 5870 4337 5894
rect 4287 5841 4337 5870
rect 4500 5889 4550 5918
rect 4500 5869 4517 5889
rect 4537 5869 4550 5889
rect 4500 5841 4550 5869
rect 384 5769 434 5797
rect 384 5749 397 5769
rect 417 5749 434 5769
rect 384 5720 434 5749
rect 597 5768 647 5797
rect 597 5744 608 5768
rect 632 5744 647 5768
rect 597 5720 647 5744
rect 805 5773 855 5797
rect 805 5749 817 5773
rect 841 5749 855 5773
rect 805 5720 855 5749
rect 1013 5771 1063 5797
rect 1013 5745 1031 5771
rect 1057 5745 1063 5771
rect 1013 5720 1063 5745
rect 8927 5934 8977 5959
rect 8927 5908 8933 5934
rect 8959 5908 8977 5934
rect 8927 5882 8977 5908
rect 9135 5930 9185 5959
rect 9135 5906 9149 5930
rect 9173 5906 9185 5930
rect 9135 5882 9185 5906
rect 9343 5935 9393 5959
rect 9343 5911 9358 5935
rect 9382 5911 9393 5935
rect 9343 5882 9393 5911
rect 9556 5930 9606 5959
rect 9556 5910 9573 5930
rect 9593 5910 9606 5930
rect 13902 5965 13952 5981
rect 14110 5965 14160 5981
rect 14318 5965 14368 5981
rect 14531 5965 14581 5981
rect 11493 5934 11543 5950
rect 11706 5934 11756 5950
rect 11914 5934 11964 5950
rect 12122 5934 12172 5950
rect 18958 6006 19008 6022
rect 19166 6006 19216 6022
rect 19374 6006 19424 6022
rect 19587 6006 19637 6022
rect 16549 5975 16599 5991
rect 16762 5975 16812 5991
rect 16970 5975 17020 5991
rect 17178 5975 17228 5991
rect 15471 5943 15521 5956
rect 15684 5943 15734 5956
rect 15892 5943 15942 5956
rect 16100 5943 16150 5956
rect 9556 5882 9606 5910
rect 10415 5902 10465 5915
rect 10628 5902 10678 5915
rect 10836 5902 10886 5915
rect 11044 5902 11094 5915
rect 5440 5810 5490 5838
rect 5440 5790 5453 5810
rect 5473 5790 5490 5810
rect 3871 5728 3921 5741
rect 4079 5728 4129 5741
rect 4287 5728 4337 5741
rect 4500 5728 4550 5741
rect 5440 5761 5490 5790
rect 5653 5809 5703 5838
rect 5653 5785 5664 5809
rect 5688 5785 5703 5809
rect 5653 5761 5703 5785
rect 5861 5814 5911 5838
rect 5861 5790 5873 5814
rect 5897 5790 5911 5814
rect 5861 5761 5911 5790
rect 6069 5812 6119 5838
rect 6069 5786 6087 5812
rect 6113 5786 6119 5812
rect 6069 5761 6119 5786
rect 8927 5769 8977 5782
rect 9135 5769 9185 5782
rect 9343 5769 9393 5782
rect 9556 5769 9606 5782
rect 13902 5898 13952 5923
rect 13902 5872 13908 5898
rect 13934 5872 13952 5898
rect 13902 5846 13952 5872
rect 14110 5894 14160 5923
rect 14110 5870 14124 5894
rect 14148 5870 14160 5894
rect 14110 5846 14160 5870
rect 14318 5899 14368 5923
rect 14318 5875 14333 5899
rect 14357 5875 14368 5899
rect 14318 5846 14368 5875
rect 14531 5894 14581 5923
rect 14531 5874 14548 5894
rect 14568 5874 14581 5894
rect 14531 5846 14581 5874
rect 10415 5774 10465 5802
rect 5440 5703 5490 5719
rect 5653 5703 5703 5719
rect 5861 5703 5911 5719
rect 6069 5703 6119 5719
rect 10415 5754 10428 5774
rect 10448 5754 10465 5774
rect 384 5662 434 5678
rect 597 5662 647 5678
rect 805 5662 855 5678
rect 1013 5662 1063 5678
rect 6378 5694 6428 5707
rect 6591 5694 6641 5707
rect 6799 5694 6849 5707
rect 7007 5694 7057 5707
rect 1322 5653 1372 5666
rect 1535 5653 1585 5666
rect 1743 5653 1793 5666
rect 1951 5653 2001 5666
rect 2932 5650 2982 5666
rect 3140 5650 3190 5666
rect 3348 5650 3398 5666
rect 3561 5650 3611 5666
rect 2932 5583 2982 5608
rect 2932 5557 2938 5583
rect 2964 5557 2982 5583
rect 1322 5525 1372 5553
rect 1322 5505 1335 5525
rect 1355 5505 1372 5525
rect 1322 5476 1372 5505
rect 1535 5524 1585 5553
rect 1535 5500 1546 5524
rect 1570 5500 1585 5524
rect 1535 5476 1585 5500
rect 1743 5529 1793 5553
rect 1743 5505 1755 5529
rect 1779 5505 1793 5529
rect 1743 5476 1793 5505
rect 1951 5527 2001 5553
rect 2932 5531 2982 5557
rect 3140 5579 3190 5608
rect 3140 5555 3154 5579
rect 3178 5555 3190 5579
rect 3140 5531 3190 5555
rect 3348 5584 3398 5608
rect 3348 5560 3363 5584
rect 3387 5560 3398 5584
rect 3348 5531 3398 5560
rect 3561 5579 3611 5608
rect 3561 5559 3578 5579
rect 3598 5559 3611 5579
rect 3561 5531 3611 5559
rect 1951 5501 1969 5527
rect 1995 5501 2001 5527
rect 1951 5476 2001 5501
rect 1322 5418 1372 5434
rect 1535 5418 1585 5434
rect 1743 5418 1793 5434
rect 1951 5418 2001 5434
rect 7988 5691 8038 5707
rect 8196 5691 8246 5707
rect 8404 5691 8454 5707
rect 8617 5691 8667 5707
rect 10415 5725 10465 5754
rect 10628 5773 10678 5802
rect 10628 5749 10639 5773
rect 10663 5749 10678 5773
rect 10628 5725 10678 5749
rect 10836 5778 10886 5802
rect 10836 5754 10848 5778
rect 10872 5754 10886 5778
rect 10836 5725 10886 5754
rect 11044 5776 11094 5802
rect 11044 5750 11062 5776
rect 11088 5750 11094 5776
rect 11044 5725 11094 5750
rect 18958 5939 19008 5964
rect 18958 5913 18964 5939
rect 18990 5913 19008 5939
rect 18958 5887 19008 5913
rect 19166 5935 19216 5964
rect 19166 5911 19180 5935
rect 19204 5911 19216 5935
rect 19166 5887 19216 5911
rect 19374 5940 19424 5964
rect 19374 5916 19389 5940
rect 19413 5916 19424 5940
rect 19374 5887 19424 5916
rect 19587 5935 19637 5964
rect 19587 5915 19604 5935
rect 19624 5915 19637 5935
rect 19587 5887 19637 5915
rect 15471 5815 15521 5843
rect 15471 5795 15484 5815
rect 15504 5795 15521 5815
rect 13902 5733 13952 5746
rect 14110 5733 14160 5746
rect 14318 5733 14368 5746
rect 14531 5733 14581 5746
rect 15471 5766 15521 5795
rect 15684 5814 15734 5843
rect 15684 5790 15695 5814
rect 15719 5790 15734 5814
rect 15684 5766 15734 5790
rect 15892 5819 15942 5843
rect 15892 5795 15904 5819
rect 15928 5795 15942 5819
rect 15892 5766 15942 5795
rect 16100 5817 16150 5843
rect 16100 5791 16118 5817
rect 16144 5791 16150 5817
rect 16100 5766 16150 5791
rect 18958 5774 19008 5787
rect 19166 5774 19216 5787
rect 19374 5774 19424 5787
rect 19587 5774 19637 5787
rect 15471 5708 15521 5724
rect 15684 5708 15734 5724
rect 15892 5708 15942 5724
rect 16100 5708 16150 5724
rect 10415 5667 10465 5683
rect 10628 5667 10678 5683
rect 10836 5667 10886 5683
rect 11044 5667 11094 5683
rect 16409 5699 16459 5712
rect 16622 5699 16672 5712
rect 16830 5699 16880 5712
rect 17038 5699 17088 5712
rect 7988 5624 8038 5649
rect 7988 5598 7994 5624
rect 8020 5598 8038 5624
rect 6378 5566 6428 5594
rect 6378 5546 6391 5566
rect 6411 5546 6428 5566
rect 6378 5517 6428 5546
rect 6591 5565 6641 5594
rect 6591 5541 6602 5565
rect 6626 5541 6641 5565
rect 6591 5517 6641 5541
rect 6799 5570 6849 5594
rect 6799 5546 6811 5570
rect 6835 5546 6849 5570
rect 6799 5517 6849 5546
rect 7007 5568 7057 5594
rect 7988 5572 8038 5598
rect 8196 5620 8246 5649
rect 8196 5596 8210 5620
rect 8234 5596 8246 5620
rect 8196 5572 8246 5596
rect 8404 5625 8454 5649
rect 8404 5601 8419 5625
rect 8443 5601 8454 5625
rect 8404 5572 8454 5601
rect 8617 5620 8667 5649
rect 11353 5658 11403 5671
rect 11566 5658 11616 5671
rect 11774 5658 11824 5671
rect 11982 5658 12032 5671
rect 8617 5600 8634 5620
rect 8654 5600 8667 5620
rect 8617 5572 8667 5600
rect 7007 5542 7025 5568
rect 7051 5542 7057 5568
rect 7007 5517 7057 5542
rect 6378 5459 6428 5475
rect 6591 5459 6641 5475
rect 6799 5459 6849 5475
rect 7007 5459 7057 5475
rect 12963 5655 13013 5671
rect 13171 5655 13221 5671
rect 13379 5655 13429 5671
rect 13592 5655 13642 5671
rect 12963 5588 13013 5613
rect 12963 5562 12969 5588
rect 12995 5562 13013 5588
rect 11353 5530 11403 5558
rect 11353 5510 11366 5530
rect 11386 5510 11403 5530
rect 7988 5459 8038 5472
rect 8196 5459 8246 5472
rect 8404 5459 8454 5472
rect 8617 5459 8667 5472
rect 11353 5481 11403 5510
rect 11566 5529 11616 5558
rect 11566 5505 11577 5529
rect 11601 5505 11616 5529
rect 11566 5481 11616 5505
rect 11774 5534 11824 5558
rect 11774 5510 11786 5534
rect 11810 5510 11824 5534
rect 11774 5481 11824 5510
rect 11982 5532 12032 5558
rect 12963 5536 13013 5562
rect 13171 5584 13221 5613
rect 13171 5560 13185 5584
rect 13209 5560 13221 5584
rect 13171 5536 13221 5560
rect 13379 5589 13429 5613
rect 13379 5565 13394 5589
rect 13418 5565 13429 5589
rect 13379 5536 13429 5565
rect 13592 5584 13642 5613
rect 13592 5564 13609 5584
rect 13629 5564 13642 5584
rect 13592 5536 13642 5564
rect 11982 5506 12000 5532
rect 12026 5506 12032 5532
rect 11982 5481 12032 5506
rect 2932 5418 2982 5431
rect 3140 5418 3190 5431
rect 3348 5418 3398 5431
rect 3561 5418 3611 5431
rect 8926 5447 8976 5463
rect 9134 5447 9184 5463
rect 9342 5447 9392 5463
rect 9555 5447 9605 5463
rect 3870 5406 3920 5422
rect 4078 5406 4128 5422
rect 4286 5406 4336 5422
rect 4499 5406 4549 5422
rect 383 5343 433 5356
rect 596 5343 646 5356
rect 804 5343 854 5356
rect 1012 5343 1062 5356
rect 3870 5339 3920 5364
rect 3870 5313 3876 5339
rect 3902 5313 3920 5339
rect 3870 5287 3920 5313
rect 4078 5335 4128 5364
rect 4078 5311 4092 5335
rect 4116 5311 4128 5335
rect 4078 5287 4128 5311
rect 4286 5340 4336 5364
rect 4286 5316 4301 5340
rect 4325 5316 4336 5340
rect 4286 5287 4336 5316
rect 4499 5335 4549 5364
rect 5439 5384 5489 5397
rect 5652 5384 5702 5397
rect 5860 5384 5910 5397
rect 6068 5384 6118 5397
rect 4499 5315 4516 5335
rect 4536 5315 4549 5335
rect 4499 5287 4549 5315
rect 383 5215 433 5243
rect 383 5195 396 5215
rect 416 5195 433 5215
rect 383 5166 433 5195
rect 596 5214 646 5243
rect 596 5190 607 5214
rect 631 5190 646 5214
rect 596 5166 646 5190
rect 804 5219 854 5243
rect 804 5195 816 5219
rect 840 5195 854 5219
rect 804 5166 854 5195
rect 1012 5217 1062 5243
rect 1012 5191 1030 5217
rect 1056 5191 1062 5217
rect 1012 5166 1062 5191
rect 8926 5380 8976 5405
rect 8926 5354 8932 5380
rect 8958 5354 8976 5380
rect 8926 5328 8976 5354
rect 9134 5376 9184 5405
rect 9134 5352 9148 5376
rect 9172 5352 9184 5376
rect 9134 5328 9184 5352
rect 9342 5381 9392 5405
rect 9342 5357 9357 5381
rect 9381 5357 9392 5381
rect 9342 5328 9392 5357
rect 9555 5376 9605 5405
rect 11353 5423 11403 5439
rect 11566 5423 11616 5439
rect 11774 5423 11824 5439
rect 11982 5423 12032 5439
rect 18019 5696 18069 5712
rect 18227 5696 18277 5712
rect 18435 5696 18485 5712
rect 18648 5696 18698 5712
rect 18019 5629 18069 5654
rect 18019 5603 18025 5629
rect 18051 5603 18069 5629
rect 16409 5571 16459 5599
rect 16409 5551 16422 5571
rect 16442 5551 16459 5571
rect 16409 5522 16459 5551
rect 16622 5570 16672 5599
rect 16622 5546 16633 5570
rect 16657 5546 16672 5570
rect 16622 5522 16672 5546
rect 16830 5575 16880 5599
rect 16830 5551 16842 5575
rect 16866 5551 16880 5575
rect 16830 5522 16880 5551
rect 17038 5573 17088 5599
rect 18019 5577 18069 5603
rect 18227 5625 18277 5654
rect 18227 5601 18241 5625
rect 18265 5601 18277 5625
rect 18227 5577 18277 5601
rect 18435 5630 18485 5654
rect 18435 5606 18450 5630
rect 18474 5606 18485 5630
rect 18435 5577 18485 5606
rect 18648 5625 18698 5654
rect 18648 5605 18665 5625
rect 18685 5605 18698 5625
rect 18648 5577 18698 5605
rect 17038 5547 17056 5573
rect 17082 5547 17088 5573
rect 17038 5522 17088 5547
rect 16409 5464 16459 5480
rect 16622 5464 16672 5480
rect 16830 5464 16880 5480
rect 17038 5464 17088 5480
rect 18019 5464 18069 5477
rect 18227 5464 18277 5477
rect 18435 5464 18485 5477
rect 18648 5464 18698 5477
rect 12963 5423 13013 5436
rect 13171 5423 13221 5436
rect 13379 5423 13429 5436
rect 13592 5423 13642 5436
rect 18957 5452 19007 5468
rect 19165 5452 19215 5468
rect 19373 5452 19423 5468
rect 19586 5452 19636 5468
rect 9555 5356 9572 5376
rect 9592 5356 9605 5376
rect 13901 5411 13951 5427
rect 14109 5411 14159 5427
rect 14317 5411 14367 5427
rect 14530 5411 14580 5427
rect 9555 5328 9605 5356
rect 5439 5256 5489 5284
rect 5439 5236 5452 5256
rect 5472 5236 5489 5256
rect 5439 5207 5489 5236
rect 5652 5255 5702 5284
rect 5652 5231 5663 5255
rect 5687 5231 5702 5255
rect 5652 5207 5702 5231
rect 5860 5260 5910 5284
rect 5860 5236 5872 5260
rect 5896 5236 5910 5260
rect 5860 5207 5910 5236
rect 6068 5258 6118 5284
rect 6068 5232 6086 5258
rect 6112 5232 6118 5258
rect 6068 5207 6118 5232
rect 10414 5348 10464 5361
rect 10627 5348 10677 5361
rect 10835 5348 10885 5361
rect 11043 5348 11093 5361
rect 13901 5344 13951 5369
rect 13901 5318 13907 5344
rect 13933 5318 13951 5344
rect 13901 5292 13951 5318
rect 14109 5340 14159 5369
rect 14109 5316 14123 5340
rect 14147 5316 14159 5340
rect 14109 5292 14159 5316
rect 14317 5345 14367 5369
rect 14317 5321 14332 5345
rect 14356 5321 14367 5345
rect 14317 5292 14367 5321
rect 14530 5340 14580 5369
rect 15470 5389 15520 5402
rect 15683 5389 15733 5402
rect 15891 5389 15941 5402
rect 16099 5389 16149 5402
rect 14530 5320 14547 5340
rect 14567 5320 14580 5340
rect 14530 5292 14580 5320
rect 3870 5174 3920 5187
rect 4078 5174 4128 5187
rect 4286 5174 4336 5187
rect 4499 5174 4549 5187
rect 383 5108 433 5124
rect 596 5108 646 5124
rect 804 5108 854 5124
rect 1012 5108 1062 5124
rect 2823 5120 2873 5136
rect 3031 5120 3081 5136
rect 3239 5120 3289 5136
rect 3452 5120 3502 5136
rect 1431 5080 1481 5093
rect 1644 5080 1694 5093
rect 1852 5080 1902 5093
rect 2060 5080 2110 5093
rect 8926 5215 8976 5228
rect 9134 5215 9184 5228
rect 9342 5215 9392 5228
rect 9555 5215 9605 5228
rect 10414 5220 10464 5248
rect 5439 5149 5489 5165
rect 5652 5149 5702 5165
rect 5860 5149 5910 5165
rect 6068 5149 6118 5165
rect 7879 5161 7929 5177
rect 8087 5161 8137 5177
rect 8295 5161 8345 5177
rect 8508 5161 8558 5177
rect 6487 5121 6537 5134
rect 6700 5121 6750 5134
rect 6908 5121 6958 5134
rect 7116 5121 7166 5134
rect 2823 5053 2873 5078
rect 2823 5027 2829 5053
rect 2855 5027 2873 5053
rect 2823 5001 2873 5027
rect 3031 5049 3081 5078
rect 3031 5025 3045 5049
rect 3069 5025 3081 5049
rect 3031 5001 3081 5025
rect 3239 5054 3289 5078
rect 3239 5030 3254 5054
rect 3278 5030 3289 5054
rect 3239 5001 3289 5030
rect 3452 5049 3502 5078
rect 3452 5029 3469 5049
rect 3489 5029 3502 5049
rect 3452 5001 3502 5029
rect 10414 5200 10427 5220
rect 10447 5200 10464 5220
rect 10414 5171 10464 5200
rect 10627 5219 10677 5248
rect 10627 5195 10638 5219
rect 10662 5195 10677 5219
rect 10627 5171 10677 5195
rect 10835 5224 10885 5248
rect 10835 5200 10847 5224
rect 10871 5200 10885 5224
rect 10835 5171 10885 5200
rect 11043 5222 11093 5248
rect 11043 5196 11061 5222
rect 11087 5196 11093 5222
rect 11043 5171 11093 5196
rect 18957 5385 19007 5410
rect 18957 5359 18963 5385
rect 18989 5359 19007 5385
rect 18957 5333 19007 5359
rect 19165 5381 19215 5410
rect 19165 5357 19179 5381
rect 19203 5357 19215 5381
rect 19165 5333 19215 5357
rect 19373 5386 19423 5410
rect 19373 5362 19388 5386
rect 19412 5362 19423 5386
rect 19373 5333 19423 5362
rect 19586 5381 19636 5410
rect 19586 5361 19603 5381
rect 19623 5361 19636 5381
rect 19586 5333 19636 5361
rect 15470 5261 15520 5289
rect 15470 5241 15483 5261
rect 15503 5241 15520 5261
rect 15470 5212 15520 5241
rect 15683 5260 15733 5289
rect 15683 5236 15694 5260
rect 15718 5236 15733 5260
rect 15683 5212 15733 5236
rect 15891 5265 15941 5289
rect 15891 5241 15903 5265
rect 15927 5241 15941 5265
rect 15891 5212 15941 5241
rect 16099 5263 16149 5289
rect 16099 5237 16117 5263
rect 16143 5237 16149 5263
rect 16099 5212 16149 5237
rect 7879 5094 7929 5119
rect 7879 5068 7885 5094
rect 7911 5068 7929 5094
rect 7879 5042 7929 5068
rect 8087 5090 8137 5119
rect 8087 5066 8101 5090
rect 8125 5066 8137 5090
rect 8087 5042 8137 5066
rect 8295 5095 8345 5119
rect 8295 5071 8310 5095
rect 8334 5071 8345 5095
rect 8295 5042 8345 5071
rect 8508 5090 8558 5119
rect 13901 5179 13951 5192
rect 14109 5179 14159 5192
rect 14317 5179 14367 5192
rect 14530 5179 14580 5192
rect 10414 5113 10464 5129
rect 10627 5113 10677 5129
rect 10835 5113 10885 5129
rect 11043 5113 11093 5129
rect 12854 5125 12904 5141
rect 13062 5125 13112 5141
rect 13270 5125 13320 5141
rect 13483 5125 13533 5141
rect 8508 5070 8525 5090
rect 8545 5070 8558 5090
rect 8508 5042 8558 5070
rect 11462 5085 11512 5098
rect 11675 5085 11725 5098
rect 11883 5085 11933 5098
rect 12091 5085 12141 5098
rect 1431 4952 1481 4980
rect 1431 4932 1444 4952
rect 1464 4932 1481 4952
rect 1431 4903 1481 4932
rect 1644 4951 1694 4980
rect 1644 4927 1655 4951
rect 1679 4927 1694 4951
rect 1644 4903 1694 4927
rect 1852 4956 1902 4980
rect 1852 4932 1864 4956
rect 1888 4932 1902 4956
rect 1852 4903 1902 4932
rect 2060 4954 2110 4980
rect 2060 4928 2078 4954
rect 2104 4928 2110 4954
rect 2060 4903 2110 4928
rect 6487 4993 6537 5021
rect 6487 4973 6500 4993
rect 6520 4973 6537 4993
rect 6487 4944 6537 4973
rect 6700 4992 6750 5021
rect 6700 4968 6711 4992
rect 6735 4968 6750 4992
rect 6700 4944 6750 4968
rect 6908 4997 6958 5021
rect 6908 4973 6920 4997
rect 6944 4973 6958 4997
rect 6908 4944 6958 4973
rect 7116 4995 7166 5021
rect 7116 4969 7134 4995
rect 7160 4969 7166 4995
rect 7116 4944 7166 4969
rect 2823 4888 2873 4901
rect 3031 4888 3081 4901
rect 3239 4888 3289 4901
rect 3452 4888 3502 4901
rect 1431 4845 1481 4861
rect 1644 4845 1694 4861
rect 1852 4845 1902 4861
rect 2060 4845 2110 4861
rect 3871 4857 3921 4873
rect 4079 4857 4129 4873
rect 4287 4857 4337 4873
rect 4500 4857 4550 4873
rect 384 4794 434 4807
rect 597 4794 647 4807
rect 805 4794 855 4807
rect 1013 4794 1063 4807
rect 18957 5220 19007 5233
rect 19165 5220 19215 5233
rect 19373 5220 19423 5233
rect 19586 5220 19636 5233
rect 15470 5154 15520 5170
rect 15683 5154 15733 5170
rect 15891 5154 15941 5170
rect 16099 5154 16149 5170
rect 17910 5166 17960 5182
rect 18118 5166 18168 5182
rect 18326 5166 18376 5182
rect 18539 5166 18589 5182
rect 16518 5126 16568 5139
rect 16731 5126 16781 5139
rect 16939 5126 16989 5139
rect 17147 5126 17197 5139
rect 12854 5058 12904 5083
rect 12854 5032 12860 5058
rect 12886 5032 12904 5058
rect 12854 5006 12904 5032
rect 13062 5054 13112 5083
rect 13062 5030 13076 5054
rect 13100 5030 13112 5054
rect 13062 5006 13112 5030
rect 13270 5059 13320 5083
rect 13270 5035 13285 5059
rect 13309 5035 13320 5059
rect 13270 5006 13320 5035
rect 13483 5054 13533 5083
rect 13483 5034 13500 5054
rect 13520 5034 13533 5054
rect 13483 5006 13533 5034
rect 17910 5099 17960 5124
rect 17910 5073 17916 5099
rect 17942 5073 17960 5099
rect 17910 5047 17960 5073
rect 18118 5095 18168 5124
rect 18118 5071 18132 5095
rect 18156 5071 18168 5095
rect 18118 5047 18168 5071
rect 18326 5100 18376 5124
rect 18326 5076 18341 5100
rect 18365 5076 18376 5100
rect 18326 5047 18376 5076
rect 18539 5095 18589 5124
rect 18539 5075 18556 5095
rect 18576 5075 18589 5095
rect 18539 5047 18589 5075
rect 7879 4929 7929 4942
rect 8087 4929 8137 4942
rect 8295 4929 8345 4942
rect 8508 4929 8558 4942
rect 11462 4957 11512 4985
rect 11462 4937 11475 4957
rect 11495 4937 11512 4957
rect 6487 4886 6537 4902
rect 6700 4886 6750 4902
rect 6908 4886 6958 4902
rect 7116 4886 7166 4902
rect 8927 4898 8977 4914
rect 9135 4898 9185 4914
rect 9343 4898 9393 4914
rect 9556 4898 9606 4914
rect 5440 4835 5490 4848
rect 5653 4835 5703 4848
rect 5861 4835 5911 4848
rect 6069 4835 6119 4848
rect 11462 4908 11512 4937
rect 11675 4956 11725 4985
rect 11675 4932 11686 4956
rect 11710 4932 11725 4956
rect 11675 4908 11725 4932
rect 11883 4961 11933 4985
rect 11883 4937 11895 4961
rect 11919 4937 11933 4961
rect 11883 4908 11933 4937
rect 12091 4959 12141 4985
rect 12091 4933 12109 4959
rect 12135 4933 12141 4959
rect 12091 4908 12141 4933
rect 3871 4790 3921 4815
rect 3871 4764 3877 4790
rect 3903 4764 3921 4790
rect 3871 4738 3921 4764
rect 4079 4786 4129 4815
rect 4079 4762 4093 4786
rect 4117 4762 4129 4786
rect 4079 4738 4129 4762
rect 4287 4791 4337 4815
rect 4287 4767 4302 4791
rect 4326 4767 4337 4791
rect 4287 4738 4337 4767
rect 4500 4786 4550 4815
rect 4500 4766 4517 4786
rect 4537 4766 4550 4786
rect 4500 4738 4550 4766
rect 384 4666 434 4694
rect 384 4646 397 4666
rect 417 4646 434 4666
rect 384 4617 434 4646
rect 597 4665 647 4694
rect 597 4641 608 4665
rect 632 4641 647 4665
rect 597 4617 647 4641
rect 805 4670 855 4694
rect 805 4646 817 4670
rect 841 4646 855 4670
rect 805 4617 855 4646
rect 1013 4668 1063 4694
rect 1013 4642 1031 4668
rect 1057 4642 1063 4668
rect 1013 4617 1063 4642
rect 8927 4831 8977 4856
rect 8927 4805 8933 4831
rect 8959 4805 8977 4831
rect 8927 4779 8977 4805
rect 9135 4827 9185 4856
rect 9135 4803 9149 4827
rect 9173 4803 9185 4827
rect 9135 4779 9185 4803
rect 9343 4832 9393 4856
rect 9343 4808 9358 4832
rect 9382 4808 9393 4832
rect 9343 4779 9393 4808
rect 9556 4827 9606 4856
rect 9556 4807 9573 4827
rect 9593 4807 9606 4827
rect 16518 4998 16568 5026
rect 16518 4978 16531 4998
rect 16551 4978 16568 4998
rect 16518 4949 16568 4978
rect 16731 4997 16781 5026
rect 16731 4973 16742 4997
rect 16766 4973 16781 4997
rect 16731 4949 16781 4973
rect 16939 5002 16989 5026
rect 16939 4978 16951 5002
rect 16975 4978 16989 5002
rect 16939 4949 16989 4978
rect 17147 5000 17197 5026
rect 17147 4974 17165 5000
rect 17191 4974 17197 5000
rect 17147 4949 17197 4974
rect 12854 4893 12904 4906
rect 13062 4893 13112 4906
rect 13270 4893 13320 4906
rect 13483 4893 13533 4906
rect 11462 4850 11512 4866
rect 11675 4850 11725 4866
rect 11883 4850 11933 4866
rect 12091 4850 12141 4866
rect 13902 4862 13952 4878
rect 14110 4862 14160 4878
rect 14318 4862 14368 4878
rect 14531 4862 14581 4878
rect 9556 4779 9606 4807
rect 10415 4799 10465 4812
rect 10628 4799 10678 4812
rect 10836 4799 10886 4812
rect 11044 4799 11094 4812
rect 17910 4934 17960 4947
rect 18118 4934 18168 4947
rect 18326 4934 18376 4947
rect 18539 4934 18589 4947
rect 16518 4891 16568 4907
rect 16731 4891 16781 4907
rect 16939 4891 16989 4907
rect 17147 4891 17197 4907
rect 18958 4903 19008 4919
rect 19166 4903 19216 4919
rect 19374 4903 19424 4919
rect 19587 4903 19637 4919
rect 15471 4840 15521 4853
rect 15684 4840 15734 4853
rect 15892 4840 15942 4853
rect 16100 4840 16150 4853
rect 5440 4707 5490 4735
rect 5440 4687 5453 4707
rect 5473 4687 5490 4707
rect 3871 4625 3921 4638
rect 4079 4625 4129 4638
rect 4287 4625 4337 4638
rect 4500 4625 4550 4638
rect 5440 4658 5490 4687
rect 5653 4706 5703 4735
rect 5653 4682 5664 4706
rect 5688 4682 5703 4706
rect 5653 4658 5703 4682
rect 5861 4711 5911 4735
rect 5861 4687 5873 4711
rect 5897 4687 5911 4711
rect 5861 4658 5911 4687
rect 6069 4709 6119 4735
rect 6069 4683 6087 4709
rect 6113 4683 6119 4709
rect 6069 4658 6119 4683
rect 8927 4666 8977 4679
rect 9135 4666 9185 4679
rect 9343 4666 9393 4679
rect 9556 4666 9606 4679
rect 13902 4795 13952 4820
rect 13902 4769 13908 4795
rect 13934 4769 13952 4795
rect 13902 4743 13952 4769
rect 14110 4791 14160 4820
rect 14110 4767 14124 4791
rect 14148 4767 14160 4791
rect 14110 4743 14160 4767
rect 14318 4796 14368 4820
rect 14318 4772 14333 4796
rect 14357 4772 14368 4796
rect 14318 4743 14368 4772
rect 14531 4791 14581 4820
rect 14531 4771 14548 4791
rect 14568 4771 14581 4791
rect 14531 4743 14581 4771
rect 10415 4671 10465 4699
rect 5440 4600 5490 4616
rect 5653 4600 5703 4616
rect 5861 4600 5911 4616
rect 6069 4600 6119 4616
rect 10415 4651 10428 4671
rect 10448 4651 10465 4671
rect 384 4559 434 4575
rect 597 4559 647 4575
rect 805 4559 855 4575
rect 1013 4559 1063 4575
rect 6378 4591 6428 4604
rect 6591 4591 6641 4604
rect 6799 4591 6849 4604
rect 7007 4591 7057 4604
rect 1322 4550 1372 4563
rect 1535 4550 1585 4563
rect 1743 4550 1793 4563
rect 1951 4550 2001 4563
rect 2932 4547 2982 4563
rect 3140 4547 3190 4563
rect 3348 4547 3398 4563
rect 3561 4547 3611 4563
rect 2932 4480 2982 4505
rect 2932 4454 2938 4480
rect 2964 4454 2982 4480
rect 1322 4422 1372 4450
rect 1322 4402 1335 4422
rect 1355 4402 1372 4422
rect 1322 4373 1372 4402
rect 1535 4421 1585 4450
rect 1535 4397 1546 4421
rect 1570 4397 1585 4421
rect 1535 4373 1585 4397
rect 1743 4426 1793 4450
rect 1743 4402 1755 4426
rect 1779 4402 1793 4426
rect 1743 4373 1793 4402
rect 1951 4424 2001 4450
rect 2932 4428 2982 4454
rect 3140 4476 3190 4505
rect 3140 4452 3154 4476
rect 3178 4452 3190 4476
rect 3140 4428 3190 4452
rect 3348 4481 3398 4505
rect 3348 4457 3363 4481
rect 3387 4457 3398 4481
rect 3348 4428 3398 4457
rect 3561 4476 3611 4505
rect 3561 4456 3578 4476
rect 3598 4456 3611 4476
rect 3561 4428 3611 4456
rect 1951 4398 1969 4424
rect 1995 4398 2001 4424
rect 1951 4373 2001 4398
rect 1322 4315 1372 4331
rect 1535 4315 1585 4331
rect 1743 4315 1793 4331
rect 1951 4315 2001 4331
rect 7988 4588 8038 4604
rect 8196 4588 8246 4604
rect 8404 4588 8454 4604
rect 8617 4588 8667 4604
rect 10415 4622 10465 4651
rect 10628 4670 10678 4699
rect 10628 4646 10639 4670
rect 10663 4646 10678 4670
rect 10628 4622 10678 4646
rect 10836 4675 10886 4699
rect 10836 4651 10848 4675
rect 10872 4651 10886 4675
rect 10836 4622 10886 4651
rect 11044 4673 11094 4699
rect 11044 4647 11062 4673
rect 11088 4647 11094 4673
rect 11044 4622 11094 4647
rect 18958 4836 19008 4861
rect 18958 4810 18964 4836
rect 18990 4810 19008 4836
rect 18958 4784 19008 4810
rect 19166 4832 19216 4861
rect 19166 4808 19180 4832
rect 19204 4808 19216 4832
rect 19166 4784 19216 4808
rect 19374 4837 19424 4861
rect 19374 4813 19389 4837
rect 19413 4813 19424 4837
rect 19374 4784 19424 4813
rect 19587 4832 19637 4861
rect 19587 4812 19604 4832
rect 19624 4812 19637 4832
rect 19587 4784 19637 4812
rect 15471 4712 15521 4740
rect 15471 4692 15484 4712
rect 15504 4692 15521 4712
rect 13902 4630 13952 4643
rect 14110 4630 14160 4643
rect 14318 4630 14368 4643
rect 14531 4630 14581 4643
rect 15471 4663 15521 4692
rect 15684 4711 15734 4740
rect 15684 4687 15695 4711
rect 15719 4687 15734 4711
rect 15684 4663 15734 4687
rect 15892 4716 15942 4740
rect 15892 4692 15904 4716
rect 15928 4692 15942 4716
rect 15892 4663 15942 4692
rect 16100 4714 16150 4740
rect 16100 4688 16118 4714
rect 16144 4688 16150 4714
rect 16100 4663 16150 4688
rect 18958 4671 19008 4684
rect 19166 4671 19216 4684
rect 19374 4671 19424 4684
rect 19587 4671 19637 4684
rect 15471 4605 15521 4621
rect 15684 4605 15734 4621
rect 15892 4605 15942 4621
rect 16100 4605 16150 4621
rect 10415 4564 10465 4580
rect 10628 4564 10678 4580
rect 10836 4564 10886 4580
rect 11044 4564 11094 4580
rect 16409 4596 16459 4609
rect 16622 4596 16672 4609
rect 16830 4596 16880 4609
rect 17038 4596 17088 4609
rect 7988 4521 8038 4546
rect 7988 4495 7994 4521
rect 8020 4495 8038 4521
rect 6378 4463 6428 4491
rect 6378 4443 6391 4463
rect 6411 4443 6428 4463
rect 6378 4414 6428 4443
rect 6591 4462 6641 4491
rect 6591 4438 6602 4462
rect 6626 4438 6641 4462
rect 6591 4414 6641 4438
rect 6799 4467 6849 4491
rect 6799 4443 6811 4467
rect 6835 4443 6849 4467
rect 6799 4414 6849 4443
rect 7007 4465 7057 4491
rect 7988 4469 8038 4495
rect 8196 4517 8246 4546
rect 8196 4493 8210 4517
rect 8234 4493 8246 4517
rect 8196 4469 8246 4493
rect 8404 4522 8454 4546
rect 8404 4498 8419 4522
rect 8443 4498 8454 4522
rect 8404 4469 8454 4498
rect 8617 4517 8667 4546
rect 11353 4555 11403 4568
rect 11566 4555 11616 4568
rect 11774 4555 11824 4568
rect 11982 4555 12032 4568
rect 8617 4497 8634 4517
rect 8654 4497 8667 4517
rect 8617 4469 8667 4497
rect 7007 4439 7025 4465
rect 7051 4439 7057 4465
rect 7007 4414 7057 4439
rect 6378 4356 6428 4372
rect 6591 4356 6641 4372
rect 6799 4356 6849 4372
rect 7007 4356 7057 4372
rect 12963 4552 13013 4568
rect 13171 4552 13221 4568
rect 13379 4552 13429 4568
rect 13592 4552 13642 4568
rect 12963 4485 13013 4510
rect 12963 4459 12969 4485
rect 12995 4459 13013 4485
rect 11353 4427 11403 4455
rect 11353 4407 11366 4427
rect 11386 4407 11403 4427
rect 7988 4356 8038 4369
rect 8196 4356 8246 4369
rect 8404 4356 8454 4369
rect 8617 4356 8667 4369
rect 11353 4378 11403 4407
rect 11566 4426 11616 4455
rect 11566 4402 11577 4426
rect 11601 4402 11616 4426
rect 11566 4378 11616 4402
rect 11774 4431 11824 4455
rect 11774 4407 11786 4431
rect 11810 4407 11824 4431
rect 11774 4378 11824 4407
rect 11982 4429 12032 4455
rect 12963 4433 13013 4459
rect 13171 4481 13221 4510
rect 13171 4457 13185 4481
rect 13209 4457 13221 4481
rect 13171 4433 13221 4457
rect 13379 4486 13429 4510
rect 13379 4462 13394 4486
rect 13418 4462 13429 4486
rect 13379 4433 13429 4462
rect 13592 4481 13642 4510
rect 13592 4461 13609 4481
rect 13629 4461 13642 4481
rect 13592 4433 13642 4461
rect 11982 4403 12000 4429
rect 12026 4403 12032 4429
rect 11982 4378 12032 4403
rect 2932 4315 2982 4328
rect 3140 4315 3190 4328
rect 3348 4315 3398 4328
rect 3561 4315 3611 4328
rect 8926 4344 8976 4360
rect 9134 4344 9184 4360
rect 9342 4344 9392 4360
rect 9555 4344 9605 4360
rect 3870 4303 3920 4319
rect 4078 4303 4128 4319
rect 4286 4303 4336 4319
rect 4499 4303 4549 4319
rect 383 4240 433 4253
rect 596 4240 646 4253
rect 804 4240 854 4253
rect 1012 4240 1062 4253
rect 3870 4236 3920 4261
rect 3870 4210 3876 4236
rect 3902 4210 3920 4236
rect 3870 4184 3920 4210
rect 4078 4232 4128 4261
rect 4078 4208 4092 4232
rect 4116 4208 4128 4232
rect 4078 4184 4128 4208
rect 4286 4237 4336 4261
rect 4286 4213 4301 4237
rect 4325 4213 4336 4237
rect 4286 4184 4336 4213
rect 4499 4232 4549 4261
rect 5439 4281 5489 4294
rect 5652 4281 5702 4294
rect 5860 4281 5910 4294
rect 6068 4281 6118 4294
rect 4499 4212 4516 4232
rect 4536 4212 4549 4232
rect 4499 4184 4549 4212
rect 383 4112 433 4140
rect 383 4092 396 4112
rect 416 4092 433 4112
rect 383 4063 433 4092
rect 596 4111 646 4140
rect 596 4087 607 4111
rect 631 4087 646 4111
rect 596 4063 646 4087
rect 804 4116 854 4140
rect 804 4092 816 4116
rect 840 4092 854 4116
rect 804 4063 854 4092
rect 1012 4114 1062 4140
rect 1012 4088 1030 4114
rect 1056 4088 1062 4114
rect 1012 4063 1062 4088
rect 8926 4277 8976 4302
rect 8926 4251 8932 4277
rect 8958 4251 8976 4277
rect 8926 4225 8976 4251
rect 9134 4273 9184 4302
rect 9134 4249 9148 4273
rect 9172 4249 9184 4273
rect 9134 4225 9184 4249
rect 9342 4278 9392 4302
rect 9342 4254 9357 4278
rect 9381 4254 9392 4278
rect 9342 4225 9392 4254
rect 9555 4273 9605 4302
rect 11353 4320 11403 4336
rect 11566 4320 11616 4336
rect 11774 4320 11824 4336
rect 11982 4320 12032 4336
rect 18019 4593 18069 4609
rect 18227 4593 18277 4609
rect 18435 4593 18485 4609
rect 18648 4593 18698 4609
rect 18019 4526 18069 4551
rect 18019 4500 18025 4526
rect 18051 4500 18069 4526
rect 16409 4468 16459 4496
rect 16409 4448 16422 4468
rect 16442 4448 16459 4468
rect 16409 4419 16459 4448
rect 16622 4467 16672 4496
rect 16622 4443 16633 4467
rect 16657 4443 16672 4467
rect 16622 4419 16672 4443
rect 16830 4472 16880 4496
rect 16830 4448 16842 4472
rect 16866 4448 16880 4472
rect 16830 4419 16880 4448
rect 17038 4470 17088 4496
rect 18019 4474 18069 4500
rect 18227 4522 18277 4551
rect 18227 4498 18241 4522
rect 18265 4498 18277 4522
rect 18227 4474 18277 4498
rect 18435 4527 18485 4551
rect 18435 4503 18450 4527
rect 18474 4503 18485 4527
rect 18435 4474 18485 4503
rect 18648 4522 18698 4551
rect 18648 4502 18665 4522
rect 18685 4502 18698 4522
rect 18648 4474 18698 4502
rect 17038 4444 17056 4470
rect 17082 4444 17088 4470
rect 17038 4419 17088 4444
rect 16409 4361 16459 4377
rect 16622 4361 16672 4377
rect 16830 4361 16880 4377
rect 17038 4361 17088 4377
rect 18019 4361 18069 4374
rect 18227 4361 18277 4374
rect 18435 4361 18485 4374
rect 18648 4361 18698 4374
rect 12963 4320 13013 4333
rect 13171 4320 13221 4333
rect 13379 4320 13429 4333
rect 13592 4320 13642 4333
rect 18957 4349 19007 4365
rect 19165 4349 19215 4365
rect 19373 4349 19423 4365
rect 19586 4349 19636 4365
rect 9555 4253 9572 4273
rect 9592 4253 9605 4273
rect 13901 4308 13951 4324
rect 14109 4308 14159 4324
rect 14317 4308 14367 4324
rect 14530 4308 14580 4324
rect 9555 4225 9605 4253
rect 5439 4153 5489 4181
rect 5439 4133 5452 4153
rect 5472 4133 5489 4153
rect 5439 4104 5489 4133
rect 5652 4152 5702 4181
rect 5652 4128 5663 4152
rect 5687 4128 5702 4152
rect 5652 4104 5702 4128
rect 5860 4157 5910 4181
rect 5860 4133 5872 4157
rect 5896 4133 5910 4157
rect 5860 4104 5910 4133
rect 6068 4155 6118 4181
rect 6068 4129 6086 4155
rect 6112 4129 6118 4155
rect 6068 4104 6118 4129
rect 10414 4245 10464 4258
rect 10627 4245 10677 4258
rect 10835 4245 10885 4258
rect 11043 4245 11093 4258
rect 13901 4241 13951 4266
rect 13901 4215 13907 4241
rect 13933 4215 13951 4241
rect 13901 4189 13951 4215
rect 14109 4237 14159 4266
rect 14109 4213 14123 4237
rect 14147 4213 14159 4237
rect 14109 4189 14159 4213
rect 14317 4242 14367 4266
rect 14317 4218 14332 4242
rect 14356 4218 14367 4242
rect 14317 4189 14367 4218
rect 14530 4237 14580 4266
rect 15470 4286 15520 4299
rect 15683 4286 15733 4299
rect 15891 4286 15941 4299
rect 16099 4286 16149 4299
rect 14530 4217 14547 4237
rect 14567 4217 14580 4237
rect 14530 4189 14580 4217
rect 8926 4112 8976 4125
rect 9134 4112 9184 4125
rect 9342 4112 9392 4125
rect 9555 4112 9605 4125
rect 10414 4117 10464 4145
rect 3870 4071 3920 4084
rect 4078 4071 4128 4084
rect 4286 4071 4336 4084
rect 4499 4071 4549 4084
rect 2792 4036 2842 4052
rect 3000 4036 3050 4052
rect 3208 4036 3258 4052
rect 3421 4036 3471 4052
rect 383 4005 433 4021
rect 596 4005 646 4021
rect 804 4005 854 4021
rect 1012 4005 1062 4021
rect 7848 4077 7898 4093
rect 8056 4077 8106 4093
rect 8264 4077 8314 4093
rect 8477 4077 8527 4093
rect 5439 4046 5489 4062
rect 5652 4046 5702 4062
rect 5860 4046 5910 4062
rect 6068 4046 6118 4062
rect 10414 4097 10427 4117
rect 10447 4097 10464 4117
rect 10414 4068 10464 4097
rect 10627 4116 10677 4145
rect 10627 4092 10638 4116
rect 10662 4092 10677 4116
rect 10627 4068 10677 4092
rect 10835 4121 10885 4145
rect 10835 4097 10847 4121
rect 10871 4097 10885 4121
rect 10835 4068 10885 4097
rect 11043 4119 11093 4145
rect 11043 4093 11061 4119
rect 11087 4093 11093 4119
rect 11043 4068 11093 4093
rect 18957 4282 19007 4307
rect 18957 4256 18963 4282
rect 18989 4256 19007 4282
rect 18957 4230 19007 4256
rect 19165 4278 19215 4307
rect 19165 4254 19179 4278
rect 19203 4254 19215 4278
rect 19165 4230 19215 4254
rect 19373 4283 19423 4307
rect 19373 4259 19388 4283
rect 19412 4259 19423 4283
rect 19373 4230 19423 4259
rect 19586 4278 19636 4307
rect 19586 4258 19603 4278
rect 19623 4258 19636 4278
rect 19586 4230 19636 4258
rect 15470 4158 15520 4186
rect 15470 4138 15483 4158
rect 15503 4138 15520 4158
rect 15470 4109 15520 4138
rect 15683 4157 15733 4186
rect 15683 4133 15694 4157
rect 15718 4133 15733 4157
rect 15683 4109 15733 4133
rect 15891 4162 15941 4186
rect 15891 4138 15903 4162
rect 15927 4138 15941 4162
rect 15891 4109 15941 4138
rect 16099 4160 16149 4186
rect 16099 4134 16117 4160
rect 16143 4134 16149 4160
rect 16099 4109 16149 4134
rect 18957 4117 19007 4130
rect 19165 4117 19215 4130
rect 19373 4117 19423 4130
rect 19586 4117 19636 4130
rect 13901 4076 13951 4089
rect 14109 4076 14159 4089
rect 14317 4076 14367 4089
rect 14530 4076 14580 4089
rect 1463 3958 1513 3971
rect 1676 3958 1726 3971
rect 1884 3958 1934 3971
rect 2092 3958 2142 3971
rect 2792 3969 2842 3994
rect 2792 3943 2798 3969
rect 2824 3943 2842 3969
rect 2792 3917 2842 3943
rect 3000 3965 3050 3994
rect 3000 3941 3014 3965
rect 3038 3941 3050 3965
rect 3000 3917 3050 3941
rect 3208 3970 3258 3994
rect 3208 3946 3223 3970
rect 3247 3946 3258 3970
rect 3208 3917 3258 3946
rect 3421 3965 3471 3994
rect 6519 3999 6569 4012
rect 6732 3999 6782 4012
rect 6940 3999 6990 4012
rect 7148 3999 7198 4012
rect 7848 4010 7898 4035
rect 3421 3945 3438 3965
rect 3458 3945 3471 3965
rect 3421 3917 3471 3945
rect 1463 3830 1513 3858
rect 1463 3810 1476 3830
rect 1496 3810 1513 3830
rect 1463 3781 1513 3810
rect 1676 3829 1726 3858
rect 1676 3805 1687 3829
rect 1711 3805 1726 3829
rect 1676 3781 1726 3805
rect 1884 3834 1934 3858
rect 1884 3810 1896 3834
rect 1920 3810 1934 3834
rect 1884 3781 1934 3810
rect 2092 3832 2142 3858
rect 2092 3806 2110 3832
rect 2136 3806 2142 3832
rect 7848 3984 7854 4010
rect 7880 3984 7898 4010
rect 7848 3958 7898 3984
rect 8056 4006 8106 4035
rect 8056 3982 8070 4006
rect 8094 3982 8106 4006
rect 8056 3958 8106 3982
rect 8264 4011 8314 4035
rect 8264 3987 8279 4011
rect 8303 3987 8314 4011
rect 8264 3958 8314 3987
rect 8477 4006 8527 4035
rect 12823 4041 12873 4057
rect 13031 4041 13081 4057
rect 13239 4041 13289 4057
rect 13452 4041 13502 4057
rect 10414 4010 10464 4026
rect 10627 4010 10677 4026
rect 10835 4010 10885 4026
rect 11043 4010 11093 4026
rect 8477 3986 8494 4006
rect 8514 3986 8527 4006
rect 17879 4082 17929 4098
rect 18087 4082 18137 4098
rect 18295 4082 18345 4098
rect 18508 4082 18558 4098
rect 15470 4051 15520 4067
rect 15683 4051 15733 4067
rect 15891 4051 15941 4067
rect 16099 4051 16149 4067
rect 8477 3958 8527 3986
rect 6519 3871 6569 3899
rect 6519 3851 6532 3871
rect 6552 3851 6569 3871
rect 2092 3781 2142 3806
rect 2792 3804 2842 3817
rect 3000 3804 3050 3817
rect 3208 3804 3258 3817
rect 3421 3804 3471 3817
rect 6519 3822 6569 3851
rect 6732 3870 6782 3899
rect 6732 3846 6743 3870
rect 6767 3846 6782 3870
rect 6732 3822 6782 3846
rect 6940 3875 6990 3899
rect 6940 3851 6952 3875
rect 6976 3851 6990 3875
rect 6940 3822 6990 3851
rect 7148 3873 7198 3899
rect 7148 3847 7166 3873
rect 7192 3847 7198 3873
rect 11494 3963 11544 3976
rect 11707 3963 11757 3976
rect 11915 3963 11965 3976
rect 12123 3963 12173 3976
rect 12823 3974 12873 3999
rect 7148 3822 7198 3847
rect 7848 3845 7898 3858
rect 8056 3845 8106 3858
rect 8264 3845 8314 3858
rect 8477 3845 8527 3858
rect 12823 3948 12829 3974
rect 12855 3948 12873 3974
rect 12823 3922 12873 3948
rect 13031 3970 13081 3999
rect 13031 3946 13045 3970
rect 13069 3946 13081 3970
rect 13031 3922 13081 3946
rect 13239 3975 13289 3999
rect 13239 3951 13254 3975
rect 13278 3951 13289 3975
rect 13239 3922 13289 3951
rect 13452 3970 13502 3999
rect 16550 4004 16600 4017
rect 16763 4004 16813 4017
rect 16971 4004 17021 4017
rect 17179 4004 17229 4017
rect 17879 4015 17929 4040
rect 13452 3950 13469 3970
rect 13489 3950 13502 3970
rect 13452 3922 13502 3950
rect 11494 3835 11544 3863
rect 3872 3754 3922 3770
rect 4080 3754 4130 3770
rect 4288 3754 4338 3770
rect 4501 3754 4551 3770
rect 1463 3723 1513 3739
rect 1676 3723 1726 3739
rect 1884 3723 1934 3739
rect 2092 3723 2142 3739
rect 11494 3815 11507 3835
rect 11527 3815 11544 3835
rect 8928 3795 8978 3811
rect 9136 3795 9186 3811
rect 9344 3795 9394 3811
rect 9557 3795 9607 3811
rect 6519 3764 6569 3780
rect 6732 3764 6782 3780
rect 6940 3764 6990 3780
rect 7148 3764 7198 3780
rect 11494 3786 11544 3815
rect 11707 3834 11757 3863
rect 11707 3810 11718 3834
rect 11742 3810 11757 3834
rect 11707 3786 11757 3810
rect 11915 3839 11965 3863
rect 11915 3815 11927 3839
rect 11951 3815 11965 3839
rect 11915 3786 11965 3815
rect 12123 3837 12173 3863
rect 12123 3811 12141 3837
rect 12167 3811 12173 3837
rect 17879 3989 17885 4015
rect 17911 3989 17929 4015
rect 17879 3963 17929 3989
rect 18087 4011 18137 4040
rect 18087 3987 18101 4011
rect 18125 3987 18137 4011
rect 18087 3963 18137 3987
rect 18295 4016 18345 4040
rect 18295 3992 18310 4016
rect 18334 3992 18345 4016
rect 18295 3963 18345 3992
rect 18508 4011 18558 4040
rect 18508 3991 18525 4011
rect 18545 3991 18558 4011
rect 18508 3963 18558 3991
rect 16550 3876 16600 3904
rect 16550 3856 16563 3876
rect 16583 3856 16600 3876
rect 12123 3786 12173 3811
rect 12823 3809 12873 3822
rect 13031 3809 13081 3822
rect 13239 3809 13289 3822
rect 13452 3809 13502 3822
rect 16550 3827 16600 3856
rect 16763 3875 16813 3904
rect 16763 3851 16774 3875
rect 16798 3851 16813 3875
rect 16763 3827 16813 3851
rect 16971 3880 17021 3904
rect 16971 3856 16983 3880
rect 17007 3856 17021 3880
rect 16971 3827 17021 3856
rect 17179 3878 17229 3904
rect 17179 3852 17197 3878
rect 17223 3852 17229 3878
rect 17179 3827 17229 3852
rect 17879 3850 17929 3863
rect 18087 3850 18137 3863
rect 18295 3850 18345 3863
rect 18508 3850 18558 3863
rect 5441 3732 5491 3745
rect 5654 3732 5704 3745
rect 5862 3732 5912 3745
rect 6070 3732 6120 3745
rect 385 3691 435 3704
rect 598 3691 648 3704
rect 806 3691 856 3704
rect 1014 3691 1064 3704
rect 3872 3687 3922 3712
rect 3872 3661 3878 3687
rect 3904 3661 3922 3687
rect 3872 3635 3922 3661
rect 4080 3683 4130 3712
rect 4080 3659 4094 3683
rect 4118 3659 4130 3683
rect 4080 3635 4130 3659
rect 4288 3688 4338 3712
rect 4288 3664 4303 3688
rect 4327 3664 4338 3688
rect 4288 3635 4338 3664
rect 4501 3683 4551 3712
rect 4501 3663 4518 3683
rect 4538 3663 4551 3683
rect 4501 3635 4551 3663
rect 385 3563 435 3591
rect 385 3543 398 3563
rect 418 3543 435 3563
rect 385 3514 435 3543
rect 598 3562 648 3591
rect 598 3538 609 3562
rect 633 3538 648 3562
rect 598 3514 648 3538
rect 806 3567 856 3591
rect 806 3543 818 3567
rect 842 3543 856 3567
rect 806 3514 856 3543
rect 1014 3565 1064 3591
rect 1014 3539 1032 3565
rect 1058 3539 1064 3565
rect 1014 3514 1064 3539
rect 8928 3728 8978 3753
rect 8928 3702 8934 3728
rect 8960 3702 8978 3728
rect 8928 3676 8978 3702
rect 9136 3724 9186 3753
rect 9136 3700 9150 3724
rect 9174 3700 9186 3724
rect 9136 3676 9186 3700
rect 9344 3729 9394 3753
rect 9344 3705 9359 3729
rect 9383 3705 9394 3729
rect 9344 3676 9394 3705
rect 9557 3724 9607 3753
rect 9557 3704 9574 3724
rect 9594 3704 9607 3724
rect 13903 3759 13953 3775
rect 14111 3759 14161 3775
rect 14319 3759 14369 3775
rect 14532 3759 14582 3775
rect 11494 3728 11544 3744
rect 11707 3728 11757 3744
rect 11915 3728 11965 3744
rect 12123 3728 12173 3744
rect 18959 3800 19009 3816
rect 19167 3800 19217 3816
rect 19375 3800 19425 3816
rect 19588 3800 19638 3816
rect 16550 3769 16600 3785
rect 16763 3769 16813 3785
rect 16971 3769 17021 3785
rect 17179 3769 17229 3785
rect 15472 3737 15522 3750
rect 15685 3737 15735 3750
rect 15893 3737 15943 3750
rect 16101 3737 16151 3750
rect 9557 3676 9607 3704
rect 10416 3696 10466 3709
rect 10629 3696 10679 3709
rect 10837 3696 10887 3709
rect 11045 3696 11095 3709
rect 5441 3604 5491 3632
rect 5441 3584 5454 3604
rect 5474 3584 5491 3604
rect 3872 3522 3922 3535
rect 4080 3522 4130 3535
rect 4288 3522 4338 3535
rect 4501 3522 4551 3535
rect 5441 3555 5491 3584
rect 5654 3603 5704 3632
rect 5654 3579 5665 3603
rect 5689 3579 5704 3603
rect 5654 3555 5704 3579
rect 5862 3608 5912 3632
rect 5862 3584 5874 3608
rect 5898 3584 5912 3608
rect 5862 3555 5912 3584
rect 6070 3606 6120 3632
rect 6070 3580 6088 3606
rect 6114 3580 6120 3606
rect 6070 3555 6120 3580
rect 8928 3563 8978 3576
rect 9136 3563 9186 3576
rect 9344 3563 9394 3576
rect 9557 3563 9607 3576
rect 13903 3692 13953 3717
rect 13903 3666 13909 3692
rect 13935 3666 13953 3692
rect 13903 3640 13953 3666
rect 14111 3688 14161 3717
rect 14111 3664 14125 3688
rect 14149 3664 14161 3688
rect 14111 3640 14161 3664
rect 14319 3693 14369 3717
rect 14319 3669 14334 3693
rect 14358 3669 14369 3693
rect 14319 3640 14369 3669
rect 14532 3688 14582 3717
rect 14532 3668 14549 3688
rect 14569 3668 14582 3688
rect 14532 3640 14582 3668
rect 10416 3568 10466 3596
rect 5441 3497 5491 3513
rect 5654 3497 5704 3513
rect 5862 3497 5912 3513
rect 6070 3497 6120 3513
rect 10416 3548 10429 3568
rect 10449 3548 10466 3568
rect 385 3456 435 3472
rect 598 3456 648 3472
rect 806 3456 856 3472
rect 1014 3456 1064 3472
rect 6379 3488 6429 3501
rect 6592 3488 6642 3501
rect 6800 3488 6850 3501
rect 7008 3488 7058 3501
rect 1323 3447 1373 3460
rect 1536 3447 1586 3460
rect 1744 3447 1794 3460
rect 1952 3447 2002 3460
rect 2933 3444 2983 3460
rect 3141 3444 3191 3460
rect 3349 3444 3399 3460
rect 3562 3444 3612 3460
rect 2933 3377 2983 3402
rect 2933 3351 2939 3377
rect 2965 3351 2983 3377
rect 1323 3319 1373 3347
rect 1323 3299 1336 3319
rect 1356 3299 1373 3319
rect 1323 3270 1373 3299
rect 1536 3318 1586 3347
rect 1536 3294 1547 3318
rect 1571 3294 1586 3318
rect 1536 3270 1586 3294
rect 1744 3323 1794 3347
rect 1744 3299 1756 3323
rect 1780 3299 1794 3323
rect 1744 3270 1794 3299
rect 1952 3321 2002 3347
rect 2933 3325 2983 3351
rect 3141 3373 3191 3402
rect 3141 3349 3155 3373
rect 3179 3349 3191 3373
rect 3141 3325 3191 3349
rect 3349 3378 3399 3402
rect 3349 3354 3364 3378
rect 3388 3354 3399 3378
rect 3349 3325 3399 3354
rect 3562 3373 3612 3402
rect 3562 3353 3579 3373
rect 3599 3353 3612 3373
rect 3562 3325 3612 3353
rect 1952 3295 1970 3321
rect 1996 3295 2002 3321
rect 1952 3270 2002 3295
rect 1323 3212 1373 3228
rect 1536 3212 1586 3228
rect 1744 3212 1794 3228
rect 1952 3212 2002 3228
rect 7989 3485 8039 3501
rect 8197 3485 8247 3501
rect 8405 3485 8455 3501
rect 8618 3485 8668 3501
rect 10416 3519 10466 3548
rect 10629 3567 10679 3596
rect 10629 3543 10640 3567
rect 10664 3543 10679 3567
rect 10629 3519 10679 3543
rect 10837 3572 10887 3596
rect 10837 3548 10849 3572
rect 10873 3548 10887 3572
rect 10837 3519 10887 3548
rect 11045 3570 11095 3596
rect 11045 3544 11063 3570
rect 11089 3544 11095 3570
rect 11045 3519 11095 3544
rect 18959 3733 19009 3758
rect 18959 3707 18965 3733
rect 18991 3707 19009 3733
rect 18959 3681 19009 3707
rect 19167 3729 19217 3758
rect 19167 3705 19181 3729
rect 19205 3705 19217 3729
rect 19167 3681 19217 3705
rect 19375 3734 19425 3758
rect 19375 3710 19390 3734
rect 19414 3710 19425 3734
rect 19375 3681 19425 3710
rect 19588 3729 19638 3758
rect 19588 3709 19605 3729
rect 19625 3709 19638 3729
rect 19588 3681 19638 3709
rect 15472 3609 15522 3637
rect 15472 3589 15485 3609
rect 15505 3589 15522 3609
rect 13903 3527 13953 3540
rect 14111 3527 14161 3540
rect 14319 3527 14369 3540
rect 14532 3527 14582 3540
rect 15472 3560 15522 3589
rect 15685 3608 15735 3637
rect 15685 3584 15696 3608
rect 15720 3584 15735 3608
rect 15685 3560 15735 3584
rect 15893 3613 15943 3637
rect 15893 3589 15905 3613
rect 15929 3589 15943 3613
rect 15893 3560 15943 3589
rect 16101 3611 16151 3637
rect 16101 3585 16119 3611
rect 16145 3585 16151 3611
rect 16101 3560 16151 3585
rect 18959 3568 19009 3581
rect 19167 3568 19217 3581
rect 19375 3568 19425 3581
rect 19588 3568 19638 3581
rect 15472 3502 15522 3518
rect 15685 3502 15735 3518
rect 15893 3502 15943 3518
rect 16101 3502 16151 3518
rect 10416 3461 10466 3477
rect 10629 3461 10679 3477
rect 10837 3461 10887 3477
rect 11045 3461 11095 3477
rect 16410 3493 16460 3506
rect 16623 3493 16673 3506
rect 16831 3493 16881 3506
rect 17039 3493 17089 3506
rect 7989 3418 8039 3443
rect 7989 3392 7995 3418
rect 8021 3392 8039 3418
rect 6379 3360 6429 3388
rect 6379 3340 6392 3360
rect 6412 3340 6429 3360
rect 6379 3311 6429 3340
rect 6592 3359 6642 3388
rect 6592 3335 6603 3359
rect 6627 3335 6642 3359
rect 6592 3311 6642 3335
rect 6800 3364 6850 3388
rect 6800 3340 6812 3364
rect 6836 3340 6850 3364
rect 6800 3311 6850 3340
rect 7008 3362 7058 3388
rect 7989 3366 8039 3392
rect 8197 3414 8247 3443
rect 8197 3390 8211 3414
rect 8235 3390 8247 3414
rect 8197 3366 8247 3390
rect 8405 3419 8455 3443
rect 8405 3395 8420 3419
rect 8444 3395 8455 3419
rect 8405 3366 8455 3395
rect 8618 3414 8668 3443
rect 11354 3452 11404 3465
rect 11567 3452 11617 3465
rect 11775 3452 11825 3465
rect 11983 3452 12033 3465
rect 8618 3394 8635 3414
rect 8655 3394 8668 3414
rect 8618 3366 8668 3394
rect 7008 3336 7026 3362
rect 7052 3336 7058 3362
rect 7008 3311 7058 3336
rect 6379 3253 6429 3269
rect 6592 3253 6642 3269
rect 6800 3253 6850 3269
rect 7008 3253 7058 3269
rect 12964 3449 13014 3465
rect 13172 3449 13222 3465
rect 13380 3449 13430 3465
rect 13593 3449 13643 3465
rect 12964 3382 13014 3407
rect 12964 3356 12970 3382
rect 12996 3356 13014 3382
rect 11354 3324 11404 3352
rect 11354 3304 11367 3324
rect 11387 3304 11404 3324
rect 7989 3253 8039 3266
rect 8197 3253 8247 3266
rect 8405 3253 8455 3266
rect 8618 3253 8668 3266
rect 11354 3275 11404 3304
rect 11567 3323 11617 3352
rect 11567 3299 11578 3323
rect 11602 3299 11617 3323
rect 11567 3275 11617 3299
rect 11775 3328 11825 3352
rect 11775 3304 11787 3328
rect 11811 3304 11825 3328
rect 11775 3275 11825 3304
rect 11983 3326 12033 3352
rect 12964 3330 13014 3356
rect 13172 3378 13222 3407
rect 13172 3354 13186 3378
rect 13210 3354 13222 3378
rect 13172 3330 13222 3354
rect 13380 3383 13430 3407
rect 13380 3359 13395 3383
rect 13419 3359 13430 3383
rect 13380 3330 13430 3359
rect 13593 3378 13643 3407
rect 13593 3358 13610 3378
rect 13630 3358 13643 3378
rect 13593 3330 13643 3358
rect 11983 3300 12001 3326
rect 12027 3300 12033 3326
rect 11983 3275 12033 3300
rect 2933 3212 2983 3225
rect 3141 3212 3191 3225
rect 3349 3212 3399 3225
rect 3562 3212 3612 3225
rect 8927 3241 8977 3257
rect 9135 3241 9185 3257
rect 9343 3241 9393 3257
rect 9556 3241 9606 3257
rect 3871 3200 3921 3216
rect 4079 3200 4129 3216
rect 4287 3200 4337 3216
rect 4500 3200 4550 3216
rect 384 3137 434 3150
rect 597 3137 647 3150
rect 805 3137 855 3150
rect 1013 3137 1063 3150
rect 3871 3133 3921 3158
rect 3871 3107 3877 3133
rect 3903 3107 3921 3133
rect 3871 3081 3921 3107
rect 4079 3129 4129 3158
rect 4079 3105 4093 3129
rect 4117 3105 4129 3129
rect 4079 3081 4129 3105
rect 4287 3134 4337 3158
rect 4287 3110 4302 3134
rect 4326 3110 4337 3134
rect 4287 3081 4337 3110
rect 4500 3129 4550 3158
rect 5440 3178 5490 3191
rect 5653 3178 5703 3191
rect 5861 3178 5911 3191
rect 6069 3178 6119 3191
rect 4500 3109 4517 3129
rect 4537 3109 4550 3129
rect 4500 3081 4550 3109
rect 384 3009 434 3037
rect 384 2989 397 3009
rect 417 2989 434 3009
rect 384 2960 434 2989
rect 597 3008 647 3037
rect 597 2984 608 3008
rect 632 2984 647 3008
rect 597 2960 647 2984
rect 805 3013 855 3037
rect 805 2989 817 3013
rect 841 2989 855 3013
rect 805 2960 855 2989
rect 1013 3011 1063 3037
rect 1013 2985 1031 3011
rect 1057 2985 1063 3011
rect 1013 2960 1063 2985
rect 8927 3174 8977 3199
rect 8927 3148 8933 3174
rect 8959 3148 8977 3174
rect 8927 3122 8977 3148
rect 9135 3170 9185 3199
rect 9135 3146 9149 3170
rect 9173 3146 9185 3170
rect 9135 3122 9185 3146
rect 9343 3175 9393 3199
rect 9343 3151 9358 3175
rect 9382 3151 9393 3175
rect 9343 3122 9393 3151
rect 9556 3170 9606 3199
rect 11354 3217 11404 3233
rect 11567 3217 11617 3233
rect 11775 3217 11825 3233
rect 11983 3217 12033 3233
rect 18020 3490 18070 3506
rect 18228 3490 18278 3506
rect 18436 3490 18486 3506
rect 18649 3490 18699 3506
rect 18020 3423 18070 3448
rect 18020 3397 18026 3423
rect 18052 3397 18070 3423
rect 16410 3365 16460 3393
rect 16410 3345 16423 3365
rect 16443 3345 16460 3365
rect 16410 3316 16460 3345
rect 16623 3364 16673 3393
rect 16623 3340 16634 3364
rect 16658 3340 16673 3364
rect 16623 3316 16673 3340
rect 16831 3369 16881 3393
rect 16831 3345 16843 3369
rect 16867 3345 16881 3369
rect 16831 3316 16881 3345
rect 17039 3367 17089 3393
rect 18020 3371 18070 3397
rect 18228 3419 18278 3448
rect 18228 3395 18242 3419
rect 18266 3395 18278 3419
rect 18228 3371 18278 3395
rect 18436 3424 18486 3448
rect 18436 3400 18451 3424
rect 18475 3400 18486 3424
rect 18436 3371 18486 3400
rect 18649 3419 18699 3448
rect 18649 3399 18666 3419
rect 18686 3399 18699 3419
rect 18649 3371 18699 3399
rect 17039 3341 17057 3367
rect 17083 3341 17089 3367
rect 17039 3316 17089 3341
rect 16410 3258 16460 3274
rect 16623 3258 16673 3274
rect 16831 3258 16881 3274
rect 17039 3258 17089 3274
rect 18020 3258 18070 3271
rect 18228 3258 18278 3271
rect 18436 3258 18486 3271
rect 18649 3258 18699 3271
rect 12964 3217 13014 3230
rect 13172 3217 13222 3230
rect 13380 3217 13430 3230
rect 13593 3217 13643 3230
rect 18958 3246 19008 3262
rect 19166 3246 19216 3262
rect 19374 3246 19424 3262
rect 19587 3246 19637 3262
rect 9556 3150 9573 3170
rect 9593 3150 9606 3170
rect 13902 3205 13952 3221
rect 14110 3205 14160 3221
rect 14318 3205 14368 3221
rect 14531 3205 14581 3221
rect 9556 3122 9606 3150
rect 5440 3050 5490 3078
rect 5440 3030 5453 3050
rect 5473 3030 5490 3050
rect 5440 3001 5490 3030
rect 5653 3049 5703 3078
rect 5653 3025 5664 3049
rect 5688 3025 5703 3049
rect 5653 3001 5703 3025
rect 5861 3054 5911 3078
rect 5861 3030 5873 3054
rect 5897 3030 5911 3054
rect 5861 3001 5911 3030
rect 6069 3052 6119 3078
rect 6069 3026 6087 3052
rect 6113 3026 6119 3052
rect 6069 3001 6119 3026
rect 10415 3142 10465 3155
rect 10628 3142 10678 3155
rect 10836 3142 10886 3155
rect 11044 3142 11094 3155
rect 13902 3138 13952 3163
rect 13902 3112 13908 3138
rect 13934 3112 13952 3138
rect 13902 3086 13952 3112
rect 14110 3134 14160 3163
rect 14110 3110 14124 3134
rect 14148 3110 14160 3134
rect 14110 3086 14160 3110
rect 14318 3139 14368 3163
rect 14318 3115 14333 3139
rect 14357 3115 14368 3139
rect 14318 3086 14368 3115
rect 14531 3134 14581 3163
rect 15471 3183 15521 3196
rect 15684 3183 15734 3196
rect 15892 3183 15942 3196
rect 16100 3183 16150 3196
rect 14531 3114 14548 3134
rect 14568 3114 14581 3134
rect 14531 3086 14581 3114
rect 8927 3009 8977 3022
rect 9135 3009 9185 3022
rect 9343 3009 9393 3022
rect 9556 3009 9606 3022
rect 10415 3014 10465 3042
rect 3871 2968 3921 2981
rect 4079 2968 4129 2981
rect 4287 2968 4337 2981
rect 4500 2968 4550 2981
rect 384 2902 434 2918
rect 597 2902 647 2918
rect 805 2902 855 2918
rect 1013 2902 1063 2918
rect 2823 2920 2873 2936
rect 3031 2920 3081 2936
rect 3239 2920 3289 2936
rect 3452 2920 3502 2936
rect 1433 2868 1483 2881
rect 1646 2868 1696 2881
rect 1854 2868 1904 2881
rect 2062 2868 2112 2881
rect 5440 2943 5490 2959
rect 5653 2943 5703 2959
rect 5861 2943 5911 2959
rect 6069 2943 6119 2959
rect 7879 2961 7929 2977
rect 8087 2961 8137 2977
rect 8295 2961 8345 2977
rect 8508 2961 8558 2977
rect 6489 2909 6539 2922
rect 6702 2909 6752 2922
rect 6910 2909 6960 2922
rect 7118 2909 7168 2922
rect 10415 2994 10428 3014
rect 10448 2994 10465 3014
rect 10415 2965 10465 2994
rect 10628 3013 10678 3042
rect 10628 2989 10639 3013
rect 10663 2989 10678 3013
rect 10628 2965 10678 2989
rect 10836 3018 10886 3042
rect 10836 2994 10848 3018
rect 10872 2994 10886 3018
rect 10836 2965 10886 2994
rect 11044 3016 11094 3042
rect 11044 2990 11062 3016
rect 11088 2990 11094 3016
rect 11044 2965 11094 2990
rect 18958 3179 19008 3204
rect 18958 3153 18964 3179
rect 18990 3153 19008 3179
rect 18958 3127 19008 3153
rect 19166 3175 19216 3204
rect 19166 3151 19180 3175
rect 19204 3151 19216 3175
rect 19166 3127 19216 3151
rect 19374 3180 19424 3204
rect 19374 3156 19389 3180
rect 19413 3156 19424 3180
rect 19374 3127 19424 3156
rect 19587 3175 19637 3204
rect 19587 3155 19604 3175
rect 19624 3155 19637 3175
rect 19587 3127 19637 3155
rect 15471 3055 15521 3083
rect 15471 3035 15484 3055
rect 15504 3035 15521 3055
rect 15471 3006 15521 3035
rect 15684 3054 15734 3083
rect 15684 3030 15695 3054
rect 15719 3030 15734 3054
rect 15684 3006 15734 3030
rect 15892 3059 15942 3083
rect 15892 3035 15904 3059
rect 15928 3035 15942 3059
rect 15892 3006 15942 3035
rect 16100 3057 16150 3083
rect 16100 3031 16118 3057
rect 16144 3031 16150 3057
rect 16100 3006 16150 3031
rect 18958 3014 19008 3027
rect 19166 3014 19216 3027
rect 19374 3014 19424 3027
rect 19587 3014 19637 3027
rect 13902 2973 13952 2986
rect 14110 2973 14160 2986
rect 14318 2973 14368 2986
rect 14531 2973 14581 2986
rect 2823 2853 2873 2878
rect 2823 2827 2829 2853
rect 2855 2827 2873 2853
rect 2823 2801 2873 2827
rect 3031 2849 3081 2878
rect 3031 2825 3045 2849
rect 3069 2825 3081 2849
rect 3031 2801 3081 2825
rect 3239 2854 3289 2878
rect 3239 2830 3254 2854
rect 3278 2830 3289 2854
rect 3239 2801 3289 2830
rect 3452 2849 3502 2878
rect 3452 2829 3469 2849
rect 3489 2829 3502 2849
rect 3452 2801 3502 2829
rect 7879 2894 7929 2919
rect 7879 2868 7885 2894
rect 7911 2868 7929 2894
rect 7879 2842 7929 2868
rect 8087 2890 8137 2919
rect 8087 2866 8101 2890
rect 8125 2866 8137 2890
rect 8087 2842 8137 2866
rect 8295 2895 8345 2919
rect 8295 2871 8310 2895
rect 8334 2871 8345 2895
rect 8295 2842 8345 2871
rect 8508 2890 8558 2919
rect 10415 2907 10465 2923
rect 10628 2907 10678 2923
rect 10836 2907 10886 2923
rect 11044 2907 11094 2923
rect 12854 2925 12904 2941
rect 13062 2925 13112 2941
rect 13270 2925 13320 2941
rect 13483 2925 13533 2941
rect 8508 2870 8525 2890
rect 8545 2870 8558 2890
rect 8508 2842 8558 2870
rect 11464 2873 11514 2886
rect 11677 2873 11727 2886
rect 11885 2873 11935 2886
rect 12093 2873 12143 2886
rect 15471 2948 15521 2964
rect 15684 2948 15734 2964
rect 15892 2948 15942 2964
rect 16100 2948 16150 2964
rect 17910 2966 17960 2982
rect 18118 2966 18168 2982
rect 18326 2966 18376 2982
rect 18539 2966 18589 2982
rect 16520 2914 16570 2927
rect 16733 2914 16783 2927
rect 16941 2914 16991 2927
rect 17149 2914 17199 2927
rect 1433 2740 1483 2768
rect 1433 2720 1446 2740
rect 1466 2720 1483 2740
rect 1433 2691 1483 2720
rect 1646 2739 1696 2768
rect 1646 2715 1657 2739
rect 1681 2715 1696 2739
rect 1646 2691 1696 2715
rect 1854 2744 1904 2768
rect 1854 2720 1866 2744
rect 1890 2720 1904 2744
rect 1854 2691 1904 2720
rect 2062 2742 2112 2768
rect 2062 2716 2080 2742
rect 2106 2716 2112 2742
rect 2062 2691 2112 2716
rect 6489 2781 6539 2809
rect 6489 2761 6502 2781
rect 6522 2761 6539 2781
rect 6489 2732 6539 2761
rect 6702 2780 6752 2809
rect 6702 2756 6713 2780
rect 6737 2756 6752 2780
rect 6702 2732 6752 2756
rect 6910 2785 6960 2809
rect 6910 2761 6922 2785
rect 6946 2761 6960 2785
rect 6910 2732 6960 2761
rect 7118 2783 7168 2809
rect 7118 2757 7136 2783
rect 7162 2757 7168 2783
rect 7118 2732 7168 2757
rect 12854 2858 12904 2883
rect 12854 2832 12860 2858
rect 12886 2832 12904 2858
rect 12854 2806 12904 2832
rect 13062 2854 13112 2883
rect 13062 2830 13076 2854
rect 13100 2830 13112 2854
rect 13062 2806 13112 2830
rect 13270 2859 13320 2883
rect 13270 2835 13285 2859
rect 13309 2835 13320 2859
rect 13270 2806 13320 2835
rect 13483 2854 13533 2883
rect 13483 2834 13500 2854
rect 13520 2834 13533 2854
rect 13483 2806 13533 2834
rect 17910 2899 17960 2924
rect 17910 2873 17916 2899
rect 17942 2873 17960 2899
rect 17910 2847 17960 2873
rect 18118 2895 18168 2924
rect 18118 2871 18132 2895
rect 18156 2871 18168 2895
rect 18118 2847 18168 2871
rect 18326 2900 18376 2924
rect 18326 2876 18341 2900
rect 18365 2876 18376 2900
rect 18326 2847 18376 2876
rect 18539 2895 18589 2924
rect 18539 2875 18556 2895
rect 18576 2875 18589 2895
rect 18539 2847 18589 2875
rect 2823 2688 2873 2701
rect 3031 2688 3081 2701
rect 3239 2688 3289 2701
rect 3452 2688 3502 2701
rect 1433 2633 1483 2649
rect 1646 2633 1696 2649
rect 1854 2633 1904 2649
rect 2062 2633 2112 2649
rect 3872 2651 3922 2667
rect 4080 2651 4130 2667
rect 4288 2651 4338 2667
rect 4501 2651 4551 2667
rect 7879 2729 7929 2742
rect 8087 2729 8137 2742
rect 8295 2729 8345 2742
rect 8508 2729 8558 2742
rect 11464 2745 11514 2773
rect 11464 2725 11477 2745
rect 11497 2725 11514 2745
rect 6489 2674 6539 2690
rect 6702 2674 6752 2690
rect 6910 2674 6960 2690
rect 7118 2674 7168 2690
rect 8928 2692 8978 2708
rect 9136 2692 9186 2708
rect 9344 2692 9394 2708
rect 9557 2692 9607 2708
rect 11464 2696 11514 2725
rect 11677 2744 11727 2773
rect 11677 2720 11688 2744
rect 11712 2720 11727 2744
rect 11677 2696 11727 2720
rect 11885 2749 11935 2773
rect 11885 2725 11897 2749
rect 11921 2725 11935 2749
rect 11885 2696 11935 2725
rect 12093 2747 12143 2773
rect 12093 2721 12111 2747
rect 12137 2721 12143 2747
rect 12093 2696 12143 2721
rect 16520 2786 16570 2814
rect 16520 2766 16533 2786
rect 16553 2766 16570 2786
rect 16520 2737 16570 2766
rect 16733 2785 16783 2814
rect 16733 2761 16744 2785
rect 16768 2761 16783 2785
rect 16733 2737 16783 2761
rect 16941 2790 16991 2814
rect 16941 2766 16953 2790
rect 16977 2766 16991 2790
rect 16941 2737 16991 2766
rect 17149 2788 17199 2814
rect 17149 2762 17167 2788
rect 17193 2762 17199 2788
rect 17149 2737 17199 2762
rect 5441 2629 5491 2642
rect 5654 2629 5704 2642
rect 5862 2629 5912 2642
rect 6070 2629 6120 2642
rect 385 2588 435 2601
rect 598 2588 648 2601
rect 806 2588 856 2601
rect 1014 2588 1064 2601
rect 3872 2584 3922 2609
rect 3872 2558 3878 2584
rect 3904 2558 3922 2584
rect 3872 2532 3922 2558
rect 4080 2580 4130 2609
rect 4080 2556 4094 2580
rect 4118 2556 4130 2580
rect 4080 2532 4130 2556
rect 4288 2585 4338 2609
rect 4288 2561 4303 2585
rect 4327 2561 4338 2585
rect 4288 2532 4338 2561
rect 4501 2580 4551 2609
rect 4501 2560 4518 2580
rect 4538 2560 4551 2580
rect 4501 2532 4551 2560
rect 385 2460 435 2488
rect 385 2440 398 2460
rect 418 2440 435 2460
rect 385 2411 435 2440
rect 598 2459 648 2488
rect 598 2435 609 2459
rect 633 2435 648 2459
rect 598 2411 648 2435
rect 806 2464 856 2488
rect 806 2440 818 2464
rect 842 2440 856 2464
rect 806 2411 856 2440
rect 1014 2462 1064 2488
rect 1014 2436 1032 2462
rect 1058 2436 1064 2462
rect 1014 2411 1064 2436
rect 8928 2625 8978 2650
rect 8928 2599 8934 2625
rect 8960 2599 8978 2625
rect 8928 2573 8978 2599
rect 9136 2621 9186 2650
rect 9136 2597 9150 2621
rect 9174 2597 9186 2621
rect 9136 2573 9186 2597
rect 9344 2626 9394 2650
rect 9344 2602 9359 2626
rect 9383 2602 9394 2626
rect 9344 2573 9394 2602
rect 9557 2621 9607 2650
rect 9557 2601 9574 2621
rect 9594 2601 9607 2621
rect 12854 2693 12904 2706
rect 13062 2693 13112 2706
rect 13270 2693 13320 2706
rect 13483 2693 13533 2706
rect 11464 2638 11514 2654
rect 11677 2638 11727 2654
rect 11885 2638 11935 2654
rect 12093 2638 12143 2654
rect 13903 2656 13953 2672
rect 14111 2656 14161 2672
rect 14319 2656 14369 2672
rect 14532 2656 14582 2672
rect 17910 2734 17960 2747
rect 18118 2734 18168 2747
rect 18326 2734 18376 2747
rect 18539 2734 18589 2747
rect 16520 2679 16570 2695
rect 16733 2679 16783 2695
rect 16941 2679 16991 2695
rect 17149 2679 17199 2695
rect 18959 2697 19009 2713
rect 19167 2697 19217 2713
rect 19375 2697 19425 2713
rect 19588 2697 19638 2713
rect 15472 2634 15522 2647
rect 15685 2634 15735 2647
rect 15893 2634 15943 2647
rect 16101 2634 16151 2647
rect 9557 2573 9607 2601
rect 10416 2593 10466 2606
rect 10629 2593 10679 2606
rect 10837 2593 10887 2606
rect 11045 2593 11095 2606
rect 5441 2501 5491 2529
rect 5441 2481 5454 2501
rect 5474 2481 5491 2501
rect 3872 2419 3922 2432
rect 4080 2419 4130 2432
rect 4288 2419 4338 2432
rect 4501 2419 4551 2432
rect 5441 2452 5491 2481
rect 5654 2500 5704 2529
rect 5654 2476 5665 2500
rect 5689 2476 5704 2500
rect 5654 2452 5704 2476
rect 5862 2505 5912 2529
rect 5862 2481 5874 2505
rect 5898 2481 5912 2505
rect 5862 2452 5912 2481
rect 6070 2503 6120 2529
rect 6070 2477 6088 2503
rect 6114 2477 6120 2503
rect 6070 2452 6120 2477
rect 8928 2460 8978 2473
rect 9136 2460 9186 2473
rect 9344 2460 9394 2473
rect 9557 2460 9607 2473
rect 13903 2589 13953 2614
rect 13903 2563 13909 2589
rect 13935 2563 13953 2589
rect 13903 2537 13953 2563
rect 14111 2585 14161 2614
rect 14111 2561 14125 2585
rect 14149 2561 14161 2585
rect 14111 2537 14161 2561
rect 14319 2590 14369 2614
rect 14319 2566 14334 2590
rect 14358 2566 14369 2590
rect 14319 2537 14369 2566
rect 14532 2585 14582 2614
rect 14532 2565 14549 2585
rect 14569 2565 14582 2585
rect 14532 2537 14582 2565
rect 10416 2465 10466 2493
rect 5441 2394 5491 2410
rect 5654 2394 5704 2410
rect 5862 2394 5912 2410
rect 6070 2394 6120 2410
rect 10416 2445 10429 2465
rect 10449 2445 10466 2465
rect 385 2353 435 2369
rect 598 2353 648 2369
rect 806 2353 856 2369
rect 1014 2353 1064 2369
rect 6379 2385 6429 2398
rect 6592 2385 6642 2398
rect 6800 2385 6850 2398
rect 7008 2385 7058 2398
rect 1323 2344 1373 2357
rect 1536 2344 1586 2357
rect 1744 2344 1794 2357
rect 1952 2344 2002 2357
rect 2933 2341 2983 2357
rect 3141 2341 3191 2357
rect 3349 2341 3399 2357
rect 3562 2341 3612 2357
rect 2933 2274 2983 2299
rect 2933 2248 2939 2274
rect 2965 2248 2983 2274
rect 1323 2216 1373 2244
rect 1323 2196 1336 2216
rect 1356 2196 1373 2216
rect 1323 2167 1373 2196
rect 1536 2215 1586 2244
rect 1536 2191 1547 2215
rect 1571 2191 1586 2215
rect 1536 2167 1586 2191
rect 1744 2220 1794 2244
rect 1744 2196 1756 2220
rect 1780 2196 1794 2220
rect 1744 2167 1794 2196
rect 1952 2218 2002 2244
rect 2933 2222 2983 2248
rect 3141 2270 3191 2299
rect 3141 2246 3155 2270
rect 3179 2246 3191 2270
rect 3141 2222 3191 2246
rect 3349 2275 3399 2299
rect 3349 2251 3364 2275
rect 3388 2251 3399 2275
rect 3349 2222 3399 2251
rect 3562 2270 3612 2299
rect 3562 2250 3579 2270
rect 3599 2250 3612 2270
rect 3562 2222 3612 2250
rect 1952 2192 1970 2218
rect 1996 2192 2002 2218
rect 1952 2167 2002 2192
rect 1323 2109 1373 2125
rect 1536 2109 1586 2125
rect 1744 2109 1794 2125
rect 1952 2109 2002 2125
rect 7989 2382 8039 2398
rect 8197 2382 8247 2398
rect 8405 2382 8455 2398
rect 8618 2382 8668 2398
rect 10416 2416 10466 2445
rect 10629 2464 10679 2493
rect 10629 2440 10640 2464
rect 10664 2440 10679 2464
rect 10629 2416 10679 2440
rect 10837 2469 10887 2493
rect 10837 2445 10849 2469
rect 10873 2445 10887 2469
rect 10837 2416 10887 2445
rect 11045 2467 11095 2493
rect 11045 2441 11063 2467
rect 11089 2441 11095 2467
rect 11045 2416 11095 2441
rect 18959 2630 19009 2655
rect 18959 2604 18965 2630
rect 18991 2604 19009 2630
rect 18959 2578 19009 2604
rect 19167 2626 19217 2655
rect 19167 2602 19181 2626
rect 19205 2602 19217 2626
rect 19167 2578 19217 2602
rect 19375 2631 19425 2655
rect 19375 2607 19390 2631
rect 19414 2607 19425 2631
rect 19375 2578 19425 2607
rect 19588 2626 19638 2655
rect 19588 2606 19605 2626
rect 19625 2606 19638 2626
rect 19588 2578 19638 2606
rect 15472 2506 15522 2534
rect 15472 2486 15485 2506
rect 15505 2486 15522 2506
rect 13903 2424 13953 2437
rect 14111 2424 14161 2437
rect 14319 2424 14369 2437
rect 14532 2424 14582 2437
rect 15472 2457 15522 2486
rect 15685 2505 15735 2534
rect 15685 2481 15696 2505
rect 15720 2481 15735 2505
rect 15685 2457 15735 2481
rect 15893 2510 15943 2534
rect 15893 2486 15905 2510
rect 15929 2486 15943 2510
rect 15893 2457 15943 2486
rect 16101 2508 16151 2534
rect 16101 2482 16119 2508
rect 16145 2482 16151 2508
rect 16101 2457 16151 2482
rect 18959 2465 19009 2478
rect 19167 2465 19217 2478
rect 19375 2465 19425 2478
rect 19588 2465 19638 2478
rect 15472 2399 15522 2415
rect 15685 2399 15735 2415
rect 15893 2399 15943 2415
rect 16101 2399 16151 2415
rect 10416 2358 10466 2374
rect 10629 2358 10679 2374
rect 10837 2358 10887 2374
rect 11045 2358 11095 2374
rect 16410 2390 16460 2403
rect 16623 2390 16673 2403
rect 16831 2390 16881 2403
rect 17039 2390 17089 2403
rect 7989 2315 8039 2340
rect 7989 2289 7995 2315
rect 8021 2289 8039 2315
rect 6379 2257 6429 2285
rect 6379 2237 6392 2257
rect 6412 2237 6429 2257
rect 6379 2208 6429 2237
rect 6592 2256 6642 2285
rect 6592 2232 6603 2256
rect 6627 2232 6642 2256
rect 6592 2208 6642 2232
rect 6800 2261 6850 2285
rect 6800 2237 6812 2261
rect 6836 2237 6850 2261
rect 6800 2208 6850 2237
rect 7008 2259 7058 2285
rect 7989 2263 8039 2289
rect 8197 2311 8247 2340
rect 8197 2287 8211 2311
rect 8235 2287 8247 2311
rect 8197 2263 8247 2287
rect 8405 2316 8455 2340
rect 8405 2292 8420 2316
rect 8444 2292 8455 2316
rect 8405 2263 8455 2292
rect 8618 2311 8668 2340
rect 11354 2349 11404 2362
rect 11567 2349 11617 2362
rect 11775 2349 11825 2362
rect 11983 2349 12033 2362
rect 8618 2291 8635 2311
rect 8655 2291 8668 2311
rect 8618 2263 8668 2291
rect 7008 2233 7026 2259
rect 7052 2233 7058 2259
rect 7008 2208 7058 2233
rect 6379 2150 6429 2166
rect 6592 2150 6642 2166
rect 6800 2150 6850 2166
rect 7008 2150 7058 2166
rect 12964 2346 13014 2362
rect 13172 2346 13222 2362
rect 13380 2346 13430 2362
rect 13593 2346 13643 2362
rect 12964 2279 13014 2304
rect 12964 2253 12970 2279
rect 12996 2253 13014 2279
rect 11354 2221 11404 2249
rect 11354 2201 11367 2221
rect 11387 2201 11404 2221
rect 7989 2150 8039 2163
rect 8197 2150 8247 2163
rect 8405 2150 8455 2163
rect 8618 2150 8668 2163
rect 11354 2172 11404 2201
rect 11567 2220 11617 2249
rect 11567 2196 11578 2220
rect 11602 2196 11617 2220
rect 11567 2172 11617 2196
rect 11775 2225 11825 2249
rect 11775 2201 11787 2225
rect 11811 2201 11825 2225
rect 11775 2172 11825 2201
rect 11983 2223 12033 2249
rect 12964 2227 13014 2253
rect 13172 2275 13222 2304
rect 13172 2251 13186 2275
rect 13210 2251 13222 2275
rect 13172 2227 13222 2251
rect 13380 2280 13430 2304
rect 13380 2256 13395 2280
rect 13419 2256 13430 2280
rect 13380 2227 13430 2256
rect 13593 2275 13643 2304
rect 13593 2255 13610 2275
rect 13630 2255 13643 2275
rect 13593 2227 13643 2255
rect 11983 2197 12001 2223
rect 12027 2197 12033 2223
rect 11983 2172 12033 2197
rect 2933 2109 2983 2122
rect 3141 2109 3191 2122
rect 3349 2109 3399 2122
rect 3562 2109 3612 2122
rect 8927 2138 8977 2154
rect 9135 2138 9185 2154
rect 9343 2138 9393 2154
rect 9556 2138 9606 2154
rect 3871 2097 3921 2113
rect 4079 2097 4129 2113
rect 4287 2097 4337 2113
rect 4500 2097 4550 2113
rect 384 2034 434 2047
rect 597 2034 647 2047
rect 805 2034 855 2047
rect 1013 2034 1063 2047
rect 3871 2030 3921 2055
rect 3871 2004 3877 2030
rect 3903 2004 3921 2030
rect 3871 1978 3921 2004
rect 4079 2026 4129 2055
rect 4079 2002 4093 2026
rect 4117 2002 4129 2026
rect 4079 1978 4129 2002
rect 4287 2031 4337 2055
rect 4287 2007 4302 2031
rect 4326 2007 4337 2031
rect 4287 1978 4337 2007
rect 4500 2026 4550 2055
rect 5440 2075 5490 2088
rect 5653 2075 5703 2088
rect 5861 2075 5911 2088
rect 6069 2075 6119 2088
rect 4500 2006 4517 2026
rect 4537 2006 4550 2026
rect 4500 1978 4550 2006
rect 384 1906 434 1934
rect 384 1886 397 1906
rect 417 1886 434 1906
rect 384 1857 434 1886
rect 597 1905 647 1934
rect 597 1881 608 1905
rect 632 1881 647 1905
rect 597 1857 647 1881
rect 805 1910 855 1934
rect 805 1886 817 1910
rect 841 1886 855 1910
rect 805 1857 855 1886
rect 1013 1908 1063 1934
rect 1013 1882 1031 1908
rect 1057 1882 1063 1908
rect 1013 1857 1063 1882
rect 8927 2071 8977 2096
rect 8927 2045 8933 2071
rect 8959 2045 8977 2071
rect 8927 2019 8977 2045
rect 9135 2067 9185 2096
rect 9135 2043 9149 2067
rect 9173 2043 9185 2067
rect 9135 2019 9185 2043
rect 9343 2072 9393 2096
rect 9343 2048 9358 2072
rect 9382 2048 9393 2072
rect 9343 2019 9393 2048
rect 9556 2067 9606 2096
rect 11354 2114 11404 2130
rect 11567 2114 11617 2130
rect 11775 2114 11825 2130
rect 11983 2114 12033 2130
rect 18020 2387 18070 2403
rect 18228 2387 18278 2403
rect 18436 2387 18486 2403
rect 18649 2387 18699 2403
rect 18020 2320 18070 2345
rect 18020 2294 18026 2320
rect 18052 2294 18070 2320
rect 16410 2262 16460 2290
rect 16410 2242 16423 2262
rect 16443 2242 16460 2262
rect 16410 2213 16460 2242
rect 16623 2261 16673 2290
rect 16623 2237 16634 2261
rect 16658 2237 16673 2261
rect 16623 2213 16673 2237
rect 16831 2266 16881 2290
rect 16831 2242 16843 2266
rect 16867 2242 16881 2266
rect 16831 2213 16881 2242
rect 17039 2264 17089 2290
rect 18020 2268 18070 2294
rect 18228 2316 18278 2345
rect 18228 2292 18242 2316
rect 18266 2292 18278 2316
rect 18228 2268 18278 2292
rect 18436 2321 18486 2345
rect 18436 2297 18451 2321
rect 18475 2297 18486 2321
rect 18436 2268 18486 2297
rect 18649 2316 18699 2345
rect 18649 2296 18666 2316
rect 18686 2296 18699 2316
rect 18649 2268 18699 2296
rect 17039 2238 17057 2264
rect 17083 2238 17089 2264
rect 17039 2213 17089 2238
rect 16410 2155 16460 2171
rect 16623 2155 16673 2171
rect 16831 2155 16881 2171
rect 17039 2155 17089 2171
rect 18020 2155 18070 2168
rect 18228 2155 18278 2168
rect 18436 2155 18486 2168
rect 18649 2155 18699 2168
rect 12964 2114 13014 2127
rect 13172 2114 13222 2127
rect 13380 2114 13430 2127
rect 13593 2114 13643 2127
rect 18958 2143 19008 2159
rect 19166 2143 19216 2159
rect 19374 2143 19424 2159
rect 19587 2143 19637 2159
rect 9556 2047 9573 2067
rect 9593 2047 9606 2067
rect 13902 2102 13952 2118
rect 14110 2102 14160 2118
rect 14318 2102 14368 2118
rect 14531 2102 14581 2118
rect 9556 2019 9606 2047
rect 5440 1947 5490 1975
rect 5440 1927 5453 1947
rect 5473 1927 5490 1947
rect 5440 1898 5490 1927
rect 5653 1946 5703 1975
rect 5653 1922 5664 1946
rect 5688 1922 5703 1946
rect 5653 1898 5703 1922
rect 5861 1951 5911 1975
rect 5861 1927 5873 1951
rect 5897 1927 5911 1951
rect 5861 1898 5911 1927
rect 6069 1949 6119 1975
rect 6069 1923 6087 1949
rect 6113 1923 6119 1949
rect 6069 1898 6119 1923
rect 10415 2039 10465 2052
rect 10628 2039 10678 2052
rect 10836 2039 10886 2052
rect 11044 2039 11094 2052
rect 13902 2035 13952 2060
rect 13902 2009 13908 2035
rect 13934 2009 13952 2035
rect 13902 1983 13952 2009
rect 14110 2031 14160 2060
rect 14110 2007 14124 2031
rect 14148 2007 14160 2031
rect 14110 1983 14160 2007
rect 14318 2036 14368 2060
rect 14318 2012 14333 2036
rect 14357 2012 14368 2036
rect 14318 1983 14368 2012
rect 14531 2031 14581 2060
rect 15471 2080 15521 2093
rect 15684 2080 15734 2093
rect 15892 2080 15942 2093
rect 16100 2080 16150 2093
rect 14531 2011 14548 2031
rect 14568 2011 14581 2031
rect 14531 1983 14581 2011
rect 8927 1906 8977 1919
rect 9135 1906 9185 1919
rect 9343 1906 9393 1919
rect 9556 1906 9606 1919
rect 10415 1911 10465 1939
rect 3871 1865 3921 1878
rect 4079 1865 4129 1878
rect 4287 1865 4337 1878
rect 4500 1865 4550 1878
rect 2793 1830 2843 1846
rect 3001 1830 3051 1846
rect 3209 1830 3259 1846
rect 3422 1830 3472 1846
rect 384 1799 434 1815
rect 597 1799 647 1815
rect 805 1799 855 1815
rect 1013 1799 1063 1815
rect 7849 1871 7899 1887
rect 8057 1871 8107 1887
rect 8265 1871 8315 1887
rect 8478 1871 8528 1887
rect 5440 1840 5490 1856
rect 5653 1840 5703 1856
rect 5861 1840 5911 1856
rect 6069 1840 6119 1856
rect 10415 1891 10428 1911
rect 10448 1891 10465 1911
rect 10415 1862 10465 1891
rect 10628 1910 10678 1939
rect 10628 1886 10639 1910
rect 10663 1886 10678 1910
rect 10628 1862 10678 1886
rect 10836 1915 10886 1939
rect 10836 1891 10848 1915
rect 10872 1891 10886 1915
rect 10836 1862 10886 1891
rect 11044 1913 11094 1939
rect 11044 1887 11062 1913
rect 11088 1887 11094 1913
rect 11044 1862 11094 1887
rect 18958 2076 19008 2101
rect 18958 2050 18964 2076
rect 18990 2050 19008 2076
rect 18958 2024 19008 2050
rect 19166 2072 19216 2101
rect 19166 2048 19180 2072
rect 19204 2048 19216 2072
rect 19166 2024 19216 2048
rect 19374 2077 19424 2101
rect 19374 2053 19389 2077
rect 19413 2053 19424 2077
rect 19374 2024 19424 2053
rect 19587 2072 19637 2101
rect 19587 2052 19604 2072
rect 19624 2052 19637 2072
rect 19587 2024 19637 2052
rect 15471 1952 15521 1980
rect 15471 1932 15484 1952
rect 15504 1932 15521 1952
rect 15471 1903 15521 1932
rect 15684 1951 15734 1980
rect 15684 1927 15695 1951
rect 15719 1927 15734 1951
rect 15684 1903 15734 1927
rect 15892 1956 15942 1980
rect 15892 1932 15904 1956
rect 15928 1932 15942 1956
rect 15892 1903 15942 1932
rect 16100 1954 16150 1980
rect 16100 1928 16118 1954
rect 16144 1928 16150 1954
rect 16100 1903 16150 1928
rect 18958 1911 19008 1924
rect 19166 1911 19216 1924
rect 19374 1911 19424 1924
rect 19587 1911 19637 1924
rect 13902 1870 13952 1883
rect 14110 1870 14160 1883
rect 14318 1870 14368 1883
rect 14531 1870 14581 1883
rect 1464 1752 1514 1765
rect 1677 1752 1727 1765
rect 1885 1752 1935 1765
rect 2093 1752 2143 1765
rect 2793 1763 2843 1788
rect 2793 1737 2799 1763
rect 2825 1737 2843 1763
rect 2793 1711 2843 1737
rect 3001 1759 3051 1788
rect 3001 1735 3015 1759
rect 3039 1735 3051 1759
rect 3001 1711 3051 1735
rect 3209 1764 3259 1788
rect 3209 1740 3224 1764
rect 3248 1740 3259 1764
rect 3209 1711 3259 1740
rect 3422 1759 3472 1788
rect 6520 1793 6570 1806
rect 6733 1793 6783 1806
rect 6941 1793 6991 1806
rect 7149 1793 7199 1806
rect 7849 1804 7899 1829
rect 3422 1739 3439 1759
rect 3459 1739 3472 1759
rect 3422 1711 3472 1739
rect 1464 1624 1514 1652
rect 1464 1604 1477 1624
rect 1497 1604 1514 1624
rect 1464 1575 1514 1604
rect 1677 1623 1727 1652
rect 1677 1599 1688 1623
rect 1712 1599 1727 1623
rect 1677 1575 1727 1599
rect 1885 1628 1935 1652
rect 1885 1604 1897 1628
rect 1921 1604 1935 1628
rect 1885 1575 1935 1604
rect 2093 1626 2143 1652
rect 2093 1600 2111 1626
rect 2137 1600 2143 1626
rect 7849 1778 7855 1804
rect 7881 1778 7899 1804
rect 7849 1752 7899 1778
rect 8057 1800 8107 1829
rect 8057 1776 8071 1800
rect 8095 1776 8107 1800
rect 8057 1752 8107 1776
rect 8265 1805 8315 1829
rect 8265 1781 8280 1805
rect 8304 1781 8315 1805
rect 8265 1752 8315 1781
rect 8478 1800 8528 1829
rect 12824 1835 12874 1851
rect 13032 1835 13082 1851
rect 13240 1835 13290 1851
rect 13453 1835 13503 1851
rect 10415 1804 10465 1820
rect 10628 1804 10678 1820
rect 10836 1804 10886 1820
rect 11044 1804 11094 1820
rect 8478 1780 8495 1800
rect 8515 1780 8528 1800
rect 17880 1876 17930 1892
rect 18088 1876 18138 1892
rect 18296 1876 18346 1892
rect 18509 1876 18559 1892
rect 15471 1845 15521 1861
rect 15684 1845 15734 1861
rect 15892 1845 15942 1861
rect 16100 1845 16150 1861
rect 8478 1752 8528 1780
rect 6520 1665 6570 1693
rect 6520 1645 6533 1665
rect 6553 1645 6570 1665
rect 2093 1575 2143 1600
rect 2793 1598 2843 1611
rect 3001 1598 3051 1611
rect 3209 1598 3259 1611
rect 3422 1598 3472 1611
rect 6520 1616 6570 1645
rect 6733 1664 6783 1693
rect 6733 1640 6744 1664
rect 6768 1640 6783 1664
rect 6733 1616 6783 1640
rect 6941 1669 6991 1693
rect 6941 1645 6953 1669
rect 6977 1645 6991 1669
rect 6941 1616 6991 1645
rect 7149 1667 7199 1693
rect 7149 1641 7167 1667
rect 7193 1641 7199 1667
rect 11495 1757 11545 1770
rect 11708 1757 11758 1770
rect 11916 1757 11966 1770
rect 12124 1757 12174 1770
rect 12824 1768 12874 1793
rect 7149 1616 7199 1641
rect 7849 1639 7899 1652
rect 8057 1639 8107 1652
rect 8265 1639 8315 1652
rect 8478 1639 8528 1652
rect 12824 1742 12830 1768
rect 12856 1742 12874 1768
rect 12824 1716 12874 1742
rect 13032 1764 13082 1793
rect 13032 1740 13046 1764
rect 13070 1740 13082 1764
rect 13032 1716 13082 1740
rect 13240 1769 13290 1793
rect 13240 1745 13255 1769
rect 13279 1745 13290 1769
rect 13240 1716 13290 1745
rect 13453 1764 13503 1793
rect 16551 1798 16601 1811
rect 16764 1798 16814 1811
rect 16972 1798 17022 1811
rect 17180 1798 17230 1811
rect 17880 1809 17930 1834
rect 13453 1744 13470 1764
rect 13490 1744 13503 1764
rect 13453 1716 13503 1744
rect 11495 1629 11545 1657
rect 3873 1548 3923 1564
rect 4081 1548 4131 1564
rect 4289 1548 4339 1564
rect 4502 1548 4552 1564
rect 1464 1517 1514 1533
rect 1677 1517 1727 1533
rect 1885 1517 1935 1533
rect 2093 1517 2143 1533
rect 11495 1609 11508 1629
rect 11528 1609 11545 1629
rect 8929 1589 8979 1605
rect 9137 1589 9187 1605
rect 9345 1589 9395 1605
rect 9558 1589 9608 1605
rect 6520 1558 6570 1574
rect 6733 1558 6783 1574
rect 6941 1558 6991 1574
rect 7149 1558 7199 1574
rect 11495 1580 11545 1609
rect 11708 1628 11758 1657
rect 11708 1604 11719 1628
rect 11743 1604 11758 1628
rect 11708 1580 11758 1604
rect 11916 1633 11966 1657
rect 11916 1609 11928 1633
rect 11952 1609 11966 1633
rect 11916 1580 11966 1609
rect 12124 1631 12174 1657
rect 12124 1605 12142 1631
rect 12168 1605 12174 1631
rect 17880 1783 17886 1809
rect 17912 1783 17930 1809
rect 17880 1757 17930 1783
rect 18088 1805 18138 1834
rect 18088 1781 18102 1805
rect 18126 1781 18138 1805
rect 18088 1757 18138 1781
rect 18296 1810 18346 1834
rect 18296 1786 18311 1810
rect 18335 1786 18346 1810
rect 18296 1757 18346 1786
rect 18509 1805 18559 1834
rect 18509 1785 18526 1805
rect 18546 1785 18559 1805
rect 18509 1757 18559 1785
rect 16551 1670 16601 1698
rect 16551 1650 16564 1670
rect 16584 1650 16601 1670
rect 12124 1580 12174 1605
rect 12824 1603 12874 1616
rect 13032 1603 13082 1616
rect 13240 1603 13290 1616
rect 13453 1603 13503 1616
rect 16551 1621 16601 1650
rect 16764 1669 16814 1698
rect 16764 1645 16775 1669
rect 16799 1645 16814 1669
rect 16764 1621 16814 1645
rect 16972 1674 17022 1698
rect 16972 1650 16984 1674
rect 17008 1650 17022 1674
rect 16972 1621 17022 1650
rect 17180 1672 17230 1698
rect 17180 1646 17198 1672
rect 17224 1646 17230 1672
rect 17180 1621 17230 1646
rect 17880 1644 17930 1657
rect 18088 1644 18138 1657
rect 18296 1644 18346 1657
rect 18509 1644 18559 1657
rect 5442 1526 5492 1539
rect 5655 1526 5705 1539
rect 5863 1526 5913 1539
rect 6071 1526 6121 1539
rect 386 1485 436 1498
rect 599 1485 649 1498
rect 807 1485 857 1498
rect 1015 1485 1065 1498
rect 3873 1481 3923 1506
rect 3873 1455 3879 1481
rect 3905 1455 3923 1481
rect 3873 1429 3923 1455
rect 4081 1477 4131 1506
rect 4081 1453 4095 1477
rect 4119 1453 4131 1477
rect 4081 1429 4131 1453
rect 4289 1482 4339 1506
rect 4289 1458 4304 1482
rect 4328 1458 4339 1482
rect 4289 1429 4339 1458
rect 4502 1477 4552 1506
rect 4502 1457 4519 1477
rect 4539 1457 4552 1477
rect 4502 1429 4552 1457
rect 386 1357 436 1385
rect 386 1337 399 1357
rect 419 1337 436 1357
rect 386 1308 436 1337
rect 599 1356 649 1385
rect 599 1332 610 1356
rect 634 1332 649 1356
rect 599 1308 649 1332
rect 807 1361 857 1385
rect 807 1337 819 1361
rect 843 1337 857 1361
rect 807 1308 857 1337
rect 1015 1359 1065 1385
rect 1015 1333 1033 1359
rect 1059 1333 1065 1359
rect 1015 1308 1065 1333
rect 8929 1522 8979 1547
rect 8929 1496 8935 1522
rect 8961 1496 8979 1522
rect 8929 1470 8979 1496
rect 9137 1518 9187 1547
rect 9137 1494 9151 1518
rect 9175 1494 9187 1518
rect 9137 1470 9187 1494
rect 9345 1523 9395 1547
rect 9345 1499 9360 1523
rect 9384 1499 9395 1523
rect 9345 1470 9395 1499
rect 9558 1518 9608 1547
rect 9558 1498 9575 1518
rect 9595 1498 9608 1518
rect 13904 1553 13954 1569
rect 14112 1553 14162 1569
rect 14320 1553 14370 1569
rect 14533 1553 14583 1569
rect 11495 1522 11545 1538
rect 11708 1522 11758 1538
rect 11916 1522 11966 1538
rect 12124 1522 12174 1538
rect 18960 1594 19010 1610
rect 19168 1594 19218 1610
rect 19376 1594 19426 1610
rect 19589 1594 19639 1610
rect 16551 1563 16601 1579
rect 16764 1563 16814 1579
rect 16972 1563 17022 1579
rect 17180 1563 17230 1579
rect 15473 1531 15523 1544
rect 15686 1531 15736 1544
rect 15894 1531 15944 1544
rect 16102 1531 16152 1544
rect 9558 1470 9608 1498
rect 10417 1490 10467 1503
rect 10630 1490 10680 1503
rect 10838 1490 10888 1503
rect 11046 1490 11096 1503
rect 5442 1398 5492 1426
rect 5442 1378 5455 1398
rect 5475 1378 5492 1398
rect 3873 1316 3923 1329
rect 4081 1316 4131 1329
rect 4289 1316 4339 1329
rect 4502 1316 4552 1329
rect 5442 1349 5492 1378
rect 5655 1397 5705 1426
rect 5655 1373 5666 1397
rect 5690 1373 5705 1397
rect 5655 1349 5705 1373
rect 5863 1402 5913 1426
rect 5863 1378 5875 1402
rect 5899 1378 5913 1402
rect 5863 1349 5913 1378
rect 6071 1400 6121 1426
rect 6071 1374 6089 1400
rect 6115 1374 6121 1400
rect 6071 1349 6121 1374
rect 8929 1357 8979 1370
rect 9137 1357 9187 1370
rect 9345 1357 9395 1370
rect 9558 1357 9608 1370
rect 13904 1486 13954 1511
rect 13904 1460 13910 1486
rect 13936 1460 13954 1486
rect 13904 1434 13954 1460
rect 14112 1482 14162 1511
rect 14112 1458 14126 1482
rect 14150 1458 14162 1482
rect 14112 1434 14162 1458
rect 14320 1487 14370 1511
rect 14320 1463 14335 1487
rect 14359 1463 14370 1487
rect 14320 1434 14370 1463
rect 14533 1482 14583 1511
rect 14533 1462 14550 1482
rect 14570 1462 14583 1482
rect 14533 1434 14583 1462
rect 10417 1362 10467 1390
rect 5442 1291 5492 1307
rect 5655 1291 5705 1307
rect 5863 1291 5913 1307
rect 6071 1291 6121 1307
rect 10417 1342 10430 1362
rect 10450 1342 10467 1362
rect 386 1250 436 1266
rect 599 1250 649 1266
rect 807 1250 857 1266
rect 1015 1250 1065 1266
rect 6380 1282 6430 1295
rect 6593 1282 6643 1295
rect 6801 1282 6851 1295
rect 7009 1282 7059 1295
rect 1324 1241 1374 1254
rect 1537 1241 1587 1254
rect 1745 1241 1795 1254
rect 1953 1241 2003 1254
rect 2934 1238 2984 1254
rect 3142 1238 3192 1254
rect 3350 1238 3400 1254
rect 3563 1238 3613 1254
rect 2934 1171 2984 1196
rect 2934 1145 2940 1171
rect 2966 1145 2984 1171
rect 1324 1113 1374 1141
rect 1324 1093 1337 1113
rect 1357 1093 1374 1113
rect 1324 1064 1374 1093
rect 1537 1112 1587 1141
rect 1537 1088 1548 1112
rect 1572 1088 1587 1112
rect 1537 1064 1587 1088
rect 1745 1117 1795 1141
rect 1745 1093 1757 1117
rect 1781 1093 1795 1117
rect 1745 1064 1795 1093
rect 1953 1115 2003 1141
rect 2934 1119 2984 1145
rect 3142 1167 3192 1196
rect 3142 1143 3156 1167
rect 3180 1143 3192 1167
rect 3142 1119 3192 1143
rect 3350 1172 3400 1196
rect 3350 1148 3365 1172
rect 3389 1148 3400 1172
rect 3350 1119 3400 1148
rect 3563 1167 3613 1196
rect 3563 1147 3580 1167
rect 3600 1147 3613 1167
rect 3563 1119 3613 1147
rect 1953 1089 1971 1115
rect 1997 1089 2003 1115
rect 1953 1064 2003 1089
rect 1324 1006 1374 1022
rect 1537 1006 1587 1022
rect 1745 1006 1795 1022
rect 1953 1006 2003 1022
rect 7990 1279 8040 1295
rect 8198 1279 8248 1295
rect 8406 1279 8456 1295
rect 8619 1279 8669 1295
rect 10417 1313 10467 1342
rect 10630 1361 10680 1390
rect 10630 1337 10641 1361
rect 10665 1337 10680 1361
rect 10630 1313 10680 1337
rect 10838 1366 10888 1390
rect 10838 1342 10850 1366
rect 10874 1342 10888 1366
rect 10838 1313 10888 1342
rect 11046 1364 11096 1390
rect 11046 1338 11064 1364
rect 11090 1338 11096 1364
rect 11046 1313 11096 1338
rect 18960 1527 19010 1552
rect 18960 1501 18966 1527
rect 18992 1501 19010 1527
rect 18960 1475 19010 1501
rect 19168 1523 19218 1552
rect 19168 1499 19182 1523
rect 19206 1499 19218 1523
rect 19168 1475 19218 1499
rect 19376 1528 19426 1552
rect 19376 1504 19391 1528
rect 19415 1504 19426 1528
rect 19376 1475 19426 1504
rect 19589 1523 19639 1552
rect 19589 1503 19606 1523
rect 19626 1503 19639 1523
rect 19589 1475 19639 1503
rect 15473 1403 15523 1431
rect 15473 1383 15486 1403
rect 15506 1383 15523 1403
rect 13904 1321 13954 1334
rect 14112 1321 14162 1334
rect 14320 1321 14370 1334
rect 14533 1321 14583 1334
rect 15473 1354 15523 1383
rect 15686 1402 15736 1431
rect 15686 1378 15697 1402
rect 15721 1378 15736 1402
rect 15686 1354 15736 1378
rect 15894 1407 15944 1431
rect 15894 1383 15906 1407
rect 15930 1383 15944 1407
rect 15894 1354 15944 1383
rect 16102 1405 16152 1431
rect 16102 1379 16120 1405
rect 16146 1379 16152 1405
rect 16102 1354 16152 1379
rect 18960 1362 19010 1375
rect 19168 1362 19218 1375
rect 19376 1362 19426 1375
rect 19589 1362 19639 1375
rect 15473 1296 15523 1312
rect 15686 1296 15736 1312
rect 15894 1296 15944 1312
rect 16102 1296 16152 1312
rect 10417 1255 10467 1271
rect 10630 1255 10680 1271
rect 10838 1255 10888 1271
rect 11046 1255 11096 1271
rect 16411 1287 16461 1300
rect 16624 1287 16674 1300
rect 16832 1287 16882 1300
rect 17040 1287 17090 1300
rect 7990 1212 8040 1237
rect 7990 1186 7996 1212
rect 8022 1186 8040 1212
rect 6380 1154 6430 1182
rect 6380 1134 6393 1154
rect 6413 1134 6430 1154
rect 6380 1105 6430 1134
rect 6593 1153 6643 1182
rect 6593 1129 6604 1153
rect 6628 1129 6643 1153
rect 6593 1105 6643 1129
rect 6801 1158 6851 1182
rect 6801 1134 6813 1158
rect 6837 1134 6851 1158
rect 6801 1105 6851 1134
rect 7009 1156 7059 1182
rect 7990 1160 8040 1186
rect 8198 1208 8248 1237
rect 8198 1184 8212 1208
rect 8236 1184 8248 1208
rect 8198 1160 8248 1184
rect 8406 1213 8456 1237
rect 8406 1189 8421 1213
rect 8445 1189 8456 1213
rect 8406 1160 8456 1189
rect 8619 1208 8669 1237
rect 11355 1246 11405 1259
rect 11568 1246 11618 1259
rect 11776 1246 11826 1259
rect 11984 1246 12034 1259
rect 8619 1188 8636 1208
rect 8656 1188 8669 1208
rect 8619 1160 8669 1188
rect 7009 1130 7027 1156
rect 7053 1130 7059 1156
rect 7009 1105 7059 1130
rect 6380 1047 6430 1063
rect 6593 1047 6643 1063
rect 6801 1047 6851 1063
rect 7009 1047 7059 1063
rect 12965 1243 13015 1259
rect 13173 1243 13223 1259
rect 13381 1243 13431 1259
rect 13594 1243 13644 1259
rect 12965 1176 13015 1201
rect 12965 1150 12971 1176
rect 12997 1150 13015 1176
rect 11355 1118 11405 1146
rect 11355 1098 11368 1118
rect 11388 1098 11405 1118
rect 7990 1047 8040 1060
rect 8198 1047 8248 1060
rect 8406 1047 8456 1060
rect 8619 1047 8669 1060
rect 11355 1069 11405 1098
rect 11568 1117 11618 1146
rect 11568 1093 11579 1117
rect 11603 1093 11618 1117
rect 11568 1069 11618 1093
rect 11776 1122 11826 1146
rect 11776 1098 11788 1122
rect 11812 1098 11826 1122
rect 11776 1069 11826 1098
rect 11984 1120 12034 1146
rect 12965 1124 13015 1150
rect 13173 1172 13223 1201
rect 13173 1148 13187 1172
rect 13211 1148 13223 1172
rect 13173 1124 13223 1148
rect 13381 1177 13431 1201
rect 13381 1153 13396 1177
rect 13420 1153 13431 1177
rect 13381 1124 13431 1153
rect 13594 1172 13644 1201
rect 13594 1152 13611 1172
rect 13631 1152 13644 1172
rect 13594 1124 13644 1152
rect 11984 1094 12002 1120
rect 12028 1094 12034 1120
rect 11984 1069 12034 1094
rect 2934 1006 2984 1019
rect 3142 1006 3192 1019
rect 3350 1006 3400 1019
rect 3563 1006 3613 1019
rect 8928 1035 8978 1051
rect 9136 1035 9186 1051
rect 9344 1035 9394 1051
rect 9557 1035 9607 1051
rect 3872 994 3922 1010
rect 4080 994 4130 1010
rect 4288 994 4338 1010
rect 4501 994 4551 1010
rect 385 931 435 944
rect 598 931 648 944
rect 806 931 856 944
rect 1014 931 1064 944
rect 3872 927 3922 952
rect 3872 901 3878 927
rect 3904 901 3922 927
rect 3872 875 3922 901
rect 4080 923 4130 952
rect 4080 899 4094 923
rect 4118 899 4130 923
rect 4080 875 4130 899
rect 4288 928 4338 952
rect 4288 904 4303 928
rect 4327 904 4338 928
rect 4288 875 4338 904
rect 4501 923 4551 952
rect 5441 972 5491 985
rect 5654 972 5704 985
rect 5862 972 5912 985
rect 6070 972 6120 985
rect 4501 903 4518 923
rect 4538 903 4551 923
rect 4501 875 4551 903
rect 385 803 435 831
rect 385 783 398 803
rect 418 783 435 803
rect 385 754 435 783
rect 598 802 648 831
rect 598 778 609 802
rect 633 778 648 802
rect 598 754 648 778
rect 806 807 856 831
rect 806 783 818 807
rect 842 783 856 807
rect 806 754 856 783
rect 1014 805 1064 831
rect 1014 779 1032 805
rect 1058 779 1064 805
rect 1014 754 1064 779
rect 8928 968 8978 993
rect 8928 942 8934 968
rect 8960 942 8978 968
rect 8928 916 8978 942
rect 9136 964 9186 993
rect 9136 940 9150 964
rect 9174 940 9186 964
rect 9136 916 9186 940
rect 9344 969 9394 993
rect 9344 945 9359 969
rect 9383 945 9394 969
rect 9344 916 9394 945
rect 9557 964 9607 993
rect 11355 1011 11405 1027
rect 11568 1011 11618 1027
rect 11776 1011 11826 1027
rect 11984 1011 12034 1027
rect 18021 1284 18071 1300
rect 18229 1284 18279 1300
rect 18437 1284 18487 1300
rect 18650 1284 18700 1300
rect 18021 1217 18071 1242
rect 18021 1191 18027 1217
rect 18053 1191 18071 1217
rect 16411 1159 16461 1187
rect 16411 1139 16424 1159
rect 16444 1139 16461 1159
rect 16411 1110 16461 1139
rect 16624 1158 16674 1187
rect 16624 1134 16635 1158
rect 16659 1134 16674 1158
rect 16624 1110 16674 1134
rect 16832 1163 16882 1187
rect 16832 1139 16844 1163
rect 16868 1139 16882 1163
rect 16832 1110 16882 1139
rect 17040 1161 17090 1187
rect 18021 1165 18071 1191
rect 18229 1213 18279 1242
rect 18229 1189 18243 1213
rect 18267 1189 18279 1213
rect 18229 1165 18279 1189
rect 18437 1218 18487 1242
rect 18437 1194 18452 1218
rect 18476 1194 18487 1218
rect 18437 1165 18487 1194
rect 18650 1213 18700 1242
rect 18650 1193 18667 1213
rect 18687 1193 18700 1213
rect 18650 1165 18700 1193
rect 17040 1135 17058 1161
rect 17084 1135 17090 1161
rect 17040 1110 17090 1135
rect 16411 1052 16461 1068
rect 16624 1052 16674 1068
rect 16832 1052 16882 1068
rect 17040 1052 17090 1068
rect 18021 1052 18071 1065
rect 18229 1052 18279 1065
rect 18437 1052 18487 1065
rect 18650 1052 18700 1065
rect 12965 1011 13015 1024
rect 13173 1011 13223 1024
rect 13381 1011 13431 1024
rect 13594 1011 13644 1024
rect 18959 1040 19009 1056
rect 19167 1040 19217 1056
rect 19375 1040 19425 1056
rect 19588 1040 19638 1056
rect 9557 944 9574 964
rect 9594 944 9607 964
rect 13903 999 13953 1015
rect 14111 999 14161 1015
rect 14319 999 14369 1015
rect 14532 999 14582 1015
rect 9557 916 9607 944
rect 5441 844 5491 872
rect 5441 824 5454 844
rect 5474 824 5491 844
rect 5441 795 5491 824
rect 5654 843 5704 872
rect 5654 819 5665 843
rect 5689 819 5704 843
rect 5654 795 5704 819
rect 5862 848 5912 872
rect 5862 824 5874 848
rect 5898 824 5912 848
rect 5862 795 5912 824
rect 6070 846 6120 872
rect 6070 820 6088 846
rect 6114 820 6120 846
rect 6070 795 6120 820
rect 10416 936 10466 949
rect 10629 936 10679 949
rect 10837 936 10887 949
rect 11045 936 11095 949
rect 13903 932 13953 957
rect 13903 906 13909 932
rect 13935 906 13953 932
rect 13903 880 13953 906
rect 14111 928 14161 957
rect 14111 904 14125 928
rect 14149 904 14161 928
rect 14111 880 14161 904
rect 14319 933 14369 957
rect 14319 909 14334 933
rect 14358 909 14369 933
rect 14319 880 14369 909
rect 14532 928 14582 957
rect 15472 977 15522 990
rect 15685 977 15735 990
rect 15893 977 15943 990
rect 16101 977 16151 990
rect 14532 908 14549 928
rect 14569 908 14582 928
rect 14532 880 14582 908
rect 8928 803 8978 816
rect 9136 803 9186 816
rect 9344 803 9394 816
rect 9557 803 9607 816
rect 10416 808 10466 836
rect 3872 762 3922 775
rect 4080 762 4130 775
rect 4288 762 4338 775
rect 4501 762 4551 775
rect 385 696 435 712
rect 598 696 648 712
rect 806 696 856 712
rect 1014 696 1064 712
rect 5441 737 5491 753
rect 5654 737 5704 753
rect 5862 737 5912 753
rect 6070 737 6120 753
rect 10416 788 10429 808
rect 10449 788 10466 808
rect 10416 759 10466 788
rect 10629 807 10679 836
rect 10629 783 10640 807
rect 10664 783 10679 807
rect 10629 759 10679 783
rect 10837 812 10887 836
rect 10837 788 10849 812
rect 10873 788 10887 812
rect 10837 759 10887 788
rect 11045 810 11095 836
rect 11045 784 11063 810
rect 11089 784 11095 810
rect 11045 759 11095 784
rect 18959 973 19009 998
rect 18959 947 18965 973
rect 18991 947 19009 973
rect 18959 921 19009 947
rect 19167 969 19217 998
rect 19167 945 19181 969
rect 19205 945 19217 969
rect 19167 921 19217 945
rect 19375 974 19425 998
rect 19375 950 19390 974
rect 19414 950 19425 974
rect 19375 921 19425 950
rect 19588 969 19638 998
rect 19588 949 19605 969
rect 19625 949 19638 969
rect 19588 921 19638 949
rect 15472 849 15522 877
rect 15472 829 15485 849
rect 15505 829 15522 849
rect 15472 800 15522 829
rect 15685 848 15735 877
rect 15685 824 15696 848
rect 15720 824 15735 848
rect 15685 800 15735 824
rect 15893 853 15943 877
rect 15893 829 15905 853
rect 15929 829 15943 853
rect 15893 800 15943 829
rect 16101 851 16151 877
rect 16101 825 16119 851
rect 16145 825 16151 851
rect 16101 800 16151 825
rect 18959 808 19009 821
rect 19167 808 19217 821
rect 19375 808 19425 821
rect 19588 808 19638 821
rect 13903 767 13953 780
rect 14111 767 14161 780
rect 14319 767 14369 780
rect 14532 767 14582 780
rect 10416 701 10466 717
rect 10629 701 10679 717
rect 10837 701 10887 717
rect 11045 701 11095 717
rect 15472 742 15522 758
rect 15685 742 15735 758
rect 15893 742 15943 758
rect 16101 742 16151 758
rect 6688 413 6738 426
rect 6901 413 6951 426
rect 7109 413 7159 426
rect 7317 413 7367 426
rect 1632 372 1682 385
rect 1845 372 1895 385
rect 2053 372 2103 385
rect 2261 372 2311 385
rect 4582 352 4632 365
rect 4795 352 4845 365
rect 5003 352 5053 365
rect 5211 352 5261 365
rect 1632 244 1682 272
rect 1632 224 1645 244
rect 1665 224 1682 244
rect 1632 195 1682 224
rect 1845 243 1895 272
rect 1845 219 1856 243
rect 1880 219 1895 243
rect 1845 195 1895 219
rect 2053 248 2103 272
rect 2053 224 2065 248
rect 2089 224 2103 248
rect 2053 195 2103 224
rect 2261 246 2311 272
rect 16719 418 16769 431
rect 16932 418 16982 431
rect 17140 418 17190 431
rect 17348 418 17398 431
rect 11663 377 11713 390
rect 11876 377 11926 390
rect 12084 377 12134 390
rect 12292 377 12342 390
rect 6688 285 6738 313
rect 6688 265 6701 285
rect 6721 265 6738 285
rect 2261 220 2279 246
rect 2305 220 2311 246
rect 2261 195 2311 220
rect 4582 224 4632 252
rect 4582 204 4595 224
rect 4615 204 4632 224
rect 4582 175 4632 204
rect 4795 223 4845 252
rect 4795 199 4806 223
rect 4830 199 4845 223
rect 4795 175 4845 199
rect 5003 228 5053 252
rect 5003 204 5015 228
rect 5039 204 5053 228
rect 5003 175 5053 204
rect 5211 226 5261 252
rect 6688 236 6738 265
rect 6901 284 6951 313
rect 6901 260 6912 284
rect 6936 260 6951 284
rect 6901 236 6951 260
rect 7109 289 7159 313
rect 7109 265 7121 289
rect 7145 265 7159 289
rect 7109 236 7159 265
rect 7317 287 7367 313
rect 7317 261 7335 287
rect 7361 261 7367 287
rect 14613 357 14663 370
rect 14826 357 14876 370
rect 15034 357 15084 370
rect 15242 357 15292 370
rect 7317 236 7367 261
rect 11663 249 11713 277
rect 9516 236 9566 249
rect 9729 236 9779 249
rect 9937 236 9987 249
rect 10145 236 10195 249
rect 5211 200 5229 226
rect 5255 200 5261 226
rect 5211 175 5261 200
rect 6688 178 6738 194
rect 6901 178 6951 194
rect 7109 178 7159 194
rect 7317 178 7367 194
rect 1632 137 1682 153
rect 1845 137 1895 153
rect 2053 137 2103 153
rect 2261 137 2311 153
rect 4582 117 4632 133
rect 4795 117 4845 133
rect 5003 117 5053 133
rect 5211 117 5261 133
rect 11663 229 11676 249
rect 11696 229 11713 249
rect 11663 200 11713 229
rect 11876 248 11926 277
rect 11876 224 11887 248
rect 11911 224 11926 248
rect 11876 200 11926 224
rect 12084 253 12134 277
rect 12084 229 12096 253
rect 12120 229 12134 253
rect 12084 200 12134 229
rect 12292 251 12342 277
rect 16719 290 16769 318
rect 16719 270 16732 290
rect 16752 270 16769 290
rect 12292 225 12310 251
rect 12336 225 12342 251
rect 12292 200 12342 225
rect 14613 229 14663 257
rect 14613 209 14626 229
rect 14646 209 14663 229
rect 14613 180 14663 209
rect 14826 228 14876 257
rect 14826 204 14837 228
rect 14861 204 14876 228
rect 14826 180 14876 204
rect 15034 233 15084 257
rect 15034 209 15046 233
rect 15070 209 15084 233
rect 15034 180 15084 209
rect 15242 231 15292 257
rect 16719 241 16769 270
rect 16932 289 16982 318
rect 16932 265 16943 289
rect 16967 265 16982 289
rect 16932 241 16982 265
rect 17140 294 17190 318
rect 17140 270 17152 294
rect 17176 270 17190 294
rect 17140 241 17190 270
rect 17348 292 17398 318
rect 17348 266 17366 292
rect 17392 266 17398 292
rect 17348 241 17398 266
rect 15242 205 15260 231
rect 15286 205 15292 231
rect 15242 180 15292 205
rect 16719 183 16769 199
rect 16932 183 16982 199
rect 17140 183 17190 199
rect 17348 183 17398 199
rect 11663 142 11713 158
rect 11876 142 11926 158
rect 12084 142 12134 158
rect 12292 142 12342 158
rect 9516 108 9566 136
rect 9516 88 9529 108
rect 9549 88 9566 108
rect 9516 59 9566 88
rect 9729 107 9779 136
rect 9729 83 9740 107
rect 9764 83 9779 107
rect 9729 59 9779 83
rect 9937 112 9987 136
rect 9937 88 9949 112
rect 9973 88 9987 112
rect 9937 59 9987 88
rect 10145 110 10195 136
rect 14613 122 14663 138
rect 14826 122 14876 138
rect 15034 122 15084 138
rect 15242 122 15292 138
rect 10145 84 10163 110
rect 10189 84 10195 110
rect 10145 59 10195 84
rect 9516 1 9566 17
rect 9729 1 9779 17
rect 9937 1 9987 17
rect 10145 1 10195 17
<< polycont >>
rect 3875 9176 3901 9202
rect 4091 9174 4115 9198
rect 4300 9179 4324 9203
rect 4515 9178 4535 9198
rect 395 9058 415 9078
rect 606 9053 630 9077
rect 815 9058 839 9082
rect 1029 9054 1055 9080
rect 8931 9217 8957 9243
rect 9147 9215 9171 9239
rect 9356 9220 9380 9244
rect 9571 9219 9591 9239
rect 5451 9099 5471 9119
rect 5662 9094 5686 9118
rect 5871 9099 5895 9123
rect 6085 9095 6111 9121
rect 13906 9181 13932 9207
rect 14122 9179 14146 9203
rect 14331 9184 14355 9208
rect 14546 9183 14566 9203
rect 10426 9063 10446 9083
rect 2936 8866 2962 8892
rect 1333 8814 1353 8834
rect 1544 8809 1568 8833
rect 1753 8814 1777 8838
rect 3152 8864 3176 8888
rect 3361 8869 3385 8893
rect 3576 8868 3596 8888
rect 1967 8810 1993 8836
rect 10637 9058 10661 9082
rect 10846 9063 10870 9087
rect 11060 9059 11086 9085
rect 18962 9222 18988 9248
rect 19178 9220 19202 9244
rect 19387 9225 19411 9249
rect 19602 9224 19622 9244
rect 15482 9104 15502 9124
rect 15693 9099 15717 9123
rect 15902 9104 15926 9128
rect 16116 9100 16142 9126
rect 7992 8907 8018 8933
rect 6389 8855 6409 8875
rect 6600 8850 6624 8874
rect 6809 8855 6833 8879
rect 8208 8905 8232 8929
rect 8417 8910 8441 8934
rect 8632 8909 8652 8929
rect 7023 8851 7049 8877
rect 12967 8871 12993 8897
rect 11364 8819 11384 8839
rect 11575 8814 11599 8838
rect 11784 8819 11808 8843
rect 13183 8869 13207 8893
rect 13392 8874 13416 8898
rect 13607 8873 13627 8893
rect 11998 8815 12024 8841
rect 3874 8622 3900 8648
rect 4090 8620 4114 8644
rect 4299 8625 4323 8649
rect 4514 8624 4534 8644
rect 394 8504 414 8524
rect 605 8499 629 8523
rect 814 8504 838 8528
rect 1028 8500 1054 8526
rect 8930 8663 8956 8689
rect 9146 8661 9170 8685
rect 9355 8666 9379 8690
rect 18023 8912 18049 8938
rect 16420 8860 16440 8880
rect 16631 8855 16655 8879
rect 16840 8860 16864 8884
rect 18239 8910 18263 8934
rect 18448 8915 18472 8939
rect 18663 8914 18683 8934
rect 17054 8856 17080 8882
rect 9570 8665 9590 8685
rect 5450 8545 5470 8565
rect 5661 8540 5685 8564
rect 5870 8545 5894 8569
rect 6084 8541 6110 8567
rect 13905 8627 13931 8653
rect 14121 8625 14145 8649
rect 14330 8630 14354 8654
rect 14545 8629 14565 8649
rect 10425 8509 10445 8529
rect 10636 8504 10660 8528
rect 10845 8509 10869 8533
rect 11059 8505 11085 8531
rect 18961 8668 18987 8694
rect 19177 8666 19201 8690
rect 19386 8671 19410 8695
rect 19601 8670 19621 8690
rect 15481 8550 15501 8570
rect 15692 8545 15716 8569
rect 15901 8550 15925 8574
rect 16115 8546 16141 8572
rect 2796 8355 2822 8381
rect 3012 8353 3036 8377
rect 3221 8358 3245 8382
rect 3436 8357 3456 8377
rect 1474 8222 1494 8242
rect 1685 8217 1709 8241
rect 1894 8222 1918 8246
rect 2108 8218 2134 8244
rect 7852 8396 7878 8422
rect 8068 8394 8092 8418
rect 8277 8399 8301 8423
rect 8492 8398 8512 8418
rect 6530 8263 6550 8283
rect 6741 8258 6765 8282
rect 6950 8263 6974 8287
rect 7164 8259 7190 8285
rect 12827 8360 12853 8386
rect 13043 8358 13067 8382
rect 13252 8363 13276 8387
rect 13467 8362 13487 8382
rect 11505 8227 11525 8247
rect 11716 8222 11740 8246
rect 11925 8227 11949 8251
rect 12139 8223 12165 8249
rect 17883 8401 17909 8427
rect 18099 8399 18123 8423
rect 18308 8404 18332 8428
rect 18523 8403 18543 8423
rect 16561 8268 16581 8288
rect 16772 8263 16796 8287
rect 16981 8268 17005 8292
rect 17195 8264 17221 8290
rect 3876 8073 3902 8099
rect 4092 8071 4116 8095
rect 4301 8076 4325 8100
rect 4516 8075 4536 8095
rect 396 7955 416 7975
rect 607 7950 631 7974
rect 816 7955 840 7979
rect 1030 7951 1056 7977
rect 8932 8114 8958 8140
rect 9148 8112 9172 8136
rect 9357 8117 9381 8141
rect 9572 8116 9592 8136
rect 5452 7996 5472 8016
rect 5663 7991 5687 8015
rect 5872 7996 5896 8020
rect 6086 7992 6112 8018
rect 13907 8078 13933 8104
rect 14123 8076 14147 8100
rect 14332 8081 14356 8105
rect 14547 8080 14567 8100
rect 10427 7960 10447 7980
rect 2937 7763 2963 7789
rect 1334 7711 1354 7731
rect 1545 7706 1569 7730
rect 1754 7711 1778 7735
rect 3153 7761 3177 7785
rect 3362 7766 3386 7790
rect 3577 7765 3597 7785
rect 1968 7707 1994 7733
rect 10638 7955 10662 7979
rect 10847 7960 10871 7984
rect 11061 7956 11087 7982
rect 18963 8119 18989 8145
rect 19179 8117 19203 8141
rect 19388 8122 19412 8146
rect 19603 8121 19623 8141
rect 15483 8001 15503 8021
rect 15694 7996 15718 8020
rect 15903 8001 15927 8025
rect 16117 7997 16143 8023
rect 7993 7804 8019 7830
rect 6390 7752 6410 7772
rect 6601 7747 6625 7771
rect 6810 7752 6834 7776
rect 8209 7802 8233 7826
rect 8418 7807 8442 7831
rect 8633 7806 8653 7826
rect 7024 7748 7050 7774
rect 12968 7768 12994 7794
rect 11365 7716 11385 7736
rect 11576 7711 11600 7735
rect 11785 7716 11809 7740
rect 13184 7766 13208 7790
rect 13393 7771 13417 7795
rect 13608 7770 13628 7790
rect 11999 7712 12025 7738
rect 3875 7519 3901 7545
rect 4091 7517 4115 7541
rect 4300 7522 4324 7546
rect 4515 7521 4535 7541
rect 395 7401 415 7421
rect 606 7396 630 7420
rect 815 7401 839 7425
rect 1029 7397 1055 7423
rect 8931 7560 8957 7586
rect 9147 7558 9171 7582
rect 9356 7563 9380 7587
rect 18024 7809 18050 7835
rect 16421 7757 16441 7777
rect 16632 7752 16656 7776
rect 16841 7757 16865 7781
rect 18240 7807 18264 7831
rect 18449 7812 18473 7836
rect 18664 7811 18684 7831
rect 17055 7753 17081 7779
rect 9571 7562 9591 7582
rect 5451 7442 5471 7462
rect 5662 7437 5686 7461
rect 5871 7442 5895 7466
rect 6085 7438 6111 7464
rect 13906 7524 13932 7550
rect 14122 7522 14146 7546
rect 14331 7527 14355 7551
rect 14546 7526 14566 7546
rect 10426 7406 10446 7426
rect 10637 7401 10661 7425
rect 10846 7406 10870 7430
rect 11060 7402 11086 7428
rect 18962 7565 18988 7591
rect 19178 7563 19202 7587
rect 19387 7568 19411 7592
rect 19602 7567 19622 7587
rect 15482 7447 15502 7467
rect 15693 7442 15717 7466
rect 15902 7447 15926 7471
rect 16116 7443 16142 7469
rect 2827 7239 2853 7265
rect 3043 7237 3067 7261
rect 3252 7242 3276 7266
rect 3467 7241 3487 7261
rect 7883 7280 7909 7306
rect 8099 7278 8123 7302
rect 8308 7283 8332 7307
rect 8523 7282 8543 7302
rect 1444 7132 1464 7152
rect 1655 7127 1679 7151
rect 1864 7132 1888 7156
rect 2078 7128 2104 7154
rect 6500 7173 6520 7193
rect 6711 7168 6735 7192
rect 6920 7173 6944 7197
rect 7134 7169 7160 7195
rect 12858 7244 12884 7270
rect 13074 7242 13098 7266
rect 13283 7247 13307 7271
rect 13498 7246 13518 7266
rect 17914 7285 17940 7311
rect 18130 7283 18154 7307
rect 18339 7288 18363 7312
rect 18554 7287 18574 7307
rect 11475 7137 11495 7157
rect 11686 7132 11710 7156
rect 11895 7137 11919 7161
rect 12109 7133 12135 7159
rect 16531 7178 16551 7198
rect 16742 7173 16766 7197
rect 16951 7178 16975 7202
rect 17165 7174 17191 7200
rect 3876 6970 3902 6996
rect 4092 6968 4116 6992
rect 4301 6973 4325 6997
rect 4516 6972 4536 6992
rect 396 6852 416 6872
rect 607 6847 631 6871
rect 816 6852 840 6876
rect 1030 6848 1056 6874
rect 8932 7011 8958 7037
rect 9148 7009 9172 7033
rect 9357 7014 9381 7038
rect 9572 7013 9592 7033
rect 5452 6893 5472 6913
rect 5663 6888 5687 6912
rect 5872 6893 5896 6917
rect 6086 6889 6112 6915
rect 13907 6975 13933 7001
rect 14123 6973 14147 6997
rect 14332 6978 14356 7002
rect 14547 6977 14567 6997
rect 10427 6857 10447 6877
rect 2937 6660 2963 6686
rect 1334 6608 1354 6628
rect 1545 6603 1569 6627
rect 1754 6608 1778 6632
rect 3153 6658 3177 6682
rect 3362 6663 3386 6687
rect 3577 6662 3597 6682
rect 1968 6604 1994 6630
rect 10638 6852 10662 6876
rect 10847 6857 10871 6881
rect 11061 6853 11087 6879
rect 18963 7016 18989 7042
rect 19179 7014 19203 7038
rect 19388 7019 19412 7043
rect 19603 7018 19623 7038
rect 15483 6898 15503 6918
rect 15694 6893 15718 6917
rect 15903 6898 15927 6922
rect 16117 6894 16143 6920
rect 7993 6701 8019 6727
rect 6390 6649 6410 6669
rect 6601 6644 6625 6668
rect 6810 6649 6834 6673
rect 8209 6699 8233 6723
rect 8418 6704 8442 6728
rect 8633 6703 8653 6723
rect 7024 6645 7050 6671
rect 12968 6665 12994 6691
rect 11365 6613 11385 6633
rect 11576 6608 11600 6632
rect 11785 6613 11809 6637
rect 13184 6663 13208 6687
rect 13393 6668 13417 6692
rect 13608 6667 13628 6687
rect 11999 6609 12025 6635
rect 3875 6416 3901 6442
rect 4091 6414 4115 6438
rect 4300 6419 4324 6443
rect 4515 6418 4535 6438
rect 395 6298 415 6318
rect 606 6293 630 6317
rect 815 6298 839 6322
rect 1029 6294 1055 6320
rect 8931 6457 8957 6483
rect 9147 6455 9171 6479
rect 9356 6460 9380 6484
rect 18024 6706 18050 6732
rect 16421 6654 16441 6674
rect 16632 6649 16656 6673
rect 16841 6654 16865 6678
rect 18240 6704 18264 6728
rect 18449 6709 18473 6733
rect 18664 6708 18684 6728
rect 17055 6650 17081 6676
rect 9571 6459 9591 6479
rect 5451 6339 5471 6359
rect 5662 6334 5686 6358
rect 5871 6339 5895 6363
rect 6085 6335 6111 6361
rect 13906 6421 13932 6447
rect 14122 6419 14146 6443
rect 14331 6424 14355 6448
rect 14546 6423 14566 6443
rect 10426 6303 10446 6323
rect 10637 6298 10661 6322
rect 10846 6303 10870 6327
rect 11060 6299 11086 6325
rect 18962 6462 18988 6488
rect 19178 6460 19202 6484
rect 19387 6465 19411 6489
rect 19602 6464 19622 6484
rect 15482 6344 15502 6364
rect 15693 6339 15717 6363
rect 15902 6344 15926 6368
rect 16116 6340 16142 6366
rect 2797 6149 2823 6175
rect 3013 6147 3037 6171
rect 3222 6152 3246 6176
rect 3437 6151 3457 6171
rect 1475 6016 1495 6036
rect 1686 6011 1710 6035
rect 1895 6016 1919 6040
rect 2109 6012 2135 6038
rect 7853 6190 7879 6216
rect 8069 6188 8093 6212
rect 8278 6193 8302 6217
rect 8493 6192 8513 6212
rect 6531 6057 6551 6077
rect 6742 6052 6766 6076
rect 6951 6057 6975 6081
rect 7165 6053 7191 6079
rect 12828 6154 12854 6180
rect 13044 6152 13068 6176
rect 13253 6157 13277 6181
rect 13468 6156 13488 6176
rect 11506 6021 11526 6041
rect 11717 6016 11741 6040
rect 11926 6021 11950 6045
rect 12140 6017 12166 6043
rect 17884 6195 17910 6221
rect 18100 6193 18124 6217
rect 18309 6198 18333 6222
rect 18524 6197 18544 6217
rect 16562 6062 16582 6082
rect 16773 6057 16797 6081
rect 16982 6062 17006 6086
rect 17196 6058 17222 6084
rect 3877 5867 3903 5893
rect 4093 5865 4117 5889
rect 4302 5870 4326 5894
rect 4517 5869 4537 5889
rect 397 5749 417 5769
rect 608 5744 632 5768
rect 817 5749 841 5773
rect 1031 5745 1057 5771
rect 8933 5908 8959 5934
rect 9149 5906 9173 5930
rect 9358 5911 9382 5935
rect 9573 5910 9593 5930
rect 5453 5790 5473 5810
rect 5664 5785 5688 5809
rect 5873 5790 5897 5814
rect 6087 5786 6113 5812
rect 13908 5872 13934 5898
rect 14124 5870 14148 5894
rect 14333 5875 14357 5899
rect 14548 5874 14568 5894
rect 10428 5754 10448 5774
rect 2938 5557 2964 5583
rect 1335 5505 1355 5525
rect 1546 5500 1570 5524
rect 1755 5505 1779 5529
rect 3154 5555 3178 5579
rect 3363 5560 3387 5584
rect 3578 5559 3598 5579
rect 1969 5501 1995 5527
rect 10639 5749 10663 5773
rect 10848 5754 10872 5778
rect 11062 5750 11088 5776
rect 18964 5913 18990 5939
rect 19180 5911 19204 5935
rect 19389 5916 19413 5940
rect 19604 5915 19624 5935
rect 15484 5795 15504 5815
rect 15695 5790 15719 5814
rect 15904 5795 15928 5819
rect 16118 5791 16144 5817
rect 7994 5598 8020 5624
rect 6391 5546 6411 5566
rect 6602 5541 6626 5565
rect 6811 5546 6835 5570
rect 8210 5596 8234 5620
rect 8419 5601 8443 5625
rect 8634 5600 8654 5620
rect 7025 5542 7051 5568
rect 12969 5562 12995 5588
rect 11366 5510 11386 5530
rect 11577 5505 11601 5529
rect 11786 5510 11810 5534
rect 13185 5560 13209 5584
rect 13394 5565 13418 5589
rect 13609 5564 13629 5584
rect 12000 5506 12026 5532
rect 3876 5313 3902 5339
rect 4092 5311 4116 5335
rect 4301 5316 4325 5340
rect 4516 5315 4536 5335
rect 396 5195 416 5215
rect 607 5190 631 5214
rect 816 5195 840 5219
rect 1030 5191 1056 5217
rect 8932 5354 8958 5380
rect 9148 5352 9172 5376
rect 9357 5357 9381 5381
rect 18025 5603 18051 5629
rect 16422 5551 16442 5571
rect 16633 5546 16657 5570
rect 16842 5551 16866 5575
rect 18241 5601 18265 5625
rect 18450 5606 18474 5630
rect 18665 5605 18685 5625
rect 17056 5547 17082 5573
rect 9572 5356 9592 5376
rect 5452 5236 5472 5256
rect 5663 5231 5687 5255
rect 5872 5236 5896 5260
rect 6086 5232 6112 5258
rect 13907 5318 13933 5344
rect 14123 5316 14147 5340
rect 14332 5321 14356 5345
rect 14547 5320 14567 5340
rect 2829 5027 2855 5053
rect 3045 5025 3069 5049
rect 3254 5030 3278 5054
rect 3469 5029 3489 5049
rect 10427 5200 10447 5220
rect 10638 5195 10662 5219
rect 10847 5200 10871 5224
rect 11061 5196 11087 5222
rect 18963 5359 18989 5385
rect 19179 5357 19203 5381
rect 19388 5362 19412 5386
rect 19603 5361 19623 5381
rect 15483 5241 15503 5261
rect 15694 5236 15718 5260
rect 15903 5241 15927 5265
rect 16117 5237 16143 5263
rect 7885 5068 7911 5094
rect 8101 5066 8125 5090
rect 8310 5071 8334 5095
rect 8525 5070 8545 5090
rect 1444 4932 1464 4952
rect 1655 4927 1679 4951
rect 1864 4932 1888 4956
rect 2078 4928 2104 4954
rect 6500 4973 6520 4993
rect 6711 4968 6735 4992
rect 6920 4973 6944 4997
rect 7134 4969 7160 4995
rect 12860 5032 12886 5058
rect 13076 5030 13100 5054
rect 13285 5035 13309 5059
rect 13500 5034 13520 5054
rect 17916 5073 17942 5099
rect 18132 5071 18156 5095
rect 18341 5076 18365 5100
rect 18556 5075 18576 5095
rect 11475 4937 11495 4957
rect 11686 4932 11710 4956
rect 11895 4937 11919 4961
rect 12109 4933 12135 4959
rect 3877 4764 3903 4790
rect 4093 4762 4117 4786
rect 4302 4767 4326 4791
rect 4517 4766 4537 4786
rect 397 4646 417 4666
rect 608 4641 632 4665
rect 817 4646 841 4670
rect 1031 4642 1057 4668
rect 8933 4805 8959 4831
rect 9149 4803 9173 4827
rect 9358 4808 9382 4832
rect 9573 4807 9593 4827
rect 16531 4978 16551 4998
rect 16742 4973 16766 4997
rect 16951 4978 16975 5002
rect 17165 4974 17191 5000
rect 5453 4687 5473 4707
rect 5664 4682 5688 4706
rect 5873 4687 5897 4711
rect 6087 4683 6113 4709
rect 13908 4769 13934 4795
rect 14124 4767 14148 4791
rect 14333 4772 14357 4796
rect 14548 4771 14568 4791
rect 10428 4651 10448 4671
rect 2938 4454 2964 4480
rect 1335 4402 1355 4422
rect 1546 4397 1570 4421
rect 1755 4402 1779 4426
rect 3154 4452 3178 4476
rect 3363 4457 3387 4481
rect 3578 4456 3598 4476
rect 1969 4398 1995 4424
rect 10639 4646 10663 4670
rect 10848 4651 10872 4675
rect 11062 4647 11088 4673
rect 18964 4810 18990 4836
rect 19180 4808 19204 4832
rect 19389 4813 19413 4837
rect 19604 4812 19624 4832
rect 15484 4692 15504 4712
rect 15695 4687 15719 4711
rect 15904 4692 15928 4716
rect 16118 4688 16144 4714
rect 7994 4495 8020 4521
rect 6391 4443 6411 4463
rect 6602 4438 6626 4462
rect 6811 4443 6835 4467
rect 8210 4493 8234 4517
rect 8419 4498 8443 4522
rect 8634 4497 8654 4517
rect 7025 4439 7051 4465
rect 12969 4459 12995 4485
rect 11366 4407 11386 4427
rect 11577 4402 11601 4426
rect 11786 4407 11810 4431
rect 13185 4457 13209 4481
rect 13394 4462 13418 4486
rect 13609 4461 13629 4481
rect 12000 4403 12026 4429
rect 3876 4210 3902 4236
rect 4092 4208 4116 4232
rect 4301 4213 4325 4237
rect 4516 4212 4536 4232
rect 396 4092 416 4112
rect 607 4087 631 4111
rect 816 4092 840 4116
rect 1030 4088 1056 4114
rect 8932 4251 8958 4277
rect 9148 4249 9172 4273
rect 9357 4254 9381 4278
rect 18025 4500 18051 4526
rect 16422 4448 16442 4468
rect 16633 4443 16657 4467
rect 16842 4448 16866 4472
rect 18241 4498 18265 4522
rect 18450 4503 18474 4527
rect 18665 4502 18685 4522
rect 17056 4444 17082 4470
rect 9572 4253 9592 4273
rect 5452 4133 5472 4153
rect 5663 4128 5687 4152
rect 5872 4133 5896 4157
rect 6086 4129 6112 4155
rect 13907 4215 13933 4241
rect 14123 4213 14147 4237
rect 14332 4218 14356 4242
rect 14547 4217 14567 4237
rect 10427 4097 10447 4117
rect 10638 4092 10662 4116
rect 10847 4097 10871 4121
rect 11061 4093 11087 4119
rect 18963 4256 18989 4282
rect 19179 4254 19203 4278
rect 19388 4259 19412 4283
rect 19603 4258 19623 4278
rect 15483 4138 15503 4158
rect 15694 4133 15718 4157
rect 15903 4138 15927 4162
rect 16117 4134 16143 4160
rect 2798 3943 2824 3969
rect 3014 3941 3038 3965
rect 3223 3946 3247 3970
rect 3438 3945 3458 3965
rect 1476 3810 1496 3830
rect 1687 3805 1711 3829
rect 1896 3810 1920 3834
rect 2110 3806 2136 3832
rect 7854 3984 7880 4010
rect 8070 3982 8094 4006
rect 8279 3987 8303 4011
rect 8494 3986 8514 4006
rect 6532 3851 6552 3871
rect 6743 3846 6767 3870
rect 6952 3851 6976 3875
rect 7166 3847 7192 3873
rect 12829 3948 12855 3974
rect 13045 3946 13069 3970
rect 13254 3951 13278 3975
rect 13469 3950 13489 3970
rect 11507 3815 11527 3835
rect 11718 3810 11742 3834
rect 11927 3815 11951 3839
rect 12141 3811 12167 3837
rect 17885 3989 17911 4015
rect 18101 3987 18125 4011
rect 18310 3992 18334 4016
rect 18525 3991 18545 4011
rect 16563 3856 16583 3876
rect 16774 3851 16798 3875
rect 16983 3856 17007 3880
rect 17197 3852 17223 3878
rect 3878 3661 3904 3687
rect 4094 3659 4118 3683
rect 4303 3664 4327 3688
rect 4518 3663 4538 3683
rect 398 3543 418 3563
rect 609 3538 633 3562
rect 818 3543 842 3567
rect 1032 3539 1058 3565
rect 8934 3702 8960 3728
rect 9150 3700 9174 3724
rect 9359 3705 9383 3729
rect 9574 3704 9594 3724
rect 5454 3584 5474 3604
rect 5665 3579 5689 3603
rect 5874 3584 5898 3608
rect 6088 3580 6114 3606
rect 13909 3666 13935 3692
rect 14125 3664 14149 3688
rect 14334 3669 14358 3693
rect 14549 3668 14569 3688
rect 10429 3548 10449 3568
rect 2939 3351 2965 3377
rect 1336 3299 1356 3319
rect 1547 3294 1571 3318
rect 1756 3299 1780 3323
rect 3155 3349 3179 3373
rect 3364 3354 3388 3378
rect 3579 3353 3599 3373
rect 1970 3295 1996 3321
rect 10640 3543 10664 3567
rect 10849 3548 10873 3572
rect 11063 3544 11089 3570
rect 18965 3707 18991 3733
rect 19181 3705 19205 3729
rect 19390 3710 19414 3734
rect 19605 3709 19625 3729
rect 15485 3589 15505 3609
rect 15696 3584 15720 3608
rect 15905 3589 15929 3613
rect 16119 3585 16145 3611
rect 7995 3392 8021 3418
rect 6392 3340 6412 3360
rect 6603 3335 6627 3359
rect 6812 3340 6836 3364
rect 8211 3390 8235 3414
rect 8420 3395 8444 3419
rect 8635 3394 8655 3414
rect 7026 3336 7052 3362
rect 12970 3356 12996 3382
rect 11367 3304 11387 3324
rect 11578 3299 11602 3323
rect 11787 3304 11811 3328
rect 13186 3354 13210 3378
rect 13395 3359 13419 3383
rect 13610 3358 13630 3378
rect 12001 3300 12027 3326
rect 3877 3107 3903 3133
rect 4093 3105 4117 3129
rect 4302 3110 4326 3134
rect 4517 3109 4537 3129
rect 397 2989 417 3009
rect 608 2984 632 3008
rect 817 2989 841 3013
rect 1031 2985 1057 3011
rect 8933 3148 8959 3174
rect 9149 3146 9173 3170
rect 9358 3151 9382 3175
rect 18026 3397 18052 3423
rect 16423 3345 16443 3365
rect 16634 3340 16658 3364
rect 16843 3345 16867 3369
rect 18242 3395 18266 3419
rect 18451 3400 18475 3424
rect 18666 3399 18686 3419
rect 17057 3341 17083 3367
rect 9573 3150 9593 3170
rect 5453 3030 5473 3050
rect 5664 3025 5688 3049
rect 5873 3030 5897 3054
rect 6087 3026 6113 3052
rect 13908 3112 13934 3138
rect 14124 3110 14148 3134
rect 14333 3115 14357 3139
rect 14548 3114 14568 3134
rect 10428 2994 10448 3014
rect 10639 2989 10663 3013
rect 10848 2994 10872 3018
rect 11062 2990 11088 3016
rect 18964 3153 18990 3179
rect 19180 3151 19204 3175
rect 19389 3156 19413 3180
rect 19604 3155 19624 3175
rect 15484 3035 15504 3055
rect 15695 3030 15719 3054
rect 15904 3035 15928 3059
rect 16118 3031 16144 3057
rect 2829 2827 2855 2853
rect 3045 2825 3069 2849
rect 3254 2830 3278 2854
rect 3469 2829 3489 2849
rect 7885 2868 7911 2894
rect 8101 2866 8125 2890
rect 8310 2871 8334 2895
rect 8525 2870 8545 2890
rect 1446 2720 1466 2740
rect 1657 2715 1681 2739
rect 1866 2720 1890 2744
rect 2080 2716 2106 2742
rect 6502 2761 6522 2781
rect 6713 2756 6737 2780
rect 6922 2761 6946 2785
rect 7136 2757 7162 2783
rect 12860 2832 12886 2858
rect 13076 2830 13100 2854
rect 13285 2835 13309 2859
rect 13500 2834 13520 2854
rect 17916 2873 17942 2899
rect 18132 2871 18156 2895
rect 18341 2876 18365 2900
rect 18556 2875 18576 2895
rect 11477 2725 11497 2745
rect 11688 2720 11712 2744
rect 11897 2725 11921 2749
rect 12111 2721 12137 2747
rect 16533 2766 16553 2786
rect 16744 2761 16768 2785
rect 16953 2766 16977 2790
rect 17167 2762 17193 2788
rect 3878 2558 3904 2584
rect 4094 2556 4118 2580
rect 4303 2561 4327 2585
rect 4518 2560 4538 2580
rect 398 2440 418 2460
rect 609 2435 633 2459
rect 818 2440 842 2464
rect 1032 2436 1058 2462
rect 8934 2599 8960 2625
rect 9150 2597 9174 2621
rect 9359 2602 9383 2626
rect 9574 2601 9594 2621
rect 5454 2481 5474 2501
rect 5665 2476 5689 2500
rect 5874 2481 5898 2505
rect 6088 2477 6114 2503
rect 13909 2563 13935 2589
rect 14125 2561 14149 2585
rect 14334 2566 14358 2590
rect 14549 2565 14569 2585
rect 10429 2445 10449 2465
rect 2939 2248 2965 2274
rect 1336 2196 1356 2216
rect 1547 2191 1571 2215
rect 1756 2196 1780 2220
rect 3155 2246 3179 2270
rect 3364 2251 3388 2275
rect 3579 2250 3599 2270
rect 1970 2192 1996 2218
rect 10640 2440 10664 2464
rect 10849 2445 10873 2469
rect 11063 2441 11089 2467
rect 18965 2604 18991 2630
rect 19181 2602 19205 2626
rect 19390 2607 19414 2631
rect 19605 2606 19625 2626
rect 15485 2486 15505 2506
rect 15696 2481 15720 2505
rect 15905 2486 15929 2510
rect 16119 2482 16145 2508
rect 7995 2289 8021 2315
rect 6392 2237 6412 2257
rect 6603 2232 6627 2256
rect 6812 2237 6836 2261
rect 8211 2287 8235 2311
rect 8420 2292 8444 2316
rect 8635 2291 8655 2311
rect 7026 2233 7052 2259
rect 12970 2253 12996 2279
rect 11367 2201 11387 2221
rect 11578 2196 11602 2220
rect 11787 2201 11811 2225
rect 13186 2251 13210 2275
rect 13395 2256 13419 2280
rect 13610 2255 13630 2275
rect 12001 2197 12027 2223
rect 3877 2004 3903 2030
rect 4093 2002 4117 2026
rect 4302 2007 4326 2031
rect 4517 2006 4537 2026
rect 397 1886 417 1906
rect 608 1881 632 1905
rect 817 1886 841 1910
rect 1031 1882 1057 1908
rect 8933 2045 8959 2071
rect 9149 2043 9173 2067
rect 9358 2048 9382 2072
rect 18026 2294 18052 2320
rect 16423 2242 16443 2262
rect 16634 2237 16658 2261
rect 16843 2242 16867 2266
rect 18242 2292 18266 2316
rect 18451 2297 18475 2321
rect 18666 2296 18686 2316
rect 17057 2238 17083 2264
rect 9573 2047 9593 2067
rect 5453 1927 5473 1947
rect 5664 1922 5688 1946
rect 5873 1927 5897 1951
rect 6087 1923 6113 1949
rect 13908 2009 13934 2035
rect 14124 2007 14148 2031
rect 14333 2012 14357 2036
rect 14548 2011 14568 2031
rect 10428 1891 10448 1911
rect 10639 1886 10663 1910
rect 10848 1891 10872 1915
rect 11062 1887 11088 1913
rect 18964 2050 18990 2076
rect 19180 2048 19204 2072
rect 19389 2053 19413 2077
rect 19604 2052 19624 2072
rect 15484 1932 15504 1952
rect 15695 1927 15719 1951
rect 15904 1932 15928 1956
rect 16118 1928 16144 1954
rect 2799 1737 2825 1763
rect 3015 1735 3039 1759
rect 3224 1740 3248 1764
rect 3439 1739 3459 1759
rect 1477 1604 1497 1624
rect 1688 1599 1712 1623
rect 1897 1604 1921 1628
rect 2111 1600 2137 1626
rect 7855 1778 7881 1804
rect 8071 1776 8095 1800
rect 8280 1781 8304 1805
rect 8495 1780 8515 1800
rect 6533 1645 6553 1665
rect 6744 1640 6768 1664
rect 6953 1645 6977 1669
rect 7167 1641 7193 1667
rect 12830 1742 12856 1768
rect 13046 1740 13070 1764
rect 13255 1745 13279 1769
rect 13470 1744 13490 1764
rect 11508 1609 11528 1629
rect 11719 1604 11743 1628
rect 11928 1609 11952 1633
rect 12142 1605 12168 1631
rect 17886 1783 17912 1809
rect 18102 1781 18126 1805
rect 18311 1786 18335 1810
rect 18526 1785 18546 1805
rect 16564 1650 16584 1670
rect 16775 1645 16799 1669
rect 16984 1650 17008 1674
rect 17198 1646 17224 1672
rect 3879 1455 3905 1481
rect 4095 1453 4119 1477
rect 4304 1458 4328 1482
rect 4519 1457 4539 1477
rect 399 1337 419 1357
rect 610 1332 634 1356
rect 819 1337 843 1361
rect 1033 1333 1059 1359
rect 8935 1496 8961 1522
rect 9151 1494 9175 1518
rect 9360 1499 9384 1523
rect 9575 1498 9595 1518
rect 5455 1378 5475 1398
rect 5666 1373 5690 1397
rect 5875 1378 5899 1402
rect 6089 1374 6115 1400
rect 13910 1460 13936 1486
rect 14126 1458 14150 1482
rect 14335 1463 14359 1487
rect 14550 1462 14570 1482
rect 10430 1342 10450 1362
rect 2940 1145 2966 1171
rect 1337 1093 1357 1113
rect 1548 1088 1572 1112
rect 1757 1093 1781 1117
rect 3156 1143 3180 1167
rect 3365 1148 3389 1172
rect 3580 1147 3600 1167
rect 1971 1089 1997 1115
rect 10641 1337 10665 1361
rect 10850 1342 10874 1366
rect 11064 1338 11090 1364
rect 18966 1501 18992 1527
rect 19182 1499 19206 1523
rect 19391 1504 19415 1528
rect 19606 1503 19626 1523
rect 15486 1383 15506 1403
rect 15697 1378 15721 1402
rect 15906 1383 15930 1407
rect 16120 1379 16146 1405
rect 7996 1186 8022 1212
rect 6393 1134 6413 1154
rect 6604 1129 6628 1153
rect 6813 1134 6837 1158
rect 8212 1184 8236 1208
rect 8421 1189 8445 1213
rect 8636 1188 8656 1208
rect 7027 1130 7053 1156
rect 12971 1150 12997 1176
rect 11368 1098 11388 1118
rect 11579 1093 11603 1117
rect 11788 1098 11812 1122
rect 13187 1148 13211 1172
rect 13396 1153 13420 1177
rect 13611 1152 13631 1172
rect 12002 1094 12028 1120
rect 3878 901 3904 927
rect 4094 899 4118 923
rect 4303 904 4327 928
rect 4518 903 4538 923
rect 398 783 418 803
rect 609 778 633 802
rect 818 783 842 807
rect 1032 779 1058 805
rect 8934 942 8960 968
rect 9150 940 9174 964
rect 9359 945 9383 969
rect 18027 1191 18053 1217
rect 16424 1139 16444 1159
rect 16635 1134 16659 1158
rect 16844 1139 16868 1163
rect 18243 1189 18267 1213
rect 18452 1194 18476 1218
rect 18667 1193 18687 1213
rect 17058 1135 17084 1161
rect 9574 944 9594 964
rect 5454 824 5474 844
rect 5665 819 5689 843
rect 5874 824 5898 848
rect 6088 820 6114 846
rect 13909 906 13935 932
rect 14125 904 14149 928
rect 14334 909 14358 933
rect 14549 908 14569 928
rect 10429 788 10449 808
rect 10640 783 10664 807
rect 10849 788 10873 812
rect 11063 784 11089 810
rect 18965 947 18991 973
rect 19181 945 19205 969
rect 19390 950 19414 974
rect 19605 949 19625 969
rect 15485 829 15505 849
rect 15696 824 15720 848
rect 15905 829 15929 853
rect 16119 825 16145 851
rect 1645 224 1665 244
rect 1856 219 1880 243
rect 2065 224 2089 248
rect 6701 265 6721 285
rect 2279 220 2305 246
rect 4595 204 4615 224
rect 4806 199 4830 223
rect 5015 204 5039 228
rect 6912 260 6936 284
rect 7121 265 7145 289
rect 7335 261 7361 287
rect 5229 200 5255 226
rect 11676 229 11696 249
rect 11887 224 11911 248
rect 12096 229 12120 253
rect 16732 270 16752 290
rect 12310 225 12336 251
rect 14626 209 14646 229
rect 14837 204 14861 228
rect 15046 209 15070 233
rect 16943 265 16967 289
rect 17152 270 17176 294
rect 17366 266 17392 292
rect 15260 205 15286 231
rect 9529 88 9549 108
rect 9740 83 9764 107
rect 9949 88 9973 112
rect 10163 84 10189 110
<< ndiffres >>
rect 5151 9343 5208 9362
rect 5151 9340 5172 9343
rect 95 9302 152 9321
rect 5057 9325 5172 9340
rect 5190 9325 5208 9343
rect 95 9299 116 9302
rect 1 9284 116 9299
rect 134 9284 152 9302
rect 5057 9302 5208 9325
rect 15182 9348 15239 9367
rect 15182 9345 15203 9348
rect 1 9261 152 9284
rect 1 9225 43 9261
rect 5057 9266 5099 9302
rect 10126 9307 10183 9326
rect 15088 9330 15203 9345
rect 15221 9330 15239 9348
rect 10126 9304 10147 9307
rect 10032 9289 10147 9304
rect 10165 9289 10183 9307
rect 15088 9307 15239 9330
rect 5056 9265 5156 9266
rect 5056 9244 5212 9265
rect 0 9224 100 9225
rect 0 9203 156 9224
rect 0 9185 118 9203
rect 136 9185 156 9203
rect 0 9181 156 9185
rect 95 9165 156 9181
rect 95 9115 152 9134
rect 95 9112 116 9115
rect 1 9097 116 9112
rect 134 9097 152 9115
rect 5056 9226 5174 9244
rect 5192 9226 5212 9244
rect 5056 9222 5212 9226
rect 5151 9206 5212 9222
rect 4773 9167 4834 9183
rect 4773 9163 4929 9167
rect 1 9074 152 9097
rect 1 9038 43 9074
rect 0 9037 100 9038
rect 0 9016 156 9037
rect 0 8998 118 9016
rect 136 8998 156 9016
rect 0 8994 156 8998
rect 95 8978 156 8994
rect 4773 9145 4793 9163
rect 4811 9145 4929 9163
rect 5151 9156 5208 9175
rect 5151 9153 5172 9156
rect 4773 9124 4929 9145
rect 4829 9123 4929 9124
rect 5057 9138 5172 9153
rect 5190 9138 5208 9156
rect 10032 9266 10183 9289
rect 10032 9230 10074 9266
rect 15088 9271 15130 9307
rect 15087 9270 15187 9271
rect 15087 9249 15243 9270
rect 10031 9229 10131 9230
rect 9829 9208 9890 9224
rect 10031 9208 10187 9229
rect 9829 9204 9985 9208
rect 4886 9087 4928 9123
rect 4777 9064 4928 9087
rect 5057 9115 5208 9138
rect 5057 9079 5099 9115
rect 4777 9046 4795 9064
rect 4813 9049 4928 9064
rect 5056 9078 5156 9079
rect 5056 9057 5212 9078
rect 4813 9046 4834 9049
rect 4777 9027 4834 9046
rect 5056 9039 5174 9057
rect 5192 9039 5212 9057
rect 5056 9035 5212 9039
rect 5151 9019 5212 9035
rect 9829 9186 9849 9204
rect 9867 9186 9985 9204
rect 10031 9190 10149 9208
rect 10167 9190 10187 9208
rect 10031 9186 10187 9190
rect 9829 9165 9985 9186
rect 10126 9170 10187 9186
rect 9885 9164 9985 9165
rect 9942 9128 9984 9164
rect 9833 9105 9984 9128
rect 10126 9120 10183 9139
rect 10126 9117 10147 9120
rect 9833 9087 9851 9105
rect 9869 9090 9984 9105
rect 10032 9102 10147 9117
rect 10165 9102 10183 9120
rect 15087 9231 15205 9249
rect 15223 9231 15243 9249
rect 15087 9227 15243 9231
rect 15182 9211 15243 9227
rect 14804 9172 14865 9188
rect 14804 9168 14960 9172
rect 9869 9087 9890 9090
rect 9833 9068 9890 9087
rect 10032 9079 10183 9102
rect 10032 9043 10074 9079
rect 95 8886 152 8905
rect 95 8883 116 8886
rect 1 8868 116 8883
rect 134 8868 152 8886
rect 1 8845 152 8868
rect 4773 8937 4834 8953
rect 4773 8933 4929 8937
rect 1 8809 43 8845
rect 0 8808 100 8809
rect 0 8787 156 8808
rect 0 8769 118 8787
rect 136 8769 156 8787
rect 4773 8915 4793 8933
rect 4811 8915 4929 8933
rect 5151 8927 5208 8946
rect 5151 8924 5172 8927
rect 4773 8894 4929 8915
rect 4829 8893 4929 8894
rect 5057 8909 5172 8924
rect 5190 8909 5208 8927
rect 4886 8857 4928 8893
rect 0 8765 156 8769
rect 95 8749 156 8765
rect 4777 8834 4928 8857
rect 5057 8886 5208 8909
rect 10031 9042 10131 9043
rect 10031 9021 10187 9042
rect 10031 9003 10149 9021
rect 10167 9003 10187 9021
rect 10031 8999 10187 9003
rect 9829 8978 9890 8994
rect 10126 8983 10187 8999
rect 14804 9150 14824 9168
rect 14842 9150 14960 9168
rect 15182 9161 15239 9180
rect 15182 9158 15203 9161
rect 14804 9129 14960 9150
rect 14860 9128 14960 9129
rect 15088 9143 15203 9158
rect 15221 9143 15239 9161
rect 19860 9213 19921 9229
rect 19860 9209 20016 9213
rect 14917 9092 14959 9128
rect 14808 9069 14959 9092
rect 15088 9120 15239 9143
rect 15088 9084 15130 9120
rect 14808 9051 14826 9069
rect 14844 9054 14959 9069
rect 15087 9083 15187 9084
rect 15087 9062 15243 9083
rect 14844 9051 14865 9054
rect 14808 9032 14865 9051
rect 15087 9044 15205 9062
rect 15223 9044 15243 9062
rect 15087 9040 15243 9044
rect 15182 9024 15243 9040
rect 19860 9191 19880 9209
rect 19898 9191 20016 9209
rect 19860 9170 20016 9191
rect 19916 9169 20016 9170
rect 19973 9133 20015 9169
rect 19864 9110 20015 9133
rect 19864 9092 19882 9110
rect 19900 9095 20015 9110
rect 19900 9092 19921 9095
rect 19864 9073 19921 9092
rect 9829 8974 9985 8978
rect 5057 8850 5099 8886
rect 4777 8816 4795 8834
rect 4813 8819 4928 8834
rect 5056 8849 5156 8850
rect 5056 8828 5212 8849
rect 4813 8816 4834 8819
rect 4777 8797 4834 8816
rect 5056 8810 5174 8828
rect 5192 8810 5212 8828
rect 9829 8956 9849 8974
rect 9867 8956 9985 8974
rect 9829 8935 9985 8956
rect 9885 8934 9985 8935
rect 9942 8898 9984 8934
rect 5056 8806 5212 8810
rect 5151 8790 5212 8806
rect 9833 8875 9984 8898
rect 10126 8891 10183 8910
rect 10126 8888 10147 8891
rect 9833 8857 9851 8875
rect 9869 8860 9984 8875
rect 10032 8873 10147 8888
rect 10165 8873 10183 8891
rect 9869 8857 9890 8860
rect 9833 8838 9890 8857
rect 10032 8850 10183 8873
rect 14804 8942 14865 8958
rect 14804 8938 14960 8942
rect 10032 8814 10074 8850
rect 10031 8813 10131 8814
rect 10031 8792 10187 8813
rect 10031 8774 10149 8792
rect 10167 8774 10187 8792
rect 14804 8920 14824 8938
rect 14842 8920 14960 8938
rect 15182 8932 15239 8951
rect 15182 8929 15203 8932
rect 14804 8899 14960 8920
rect 14860 8898 14960 8899
rect 15088 8914 15203 8929
rect 15221 8914 15239 8932
rect 14917 8862 14959 8898
rect 10031 8770 10187 8774
rect 95 8656 152 8675
rect 95 8653 116 8656
rect 1 8638 116 8653
rect 134 8638 152 8656
rect 1 8615 152 8638
rect 1 8579 43 8615
rect 0 8578 100 8579
rect 0 8557 156 8578
rect 0 8539 118 8557
rect 136 8539 156 8557
rect 4773 8708 4834 8724
rect 4773 8704 4929 8708
rect 4773 8686 4793 8704
rect 4811 8686 4929 8704
rect 5151 8697 5208 8716
rect 5151 8694 5172 8697
rect 4773 8665 4929 8686
rect 4829 8664 4929 8665
rect 5057 8679 5172 8694
rect 5190 8679 5208 8697
rect 4886 8628 4928 8664
rect 4777 8605 4928 8628
rect 5057 8656 5208 8679
rect 5057 8620 5099 8656
rect 0 8535 156 8539
rect 95 8519 156 8535
rect 4777 8587 4795 8605
rect 4813 8590 4928 8605
rect 5056 8619 5156 8620
rect 5056 8598 5212 8619
rect 4813 8587 4834 8590
rect 4777 8568 4834 8587
rect 5056 8580 5174 8598
rect 5192 8580 5212 8598
rect 9829 8749 9890 8765
rect 10126 8754 10187 8770
rect 9829 8745 9985 8749
rect 9829 8727 9849 8745
rect 9867 8727 9985 8745
rect 9829 8706 9985 8727
rect 9885 8705 9985 8706
rect 14808 8839 14959 8862
rect 15088 8891 15239 8914
rect 19860 8983 19921 8999
rect 19860 8979 20016 8983
rect 15088 8855 15130 8891
rect 14808 8821 14826 8839
rect 14844 8824 14959 8839
rect 15087 8854 15187 8855
rect 15087 8833 15243 8854
rect 14844 8821 14865 8824
rect 14808 8802 14865 8821
rect 15087 8815 15205 8833
rect 15223 8815 15243 8833
rect 19860 8961 19880 8979
rect 19898 8961 20016 8979
rect 19860 8940 20016 8961
rect 19916 8939 20016 8940
rect 19973 8903 20015 8939
rect 15087 8811 15243 8815
rect 15182 8795 15243 8811
rect 19864 8880 20015 8903
rect 19864 8862 19882 8880
rect 19900 8865 20015 8880
rect 19900 8862 19921 8865
rect 19864 8843 19921 8862
rect 9942 8669 9984 8705
rect 9833 8646 9984 8669
rect 10126 8661 10183 8680
rect 10126 8658 10147 8661
rect 5056 8576 5212 8580
rect 5151 8560 5212 8576
rect 4773 8521 4834 8537
rect 4773 8517 4929 8521
rect 4773 8499 4793 8517
rect 4811 8499 4929 8517
rect 9833 8628 9851 8646
rect 9869 8631 9984 8646
rect 10032 8643 10147 8658
rect 10165 8643 10183 8661
rect 9869 8628 9890 8631
rect 9833 8609 9890 8628
rect 10032 8620 10183 8643
rect 10032 8584 10074 8620
rect 10031 8583 10131 8584
rect 9829 8562 9890 8578
rect 10031 8562 10187 8583
rect 9829 8558 9985 8562
rect 9829 8540 9849 8558
rect 9867 8540 9985 8558
rect 10031 8544 10149 8562
rect 10167 8544 10187 8562
rect 14804 8713 14865 8729
rect 14804 8709 14960 8713
rect 14804 8691 14824 8709
rect 14842 8691 14960 8709
rect 15182 8702 15239 8721
rect 15182 8699 15203 8702
rect 14804 8670 14960 8691
rect 14860 8669 14960 8670
rect 15088 8684 15203 8699
rect 15221 8684 15239 8702
rect 14917 8633 14959 8669
rect 14808 8610 14959 8633
rect 15088 8661 15239 8684
rect 15088 8625 15130 8661
rect 10031 8540 10187 8544
rect 9829 8519 9985 8540
rect 10126 8524 10187 8540
rect 9885 8518 9985 8519
rect 4773 8478 4929 8499
rect 4829 8477 4929 8478
rect 4886 8441 4928 8477
rect 4777 8418 4928 8441
rect 9942 8482 9984 8518
rect 9833 8459 9984 8482
rect 14808 8592 14826 8610
rect 14844 8595 14959 8610
rect 15087 8624 15187 8625
rect 15087 8603 15243 8624
rect 14844 8592 14865 8595
rect 14808 8573 14865 8592
rect 15087 8585 15205 8603
rect 15223 8585 15243 8603
rect 19860 8754 19921 8770
rect 19860 8750 20016 8754
rect 19860 8732 19880 8750
rect 19898 8732 20016 8750
rect 19860 8711 20016 8732
rect 19916 8710 20016 8711
rect 19973 8674 20015 8710
rect 19864 8651 20015 8674
rect 15087 8581 15243 8585
rect 15182 8565 15243 8581
rect 14804 8526 14865 8542
rect 14804 8522 14960 8526
rect 14804 8504 14824 8522
rect 14842 8504 14960 8522
rect 19864 8633 19882 8651
rect 19900 8636 20015 8651
rect 19900 8633 19921 8636
rect 19864 8614 19921 8633
rect 19860 8567 19921 8583
rect 19860 8563 20016 8567
rect 19860 8545 19880 8563
rect 19898 8545 20016 8563
rect 19860 8524 20016 8545
rect 19916 8523 20016 8524
rect 14804 8483 14960 8504
rect 14860 8482 14960 8483
rect 4777 8400 4795 8418
rect 4813 8403 4928 8418
rect 4813 8400 4834 8403
rect 4777 8381 4834 8400
rect 96 8199 153 8218
rect 96 8196 117 8199
rect 2 8181 117 8196
rect 135 8181 153 8199
rect 9833 8441 9851 8459
rect 9869 8444 9984 8459
rect 9869 8441 9890 8444
rect 9833 8422 9890 8441
rect 14917 8446 14959 8482
rect 14808 8423 14959 8446
rect 19973 8487 20015 8523
rect 19864 8464 20015 8487
rect 5152 8240 5209 8259
rect 5152 8237 5173 8240
rect 5058 8222 5173 8237
rect 5191 8222 5209 8240
rect 14808 8405 14826 8423
rect 14844 8408 14959 8423
rect 14844 8405 14865 8408
rect 14808 8386 14865 8405
rect 2 8158 153 8181
rect 2 8122 44 8158
rect 5058 8199 5209 8222
rect 5058 8163 5100 8199
rect 10127 8204 10184 8223
rect 10127 8201 10148 8204
rect 10033 8186 10148 8201
rect 10166 8186 10184 8204
rect 19864 8446 19882 8464
rect 19900 8449 20015 8464
rect 19900 8446 19921 8449
rect 19864 8427 19921 8446
rect 15183 8245 15240 8264
rect 15183 8242 15204 8245
rect 15089 8227 15204 8242
rect 15222 8227 15240 8245
rect 5057 8162 5157 8163
rect 5057 8141 5213 8162
rect 1 8121 101 8122
rect 1 8100 157 8121
rect 1 8082 119 8100
rect 137 8082 157 8100
rect 1 8078 157 8082
rect 96 8062 157 8078
rect 96 8012 153 8031
rect 96 8009 117 8012
rect 2 7994 117 8009
rect 135 7994 153 8012
rect 5057 8123 5175 8141
rect 5193 8123 5213 8141
rect 5057 8119 5213 8123
rect 5152 8103 5213 8119
rect 4774 8064 4835 8080
rect 4774 8060 4930 8064
rect 2 7971 153 7994
rect 2 7935 44 7971
rect 1 7934 101 7935
rect 1 7913 157 7934
rect 1 7895 119 7913
rect 137 7895 157 7913
rect 1 7891 157 7895
rect 96 7875 157 7891
rect 4774 8042 4794 8060
rect 4812 8042 4930 8060
rect 5152 8053 5209 8072
rect 5152 8050 5173 8053
rect 4774 8021 4930 8042
rect 4830 8020 4930 8021
rect 5058 8035 5173 8050
rect 5191 8035 5209 8053
rect 10033 8163 10184 8186
rect 10033 8127 10075 8163
rect 15089 8204 15240 8227
rect 15089 8168 15131 8204
rect 15088 8167 15188 8168
rect 15088 8146 15244 8167
rect 10032 8126 10132 8127
rect 9830 8105 9891 8121
rect 10032 8105 10188 8126
rect 9830 8101 9986 8105
rect 4887 7984 4929 8020
rect 4778 7961 4929 7984
rect 5058 8012 5209 8035
rect 5058 7976 5100 8012
rect 4778 7943 4796 7961
rect 4814 7946 4929 7961
rect 5057 7975 5157 7976
rect 5057 7954 5213 7975
rect 4814 7943 4835 7946
rect 4778 7924 4835 7943
rect 5057 7936 5175 7954
rect 5193 7936 5213 7954
rect 5057 7932 5213 7936
rect 5152 7916 5213 7932
rect 9830 8083 9850 8101
rect 9868 8083 9986 8101
rect 10032 8087 10150 8105
rect 10168 8087 10188 8105
rect 10032 8083 10188 8087
rect 9830 8062 9986 8083
rect 10127 8067 10188 8083
rect 9886 8061 9986 8062
rect 9943 8025 9985 8061
rect 9834 8002 9985 8025
rect 10127 8017 10184 8036
rect 10127 8014 10148 8017
rect 9834 7984 9852 8002
rect 9870 7987 9985 8002
rect 10033 7999 10148 8014
rect 10166 7999 10184 8017
rect 15088 8128 15206 8146
rect 15224 8128 15244 8146
rect 15088 8124 15244 8128
rect 15183 8108 15244 8124
rect 14805 8069 14866 8085
rect 14805 8065 14961 8069
rect 9870 7984 9891 7987
rect 9834 7965 9891 7984
rect 10033 7976 10184 7999
rect 10033 7940 10075 7976
rect 96 7783 153 7802
rect 96 7780 117 7783
rect 2 7765 117 7780
rect 135 7765 153 7783
rect 2 7742 153 7765
rect 4774 7834 4835 7850
rect 4774 7830 4930 7834
rect 2 7706 44 7742
rect 1 7705 101 7706
rect 1 7684 157 7705
rect 1 7666 119 7684
rect 137 7666 157 7684
rect 4774 7812 4794 7830
rect 4812 7812 4930 7830
rect 5152 7824 5209 7843
rect 5152 7821 5173 7824
rect 4774 7791 4930 7812
rect 4830 7790 4930 7791
rect 5058 7806 5173 7821
rect 5191 7806 5209 7824
rect 4887 7754 4929 7790
rect 1 7662 157 7666
rect 96 7646 157 7662
rect 4778 7731 4929 7754
rect 5058 7783 5209 7806
rect 10032 7939 10132 7940
rect 10032 7918 10188 7939
rect 10032 7900 10150 7918
rect 10168 7900 10188 7918
rect 10032 7896 10188 7900
rect 9830 7875 9891 7891
rect 10127 7880 10188 7896
rect 14805 8047 14825 8065
rect 14843 8047 14961 8065
rect 15183 8058 15240 8077
rect 15183 8055 15204 8058
rect 14805 8026 14961 8047
rect 14861 8025 14961 8026
rect 15089 8040 15204 8055
rect 15222 8040 15240 8058
rect 19861 8110 19922 8126
rect 19861 8106 20017 8110
rect 14918 7989 14960 8025
rect 14809 7966 14960 7989
rect 15089 8017 15240 8040
rect 15089 7981 15131 8017
rect 14809 7948 14827 7966
rect 14845 7951 14960 7966
rect 15088 7980 15188 7981
rect 15088 7959 15244 7980
rect 14845 7948 14866 7951
rect 14809 7929 14866 7948
rect 15088 7941 15206 7959
rect 15224 7941 15244 7959
rect 15088 7937 15244 7941
rect 15183 7921 15244 7937
rect 19861 8088 19881 8106
rect 19899 8088 20017 8106
rect 19861 8067 20017 8088
rect 19917 8066 20017 8067
rect 19974 8030 20016 8066
rect 19865 8007 20016 8030
rect 19865 7989 19883 8007
rect 19901 7992 20016 8007
rect 19901 7989 19922 7992
rect 19865 7970 19922 7989
rect 9830 7871 9986 7875
rect 5058 7747 5100 7783
rect 4778 7713 4796 7731
rect 4814 7716 4929 7731
rect 5057 7746 5157 7747
rect 5057 7725 5213 7746
rect 4814 7713 4835 7716
rect 4778 7694 4835 7713
rect 5057 7707 5175 7725
rect 5193 7707 5213 7725
rect 9830 7853 9850 7871
rect 9868 7853 9986 7871
rect 9830 7832 9986 7853
rect 9886 7831 9986 7832
rect 9943 7795 9985 7831
rect 5057 7703 5213 7707
rect 5152 7687 5213 7703
rect 9834 7772 9985 7795
rect 10127 7788 10184 7807
rect 10127 7785 10148 7788
rect 9834 7754 9852 7772
rect 9870 7757 9985 7772
rect 10033 7770 10148 7785
rect 10166 7770 10184 7788
rect 9870 7754 9891 7757
rect 9834 7735 9891 7754
rect 10033 7747 10184 7770
rect 14805 7839 14866 7855
rect 14805 7835 14961 7839
rect 10033 7711 10075 7747
rect 10032 7710 10132 7711
rect 10032 7689 10188 7710
rect 10032 7671 10150 7689
rect 10168 7671 10188 7689
rect 14805 7817 14825 7835
rect 14843 7817 14961 7835
rect 15183 7829 15240 7848
rect 15183 7826 15204 7829
rect 14805 7796 14961 7817
rect 14861 7795 14961 7796
rect 15089 7811 15204 7826
rect 15222 7811 15240 7829
rect 14918 7759 14960 7795
rect 10032 7667 10188 7671
rect 96 7553 153 7572
rect 96 7550 117 7553
rect 2 7535 117 7550
rect 135 7535 153 7553
rect 2 7512 153 7535
rect 2 7476 44 7512
rect 1 7475 101 7476
rect 1 7454 157 7475
rect 1 7436 119 7454
rect 137 7436 157 7454
rect 4774 7605 4835 7621
rect 4774 7601 4930 7605
rect 4774 7583 4794 7601
rect 4812 7583 4930 7601
rect 5152 7594 5209 7613
rect 5152 7591 5173 7594
rect 4774 7562 4930 7583
rect 4830 7561 4930 7562
rect 5058 7576 5173 7591
rect 5191 7576 5209 7594
rect 4887 7525 4929 7561
rect 4778 7502 4929 7525
rect 5058 7553 5209 7576
rect 5058 7517 5100 7553
rect 1 7432 157 7436
rect 96 7416 157 7432
rect 4778 7484 4796 7502
rect 4814 7487 4929 7502
rect 5057 7516 5157 7517
rect 5057 7495 5213 7516
rect 4814 7484 4835 7487
rect 4778 7465 4835 7484
rect 5057 7477 5175 7495
rect 5193 7477 5213 7495
rect 9830 7646 9891 7662
rect 10127 7651 10188 7667
rect 9830 7642 9986 7646
rect 9830 7624 9850 7642
rect 9868 7624 9986 7642
rect 9830 7603 9986 7624
rect 9886 7602 9986 7603
rect 14809 7736 14960 7759
rect 15089 7788 15240 7811
rect 19861 7880 19922 7896
rect 19861 7876 20017 7880
rect 15089 7752 15131 7788
rect 14809 7718 14827 7736
rect 14845 7721 14960 7736
rect 15088 7751 15188 7752
rect 15088 7730 15244 7751
rect 14845 7718 14866 7721
rect 14809 7699 14866 7718
rect 15088 7712 15206 7730
rect 15224 7712 15244 7730
rect 19861 7858 19881 7876
rect 19899 7858 20017 7876
rect 19861 7837 20017 7858
rect 19917 7836 20017 7837
rect 19974 7800 20016 7836
rect 15088 7708 15244 7712
rect 15183 7692 15244 7708
rect 19865 7777 20016 7800
rect 19865 7759 19883 7777
rect 19901 7762 20016 7777
rect 19901 7759 19922 7762
rect 19865 7740 19922 7759
rect 9943 7566 9985 7602
rect 9834 7543 9985 7566
rect 10127 7558 10184 7577
rect 10127 7555 10148 7558
rect 5057 7473 5213 7477
rect 5152 7457 5213 7473
rect 4774 7418 4835 7434
rect 4774 7414 4930 7418
rect 4774 7396 4794 7414
rect 4812 7396 4930 7414
rect 9834 7525 9852 7543
rect 9870 7528 9985 7543
rect 10033 7540 10148 7555
rect 10166 7540 10184 7558
rect 9870 7525 9891 7528
rect 9834 7506 9891 7525
rect 10033 7517 10184 7540
rect 10033 7481 10075 7517
rect 10032 7480 10132 7481
rect 9830 7459 9891 7475
rect 10032 7459 10188 7480
rect 9830 7455 9986 7459
rect 9830 7437 9850 7455
rect 9868 7437 9986 7455
rect 10032 7441 10150 7459
rect 10168 7441 10188 7459
rect 14805 7610 14866 7626
rect 14805 7606 14961 7610
rect 14805 7588 14825 7606
rect 14843 7588 14961 7606
rect 15183 7599 15240 7618
rect 15183 7596 15204 7599
rect 14805 7567 14961 7588
rect 14861 7566 14961 7567
rect 15089 7581 15204 7596
rect 15222 7581 15240 7599
rect 14918 7530 14960 7566
rect 14809 7507 14960 7530
rect 15089 7558 15240 7581
rect 15089 7522 15131 7558
rect 10032 7437 10188 7441
rect 9830 7416 9986 7437
rect 10127 7421 10188 7437
rect 9886 7415 9986 7416
rect 4774 7375 4930 7396
rect 4830 7374 4930 7375
rect 4887 7338 4929 7374
rect 4778 7315 4929 7338
rect 4778 7297 4796 7315
rect 4814 7300 4929 7315
rect 9943 7379 9985 7415
rect 9834 7356 9985 7379
rect 14809 7489 14827 7507
rect 14845 7492 14960 7507
rect 15088 7521 15188 7522
rect 15088 7500 15244 7521
rect 14845 7489 14866 7492
rect 14809 7470 14866 7489
rect 15088 7482 15206 7500
rect 15224 7482 15244 7500
rect 19861 7651 19922 7667
rect 19861 7647 20017 7651
rect 19861 7629 19881 7647
rect 19899 7629 20017 7647
rect 19861 7608 20017 7629
rect 19917 7607 20017 7608
rect 19974 7571 20016 7607
rect 19865 7548 20016 7571
rect 15088 7478 15244 7482
rect 15183 7462 15244 7478
rect 14805 7423 14866 7439
rect 14805 7419 14961 7423
rect 14805 7401 14825 7419
rect 14843 7401 14961 7419
rect 19865 7530 19883 7548
rect 19901 7533 20016 7548
rect 19901 7530 19922 7533
rect 19865 7511 19922 7530
rect 19861 7464 19922 7480
rect 19861 7460 20017 7464
rect 19861 7442 19881 7460
rect 19899 7442 20017 7460
rect 19861 7421 20017 7442
rect 19917 7420 20017 7421
rect 14805 7380 14961 7401
rect 14861 7379 14961 7380
rect 9834 7338 9852 7356
rect 9870 7341 9985 7356
rect 9870 7338 9891 7341
rect 4814 7297 4835 7300
rect 4778 7278 4835 7297
rect 9834 7319 9891 7338
rect 14918 7343 14960 7379
rect 14809 7320 14960 7343
rect 14809 7302 14827 7320
rect 14845 7305 14960 7320
rect 19974 7384 20016 7420
rect 19865 7361 20016 7384
rect 19865 7343 19883 7361
rect 19901 7346 20016 7361
rect 19901 7343 19922 7346
rect 14845 7302 14866 7305
rect 96 7096 153 7115
rect 5152 7137 5209 7156
rect 14809 7283 14866 7302
rect 19865 7324 19922 7343
rect 5152 7134 5173 7137
rect 96 7093 117 7096
rect 2 7078 117 7093
rect 135 7078 153 7096
rect 2 7055 153 7078
rect 2 7019 44 7055
rect 5058 7119 5173 7134
rect 5191 7119 5209 7137
rect 5058 7096 5209 7119
rect 5058 7060 5100 7096
rect 10127 7101 10184 7120
rect 15183 7142 15240 7161
rect 15183 7139 15204 7142
rect 10127 7098 10148 7101
rect 10033 7083 10148 7098
rect 10166 7083 10184 7101
rect 5057 7059 5157 7060
rect 5057 7038 5213 7059
rect 1 7018 101 7019
rect 1 6997 157 7018
rect 1 6979 119 6997
rect 137 6979 157 6997
rect 1 6975 157 6979
rect 96 6959 157 6975
rect 96 6909 153 6928
rect 96 6906 117 6909
rect 2 6891 117 6906
rect 135 6891 153 6909
rect 5057 7020 5175 7038
rect 5193 7020 5213 7038
rect 5057 7016 5213 7020
rect 5152 7000 5213 7016
rect 4774 6961 4835 6977
rect 4774 6957 4930 6961
rect 2 6868 153 6891
rect 2 6832 44 6868
rect 1 6831 101 6832
rect 1 6810 157 6831
rect 1 6792 119 6810
rect 137 6792 157 6810
rect 1 6788 157 6792
rect 96 6772 157 6788
rect 4774 6939 4794 6957
rect 4812 6939 4930 6957
rect 5152 6950 5209 6969
rect 5152 6947 5173 6950
rect 4774 6918 4930 6939
rect 4830 6917 4930 6918
rect 5058 6932 5173 6947
rect 5191 6932 5209 6950
rect 10033 7060 10184 7083
rect 10033 7024 10075 7060
rect 15089 7124 15204 7139
rect 15222 7124 15240 7142
rect 15089 7101 15240 7124
rect 15089 7065 15131 7101
rect 15088 7064 15188 7065
rect 15088 7043 15244 7064
rect 10032 7023 10132 7024
rect 9830 7002 9891 7018
rect 10032 7002 10188 7023
rect 9830 6998 9986 7002
rect 4887 6881 4929 6917
rect 4778 6858 4929 6881
rect 5058 6909 5209 6932
rect 5058 6873 5100 6909
rect 4778 6840 4796 6858
rect 4814 6843 4929 6858
rect 5057 6872 5157 6873
rect 5057 6851 5213 6872
rect 4814 6840 4835 6843
rect 4778 6821 4835 6840
rect 5057 6833 5175 6851
rect 5193 6833 5213 6851
rect 5057 6829 5213 6833
rect 5152 6813 5213 6829
rect 9830 6980 9850 6998
rect 9868 6980 9986 6998
rect 10032 6984 10150 7002
rect 10168 6984 10188 7002
rect 10032 6980 10188 6984
rect 9830 6959 9986 6980
rect 10127 6964 10188 6980
rect 9886 6958 9986 6959
rect 9943 6922 9985 6958
rect 9834 6899 9985 6922
rect 10127 6914 10184 6933
rect 10127 6911 10148 6914
rect 9834 6881 9852 6899
rect 9870 6884 9985 6899
rect 10033 6896 10148 6911
rect 10166 6896 10184 6914
rect 15088 7025 15206 7043
rect 15224 7025 15244 7043
rect 15088 7021 15244 7025
rect 15183 7005 15244 7021
rect 14805 6966 14866 6982
rect 14805 6962 14961 6966
rect 9870 6881 9891 6884
rect 9834 6862 9891 6881
rect 10033 6873 10184 6896
rect 10033 6837 10075 6873
rect 96 6680 153 6699
rect 96 6677 117 6680
rect 2 6662 117 6677
rect 135 6662 153 6680
rect 2 6639 153 6662
rect 4774 6731 4835 6747
rect 4774 6727 4930 6731
rect 2 6603 44 6639
rect 1 6602 101 6603
rect 1 6581 157 6602
rect 1 6563 119 6581
rect 137 6563 157 6581
rect 4774 6709 4794 6727
rect 4812 6709 4930 6727
rect 5152 6721 5209 6740
rect 5152 6718 5173 6721
rect 4774 6688 4930 6709
rect 4830 6687 4930 6688
rect 5058 6703 5173 6718
rect 5191 6703 5209 6721
rect 4887 6651 4929 6687
rect 1 6559 157 6563
rect 96 6543 157 6559
rect 4778 6628 4929 6651
rect 5058 6680 5209 6703
rect 10032 6836 10132 6837
rect 10032 6815 10188 6836
rect 10032 6797 10150 6815
rect 10168 6797 10188 6815
rect 10032 6793 10188 6797
rect 9830 6772 9891 6788
rect 10127 6777 10188 6793
rect 14805 6944 14825 6962
rect 14843 6944 14961 6962
rect 15183 6955 15240 6974
rect 15183 6952 15204 6955
rect 14805 6923 14961 6944
rect 14861 6922 14961 6923
rect 15089 6937 15204 6952
rect 15222 6937 15240 6955
rect 19861 7007 19922 7023
rect 19861 7003 20017 7007
rect 14918 6886 14960 6922
rect 14809 6863 14960 6886
rect 15089 6914 15240 6937
rect 15089 6878 15131 6914
rect 14809 6845 14827 6863
rect 14845 6848 14960 6863
rect 15088 6877 15188 6878
rect 15088 6856 15244 6877
rect 14845 6845 14866 6848
rect 14809 6826 14866 6845
rect 15088 6838 15206 6856
rect 15224 6838 15244 6856
rect 15088 6834 15244 6838
rect 15183 6818 15244 6834
rect 19861 6985 19881 7003
rect 19899 6985 20017 7003
rect 19861 6964 20017 6985
rect 19917 6963 20017 6964
rect 19974 6927 20016 6963
rect 19865 6904 20016 6927
rect 19865 6886 19883 6904
rect 19901 6889 20016 6904
rect 19901 6886 19922 6889
rect 19865 6867 19922 6886
rect 9830 6768 9986 6772
rect 5058 6644 5100 6680
rect 4778 6610 4796 6628
rect 4814 6613 4929 6628
rect 5057 6643 5157 6644
rect 5057 6622 5213 6643
rect 4814 6610 4835 6613
rect 4778 6591 4835 6610
rect 5057 6604 5175 6622
rect 5193 6604 5213 6622
rect 9830 6750 9850 6768
rect 9868 6750 9986 6768
rect 9830 6729 9986 6750
rect 9886 6728 9986 6729
rect 9943 6692 9985 6728
rect 5057 6600 5213 6604
rect 5152 6584 5213 6600
rect 9834 6669 9985 6692
rect 10127 6685 10184 6704
rect 10127 6682 10148 6685
rect 9834 6651 9852 6669
rect 9870 6654 9985 6669
rect 10033 6667 10148 6682
rect 10166 6667 10184 6685
rect 9870 6651 9891 6654
rect 9834 6632 9891 6651
rect 10033 6644 10184 6667
rect 14805 6736 14866 6752
rect 14805 6732 14961 6736
rect 10033 6608 10075 6644
rect 10032 6607 10132 6608
rect 10032 6586 10188 6607
rect 10032 6568 10150 6586
rect 10168 6568 10188 6586
rect 14805 6714 14825 6732
rect 14843 6714 14961 6732
rect 15183 6726 15240 6745
rect 15183 6723 15204 6726
rect 14805 6693 14961 6714
rect 14861 6692 14961 6693
rect 15089 6708 15204 6723
rect 15222 6708 15240 6726
rect 14918 6656 14960 6692
rect 10032 6564 10188 6568
rect 96 6450 153 6469
rect 96 6447 117 6450
rect 2 6432 117 6447
rect 135 6432 153 6450
rect 2 6409 153 6432
rect 2 6373 44 6409
rect 1 6372 101 6373
rect 1 6351 157 6372
rect 1 6333 119 6351
rect 137 6333 157 6351
rect 4774 6502 4835 6518
rect 4774 6498 4930 6502
rect 4774 6480 4794 6498
rect 4812 6480 4930 6498
rect 5152 6491 5209 6510
rect 5152 6488 5173 6491
rect 4774 6459 4930 6480
rect 4830 6458 4930 6459
rect 5058 6473 5173 6488
rect 5191 6473 5209 6491
rect 4887 6422 4929 6458
rect 4778 6399 4929 6422
rect 5058 6450 5209 6473
rect 5058 6414 5100 6450
rect 1 6329 157 6333
rect 96 6313 157 6329
rect 4778 6381 4796 6399
rect 4814 6384 4929 6399
rect 5057 6413 5157 6414
rect 5057 6392 5213 6413
rect 4814 6381 4835 6384
rect 4778 6362 4835 6381
rect 5057 6374 5175 6392
rect 5193 6374 5213 6392
rect 9830 6543 9891 6559
rect 10127 6548 10188 6564
rect 9830 6539 9986 6543
rect 9830 6521 9850 6539
rect 9868 6521 9986 6539
rect 9830 6500 9986 6521
rect 9886 6499 9986 6500
rect 14809 6633 14960 6656
rect 15089 6685 15240 6708
rect 19861 6777 19922 6793
rect 19861 6773 20017 6777
rect 15089 6649 15131 6685
rect 14809 6615 14827 6633
rect 14845 6618 14960 6633
rect 15088 6648 15188 6649
rect 15088 6627 15244 6648
rect 14845 6615 14866 6618
rect 14809 6596 14866 6615
rect 15088 6609 15206 6627
rect 15224 6609 15244 6627
rect 19861 6755 19881 6773
rect 19899 6755 20017 6773
rect 19861 6734 20017 6755
rect 19917 6733 20017 6734
rect 19974 6697 20016 6733
rect 15088 6605 15244 6609
rect 15183 6589 15244 6605
rect 19865 6674 20016 6697
rect 19865 6656 19883 6674
rect 19901 6659 20016 6674
rect 19901 6656 19922 6659
rect 19865 6637 19922 6656
rect 9943 6463 9985 6499
rect 9834 6440 9985 6463
rect 10127 6455 10184 6474
rect 10127 6452 10148 6455
rect 5057 6370 5213 6374
rect 5152 6354 5213 6370
rect 4774 6315 4835 6331
rect 4774 6311 4930 6315
rect 4774 6293 4794 6311
rect 4812 6293 4930 6311
rect 9834 6422 9852 6440
rect 9870 6425 9985 6440
rect 10033 6437 10148 6452
rect 10166 6437 10184 6455
rect 9870 6422 9891 6425
rect 9834 6403 9891 6422
rect 10033 6414 10184 6437
rect 10033 6378 10075 6414
rect 10032 6377 10132 6378
rect 9830 6356 9891 6372
rect 10032 6356 10188 6377
rect 9830 6352 9986 6356
rect 9830 6334 9850 6352
rect 9868 6334 9986 6352
rect 10032 6338 10150 6356
rect 10168 6338 10188 6356
rect 14805 6507 14866 6523
rect 14805 6503 14961 6507
rect 14805 6485 14825 6503
rect 14843 6485 14961 6503
rect 15183 6496 15240 6515
rect 15183 6493 15204 6496
rect 14805 6464 14961 6485
rect 14861 6463 14961 6464
rect 15089 6478 15204 6493
rect 15222 6478 15240 6496
rect 14918 6427 14960 6463
rect 14809 6404 14960 6427
rect 15089 6455 15240 6478
rect 15089 6419 15131 6455
rect 10032 6334 10188 6338
rect 9830 6313 9986 6334
rect 10127 6318 10188 6334
rect 9886 6312 9986 6313
rect 4774 6272 4930 6293
rect 4830 6271 4930 6272
rect 4887 6235 4929 6271
rect 4778 6212 4929 6235
rect 9943 6276 9985 6312
rect 9834 6253 9985 6276
rect 14809 6386 14827 6404
rect 14845 6389 14960 6404
rect 15088 6418 15188 6419
rect 15088 6397 15244 6418
rect 14845 6386 14866 6389
rect 14809 6367 14866 6386
rect 15088 6379 15206 6397
rect 15224 6379 15244 6397
rect 19861 6548 19922 6564
rect 19861 6544 20017 6548
rect 19861 6526 19881 6544
rect 19899 6526 20017 6544
rect 19861 6505 20017 6526
rect 19917 6504 20017 6505
rect 19974 6468 20016 6504
rect 19865 6445 20016 6468
rect 15088 6375 15244 6379
rect 15183 6359 15244 6375
rect 14805 6320 14866 6336
rect 14805 6316 14961 6320
rect 14805 6298 14825 6316
rect 14843 6298 14961 6316
rect 19865 6427 19883 6445
rect 19901 6430 20016 6445
rect 19901 6427 19922 6430
rect 19865 6408 19922 6427
rect 19861 6361 19922 6377
rect 19861 6357 20017 6361
rect 19861 6339 19881 6357
rect 19899 6339 20017 6357
rect 19861 6318 20017 6339
rect 19917 6317 20017 6318
rect 14805 6277 14961 6298
rect 14861 6276 14961 6277
rect 4778 6194 4796 6212
rect 4814 6197 4929 6212
rect 4814 6194 4835 6197
rect 4778 6175 4835 6194
rect 97 5993 154 6012
rect 97 5990 118 5993
rect 3 5975 118 5990
rect 136 5975 154 5993
rect 9834 6235 9852 6253
rect 9870 6238 9985 6253
rect 9870 6235 9891 6238
rect 9834 6216 9891 6235
rect 14918 6240 14960 6276
rect 14809 6217 14960 6240
rect 19974 6281 20016 6317
rect 19865 6258 20016 6281
rect 5153 6034 5210 6053
rect 5153 6031 5174 6034
rect 5059 6016 5174 6031
rect 5192 6016 5210 6034
rect 14809 6199 14827 6217
rect 14845 6202 14960 6217
rect 14845 6199 14866 6202
rect 14809 6180 14866 6199
rect 3 5952 154 5975
rect 3 5916 45 5952
rect 5059 5993 5210 6016
rect 5059 5957 5101 5993
rect 10128 5998 10185 6017
rect 10128 5995 10149 5998
rect 10034 5980 10149 5995
rect 10167 5980 10185 5998
rect 19865 6240 19883 6258
rect 19901 6243 20016 6258
rect 19901 6240 19922 6243
rect 19865 6221 19922 6240
rect 15184 6039 15241 6058
rect 15184 6036 15205 6039
rect 15090 6021 15205 6036
rect 15223 6021 15241 6039
rect 5058 5956 5158 5957
rect 5058 5935 5214 5956
rect 2 5915 102 5916
rect 2 5894 158 5915
rect 2 5876 120 5894
rect 138 5876 158 5894
rect 2 5872 158 5876
rect 97 5856 158 5872
rect 97 5806 154 5825
rect 97 5803 118 5806
rect 3 5788 118 5803
rect 136 5788 154 5806
rect 5058 5917 5176 5935
rect 5194 5917 5214 5935
rect 5058 5913 5214 5917
rect 5153 5897 5214 5913
rect 4775 5858 4836 5874
rect 4775 5854 4931 5858
rect 3 5765 154 5788
rect 3 5729 45 5765
rect 2 5728 102 5729
rect 2 5707 158 5728
rect 2 5689 120 5707
rect 138 5689 158 5707
rect 2 5685 158 5689
rect 97 5669 158 5685
rect 4775 5836 4795 5854
rect 4813 5836 4931 5854
rect 5153 5847 5210 5866
rect 5153 5844 5174 5847
rect 4775 5815 4931 5836
rect 4831 5814 4931 5815
rect 5059 5829 5174 5844
rect 5192 5829 5210 5847
rect 10034 5957 10185 5980
rect 10034 5921 10076 5957
rect 15090 5998 15241 6021
rect 15090 5962 15132 5998
rect 15089 5961 15189 5962
rect 15089 5940 15245 5961
rect 10033 5920 10133 5921
rect 9831 5899 9892 5915
rect 10033 5899 10189 5920
rect 9831 5895 9987 5899
rect 4888 5778 4930 5814
rect 4779 5755 4930 5778
rect 5059 5806 5210 5829
rect 5059 5770 5101 5806
rect 4779 5737 4797 5755
rect 4815 5740 4930 5755
rect 5058 5769 5158 5770
rect 5058 5748 5214 5769
rect 4815 5737 4836 5740
rect 4779 5718 4836 5737
rect 5058 5730 5176 5748
rect 5194 5730 5214 5748
rect 5058 5726 5214 5730
rect 5153 5710 5214 5726
rect 9831 5877 9851 5895
rect 9869 5877 9987 5895
rect 10033 5881 10151 5899
rect 10169 5881 10189 5899
rect 10033 5877 10189 5881
rect 9831 5856 9987 5877
rect 10128 5861 10189 5877
rect 9887 5855 9987 5856
rect 9944 5819 9986 5855
rect 9835 5796 9986 5819
rect 10128 5811 10185 5830
rect 10128 5808 10149 5811
rect 9835 5778 9853 5796
rect 9871 5781 9986 5796
rect 10034 5793 10149 5808
rect 10167 5793 10185 5811
rect 15089 5922 15207 5940
rect 15225 5922 15245 5940
rect 15089 5918 15245 5922
rect 15184 5902 15245 5918
rect 14806 5863 14867 5879
rect 14806 5859 14962 5863
rect 9871 5778 9892 5781
rect 9835 5759 9892 5778
rect 10034 5770 10185 5793
rect 10034 5734 10076 5770
rect 97 5577 154 5596
rect 97 5574 118 5577
rect 3 5559 118 5574
rect 136 5559 154 5577
rect 3 5536 154 5559
rect 4775 5628 4836 5644
rect 4775 5624 4931 5628
rect 3 5500 45 5536
rect 2 5499 102 5500
rect 2 5478 158 5499
rect 2 5460 120 5478
rect 138 5460 158 5478
rect 4775 5606 4795 5624
rect 4813 5606 4931 5624
rect 5153 5618 5210 5637
rect 5153 5615 5174 5618
rect 4775 5585 4931 5606
rect 4831 5584 4931 5585
rect 5059 5600 5174 5615
rect 5192 5600 5210 5618
rect 4888 5548 4930 5584
rect 2 5456 158 5460
rect 97 5440 158 5456
rect 4779 5525 4930 5548
rect 5059 5577 5210 5600
rect 10033 5733 10133 5734
rect 10033 5712 10189 5733
rect 10033 5694 10151 5712
rect 10169 5694 10189 5712
rect 10033 5690 10189 5694
rect 9831 5669 9892 5685
rect 10128 5674 10189 5690
rect 14806 5841 14826 5859
rect 14844 5841 14962 5859
rect 15184 5852 15241 5871
rect 15184 5849 15205 5852
rect 14806 5820 14962 5841
rect 14862 5819 14962 5820
rect 15090 5834 15205 5849
rect 15223 5834 15241 5852
rect 19862 5904 19923 5920
rect 19862 5900 20018 5904
rect 14919 5783 14961 5819
rect 14810 5760 14961 5783
rect 15090 5811 15241 5834
rect 15090 5775 15132 5811
rect 14810 5742 14828 5760
rect 14846 5745 14961 5760
rect 15089 5774 15189 5775
rect 15089 5753 15245 5774
rect 14846 5742 14867 5745
rect 14810 5723 14867 5742
rect 15089 5735 15207 5753
rect 15225 5735 15245 5753
rect 15089 5731 15245 5735
rect 15184 5715 15245 5731
rect 19862 5882 19882 5900
rect 19900 5882 20018 5900
rect 19862 5861 20018 5882
rect 19918 5860 20018 5861
rect 19975 5824 20017 5860
rect 19866 5801 20017 5824
rect 19866 5783 19884 5801
rect 19902 5786 20017 5801
rect 19902 5783 19923 5786
rect 19866 5764 19923 5783
rect 9831 5665 9987 5669
rect 5059 5541 5101 5577
rect 4779 5507 4797 5525
rect 4815 5510 4930 5525
rect 5058 5540 5158 5541
rect 5058 5519 5214 5540
rect 4815 5507 4836 5510
rect 4779 5488 4836 5507
rect 5058 5501 5176 5519
rect 5194 5501 5214 5519
rect 9831 5647 9851 5665
rect 9869 5647 9987 5665
rect 9831 5626 9987 5647
rect 9887 5625 9987 5626
rect 9944 5589 9986 5625
rect 5058 5497 5214 5501
rect 5153 5481 5214 5497
rect 9835 5566 9986 5589
rect 10128 5582 10185 5601
rect 10128 5579 10149 5582
rect 9835 5548 9853 5566
rect 9871 5551 9986 5566
rect 10034 5564 10149 5579
rect 10167 5564 10185 5582
rect 9871 5548 9892 5551
rect 9835 5529 9892 5548
rect 10034 5541 10185 5564
rect 14806 5633 14867 5649
rect 14806 5629 14962 5633
rect 10034 5505 10076 5541
rect 10033 5504 10133 5505
rect 10033 5483 10189 5504
rect 10033 5465 10151 5483
rect 10169 5465 10189 5483
rect 14806 5611 14826 5629
rect 14844 5611 14962 5629
rect 15184 5623 15241 5642
rect 15184 5620 15205 5623
rect 14806 5590 14962 5611
rect 14862 5589 14962 5590
rect 15090 5605 15205 5620
rect 15223 5605 15241 5623
rect 14919 5553 14961 5589
rect 10033 5461 10189 5465
rect 97 5347 154 5366
rect 97 5344 118 5347
rect 3 5329 118 5344
rect 136 5329 154 5347
rect 3 5306 154 5329
rect 3 5270 45 5306
rect 2 5269 102 5270
rect 2 5248 158 5269
rect 2 5230 120 5248
rect 138 5230 158 5248
rect 4775 5399 4836 5415
rect 4775 5395 4931 5399
rect 4775 5377 4795 5395
rect 4813 5377 4931 5395
rect 5153 5388 5210 5407
rect 5153 5385 5174 5388
rect 4775 5356 4931 5377
rect 4831 5355 4931 5356
rect 5059 5370 5174 5385
rect 5192 5370 5210 5388
rect 4888 5319 4930 5355
rect 4779 5296 4930 5319
rect 5059 5347 5210 5370
rect 5059 5311 5101 5347
rect 2 5226 158 5230
rect 97 5210 158 5226
rect 4779 5278 4797 5296
rect 4815 5281 4930 5296
rect 5058 5310 5158 5311
rect 5058 5289 5214 5310
rect 4815 5278 4836 5281
rect 4779 5259 4836 5278
rect 5058 5271 5176 5289
rect 5194 5271 5214 5289
rect 9831 5440 9892 5456
rect 10128 5445 10189 5461
rect 9831 5436 9987 5440
rect 9831 5418 9851 5436
rect 9869 5418 9987 5436
rect 9831 5397 9987 5418
rect 9887 5396 9987 5397
rect 14810 5530 14961 5553
rect 15090 5582 15241 5605
rect 19862 5674 19923 5690
rect 19862 5670 20018 5674
rect 15090 5546 15132 5582
rect 14810 5512 14828 5530
rect 14846 5515 14961 5530
rect 15089 5545 15189 5546
rect 15089 5524 15245 5545
rect 14846 5512 14867 5515
rect 14810 5493 14867 5512
rect 15089 5506 15207 5524
rect 15225 5506 15245 5524
rect 19862 5652 19882 5670
rect 19900 5652 20018 5670
rect 19862 5631 20018 5652
rect 19918 5630 20018 5631
rect 19975 5594 20017 5630
rect 15089 5502 15245 5506
rect 15184 5486 15245 5502
rect 19866 5571 20017 5594
rect 19866 5553 19884 5571
rect 19902 5556 20017 5571
rect 19902 5553 19923 5556
rect 19866 5534 19923 5553
rect 9944 5360 9986 5396
rect 9835 5337 9986 5360
rect 10128 5352 10185 5371
rect 10128 5349 10149 5352
rect 5058 5267 5214 5271
rect 5153 5251 5214 5267
rect 4775 5212 4836 5228
rect 4775 5208 4931 5212
rect 4775 5190 4795 5208
rect 4813 5190 4931 5208
rect 9835 5319 9853 5337
rect 9871 5322 9986 5337
rect 10034 5334 10149 5349
rect 10167 5334 10185 5352
rect 9871 5319 9892 5322
rect 9835 5300 9892 5319
rect 10034 5311 10185 5334
rect 10034 5275 10076 5311
rect 10033 5274 10133 5275
rect 9831 5253 9892 5269
rect 10033 5253 10189 5274
rect 9831 5249 9987 5253
rect 9831 5231 9851 5249
rect 9869 5231 9987 5249
rect 10033 5235 10151 5253
rect 10169 5235 10189 5253
rect 14806 5404 14867 5420
rect 14806 5400 14962 5404
rect 14806 5382 14826 5400
rect 14844 5382 14962 5400
rect 15184 5393 15241 5412
rect 15184 5390 15205 5393
rect 14806 5361 14962 5382
rect 14862 5360 14962 5361
rect 15090 5375 15205 5390
rect 15223 5375 15241 5393
rect 14919 5324 14961 5360
rect 14810 5301 14961 5324
rect 15090 5352 15241 5375
rect 15090 5316 15132 5352
rect 10033 5231 10189 5235
rect 4775 5169 4931 5190
rect 4831 5168 4931 5169
rect 4888 5132 4930 5168
rect 9831 5210 9987 5231
rect 10128 5215 10189 5231
rect 9887 5209 9987 5210
rect 4779 5109 4930 5132
rect 4779 5091 4797 5109
rect 4815 5094 4930 5109
rect 4815 5091 4836 5094
rect 4779 5072 4836 5091
rect 9944 5173 9986 5209
rect 9835 5150 9986 5173
rect 14810 5283 14828 5301
rect 14846 5286 14961 5301
rect 15089 5315 15189 5316
rect 15089 5294 15245 5315
rect 14846 5283 14867 5286
rect 14810 5264 14867 5283
rect 15089 5276 15207 5294
rect 15225 5276 15245 5294
rect 19862 5445 19923 5461
rect 19862 5441 20018 5445
rect 19862 5423 19882 5441
rect 19900 5423 20018 5441
rect 19862 5402 20018 5423
rect 19918 5401 20018 5402
rect 19975 5365 20017 5401
rect 19866 5342 20017 5365
rect 15089 5272 15245 5276
rect 15184 5256 15245 5272
rect 14806 5217 14867 5233
rect 14806 5213 14962 5217
rect 14806 5195 14826 5213
rect 14844 5195 14962 5213
rect 19866 5324 19884 5342
rect 19902 5327 20017 5342
rect 19902 5324 19923 5327
rect 19866 5305 19923 5324
rect 19862 5258 19923 5274
rect 19862 5254 20018 5258
rect 19862 5236 19882 5254
rect 19900 5236 20018 5254
rect 9835 5132 9853 5150
rect 9871 5135 9986 5150
rect 9871 5132 9892 5135
rect 9835 5113 9892 5132
rect 14806 5174 14962 5195
rect 14862 5173 14962 5174
rect 97 4890 154 4909
rect 97 4887 118 4890
rect 3 4872 118 4887
rect 136 4872 154 4890
rect 3 4849 154 4872
rect 3 4813 45 4849
rect 5153 4931 5210 4950
rect 5153 4928 5174 4931
rect 5059 4913 5174 4928
rect 5192 4913 5210 4931
rect 5059 4890 5210 4913
rect 2 4812 102 4813
rect 2 4791 158 4812
rect 5059 4854 5101 4890
rect 14919 5137 14961 5173
rect 19862 5215 20018 5236
rect 19918 5214 20018 5215
rect 14810 5114 14961 5137
rect 14810 5096 14828 5114
rect 14846 5099 14961 5114
rect 14846 5096 14867 5099
rect 14810 5077 14867 5096
rect 19975 5178 20017 5214
rect 19866 5155 20017 5178
rect 19866 5137 19884 5155
rect 19902 5140 20017 5155
rect 19902 5137 19923 5140
rect 19866 5118 19923 5137
rect 5058 4853 5158 4854
rect 5058 4832 5214 4853
rect 10128 4895 10185 4914
rect 10128 4892 10149 4895
rect 10034 4877 10149 4892
rect 10167 4877 10185 4895
rect 2 4773 120 4791
rect 138 4773 158 4791
rect 2 4769 158 4773
rect 97 4753 158 4769
rect 97 4703 154 4722
rect 97 4700 118 4703
rect 3 4685 118 4700
rect 136 4685 154 4703
rect 5058 4814 5176 4832
rect 5194 4814 5214 4832
rect 5058 4810 5214 4814
rect 5153 4794 5214 4810
rect 4775 4755 4836 4771
rect 4775 4751 4931 4755
rect 3 4662 154 4685
rect 3 4626 45 4662
rect 2 4625 102 4626
rect 2 4604 158 4625
rect 2 4586 120 4604
rect 138 4586 158 4604
rect 2 4582 158 4586
rect 97 4566 158 4582
rect 4775 4733 4795 4751
rect 4813 4733 4931 4751
rect 5153 4744 5210 4763
rect 5153 4741 5174 4744
rect 4775 4712 4931 4733
rect 4831 4711 4931 4712
rect 5059 4726 5174 4741
rect 5192 4726 5210 4744
rect 10034 4854 10185 4877
rect 10034 4818 10076 4854
rect 15184 4936 15241 4955
rect 15184 4933 15205 4936
rect 15090 4918 15205 4933
rect 15223 4918 15241 4936
rect 15090 4895 15241 4918
rect 10033 4817 10133 4818
rect 9831 4796 9892 4812
rect 10033 4796 10189 4817
rect 15090 4859 15132 4895
rect 15089 4858 15189 4859
rect 15089 4837 15245 4858
rect 9831 4792 9987 4796
rect 4888 4675 4930 4711
rect 4779 4652 4930 4675
rect 5059 4703 5210 4726
rect 5059 4667 5101 4703
rect 4779 4634 4797 4652
rect 4815 4637 4930 4652
rect 5058 4666 5158 4667
rect 5058 4645 5214 4666
rect 4815 4634 4836 4637
rect 4779 4615 4836 4634
rect 5058 4627 5176 4645
rect 5194 4627 5214 4645
rect 5058 4623 5214 4627
rect 5153 4607 5214 4623
rect 9831 4774 9851 4792
rect 9869 4774 9987 4792
rect 10033 4778 10151 4796
rect 10169 4778 10189 4796
rect 10033 4774 10189 4778
rect 9831 4753 9987 4774
rect 10128 4758 10189 4774
rect 9887 4752 9987 4753
rect 9944 4716 9986 4752
rect 9835 4693 9986 4716
rect 10128 4708 10185 4727
rect 10128 4705 10149 4708
rect 9835 4675 9853 4693
rect 9871 4678 9986 4693
rect 10034 4690 10149 4705
rect 10167 4690 10185 4708
rect 15089 4819 15207 4837
rect 15225 4819 15245 4837
rect 15089 4815 15245 4819
rect 15184 4799 15245 4815
rect 14806 4760 14867 4776
rect 14806 4756 14962 4760
rect 9871 4675 9892 4678
rect 9835 4656 9892 4675
rect 10034 4667 10185 4690
rect 10034 4631 10076 4667
rect 97 4474 154 4493
rect 97 4471 118 4474
rect 3 4456 118 4471
rect 136 4456 154 4474
rect 3 4433 154 4456
rect 4775 4525 4836 4541
rect 4775 4521 4931 4525
rect 3 4397 45 4433
rect 2 4396 102 4397
rect 2 4375 158 4396
rect 2 4357 120 4375
rect 138 4357 158 4375
rect 4775 4503 4795 4521
rect 4813 4503 4931 4521
rect 5153 4515 5210 4534
rect 5153 4512 5174 4515
rect 4775 4482 4931 4503
rect 4831 4481 4931 4482
rect 5059 4497 5174 4512
rect 5192 4497 5210 4515
rect 4888 4445 4930 4481
rect 2 4353 158 4357
rect 97 4337 158 4353
rect 4779 4422 4930 4445
rect 5059 4474 5210 4497
rect 10033 4630 10133 4631
rect 10033 4609 10189 4630
rect 10033 4591 10151 4609
rect 10169 4591 10189 4609
rect 10033 4587 10189 4591
rect 9831 4566 9892 4582
rect 10128 4571 10189 4587
rect 14806 4738 14826 4756
rect 14844 4738 14962 4756
rect 15184 4749 15241 4768
rect 15184 4746 15205 4749
rect 14806 4717 14962 4738
rect 14862 4716 14962 4717
rect 15090 4731 15205 4746
rect 15223 4731 15241 4749
rect 19862 4801 19923 4817
rect 19862 4797 20018 4801
rect 14919 4680 14961 4716
rect 14810 4657 14961 4680
rect 15090 4708 15241 4731
rect 15090 4672 15132 4708
rect 14810 4639 14828 4657
rect 14846 4642 14961 4657
rect 15089 4671 15189 4672
rect 15089 4650 15245 4671
rect 14846 4639 14867 4642
rect 14810 4620 14867 4639
rect 15089 4632 15207 4650
rect 15225 4632 15245 4650
rect 15089 4628 15245 4632
rect 15184 4612 15245 4628
rect 19862 4779 19882 4797
rect 19900 4779 20018 4797
rect 19862 4758 20018 4779
rect 19918 4757 20018 4758
rect 19975 4721 20017 4757
rect 19866 4698 20017 4721
rect 19866 4680 19884 4698
rect 19902 4683 20017 4698
rect 19902 4680 19923 4683
rect 19866 4661 19923 4680
rect 9831 4562 9987 4566
rect 5059 4438 5101 4474
rect 4779 4404 4797 4422
rect 4815 4407 4930 4422
rect 5058 4437 5158 4438
rect 5058 4416 5214 4437
rect 4815 4404 4836 4407
rect 4779 4385 4836 4404
rect 5058 4398 5176 4416
rect 5194 4398 5214 4416
rect 9831 4544 9851 4562
rect 9869 4544 9987 4562
rect 9831 4523 9987 4544
rect 9887 4522 9987 4523
rect 9944 4486 9986 4522
rect 5058 4394 5214 4398
rect 5153 4378 5214 4394
rect 9835 4463 9986 4486
rect 10128 4479 10185 4498
rect 10128 4476 10149 4479
rect 9835 4445 9853 4463
rect 9871 4448 9986 4463
rect 10034 4461 10149 4476
rect 10167 4461 10185 4479
rect 9871 4445 9892 4448
rect 9835 4426 9892 4445
rect 10034 4438 10185 4461
rect 14806 4530 14867 4546
rect 14806 4526 14962 4530
rect 10034 4402 10076 4438
rect 10033 4401 10133 4402
rect 10033 4380 10189 4401
rect 10033 4362 10151 4380
rect 10169 4362 10189 4380
rect 14806 4508 14826 4526
rect 14844 4508 14962 4526
rect 15184 4520 15241 4539
rect 15184 4517 15205 4520
rect 14806 4487 14962 4508
rect 14862 4486 14962 4487
rect 15090 4502 15205 4517
rect 15223 4502 15241 4520
rect 14919 4450 14961 4486
rect 10033 4358 10189 4362
rect 97 4244 154 4263
rect 97 4241 118 4244
rect 3 4226 118 4241
rect 136 4226 154 4244
rect 3 4203 154 4226
rect 3 4167 45 4203
rect 2 4166 102 4167
rect 2 4145 158 4166
rect 2 4127 120 4145
rect 138 4127 158 4145
rect 4775 4296 4836 4312
rect 4775 4292 4931 4296
rect 4775 4274 4795 4292
rect 4813 4274 4931 4292
rect 5153 4285 5210 4304
rect 5153 4282 5174 4285
rect 4775 4253 4931 4274
rect 4831 4252 4931 4253
rect 5059 4267 5174 4282
rect 5192 4267 5210 4285
rect 4888 4216 4930 4252
rect 4779 4193 4930 4216
rect 5059 4244 5210 4267
rect 5059 4208 5101 4244
rect 2 4123 158 4127
rect 97 4107 158 4123
rect 4779 4175 4797 4193
rect 4815 4178 4930 4193
rect 5058 4207 5158 4208
rect 5058 4186 5214 4207
rect 4815 4175 4836 4178
rect 4779 4156 4836 4175
rect 5058 4168 5176 4186
rect 5194 4168 5214 4186
rect 9831 4337 9892 4353
rect 10128 4342 10189 4358
rect 9831 4333 9987 4337
rect 9831 4315 9851 4333
rect 9869 4315 9987 4333
rect 9831 4294 9987 4315
rect 9887 4293 9987 4294
rect 14810 4427 14961 4450
rect 15090 4479 15241 4502
rect 19862 4571 19923 4587
rect 19862 4567 20018 4571
rect 15090 4443 15132 4479
rect 14810 4409 14828 4427
rect 14846 4412 14961 4427
rect 15089 4442 15189 4443
rect 15089 4421 15245 4442
rect 14846 4409 14867 4412
rect 14810 4390 14867 4409
rect 15089 4403 15207 4421
rect 15225 4403 15245 4421
rect 19862 4549 19882 4567
rect 19900 4549 20018 4567
rect 19862 4528 20018 4549
rect 19918 4527 20018 4528
rect 19975 4491 20017 4527
rect 15089 4399 15245 4403
rect 15184 4383 15245 4399
rect 19866 4468 20017 4491
rect 19866 4450 19884 4468
rect 19902 4453 20017 4468
rect 19902 4450 19923 4453
rect 19866 4431 19923 4450
rect 9944 4257 9986 4293
rect 9835 4234 9986 4257
rect 10128 4249 10185 4268
rect 10128 4246 10149 4249
rect 5058 4164 5214 4168
rect 5153 4148 5214 4164
rect 4775 4109 4836 4125
rect 4775 4105 4931 4109
rect 4775 4087 4795 4105
rect 4813 4087 4931 4105
rect 9835 4216 9853 4234
rect 9871 4219 9986 4234
rect 10034 4231 10149 4246
rect 10167 4231 10185 4249
rect 9871 4216 9892 4219
rect 9835 4197 9892 4216
rect 10034 4208 10185 4231
rect 10034 4172 10076 4208
rect 10033 4171 10133 4172
rect 9831 4150 9892 4166
rect 10033 4150 10189 4171
rect 9831 4146 9987 4150
rect 9831 4128 9851 4146
rect 9869 4128 9987 4146
rect 10033 4132 10151 4150
rect 10169 4132 10189 4150
rect 14806 4301 14867 4317
rect 14806 4297 14962 4301
rect 14806 4279 14826 4297
rect 14844 4279 14962 4297
rect 15184 4290 15241 4309
rect 15184 4287 15205 4290
rect 14806 4258 14962 4279
rect 14862 4257 14962 4258
rect 15090 4272 15205 4287
rect 15223 4272 15241 4290
rect 14919 4221 14961 4257
rect 14810 4198 14961 4221
rect 15090 4249 15241 4272
rect 15090 4213 15132 4249
rect 10033 4128 10189 4132
rect 9831 4107 9987 4128
rect 10128 4112 10189 4128
rect 9887 4106 9987 4107
rect 4775 4066 4931 4087
rect 4831 4065 4931 4066
rect 4888 4029 4930 4065
rect 4779 4006 4930 4029
rect 9944 4070 9986 4106
rect 9835 4047 9986 4070
rect 14810 4180 14828 4198
rect 14846 4183 14961 4198
rect 15089 4212 15189 4213
rect 15089 4191 15245 4212
rect 14846 4180 14867 4183
rect 14810 4161 14867 4180
rect 15089 4173 15207 4191
rect 15225 4173 15245 4191
rect 19862 4342 19923 4358
rect 19862 4338 20018 4342
rect 19862 4320 19882 4338
rect 19900 4320 20018 4338
rect 19862 4299 20018 4320
rect 19918 4298 20018 4299
rect 19975 4262 20017 4298
rect 19866 4239 20017 4262
rect 15089 4169 15245 4173
rect 15184 4153 15245 4169
rect 14806 4114 14867 4130
rect 14806 4110 14962 4114
rect 14806 4092 14826 4110
rect 14844 4092 14962 4110
rect 19866 4221 19884 4239
rect 19902 4224 20017 4239
rect 19902 4221 19923 4224
rect 19866 4202 19923 4221
rect 19862 4155 19923 4171
rect 19862 4151 20018 4155
rect 19862 4133 19882 4151
rect 19900 4133 20018 4151
rect 19862 4112 20018 4133
rect 19918 4111 20018 4112
rect 14806 4071 14962 4092
rect 14862 4070 14962 4071
rect 4779 3988 4797 4006
rect 4815 3991 4930 4006
rect 4815 3988 4836 3991
rect 4779 3969 4836 3988
rect 98 3787 155 3806
rect 98 3784 119 3787
rect 4 3769 119 3784
rect 137 3769 155 3787
rect 9835 4029 9853 4047
rect 9871 4032 9986 4047
rect 9871 4029 9892 4032
rect 9835 4010 9892 4029
rect 14919 4034 14961 4070
rect 14810 4011 14961 4034
rect 19975 4075 20017 4111
rect 19866 4052 20017 4075
rect 5154 3828 5211 3847
rect 5154 3825 5175 3828
rect 5060 3810 5175 3825
rect 5193 3810 5211 3828
rect 14810 3993 14828 4011
rect 14846 3996 14961 4011
rect 14846 3993 14867 3996
rect 14810 3974 14867 3993
rect 4 3746 155 3769
rect 4 3710 46 3746
rect 5060 3787 5211 3810
rect 5060 3751 5102 3787
rect 10129 3792 10186 3811
rect 10129 3789 10150 3792
rect 10035 3774 10150 3789
rect 10168 3774 10186 3792
rect 19866 4034 19884 4052
rect 19902 4037 20017 4052
rect 19902 4034 19923 4037
rect 19866 4015 19923 4034
rect 15185 3833 15242 3852
rect 15185 3830 15206 3833
rect 15091 3815 15206 3830
rect 15224 3815 15242 3833
rect 5059 3750 5159 3751
rect 5059 3729 5215 3750
rect 3 3709 103 3710
rect 3 3688 159 3709
rect 3 3670 121 3688
rect 139 3670 159 3688
rect 3 3666 159 3670
rect 98 3650 159 3666
rect 98 3600 155 3619
rect 98 3597 119 3600
rect 4 3582 119 3597
rect 137 3582 155 3600
rect 5059 3711 5177 3729
rect 5195 3711 5215 3729
rect 5059 3707 5215 3711
rect 5154 3691 5215 3707
rect 4776 3652 4837 3668
rect 4776 3648 4932 3652
rect 4 3559 155 3582
rect 4 3523 46 3559
rect 3 3522 103 3523
rect 3 3501 159 3522
rect 3 3483 121 3501
rect 139 3483 159 3501
rect 3 3479 159 3483
rect 98 3463 159 3479
rect 4776 3630 4796 3648
rect 4814 3630 4932 3648
rect 5154 3641 5211 3660
rect 5154 3638 5175 3641
rect 4776 3609 4932 3630
rect 4832 3608 4932 3609
rect 5060 3623 5175 3638
rect 5193 3623 5211 3641
rect 10035 3751 10186 3774
rect 10035 3715 10077 3751
rect 15091 3792 15242 3815
rect 15091 3756 15133 3792
rect 15090 3755 15190 3756
rect 15090 3734 15246 3755
rect 10034 3714 10134 3715
rect 9832 3693 9893 3709
rect 10034 3693 10190 3714
rect 9832 3689 9988 3693
rect 4889 3572 4931 3608
rect 4780 3549 4931 3572
rect 5060 3600 5211 3623
rect 5060 3564 5102 3600
rect 4780 3531 4798 3549
rect 4816 3534 4931 3549
rect 5059 3563 5159 3564
rect 5059 3542 5215 3563
rect 4816 3531 4837 3534
rect 4780 3512 4837 3531
rect 5059 3524 5177 3542
rect 5195 3524 5215 3542
rect 5059 3520 5215 3524
rect 5154 3504 5215 3520
rect 9832 3671 9852 3689
rect 9870 3671 9988 3689
rect 10034 3675 10152 3693
rect 10170 3675 10190 3693
rect 10034 3671 10190 3675
rect 9832 3650 9988 3671
rect 10129 3655 10190 3671
rect 9888 3649 9988 3650
rect 9945 3613 9987 3649
rect 9836 3590 9987 3613
rect 10129 3605 10186 3624
rect 10129 3602 10150 3605
rect 9836 3572 9854 3590
rect 9872 3575 9987 3590
rect 10035 3587 10150 3602
rect 10168 3587 10186 3605
rect 15090 3716 15208 3734
rect 15226 3716 15246 3734
rect 15090 3712 15246 3716
rect 15185 3696 15246 3712
rect 14807 3657 14868 3673
rect 14807 3653 14963 3657
rect 9872 3572 9893 3575
rect 9836 3553 9893 3572
rect 10035 3564 10186 3587
rect 10035 3528 10077 3564
rect 98 3371 155 3390
rect 98 3368 119 3371
rect 4 3353 119 3368
rect 137 3353 155 3371
rect 4 3330 155 3353
rect 4776 3422 4837 3438
rect 4776 3418 4932 3422
rect 4 3294 46 3330
rect 3 3293 103 3294
rect 3 3272 159 3293
rect 3 3254 121 3272
rect 139 3254 159 3272
rect 4776 3400 4796 3418
rect 4814 3400 4932 3418
rect 5154 3412 5211 3431
rect 5154 3409 5175 3412
rect 4776 3379 4932 3400
rect 4832 3378 4932 3379
rect 5060 3394 5175 3409
rect 5193 3394 5211 3412
rect 4889 3342 4931 3378
rect 3 3250 159 3254
rect 98 3234 159 3250
rect 4780 3319 4931 3342
rect 5060 3371 5211 3394
rect 10034 3527 10134 3528
rect 10034 3506 10190 3527
rect 10034 3488 10152 3506
rect 10170 3488 10190 3506
rect 10034 3484 10190 3488
rect 9832 3463 9893 3479
rect 10129 3468 10190 3484
rect 14807 3635 14827 3653
rect 14845 3635 14963 3653
rect 15185 3646 15242 3665
rect 15185 3643 15206 3646
rect 14807 3614 14963 3635
rect 14863 3613 14963 3614
rect 15091 3628 15206 3643
rect 15224 3628 15242 3646
rect 19863 3698 19924 3714
rect 19863 3694 20019 3698
rect 14920 3577 14962 3613
rect 14811 3554 14962 3577
rect 15091 3605 15242 3628
rect 15091 3569 15133 3605
rect 14811 3536 14829 3554
rect 14847 3539 14962 3554
rect 15090 3568 15190 3569
rect 15090 3547 15246 3568
rect 14847 3536 14868 3539
rect 14811 3517 14868 3536
rect 15090 3529 15208 3547
rect 15226 3529 15246 3547
rect 15090 3525 15246 3529
rect 15185 3509 15246 3525
rect 19863 3676 19883 3694
rect 19901 3676 20019 3694
rect 19863 3655 20019 3676
rect 19919 3654 20019 3655
rect 19976 3618 20018 3654
rect 19867 3595 20018 3618
rect 19867 3577 19885 3595
rect 19903 3580 20018 3595
rect 19903 3577 19924 3580
rect 19867 3558 19924 3577
rect 9832 3459 9988 3463
rect 5060 3335 5102 3371
rect 4780 3301 4798 3319
rect 4816 3304 4931 3319
rect 5059 3334 5159 3335
rect 5059 3313 5215 3334
rect 4816 3301 4837 3304
rect 4780 3282 4837 3301
rect 5059 3295 5177 3313
rect 5195 3295 5215 3313
rect 9832 3441 9852 3459
rect 9870 3441 9988 3459
rect 9832 3420 9988 3441
rect 9888 3419 9988 3420
rect 9945 3383 9987 3419
rect 5059 3291 5215 3295
rect 5154 3275 5215 3291
rect 9836 3360 9987 3383
rect 10129 3376 10186 3395
rect 10129 3373 10150 3376
rect 9836 3342 9854 3360
rect 9872 3345 9987 3360
rect 10035 3358 10150 3373
rect 10168 3358 10186 3376
rect 9872 3342 9893 3345
rect 9836 3323 9893 3342
rect 10035 3335 10186 3358
rect 14807 3427 14868 3443
rect 14807 3423 14963 3427
rect 10035 3299 10077 3335
rect 10034 3298 10134 3299
rect 10034 3277 10190 3298
rect 10034 3259 10152 3277
rect 10170 3259 10190 3277
rect 14807 3405 14827 3423
rect 14845 3405 14963 3423
rect 15185 3417 15242 3436
rect 15185 3414 15206 3417
rect 14807 3384 14963 3405
rect 14863 3383 14963 3384
rect 15091 3399 15206 3414
rect 15224 3399 15242 3417
rect 14920 3347 14962 3383
rect 10034 3255 10190 3259
rect 98 3141 155 3160
rect 98 3138 119 3141
rect 4 3123 119 3138
rect 137 3123 155 3141
rect 4 3100 155 3123
rect 4 3064 46 3100
rect 3 3063 103 3064
rect 3 3042 159 3063
rect 3 3024 121 3042
rect 139 3024 159 3042
rect 4776 3193 4837 3209
rect 4776 3189 4932 3193
rect 4776 3171 4796 3189
rect 4814 3171 4932 3189
rect 5154 3182 5211 3201
rect 5154 3179 5175 3182
rect 4776 3150 4932 3171
rect 4832 3149 4932 3150
rect 5060 3164 5175 3179
rect 5193 3164 5211 3182
rect 4889 3113 4931 3149
rect 4780 3090 4931 3113
rect 5060 3141 5211 3164
rect 5060 3105 5102 3141
rect 3 3020 159 3024
rect 98 3004 159 3020
rect 4780 3072 4798 3090
rect 4816 3075 4931 3090
rect 5059 3104 5159 3105
rect 5059 3083 5215 3104
rect 4816 3072 4837 3075
rect 4780 3053 4837 3072
rect 5059 3065 5177 3083
rect 5195 3065 5215 3083
rect 9832 3234 9893 3250
rect 10129 3239 10190 3255
rect 9832 3230 9988 3234
rect 9832 3212 9852 3230
rect 9870 3212 9988 3230
rect 9832 3191 9988 3212
rect 9888 3190 9988 3191
rect 14811 3324 14962 3347
rect 15091 3376 15242 3399
rect 19863 3468 19924 3484
rect 19863 3464 20019 3468
rect 15091 3340 15133 3376
rect 14811 3306 14829 3324
rect 14847 3309 14962 3324
rect 15090 3339 15190 3340
rect 15090 3318 15246 3339
rect 14847 3306 14868 3309
rect 14811 3287 14868 3306
rect 15090 3300 15208 3318
rect 15226 3300 15246 3318
rect 19863 3446 19883 3464
rect 19901 3446 20019 3464
rect 19863 3425 20019 3446
rect 19919 3424 20019 3425
rect 19976 3388 20018 3424
rect 15090 3296 15246 3300
rect 15185 3280 15246 3296
rect 19867 3365 20018 3388
rect 19867 3347 19885 3365
rect 19903 3350 20018 3365
rect 19903 3347 19924 3350
rect 19867 3328 19924 3347
rect 9945 3154 9987 3190
rect 9836 3131 9987 3154
rect 10129 3146 10186 3165
rect 10129 3143 10150 3146
rect 5059 3061 5215 3065
rect 5154 3045 5215 3061
rect 4776 3006 4837 3022
rect 4776 3002 4932 3006
rect 4776 2984 4796 3002
rect 4814 2984 4932 3002
rect 9836 3113 9854 3131
rect 9872 3116 9987 3131
rect 10035 3128 10150 3143
rect 10168 3128 10186 3146
rect 9872 3113 9893 3116
rect 9836 3094 9893 3113
rect 10035 3105 10186 3128
rect 10035 3069 10077 3105
rect 10034 3068 10134 3069
rect 9832 3047 9893 3063
rect 10034 3047 10190 3068
rect 9832 3043 9988 3047
rect 9832 3025 9852 3043
rect 9870 3025 9988 3043
rect 10034 3029 10152 3047
rect 10170 3029 10190 3047
rect 14807 3198 14868 3214
rect 14807 3194 14963 3198
rect 14807 3176 14827 3194
rect 14845 3176 14963 3194
rect 15185 3187 15242 3206
rect 15185 3184 15206 3187
rect 14807 3155 14963 3176
rect 14863 3154 14963 3155
rect 15091 3169 15206 3184
rect 15224 3169 15242 3187
rect 14920 3118 14962 3154
rect 14811 3095 14962 3118
rect 15091 3146 15242 3169
rect 15091 3110 15133 3146
rect 10034 3025 10190 3029
rect 9832 3004 9988 3025
rect 10129 3009 10190 3025
rect 9888 3003 9988 3004
rect 4776 2963 4932 2984
rect 4832 2962 4932 2963
rect 4889 2926 4931 2962
rect 4780 2903 4931 2926
rect 4780 2885 4798 2903
rect 4816 2888 4931 2903
rect 9945 2967 9987 3003
rect 9836 2944 9987 2967
rect 14811 3077 14829 3095
rect 14847 3080 14962 3095
rect 15090 3109 15190 3110
rect 15090 3088 15246 3109
rect 14847 3077 14868 3080
rect 14811 3058 14868 3077
rect 15090 3070 15208 3088
rect 15226 3070 15246 3088
rect 19863 3239 19924 3255
rect 19863 3235 20019 3239
rect 19863 3217 19883 3235
rect 19901 3217 20019 3235
rect 19863 3196 20019 3217
rect 19919 3195 20019 3196
rect 19976 3159 20018 3195
rect 19867 3136 20018 3159
rect 15090 3066 15246 3070
rect 15185 3050 15246 3066
rect 14807 3011 14868 3027
rect 14807 3007 14963 3011
rect 14807 2989 14827 3007
rect 14845 2989 14963 3007
rect 19867 3118 19885 3136
rect 19903 3121 20018 3136
rect 19903 3118 19924 3121
rect 19867 3099 19924 3118
rect 19863 3052 19924 3068
rect 19863 3048 20019 3052
rect 19863 3030 19883 3048
rect 19901 3030 20019 3048
rect 19863 3009 20019 3030
rect 19919 3008 20019 3009
rect 14807 2968 14963 2989
rect 14863 2967 14963 2968
rect 9836 2926 9854 2944
rect 9872 2929 9987 2944
rect 9872 2926 9893 2929
rect 4816 2885 4837 2888
rect 4780 2866 4837 2885
rect 9836 2907 9893 2926
rect 14920 2931 14962 2967
rect 14811 2908 14962 2931
rect 14811 2890 14829 2908
rect 14847 2893 14962 2908
rect 19976 2972 20018 3008
rect 19867 2949 20018 2972
rect 19867 2931 19885 2949
rect 19903 2934 20018 2949
rect 19903 2931 19924 2934
rect 14847 2890 14868 2893
rect 98 2684 155 2703
rect 5154 2725 5211 2744
rect 14811 2871 14868 2890
rect 19867 2912 19924 2931
rect 5154 2722 5175 2725
rect 98 2681 119 2684
rect 4 2666 119 2681
rect 137 2666 155 2684
rect 4 2643 155 2666
rect 4 2607 46 2643
rect 5060 2707 5175 2722
rect 5193 2707 5211 2725
rect 5060 2684 5211 2707
rect 5060 2648 5102 2684
rect 10129 2689 10186 2708
rect 15185 2730 15242 2749
rect 15185 2727 15206 2730
rect 10129 2686 10150 2689
rect 10035 2671 10150 2686
rect 10168 2671 10186 2689
rect 5059 2647 5159 2648
rect 5059 2626 5215 2647
rect 3 2606 103 2607
rect 3 2585 159 2606
rect 3 2567 121 2585
rect 139 2567 159 2585
rect 3 2563 159 2567
rect 98 2547 159 2563
rect 98 2497 155 2516
rect 98 2494 119 2497
rect 4 2479 119 2494
rect 137 2479 155 2497
rect 5059 2608 5177 2626
rect 5195 2608 5215 2626
rect 5059 2604 5215 2608
rect 5154 2588 5215 2604
rect 4776 2549 4837 2565
rect 4776 2545 4932 2549
rect 4 2456 155 2479
rect 4 2420 46 2456
rect 3 2419 103 2420
rect 3 2398 159 2419
rect 3 2380 121 2398
rect 139 2380 159 2398
rect 3 2376 159 2380
rect 98 2360 159 2376
rect 4776 2527 4796 2545
rect 4814 2527 4932 2545
rect 5154 2538 5211 2557
rect 5154 2535 5175 2538
rect 4776 2506 4932 2527
rect 4832 2505 4932 2506
rect 5060 2520 5175 2535
rect 5193 2520 5211 2538
rect 10035 2648 10186 2671
rect 10035 2612 10077 2648
rect 15091 2712 15206 2727
rect 15224 2712 15242 2730
rect 15091 2689 15242 2712
rect 15091 2653 15133 2689
rect 15090 2652 15190 2653
rect 15090 2631 15246 2652
rect 10034 2611 10134 2612
rect 9832 2590 9893 2606
rect 10034 2590 10190 2611
rect 9832 2586 9988 2590
rect 4889 2469 4931 2505
rect 4780 2446 4931 2469
rect 5060 2497 5211 2520
rect 5060 2461 5102 2497
rect 4780 2428 4798 2446
rect 4816 2431 4931 2446
rect 5059 2460 5159 2461
rect 5059 2439 5215 2460
rect 4816 2428 4837 2431
rect 4780 2409 4837 2428
rect 5059 2421 5177 2439
rect 5195 2421 5215 2439
rect 5059 2417 5215 2421
rect 5154 2401 5215 2417
rect 9832 2568 9852 2586
rect 9870 2568 9988 2586
rect 10034 2572 10152 2590
rect 10170 2572 10190 2590
rect 10034 2568 10190 2572
rect 9832 2547 9988 2568
rect 10129 2552 10190 2568
rect 9888 2546 9988 2547
rect 9945 2510 9987 2546
rect 9836 2487 9987 2510
rect 10129 2502 10186 2521
rect 10129 2499 10150 2502
rect 9836 2469 9854 2487
rect 9872 2472 9987 2487
rect 10035 2484 10150 2499
rect 10168 2484 10186 2502
rect 15090 2613 15208 2631
rect 15226 2613 15246 2631
rect 15090 2609 15246 2613
rect 15185 2593 15246 2609
rect 14807 2554 14868 2570
rect 14807 2550 14963 2554
rect 9872 2469 9893 2472
rect 9836 2450 9893 2469
rect 10035 2461 10186 2484
rect 10035 2425 10077 2461
rect 98 2268 155 2287
rect 98 2265 119 2268
rect 4 2250 119 2265
rect 137 2250 155 2268
rect 4 2227 155 2250
rect 4776 2319 4837 2335
rect 4776 2315 4932 2319
rect 4 2191 46 2227
rect 3 2190 103 2191
rect 3 2169 159 2190
rect 3 2151 121 2169
rect 139 2151 159 2169
rect 4776 2297 4796 2315
rect 4814 2297 4932 2315
rect 5154 2309 5211 2328
rect 5154 2306 5175 2309
rect 4776 2276 4932 2297
rect 4832 2275 4932 2276
rect 5060 2291 5175 2306
rect 5193 2291 5211 2309
rect 4889 2239 4931 2275
rect 3 2147 159 2151
rect 98 2131 159 2147
rect 4780 2216 4931 2239
rect 5060 2268 5211 2291
rect 10034 2424 10134 2425
rect 10034 2403 10190 2424
rect 10034 2385 10152 2403
rect 10170 2385 10190 2403
rect 10034 2381 10190 2385
rect 9832 2360 9893 2376
rect 10129 2365 10190 2381
rect 14807 2532 14827 2550
rect 14845 2532 14963 2550
rect 15185 2543 15242 2562
rect 15185 2540 15206 2543
rect 14807 2511 14963 2532
rect 14863 2510 14963 2511
rect 15091 2525 15206 2540
rect 15224 2525 15242 2543
rect 19863 2595 19924 2611
rect 19863 2591 20019 2595
rect 14920 2474 14962 2510
rect 14811 2451 14962 2474
rect 15091 2502 15242 2525
rect 15091 2466 15133 2502
rect 14811 2433 14829 2451
rect 14847 2436 14962 2451
rect 15090 2465 15190 2466
rect 15090 2444 15246 2465
rect 14847 2433 14868 2436
rect 14811 2414 14868 2433
rect 15090 2426 15208 2444
rect 15226 2426 15246 2444
rect 15090 2422 15246 2426
rect 15185 2406 15246 2422
rect 19863 2573 19883 2591
rect 19901 2573 20019 2591
rect 19863 2552 20019 2573
rect 19919 2551 20019 2552
rect 19976 2515 20018 2551
rect 19867 2492 20018 2515
rect 19867 2474 19885 2492
rect 19903 2477 20018 2492
rect 19903 2474 19924 2477
rect 19867 2455 19924 2474
rect 9832 2356 9988 2360
rect 5060 2232 5102 2268
rect 4780 2198 4798 2216
rect 4816 2201 4931 2216
rect 5059 2231 5159 2232
rect 5059 2210 5215 2231
rect 4816 2198 4837 2201
rect 4780 2179 4837 2198
rect 5059 2192 5177 2210
rect 5195 2192 5215 2210
rect 9832 2338 9852 2356
rect 9870 2338 9988 2356
rect 9832 2317 9988 2338
rect 9888 2316 9988 2317
rect 9945 2280 9987 2316
rect 5059 2188 5215 2192
rect 5154 2172 5215 2188
rect 9836 2257 9987 2280
rect 10129 2273 10186 2292
rect 10129 2270 10150 2273
rect 9836 2239 9854 2257
rect 9872 2242 9987 2257
rect 10035 2255 10150 2270
rect 10168 2255 10186 2273
rect 9872 2239 9893 2242
rect 9836 2220 9893 2239
rect 10035 2232 10186 2255
rect 14807 2324 14868 2340
rect 14807 2320 14963 2324
rect 10035 2196 10077 2232
rect 10034 2195 10134 2196
rect 10034 2174 10190 2195
rect 10034 2156 10152 2174
rect 10170 2156 10190 2174
rect 14807 2302 14827 2320
rect 14845 2302 14963 2320
rect 15185 2314 15242 2333
rect 15185 2311 15206 2314
rect 14807 2281 14963 2302
rect 14863 2280 14963 2281
rect 15091 2296 15206 2311
rect 15224 2296 15242 2314
rect 14920 2244 14962 2280
rect 10034 2152 10190 2156
rect 98 2038 155 2057
rect 98 2035 119 2038
rect 4 2020 119 2035
rect 137 2020 155 2038
rect 4 1997 155 2020
rect 4 1961 46 1997
rect 3 1960 103 1961
rect 3 1939 159 1960
rect 3 1921 121 1939
rect 139 1921 159 1939
rect 4776 2090 4837 2106
rect 4776 2086 4932 2090
rect 4776 2068 4796 2086
rect 4814 2068 4932 2086
rect 5154 2079 5211 2098
rect 5154 2076 5175 2079
rect 4776 2047 4932 2068
rect 4832 2046 4932 2047
rect 5060 2061 5175 2076
rect 5193 2061 5211 2079
rect 4889 2010 4931 2046
rect 4780 1987 4931 2010
rect 5060 2038 5211 2061
rect 5060 2002 5102 2038
rect 3 1917 159 1921
rect 98 1901 159 1917
rect 4780 1969 4798 1987
rect 4816 1972 4931 1987
rect 5059 2001 5159 2002
rect 5059 1980 5215 2001
rect 4816 1969 4837 1972
rect 4780 1950 4837 1969
rect 5059 1962 5177 1980
rect 5195 1962 5215 1980
rect 9832 2131 9893 2147
rect 10129 2136 10190 2152
rect 9832 2127 9988 2131
rect 9832 2109 9852 2127
rect 9870 2109 9988 2127
rect 9832 2088 9988 2109
rect 9888 2087 9988 2088
rect 14811 2221 14962 2244
rect 15091 2273 15242 2296
rect 19863 2365 19924 2381
rect 19863 2361 20019 2365
rect 15091 2237 15133 2273
rect 14811 2203 14829 2221
rect 14847 2206 14962 2221
rect 15090 2236 15190 2237
rect 15090 2215 15246 2236
rect 14847 2203 14868 2206
rect 14811 2184 14868 2203
rect 15090 2197 15208 2215
rect 15226 2197 15246 2215
rect 19863 2343 19883 2361
rect 19901 2343 20019 2361
rect 19863 2322 20019 2343
rect 19919 2321 20019 2322
rect 19976 2285 20018 2321
rect 15090 2193 15246 2197
rect 15185 2177 15246 2193
rect 19867 2262 20018 2285
rect 19867 2244 19885 2262
rect 19903 2247 20018 2262
rect 19903 2244 19924 2247
rect 19867 2225 19924 2244
rect 9945 2051 9987 2087
rect 9836 2028 9987 2051
rect 10129 2043 10186 2062
rect 10129 2040 10150 2043
rect 5059 1958 5215 1962
rect 5154 1942 5215 1958
rect 4776 1903 4837 1919
rect 4776 1899 4932 1903
rect 4776 1881 4796 1899
rect 4814 1881 4932 1899
rect 9836 2010 9854 2028
rect 9872 2013 9987 2028
rect 10035 2025 10150 2040
rect 10168 2025 10186 2043
rect 9872 2010 9893 2013
rect 9836 1991 9893 2010
rect 10035 2002 10186 2025
rect 10035 1966 10077 2002
rect 10034 1965 10134 1966
rect 9832 1944 9893 1960
rect 10034 1944 10190 1965
rect 9832 1940 9988 1944
rect 9832 1922 9852 1940
rect 9870 1922 9988 1940
rect 10034 1926 10152 1944
rect 10170 1926 10190 1944
rect 14807 2095 14868 2111
rect 14807 2091 14963 2095
rect 14807 2073 14827 2091
rect 14845 2073 14963 2091
rect 15185 2084 15242 2103
rect 15185 2081 15206 2084
rect 14807 2052 14963 2073
rect 14863 2051 14963 2052
rect 15091 2066 15206 2081
rect 15224 2066 15242 2084
rect 14920 2015 14962 2051
rect 14811 1992 14962 2015
rect 15091 2043 15242 2066
rect 15091 2007 15133 2043
rect 10034 1922 10190 1926
rect 9832 1901 9988 1922
rect 10129 1906 10190 1922
rect 9888 1900 9988 1901
rect 4776 1860 4932 1881
rect 4832 1859 4932 1860
rect 4889 1823 4931 1859
rect 4780 1800 4931 1823
rect 9945 1864 9987 1900
rect 9836 1841 9987 1864
rect 14811 1974 14829 1992
rect 14847 1977 14962 1992
rect 15090 2006 15190 2007
rect 15090 1985 15246 2006
rect 14847 1974 14868 1977
rect 14811 1955 14868 1974
rect 15090 1967 15208 1985
rect 15226 1967 15246 1985
rect 19863 2136 19924 2152
rect 19863 2132 20019 2136
rect 19863 2114 19883 2132
rect 19901 2114 20019 2132
rect 19863 2093 20019 2114
rect 19919 2092 20019 2093
rect 19976 2056 20018 2092
rect 19867 2033 20018 2056
rect 15090 1963 15246 1967
rect 15185 1947 15246 1963
rect 14807 1908 14868 1924
rect 14807 1904 14963 1908
rect 14807 1886 14827 1904
rect 14845 1886 14963 1904
rect 19867 2015 19885 2033
rect 19903 2018 20018 2033
rect 19903 2015 19924 2018
rect 19867 1996 19924 2015
rect 19863 1949 19924 1965
rect 19863 1945 20019 1949
rect 19863 1927 19883 1945
rect 19901 1927 20019 1945
rect 19863 1906 20019 1927
rect 19919 1905 20019 1906
rect 14807 1865 14963 1886
rect 14863 1864 14963 1865
rect 4780 1782 4798 1800
rect 4816 1785 4931 1800
rect 4816 1782 4837 1785
rect 4780 1763 4837 1782
rect 99 1581 156 1600
rect 99 1578 120 1581
rect 5 1563 120 1578
rect 138 1563 156 1581
rect 9836 1823 9854 1841
rect 9872 1826 9987 1841
rect 9872 1823 9893 1826
rect 9836 1804 9893 1823
rect 14920 1828 14962 1864
rect 14811 1805 14962 1828
rect 19976 1869 20018 1905
rect 19867 1846 20018 1869
rect 5155 1622 5212 1641
rect 5155 1619 5176 1622
rect 5061 1604 5176 1619
rect 5194 1604 5212 1622
rect 14811 1787 14829 1805
rect 14847 1790 14962 1805
rect 14847 1787 14868 1790
rect 14811 1768 14868 1787
rect 5 1540 156 1563
rect 5 1504 47 1540
rect 5061 1581 5212 1604
rect 5061 1545 5103 1581
rect 10130 1586 10187 1605
rect 10130 1583 10151 1586
rect 10036 1568 10151 1583
rect 10169 1568 10187 1586
rect 19867 1828 19885 1846
rect 19903 1831 20018 1846
rect 19903 1828 19924 1831
rect 19867 1809 19924 1828
rect 15186 1627 15243 1646
rect 15186 1624 15207 1627
rect 15092 1609 15207 1624
rect 15225 1609 15243 1627
rect 5060 1544 5160 1545
rect 5060 1523 5216 1544
rect 4 1503 104 1504
rect 4 1482 160 1503
rect 4 1464 122 1482
rect 140 1464 160 1482
rect 4 1460 160 1464
rect 99 1444 160 1460
rect 99 1394 156 1413
rect 99 1391 120 1394
rect 5 1376 120 1391
rect 138 1376 156 1394
rect 5060 1505 5178 1523
rect 5196 1505 5216 1523
rect 5060 1501 5216 1505
rect 5155 1485 5216 1501
rect 4777 1446 4838 1462
rect 4777 1442 4933 1446
rect 5 1353 156 1376
rect 5 1317 47 1353
rect 4 1316 104 1317
rect 4 1295 160 1316
rect 4 1277 122 1295
rect 140 1277 160 1295
rect 4 1273 160 1277
rect 99 1257 160 1273
rect 4777 1424 4797 1442
rect 4815 1424 4933 1442
rect 5155 1435 5212 1454
rect 5155 1432 5176 1435
rect 4777 1403 4933 1424
rect 4833 1402 4933 1403
rect 5061 1417 5176 1432
rect 5194 1417 5212 1435
rect 10036 1545 10187 1568
rect 10036 1509 10078 1545
rect 15092 1586 15243 1609
rect 15092 1550 15134 1586
rect 15091 1549 15191 1550
rect 15091 1528 15247 1549
rect 10035 1508 10135 1509
rect 9833 1487 9894 1503
rect 10035 1487 10191 1508
rect 9833 1483 9989 1487
rect 4890 1366 4932 1402
rect 4781 1343 4932 1366
rect 5061 1394 5212 1417
rect 5061 1358 5103 1394
rect 4781 1325 4799 1343
rect 4817 1328 4932 1343
rect 5060 1357 5160 1358
rect 5060 1336 5216 1357
rect 4817 1325 4838 1328
rect 4781 1306 4838 1325
rect 5060 1318 5178 1336
rect 5196 1318 5216 1336
rect 5060 1314 5216 1318
rect 5155 1298 5216 1314
rect 9833 1465 9853 1483
rect 9871 1465 9989 1483
rect 10035 1469 10153 1487
rect 10171 1469 10191 1487
rect 10035 1465 10191 1469
rect 9833 1444 9989 1465
rect 10130 1449 10191 1465
rect 9889 1443 9989 1444
rect 9946 1407 9988 1443
rect 9837 1384 9988 1407
rect 10130 1399 10187 1418
rect 10130 1396 10151 1399
rect 9837 1366 9855 1384
rect 9873 1369 9988 1384
rect 10036 1381 10151 1396
rect 10169 1381 10187 1399
rect 15091 1510 15209 1528
rect 15227 1510 15247 1528
rect 15091 1506 15247 1510
rect 15186 1490 15247 1506
rect 14808 1451 14869 1467
rect 14808 1447 14964 1451
rect 9873 1366 9894 1369
rect 9837 1347 9894 1366
rect 10036 1358 10187 1381
rect 10036 1322 10078 1358
rect 99 1165 156 1184
rect 99 1162 120 1165
rect 5 1147 120 1162
rect 138 1147 156 1165
rect 5 1124 156 1147
rect 4777 1216 4838 1232
rect 4777 1212 4933 1216
rect 5 1088 47 1124
rect 4 1087 104 1088
rect 4 1066 160 1087
rect 4 1048 122 1066
rect 140 1048 160 1066
rect 4777 1194 4797 1212
rect 4815 1194 4933 1212
rect 5155 1206 5212 1225
rect 5155 1203 5176 1206
rect 4777 1173 4933 1194
rect 4833 1172 4933 1173
rect 5061 1188 5176 1203
rect 5194 1188 5212 1206
rect 4890 1136 4932 1172
rect 4 1044 160 1048
rect 99 1028 160 1044
rect 4781 1113 4932 1136
rect 5061 1165 5212 1188
rect 10035 1321 10135 1322
rect 10035 1300 10191 1321
rect 10035 1282 10153 1300
rect 10171 1282 10191 1300
rect 10035 1278 10191 1282
rect 9833 1257 9894 1273
rect 10130 1262 10191 1278
rect 14808 1429 14828 1447
rect 14846 1429 14964 1447
rect 15186 1440 15243 1459
rect 15186 1437 15207 1440
rect 14808 1408 14964 1429
rect 14864 1407 14964 1408
rect 15092 1422 15207 1437
rect 15225 1422 15243 1440
rect 19864 1492 19925 1508
rect 19864 1488 20020 1492
rect 14921 1371 14963 1407
rect 14812 1348 14963 1371
rect 15092 1399 15243 1422
rect 15092 1363 15134 1399
rect 14812 1330 14830 1348
rect 14848 1333 14963 1348
rect 15091 1362 15191 1363
rect 15091 1341 15247 1362
rect 14848 1330 14869 1333
rect 14812 1311 14869 1330
rect 15091 1323 15209 1341
rect 15227 1323 15247 1341
rect 15091 1319 15247 1323
rect 15186 1303 15247 1319
rect 19864 1470 19884 1488
rect 19902 1470 20020 1488
rect 19864 1449 20020 1470
rect 19920 1448 20020 1449
rect 19977 1412 20019 1448
rect 19868 1389 20019 1412
rect 19868 1371 19886 1389
rect 19904 1374 20019 1389
rect 19904 1371 19925 1374
rect 19868 1352 19925 1371
rect 9833 1253 9989 1257
rect 5061 1129 5103 1165
rect 4781 1095 4799 1113
rect 4817 1098 4932 1113
rect 5060 1128 5160 1129
rect 5060 1107 5216 1128
rect 4817 1095 4838 1098
rect 4781 1076 4838 1095
rect 5060 1089 5178 1107
rect 5196 1089 5216 1107
rect 9833 1235 9853 1253
rect 9871 1235 9989 1253
rect 9833 1214 9989 1235
rect 9889 1213 9989 1214
rect 9946 1177 9988 1213
rect 5060 1085 5216 1089
rect 5155 1069 5216 1085
rect 9837 1154 9988 1177
rect 10130 1170 10187 1189
rect 10130 1167 10151 1170
rect 9837 1136 9855 1154
rect 9873 1139 9988 1154
rect 10036 1152 10151 1167
rect 10169 1152 10187 1170
rect 9873 1136 9894 1139
rect 9837 1117 9894 1136
rect 10036 1129 10187 1152
rect 14808 1221 14869 1237
rect 14808 1217 14964 1221
rect 10036 1093 10078 1129
rect 10035 1092 10135 1093
rect 10035 1071 10191 1092
rect 10035 1053 10153 1071
rect 10171 1053 10191 1071
rect 14808 1199 14828 1217
rect 14846 1199 14964 1217
rect 15186 1211 15243 1230
rect 15186 1208 15207 1211
rect 14808 1178 14964 1199
rect 14864 1177 14964 1178
rect 15092 1193 15207 1208
rect 15225 1193 15243 1211
rect 14921 1141 14963 1177
rect 10035 1049 10191 1053
rect 99 935 156 954
rect 99 932 120 935
rect 5 917 120 932
rect 138 917 156 935
rect 5 894 156 917
rect 5 858 47 894
rect 4 857 104 858
rect 4 836 160 857
rect 4 818 122 836
rect 140 818 160 836
rect 4777 987 4838 1003
rect 4777 983 4933 987
rect 4777 965 4797 983
rect 4815 965 4933 983
rect 5155 976 5212 995
rect 5155 973 5176 976
rect 4777 944 4933 965
rect 4833 943 4933 944
rect 5061 958 5176 973
rect 5194 958 5212 976
rect 4890 907 4932 943
rect 4781 884 4932 907
rect 5061 935 5212 958
rect 5061 899 5103 935
rect 4 814 160 818
rect 99 798 160 814
rect 4781 866 4799 884
rect 4817 869 4932 884
rect 5060 898 5160 899
rect 5060 877 5216 898
rect 4817 866 4838 869
rect 4781 847 4838 866
rect 5060 859 5178 877
rect 5196 859 5216 877
rect 9833 1028 9894 1044
rect 10130 1033 10191 1049
rect 9833 1024 9989 1028
rect 9833 1006 9853 1024
rect 9871 1006 9989 1024
rect 9833 985 9989 1006
rect 9889 984 9989 985
rect 14812 1118 14963 1141
rect 15092 1170 15243 1193
rect 19864 1262 19925 1278
rect 19864 1258 20020 1262
rect 15092 1134 15134 1170
rect 14812 1100 14830 1118
rect 14848 1103 14963 1118
rect 15091 1133 15191 1134
rect 15091 1112 15247 1133
rect 14848 1100 14869 1103
rect 14812 1081 14869 1100
rect 15091 1094 15209 1112
rect 15227 1094 15247 1112
rect 19864 1240 19884 1258
rect 19902 1240 20020 1258
rect 19864 1219 20020 1240
rect 19920 1218 20020 1219
rect 19977 1182 20019 1218
rect 15091 1090 15247 1094
rect 15186 1074 15247 1090
rect 19868 1159 20019 1182
rect 19868 1141 19886 1159
rect 19904 1144 20019 1159
rect 19904 1141 19925 1144
rect 19868 1122 19925 1141
rect 9946 948 9988 984
rect 9837 925 9988 948
rect 10130 940 10187 959
rect 10130 937 10151 940
rect 5060 855 5216 859
rect 5155 839 5216 855
rect 4777 800 4838 816
rect 4777 796 4933 800
rect 4777 778 4797 796
rect 4815 778 4933 796
rect 9837 907 9855 925
rect 9873 910 9988 925
rect 10036 922 10151 937
rect 10169 922 10187 940
rect 9873 907 9894 910
rect 9837 888 9894 907
rect 10036 899 10187 922
rect 10036 863 10078 899
rect 10035 862 10135 863
rect 9833 841 9894 857
rect 10035 841 10191 862
rect 9833 837 9989 841
rect 9833 819 9853 837
rect 9871 819 9989 837
rect 10035 823 10153 841
rect 10171 823 10191 841
rect 14808 992 14869 1008
rect 14808 988 14964 992
rect 14808 970 14828 988
rect 14846 970 14964 988
rect 15186 981 15243 1000
rect 15186 978 15207 981
rect 14808 949 14964 970
rect 14864 948 14964 949
rect 15092 963 15207 978
rect 15225 963 15243 981
rect 14921 912 14963 948
rect 14812 889 14963 912
rect 15092 940 15243 963
rect 15092 904 15134 940
rect 10035 819 10191 823
rect 9833 798 9989 819
rect 10130 803 10191 819
rect 9889 797 9989 798
rect 4777 757 4933 778
rect 4833 756 4933 757
rect 4890 720 4932 756
rect 9946 761 9988 797
rect 9837 738 9988 761
rect 14812 871 14830 889
rect 14848 874 14963 889
rect 15091 903 15191 904
rect 15091 882 15247 903
rect 14848 871 14869 874
rect 14812 852 14869 871
rect 15091 864 15209 882
rect 15227 864 15247 882
rect 19864 1033 19925 1049
rect 19864 1029 20020 1033
rect 19864 1011 19884 1029
rect 19902 1011 20020 1029
rect 19864 990 20020 1011
rect 19920 989 20020 990
rect 19977 953 20019 989
rect 19868 930 20019 953
rect 15091 860 15247 864
rect 15186 844 15247 860
rect 14808 805 14869 821
rect 14808 801 14964 805
rect 14808 783 14828 801
rect 14846 783 14964 801
rect 19868 912 19886 930
rect 19904 915 20019 930
rect 19904 912 19925 915
rect 19868 893 19925 912
rect 19864 846 19925 862
rect 19864 842 20020 846
rect 19864 824 19884 842
rect 19902 824 20020 842
rect 19864 803 20020 824
rect 19920 802 20020 803
rect 14808 762 14964 783
rect 14864 761 14964 762
rect 4781 697 4932 720
rect 9837 720 9855 738
rect 9873 723 9988 738
rect 9873 720 9894 723
rect 4781 679 4799 697
rect 4817 682 4932 697
rect 9837 701 9894 720
rect 14921 725 14963 761
rect 19977 766 20019 802
rect 19868 743 20019 766
rect 4817 679 4838 682
rect 4781 660 4838 679
rect 14812 702 14963 725
rect 19868 725 19886 743
rect 19904 728 20019 743
rect 19904 725 19925 728
rect 14812 684 14830 702
rect 14848 687 14963 702
rect 19868 706 19925 725
rect 14848 684 14869 687
rect 14812 665 14869 684
<< locali >>
rect 19224 9490 19262 9492
rect 9193 9485 9231 9487
rect 9193 9452 9879 9485
rect 4137 9444 4175 9446
rect 4780 9444 5205 9446
rect 4137 9413 5214 9444
rect 4137 9411 4386 9413
rect 4542 9411 5214 9413
rect 105 9304 144 9361
rect 3729 9323 3897 9324
rect 4137 9323 4175 9411
rect 4780 9410 5215 9411
rect 4783 9387 4823 9410
rect 5135 9406 5215 9410
rect 4400 9354 4512 9372
rect 4400 9353 4443 9354
rect 105 9302 153 9304
rect 105 9284 116 9302
rect 134 9284 153 9302
rect 3729 9300 4175 9323
rect 4401 9352 4443 9353
rect 4401 9332 4408 9352
rect 4427 9332 4443 9352
rect 4401 9324 4443 9332
rect 4471 9352 4512 9354
rect 4471 9332 4485 9352
rect 4504 9332 4512 9352
rect 4784 9343 4823 9387
rect 5157 9362 5215 9406
rect 5159 9348 5215 9362
rect 4471 9324 4512 9332
rect 4401 9318 4512 9324
rect 3729 9297 4173 9300
rect 3729 9295 3897 9297
rect 105 9275 153 9284
rect 106 9274 153 9275
rect 419 9279 529 9293
rect 419 9276 462 9279
rect 419 9271 423 9276
rect 341 9249 423 9271
rect 452 9249 462 9276
rect 490 9252 497 9279
rect 526 9271 529 9279
rect 526 9252 591 9271
rect 490 9249 591 9252
rect 341 9247 591 9249
rect 109 9211 146 9212
rect 105 9208 146 9211
rect 105 9203 147 9208
rect 105 9185 118 9203
rect 136 9185 147 9203
rect 105 9171 147 9185
rect 185 9171 232 9175
rect 105 9165 232 9171
rect 105 9136 193 9165
rect 222 9136 232 9165
rect 341 9168 378 9247
rect 419 9234 529 9247
rect 493 9178 524 9179
rect 341 9148 350 9168
rect 370 9148 378 9168
rect 341 9138 378 9148
rect 437 9168 524 9178
rect 437 9148 446 9168
rect 466 9148 524 9168
rect 437 9139 524 9148
rect 437 9138 474 9139
rect 105 9132 232 9136
rect 105 9115 144 9132
rect 185 9131 232 9132
rect 105 9097 116 9115
rect 134 9097 144 9115
rect 105 9088 144 9097
rect 106 9087 143 9088
rect 493 9086 524 9139
rect 554 9168 591 9247
rect 762 9244 1155 9264
rect 1175 9244 1178 9264
rect 762 9239 1178 9244
rect 762 9238 1103 9239
rect 706 9178 737 9179
rect 554 9148 563 9168
rect 583 9148 591 9168
rect 554 9138 591 9148
rect 650 9171 737 9178
rect 650 9168 711 9171
rect 650 9148 659 9168
rect 679 9151 711 9168
rect 732 9151 737 9171
rect 679 9148 737 9151
rect 650 9141 737 9148
rect 762 9168 799 9238
rect 1065 9237 1102 9238
rect 914 9178 950 9179
rect 762 9148 771 9168
rect 791 9148 799 9168
rect 650 9139 706 9141
rect 650 9138 687 9139
rect 762 9138 799 9148
rect 858 9168 1006 9178
rect 1106 9175 1202 9177
rect 858 9148 867 9168
rect 887 9148 977 9168
rect 997 9148 1006 9168
rect 858 9139 1006 9148
rect 1064 9168 1202 9175
rect 1064 9148 1073 9168
rect 1093 9148 1202 9168
rect 1064 9139 1202 9148
rect 858 9138 895 9139
rect 914 9087 950 9139
rect 969 9138 1006 9139
rect 1065 9138 1102 9139
rect 385 9085 426 9086
rect 277 9078 426 9085
rect 277 9058 395 9078
rect 415 9058 426 9078
rect 277 9050 426 9058
rect 493 9082 852 9086
rect 493 9077 815 9082
rect 493 9053 606 9077
rect 630 9058 815 9077
rect 839 9058 852 9082
rect 630 9053 852 9058
rect 493 9050 852 9053
rect 914 9050 949 9087
rect 1017 9084 1117 9087
rect 1017 9080 1084 9084
rect 1017 9054 1029 9080
rect 1055 9058 1084 9080
rect 1110 9058 1117 9084
rect 1055 9054 1117 9058
rect 1017 9050 1117 9054
rect 493 9029 524 9050
rect 914 9029 950 9050
rect 336 9028 373 9029
rect 110 9025 144 9026
rect 109 9016 146 9025
rect 109 8998 118 9016
rect 136 8998 146 9016
rect 109 8988 146 8998
rect 335 9019 373 9028
rect 335 8999 344 9019
rect 364 8999 373 9019
rect 335 8991 373 8999
rect 439 9023 524 9029
rect 549 9028 586 9029
rect 439 9003 447 9023
rect 467 9003 524 9023
rect 439 8995 524 9003
rect 548 9019 586 9028
rect 548 8999 557 9019
rect 577 8999 586 9019
rect 439 8994 475 8995
rect 548 8991 586 8999
rect 652 9023 737 9029
rect 757 9028 794 9029
rect 652 9003 660 9023
rect 680 9022 737 9023
rect 680 9003 709 9022
rect 652 9002 709 9003
rect 730 9002 737 9022
rect 652 8995 737 9002
rect 756 9019 794 9028
rect 756 8999 765 9019
rect 785 8999 794 9019
rect 652 8994 688 8995
rect 756 8991 794 8999
rect 860 9023 1004 9029
rect 860 9003 868 9023
rect 888 9022 976 9023
rect 888 9003 919 9022
rect 860 9002 919 9003
rect 944 9003 976 9022
rect 996 9003 1004 9023
rect 944 9002 1004 9003
rect 860 8995 1004 9002
rect 860 8994 896 8995
rect 968 8994 1004 8995
rect 1070 9028 1107 9029
rect 1070 9027 1108 9028
rect 1070 9019 1134 9027
rect 1070 8999 1079 9019
rect 1099 9005 1134 9019
rect 1154 9005 1157 9025
rect 1099 9000 1157 9005
rect 1099 8999 1134 9000
rect 110 8960 144 8988
rect 336 8962 373 8991
rect 337 8960 373 8962
rect 549 8960 586 8991
rect 110 8959 282 8960
rect 110 8927 296 8959
rect 337 8938 586 8960
rect 757 8959 794 8991
rect 1070 8987 1134 8999
rect 1174 8961 1201 9139
rect 3729 9117 3756 9295
rect 3796 9257 3860 9269
rect 4136 9265 4173 9297
rect 4344 9296 4593 9318
rect 4344 9265 4381 9296
rect 4557 9294 4593 9296
rect 4557 9265 4594 9294
rect 3796 9256 3831 9257
rect 3773 9251 3831 9256
rect 3773 9231 3776 9251
rect 3796 9237 3831 9251
rect 3851 9237 3860 9257
rect 3796 9229 3860 9237
rect 3822 9228 3860 9229
rect 3823 9227 3860 9228
rect 3926 9261 3962 9262
rect 4034 9261 4070 9262
rect 3926 9256 4070 9261
rect 3926 9253 3988 9256
rect 3926 9233 3934 9253
rect 3954 9236 3988 9253
rect 4011 9253 4070 9256
rect 4011 9236 4042 9253
rect 3954 9233 4042 9236
rect 4062 9233 4070 9253
rect 3926 9227 4070 9233
rect 4136 9257 4174 9265
rect 4242 9261 4278 9262
rect 4136 9237 4145 9257
rect 4165 9237 4174 9257
rect 4136 9228 4174 9237
rect 4193 9254 4278 9261
rect 4193 9234 4200 9254
rect 4221 9253 4278 9254
rect 4221 9234 4250 9253
rect 4193 9233 4250 9234
rect 4270 9233 4278 9253
rect 4136 9227 4173 9228
rect 4193 9227 4278 9233
rect 4344 9257 4382 9265
rect 4455 9261 4491 9262
rect 4344 9237 4353 9257
rect 4373 9237 4382 9257
rect 4344 9228 4382 9237
rect 4406 9253 4491 9261
rect 4406 9233 4463 9253
rect 4483 9233 4491 9253
rect 4344 9227 4381 9228
rect 4406 9227 4491 9233
rect 4557 9257 4595 9265
rect 4557 9237 4566 9257
rect 4586 9237 4595 9257
rect 4557 9228 4595 9237
rect 4557 9227 4594 9228
rect 3980 9206 4016 9227
rect 4406 9206 4437 9227
rect 3813 9202 3913 9206
rect 3813 9198 3875 9202
rect 3813 9172 3820 9198
rect 3846 9176 3875 9198
rect 3901 9176 3913 9202
rect 3846 9172 3913 9176
rect 3813 9169 3913 9172
rect 3981 9169 4016 9206
rect 4078 9203 4437 9206
rect 4078 9198 4300 9203
rect 4078 9174 4091 9198
rect 4115 9179 4300 9198
rect 4324 9179 4437 9203
rect 4115 9174 4437 9179
rect 4078 9170 4437 9174
rect 4504 9198 4653 9206
rect 4504 9178 4515 9198
rect 4535 9178 4653 9198
rect 4504 9171 4653 9178
rect 4504 9170 4545 9171
rect 3828 9117 3865 9118
rect 3924 9117 3961 9118
rect 3980 9117 4016 9169
rect 4035 9117 4072 9118
rect 3728 9108 3866 9117
rect 3728 9088 3837 9108
rect 3857 9088 3866 9108
rect 3728 9081 3866 9088
rect 3924 9108 4072 9117
rect 3924 9088 3933 9108
rect 3953 9088 4043 9108
rect 4063 9088 4072 9108
rect 3728 9079 3824 9081
rect 3924 9078 4072 9088
rect 4131 9108 4168 9118
rect 4243 9117 4280 9118
rect 4224 9115 4280 9117
rect 4131 9088 4139 9108
rect 4159 9088 4168 9108
rect 3980 9077 4016 9078
rect 1357 9035 1467 9049
rect 1357 9032 1400 9035
rect 1357 9027 1361 9032
rect 1033 8959 1201 8961
rect 757 8953 1201 8959
rect 110 8895 144 8927
rect 106 8886 144 8895
rect 106 8868 116 8886
rect 134 8868 144 8886
rect 106 8862 144 8868
rect 262 8864 296 8927
rect 418 8932 529 8938
rect 418 8924 459 8932
rect 418 8904 426 8924
rect 445 8904 459 8924
rect 418 8902 459 8904
rect 487 8924 529 8932
rect 487 8904 503 8924
rect 522 8904 529 8924
rect 487 8902 529 8904
rect 418 8887 529 8902
rect 756 8933 1201 8953
rect 756 8864 794 8933
rect 1033 8932 1201 8933
rect 1279 9005 1361 9027
rect 1390 9005 1400 9032
rect 1428 9008 1435 9035
rect 1464 9027 1467 9035
rect 3462 9044 3573 9059
rect 3462 9042 3504 9044
rect 1464 9008 1529 9027
rect 1428 9005 1529 9008
rect 1279 9003 1529 9005
rect 1279 8924 1316 9003
rect 1357 8990 1467 9003
rect 1431 8934 1462 8935
rect 1279 8904 1288 8924
rect 1308 8904 1316 8924
rect 1279 8894 1316 8904
rect 1375 8924 1462 8934
rect 1375 8904 1384 8924
rect 1404 8904 1462 8924
rect 1375 8895 1462 8904
rect 1375 8894 1412 8895
rect 106 8858 143 8862
rect 262 8853 794 8864
rect 261 8837 794 8853
rect 1431 8842 1462 8895
rect 1492 8924 1529 9003
rect 1700 9000 2093 9020
rect 2113 9000 2116 9020
rect 3195 9015 3236 9024
rect 1700 8995 2116 9000
rect 2790 9013 2958 9014
rect 3195 9013 3204 9015
rect 1700 8994 2041 8995
rect 1644 8934 1675 8935
rect 1492 8904 1501 8924
rect 1521 8904 1529 8924
rect 1492 8894 1529 8904
rect 1588 8927 1675 8934
rect 1588 8924 1649 8927
rect 1588 8904 1597 8924
rect 1617 8907 1649 8924
rect 1670 8907 1675 8927
rect 1617 8904 1675 8907
rect 1588 8897 1675 8904
rect 1700 8924 1737 8994
rect 2003 8993 2040 8994
rect 2790 8993 3204 9013
rect 3230 8993 3236 9015
rect 3462 9022 3469 9042
rect 3488 9022 3504 9042
rect 3462 9014 3504 9022
rect 3532 9042 3573 9044
rect 3532 9022 3546 9042
rect 3565 9022 3573 9042
rect 3532 9014 3573 9022
rect 3828 9018 3865 9019
rect 4131 9018 4168 9088
rect 4193 9108 4280 9115
rect 4193 9105 4251 9108
rect 4193 9085 4198 9105
rect 4219 9088 4251 9105
rect 4271 9088 4280 9108
rect 4219 9085 4280 9088
rect 4193 9078 4280 9085
rect 4339 9108 4376 9118
rect 4339 9088 4347 9108
rect 4367 9088 4376 9108
rect 4193 9077 4224 9078
rect 3827 9017 4168 9018
rect 3462 9008 3573 9014
rect 3752 9012 4168 9017
rect 2790 8987 3236 8993
rect 2790 8985 2958 8987
rect 1852 8934 1888 8935
rect 1700 8904 1709 8924
rect 1729 8904 1737 8924
rect 1588 8895 1644 8897
rect 1588 8894 1625 8895
rect 1700 8894 1737 8904
rect 1796 8924 1944 8934
rect 2044 8931 2140 8933
rect 1796 8904 1805 8924
rect 1825 8904 1915 8924
rect 1935 8904 1944 8924
rect 1796 8895 1944 8904
rect 2002 8924 2140 8931
rect 2002 8904 2011 8924
rect 2031 8904 2140 8924
rect 2002 8895 2140 8904
rect 1796 8894 1833 8895
rect 1852 8843 1888 8895
rect 1907 8894 1944 8895
rect 2003 8894 2040 8895
rect 1323 8841 1364 8842
rect 261 8836 775 8837
rect 1215 8834 1364 8841
rect 1215 8814 1333 8834
rect 1353 8814 1364 8834
rect 1215 8806 1364 8814
rect 1431 8838 1790 8842
rect 1431 8833 1753 8838
rect 1431 8809 1544 8833
rect 1568 8814 1753 8833
rect 1777 8814 1790 8838
rect 1568 8809 1790 8814
rect 1431 8806 1790 8809
rect 1852 8806 1887 8843
rect 1955 8840 2055 8843
rect 1955 8836 2022 8840
rect 1955 8810 1967 8836
rect 1993 8814 2022 8836
rect 2048 8814 2055 8840
rect 1993 8810 2055 8814
rect 1955 8806 2055 8810
rect 109 8795 146 8796
rect 107 8787 147 8795
rect 107 8769 118 8787
rect 136 8769 147 8787
rect 1431 8785 1462 8806
rect 1852 8785 1888 8806
rect 1274 8784 1311 8785
rect 107 8721 147 8769
rect 1273 8775 1311 8784
rect 1273 8755 1282 8775
rect 1302 8755 1311 8775
rect 1273 8747 1311 8755
rect 1377 8779 1462 8785
rect 1487 8784 1524 8785
rect 1377 8759 1385 8779
rect 1405 8759 1462 8779
rect 1377 8751 1462 8759
rect 1486 8775 1524 8784
rect 1486 8755 1495 8775
rect 1515 8755 1524 8775
rect 1377 8750 1413 8751
rect 1486 8747 1524 8755
rect 1590 8779 1675 8785
rect 1695 8784 1732 8785
rect 1590 8759 1598 8779
rect 1618 8778 1675 8779
rect 1618 8759 1647 8778
rect 1590 8758 1647 8759
rect 1668 8758 1675 8778
rect 1590 8751 1675 8758
rect 1694 8775 1732 8784
rect 1694 8755 1703 8775
rect 1723 8755 1732 8775
rect 1590 8750 1626 8751
rect 1694 8747 1732 8755
rect 1798 8779 1942 8785
rect 1798 8759 1806 8779
rect 1826 8762 1862 8779
rect 1882 8762 1914 8779
rect 1826 8759 1914 8762
rect 1934 8759 1942 8779
rect 1798 8751 1942 8759
rect 1798 8750 1834 8751
rect 1906 8750 1942 8751
rect 2008 8784 2045 8785
rect 2008 8783 2046 8784
rect 2008 8775 2072 8783
rect 2008 8755 2017 8775
rect 2037 8761 2072 8775
rect 2092 8761 2095 8781
rect 2037 8756 2095 8761
rect 2037 8755 2072 8756
rect 418 8725 528 8739
rect 418 8722 461 8725
rect 107 8714 232 8721
rect 418 8717 422 8722
rect 107 8695 199 8714
rect 224 8695 232 8714
rect 107 8685 232 8695
rect 340 8695 422 8717
rect 451 8695 461 8722
rect 489 8698 496 8725
rect 525 8717 528 8725
rect 1274 8718 1311 8747
rect 525 8698 590 8717
rect 1275 8716 1311 8718
rect 1487 8716 1524 8747
rect 1695 8720 1732 8747
rect 2008 8743 2072 8755
rect 489 8695 590 8698
rect 340 8693 590 8695
rect 107 8665 147 8685
rect 106 8656 147 8665
rect 106 8638 116 8656
rect 134 8638 147 8656
rect 106 8629 147 8638
rect 106 8628 143 8629
rect 340 8614 377 8693
rect 418 8680 528 8693
rect 492 8624 523 8625
rect 340 8594 349 8614
rect 369 8594 377 8614
rect 340 8584 377 8594
rect 436 8614 523 8624
rect 436 8594 445 8614
rect 465 8594 523 8614
rect 436 8585 523 8594
rect 436 8584 473 8585
rect 109 8562 146 8566
rect 106 8557 146 8562
rect 106 8539 118 8557
rect 136 8539 146 8557
rect 106 8359 146 8539
rect 492 8532 523 8585
rect 553 8614 590 8693
rect 761 8690 1154 8710
rect 1174 8690 1177 8710
rect 1275 8694 1524 8716
rect 1693 8715 1734 8720
rect 2112 8717 2139 8895
rect 2790 8807 2817 8985
rect 3195 8982 3236 8987
rect 3405 8986 3654 9008
rect 3752 8992 3755 9012
rect 3775 8992 4168 9012
rect 4339 9009 4376 9088
rect 4406 9117 4437 9170
rect 4783 9163 4823 9343
rect 5161 9343 5215 9348
rect 5161 9325 5172 9343
rect 5190 9325 5215 9343
rect 8785 9364 8953 9365
rect 9193 9364 9231 9452
rect 9492 9450 9539 9452
rect 9839 9428 9879 9452
rect 19224 9457 19910 9490
rect 8785 9341 9231 9364
rect 9457 9395 9568 9408
rect 9457 9393 9499 9395
rect 9457 9373 9464 9393
rect 9483 9373 9499 9393
rect 9457 9365 9499 9373
rect 9527 9393 9568 9395
rect 9527 9373 9541 9393
rect 9560 9373 9568 9393
rect 9840 9384 9879 9428
rect 9527 9365 9568 9373
rect 9839 9368 9879 9384
rect 14168 9449 14206 9451
rect 14811 9449 15236 9451
rect 14168 9418 15245 9449
rect 14168 9416 14417 9418
rect 14573 9416 15245 9418
rect 9457 9359 9568 9365
rect 8785 9338 9229 9341
rect 8785 9336 8953 9338
rect 5161 9316 5215 9325
rect 5162 9315 5215 9316
rect 5475 9320 5585 9334
rect 5475 9317 5518 9320
rect 5475 9312 5479 9317
rect 5397 9290 5479 9312
rect 5508 9290 5518 9317
rect 5546 9293 5553 9320
rect 5582 9312 5585 9320
rect 5582 9293 5647 9312
rect 5546 9290 5647 9293
rect 5397 9288 5647 9290
rect 5165 9252 5202 9253
rect 4783 9145 4793 9163
rect 4811 9145 4823 9163
rect 4783 9140 4823 9145
rect 5161 9249 5202 9252
rect 5161 9244 5203 9249
rect 5161 9226 5174 9244
rect 5192 9226 5203 9244
rect 5161 9212 5203 9226
rect 5241 9212 5288 9216
rect 5161 9206 5288 9212
rect 5161 9177 5249 9206
rect 5278 9177 5288 9206
rect 5397 9209 5434 9288
rect 5475 9275 5585 9288
rect 5549 9219 5580 9220
rect 5397 9189 5406 9209
rect 5426 9189 5434 9209
rect 5397 9179 5434 9189
rect 5493 9209 5580 9219
rect 5493 9189 5502 9209
rect 5522 9189 5580 9209
rect 5493 9180 5580 9189
rect 5493 9179 5530 9180
rect 5161 9173 5288 9177
rect 5161 9156 5200 9173
rect 5241 9172 5288 9173
rect 4783 9136 4820 9140
rect 5161 9138 5172 9156
rect 5190 9138 5200 9156
rect 5161 9129 5200 9138
rect 5162 9128 5199 9129
rect 5549 9127 5580 9180
rect 5610 9209 5647 9288
rect 5818 9285 6211 9305
rect 6231 9285 6234 9305
rect 5818 9280 6234 9285
rect 5818 9279 6159 9280
rect 5762 9219 5793 9220
rect 5610 9189 5619 9209
rect 5639 9189 5647 9209
rect 5610 9179 5647 9189
rect 5706 9212 5793 9219
rect 5706 9209 5767 9212
rect 5706 9189 5715 9209
rect 5735 9192 5767 9209
rect 5788 9192 5793 9212
rect 5735 9189 5793 9192
rect 5706 9182 5793 9189
rect 5818 9209 5855 9279
rect 6121 9278 6158 9279
rect 5970 9219 6006 9220
rect 5818 9189 5827 9209
rect 5847 9189 5855 9209
rect 5706 9180 5762 9182
rect 5706 9179 5743 9180
rect 5818 9179 5855 9189
rect 5914 9209 6062 9219
rect 6162 9216 6258 9218
rect 5914 9189 5923 9209
rect 5943 9189 6033 9209
rect 6053 9189 6062 9209
rect 5914 9180 6062 9189
rect 6120 9209 6258 9216
rect 6120 9189 6129 9209
rect 6149 9189 6258 9209
rect 6120 9180 6258 9189
rect 5914 9179 5951 9180
rect 5970 9128 6006 9180
rect 6025 9179 6062 9180
rect 6121 9179 6158 9180
rect 5441 9126 5482 9127
rect 5333 9119 5482 9126
rect 4456 9117 4493 9118
rect 4406 9108 4493 9117
rect 4406 9088 4464 9108
rect 4484 9088 4493 9108
rect 4406 9078 4493 9088
rect 4552 9108 4589 9118
rect 4552 9088 4560 9108
rect 4580 9088 4589 9108
rect 5333 9099 5451 9119
rect 5471 9099 5482 9119
rect 5333 9091 5482 9099
rect 5549 9123 5908 9127
rect 5549 9118 5871 9123
rect 5549 9094 5662 9118
rect 5686 9099 5871 9118
rect 5895 9099 5908 9123
rect 5686 9094 5908 9099
rect 5549 9091 5908 9094
rect 5970 9091 6005 9128
rect 6073 9125 6173 9128
rect 6073 9121 6140 9125
rect 6073 9095 6085 9121
rect 6111 9099 6140 9121
rect 6166 9099 6173 9125
rect 6111 9095 6173 9099
rect 6073 9091 6173 9095
rect 4406 9077 4437 9078
rect 4401 9009 4511 9022
rect 4552 9009 4589 9088
rect 4786 9073 4823 9074
rect 4782 9064 4823 9073
rect 5549 9070 5580 9091
rect 5970 9070 6006 9091
rect 5392 9069 5429 9070
rect 5166 9066 5200 9067
rect 4782 9046 4795 9064
rect 4813 9046 4823 9064
rect 4782 9037 4823 9046
rect 5165 9057 5202 9066
rect 5165 9039 5174 9057
rect 5192 9039 5202 9057
rect 4782 9017 4822 9037
rect 5165 9029 5202 9039
rect 5391 9060 5429 9069
rect 5391 9040 5400 9060
rect 5420 9040 5429 9060
rect 5391 9032 5429 9040
rect 5495 9064 5580 9070
rect 5605 9069 5642 9070
rect 5495 9044 5503 9064
rect 5523 9044 5580 9064
rect 5495 9036 5580 9044
rect 5604 9060 5642 9069
rect 5604 9040 5613 9060
rect 5633 9040 5642 9060
rect 5495 9035 5531 9036
rect 5604 9032 5642 9040
rect 5708 9064 5793 9070
rect 5813 9069 5850 9070
rect 5708 9044 5716 9064
rect 5736 9063 5793 9064
rect 5736 9044 5765 9063
rect 5708 9043 5765 9044
rect 5786 9043 5793 9063
rect 5708 9036 5793 9043
rect 5812 9060 5850 9069
rect 5812 9040 5821 9060
rect 5841 9040 5850 9060
rect 5708 9035 5744 9036
rect 5812 9032 5850 9040
rect 5916 9064 6060 9070
rect 5916 9044 5924 9064
rect 5944 9063 6032 9064
rect 5944 9044 5975 9063
rect 5916 9043 5975 9044
rect 6000 9044 6032 9063
rect 6052 9044 6060 9064
rect 6000 9043 6060 9044
rect 5916 9036 6060 9043
rect 5916 9035 5952 9036
rect 6024 9035 6060 9036
rect 6126 9069 6163 9070
rect 6126 9068 6164 9069
rect 6126 9060 6190 9068
rect 6126 9040 6135 9060
rect 6155 9046 6190 9060
rect 6210 9046 6213 9066
rect 6155 9041 6213 9046
rect 6155 9040 6190 9041
rect 4339 9007 4589 9009
rect 4339 9004 4440 9007
rect 2857 8947 2921 8959
rect 3197 8955 3234 8982
rect 3405 8955 3442 8986
rect 3618 8984 3654 8986
rect 4339 8985 4404 9004
rect 3618 8955 3655 8984
rect 4401 8977 4404 8985
rect 4433 8977 4440 9004
rect 4468 8980 4478 9007
rect 4507 8985 4589 9007
rect 4697 9007 4822 9017
rect 4697 8988 4705 9007
rect 4730 8988 4822 9007
rect 4507 8980 4511 8985
rect 4697 8981 4822 8988
rect 4468 8977 4511 8980
rect 4401 8963 4511 8977
rect 2857 8946 2892 8947
rect 2834 8941 2892 8946
rect 2834 8921 2837 8941
rect 2857 8927 2892 8941
rect 2912 8927 2921 8947
rect 2857 8919 2921 8927
rect 2883 8918 2921 8919
rect 2884 8917 2921 8918
rect 2987 8951 3023 8952
rect 3095 8951 3131 8952
rect 2987 8943 3131 8951
rect 2987 8923 2995 8943
rect 3015 8923 3103 8943
rect 3123 8923 3131 8943
rect 2987 8917 3131 8923
rect 3197 8947 3235 8955
rect 3303 8951 3339 8952
rect 3197 8927 3206 8947
rect 3226 8927 3235 8947
rect 3197 8918 3235 8927
rect 3254 8944 3339 8951
rect 3254 8924 3261 8944
rect 3282 8943 3339 8944
rect 3282 8924 3311 8943
rect 3254 8923 3311 8924
rect 3331 8923 3339 8943
rect 3197 8917 3234 8918
rect 3254 8917 3339 8923
rect 3405 8947 3443 8955
rect 3516 8951 3552 8952
rect 3405 8927 3414 8947
rect 3434 8927 3443 8947
rect 3405 8918 3443 8927
rect 3467 8943 3552 8951
rect 3467 8923 3524 8943
rect 3544 8923 3552 8943
rect 3405 8917 3442 8918
rect 3467 8917 3552 8923
rect 3618 8947 3656 8955
rect 3618 8927 3627 8947
rect 3647 8927 3656 8947
rect 3618 8918 3656 8927
rect 4782 8933 4822 8981
rect 5166 9001 5200 9029
rect 5392 9003 5429 9032
rect 5393 9001 5429 9003
rect 5605 9001 5642 9032
rect 5166 9000 5338 9001
rect 5166 8968 5352 9000
rect 5393 8979 5642 9001
rect 5813 9000 5850 9032
rect 6126 9028 6190 9040
rect 6230 9002 6257 9180
rect 8785 9158 8812 9336
rect 8852 9298 8916 9310
rect 9192 9306 9229 9338
rect 9400 9337 9649 9359
rect 9400 9306 9437 9337
rect 9613 9335 9649 9337
rect 9613 9306 9650 9335
rect 9837 9333 10181 9368
rect 8852 9297 8887 9298
rect 8829 9292 8887 9297
rect 8829 9272 8832 9292
rect 8852 9278 8887 9292
rect 8907 9278 8916 9298
rect 8852 9270 8916 9278
rect 8878 9269 8916 9270
rect 8879 9268 8916 9269
rect 8982 9302 9018 9303
rect 9090 9302 9126 9303
rect 8982 9297 9126 9302
rect 8982 9294 9044 9297
rect 8982 9274 8990 9294
rect 9010 9277 9044 9294
rect 9067 9294 9126 9297
rect 9067 9277 9098 9294
rect 9010 9274 9098 9277
rect 9118 9274 9126 9294
rect 8982 9268 9126 9274
rect 9192 9298 9230 9306
rect 9298 9302 9334 9303
rect 9192 9278 9201 9298
rect 9221 9278 9230 9298
rect 9192 9269 9230 9278
rect 9249 9295 9334 9302
rect 9249 9275 9256 9295
rect 9277 9294 9334 9295
rect 9277 9275 9306 9294
rect 9249 9274 9306 9275
rect 9326 9274 9334 9294
rect 9192 9268 9229 9269
rect 9249 9268 9334 9274
rect 9400 9298 9438 9306
rect 9511 9302 9547 9303
rect 9400 9278 9409 9298
rect 9429 9278 9438 9298
rect 9400 9269 9438 9278
rect 9462 9294 9547 9302
rect 9462 9274 9519 9294
rect 9539 9274 9547 9294
rect 9400 9268 9437 9269
rect 9462 9268 9547 9274
rect 9613 9298 9651 9306
rect 9613 9278 9622 9298
rect 9642 9278 9651 9298
rect 9613 9269 9651 9278
rect 9613 9268 9650 9269
rect 9036 9247 9072 9268
rect 9462 9247 9493 9268
rect 8869 9243 8969 9247
rect 8869 9239 8931 9243
rect 8869 9213 8876 9239
rect 8902 9217 8931 9239
rect 8957 9217 8969 9243
rect 8902 9213 8969 9217
rect 8869 9210 8969 9213
rect 9037 9210 9072 9247
rect 9134 9244 9493 9247
rect 9134 9239 9356 9244
rect 9134 9215 9147 9239
rect 9171 9220 9356 9239
rect 9380 9220 9493 9244
rect 9171 9215 9493 9220
rect 9134 9211 9493 9215
rect 9560 9239 9709 9247
rect 9560 9219 9571 9239
rect 9591 9219 9709 9239
rect 9560 9212 9709 9219
rect 9560 9211 9601 9212
rect 8884 9158 8921 9159
rect 8980 9158 9017 9159
rect 9036 9158 9072 9210
rect 9091 9158 9128 9159
rect 8784 9149 8922 9158
rect 8784 9129 8893 9149
rect 8913 9129 8922 9149
rect 8784 9122 8922 9129
rect 8980 9149 9128 9158
rect 8980 9129 8989 9149
rect 9009 9129 9099 9149
rect 9119 9129 9128 9149
rect 8784 9120 8880 9122
rect 8980 9119 9128 9129
rect 9187 9149 9224 9159
rect 9299 9158 9336 9159
rect 9280 9156 9336 9158
rect 9187 9129 9195 9149
rect 9215 9129 9224 9149
rect 9036 9118 9072 9119
rect 6413 9076 6523 9090
rect 6413 9073 6456 9076
rect 6413 9068 6417 9073
rect 6089 9000 6257 9002
rect 5813 8994 6257 9000
rect 5166 8936 5200 8968
rect 3618 8917 3655 8918
rect 3041 8896 3077 8917
rect 3467 8896 3498 8917
rect 4782 8915 4793 8933
rect 4811 8915 4822 8933
rect 4782 8907 4822 8915
rect 5162 8927 5200 8936
rect 5162 8909 5172 8927
rect 5190 8909 5200 8927
rect 4783 8906 4820 8907
rect 5162 8903 5200 8909
rect 5318 8905 5352 8968
rect 5474 8973 5585 8979
rect 5474 8965 5515 8973
rect 5474 8945 5482 8965
rect 5501 8945 5515 8965
rect 5474 8943 5515 8945
rect 5543 8965 5585 8973
rect 5543 8945 5559 8965
rect 5578 8945 5585 8965
rect 5543 8943 5585 8945
rect 5474 8928 5585 8943
rect 5812 8974 6257 8994
rect 5812 8905 5850 8974
rect 6089 8973 6257 8974
rect 6335 9046 6417 9068
rect 6446 9046 6456 9073
rect 6484 9049 6491 9076
rect 6520 9068 6523 9076
rect 8518 9085 8629 9100
rect 8518 9083 8560 9085
rect 6520 9049 6585 9068
rect 6484 9046 6585 9049
rect 6335 9044 6585 9046
rect 6335 8965 6372 9044
rect 6413 9031 6523 9044
rect 6487 8975 6518 8976
rect 6335 8945 6344 8965
rect 6364 8945 6372 8965
rect 6335 8935 6372 8945
rect 6431 8965 6518 8975
rect 6431 8945 6440 8965
rect 6460 8945 6518 8965
rect 6431 8936 6518 8945
rect 6431 8935 6468 8936
rect 5162 8899 5199 8903
rect 2874 8892 2974 8896
rect 2874 8888 2936 8892
rect 2874 8862 2881 8888
rect 2907 8866 2936 8888
rect 2962 8866 2974 8892
rect 2907 8862 2974 8866
rect 2874 8859 2974 8862
rect 3042 8859 3077 8896
rect 3139 8893 3498 8896
rect 3139 8888 3361 8893
rect 3139 8864 3152 8888
rect 3176 8869 3361 8888
rect 3385 8869 3498 8893
rect 3176 8864 3498 8869
rect 3139 8860 3498 8864
rect 3565 8888 3714 8896
rect 5318 8894 5850 8905
rect 3565 8868 3576 8888
rect 3596 8868 3714 8888
rect 5317 8878 5850 8894
rect 6487 8883 6518 8936
rect 6548 8965 6585 9044
rect 6756 9041 7149 9061
rect 7169 9041 7172 9061
rect 8251 9056 8292 9065
rect 6756 9036 7172 9041
rect 7846 9054 8014 9055
rect 8251 9054 8260 9056
rect 6756 9035 7097 9036
rect 6700 8975 6731 8976
rect 6548 8945 6557 8965
rect 6577 8945 6585 8965
rect 6548 8935 6585 8945
rect 6644 8968 6731 8975
rect 6644 8965 6705 8968
rect 6644 8945 6653 8965
rect 6673 8948 6705 8965
rect 6726 8948 6731 8968
rect 6673 8945 6731 8948
rect 6644 8938 6731 8945
rect 6756 8965 6793 9035
rect 7059 9034 7096 9035
rect 7846 9034 8260 9054
rect 8286 9034 8292 9056
rect 8518 9063 8525 9083
rect 8544 9063 8560 9083
rect 8518 9055 8560 9063
rect 8588 9083 8629 9085
rect 8588 9063 8602 9083
rect 8621 9063 8629 9083
rect 8588 9055 8629 9063
rect 8884 9059 8921 9060
rect 9187 9059 9224 9129
rect 9249 9149 9336 9156
rect 9249 9146 9307 9149
rect 9249 9126 9254 9146
rect 9275 9129 9307 9146
rect 9327 9129 9336 9149
rect 9275 9126 9336 9129
rect 9249 9119 9336 9126
rect 9395 9149 9432 9159
rect 9395 9129 9403 9149
rect 9423 9129 9432 9149
rect 9249 9118 9280 9119
rect 8883 9058 9224 9059
rect 8518 9049 8629 9055
rect 8808 9053 9224 9058
rect 7846 9028 8292 9034
rect 7846 9026 8014 9028
rect 6908 8975 6944 8976
rect 6756 8945 6765 8965
rect 6785 8945 6793 8965
rect 6644 8936 6700 8938
rect 6644 8935 6681 8936
rect 6756 8935 6793 8945
rect 6852 8965 7000 8975
rect 7100 8972 7196 8974
rect 6852 8945 6861 8965
rect 6881 8945 6971 8965
rect 6991 8945 7000 8965
rect 6852 8936 7000 8945
rect 7058 8965 7196 8972
rect 7058 8945 7067 8965
rect 7087 8945 7196 8965
rect 7058 8936 7196 8945
rect 6852 8935 6889 8936
rect 6908 8884 6944 8936
rect 6963 8935 7000 8936
rect 7059 8935 7096 8936
rect 6379 8882 6420 8883
rect 5317 8877 5831 8878
rect 3565 8861 3714 8868
rect 6271 8875 6420 8882
rect 4154 8865 4668 8866
rect 3565 8860 3606 8861
rect 3041 8824 3077 8859
rect 2889 8807 2926 8808
rect 2985 8807 3022 8808
rect 3041 8807 3048 8824
rect 2789 8798 2927 8807
rect 2789 8778 2898 8798
rect 2918 8778 2927 8798
rect 2789 8771 2927 8778
rect 2985 8798 3048 8807
rect 2985 8778 2994 8798
rect 3014 8783 3048 8798
rect 3069 8807 3077 8824
rect 3096 8807 3133 8808
rect 3069 8798 3133 8807
rect 3069 8783 3104 8798
rect 3014 8778 3104 8783
rect 3124 8778 3133 8798
rect 2789 8769 2885 8771
rect 2985 8768 3133 8778
rect 3192 8798 3229 8808
rect 3304 8807 3341 8808
rect 3285 8805 3341 8807
rect 3192 8778 3200 8798
rect 3220 8778 3229 8798
rect 3041 8767 3077 8768
rect 1971 8715 2139 8717
rect 1693 8709 2139 8715
rect 761 8685 1177 8690
rect 1356 8688 1467 8694
rect 761 8684 1102 8685
rect 705 8624 736 8625
rect 553 8594 562 8614
rect 582 8594 590 8614
rect 553 8584 590 8594
rect 649 8617 736 8624
rect 649 8614 710 8617
rect 649 8594 658 8614
rect 678 8597 710 8614
rect 731 8597 736 8617
rect 678 8594 736 8597
rect 649 8587 736 8594
rect 761 8614 798 8684
rect 1064 8683 1101 8684
rect 1356 8680 1397 8688
rect 1356 8660 1364 8680
rect 1383 8660 1397 8680
rect 1356 8658 1397 8660
rect 1425 8680 1467 8688
rect 1425 8660 1441 8680
rect 1460 8660 1467 8680
rect 1693 8687 1699 8709
rect 1725 8689 2139 8709
rect 2889 8708 2926 8709
rect 3192 8708 3229 8778
rect 3254 8798 3341 8805
rect 3254 8795 3312 8798
rect 3254 8775 3259 8795
rect 3280 8778 3312 8795
rect 3332 8778 3341 8798
rect 3280 8775 3341 8778
rect 3254 8768 3341 8775
rect 3400 8798 3437 8808
rect 3400 8778 3408 8798
rect 3428 8778 3437 8798
rect 3254 8767 3285 8768
rect 2888 8707 3229 8708
rect 1725 8687 1734 8689
rect 1971 8688 2139 8689
rect 2813 8706 3229 8707
rect 2813 8702 3189 8706
rect 1693 8678 1734 8687
rect 2813 8682 2816 8702
rect 2836 8689 3189 8702
rect 3221 8689 3229 8706
rect 2836 8682 3229 8689
rect 3400 8699 3437 8778
rect 3467 8807 3498 8860
rect 4135 8849 4668 8865
rect 6271 8855 6389 8875
rect 6409 8855 6420 8875
rect 4135 8838 4667 8849
rect 6271 8847 6420 8855
rect 6487 8879 6846 8883
rect 6487 8874 6809 8879
rect 6487 8850 6600 8874
rect 6624 8855 6809 8874
rect 6833 8855 6846 8879
rect 6624 8850 6846 8855
rect 6487 8847 6846 8850
rect 6908 8847 6943 8884
rect 7011 8881 7111 8884
rect 7011 8877 7078 8881
rect 7011 8851 7023 8877
rect 7049 8855 7078 8877
rect 7104 8855 7111 8881
rect 7049 8851 7111 8855
rect 7011 8847 7111 8851
rect 4786 8840 4823 8844
rect 3517 8807 3554 8808
rect 3467 8798 3554 8807
rect 3467 8778 3525 8798
rect 3545 8778 3554 8798
rect 3467 8768 3554 8778
rect 3613 8798 3650 8808
rect 3613 8778 3621 8798
rect 3641 8778 3650 8798
rect 3467 8767 3498 8768
rect 3462 8699 3572 8712
rect 3613 8699 3650 8778
rect 3400 8697 3650 8699
rect 3400 8694 3501 8697
rect 3400 8675 3465 8694
rect 1425 8658 1467 8660
rect 1356 8643 1467 8658
rect 3462 8667 3465 8675
rect 3494 8667 3501 8694
rect 3529 8670 3539 8697
rect 3568 8675 3650 8697
rect 3728 8769 3896 8770
rect 4135 8769 4173 8838
rect 3728 8749 4173 8769
rect 4400 8800 4511 8815
rect 4400 8798 4442 8800
rect 4400 8778 4407 8798
rect 4426 8778 4442 8798
rect 4400 8770 4442 8778
rect 4470 8798 4511 8800
rect 4470 8778 4484 8798
rect 4503 8778 4511 8798
rect 4470 8770 4511 8778
rect 4400 8764 4511 8770
rect 4633 8775 4667 8838
rect 4785 8834 4823 8840
rect 5165 8836 5202 8837
rect 4785 8816 4795 8834
rect 4813 8816 4823 8834
rect 4785 8807 4823 8816
rect 5163 8828 5203 8836
rect 5163 8810 5174 8828
rect 5192 8810 5203 8828
rect 6487 8826 6518 8847
rect 6908 8826 6944 8847
rect 6330 8825 6367 8826
rect 4785 8775 4819 8807
rect 3728 8743 4172 8749
rect 3728 8741 3896 8743
rect 3568 8670 3572 8675
rect 3529 8667 3572 8670
rect 3462 8653 3572 8667
rect 913 8624 949 8625
rect 761 8594 770 8614
rect 790 8594 798 8614
rect 649 8585 705 8587
rect 649 8584 686 8585
rect 761 8584 798 8594
rect 857 8614 1005 8624
rect 1105 8621 1201 8623
rect 857 8594 866 8614
rect 886 8594 976 8614
rect 996 8594 1005 8614
rect 857 8585 1005 8594
rect 1063 8614 1201 8621
rect 1063 8594 1072 8614
rect 1092 8594 1201 8614
rect 1063 8585 1201 8594
rect 857 8584 894 8585
rect 913 8533 949 8585
rect 968 8584 1005 8585
rect 1064 8584 1101 8585
rect 384 8531 425 8532
rect 276 8524 425 8531
rect 276 8504 394 8524
rect 414 8504 425 8524
rect 276 8496 425 8504
rect 492 8528 851 8532
rect 492 8523 814 8528
rect 492 8499 605 8523
rect 629 8504 814 8523
rect 838 8504 851 8528
rect 629 8499 851 8504
rect 492 8496 851 8499
rect 913 8496 948 8533
rect 1016 8530 1116 8533
rect 1016 8526 1083 8530
rect 1016 8500 1028 8526
rect 1054 8504 1083 8526
rect 1109 8504 1116 8530
rect 1054 8500 1116 8504
rect 1016 8496 1116 8500
rect 492 8475 523 8496
rect 913 8475 949 8496
rect 335 8474 372 8475
rect 334 8465 372 8474
rect 334 8445 343 8465
rect 363 8445 372 8465
rect 334 8437 372 8445
rect 438 8469 523 8475
rect 548 8474 585 8475
rect 438 8449 446 8469
rect 466 8449 523 8469
rect 438 8441 523 8449
rect 547 8465 585 8474
rect 547 8445 556 8465
rect 576 8445 585 8465
rect 438 8440 474 8441
rect 547 8437 585 8445
rect 651 8469 736 8475
rect 756 8474 793 8475
rect 651 8449 659 8469
rect 679 8468 736 8469
rect 679 8449 708 8468
rect 651 8448 708 8449
rect 729 8448 736 8468
rect 651 8441 736 8448
rect 755 8465 793 8474
rect 755 8445 764 8465
rect 784 8445 793 8465
rect 651 8440 687 8441
rect 755 8437 793 8445
rect 859 8469 1003 8475
rect 859 8449 867 8469
rect 887 8466 975 8469
rect 887 8449 918 8466
rect 859 8446 918 8449
rect 941 8449 975 8466
rect 995 8449 1003 8469
rect 941 8446 1003 8449
rect 859 8441 1003 8446
rect 859 8440 895 8441
rect 967 8440 1003 8441
rect 1069 8474 1106 8475
rect 1069 8473 1107 8474
rect 1069 8465 1133 8473
rect 1069 8445 1078 8465
rect 1098 8451 1133 8465
rect 1153 8451 1156 8471
rect 1098 8446 1156 8451
rect 1098 8445 1133 8446
rect 335 8408 372 8437
rect 336 8406 372 8408
rect 548 8406 585 8437
rect 336 8384 585 8406
rect 756 8405 793 8437
rect 1069 8433 1133 8445
rect 1173 8407 1200 8585
rect 3728 8563 3755 8741
rect 3795 8703 3859 8715
rect 4135 8711 4172 8743
rect 4343 8742 4592 8764
rect 4633 8743 4819 8775
rect 4647 8742 4819 8743
rect 4343 8711 4380 8742
rect 4556 8740 4592 8742
rect 4556 8711 4593 8740
rect 4785 8714 4819 8742
rect 5163 8762 5203 8810
rect 6329 8816 6367 8825
rect 6329 8796 6338 8816
rect 6358 8796 6367 8816
rect 6329 8788 6367 8796
rect 6433 8820 6518 8826
rect 6543 8825 6580 8826
rect 6433 8800 6441 8820
rect 6461 8800 6518 8820
rect 6433 8792 6518 8800
rect 6542 8816 6580 8825
rect 6542 8796 6551 8816
rect 6571 8796 6580 8816
rect 6433 8791 6469 8792
rect 6542 8788 6580 8796
rect 6646 8820 6731 8826
rect 6751 8825 6788 8826
rect 6646 8800 6654 8820
rect 6674 8819 6731 8820
rect 6674 8800 6703 8819
rect 6646 8799 6703 8800
rect 6724 8799 6731 8819
rect 6646 8792 6731 8799
rect 6750 8816 6788 8825
rect 6750 8796 6759 8816
rect 6779 8796 6788 8816
rect 6646 8791 6682 8792
rect 6750 8788 6788 8796
rect 6854 8820 6998 8826
rect 6854 8800 6862 8820
rect 6882 8803 6918 8820
rect 6938 8803 6970 8820
rect 6882 8800 6970 8803
rect 6990 8800 6998 8820
rect 6854 8792 6998 8800
rect 6854 8791 6890 8792
rect 6962 8791 6998 8792
rect 7064 8825 7101 8826
rect 7064 8824 7102 8825
rect 7064 8816 7128 8824
rect 7064 8796 7073 8816
rect 7093 8802 7128 8816
rect 7148 8802 7151 8822
rect 7093 8797 7151 8802
rect 7093 8796 7128 8797
rect 5474 8766 5584 8780
rect 5474 8763 5517 8766
rect 5163 8755 5288 8762
rect 5474 8758 5478 8763
rect 5163 8736 5255 8755
rect 5280 8736 5288 8755
rect 5163 8726 5288 8736
rect 5396 8736 5478 8758
rect 5507 8736 5517 8763
rect 5545 8739 5552 8766
rect 5581 8758 5584 8766
rect 6330 8759 6367 8788
rect 5581 8739 5646 8758
rect 6331 8757 6367 8759
rect 6543 8757 6580 8788
rect 6751 8761 6788 8788
rect 7064 8784 7128 8796
rect 5545 8736 5646 8739
rect 5396 8734 5646 8736
rect 3795 8702 3830 8703
rect 3772 8697 3830 8702
rect 3772 8677 3775 8697
rect 3795 8683 3830 8697
rect 3850 8683 3859 8703
rect 3795 8675 3859 8683
rect 3821 8674 3859 8675
rect 3822 8673 3859 8674
rect 3925 8707 3961 8708
rect 4033 8707 4069 8708
rect 3925 8700 4069 8707
rect 3925 8699 3985 8700
rect 3925 8679 3933 8699
rect 3953 8680 3985 8699
rect 4010 8699 4069 8700
rect 4010 8680 4041 8699
rect 3953 8679 4041 8680
rect 4061 8679 4069 8699
rect 3925 8673 4069 8679
rect 4135 8703 4173 8711
rect 4241 8707 4277 8708
rect 4135 8683 4144 8703
rect 4164 8683 4173 8703
rect 4135 8674 4173 8683
rect 4192 8700 4277 8707
rect 4192 8680 4199 8700
rect 4220 8699 4277 8700
rect 4220 8680 4249 8699
rect 4192 8679 4249 8680
rect 4269 8679 4277 8699
rect 4135 8673 4172 8674
rect 4192 8673 4277 8679
rect 4343 8703 4381 8711
rect 4454 8707 4490 8708
rect 4343 8683 4352 8703
rect 4372 8683 4381 8703
rect 4343 8674 4381 8683
rect 4405 8699 4490 8707
rect 4405 8679 4462 8699
rect 4482 8679 4490 8699
rect 4343 8673 4380 8674
rect 4405 8673 4490 8679
rect 4556 8703 4594 8711
rect 4556 8683 4565 8703
rect 4585 8683 4594 8703
rect 4556 8674 4594 8683
rect 4783 8704 4820 8714
rect 5163 8706 5203 8726
rect 4783 8686 4793 8704
rect 4811 8686 4820 8704
rect 4783 8677 4820 8686
rect 5162 8697 5203 8706
rect 5162 8679 5172 8697
rect 5190 8679 5203 8697
rect 4785 8676 4819 8677
rect 4556 8673 4593 8674
rect 3979 8652 4015 8673
rect 4405 8652 4436 8673
rect 5162 8670 5203 8679
rect 5162 8669 5199 8670
rect 5396 8655 5433 8734
rect 5474 8721 5584 8734
rect 5548 8665 5579 8666
rect 3812 8648 3912 8652
rect 3812 8644 3874 8648
rect 3812 8618 3819 8644
rect 3845 8622 3874 8644
rect 3900 8622 3912 8648
rect 3845 8618 3912 8622
rect 3812 8615 3912 8618
rect 3980 8615 4015 8652
rect 4077 8649 4436 8652
rect 4077 8644 4299 8649
rect 4077 8620 4090 8644
rect 4114 8625 4299 8644
rect 4323 8625 4436 8649
rect 4114 8620 4436 8625
rect 4077 8616 4436 8620
rect 4503 8644 4652 8652
rect 4503 8624 4514 8644
rect 4534 8624 4652 8644
rect 5396 8635 5405 8655
rect 5425 8635 5433 8655
rect 5396 8625 5433 8635
rect 5492 8655 5579 8665
rect 5492 8635 5501 8655
rect 5521 8635 5579 8655
rect 5492 8626 5579 8635
rect 5492 8625 5529 8626
rect 4503 8617 4652 8624
rect 4503 8616 4544 8617
rect 3827 8563 3864 8564
rect 3923 8563 3960 8564
rect 3979 8563 4015 8615
rect 4034 8563 4071 8564
rect 3727 8554 3865 8563
rect 3322 8533 3433 8548
rect 3322 8531 3364 8533
rect 2992 8510 3097 8512
rect 2648 8502 2818 8503
rect 2992 8502 3041 8510
rect 2648 8483 3041 8502
rect 3072 8483 3097 8510
rect 3322 8511 3329 8531
rect 3348 8511 3364 8531
rect 3322 8503 3364 8511
rect 3392 8531 3433 8533
rect 3392 8511 3406 8531
rect 3425 8511 3433 8531
rect 3727 8534 3836 8554
rect 3856 8534 3865 8554
rect 3727 8527 3865 8534
rect 3923 8554 4071 8563
rect 3923 8534 3932 8554
rect 3952 8534 4042 8554
rect 4062 8534 4071 8554
rect 3727 8525 3823 8527
rect 3923 8524 4071 8534
rect 4130 8554 4167 8564
rect 4242 8563 4279 8564
rect 4223 8561 4279 8563
rect 4130 8534 4138 8554
rect 4158 8534 4167 8554
rect 3979 8523 4015 8524
rect 3392 8503 3433 8511
rect 3322 8497 3433 8503
rect 2648 8476 3097 8483
rect 2648 8474 2818 8476
rect 1498 8443 1608 8457
rect 1498 8440 1541 8443
rect 1498 8435 1502 8440
rect 1032 8405 1200 8407
rect 756 8402 1200 8405
rect 417 8378 528 8384
rect 417 8370 458 8378
rect 106 8315 145 8359
rect 417 8350 425 8370
rect 444 8350 458 8370
rect 417 8348 458 8350
rect 486 8370 528 8378
rect 486 8350 502 8370
rect 521 8350 528 8370
rect 486 8348 528 8350
rect 417 8333 528 8348
rect 754 8379 1200 8402
rect 106 8291 146 8315
rect 446 8291 493 8293
rect 754 8291 792 8379
rect 1032 8378 1200 8379
rect 1420 8413 1502 8435
rect 1531 8413 1541 8440
rect 1569 8416 1576 8443
rect 1605 8435 1608 8443
rect 1605 8416 1670 8435
rect 1569 8413 1670 8416
rect 1420 8411 1670 8413
rect 1420 8332 1457 8411
rect 1498 8398 1608 8411
rect 1572 8342 1603 8343
rect 1420 8312 1429 8332
rect 1449 8312 1457 8332
rect 1420 8302 1457 8312
rect 1516 8332 1603 8342
rect 1516 8312 1525 8332
rect 1545 8312 1603 8332
rect 1516 8303 1603 8312
rect 1516 8302 1553 8303
rect 106 8258 792 8291
rect 106 8201 145 8258
rect 754 8256 792 8258
rect 1572 8250 1603 8303
rect 1633 8332 1670 8411
rect 1841 8424 2234 8428
rect 1841 8407 1860 8424
rect 1880 8408 2234 8424
rect 2254 8408 2257 8428
rect 1880 8407 2257 8408
rect 1841 8403 2257 8407
rect 1841 8402 2182 8403
rect 1785 8342 1816 8343
rect 1633 8312 1642 8332
rect 1662 8312 1670 8332
rect 1633 8302 1670 8312
rect 1729 8335 1816 8342
rect 1729 8332 1790 8335
rect 1729 8312 1738 8332
rect 1758 8315 1790 8332
rect 1811 8315 1816 8335
rect 1758 8312 1816 8315
rect 1729 8305 1816 8312
rect 1841 8332 1878 8402
rect 2144 8401 2181 8402
rect 1993 8342 2029 8343
rect 1841 8312 1850 8332
rect 1870 8312 1878 8332
rect 1729 8303 1785 8305
rect 1729 8302 1766 8303
rect 1841 8302 1878 8312
rect 1937 8332 2085 8342
rect 2185 8339 2281 8341
rect 1937 8312 1946 8332
rect 1966 8312 2056 8332
rect 2076 8312 2085 8332
rect 1937 8303 2085 8312
rect 2143 8332 2281 8339
rect 2143 8312 2152 8332
rect 2172 8312 2281 8332
rect 2143 8303 2281 8312
rect 1937 8302 1974 8303
rect 1993 8251 2029 8303
rect 2048 8302 2085 8303
rect 2144 8302 2181 8303
rect 1464 8249 1505 8250
rect 1356 8242 1505 8249
rect 1356 8222 1474 8242
rect 1494 8222 1505 8242
rect 1356 8214 1505 8222
rect 1572 8246 1931 8250
rect 1572 8241 1894 8246
rect 1572 8217 1685 8241
rect 1709 8222 1894 8241
rect 1918 8222 1931 8246
rect 1709 8217 1931 8222
rect 1572 8214 1931 8217
rect 1993 8214 2028 8251
rect 2096 8248 2196 8251
rect 2096 8244 2163 8248
rect 2096 8218 2108 8244
rect 2134 8222 2163 8244
rect 2189 8222 2196 8248
rect 2134 8218 2196 8222
rect 2096 8214 2196 8218
rect 106 8199 154 8201
rect 106 8181 117 8199
rect 135 8181 154 8199
rect 1572 8193 1603 8214
rect 1993 8193 2029 8214
rect 1415 8192 1452 8193
rect 106 8172 154 8181
rect 107 8171 154 8172
rect 420 8176 530 8190
rect 420 8173 463 8176
rect 420 8168 424 8173
rect 342 8146 424 8168
rect 453 8146 463 8173
rect 491 8149 498 8176
rect 527 8168 530 8176
rect 1414 8183 1452 8192
rect 527 8149 592 8168
rect 1414 8163 1423 8183
rect 1443 8163 1452 8183
rect 491 8146 592 8149
rect 342 8144 592 8146
rect 110 8108 147 8109
rect 106 8105 147 8108
rect 106 8100 148 8105
rect 106 8082 119 8100
rect 137 8082 148 8100
rect 106 8068 148 8082
rect 186 8068 233 8072
rect 106 8062 233 8068
rect 106 8033 194 8062
rect 223 8033 233 8062
rect 342 8065 379 8144
rect 420 8131 530 8144
rect 494 8075 525 8076
rect 342 8045 351 8065
rect 371 8045 379 8065
rect 342 8035 379 8045
rect 438 8065 525 8075
rect 438 8045 447 8065
rect 467 8045 525 8065
rect 438 8036 525 8045
rect 438 8035 475 8036
rect 106 8029 233 8033
rect 106 8012 145 8029
rect 186 8028 233 8029
rect 106 7994 117 8012
rect 135 7994 145 8012
rect 106 7985 145 7994
rect 107 7984 144 7985
rect 494 7983 525 8036
rect 555 8065 592 8144
rect 763 8141 1156 8161
rect 1176 8141 1179 8161
rect 1414 8155 1452 8163
rect 1518 8187 1603 8193
rect 1628 8192 1665 8193
rect 1518 8167 1526 8187
rect 1546 8167 1603 8187
rect 1518 8159 1603 8167
rect 1627 8183 1665 8192
rect 1627 8163 1636 8183
rect 1656 8163 1665 8183
rect 1518 8158 1554 8159
rect 1627 8155 1665 8163
rect 1731 8187 1816 8193
rect 1836 8192 1873 8193
rect 1731 8167 1739 8187
rect 1759 8186 1816 8187
rect 1759 8167 1788 8186
rect 1731 8166 1788 8167
rect 1809 8166 1816 8186
rect 1731 8159 1816 8166
rect 1835 8183 1873 8192
rect 1835 8163 1844 8183
rect 1864 8163 1873 8183
rect 1731 8158 1767 8159
rect 1835 8155 1873 8163
rect 1939 8187 2083 8193
rect 1939 8167 1947 8187
rect 1967 8185 2055 8187
rect 1967 8167 1996 8185
rect 1939 8164 1996 8167
rect 2023 8167 2055 8185
rect 2075 8167 2083 8187
rect 2023 8164 2083 8167
rect 1939 8159 2083 8164
rect 1939 8158 1975 8159
rect 2047 8158 2083 8159
rect 2149 8192 2186 8193
rect 2149 8191 2187 8192
rect 2149 8183 2213 8191
rect 2149 8163 2158 8183
rect 2178 8169 2213 8183
rect 2233 8169 2236 8189
rect 2178 8164 2236 8169
rect 2178 8163 2213 8164
rect 763 8136 1179 8141
rect 763 8135 1104 8136
rect 707 8075 738 8076
rect 555 8045 564 8065
rect 584 8045 592 8065
rect 555 8035 592 8045
rect 651 8068 738 8075
rect 651 8065 712 8068
rect 651 8045 660 8065
rect 680 8048 712 8065
rect 733 8048 738 8068
rect 680 8045 738 8048
rect 651 8038 738 8045
rect 763 8065 800 8135
rect 1066 8134 1103 8135
rect 1415 8126 1452 8155
rect 1416 8124 1452 8126
rect 1628 8124 1665 8155
rect 1416 8102 1665 8124
rect 1836 8123 1873 8155
rect 2149 8151 2213 8163
rect 2253 8125 2280 8303
rect 2648 8296 2677 8474
rect 2717 8436 2781 8448
rect 3057 8444 3094 8476
rect 3265 8475 3514 8497
rect 3265 8444 3302 8475
rect 3478 8473 3514 8475
rect 3478 8444 3515 8473
rect 3827 8464 3864 8465
rect 4130 8464 4167 8534
rect 4192 8554 4279 8561
rect 4192 8551 4250 8554
rect 4192 8531 4197 8551
rect 4218 8534 4250 8551
rect 4270 8534 4279 8554
rect 4218 8531 4279 8534
rect 4192 8524 4279 8531
rect 4338 8554 4375 8564
rect 4338 8534 4346 8554
rect 4366 8534 4375 8554
rect 4192 8523 4223 8524
rect 3826 8463 4167 8464
rect 3751 8458 4167 8463
rect 2717 8435 2752 8436
rect 2694 8430 2752 8435
rect 2694 8410 2697 8430
rect 2717 8416 2752 8430
rect 2772 8416 2781 8436
rect 2717 8408 2781 8416
rect 2743 8407 2781 8408
rect 2744 8406 2781 8407
rect 2847 8440 2883 8441
rect 2955 8440 2991 8441
rect 2847 8432 2991 8440
rect 2847 8412 2855 8432
rect 2875 8412 2963 8432
rect 2983 8412 2991 8432
rect 2847 8406 2991 8412
rect 3057 8436 3095 8444
rect 3163 8440 3199 8441
rect 3057 8416 3066 8436
rect 3086 8416 3095 8436
rect 3057 8407 3095 8416
rect 3114 8433 3199 8440
rect 3114 8413 3121 8433
rect 3142 8432 3199 8433
rect 3142 8413 3171 8432
rect 3114 8412 3171 8413
rect 3191 8412 3199 8432
rect 3057 8406 3094 8407
rect 3114 8406 3199 8412
rect 3265 8436 3303 8444
rect 3376 8440 3412 8441
rect 3265 8416 3274 8436
rect 3294 8416 3303 8436
rect 3265 8407 3303 8416
rect 3327 8432 3412 8440
rect 3327 8412 3384 8432
rect 3404 8412 3412 8432
rect 3265 8406 3302 8407
rect 3327 8406 3412 8412
rect 3478 8436 3516 8444
rect 3751 8438 3754 8458
rect 3774 8438 4167 8458
rect 4338 8455 4375 8534
rect 4405 8563 4436 8616
rect 4786 8614 4823 8615
rect 4785 8605 4824 8614
rect 4785 8587 4795 8605
rect 4813 8587 4824 8605
rect 5165 8603 5202 8607
rect 4697 8570 4744 8571
rect 4785 8570 4824 8587
rect 4697 8566 4824 8570
rect 4455 8563 4492 8564
rect 4405 8554 4492 8563
rect 4405 8534 4463 8554
rect 4483 8534 4492 8554
rect 4405 8524 4492 8534
rect 4551 8554 4588 8564
rect 4551 8534 4559 8554
rect 4579 8534 4588 8554
rect 4405 8523 4436 8524
rect 4400 8455 4510 8468
rect 4551 8455 4588 8534
rect 4697 8537 4707 8566
rect 4736 8537 4824 8566
rect 4697 8531 4824 8537
rect 4697 8527 4744 8531
rect 4782 8517 4824 8531
rect 4782 8499 4793 8517
rect 4811 8499 4824 8517
rect 4782 8494 4824 8499
rect 4783 8491 4824 8494
rect 5162 8598 5202 8603
rect 5162 8580 5174 8598
rect 5192 8580 5202 8598
rect 4783 8490 4820 8491
rect 4338 8453 4588 8455
rect 4338 8450 4439 8453
rect 3478 8416 3487 8436
rect 3507 8416 3516 8436
rect 4338 8431 4403 8450
rect 3478 8407 3516 8416
rect 4400 8423 4403 8431
rect 4432 8423 4439 8450
rect 4467 8426 4477 8453
rect 4506 8431 4588 8453
rect 4506 8426 4510 8431
rect 4467 8423 4510 8426
rect 4400 8409 4510 8423
rect 4776 8427 4823 8428
rect 4776 8418 4824 8427
rect 3478 8406 3515 8407
rect 2901 8385 2937 8406
rect 3327 8385 3358 8406
rect 4776 8400 4795 8418
rect 4813 8400 4824 8418
rect 4776 8398 4824 8400
rect 2734 8381 2834 8385
rect 2734 8377 2796 8381
rect 2734 8351 2741 8377
rect 2767 8355 2796 8377
rect 2822 8355 2834 8381
rect 2767 8351 2834 8355
rect 2734 8348 2834 8351
rect 2902 8348 2937 8385
rect 2999 8382 3358 8385
rect 2999 8377 3221 8382
rect 2999 8353 3012 8377
rect 3036 8358 3221 8377
rect 3245 8358 3358 8382
rect 3036 8353 3358 8358
rect 2999 8349 3358 8353
rect 3425 8377 3574 8385
rect 3425 8357 3436 8377
rect 3456 8357 3574 8377
rect 3425 8350 3574 8357
rect 3425 8349 3466 8350
rect 2901 8309 2937 8348
rect 2749 8296 2786 8297
rect 2845 8296 2882 8297
rect 2901 8296 2908 8309
rect 2648 8287 2787 8296
rect 2648 8267 2758 8287
rect 2778 8267 2787 8287
rect 2648 8260 2787 8267
rect 2845 8287 2908 8296
rect 2845 8267 2854 8287
rect 2874 8271 2908 8287
rect 2931 8296 2937 8309
rect 2956 8296 2993 8297
rect 2931 8287 2993 8296
rect 2931 8271 2964 8287
rect 2874 8267 2964 8271
rect 2984 8267 2993 8287
rect 2648 8258 2745 8260
rect 2648 8257 2677 8258
rect 2845 8257 2993 8267
rect 3052 8287 3089 8297
rect 3164 8296 3201 8297
rect 3145 8294 3201 8296
rect 3052 8267 3060 8287
rect 3080 8267 3089 8287
rect 2901 8256 2937 8257
rect 2749 8197 2786 8198
rect 3052 8197 3089 8267
rect 3114 8287 3201 8294
rect 3114 8284 3172 8287
rect 3114 8264 3119 8284
rect 3140 8267 3172 8284
rect 3192 8267 3201 8287
rect 3140 8264 3201 8267
rect 3114 8257 3201 8264
rect 3260 8287 3297 8297
rect 3260 8267 3268 8287
rect 3288 8267 3297 8287
rect 3114 8256 3145 8257
rect 2748 8196 3089 8197
rect 2673 8192 3089 8196
rect 2673 8191 3050 8192
rect 2673 8171 2676 8191
rect 2696 8175 3050 8191
rect 3070 8175 3089 8192
rect 2696 8171 3089 8175
rect 3260 8188 3297 8267
rect 3327 8296 3358 8349
rect 4138 8341 4176 8343
rect 4785 8341 4824 8398
rect 4138 8308 4824 8341
rect 3377 8296 3414 8297
rect 3327 8287 3414 8296
rect 3327 8267 3385 8287
rect 3405 8267 3414 8287
rect 3327 8257 3414 8267
rect 3473 8287 3510 8297
rect 3473 8267 3481 8287
rect 3501 8267 3510 8287
rect 3327 8256 3358 8257
rect 3322 8188 3432 8201
rect 3473 8188 3510 8267
rect 3260 8186 3510 8188
rect 3260 8183 3361 8186
rect 3260 8164 3325 8183
rect 3322 8156 3325 8164
rect 3354 8156 3361 8183
rect 3389 8159 3399 8186
rect 3428 8164 3510 8186
rect 3730 8220 3898 8221
rect 4138 8220 4176 8308
rect 4437 8306 4484 8308
rect 4784 8284 4824 8308
rect 3730 8197 4176 8220
rect 4402 8251 4513 8266
rect 4402 8249 4444 8251
rect 4402 8229 4409 8249
rect 4428 8229 4444 8249
rect 4402 8221 4444 8229
rect 4472 8249 4513 8251
rect 4472 8229 4486 8249
rect 4505 8229 4513 8249
rect 4785 8240 4824 8284
rect 4472 8221 4513 8229
rect 4402 8215 4513 8221
rect 3730 8194 4174 8197
rect 3730 8192 3898 8194
rect 3428 8159 3432 8164
rect 3389 8156 3432 8159
rect 3322 8142 3432 8156
rect 2112 8123 2280 8125
rect 1833 8116 2280 8123
rect 1497 8096 1608 8102
rect 1497 8088 1538 8096
rect 915 8075 951 8076
rect 763 8045 772 8065
rect 792 8045 800 8065
rect 651 8036 707 8038
rect 651 8035 688 8036
rect 763 8035 800 8045
rect 859 8065 1007 8075
rect 1107 8072 1203 8074
rect 859 8045 868 8065
rect 888 8045 978 8065
rect 998 8045 1007 8065
rect 859 8036 1007 8045
rect 1065 8065 1203 8072
rect 1065 8045 1074 8065
rect 1094 8045 1203 8065
rect 1497 8068 1505 8088
rect 1524 8068 1538 8088
rect 1497 8066 1538 8068
rect 1566 8088 1608 8096
rect 1566 8068 1582 8088
rect 1601 8068 1608 8088
rect 1833 8089 1858 8116
rect 1889 8097 2280 8116
rect 1889 8089 1938 8097
rect 2112 8096 2280 8097
rect 1833 8087 1938 8089
rect 1566 8066 1608 8068
rect 1497 8051 1608 8066
rect 1065 8036 1203 8045
rect 859 8035 896 8036
rect 915 7984 951 8036
rect 970 8035 1007 8036
rect 1066 8035 1103 8036
rect 386 7982 427 7983
rect 278 7975 427 7982
rect 278 7955 396 7975
rect 416 7955 427 7975
rect 278 7947 427 7955
rect 494 7979 853 7983
rect 494 7974 816 7979
rect 494 7950 607 7974
rect 631 7955 816 7974
rect 840 7955 853 7979
rect 631 7950 853 7955
rect 494 7947 853 7950
rect 915 7947 950 7984
rect 1018 7981 1118 7984
rect 1018 7977 1085 7981
rect 1018 7951 1030 7977
rect 1056 7955 1085 7977
rect 1111 7955 1118 7981
rect 1056 7951 1118 7955
rect 1018 7947 1118 7951
rect 494 7926 525 7947
rect 915 7926 951 7947
rect 337 7925 374 7926
rect 111 7922 145 7923
rect 110 7913 147 7922
rect 110 7895 119 7913
rect 137 7895 147 7913
rect 110 7885 147 7895
rect 336 7916 374 7925
rect 336 7896 345 7916
rect 365 7896 374 7916
rect 336 7888 374 7896
rect 440 7920 525 7926
rect 550 7925 587 7926
rect 440 7900 448 7920
rect 468 7900 525 7920
rect 440 7892 525 7900
rect 549 7916 587 7925
rect 549 7896 558 7916
rect 578 7896 587 7916
rect 440 7891 476 7892
rect 549 7888 587 7896
rect 653 7920 738 7926
rect 758 7925 795 7926
rect 653 7900 661 7920
rect 681 7919 738 7920
rect 681 7900 710 7919
rect 653 7899 710 7900
rect 731 7899 738 7919
rect 653 7892 738 7899
rect 757 7916 795 7925
rect 757 7896 766 7916
rect 786 7896 795 7916
rect 653 7891 689 7892
rect 757 7888 795 7896
rect 861 7920 1005 7926
rect 861 7900 869 7920
rect 889 7919 977 7920
rect 889 7900 920 7919
rect 861 7899 920 7900
rect 945 7900 977 7919
rect 997 7900 1005 7920
rect 945 7899 1005 7900
rect 861 7892 1005 7899
rect 861 7891 897 7892
rect 969 7891 1005 7892
rect 1071 7925 1108 7926
rect 1071 7924 1109 7925
rect 1071 7916 1135 7924
rect 1071 7896 1080 7916
rect 1100 7902 1135 7916
rect 1155 7902 1158 7922
rect 1100 7897 1158 7902
rect 1100 7896 1135 7897
rect 111 7857 145 7885
rect 337 7859 374 7888
rect 338 7857 374 7859
rect 550 7857 587 7888
rect 111 7856 283 7857
rect 111 7824 297 7856
rect 338 7835 587 7857
rect 758 7856 795 7888
rect 1071 7884 1135 7896
rect 1175 7858 1202 8036
rect 3730 8014 3757 8192
rect 3797 8154 3861 8166
rect 4137 8162 4174 8194
rect 4345 8193 4594 8215
rect 4345 8162 4382 8193
rect 4558 8191 4594 8193
rect 4558 8162 4595 8191
rect 3797 8153 3832 8154
rect 3774 8148 3832 8153
rect 3774 8128 3777 8148
rect 3797 8134 3832 8148
rect 3852 8134 3861 8154
rect 3797 8126 3861 8134
rect 3823 8125 3861 8126
rect 3824 8124 3861 8125
rect 3927 8158 3963 8159
rect 4035 8158 4071 8159
rect 3927 8153 4071 8158
rect 3927 8150 3989 8153
rect 3927 8130 3935 8150
rect 3955 8133 3989 8150
rect 4012 8150 4071 8153
rect 4012 8133 4043 8150
rect 3955 8130 4043 8133
rect 4063 8130 4071 8150
rect 3927 8124 4071 8130
rect 4137 8154 4175 8162
rect 4243 8158 4279 8159
rect 4137 8134 4146 8154
rect 4166 8134 4175 8154
rect 4137 8125 4175 8134
rect 4194 8151 4279 8158
rect 4194 8131 4201 8151
rect 4222 8150 4279 8151
rect 4222 8131 4251 8150
rect 4194 8130 4251 8131
rect 4271 8130 4279 8150
rect 4137 8124 4174 8125
rect 4194 8124 4279 8130
rect 4345 8154 4383 8162
rect 4456 8158 4492 8159
rect 4345 8134 4354 8154
rect 4374 8134 4383 8154
rect 4345 8125 4383 8134
rect 4407 8150 4492 8158
rect 4407 8130 4464 8150
rect 4484 8130 4492 8150
rect 4345 8124 4382 8125
rect 4407 8124 4492 8130
rect 4558 8154 4596 8162
rect 4558 8134 4567 8154
rect 4587 8134 4596 8154
rect 4558 8125 4596 8134
rect 4558 8124 4595 8125
rect 3981 8103 4017 8124
rect 4407 8103 4438 8124
rect 3814 8099 3914 8103
rect 3814 8095 3876 8099
rect 3814 8069 3821 8095
rect 3847 8073 3876 8095
rect 3902 8073 3914 8099
rect 3847 8069 3914 8073
rect 3814 8066 3914 8069
rect 3982 8066 4017 8103
rect 4079 8100 4438 8103
rect 4079 8095 4301 8100
rect 4079 8071 4092 8095
rect 4116 8076 4301 8095
rect 4325 8076 4438 8100
rect 4116 8071 4438 8076
rect 4079 8067 4438 8071
rect 4505 8095 4654 8103
rect 4505 8075 4516 8095
rect 4536 8075 4654 8095
rect 4505 8068 4654 8075
rect 4505 8067 4546 8068
rect 3829 8014 3866 8015
rect 3925 8014 3962 8015
rect 3981 8014 4017 8066
rect 4036 8014 4073 8015
rect 3729 8005 3867 8014
rect 3729 7985 3838 8005
rect 3858 7985 3867 8005
rect 3729 7978 3867 7985
rect 3925 8005 4073 8014
rect 3925 7985 3934 8005
rect 3954 7985 4044 8005
rect 4064 7985 4073 8005
rect 3729 7976 3825 7978
rect 3925 7975 4073 7985
rect 4132 8005 4169 8015
rect 4244 8014 4281 8015
rect 4225 8012 4281 8014
rect 4132 7985 4140 8005
rect 4160 7985 4169 8005
rect 3981 7974 4017 7975
rect 1358 7932 1468 7946
rect 1358 7929 1401 7932
rect 1358 7924 1362 7929
rect 1034 7856 1202 7858
rect 758 7850 1202 7856
rect 111 7792 145 7824
rect 107 7783 145 7792
rect 107 7765 117 7783
rect 135 7765 145 7783
rect 107 7759 145 7765
rect 263 7761 297 7824
rect 419 7829 530 7835
rect 419 7821 460 7829
rect 419 7801 427 7821
rect 446 7801 460 7821
rect 419 7799 460 7801
rect 488 7821 530 7829
rect 488 7801 504 7821
rect 523 7801 530 7821
rect 488 7799 530 7801
rect 419 7784 530 7799
rect 757 7830 1202 7850
rect 757 7761 795 7830
rect 1034 7829 1202 7830
rect 1280 7902 1362 7924
rect 1391 7902 1401 7929
rect 1429 7905 1436 7932
rect 1465 7924 1468 7932
rect 3463 7941 3574 7956
rect 3463 7939 3505 7941
rect 1465 7905 1530 7924
rect 1429 7902 1530 7905
rect 1280 7900 1530 7902
rect 1280 7821 1317 7900
rect 1358 7887 1468 7900
rect 1432 7831 1463 7832
rect 1280 7801 1289 7821
rect 1309 7801 1317 7821
rect 1280 7791 1317 7801
rect 1376 7821 1463 7831
rect 1376 7801 1385 7821
rect 1405 7801 1463 7821
rect 1376 7792 1463 7801
rect 1376 7791 1413 7792
rect 107 7755 144 7759
rect 263 7750 795 7761
rect 262 7734 795 7750
rect 1432 7739 1463 7792
rect 1493 7821 1530 7900
rect 1701 7910 2094 7917
rect 1701 7893 1709 7910
rect 1741 7897 2094 7910
rect 2114 7897 2117 7917
rect 3196 7912 3237 7921
rect 1741 7893 2117 7897
rect 1701 7892 2117 7893
rect 2791 7910 2959 7911
rect 3196 7910 3205 7912
rect 1701 7891 2042 7892
rect 1645 7831 1676 7832
rect 1493 7801 1502 7821
rect 1522 7801 1530 7821
rect 1493 7791 1530 7801
rect 1589 7824 1676 7831
rect 1589 7821 1650 7824
rect 1589 7801 1598 7821
rect 1618 7804 1650 7821
rect 1671 7804 1676 7824
rect 1618 7801 1676 7804
rect 1589 7794 1676 7801
rect 1701 7821 1738 7891
rect 2004 7890 2041 7891
rect 2791 7890 3205 7910
rect 3231 7890 3237 7912
rect 3463 7919 3470 7939
rect 3489 7919 3505 7939
rect 3463 7911 3505 7919
rect 3533 7939 3574 7941
rect 3533 7919 3547 7939
rect 3566 7919 3574 7939
rect 3533 7911 3574 7919
rect 3829 7915 3866 7916
rect 4132 7915 4169 7985
rect 4194 8005 4281 8012
rect 4194 8002 4252 8005
rect 4194 7982 4199 8002
rect 4220 7985 4252 8002
rect 4272 7985 4281 8005
rect 4220 7982 4281 7985
rect 4194 7975 4281 7982
rect 4340 8005 4377 8015
rect 4340 7985 4348 8005
rect 4368 7985 4377 8005
rect 4194 7974 4225 7975
rect 3828 7914 4169 7915
rect 3463 7905 3574 7911
rect 3753 7909 4169 7914
rect 2791 7884 3237 7890
rect 2791 7882 2959 7884
rect 1853 7831 1889 7832
rect 1701 7801 1710 7821
rect 1730 7801 1738 7821
rect 1589 7792 1645 7794
rect 1589 7791 1626 7792
rect 1701 7791 1738 7801
rect 1797 7821 1945 7831
rect 2045 7828 2141 7830
rect 1797 7801 1806 7821
rect 1826 7816 1916 7821
rect 1826 7801 1861 7816
rect 1797 7792 1861 7801
rect 1797 7791 1834 7792
rect 1853 7775 1861 7792
rect 1882 7801 1916 7816
rect 1936 7801 1945 7821
rect 1882 7792 1945 7801
rect 2003 7821 2141 7828
rect 2003 7801 2012 7821
rect 2032 7801 2141 7821
rect 2003 7792 2141 7801
rect 1882 7775 1889 7792
rect 1908 7791 1945 7792
rect 2004 7791 2041 7792
rect 1853 7740 1889 7775
rect 1324 7738 1365 7739
rect 262 7733 776 7734
rect 1216 7731 1365 7738
rect 1216 7711 1334 7731
rect 1354 7711 1365 7731
rect 1216 7703 1365 7711
rect 1432 7735 1791 7739
rect 1432 7730 1754 7735
rect 1432 7706 1545 7730
rect 1569 7711 1754 7730
rect 1778 7711 1791 7735
rect 1569 7706 1791 7711
rect 1432 7703 1791 7706
rect 1853 7703 1888 7740
rect 1956 7737 2056 7740
rect 1956 7733 2023 7737
rect 1956 7707 1968 7733
rect 1994 7711 2023 7733
rect 2049 7711 2056 7737
rect 1994 7707 2056 7711
rect 1956 7703 2056 7707
rect 110 7692 147 7693
rect 108 7684 148 7692
rect 108 7666 119 7684
rect 137 7666 148 7684
rect 1432 7682 1463 7703
rect 1853 7682 1889 7703
rect 1275 7681 1312 7682
rect 108 7618 148 7666
rect 1274 7672 1312 7681
rect 1274 7652 1283 7672
rect 1303 7652 1312 7672
rect 1274 7644 1312 7652
rect 1378 7676 1463 7682
rect 1488 7681 1525 7682
rect 1378 7656 1386 7676
rect 1406 7656 1463 7676
rect 1378 7648 1463 7656
rect 1487 7672 1525 7681
rect 1487 7652 1496 7672
rect 1516 7652 1525 7672
rect 1378 7647 1414 7648
rect 1487 7644 1525 7652
rect 1591 7676 1676 7682
rect 1696 7681 1733 7682
rect 1591 7656 1599 7676
rect 1619 7675 1676 7676
rect 1619 7656 1648 7675
rect 1591 7655 1648 7656
rect 1669 7655 1676 7675
rect 1591 7648 1676 7655
rect 1695 7672 1733 7681
rect 1695 7652 1704 7672
rect 1724 7652 1733 7672
rect 1591 7647 1627 7648
rect 1695 7644 1733 7652
rect 1799 7676 1943 7682
rect 1799 7656 1807 7676
rect 1827 7656 1915 7676
rect 1935 7656 1943 7676
rect 1799 7648 1943 7656
rect 1799 7647 1835 7648
rect 1907 7647 1943 7648
rect 2009 7681 2046 7682
rect 2009 7680 2047 7681
rect 2009 7672 2073 7680
rect 2009 7652 2018 7672
rect 2038 7658 2073 7672
rect 2093 7658 2096 7678
rect 2038 7653 2096 7658
rect 2038 7652 2073 7653
rect 419 7622 529 7636
rect 419 7619 462 7622
rect 108 7611 233 7618
rect 419 7614 423 7619
rect 108 7592 200 7611
rect 225 7592 233 7611
rect 108 7582 233 7592
rect 341 7592 423 7614
rect 452 7592 462 7619
rect 490 7595 497 7622
rect 526 7614 529 7622
rect 1275 7615 1312 7644
rect 526 7595 591 7614
rect 1276 7613 1312 7615
rect 1488 7613 1525 7644
rect 1696 7617 1733 7644
rect 2009 7640 2073 7652
rect 490 7592 591 7595
rect 341 7590 591 7592
rect 108 7562 148 7582
rect 107 7553 148 7562
rect 107 7535 117 7553
rect 135 7535 148 7553
rect 107 7526 148 7535
rect 107 7525 144 7526
rect 341 7511 378 7590
rect 419 7577 529 7590
rect 493 7521 524 7522
rect 341 7491 350 7511
rect 370 7491 378 7511
rect 341 7481 378 7491
rect 437 7511 524 7521
rect 437 7491 446 7511
rect 466 7491 524 7511
rect 437 7482 524 7491
rect 437 7481 474 7482
rect 110 7459 147 7463
rect 107 7454 147 7459
rect 107 7436 119 7454
rect 137 7436 147 7454
rect 107 7256 147 7436
rect 493 7429 524 7482
rect 554 7511 591 7590
rect 762 7587 1155 7607
rect 1175 7587 1178 7607
rect 1276 7591 1525 7613
rect 1694 7612 1735 7617
rect 2113 7614 2140 7792
rect 2791 7704 2818 7882
rect 3196 7879 3237 7884
rect 3406 7883 3655 7905
rect 3753 7889 3756 7909
rect 3776 7889 4169 7909
rect 4340 7906 4377 7985
rect 4407 8014 4438 8067
rect 4784 8060 4824 8240
rect 5162 8400 5202 8580
rect 5548 8573 5579 8626
rect 5609 8655 5646 8734
rect 5817 8731 6210 8751
rect 6230 8731 6233 8751
rect 6331 8735 6580 8757
rect 6749 8756 6790 8761
rect 7168 8758 7195 8936
rect 7846 8848 7873 9026
rect 8251 9023 8292 9028
rect 8461 9027 8710 9049
rect 8808 9033 8811 9053
rect 8831 9033 9224 9053
rect 9395 9050 9432 9129
rect 9462 9158 9493 9211
rect 9839 9204 9879 9333
rect 10136 9309 10175 9333
rect 13760 9328 13928 9329
rect 14168 9328 14206 9416
rect 14811 9415 15246 9416
rect 14814 9392 14854 9415
rect 15166 9411 15246 9415
rect 14431 9359 14543 9377
rect 14431 9358 14474 9359
rect 10136 9307 10184 9309
rect 10136 9289 10147 9307
rect 10165 9289 10184 9307
rect 13760 9305 14206 9328
rect 14432 9357 14474 9358
rect 14432 9337 14439 9357
rect 14458 9337 14474 9357
rect 14432 9329 14474 9337
rect 14502 9357 14543 9359
rect 14502 9337 14516 9357
rect 14535 9337 14543 9357
rect 14815 9348 14854 9392
rect 15188 9367 15246 9411
rect 15190 9353 15246 9367
rect 14502 9329 14543 9337
rect 14432 9323 14543 9329
rect 13760 9302 14204 9305
rect 13760 9300 13928 9302
rect 10136 9280 10184 9289
rect 10137 9279 10184 9280
rect 10450 9284 10560 9298
rect 10450 9281 10493 9284
rect 10450 9276 10454 9281
rect 10372 9254 10454 9276
rect 10483 9254 10493 9281
rect 10521 9257 10528 9284
rect 10557 9276 10560 9284
rect 10557 9257 10622 9276
rect 10521 9254 10622 9257
rect 10372 9252 10622 9254
rect 10140 9216 10177 9217
rect 9839 9186 9849 9204
rect 9867 9186 9879 9204
rect 9839 9181 9879 9186
rect 10136 9213 10177 9216
rect 10136 9208 10178 9213
rect 10136 9190 10149 9208
rect 10167 9190 10178 9208
rect 9839 9177 9876 9181
rect 10136 9176 10178 9190
rect 10216 9176 10263 9180
rect 10136 9170 10263 9176
rect 9512 9158 9549 9159
rect 9462 9149 9549 9158
rect 9462 9129 9520 9149
rect 9540 9129 9549 9149
rect 9462 9119 9549 9129
rect 9608 9149 9645 9159
rect 9608 9129 9616 9149
rect 9636 9129 9645 9149
rect 9462 9118 9493 9119
rect 9457 9050 9567 9063
rect 9608 9050 9645 9129
rect 10136 9141 10224 9170
rect 10253 9141 10263 9170
rect 10372 9173 10409 9252
rect 10450 9239 10560 9252
rect 10524 9183 10555 9184
rect 10372 9153 10381 9173
rect 10401 9153 10409 9173
rect 10372 9143 10409 9153
rect 10468 9173 10555 9183
rect 10468 9153 10477 9173
rect 10497 9153 10555 9173
rect 10468 9144 10555 9153
rect 10468 9143 10505 9144
rect 10136 9137 10263 9141
rect 10136 9120 10175 9137
rect 10216 9136 10263 9137
rect 9842 9114 9879 9115
rect 9838 9105 9879 9114
rect 9838 9087 9851 9105
rect 9869 9087 9879 9105
rect 10136 9102 10147 9120
rect 10165 9102 10175 9120
rect 10136 9093 10175 9102
rect 10137 9092 10174 9093
rect 10524 9091 10555 9144
rect 10585 9173 10622 9252
rect 10793 9249 11186 9269
rect 11206 9249 11209 9269
rect 10793 9244 11209 9249
rect 10793 9243 11134 9244
rect 10737 9183 10768 9184
rect 10585 9153 10594 9173
rect 10614 9153 10622 9173
rect 10585 9143 10622 9153
rect 10681 9176 10768 9183
rect 10681 9173 10742 9176
rect 10681 9153 10690 9173
rect 10710 9156 10742 9173
rect 10763 9156 10768 9176
rect 10710 9153 10768 9156
rect 10681 9146 10768 9153
rect 10793 9173 10830 9243
rect 11096 9242 11133 9243
rect 10945 9183 10981 9184
rect 10793 9153 10802 9173
rect 10822 9153 10830 9173
rect 10681 9144 10737 9146
rect 10681 9143 10718 9144
rect 10793 9143 10830 9153
rect 10889 9173 11037 9183
rect 11137 9180 11233 9182
rect 10889 9153 10898 9173
rect 10918 9153 11008 9173
rect 11028 9153 11037 9173
rect 10889 9144 11037 9153
rect 11095 9173 11233 9180
rect 11095 9153 11104 9173
rect 11124 9153 11233 9173
rect 11095 9144 11233 9153
rect 10889 9143 10926 9144
rect 10945 9092 10981 9144
rect 11000 9143 11037 9144
rect 11096 9143 11133 9144
rect 10416 9090 10457 9091
rect 9838 9078 9879 9087
rect 10308 9083 10457 9090
rect 9838 9058 9878 9078
rect 9395 9048 9645 9050
rect 9395 9045 9496 9048
rect 7913 8988 7977 9000
rect 8253 8996 8290 9023
rect 8461 8996 8498 9027
rect 8674 9025 8710 9027
rect 9395 9026 9460 9045
rect 8674 8996 8711 9025
rect 9457 9018 9460 9026
rect 9489 9018 9496 9045
rect 9524 9021 9534 9048
rect 9563 9026 9645 9048
rect 9753 9048 9878 9058
rect 10308 9063 10426 9083
rect 10446 9063 10457 9083
rect 10308 9055 10457 9063
rect 10524 9087 10883 9091
rect 10524 9082 10846 9087
rect 10524 9058 10637 9082
rect 10661 9063 10846 9082
rect 10870 9063 10883 9087
rect 10661 9058 10883 9063
rect 10524 9055 10883 9058
rect 10945 9055 10980 9092
rect 11048 9089 11148 9092
rect 11048 9085 11115 9089
rect 11048 9059 11060 9085
rect 11086 9063 11115 9085
rect 11141 9063 11148 9089
rect 11086 9059 11148 9063
rect 11048 9055 11148 9059
rect 9753 9029 9761 9048
rect 9786 9029 9878 9048
rect 10524 9034 10555 9055
rect 10945 9034 10981 9055
rect 10367 9033 10404 9034
rect 10141 9030 10175 9031
rect 9563 9021 9567 9026
rect 9753 9022 9878 9029
rect 9524 9018 9567 9021
rect 9457 9004 9567 9018
rect 7913 8987 7948 8988
rect 7890 8982 7948 8987
rect 7890 8962 7893 8982
rect 7913 8968 7948 8982
rect 7968 8968 7977 8988
rect 7913 8960 7977 8968
rect 7939 8959 7977 8960
rect 7940 8958 7977 8959
rect 8043 8992 8079 8993
rect 8151 8992 8187 8993
rect 8043 8984 8187 8992
rect 8043 8964 8051 8984
rect 8071 8964 8159 8984
rect 8179 8964 8187 8984
rect 8043 8958 8187 8964
rect 8253 8988 8291 8996
rect 8359 8992 8395 8993
rect 8253 8968 8262 8988
rect 8282 8968 8291 8988
rect 8253 8959 8291 8968
rect 8310 8985 8395 8992
rect 8310 8965 8317 8985
rect 8338 8984 8395 8985
rect 8338 8965 8367 8984
rect 8310 8964 8367 8965
rect 8387 8964 8395 8984
rect 8253 8958 8290 8959
rect 8310 8958 8395 8964
rect 8461 8988 8499 8996
rect 8572 8992 8608 8993
rect 8461 8968 8470 8988
rect 8490 8968 8499 8988
rect 8461 8959 8499 8968
rect 8523 8984 8608 8992
rect 8523 8964 8580 8984
rect 8600 8964 8608 8984
rect 8461 8958 8498 8959
rect 8523 8958 8608 8964
rect 8674 8988 8712 8996
rect 8674 8968 8683 8988
rect 8703 8968 8712 8988
rect 8674 8959 8712 8968
rect 9838 8974 9878 9022
rect 10140 9021 10177 9030
rect 10140 9003 10149 9021
rect 10167 9003 10177 9021
rect 10140 8993 10177 9003
rect 10366 9024 10404 9033
rect 10366 9004 10375 9024
rect 10395 9004 10404 9024
rect 10366 8996 10404 9004
rect 10470 9028 10555 9034
rect 10580 9033 10617 9034
rect 10470 9008 10478 9028
rect 10498 9008 10555 9028
rect 10470 9000 10555 9008
rect 10579 9024 10617 9033
rect 10579 9004 10588 9024
rect 10608 9004 10617 9024
rect 10470 8999 10506 9000
rect 10579 8996 10617 9004
rect 10683 9028 10768 9034
rect 10788 9033 10825 9034
rect 10683 9008 10691 9028
rect 10711 9027 10768 9028
rect 10711 9008 10740 9027
rect 10683 9007 10740 9008
rect 10761 9007 10768 9027
rect 10683 9000 10768 9007
rect 10787 9024 10825 9033
rect 10787 9004 10796 9024
rect 10816 9004 10825 9024
rect 10683 8999 10719 9000
rect 10787 8996 10825 9004
rect 10891 9028 11035 9034
rect 10891 9008 10899 9028
rect 10919 9027 11007 9028
rect 10919 9008 10950 9027
rect 10891 9007 10950 9008
rect 10975 9008 11007 9027
rect 11027 9008 11035 9028
rect 10975 9007 11035 9008
rect 10891 9000 11035 9007
rect 10891 8999 10927 9000
rect 10999 8999 11035 9000
rect 11101 9033 11138 9034
rect 11101 9032 11139 9033
rect 11101 9024 11165 9032
rect 11101 9004 11110 9024
rect 11130 9010 11165 9024
rect 11185 9010 11188 9030
rect 11130 9005 11188 9010
rect 11130 9004 11165 9005
rect 8674 8958 8711 8959
rect 8097 8937 8133 8958
rect 8523 8937 8554 8958
rect 9838 8956 9849 8974
rect 9867 8956 9878 8974
rect 9838 8948 9878 8956
rect 10141 8965 10175 8993
rect 10367 8967 10404 8996
rect 10368 8965 10404 8967
rect 10580 8965 10617 8996
rect 10141 8964 10313 8965
rect 9839 8947 9876 8948
rect 7930 8933 8030 8937
rect 7930 8929 7992 8933
rect 7930 8903 7937 8929
rect 7963 8907 7992 8929
rect 8018 8907 8030 8933
rect 7963 8903 8030 8907
rect 7930 8900 8030 8903
rect 8098 8900 8133 8937
rect 8195 8934 8554 8937
rect 8195 8929 8417 8934
rect 8195 8905 8208 8929
rect 8232 8910 8417 8929
rect 8441 8910 8554 8934
rect 8232 8905 8554 8910
rect 8195 8901 8554 8905
rect 8621 8929 8770 8937
rect 8621 8909 8632 8929
rect 8652 8909 8770 8929
rect 8621 8902 8770 8909
rect 10141 8932 10327 8964
rect 10368 8943 10617 8965
rect 10788 8964 10825 8996
rect 11101 8992 11165 9004
rect 11205 8966 11232 9144
rect 13760 9122 13787 9300
rect 13827 9262 13891 9274
rect 14167 9270 14204 9302
rect 14375 9301 14624 9323
rect 14375 9270 14412 9301
rect 14588 9299 14624 9301
rect 14588 9270 14625 9299
rect 13827 9261 13862 9262
rect 13804 9256 13862 9261
rect 13804 9236 13807 9256
rect 13827 9242 13862 9256
rect 13882 9242 13891 9262
rect 13827 9234 13891 9242
rect 13853 9233 13891 9234
rect 13854 9232 13891 9233
rect 13957 9266 13993 9267
rect 14065 9266 14101 9267
rect 13957 9261 14101 9266
rect 13957 9258 14019 9261
rect 13957 9238 13965 9258
rect 13985 9241 14019 9258
rect 14042 9258 14101 9261
rect 14042 9241 14073 9258
rect 13985 9238 14073 9241
rect 14093 9238 14101 9258
rect 13957 9232 14101 9238
rect 14167 9262 14205 9270
rect 14273 9266 14309 9267
rect 14167 9242 14176 9262
rect 14196 9242 14205 9262
rect 14167 9233 14205 9242
rect 14224 9259 14309 9266
rect 14224 9239 14231 9259
rect 14252 9258 14309 9259
rect 14252 9239 14281 9258
rect 14224 9238 14281 9239
rect 14301 9238 14309 9258
rect 14167 9232 14204 9233
rect 14224 9232 14309 9238
rect 14375 9262 14413 9270
rect 14486 9266 14522 9267
rect 14375 9242 14384 9262
rect 14404 9242 14413 9262
rect 14375 9233 14413 9242
rect 14437 9258 14522 9266
rect 14437 9238 14494 9258
rect 14514 9238 14522 9258
rect 14375 9232 14412 9233
rect 14437 9232 14522 9238
rect 14588 9262 14626 9270
rect 14588 9242 14597 9262
rect 14617 9242 14626 9262
rect 14588 9233 14626 9242
rect 14588 9232 14625 9233
rect 14011 9211 14047 9232
rect 14437 9211 14468 9232
rect 13844 9207 13944 9211
rect 13844 9203 13906 9207
rect 13844 9177 13851 9203
rect 13877 9181 13906 9203
rect 13932 9181 13944 9207
rect 13877 9177 13944 9181
rect 13844 9174 13944 9177
rect 14012 9174 14047 9211
rect 14109 9208 14468 9211
rect 14109 9203 14331 9208
rect 14109 9179 14122 9203
rect 14146 9184 14331 9203
rect 14355 9184 14468 9208
rect 14146 9179 14468 9184
rect 14109 9175 14468 9179
rect 14535 9203 14684 9211
rect 14535 9183 14546 9203
rect 14566 9183 14684 9203
rect 14535 9176 14684 9183
rect 14535 9175 14576 9176
rect 13859 9122 13896 9123
rect 13955 9122 13992 9123
rect 14011 9122 14047 9174
rect 14066 9122 14103 9123
rect 13759 9113 13897 9122
rect 13759 9093 13868 9113
rect 13888 9093 13897 9113
rect 13759 9086 13897 9093
rect 13955 9113 14103 9122
rect 13955 9093 13964 9113
rect 13984 9093 14074 9113
rect 14094 9093 14103 9113
rect 13759 9084 13855 9086
rect 13955 9083 14103 9093
rect 14162 9113 14199 9123
rect 14274 9122 14311 9123
rect 14255 9120 14311 9122
rect 14162 9093 14170 9113
rect 14190 9093 14199 9113
rect 14011 9082 14047 9083
rect 11388 9040 11498 9054
rect 11388 9037 11431 9040
rect 11388 9032 11392 9037
rect 11064 8964 11232 8966
rect 10788 8958 11232 8964
rect 9210 8906 9724 8907
rect 8621 8901 8662 8902
rect 8097 8865 8133 8900
rect 7945 8848 7982 8849
rect 8041 8848 8078 8849
rect 8097 8848 8104 8865
rect 7845 8839 7983 8848
rect 7845 8819 7954 8839
rect 7974 8819 7983 8839
rect 7845 8812 7983 8819
rect 8041 8839 8104 8848
rect 8041 8819 8050 8839
rect 8070 8824 8104 8839
rect 8125 8848 8133 8865
rect 8152 8848 8189 8849
rect 8125 8839 8189 8848
rect 8125 8824 8160 8839
rect 8070 8819 8160 8824
rect 8180 8819 8189 8839
rect 7845 8810 7941 8812
rect 8041 8809 8189 8819
rect 8248 8839 8285 8849
rect 8360 8848 8397 8849
rect 8341 8846 8397 8848
rect 8248 8819 8256 8839
rect 8276 8819 8285 8839
rect 8097 8808 8133 8809
rect 7027 8756 7195 8758
rect 6749 8750 7195 8756
rect 5817 8726 6233 8731
rect 6412 8729 6523 8735
rect 5817 8725 6158 8726
rect 5761 8665 5792 8666
rect 5609 8635 5618 8655
rect 5638 8635 5646 8655
rect 5609 8625 5646 8635
rect 5705 8658 5792 8665
rect 5705 8655 5766 8658
rect 5705 8635 5714 8655
rect 5734 8638 5766 8655
rect 5787 8638 5792 8658
rect 5734 8635 5792 8638
rect 5705 8628 5792 8635
rect 5817 8655 5854 8725
rect 6120 8724 6157 8725
rect 6412 8721 6453 8729
rect 6412 8701 6420 8721
rect 6439 8701 6453 8721
rect 6412 8699 6453 8701
rect 6481 8721 6523 8729
rect 6481 8701 6497 8721
rect 6516 8701 6523 8721
rect 6749 8728 6755 8750
rect 6781 8730 7195 8750
rect 7945 8749 7982 8750
rect 8248 8749 8285 8819
rect 8310 8839 8397 8846
rect 8310 8836 8368 8839
rect 8310 8816 8315 8836
rect 8336 8819 8368 8836
rect 8388 8819 8397 8839
rect 8336 8816 8397 8819
rect 8310 8809 8397 8816
rect 8456 8839 8493 8849
rect 8456 8819 8464 8839
rect 8484 8819 8493 8839
rect 8310 8808 8341 8809
rect 7944 8748 8285 8749
rect 6781 8728 6790 8730
rect 7027 8729 7195 8730
rect 7869 8747 8285 8748
rect 7869 8743 8245 8747
rect 6749 8719 6790 8728
rect 7869 8723 7872 8743
rect 7892 8730 8245 8743
rect 8277 8730 8285 8747
rect 7892 8723 8285 8730
rect 8456 8740 8493 8819
rect 8523 8848 8554 8901
rect 9191 8890 9724 8906
rect 10141 8900 10175 8932
rect 10137 8891 10175 8900
rect 9191 8879 9723 8890
rect 9842 8881 9879 8885
rect 8573 8848 8610 8849
rect 8523 8839 8610 8848
rect 8523 8819 8581 8839
rect 8601 8819 8610 8839
rect 8523 8809 8610 8819
rect 8669 8839 8706 8849
rect 8669 8819 8677 8839
rect 8697 8819 8706 8839
rect 8523 8808 8554 8809
rect 8518 8740 8628 8753
rect 8669 8740 8706 8819
rect 8456 8738 8706 8740
rect 8456 8735 8557 8738
rect 8456 8716 8521 8735
rect 6481 8699 6523 8701
rect 6412 8684 6523 8699
rect 8518 8708 8521 8716
rect 8550 8708 8557 8735
rect 8585 8711 8595 8738
rect 8624 8716 8706 8738
rect 8784 8810 8952 8811
rect 9191 8810 9229 8879
rect 8784 8790 9229 8810
rect 9456 8841 9567 8856
rect 9456 8839 9498 8841
rect 9456 8819 9463 8839
rect 9482 8819 9498 8839
rect 9456 8811 9498 8819
rect 9526 8839 9567 8841
rect 9526 8819 9540 8839
rect 9559 8819 9567 8839
rect 9526 8811 9567 8819
rect 9456 8805 9567 8811
rect 9689 8816 9723 8879
rect 9841 8875 9879 8881
rect 9841 8857 9851 8875
rect 9869 8857 9879 8875
rect 10137 8873 10147 8891
rect 10165 8873 10175 8891
rect 10137 8867 10175 8873
rect 10293 8869 10327 8932
rect 10449 8937 10560 8943
rect 10449 8929 10490 8937
rect 10449 8909 10457 8929
rect 10476 8909 10490 8929
rect 10449 8907 10490 8909
rect 10518 8929 10560 8937
rect 10518 8909 10534 8929
rect 10553 8909 10560 8929
rect 10518 8907 10560 8909
rect 10449 8892 10560 8907
rect 10787 8938 11232 8958
rect 10787 8869 10825 8938
rect 11064 8937 11232 8938
rect 11310 9010 11392 9032
rect 11421 9010 11431 9037
rect 11459 9013 11466 9040
rect 11495 9032 11498 9040
rect 13493 9049 13604 9064
rect 13493 9047 13535 9049
rect 11495 9013 11560 9032
rect 11459 9010 11560 9013
rect 11310 9008 11560 9010
rect 11310 8929 11347 9008
rect 11388 8995 11498 9008
rect 11462 8939 11493 8940
rect 11310 8909 11319 8929
rect 11339 8909 11347 8929
rect 11310 8899 11347 8909
rect 11406 8929 11493 8939
rect 11406 8909 11415 8929
rect 11435 8909 11493 8929
rect 11406 8900 11493 8909
rect 11406 8899 11443 8900
rect 10137 8863 10174 8867
rect 10293 8858 10825 8869
rect 9841 8848 9879 8857
rect 9841 8816 9875 8848
rect 10292 8842 10825 8858
rect 11462 8847 11493 8900
rect 11523 8929 11560 9008
rect 11731 9005 12124 9025
rect 12144 9005 12147 9025
rect 13226 9020 13267 9029
rect 11731 9000 12147 9005
rect 12821 9018 12989 9019
rect 13226 9018 13235 9020
rect 11731 8999 12072 9000
rect 11675 8939 11706 8940
rect 11523 8909 11532 8929
rect 11552 8909 11560 8929
rect 11523 8899 11560 8909
rect 11619 8932 11706 8939
rect 11619 8929 11680 8932
rect 11619 8909 11628 8929
rect 11648 8912 11680 8929
rect 11701 8912 11706 8932
rect 11648 8909 11706 8912
rect 11619 8902 11706 8909
rect 11731 8929 11768 8999
rect 12034 8998 12071 8999
rect 12821 8998 13235 9018
rect 13261 8998 13267 9020
rect 13493 9027 13500 9047
rect 13519 9027 13535 9047
rect 13493 9019 13535 9027
rect 13563 9047 13604 9049
rect 13563 9027 13577 9047
rect 13596 9027 13604 9047
rect 13563 9019 13604 9027
rect 13859 9023 13896 9024
rect 14162 9023 14199 9093
rect 14224 9113 14311 9120
rect 14224 9110 14282 9113
rect 14224 9090 14229 9110
rect 14250 9093 14282 9110
rect 14302 9093 14311 9113
rect 14250 9090 14311 9093
rect 14224 9083 14311 9090
rect 14370 9113 14407 9123
rect 14370 9093 14378 9113
rect 14398 9093 14407 9113
rect 14224 9082 14255 9083
rect 13858 9022 14199 9023
rect 13493 9013 13604 9019
rect 13783 9017 14199 9022
rect 12821 8992 13267 8998
rect 12821 8990 12989 8992
rect 11883 8939 11919 8940
rect 11731 8909 11740 8929
rect 11760 8909 11768 8929
rect 11619 8900 11675 8902
rect 11619 8899 11656 8900
rect 11731 8899 11768 8909
rect 11827 8929 11975 8939
rect 12075 8936 12171 8938
rect 11827 8909 11836 8929
rect 11856 8909 11946 8929
rect 11966 8909 11975 8929
rect 11827 8900 11975 8909
rect 12033 8929 12171 8936
rect 12033 8909 12042 8929
rect 12062 8909 12171 8929
rect 12033 8900 12171 8909
rect 11827 8899 11864 8900
rect 11883 8848 11919 8900
rect 11938 8899 11975 8900
rect 12034 8899 12071 8900
rect 11354 8846 11395 8847
rect 10292 8841 10806 8842
rect 8784 8784 9228 8790
rect 8784 8782 8952 8784
rect 8624 8711 8628 8716
rect 8585 8708 8628 8711
rect 8518 8694 8628 8708
rect 5969 8665 6005 8666
rect 5817 8635 5826 8655
rect 5846 8635 5854 8655
rect 5705 8626 5761 8628
rect 5705 8625 5742 8626
rect 5817 8625 5854 8635
rect 5913 8655 6061 8665
rect 6161 8662 6257 8664
rect 5913 8635 5922 8655
rect 5942 8635 6032 8655
rect 6052 8635 6061 8655
rect 5913 8626 6061 8635
rect 6119 8655 6257 8662
rect 6119 8635 6128 8655
rect 6148 8635 6257 8655
rect 6119 8626 6257 8635
rect 5913 8625 5950 8626
rect 5969 8574 6005 8626
rect 6024 8625 6061 8626
rect 6120 8625 6157 8626
rect 5440 8572 5481 8573
rect 5332 8565 5481 8572
rect 5332 8545 5450 8565
rect 5470 8545 5481 8565
rect 5332 8537 5481 8545
rect 5548 8569 5907 8573
rect 5548 8564 5870 8569
rect 5548 8540 5661 8564
rect 5685 8545 5870 8564
rect 5894 8545 5907 8569
rect 5685 8540 5907 8545
rect 5548 8537 5907 8540
rect 5969 8537 6004 8574
rect 6072 8571 6172 8574
rect 6072 8567 6139 8571
rect 6072 8541 6084 8567
rect 6110 8545 6139 8567
rect 6165 8545 6172 8571
rect 6110 8541 6172 8545
rect 6072 8537 6172 8541
rect 5548 8516 5579 8537
rect 5969 8516 6005 8537
rect 5391 8515 5428 8516
rect 5390 8506 5428 8515
rect 5390 8486 5399 8506
rect 5419 8486 5428 8506
rect 5390 8478 5428 8486
rect 5494 8510 5579 8516
rect 5604 8515 5641 8516
rect 5494 8490 5502 8510
rect 5522 8490 5579 8510
rect 5494 8482 5579 8490
rect 5603 8506 5641 8515
rect 5603 8486 5612 8506
rect 5632 8486 5641 8506
rect 5494 8481 5530 8482
rect 5603 8478 5641 8486
rect 5707 8510 5792 8516
rect 5812 8515 5849 8516
rect 5707 8490 5715 8510
rect 5735 8509 5792 8510
rect 5735 8490 5764 8509
rect 5707 8489 5764 8490
rect 5785 8489 5792 8509
rect 5707 8482 5792 8489
rect 5811 8506 5849 8515
rect 5811 8486 5820 8506
rect 5840 8486 5849 8506
rect 5707 8481 5743 8482
rect 5811 8478 5849 8486
rect 5915 8510 6059 8516
rect 5915 8490 5923 8510
rect 5943 8507 6031 8510
rect 5943 8490 5974 8507
rect 5915 8487 5974 8490
rect 5997 8490 6031 8507
rect 6051 8490 6059 8510
rect 5997 8487 6059 8490
rect 5915 8482 6059 8487
rect 5915 8481 5951 8482
rect 6023 8481 6059 8482
rect 6125 8515 6162 8516
rect 6125 8514 6163 8515
rect 6125 8506 6189 8514
rect 6125 8486 6134 8506
rect 6154 8492 6189 8506
rect 6209 8492 6212 8512
rect 6154 8487 6212 8492
rect 6154 8486 6189 8487
rect 5391 8449 5428 8478
rect 5392 8447 5428 8449
rect 5604 8447 5641 8478
rect 5392 8425 5641 8447
rect 5812 8446 5849 8478
rect 6125 8474 6189 8486
rect 6229 8448 6256 8626
rect 8784 8604 8811 8782
rect 8851 8744 8915 8756
rect 9191 8752 9228 8784
rect 9399 8783 9648 8805
rect 9689 8784 9875 8816
rect 11246 8839 11395 8846
rect 11246 8819 11364 8839
rect 11384 8819 11395 8839
rect 11246 8811 11395 8819
rect 11462 8843 11821 8847
rect 11462 8838 11784 8843
rect 11462 8814 11575 8838
rect 11599 8819 11784 8838
rect 11808 8819 11821 8843
rect 11599 8814 11821 8819
rect 11462 8811 11821 8814
rect 11883 8811 11918 8848
rect 11986 8845 12086 8848
rect 11986 8841 12053 8845
rect 11986 8815 11998 8841
rect 12024 8819 12053 8841
rect 12079 8819 12086 8845
rect 12024 8815 12086 8819
rect 11986 8811 12086 8815
rect 10140 8800 10177 8801
rect 9703 8783 9875 8784
rect 9399 8752 9436 8783
rect 9612 8781 9648 8783
rect 9612 8752 9649 8781
rect 9841 8755 9875 8783
rect 10138 8792 10178 8800
rect 10138 8774 10149 8792
rect 10167 8774 10178 8792
rect 11462 8790 11493 8811
rect 11883 8790 11919 8811
rect 11305 8789 11342 8790
rect 8851 8743 8886 8744
rect 8828 8738 8886 8743
rect 8828 8718 8831 8738
rect 8851 8724 8886 8738
rect 8906 8724 8915 8744
rect 8851 8716 8915 8724
rect 8877 8715 8915 8716
rect 8878 8714 8915 8715
rect 8981 8748 9017 8749
rect 9089 8748 9125 8749
rect 8981 8741 9125 8748
rect 8981 8740 9041 8741
rect 8981 8720 8989 8740
rect 9009 8721 9041 8740
rect 9066 8740 9125 8741
rect 9066 8721 9097 8740
rect 9009 8720 9097 8721
rect 9117 8720 9125 8740
rect 8981 8714 9125 8720
rect 9191 8744 9229 8752
rect 9297 8748 9333 8749
rect 9191 8724 9200 8744
rect 9220 8724 9229 8744
rect 9191 8715 9229 8724
rect 9248 8741 9333 8748
rect 9248 8721 9255 8741
rect 9276 8740 9333 8741
rect 9276 8721 9305 8740
rect 9248 8720 9305 8721
rect 9325 8720 9333 8740
rect 9191 8714 9228 8715
rect 9248 8714 9333 8720
rect 9399 8744 9437 8752
rect 9510 8748 9546 8749
rect 9399 8724 9408 8744
rect 9428 8724 9437 8744
rect 9399 8715 9437 8724
rect 9461 8740 9546 8748
rect 9461 8720 9518 8740
rect 9538 8720 9546 8740
rect 9399 8714 9436 8715
rect 9461 8714 9546 8720
rect 9612 8744 9650 8752
rect 9612 8724 9621 8744
rect 9641 8724 9650 8744
rect 9612 8715 9650 8724
rect 9839 8745 9876 8755
rect 9839 8727 9849 8745
rect 9867 8727 9876 8745
rect 9839 8718 9876 8727
rect 10138 8726 10178 8774
rect 11304 8780 11342 8789
rect 11304 8760 11313 8780
rect 11333 8760 11342 8780
rect 11304 8752 11342 8760
rect 11408 8784 11493 8790
rect 11518 8789 11555 8790
rect 11408 8764 11416 8784
rect 11436 8764 11493 8784
rect 11408 8756 11493 8764
rect 11517 8780 11555 8789
rect 11517 8760 11526 8780
rect 11546 8760 11555 8780
rect 11408 8755 11444 8756
rect 11517 8752 11555 8760
rect 11621 8784 11706 8790
rect 11726 8789 11763 8790
rect 11621 8764 11629 8784
rect 11649 8783 11706 8784
rect 11649 8764 11678 8783
rect 11621 8763 11678 8764
rect 11699 8763 11706 8783
rect 11621 8756 11706 8763
rect 11725 8780 11763 8789
rect 11725 8760 11734 8780
rect 11754 8760 11763 8780
rect 11621 8755 11657 8756
rect 11725 8752 11763 8760
rect 11829 8784 11973 8790
rect 11829 8764 11837 8784
rect 11857 8767 11893 8784
rect 11913 8767 11945 8784
rect 11857 8764 11945 8767
rect 11965 8764 11973 8784
rect 11829 8756 11973 8764
rect 11829 8755 11865 8756
rect 11937 8755 11973 8756
rect 12039 8789 12076 8790
rect 12039 8788 12077 8789
rect 12039 8780 12103 8788
rect 12039 8760 12048 8780
rect 12068 8766 12103 8780
rect 12123 8766 12126 8786
rect 12068 8761 12126 8766
rect 12068 8760 12103 8761
rect 10449 8730 10559 8744
rect 10449 8727 10492 8730
rect 10138 8719 10263 8726
rect 10449 8722 10453 8727
rect 9841 8717 9875 8718
rect 9612 8714 9649 8715
rect 9035 8693 9071 8714
rect 9461 8693 9492 8714
rect 10138 8700 10230 8719
rect 10255 8700 10263 8719
rect 8868 8689 8968 8693
rect 8868 8685 8930 8689
rect 8868 8659 8875 8685
rect 8901 8663 8930 8685
rect 8956 8663 8968 8689
rect 8901 8659 8968 8663
rect 8868 8656 8968 8659
rect 9036 8656 9071 8693
rect 9133 8690 9492 8693
rect 9133 8685 9355 8690
rect 9133 8661 9146 8685
rect 9170 8666 9355 8685
rect 9379 8666 9492 8690
rect 9170 8661 9492 8666
rect 9133 8657 9492 8661
rect 9559 8685 9708 8693
rect 9559 8665 9570 8685
rect 9590 8665 9708 8685
rect 10138 8690 10263 8700
rect 10371 8700 10453 8722
rect 10482 8700 10492 8727
rect 10520 8703 10527 8730
rect 10556 8722 10559 8730
rect 11305 8723 11342 8752
rect 10556 8703 10621 8722
rect 11306 8721 11342 8723
rect 11518 8721 11555 8752
rect 11726 8725 11763 8752
rect 12039 8748 12103 8760
rect 10520 8700 10621 8703
rect 10371 8698 10621 8700
rect 10138 8670 10178 8690
rect 9559 8658 9708 8665
rect 10137 8661 10178 8670
rect 9559 8657 9600 8658
rect 8883 8604 8920 8605
rect 8979 8604 9016 8605
rect 9035 8604 9071 8656
rect 9090 8604 9127 8605
rect 8783 8595 8921 8604
rect 8378 8574 8489 8589
rect 8378 8572 8420 8574
rect 8048 8551 8153 8553
rect 7704 8543 7874 8544
rect 8048 8543 8097 8551
rect 7704 8524 8097 8543
rect 8128 8524 8153 8551
rect 8378 8552 8385 8572
rect 8404 8552 8420 8572
rect 8378 8544 8420 8552
rect 8448 8572 8489 8574
rect 8448 8552 8462 8572
rect 8481 8552 8489 8572
rect 8783 8575 8892 8595
rect 8912 8575 8921 8595
rect 8783 8568 8921 8575
rect 8979 8595 9127 8604
rect 8979 8575 8988 8595
rect 9008 8575 9098 8595
rect 9118 8575 9127 8595
rect 8783 8566 8879 8568
rect 8979 8565 9127 8575
rect 9186 8595 9223 8605
rect 9298 8604 9335 8605
rect 9279 8602 9335 8604
rect 9186 8575 9194 8595
rect 9214 8575 9223 8595
rect 9035 8564 9071 8565
rect 8448 8544 8489 8552
rect 8378 8538 8489 8544
rect 7704 8517 8153 8524
rect 7704 8515 7874 8517
rect 6554 8484 6664 8498
rect 6554 8481 6597 8484
rect 6554 8476 6558 8481
rect 6088 8446 6256 8448
rect 5812 8443 6256 8446
rect 5473 8419 5584 8425
rect 5473 8411 5514 8419
rect 5162 8356 5201 8400
rect 5473 8391 5481 8411
rect 5500 8391 5514 8411
rect 5473 8389 5514 8391
rect 5542 8411 5584 8419
rect 5542 8391 5558 8411
rect 5577 8391 5584 8411
rect 5542 8389 5584 8391
rect 5473 8374 5584 8389
rect 5810 8420 6256 8443
rect 5162 8332 5202 8356
rect 5502 8332 5549 8334
rect 5810 8332 5848 8420
rect 6088 8419 6256 8420
rect 6476 8454 6558 8476
rect 6587 8454 6597 8481
rect 6625 8457 6632 8484
rect 6661 8476 6664 8484
rect 6661 8457 6726 8476
rect 6625 8454 6726 8457
rect 6476 8452 6726 8454
rect 6476 8373 6513 8452
rect 6554 8439 6664 8452
rect 6628 8383 6659 8384
rect 6476 8353 6485 8373
rect 6505 8353 6513 8373
rect 6476 8343 6513 8353
rect 6572 8373 6659 8383
rect 6572 8353 6581 8373
rect 6601 8353 6659 8373
rect 6572 8344 6659 8353
rect 6572 8343 6609 8344
rect 5162 8299 5848 8332
rect 5162 8242 5201 8299
rect 5810 8297 5848 8299
rect 6628 8291 6659 8344
rect 6689 8373 6726 8452
rect 6897 8465 7290 8469
rect 6897 8448 6916 8465
rect 6936 8449 7290 8465
rect 7310 8449 7313 8469
rect 6936 8448 7313 8449
rect 6897 8444 7313 8448
rect 6897 8443 7238 8444
rect 6841 8383 6872 8384
rect 6689 8353 6698 8373
rect 6718 8353 6726 8373
rect 6689 8343 6726 8353
rect 6785 8376 6872 8383
rect 6785 8373 6846 8376
rect 6785 8353 6794 8373
rect 6814 8356 6846 8373
rect 6867 8356 6872 8376
rect 6814 8353 6872 8356
rect 6785 8346 6872 8353
rect 6897 8373 6934 8443
rect 7200 8442 7237 8443
rect 7049 8383 7085 8384
rect 6897 8353 6906 8373
rect 6926 8353 6934 8373
rect 6785 8344 6841 8346
rect 6785 8343 6822 8344
rect 6897 8343 6934 8353
rect 6993 8373 7141 8383
rect 7241 8380 7337 8382
rect 6993 8353 7002 8373
rect 7022 8353 7112 8373
rect 7132 8353 7141 8373
rect 6993 8344 7141 8353
rect 7199 8373 7337 8380
rect 7199 8353 7208 8373
rect 7228 8353 7337 8373
rect 7199 8344 7337 8353
rect 6993 8343 7030 8344
rect 7049 8292 7085 8344
rect 7104 8343 7141 8344
rect 7200 8343 7237 8344
rect 6520 8290 6561 8291
rect 6412 8283 6561 8290
rect 6412 8263 6530 8283
rect 6550 8263 6561 8283
rect 6412 8255 6561 8263
rect 6628 8287 6987 8291
rect 6628 8282 6950 8287
rect 6628 8258 6741 8282
rect 6765 8263 6950 8282
rect 6974 8263 6987 8287
rect 6765 8258 6987 8263
rect 6628 8255 6987 8258
rect 7049 8255 7084 8292
rect 7152 8289 7252 8292
rect 7152 8285 7219 8289
rect 7152 8259 7164 8285
rect 7190 8263 7219 8285
rect 7245 8263 7252 8289
rect 7190 8259 7252 8263
rect 7152 8255 7252 8259
rect 5162 8240 5210 8242
rect 5162 8222 5173 8240
rect 5191 8222 5210 8240
rect 6628 8234 6659 8255
rect 7049 8234 7085 8255
rect 6471 8233 6508 8234
rect 5162 8213 5210 8222
rect 5163 8212 5210 8213
rect 5476 8217 5586 8231
rect 5476 8214 5519 8217
rect 5476 8209 5480 8214
rect 5398 8187 5480 8209
rect 5509 8187 5519 8214
rect 5547 8190 5554 8217
rect 5583 8209 5586 8217
rect 6470 8224 6508 8233
rect 5583 8190 5648 8209
rect 6470 8204 6479 8224
rect 6499 8204 6508 8224
rect 5547 8187 5648 8190
rect 5398 8185 5648 8187
rect 5166 8149 5203 8150
rect 4784 8042 4794 8060
rect 4812 8042 4824 8060
rect 4784 8037 4824 8042
rect 5162 8146 5203 8149
rect 5162 8141 5204 8146
rect 5162 8123 5175 8141
rect 5193 8123 5204 8141
rect 5162 8109 5204 8123
rect 5242 8109 5289 8113
rect 5162 8103 5289 8109
rect 5162 8074 5250 8103
rect 5279 8074 5289 8103
rect 5398 8106 5435 8185
rect 5476 8172 5586 8185
rect 5550 8116 5581 8117
rect 5398 8086 5407 8106
rect 5427 8086 5435 8106
rect 5398 8076 5435 8086
rect 5494 8106 5581 8116
rect 5494 8086 5503 8106
rect 5523 8086 5581 8106
rect 5494 8077 5581 8086
rect 5494 8076 5531 8077
rect 5162 8070 5289 8074
rect 5162 8053 5201 8070
rect 5242 8069 5289 8070
rect 4784 8033 4821 8037
rect 5162 8035 5173 8053
rect 5191 8035 5201 8053
rect 5162 8026 5201 8035
rect 5163 8025 5200 8026
rect 5550 8024 5581 8077
rect 5611 8106 5648 8185
rect 5819 8182 6212 8202
rect 6232 8182 6235 8202
rect 6470 8196 6508 8204
rect 6574 8228 6659 8234
rect 6684 8233 6721 8234
rect 6574 8208 6582 8228
rect 6602 8208 6659 8228
rect 6574 8200 6659 8208
rect 6683 8224 6721 8233
rect 6683 8204 6692 8224
rect 6712 8204 6721 8224
rect 6574 8199 6610 8200
rect 6683 8196 6721 8204
rect 6787 8228 6872 8234
rect 6892 8233 6929 8234
rect 6787 8208 6795 8228
rect 6815 8227 6872 8228
rect 6815 8208 6844 8227
rect 6787 8207 6844 8208
rect 6865 8207 6872 8227
rect 6787 8200 6872 8207
rect 6891 8224 6929 8233
rect 6891 8204 6900 8224
rect 6920 8204 6929 8224
rect 6787 8199 6823 8200
rect 6891 8196 6929 8204
rect 6995 8228 7139 8234
rect 6995 8208 7003 8228
rect 7023 8226 7111 8228
rect 7023 8208 7052 8226
rect 6995 8205 7052 8208
rect 7079 8208 7111 8226
rect 7131 8208 7139 8228
rect 7079 8205 7139 8208
rect 6995 8200 7139 8205
rect 6995 8199 7031 8200
rect 7103 8199 7139 8200
rect 7205 8233 7242 8234
rect 7205 8232 7243 8233
rect 7205 8224 7269 8232
rect 7205 8204 7214 8224
rect 7234 8210 7269 8224
rect 7289 8210 7292 8230
rect 7234 8205 7292 8210
rect 7234 8204 7269 8205
rect 5819 8177 6235 8182
rect 5819 8176 6160 8177
rect 5763 8116 5794 8117
rect 5611 8086 5620 8106
rect 5640 8086 5648 8106
rect 5611 8076 5648 8086
rect 5707 8109 5794 8116
rect 5707 8106 5768 8109
rect 5707 8086 5716 8106
rect 5736 8089 5768 8106
rect 5789 8089 5794 8109
rect 5736 8086 5794 8089
rect 5707 8079 5794 8086
rect 5819 8106 5856 8176
rect 6122 8175 6159 8176
rect 6471 8167 6508 8196
rect 6472 8165 6508 8167
rect 6684 8165 6721 8196
rect 6472 8143 6721 8165
rect 6892 8164 6929 8196
rect 7205 8192 7269 8204
rect 7309 8166 7336 8344
rect 7704 8337 7733 8515
rect 7773 8477 7837 8489
rect 8113 8485 8150 8517
rect 8321 8516 8570 8538
rect 8321 8485 8358 8516
rect 8534 8514 8570 8516
rect 8534 8485 8571 8514
rect 8883 8505 8920 8506
rect 9186 8505 9223 8575
rect 9248 8595 9335 8602
rect 9248 8592 9306 8595
rect 9248 8572 9253 8592
rect 9274 8575 9306 8592
rect 9326 8575 9335 8595
rect 9274 8572 9335 8575
rect 9248 8565 9335 8572
rect 9394 8595 9431 8605
rect 9394 8575 9402 8595
rect 9422 8575 9431 8595
rect 9248 8564 9279 8565
rect 8882 8504 9223 8505
rect 8807 8499 9223 8504
rect 7773 8476 7808 8477
rect 7750 8471 7808 8476
rect 7750 8451 7753 8471
rect 7773 8457 7808 8471
rect 7828 8457 7837 8477
rect 7773 8449 7837 8457
rect 7799 8448 7837 8449
rect 7800 8447 7837 8448
rect 7903 8481 7939 8482
rect 8011 8481 8047 8482
rect 7903 8473 8047 8481
rect 7903 8453 7911 8473
rect 7931 8453 8019 8473
rect 8039 8453 8047 8473
rect 7903 8447 8047 8453
rect 8113 8477 8151 8485
rect 8219 8481 8255 8482
rect 8113 8457 8122 8477
rect 8142 8457 8151 8477
rect 8113 8448 8151 8457
rect 8170 8474 8255 8481
rect 8170 8454 8177 8474
rect 8198 8473 8255 8474
rect 8198 8454 8227 8473
rect 8170 8453 8227 8454
rect 8247 8453 8255 8473
rect 8113 8447 8150 8448
rect 8170 8447 8255 8453
rect 8321 8477 8359 8485
rect 8432 8481 8468 8482
rect 8321 8457 8330 8477
rect 8350 8457 8359 8477
rect 8321 8448 8359 8457
rect 8383 8473 8468 8481
rect 8383 8453 8440 8473
rect 8460 8453 8468 8473
rect 8321 8447 8358 8448
rect 8383 8447 8468 8453
rect 8534 8477 8572 8485
rect 8807 8479 8810 8499
rect 8830 8479 9223 8499
rect 9394 8496 9431 8575
rect 9461 8604 9492 8657
rect 9842 8655 9879 8656
rect 9841 8646 9880 8655
rect 9841 8628 9851 8646
rect 9869 8628 9880 8646
rect 10137 8643 10147 8661
rect 10165 8643 10178 8661
rect 10137 8634 10178 8643
rect 10137 8633 10174 8634
rect 9753 8611 9800 8612
rect 9841 8611 9880 8628
rect 9753 8607 9880 8611
rect 9511 8604 9548 8605
rect 9461 8595 9548 8604
rect 9461 8575 9519 8595
rect 9539 8575 9548 8595
rect 9461 8565 9548 8575
rect 9607 8595 9644 8605
rect 9607 8575 9615 8595
rect 9635 8575 9644 8595
rect 9461 8564 9492 8565
rect 9456 8496 9566 8509
rect 9607 8496 9644 8575
rect 9753 8578 9763 8607
rect 9792 8578 9880 8607
rect 10371 8619 10408 8698
rect 10449 8685 10559 8698
rect 10523 8629 10554 8630
rect 10371 8599 10380 8619
rect 10400 8599 10408 8619
rect 10371 8589 10408 8599
rect 10467 8619 10554 8629
rect 10467 8599 10476 8619
rect 10496 8599 10554 8619
rect 10467 8590 10554 8599
rect 10467 8589 10504 8590
rect 9753 8572 9880 8578
rect 9753 8568 9800 8572
rect 9838 8558 9880 8572
rect 10140 8567 10177 8571
rect 9838 8540 9849 8558
rect 9867 8540 9880 8558
rect 9838 8535 9880 8540
rect 9839 8532 9880 8535
rect 10137 8562 10177 8567
rect 10137 8544 10149 8562
rect 10167 8544 10177 8562
rect 9839 8531 9876 8532
rect 9394 8494 9644 8496
rect 9394 8491 9495 8494
rect 8534 8457 8543 8477
rect 8563 8457 8572 8477
rect 9394 8472 9459 8491
rect 8534 8448 8572 8457
rect 9456 8464 9459 8472
rect 9488 8464 9495 8491
rect 9523 8467 9533 8494
rect 9562 8472 9644 8494
rect 9562 8467 9566 8472
rect 9523 8464 9566 8467
rect 9456 8450 9566 8464
rect 9832 8468 9879 8469
rect 9832 8459 9880 8468
rect 8534 8447 8571 8448
rect 7957 8426 7993 8447
rect 8383 8426 8414 8447
rect 9832 8441 9851 8459
rect 9869 8441 9880 8459
rect 9832 8439 9880 8441
rect 7790 8422 7890 8426
rect 7790 8418 7852 8422
rect 7790 8392 7797 8418
rect 7823 8396 7852 8418
rect 7878 8396 7890 8422
rect 7823 8392 7890 8396
rect 7790 8389 7890 8392
rect 7958 8389 7993 8426
rect 8055 8423 8414 8426
rect 8055 8418 8277 8423
rect 8055 8394 8068 8418
rect 8092 8399 8277 8418
rect 8301 8399 8414 8423
rect 8092 8394 8414 8399
rect 8055 8390 8414 8394
rect 8481 8418 8630 8426
rect 8481 8398 8492 8418
rect 8512 8398 8630 8418
rect 8481 8391 8630 8398
rect 8481 8390 8522 8391
rect 7957 8350 7993 8389
rect 7805 8337 7842 8338
rect 7901 8337 7938 8338
rect 7957 8337 7964 8350
rect 7704 8328 7843 8337
rect 7704 8308 7814 8328
rect 7834 8308 7843 8328
rect 7704 8301 7843 8308
rect 7901 8328 7964 8337
rect 7901 8308 7910 8328
rect 7930 8312 7964 8328
rect 7987 8337 7993 8350
rect 8012 8337 8049 8338
rect 7987 8328 8049 8337
rect 7987 8312 8020 8328
rect 7930 8308 8020 8312
rect 8040 8308 8049 8328
rect 7704 8299 7801 8301
rect 7704 8298 7733 8299
rect 7901 8298 8049 8308
rect 8108 8328 8145 8338
rect 8220 8337 8257 8338
rect 8201 8335 8257 8337
rect 8108 8308 8116 8328
rect 8136 8308 8145 8328
rect 7957 8297 7993 8298
rect 7805 8238 7842 8239
rect 8108 8238 8145 8308
rect 8170 8328 8257 8335
rect 8170 8325 8228 8328
rect 8170 8305 8175 8325
rect 8196 8308 8228 8325
rect 8248 8308 8257 8328
rect 8196 8305 8257 8308
rect 8170 8298 8257 8305
rect 8316 8328 8353 8338
rect 8316 8308 8324 8328
rect 8344 8308 8353 8328
rect 8170 8297 8201 8298
rect 7804 8237 8145 8238
rect 7729 8233 8145 8237
rect 7729 8232 8106 8233
rect 7729 8212 7732 8232
rect 7752 8216 8106 8232
rect 8126 8216 8145 8233
rect 7752 8212 8145 8216
rect 8316 8229 8353 8308
rect 8383 8337 8414 8390
rect 9194 8382 9232 8384
rect 9841 8382 9880 8439
rect 9194 8349 9880 8382
rect 8433 8337 8470 8338
rect 8383 8328 8470 8337
rect 8383 8308 8441 8328
rect 8461 8308 8470 8328
rect 8383 8298 8470 8308
rect 8529 8328 8566 8338
rect 8529 8308 8537 8328
rect 8557 8308 8566 8328
rect 8383 8297 8414 8298
rect 8378 8229 8488 8242
rect 8529 8229 8566 8308
rect 8316 8227 8566 8229
rect 8316 8224 8417 8227
rect 8316 8205 8381 8224
rect 8378 8197 8381 8205
rect 8410 8197 8417 8224
rect 8445 8200 8455 8227
rect 8484 8205 8566 8227
rect 8786 8261 8954 8262
rect 9194 8261 9232 8349
rect 9493 8347 9540 8349
rect 9840 8325 9880 8349
rect 8786 8238 9232 8261
rect 9458 8292 9569 8307
rect 9458 8290 9500 8292
rect 9458 8270 9465 8290
rect 9484 8270 9500 8290
rect 9458 8262 9500 8270
rect 9528 8290 9569 8292
rect 9528 8270 9542 8290
rect 9561 8270 9569 8290
rect 9841 8281 9880 8325
rect 9528 8262 9569 8270
rect 9458 8256 9569 8262
rect 8786 8235 9230 8238
rect 8786 8233 8954 8235
rect 8484 8200 8488 8205
rect 8445 8197 8488 8200
rect 8378 8183 8488 8197
rect 7168 8164 7336 8166
rect 6889 8157 7336 8164
rect 6553 8137 6664 8143
rect 6553 8129 6594 8137
rect 5971 8116 6007 8117
rect 5819 8086 5828 8106
rect 5848 8086 5856 8106
rect 5707 8077 5763 8079
rect 5707 8076 5744 8077
rect 5819 8076 5856 8086
rect 5915 8106 6063 8116
rect 6163 8113 6259 8115
rect 5915 8086 5924 8106
rect 5944 8086 6034 8106
rect 6054 8086 6063 8106
rect 5915 8077 6063 8086
rect 6121 8106 6259 8113
rect 6121 8086 6130 8106
rect 6150 8086 6259 8106
rect 6553 8109 6561 8129
rect 6580 8109 6594 8129
rect 6553 8107 6594 8109
rect 6622 8129 6664 8137
rect 6622 8109 6638 8129
rect 6657 8109 6664 8129
rect 6889 8130 6914 8157
rect 6945 8138 7336 8157
rect 6945 8130 6994 8138
rect 7168 8137 7336 8138
rect 6889 8128 6994 8130
rect 6622 8107 6664 8109
rect 6553 8092 6664 8107
rect 6121 8077 6259 8086
rect 5915 8076 5952 8077
rect 5971 8025 6007 8077
rect 6026 8076 6063 8077
rect 6122 8076 6159 8077
rect 5442 8023 5483 8024
rect 5334 8016 5483 8023
rect 4457 8014 4494 8015
rect 4407 8005 4494 8014
rect 4407 7985 4465 8005
rect 4485 7985 4494 8005
rect 4407 7975 4494 7985
rect 4553 8005 4590 8015
rect 4553 7985 4561 8005
rect 4581 7985 4590 8005
rect 5334 7996 5452 8016
rect 5472 7996 5483 8016
rect 5334 7988 5483 7996
rect 5550 8020 5909 8024
rect 5550 8015 5872 8020
rect 5550 7991 5663 8015
rect 5687 7996 5872 8015
rect 5896 7996 5909 8020
rect 5687 7991 5909 7996
rect 5550 7988 5909 7991
rect 5971 7988 6006 8025
rect 6074 8022 6174 8025
rect 6074 8018 6141 8022
rect 6074 7992 6086 8018
rect 6112 7996 6141 8018
rect 6167 7996 6174 8022
rect 6112 7992 6174 7996
rect 6074 7988 6174 7992
rect 4407 7974 4438 7975
rect 4402 7906 4512 7919
rect 4553 7906 4590 7985
rect 4787 7970 4824 7971
rect 4783 7961 4824 7970
rect 5550 7967 5581 7988
rect 5971 7967 6007 7988
rect 5393 7966 5430 7967
rect 5167 7963 5201 7964
rect 4783 7943 4796 7961
rect 4814 7943 4824 7961
rect 4783 7934 4824 7943
rect 5166 7954 5203 7963
rect 5166 7936 5175 7954
rect 5193 7936 5203 7954
rect 4783 7914 4823 7934
rect 5166 7926 5203 7936
rect 5392 7957 5430 7966
rect 5392 7937 5401 7957
rect 5421 7937 5430 7957
rect 5392 7929 5430 7937
rect 5496 7961 5581 7967
rect 5606 7966 5643 7967
rect 5496 7941 5504 7961
rect 5524 7941 5581 7961
rect 5496 7933 5581 7941
rect 5605 7957 5643 7966
rect 5605 7937 5614 7957
rect 5634 7937 5643 7957
rect 5496 7932 5532 7933
rect 5605 7929 5643 7937
rect 5709 7961 5794 7967
rect 5814 7966 5851 7967
rect 5709 7941 5717 7961
rect 5737 7960 5794 7961
rect 5737 7941 5766 7960
rect 5709 7940 5766 7941
rect 5787 7940 5794 7960
rect 5709 7933 5794 7940
rect 5813 7957 5851 7966
rect 5813 7937 5822 7957
rect 5842 7937 5851 7957
rect 5709 7932 5745 7933
rect 5813 7929 5851 7937
rect 5917 7961 6061 7967
rect 5917 7941 5925 7961
rect 5945 7960 6033 7961
rect 5945 7941 5976 7960
rect 5917 7940 5976 7941
rect 6001 7941 6033 7960
rect 6053 7941 6061 7961
rect 6001 7940 6061 7941
rect 5917 7933 6061 7940
rect 5917 7932 5953 7933
rect 6025 7932 6061 7933
rect 6127 7966 6164 7967
rect 6127 7965 6165 7966
rect 6127 7957 6191 7965
rect 6127 7937 6136 7957
rect 6156 7943 6191 7957
rect 6211 7943 6214 7963
rect 6156 7938 6214 7943
rect 6156 7937 6191 7938
rect 4340 7904 4590 7906
rect 4340 7901 4441 7904
rect 2858 7844 2922 7856
rect 3198 7852 3235 7879
rect 3406 7852 3443 7883
rect 3619 7881 3655 7883
rect 4340 7882 4405 7901
rect 3619 7852 3656 7881
rect 4402 7874 4405 7882
rect 4434 7874 4441 7901
rect 4469 7877 4479 7904
rect 4508 7882 4590 7904
rect 4698 7904 4823 7914
rect 4698 7885 4706 7904
rect 4731 7885 4823 7904
rect 4508 7877 4512 7882
rect 4698 7878 4823 7885
rect 4469 7874 4512 7877
rect 4402 7860 4512 7874
rect 2858 7843 2893 7844
rect 2835 7838 2893 7843
rect 2835 7818 2838 7838
rect 2858 7824 2893 7838
rect 2913 7824 2922 7844
rect 2858 7816 2922 7824
rect 2884 7815 2922 7816
rect 2885 7814 2922 7815
rect 2988 7848 3024 7849
rect 3096 7848 3132 7849
rect 2988 7840 3132 7848
rect 2988 7820 2996 7840
rect 3016 7837 3104 7840
rect 3016 7820 3048 7837
rect 3068 7820 3104 7837
rect 3124 7820 3132 7840
rect 2988 7814 3132 7820
rect 3198 7844 3236 7852
rect 3304 7848 3340 7849
rect 3198 7824 3207 7844
rect 3227 7824 3236 7844
rect 3198 7815 3236 7824
rect 3255 7841 3340 7848
rect 3255 7821 3262 7841
rect 3283 7840 3340 7841
rect 3283 7821 3312 7840
rect 3255 7820 3312 7821
rect 3332 7820 3340 7840
rect 3198 7814 3235 7815
rect 3255 7814 3340 7820
rect 3406 7844 3444 7852
rect 3517 7848 3553 7849
rect 3406 7824 3415 7844
rect 3435 7824 3444 7844
rect 3406 7815 3444 7824
rect 3468 7840 3553 7848
rect 3468 7820 3525 7840
rect 3545 7820 3553 7840
rect 3406 7814 3443 7815
rect 3468 7814 3553 7820
rect 3619 7844 3657 7852
rect 3619 7824 3628 7844
rect 3648 7824 3657 7844
rect 3619 7815 3657 7824
rect 4783 7830 4823 7878
rect 5167 7898 5201 7926
rect 5393 7900 5430 7929
rect 5394 7898 5430 7900
rect 5606 7898 5643 7929
rect 5167 7897 5339 7898
rect 5167 7865 5353 7897
rect 5394 7876 5643 7898
rect 5814 7897 5851 7929
rect 6127 7925 6191 7937
rect 6231 7899 6258 8077
rect 8786 8055 8813 8233
rect 8853 8195 8917 8207
rect 9193 8203 9230 8235
rect 9401 8234 9650 8256
rect 9401 8203 9438 8234
rect 9614 8232 9650 8234
rect 9614 8203 9651 8232
rect 8853 8194 8888 8195
rect 8830 8189 8888 8194
rect 8830 8169 8833 8189
rect 8853 8175 8888 8189
rect 8908 8175 8917 8195
rect 8853 8167 8917 8175
rect 8879 8166 8917 8167
rect 8880 8165 8917 8166
rect 8983 8199 9019 8200
rect 9091 8199 9127 8200
rect 8983 8194 9127 8199
rect 8983 8191 9045 8194
rect 8983 8171 8991 8191
rect 9011 8174 9045 8191
rect 9068 8191 9127 8194
rect 9068 8174 9099 8191
rect 9011 8171 9099 8174
rect 9119 8171 9127 8191
rect 8983 8165 9127 8171
rect 9193 8195 9231 8203
rect 9299 8199 9335 8200
rect 9193 8175 9202 8195
rect 9222 8175 9231 8195
rect 9193 8166 9231 8175
rect 9250 8192 9335 8199
rect 9250 8172 9257 8192
rect 9278 8191 9335 8192
rect 9278 8172 9307 8191
rect 9250 8171 9307 8172
rect 9327 8171 9335 8191
rect 9193 8165 9230 8166
rect 9250 8165 9335 8171
rect 9401 8195 9439 8203
rect 9512 8199 9548 8200
rect 9401 8175 9410 8195
rect 9430 8175 9439 8195
rect 9401 8166 9439 8175
rect 9463 8191 9548 8199
rect 9463 8171 9520 8191
rect 9540 8171 9548 8191
rect 9401 8165 9438 8166
rect 9463 8165 9548 8171
rect 9614 8195 9652 8203
rect 9614 8175 9623 8195
rect 9643 8175 9652 8195
rect 9614 8166 9652 8175
rect 9614 8165 9651 8166
rect 9037 8144 9073 8165
rect 9463 8144 9494 8165
rect 8870 8140 8970 8144
rect 8870 8136 8932 8140
rect 8870 8110 8877 8136
rect 8903 8114 8932 8136
rect 8958 8114 8970 8140
rect 8903 8110 8970 8114
rect 8870 8107 8970 8110
rect 9038 8107 9073 8144
rect 9135 8141 9494 8144
rect 9135 8136 9357 8141
rect 9135 8112 9148 8136
rect 9172 8117 9357 8136
rect 9381 8117 9494 8141
rect 9172 8112 9494 8117
rect 9135 8108 9494 8112
rect 9561 8136 9710 8144
rect 9561 8116 9572 8136
rect 9592 8116 9710 8136
rect 9561 8109 9710 8116
rect 9561 8108 9602 8109
rect 8885 8055 8922 8056
rect 8981 8055 9018 8056
rect 9037 8055 9073 8107
rect 9092 8055 9129 8056
rect 8785 8046 8923 8055
rect 8785 8026 8894 8046
rect 8914 8026 8923 8046
rect 8785 8019 8923 8026
rect 8981 8046 9129 8055
rect 8981 8026 8990 8046
rect 9010 8026 9100 8046
rect 9120 8026 9129 8046
rect 8785 8017 8881 8019
rect 8981 8016 9129 8026
rect 9188 8046 9225 8056
rect 9300 8055 9337 8056
rect 9281 8053 9337 8055
rect 9188 8026 9196 8046
rect 9216 8026 9225 8046
rect 9037 8015 9073 8016
rect 6414 7973 6524 7987
rect 6414 7970 6457 7973
rect 6414 7965 6418 7970
rect 6090 7897 6258 7899
rect 5814 7891 6258 7897
rect 5167 7833 5201 7865
rect 3619 7814 3656 7815
rect 3042 7793 3078 7814
rect 3468 7793 3499 7814
rect 4783 7812 4794 7830
rect 4812 7812 4823 7830
rect 4783 7804 4823 7812
rect 5163 7824 5201 7833
rect 5163 7806 5173 7824
rect 5191 7806 5201 7824
rect 4784 7803 4821 7804
rect 5163 7800 5201 7806
rect 5319 7802 5353 7865
rect 5475 7870 5586 7876
rect 5475 7862 5516 7870
rect 5475 7842 5483 7862
rect 5502 7842 5516 7862
rect 5475 7840 5516 7842
rect 5544 7862 5586 7870
rect 5544 7842 5560 7862
rect 5579 7842 5586 7862
rect 5544 7840 5586 7842
rect 5475 7825 5586 7840
rect 5813 7871 6258 7891
rect 5813 7802 5851 7871
rect 6090 7870 6258 7871
rect 6336 7943 6418 7965
rect 6447 7943 6457 7970
rect 6485 7946 6492 7973
rect 6521 7965 6524 7973
rect 8519 7982 8630 7997
rect 8519 7980 8561 7982
rect 6521 7946 6586 7965
rect 6485 7943 6586 7946
rect 6336 7941 6586 7943
rect 6336 7862 6373 7941
rect 6414 7928 6524 7941
rect 6488 7872 6519 7873
rect 6336 7842 6345 7862
rect 6365 7842 6373 7862
rect 6336 7832 6373 7842
rect 6432 7862 6519 7872
rect 6432 7842 6441 7862
rect 6461 7842 6519 7862
rect 6432 7833 6519 7842
rect 6432 7832 6469 7833
rect 5163 7796 5200 7800
rect 2875 7789 2975 7793
rect 2875 7785 2937 7789
rect 2875 7759 2882 7785
rect 2908 7763 2937 7785
rect 2963 7763 2975 7789
rect 2908 7759 2975 7763
rect 2875 7756 2975 7759
rect 3043 7756 3078 7793
rect 3140 7790 3499 7793
rect 3140 7785 3362 7790
rect 3140 7761 3153 7785
rect 3177 7766 3362 7785
rect 3386 7766 3499 7790
rect 3177 7761 3499 7766
rect 3140 7757 3499 7761
rect 3566 7785 3715 7793
rect 5319 7791 5851 7802
rect 3566 7765 3577 7785
rect 3597 7765 3715 7785
rect 5318 7775 5851 7791
rect 6488 7780 6519 7833
rect 6549 7862 6586 7941
rect 6757 7951 7150 7958
rect 6757 7934 6765 7951
rect 6797 7938 7150 7951
rect 7170 7938 7173 7958
rect 8252 7953 8293 7962
rect 6797 7934 7173 7938
rect 6757 7933 7173 7934
rect 7847 7951 8015 7952
rect 8252 7951 8261 7953
rect 6757 7932 7098 7933
rect 6701 7872 6732 7873
rect 6549 7842 6558 7862
rect 6578 7842 6586 7862
rect 6549 7832 6586 7842
rect 6645 7865 6732 7872
rect 6645 7862 6706 7865
rect 6645 7842 6654 7862
rect 6674 7845 6706 7862
rect 6727 7845 6732 7865
rect 6674 7842 6732 7845
rect 6645 7835 6732 7842
rect 6757 7862 6794 7932
rect 7060 7931 7097 7932
rect 7847 7931 8261 7951
rect 8287 7931 8293 7953
rect 8519 7960 8526 7980
rect 8545 7960 8561 7980
rect 8519 7952 8561 7960
rect 8589 7980 8630 7982
rect 8589 7960 8603 7980
rect 8622 7960 8630 7980
rect 8589 7952 8630 7960
rect 8885 7956 8922 7957
rect 9188 7956 9225 8026
rect 9250 8046 9337 8053
rect 9250 8043 9308 8046
rect 9250 8023 9255 8043
rect 9276 8026 9308 8043
rect 9328 8026 9337 8046
rect 9276 8023 9337 8026
rect 9250 8016 9337 8023
rect 9396 8046 9433 8056
rect 9396 8026 9404 8046
rect 9424 8026 9433 8046
rect 9250 8015 9281 8016
rect 8884 7955 9225 7956
rect 8519 7946 8630 7952
rect 8809 7950 9225 7955
rect 7847 7925 8293 7931
rect 7847 7923 8015 7925
rect 6909 7872 6945 7873
rect 6757 7842 6766 7862
rect 6786 7842 6794 7862
rect 6645 7833 6701 7835
rect 6645 7832 6682 7833
rect 6757 7832 6794 7842
rect 6853 7862 7001 7872
rect 7101 7869 7197 7871
rect 6853 7842 6862 7862
rect 6882 7857 6972 7862
rect 6882 7842 6917 7857
rect 6853 7833 6917 7842
rect 6853 7832 6890 7833
rect 6909 7816 6917 7833
rect 6938 7842 6972 7857
rect 6992 7842 7001 7862
rect 6938 7833 7001 7842
rect 7059 7862 7197 7869
rect 7059 7842 7068 7862
rect 7088 7842 7197 7862
rect 7059 7833 7197 7842
rect 6938 7816 6945 7833
rect 6964 7832 7001 7833
rect 7060 7832 7097 7833
rect 6909 7781 6945 7816
rect 6380 7779 6421 7780
rect 5318 7774 5832 7775
rect 3566 7758 3715 7765
rect 6272 7772 6421 7779
rect 4155 7762 4669 7763
rect 3566 7757 3607 7758
rect 2890 7704 2927 7705
rect 2986 7704 3023 7705
rect 3042 7704 3078 7756
rect 3097 7704 3134 7705
rect 2790 7695 2928 7704
rect 2790 7675 2899 7695
rect 2919 7675 2928 7695
rect 2790 7668 2928 7675
rect 2986 7695 3134 7704
rect 2986 7675 2995 7695
rect 3015 7675 3105 7695
rect 3125 7675 3134 7695
rect 2790 7666 2886 7668
rect 2986 7665 3134 7675
rect 3193 7695 3230 7705
rect 3305 7704 3342 7705
rect 3286 7702 3342 7704
rect 3193 7675 3201 7695
rect 3221 7675 3230 7695
rect 3042 7664 3078 7665
rect 1972 7612 2140 7614
rect 1694 7606 2140 7612
rect 762 7582 1178 7587
rect 1357 7585 1468 7591
rect 762 7581 1103 7582
rect 706 7521 737 7522
rect 554 7491 563 7511
rect 583 7491 591 7511
rect 554 7481 591 7491
rect 650 7514 737 7521
rect 650 7511 711 7514
rect 650 7491 659 7511
rect 679 7494 711 7511
rect 732 7494 737 7514
rect 679 7491 737 7494
rect 650 7484 737 7491
rect 762 7511 799 7581
rect 1065 7580 1102 7581
rect 1357 7577 1398 7585
rect 1357 7557 1365 7577
rect 1384 7557 1398 7577
rect 1357 7555 1398 7557
rect 1426 7577 1468 7585
rect 1426 7557 1442 7577
rect 1461 7557 1468 7577
rect 1694 7584 1700 7606
rect 1726 7586 2140 7606
rect 2890 7605 2927 7606
rect 3193 7605 3230 7675
rect 3255 7695 3342 7702
rect 3255 7692 3313 7695
rect 3255 7672 3260 7692
rect 3281 7675 3313 7692
rect 3333 7675 3342 7695
rect 3281 7672 3342 7675
rect 3255 7665 3342 7672
rect 3401 7695 3438 7705
rect 3401 7675 3409 7695
rect 3429 7675 3438 7695
rect 3255 7664 3286 7665
rect 2889 7604 3230 7605
rect 1726 7584 1735 7586
rect 1972 7585 2140 7586
rect 2814 7599 3230 7604
rect 1694 7575 1735 7584
rect 2814 7579 2817 7599
rect 2837 7579 3230 7599
rect 3401 7596 3438 7675
rect 3468 7704 3499 7757
rect 4136 7746 4669 7762
rect 6272 7752 6390 7772
rect 6410 7752 6421 7772
rect 4136 7735 4668 7746
rect 6272 7744 6421 7752
rect 6488 7776 6847 7780
rect 6488 7771 6810 7776
rect 6488 7747 6601 7771
rect 6625 7752 6810 7771
rect 6834 7752 6847 7776
rect 6625 7747 6847 7752
rect 6488 7744 6847 7747
rect 6909 7744 6944 7781
rect 7012 7778 7112 7781
rect 7012 7774 7079 7778
rect 7012 7748 7024 7774
rect 7050 7752 7079 7774
rect 7105 7752 7112 7778
rect 7050 7748 7112 7752
rect 7012 7744 7112 7748
rect 4787 7737 4824 7741
rect 3518 7704 3555 7705
rect 3468 7695 3555 7704
rect 3468 7675 3526 7695
rect 3546 7675 3555 7695
rect 3468 7665 3555 7675
rect 3614 7695 3651 7705
rect 3614 7675 3622 7695
rect 3642 7675 3651 7695
rect 3468 7664 3499 7665
rect 3463 7596 3573 7609
rect 3614 7596 3651 7675
rect 3401 7594 3651 7596
rect 3401 7591 3502 7594
rect 3401 7572 3466 7591
rect 1426 7555 1468 7557
rect 1357 7540 1468 7555
rect 3463 7564 3466 7572
rect 3495 7564 3502 7591
rect 3530 7567 3540 7594
rect 3569 7572 3651 7594
rect 3729 7666 3897 7667
rect 4136 7666 4174 7735
rect 3729 7646 4174 7666
rect 4401 7697 4512 7712
rect 4401 7695 4443 7697
rect 4401 7675 4408 7695
rect 4427 7675 4443 7695
rect 4401 7667 4443 7675
rect 4471 7695 4512 7697
rect 4471 7675 4485 7695
rect 4504 7675 4512 7695
rect 4471 7667 4512 7675
rect 4401 7661 4512 7667
rect 4634 7672 4668 7735
rect 4786 7731 4824 7737
rect 5166 7733 5203 7734
rect 4786 7713 4796 7731
rect 4814 7713 4824 7731
rect 4786 7704 4824 7713
rect 5164 7725 5204 7733
rect 5164 7707 5175 7725
rect 5193 7707 5204 7725
rect 6488 7723 6519 7744
rect 6909 7723 6945 7744
rect 6331 7722 6368 7723
rect 4786 7672 4820 7704
rect 3729 7640 4173 7646
rect 3729 7638 3897 7640
rect 3569 7567 3573 7572
rect 3530 7564 3573 7567
rect 3463 7550 3573 7564
rect 914 7521 950 7522
rect 762 7491 771 7511
rect 791 7491 799 7511
rect 650 7482 706 7484
rect 650 7481 687 7482
rect 762 7481 799 7491
rect 858 7511 1006 7521
rect 1106 7518 1202 7520
rect 858 7491 867 7511
rect 887 7491 977 7511
rect 997 7491 1006 7511
rect 858 7482 1006 7491
rect 1064 7511 1202 7518
rect 1064 7491 1073 7511
rect 1093 7491 1202 7511
rect 1064 7482 1202 7491
rect 858 7481 895 7482
rect 914 7430 950 7482
rect 969 7481 1006 7482
rect 1065 7481 1102 7482
rect 385 7428 426 7429
rect 277 7421 426 7428
rect 277 7401 395 7421
rect 415 7401 426 7421
rect 277 7393 426 7401
rect 493 7425 852 7429
rect 493 7420 815 7425
rect 493 7396 606 7420
rect 630 7401 815 7420
rect 839 7401 852 7425
rect 630 7396 852 7401
rect 493 7393 852 7396
rect 914 7393 949 7430
rect 1017 7427 1117 7430
rect 1017 7423 1084 7427
rect 1017 7397 1029 7423
rect 1055 7401 1084 7423
rect 1110 7401 1117 7427
rect 1055 7397 1117 7401
rect 1017 7393 1117 7397
rect 493 7372 524 7393
rect 914 7372 950 7393
rect 336 7371 373 7372
rect 335 7362 373 7371
rect 335 7342 344 7362
rect 364 7342 373 7362
rect 335 7334 373 7342
rect 439 7366 524 7372
rect 549 7371 586 7372
rect 439 7346 447 7366
rect 467 7346 524 7366
rect 439 7338 524 7346
rect 548 7362 586 7371
rect 548 7342 557 7362
rect 577 7342 586 7362
rect 439 7337 475 7338
rect 548 7334 586 7342
rect 652 7366 737 7372
rect 757 7371 794 7372
rect 652 7346 660 7366
rect 680 7365 737 7366
rect 680 7346 709 7365
rect 652 7345 709 7346
rect 730 7345 737 7365
rect 652 7338 737 7345
rect 756 7362 794 7371
rect 756 7342 765 7362
rect 785 7342 794 7362
rect 652 7337 688 7338
rect 756 7334 794 7342
rect 860 7366 1004 7372
rect 860 7346 868 7366
rect 888 7363 976 7366
rect 888 7346 919 7363
rect 860 7343 919 7346
rect 942 7346 976 7363
rect 996 7346 1004 7366
rect 942 7343 1004 7346
rect 860 7338 1004 7343
rect 860 7337 896 7338
rect 968 7337 1004 7338
rect 1070 7371 1107 7372
rect 1070 7370 1108 7371
rect 1070 7362 1134 7370
rect 1070 7342 1079 7362
rect 1099 7348 1134 7362
rect 1154 7348 1157 7368
rect 1099 7343 1157 7348
rect 1099 7342 1134 7343
rect 336 7305 373 7334
rect 337 7303 373 7305
rect 549 7303 586 7334
rect 337 7281 586 7303
rect 757 7302 794 7334
rect 1070 7330 1134 7342
rect 1174 7304 1201 7482
rect 3729 7460 3756 7638
rect 3796 7600 3860 7612
rect 4136 7608 4173 7640
rect 4344 7639 4593 7661
rect 4634 7640 4820 7672
rect 4648 7639 4820 7640
rect 4344 7608 4381 7639
rect 4557 7637 4593 7639
rect 4557 7608 4594 7637
rect 4786 7611 4820 7639
rect 5164 7659 5204 7707
rect 6330 7713 6368 7722
rect 6330 7693 6339 7713
rect 6359 7693 6368 7713
rect 6330 7685 6368 7693
rect 6434 7717 6519 7723
rect 6544 7722 6581 7723
rect 6434 7697 6442 7717
rect 6462 7697 6519 7717
rect 6434 7689 6519 7697
rect 6543 7713 6581 7722
rect 6543 7693 6552 7713
rect 6572 7693 6581 7713
rect 6434 7688 6470 7689
rect 6543 7685 6581 7693
rect 6647 7717 6732 7723
rect 6752 7722 6789 7723
rect 6647 7697 6655 7717
rect 6675 7716 6732 7717
rect 6675 7697 6704 7716
rect 6647 7696 6704 7697
rect 6725 7696 6732 7716
rect 6647 7689 6732 7696
rect 6751 7713 6789 7722
rect 6751 7693 6760 7713
rect 6780 7693 6789 7713
rect 6647 7688 6683 7689
rect 6751 7685 6789 7693
rect 6855 7717 6999 7723
rect 6855 7697 6863 7717
rect 6883 7697 6971 7717
rect 6991 7697 6999 7717
rect 6855 7689 6999 7697
rect 6855 7688 6891 7689
rect 6963 7688 6999 7689
rect 7065 7722 7102 7723
rect 7065 7721 7103 7722
rect 7065 7713 7129 7721
rect 7065 7693 7074 7713
rect 7094 7699 7129 7713
rect 7149 7699 7152 7719
rect 7094 7694 7152 7699
rect 7094 7693 7129 7694
rect 5475 7663 5585 7677
rect 5475 7660 5518 7663
rect 5164 7652 5289 7659
rect 5475 7655 5479 7660
rect 5164 7633 5256 7652
rect 5281 7633 5289 7652
rect 5164 7623 5289 7633
rect 5397 7633 5479 7655
rect 5508 7633 5518 7660
rect 5546 7636 5553 7663
rect 5582 7655 5585 7663
rect 6331 7656 6368 7685
rect 5582 7636 5647 7655
rect 6332 7654 6368 7656
rect 6544 7654 6581 7685
rect 6752 7658 6789 7685
rect 7065 7681 7129 7693
rect 5546 7633 5647 7636
rect 5397 7631 5647 7633
rect 3796 7599 3831 7600
rect 3773 7594 3831 7599
rect 3773 7574 3776 7594
rect 3796 7580 3831 7594
rect 3851 7580 3860 7600
rect 3796 7572 3860 7580
rect 3822 7571 3860 7572
rect 3823 7570 3860 7571
rect 3926 7604 3962 7605
rect 4034 7604 4070 7605
rect 3926 7597 4070 7604
rect 3926 7596 3986 7597
rect 3926 7576 3934 7596
rect 3954 7577 3986 7596
rect 4011 7596 4070 7597
rect 4011 7577 4042 7596
rect 3954 7576 4042 7577
rect 4062 7576 4070 7596
rect 3926 7570 4070 7576
rect 4136 7600 4174 7608
rect 4242 7604 4278 7605
rect 4136 7580 4145 7600
rect 4165 7580 4174 7600
rect 4136 7571 4174 7580
rect 4193 7597 4278 7604
rect 4193 7577 4200 7597
rect 4221 7596 4278 7597
rect 4221 7577 4250 7596
rect 4193 7576 4250 7577
rect 4270 7576 4278 7596
rect 4136 7570 4173 7571
rect 4193 7570 4278 7576
rect 4344 7600 4382 7608
rect 4455 7604 4491 7605
rect 4344 7580 4353 7600
rect 4373 7580 4382 7600
rect 4344 7571 4382 7580
rect 4406 7596 4491 7604
rect 4406 7576 4463 7596
rect 4483 7576 4491 7596
rect 4344 7570 4381 7571
rect 4406 7570 4491 7576
rect 4557 7600 4595 7608
rect 4557 7580 4566 7600
rect 4586 7580 4595 7600
rect 4557 7571 4595 7580
rect 4784 7601 4821 7611
rect 5164 7603 5204 7623
rect 4784 7583 4794 7601
rect 4812 7583 4821 7601
rect 4784 7574 4821 7583
rect 5163 7594 5204 7603
rect 5163 7576 5173 7594
rect 5191 7576 5204 7594
rect 4786 7573 4820 7574
rect 4557 7570 4594 7571
rect 3980 7549 4016 7570
rect 4406 7549 4437 7570
rect 5163 7567 5204 7576
rect 5163 7566 5200 7567
rect 5397 7552 5434 7631
rect 5475 7618 5585 7631
rect 5549 7562 5580 7563
rect 3813 7545 3913 7549
rect 3813 7541 3875 7545
rect 3813 7515 3820 7541
rect 3846 7519 3875 7541
rect 3901 7519 3913 7545
rect 3846 7515 3913 7519
rect 3813 7512 3913 7515
rect 3981 7512 4016 7549
rect 4078 7546 4437 7549
rect 4078 7541 4300 7546
rect 4078 7517 4091 7541
rect 4115 7522 4300 7541
rect 4324 7522 4437 7546
rect 4115 7517 4437 7522
rect 4078 7513 4437 7517
rect 4504 7541 4653 7549
rect 4504 7521 4515 7541
rect 4535 7521 4653 7541
rect 5397 7532 5406 7552
rect 5426 7532 5434 7552
rect 5397 7522 5434 7532
rect 5493 7552 5580 7562
rect 5493 7532 5502 7552
rect 5522 7532 5580 7552
rect 5493 7523 5580 7532
rect 5493 7522 5530 7523
rect 4504 7514 4653 7521
rect 4504 7513 4545 7514
rect 3828 7460 3865 7461
rect 3924 7460 3961 7461
rect 3980 7460 4016 7512
rect 4035 7460 4072 7461
rect 3728 7451 3866 7460
rect 3353 7417 3464 7432
rect 3728 7431 3837 7451
rect 3857 7431 3866 7451
rect 3728 7424 3866 7431
rect 3924 7451 4072 7460
rect 3924 7431 3933 7451
rect 3953 7431 4043 7451
rect 4063 7431 4072 7451
rect 3728 7422 3824 7424
rect 3924 7421 4072 7431
rect 4131 7451 4168 7461
rect 4243 7460 4280 7461
rect 4224 7458 4280 7460
rect 4131 7431 4139 7451
rect 4159 7431 4168 7451
rect 3980 7420 4016 7421
rect 3353 7415 3395 7417
rect 2690 7396 2760 7405
rect 2690 7387 2707 7396
rect 2681 7367 2707 7387
rect 2755 7387 2760 7396
rect 3353 7395 3360 7415
rect 3379 7395 3395 7415
rect 3353 7387 3395 7395
rect 3423 7415 3464 7417
rect 3423 7395 3437 7415
rect 3456 7395 3464 7415
rect 3423 7387 3464 7395
rect 2755 7386 2849 7387
rect 2755 7367 3125 7386
rect 3353 7381 3464 7387
rect 1468 7353 1578 7367
rect 1468 7350 1511 7353
rect 1468 7345 1472 7350
rect 1033 7302 1201 7304
rect 757 7299 1201 7302
rect 418 7275 529 7281
rect 418 7267 459 7275
rect 107 7212 146 7256
rect 418 7247 426 7267
rect 445 7247 459 7267
rect 418 7245 459 7247
rect 487 7267 529 7275
rect 487 7247 503 7267
rect 522 7247 529 7267
rect 487 7245 529 7247
rect 418 7231 529 7245
rect 755 7276 1201 7299
rect 107 7188 147 7212
rect 447 7188 494 7190
rect 755 7188 793 7276
rect 1033 7275 1201 7276
rect 1390 7323 1472 7345
rect 1501 7323 1511 7350
rect 1539 7326 1546 7353
rect 1575 7345 1578 7353
rect 2681 7360 3125 7367
rect 2681 7358 2849 7360
rect 2681 7350 2760 7358
rect 1575 7326 1640 7345
rect 1539 7323 1640 7326
rect 1390 7321 1640 7323
rect 1390 7242 1427 7321
rect 1468 7308 1578 7321
rect 1542 7252 1573 7253
rect 1390 7222 1399 7242
rect 1419 7222 1427 7242
rect 1390 7212 1427 7222
rect 1486 7242 1573 7252
rect 1486 7222 1495 7242
rect 1515 7222 1573 7242
rect 1486 7213 1573 7222
rect 1486 7212 1523 7213
rect 107 7155 793 7188
rect 1542 7160 1573 7213
rect 1603 7242 1640 7321
rect 1811 7318 2204 7338
rect 2224 7318 2227 7338
rect 1811 7313 2227 7318
rect 1811 7312 2152 7313
rect 1755 7252 1786 7253
rect 1603 7222 1612 7242
rect 1632 7222 1640 7242
rect 1603 7212 1640 7222
rect 1699 7245 1786 7252
rect 1699 7242 1760 7245
rect 1699 7222 1708 7242
rect 1728 7225 1760 7242
rect 1781 7225 1786 7245
rect 1728 7222 1786 7225
rect 1699 7215 1786 7222
rect 1811 7242 1848 7312
rect 2114 7311 2151 7312
rect 1963 7252 1999 7253
rect 1811 7222 1820 7242
rect 1840 7222 1848 7242
rect 1699 7213 1755 7215
rect 1699 7212 1736 7213
rect 1811 7212 1848 7222
rect 1907 7242 2055 7252
rect 2155 7249 2251 7251
rect 1907 7222 1916 7242
rect 1936 7222 2026 7242
rect 2046 7222 2055 7242
rect 1907 7213 2055 7222
rect 2113 7242 2251 7249
rect 2113 7222 2122 7242
rect 2142 7222 2251 7242
rect 2113 7213 2251 7222
rect 1907 7212 1944 7213
rect 1963 7161 1999 7213
rect 2018 7212 2055 7213
rect 2114 7212 2151 7213
rect 1434 7159 1475 7160
rect 106 7098 145 7155
rect 755 7153 793 7155
rect 1326 7152 1475 7159
rect 1326 7132 1444 7152
rect 1464 7132 1475 7152
rect 1326 7124 1475 7132
rect 1542 7156 1901 7160
rect 1542 7151 1864 7156
rect 1542 7127 1655 7151
rect 1679 7132 1864 7151
rect 1888 7132 1901 7156
rect 1679 7127 1901 7132
rect 1542 7124 1901 7127
rect 1963 7124 1998 7161
rect 2066 7158 2166 7161
rect 2066 7154 2133 7158
rect 2066 7128 2078 7154
rect 2104 7132 2133 7154
rect 2159 7132 2166 7158
rect 2104 7128 2166 7132
rect 2066 7124 2166 7128
rect 1542 7103 1573 7124
rect 1963 7103 1999 7124
rect 1385 7102 1422 7103
rect 106 7096 154 7098
rect 106 7078 117 7096
rect 135 7078 154 7096
rect 1384 7093 1422 7102
rect 106 7069 154 7078
rect 107 7068 154 7069
rect 420 7073 530 7087
rect 420 7070 463 7073
rect 420 7065 424 7070
rect 342 7043 424 7065
rect 453 7043 463 7070
rect 491 7046 498 7073
rect 527 7065 530 7073
rect 1384 7073 1393 7093
rect 1413 7073 1422 7093
rect 1384 7065 1422 7073
rect 1488 7097 1573 7103
rect 1598 7102 1635 7103
rect 1488 7077 1496 7097
rect 1516 7077 1573 7097
rect 1488 7069 1573 7077
rect 1597 7093 1635 7102
rect 1597 7073 1606 7093
rect 1626 7073 1635 7093
rect 1488 7068 1524 7069
rect 1597 7065 1635 7073
rect 1701 7097 1786 7103
rect 1806 7102 1843 7103
rect 1701 7077 1709 7097
rect 1729 7096 1786 7097
rect 1729 7077 1758 7096
rect 1701 7076 1758 7077
rect 1779 7076 1786 7096
rect 1701 7069 1786 7076
rect 1805 7093 1843 7102
rect 1805 7073 1814 7093
rect 1834 7073 1843 7093
rect 1701 7068 1737 7069
rect 1805 7065 1843 7073
rect 1909 7097 2053 7103
rect 1909 7077 1917 7097
rect 1937 7095 2025 7097
rect 1937 7077 1966 7095
rect 1909 7076 1966 7077
rect 1995 7077 2025 7095
rect 2045 7077 2053 7097
rect 1995 7076 2053 7077
rect 1909 7069 2053 7076
rect 1909 7068 1945 7069
rect 2017 7068 2053 7069
rect 2119 7102 2156 7103
rect 2119 7101 2157 7102
rect 2119 7093 2183 7101
rect 2119 7073 2128 7093
rect 2148 7079 2183 7093
rect 2203 7079 2206 7099
rect 2148 7074 2206 7079
rect 2148 7073 2183 7074
rect 527 7046 592 7065
rect 491 7043 592 7046
rect 342 7041 592 7043
rect 110 7005 147 7006
rect 106 7002 147 7005
rect 106 6997 148 7002
rect 106 6979 119 6997
rect 137 6979 148 6997
rect 106 6965 148 6979
rect 186 6965 233 6969
rect 106 6959 233 6965
rect 106 6930 194 6959
rect 223 6930 233 6959
rect 342 6962 379 7041
rect 420 7028 530 7041
rect 494 6972 525 6973
rect 342 6942 351 6962
rect 371 6942 379 6962
rect 342 6932 379 6942
rect 438 6962 525 6972
rect 438 6942 447 6962
rect 467 6942 525 6962
rect 438 6933 525 6942
rect 438 6932 475 6933
rect 106 6926 233 6930
rect 106 6909 145 6926
rect 186 6925 233 6926
rect 106 6891 117 6909
rect 135 6891 145 6909
rect 106 6882 145 6891
rect 107 6881 144 6882
rect 494 6880 525 6933
rect 555 6962 592 7041
rect 763 7038 1156 7058
rect 1176 7038 1179 7058
rect 763 7033 1179 7038
rect 1385 7036 1422 7065
rect 1386 7034 1422 7036
rect 1598 7034 1635 7065
rect 763 7032 1104 7033
rect 707 6972 738 6973
rect 555 6942 564 6962
rect 584 6942 592 6962
rect 555 6932 592 6942
rect 651 6965 738 6972
rect 651 6962 712 6965
rect 651 6942 660 6962
rect 680 6945 712 6962
rect 733 6945 738 6965
rect 680 6942 738 6945
rect 651 6935 738 6942
rect 763 6962 800 7032
rect 1066 7031 1103 7032
rect 1386 7012 1635 7034
rect 1806 7033 1843 7065
rect 2119 7061 2183 7073
rect 2223 7037 2250 7213
rect 2681 7180 2708 7350
rect 2748 7320 2812 7332
rect 3088 7328 3125 7360
rect 3296 7359 3545 7381
rect 3828 7361 3865 7362
rect 4131 7361 4168 7431
rect 4193 7451 4280 7458
rect 4193 7448 4251 7451
rect 4193 7428 4198 7448
rect 4219 7431 4251 7448
rect 4271 7431 4280 7451
rect 4219 7428 4280 7431
rect 4193 7421 4280 7428
rect 4339 7451 4376 7461
rect 4339 7431 4347 7451
rect 4367 7431 4376 7451
rect 4193 7420 4224 7421
rect 3827 7360 4168 7361
rect 3296 7328 3333 7359
rect 3509 7357 3545 7359
rect 3509 7328 3546 7357
rect 3752 7355 4168 7360
rect 3752 7335 3755 7355
rect 3775 7335 4168 7355
rect 4339 7352 4376 7431
rect 4406 7460 4437 7513
rect 4787 7511 4824 7512
rect 4786 7502 4825 7511
rect 4786 7484 4796 7502
rect 4814 7484 4825 7502
rect 5166 7500 5203 7504
rect 4698 7467 4745 7468
rect 4786 7467 4825 7484
rect 4698 7463 4825 7467
rect 4456 7460 4493 7461
rect 4406 7451 4493 7460
rect 4406 7431 4464 7451
rect 4484 7431 4493 7451
rect 4406 7421 4493 7431
rect 4552 7451 4589 7461
rect 4552 7431 4560 7451
rect 4580 7431 4589 7451
rect 4406 7420 4437 7421
rect 4401 7352 4511 7365
rect 4552 7352 4589 7431
rect 4698 7434 4708 7463
rect 4737 7434 4825 7463
rect 4698 7428 4825 7434
rect 4698 7424 4745 7428
rect 4783 7414 4825 7428
rect 4783 7396 4794 7414
rect 4812 7396 4825 7414
rect 4783 7391 4825 7396
rect 4784 7388 4825 7391
rect 5163 7495 5203 7500
rect 5163 7477 5175 7495
rect 5193 7477 5203 7495
rect 4784 7387 4821 7388
rect 4339 7350 4589 7352
rect 4339 7347 4440 7350
rect 4339 7328 4404 7347
rect 2748 7319 2783 7320
rect 2725 7314 2783 7319
rect 2725 7294 2728 7314
rect 2748 7300 2783 7314
rect 2803 7300 2812 7320
rect 2748 7292 2812 7300
rect 2774 7291 2812 7292
rect 2775 7290 2812 7291
rect 2878 7324 2914 7325
rect 2986 7324 3022 7325
rect 2878 7316 3022 7324
rect 2878 7296 2886 7316
rect 2906 7296 2994 7316
rect 3014 7296 3022 7316
rect 2878 7290 3022 7296
rect 3088 7320 3126 7328
rect 3194 7324 3230 7325
rect 3088 7300 3097 7320
rect 3117 7300 3126 7320
rect 3088 7291 3126 7300
rect 3145 7317 3230 7324
rect 3145 7297 3152 7317
rect 3173 7316 3230 7317
rect 3173 7297 3202 7316
rect 3145 7296 3202 7297
rect 3222 7296 3230 7316
rect 3088 7290 3125 7291
rect 3145 7290 3230 7296
rect 3296 7320 3334 7328
rect 3407 7324 3443 7325
rect 3296 7300 3305 7320
rect 3325 7300 3334 7320
rect 3296 7291 3334 7300
rect 3358 7316 3443 7324
rect 3358 7296 3415 7316
rect 3435 7296 3443 7316
rect 3296 7290 3333 7291
rect 3358 7290 3443 7296
rect 3509 7320 3547 7328
rect 3509 7300 3518 7320
rect 3538 7300 3547 7320
rect 4401 7320 4404 7328
rect 4433 7320 4440 7347
rect 4468 7323 4478 7350
rect 4507 7328 4589 7350
rect 4507 7323 4511 7328
rect 4468 7320 4511 7323
rect 4401 7306 4511 7320
rect 4777 7324 4824 7325
rect 4777 7315 4825 7324
rect 3509 7291 3547 7300
rect 4777 7297 4796 7315
rect 4814 7297 4825 7315
rect 4777 7295 4825 7297
rect 3509 7290 3546 7291
rect 2932 7269 2968 7290
rect 3358 7269 3389 7290
rect 2765 7265 2865 7269
rect 2765 7261 2827 7265
rect 2765 7235 2772 7261
rect 2798 7239 2827 7261
rect 2853 7239 2865 7265
rect 2798 7235 2865 7239
rect 2765 7232 2865 7235
rect 2933 7232 2968 7269
rect 3030 7266 3389 7269
rect 3030 7261 3252 7266
rect 3030 7237 3043 7261
rect 3067 7242 3252 7261
rect 3276 7242 3389 7266
rect 3067 7237 3389 7242
rect 3030 7233 3389 7237
rect 3456 7261 3605 7269
rect 3456 7241 3467 7261
rect 3487 7241 3605 7261
rect 3456 7234 3605 7241
rect 4138 7238 4176 7240
rect 4786 7238 4825 7295
rect 5163 7297 5203 7477
rect 5549 7470 5580 7523
rect 5610 7552 5647 7631
rect 5818 7628 6211 7648
rect 6231 7628 6234 7648
rect 6332 7632 6581 7654
rect 6750 7653 6791 7658
rect 7169 7655 7196 7833
rect 7847 7745 7874 7923
rect 8252 7920 8293 7925
rect 8462 7924 8711 7946
rect 8809 7930 8812 7950
rect 8832 7930 9225 7950
rect 9396 7947 9433 8026
rect 9463 8055 9494 8108
rect 9840 8101 9880 8281
rect 10137 8364 10177 8544
rect 10523 8537 10554 8590
rect 10584 8619 10621 8698
rect 10792 8695 11185 8715
rect 11205 8695 11208 8715
rect 11306 8699 11555 8721
rect 11724 8720 11765 8725
rect 12143 8722 12170 8900
rect 12821 8812 12848 8990
rect 13226 8987 13267 8992
rect 13436 8991 13685 9013
rect 13783 8997 13786 9017
rect 13806 8997 14199 9017
rect 14370 9014 14407 9093
rect 14437 9122 14468 9175
rect 14814 9168 14854 9348
rect 15192 9348 15246 9353
rect 15192 9330 15203 9348
rect 15221 9330 15246 9348
rect 18816 9369 18984 9370
rect 19224 9369 19262 9457
rect 19523 9439 19570 9457
rect 19487 9400 19599 9439
rect 19870 9433 19910 9457
rect 19487 9399 19530 9400
rect 18816 9346 19262 9369
rect 19488 9398 19530 9399
rect 19488 9378 19495 9398
rect 19514 9378 19530 9398
rect 19488 9370 19530 9378
rect 19558 9398 19599 9400
rect 19558 9378 19572 9398
rect 19591 9378 19599 9398
rect 19871 9389 19910 9433
rect 19558 9370 19599 9378
rect 19488 9364 19599 9370
rect 18816 9343 19260 9346
rect 18816 9341 18984 9343
rect 15192 9321 15246 9330
rect 15193 9320 15246 9321
rect 15506 9325 15616 9339
rect 15506 9322 15549 9325
rect 15506 9317 15510 9322
rect 15428 9295 15510 9317
rect 15539 9295 15549 9322
rect 15577 9298 15584 9325
rect 15613 9317 15616 9325
rect 15613 9298 15678 9317
rect 15577 9295 15678 9298
rect 15428 9293 15678 9295
rect 15196 9257 15233 9258
rect 14814 9150 14824 9168
rect 14842 9150 14854 9168
rect 14814 9145 14854 9150
rect 15192 9254 15233 9257
rect 15192 9249 15234 9254
rect 15192 9231 15205 9249
rect 15223 9231 15234 9249
rect 15192 9217 15234 9231
rect 15272 9217 15319 9221
rect 15192 9211 15319 9217
rect 15192 9182 15280 9211
rect 15309 9182 15319 9211
rect 15428 9214 15465 9293
rect 15506 9280 15616 9293
rect 15580 9224 15611 9225
rect 15428 9194 15437 9214
rect 15457 9194 15465 9214
rect 15428 9184 15465 9194
rect 15524 9214 15611 9224
rect 15524 9194 15533 9214
rect 15553 9194 15611 9214
rect 15524 9185 15611 9194
rect 15524 9184 15561 9185
rect 15192 9178 15319 9182
rect 15192 9161 15231 9178
rect 15272 9177 15319 9178
rect 14814 9141 14851 9145
rect 15192 9143 15203 9161
rect 15221 9143 15231 9161
rect 15192 9134 15231 9143
rect 15193 9133 15230 9134
rect 15580 9132 15611 9185
rect 15641 9214 15678 9293
rect 15849 9290 16242 9310
rect 16262 9290 16265 9310
rect 15849 9285 16265 9290
rect 15849 9284 16190 9285
rect 15793 9224 15824 9225
rect 15641 9194 15650 9214
rect 15670 9194 15678 9214
rect 15641 9184 15678 9194
rect 15737 9217 15824 9224
rect 15737 9214 15798 9217
rect 15737 9194 15746 9214
rect 15766 9197 15798 9214
rect 15819 9197 15824 9217
rect 15766 9194 15824 9197
rect 15737 9187 15824 9194
rect 15849 9214 15886 9284
rect 16152 9283 16189 9284
rect 16001 9224 16037 9225
rect 15849 9194 15858 9214
rect 15878 9194 15886 9214
rect 15737 9185 15793 9187
rect 15737 9184 15774 9185
rect 15849 9184 15886 9194
rect 15945 9214 16093 9224
rect 16193 9221 16289 9223
rect 15945 9194 15954 9214
rect 15974 9194 16064 9214
rect 16084 9194 16093 9214
rect 15945 9185 16093 9194
rect 16151 9214 16289 9221
rect 16151 9194 16160 9214
rect 16180 9194 16289 9214
rect 16151 9185 16289 9194
rect 15945 9184 15982 9185
rect 16001 9133 16037 9185
rect 16056 9184 16093 9185
rect 16152 9184 16189 9185
rect 15472 9131 15513 9132
rect 15364 9124 15513 9131
rect 14487 9122 14524 9123
rect 14437 9113 14524 9122
rect 14437 9093 14495 9113
rect 14515 9093 14524 9113
rect 14437 9083 14524 9093
rect 14583 9113 14620 9123
rect 14583 9093 14591 9113
rect 14611 9093 14620 9113
rect 15364 9104 15482 9124
rect 15502 9104 15513 9124
rect 15364 9096 15513 9104
rect 15580 9128 15939 9132
rect 15580 9123 15902 9128
rect 15580 9099 15693 9123
rect 15717 9104 15902 9123
rect 15926 9104 15939 9128
rect 15717 9099 15939 9104
rect 15580 9096 15939 9099
rect 16001 9096 16036 9133
rect 16104 9130 16204 9133
rect 16104 9126 16171 9130
rect 16104 9100 16116 9126
rect 16142 9104 16171 9126
rect 16197 9104 16204 9130
rect 16142 9100 16204 9104
rect 16104 9096 16204 9100
rect 14437 9082 14468 9083
rect 14432 9014 14542 9027
rect 14583 9014 14620 9093
rect 14817 9078 14854 9079
rect 14813 9069 14854 9078
rect 15580 9075 15611 9096
rect 16001 9075 16037 9096
rect 15423 9074 15460 9075
rect 15197 9071 15231 9072
rect 14813 9051 14826 9069
rect 14844 9051 14854 9069
rect 14813 9042 14854 9051
rect 15196 9062 15233 9071
rect 15196 9044 15205 9062
rect 15223 9044 15233 9062
rect 14813 9022 14853 9042
rect 15196 9034 15233 9044
rect 15422 9065 15460 9074
rect 15422 9045 15431 9065
rect 15451 9045 15460 9065
rect 15422 9037 15460 9045
rect 15526 9069 15611 9075
rect 15636 9074 15673 9075
rect 15526 9049 15534 9069
rect 15554 9049 15611 9069
rect 15526 9041 15611 9049
rect 15635 9065 15673 9074
rect 15635 9045 15644 9065
rect 15664 9045 15673 9065
rect 15526 9040 15562 9041
rect 15635 9037 15673 9045
rect 15739 9069 15824 9075
rect 15844 9074 15881 9075
rect 15739 9049 15747 9069
rect 15767 9068 15824 9069
rect 15767 9049 15796 9068
rect 15739 9048 15796 9049
rect 15817 9048 15824 9068
rect 15739 9041 15824 9048
rect 15843 9065 15881 9074
rect 15843 9045 15852 9065
rect 15872 9045 15881 9065
rect 15739 9040 15775 9041
rect 15843 9037 15881 9045
rect 15947 9069 16091 9075
rect 15947 9049 15955 9069
rect 15975 9068 16063 9069
rect 15975 9049 16006 9068
rect 15947 9048 16006 9049
rect 16031 9049 16063 9068
rect 16083 9049 16091 9069
rect 16031 9048 16091 9049
rect 15947 9041 16091 9048
rect 15947 9040 15983 9041
rect 16055 9040 16091 9041
rect 16157 9074 16194 9075
rect 16157 9073 16195 9074
rect 16157 9065 16221 9073
rect 16157 9045 16166 9065
rect 16186 9051 16221 9065
rect 16241 9051 16244 9071
rect 16186 9046 16244 9051
rect 16186 9045 16221 9046
rect 14370 9012 14620 9014
rect 14370 9009 14471 9012
rect 12888 8952 12952 8964
rect 13228 8960 13265 8987
rect 13436 8960 13473 8991
rect 13649 8989 13685 8991
rect 14370 8990 14435 9009
rect 13649 8960 13686 8989
rect 14432 8982 14435 8990
rect 14464 8982 14471 9009
rect 14499 8985 14509 9012
rect 14538 8990 14620 9012
rect 14728 9012 14853 9022
rect 14728 8993 14736 9012
rect 14761 8993 14853 9012
rect 14538 8985 14542 8990
rect 14728 8986 14853 8993
rect 14499 8982 14542 8985
rect 14432 8968 14542 8982
rect 12888 8951 12923 8952
rect 12865 8946 12923 8951
rect 12865 8926 12868 8946
rect 12888 8932 12923 8946
rect 12943 8932 12952 8952
rect 12888 8924 12952 8932
rect 12914 8923 12952 8924
rect 12915 8922 12952 8923
rect 13018 8956 13054 8957
rect 13126 8956 13162 8957
rect 13018 8948 13162 8956
rect 13018 8928 13026 8948
rect 13046 8928 13134 8948
rect 13154 8928 13162 8948
rect 13018 8922 13162 8928
rect 13228 8952 13266 8960
rect 13334 8956 13370 8957
rect 13228 8932 13237 8952
rect 13257 8932 13266 8952
rect 13228 8923 13266 8932
rect 13285 8949 13370 8956
rect 13285 8929 13292 8949
rect 13313 8948 13370 8949
rect 13313 8929 13342 8948
rect 13285 8928 13342 8929
rect 13362 8928 13370 8948
rect 13228 8922 13265 8923
rect 13285 8922 13370 8928
rect 13436 8952 13474 8960
rect 13547 8956 13583 8957
rect 13436 8932 13445 8952
rect 13465 8932 13474 8952
rect 13436 8923 13474 8932
rect 13498 8948 13583 8956
rect 13498 8928 13555 8948
rect 13575 8928 13583 8948
rect 13436 8922 13473 8923
rect 13498 8922 13583 8928
rect 13649 8952 13687 8960
rect 13649 8932 13658 8952
rect 13678 8932 13687 8952
rect 13649 8923 13687 8932
rect 14813 8938 14853 8986
rect 15197 9006 15231 9034
rect 15423 9008 15460 9037
rect 15424 9006 15460 9008
rect 15636 9006 15673 9037
rect 15197 9005 15369 9006
rect 15197 8973 15383 9005
rect 15424 8984 15673 9006
rect 15844 9005 15881 9037
rect 16157 9033 16221 9045
rect 16261 9007 16288 9185
rect 18816 9163 18843 9341
rect 18883 9303 18947 9315
rect 19223 9311 19260 9343
rect 19431 9342 19680 9364
rect 19431 9311 19468 9342
rect 19644 9340 19680 9342
rect 19644 9311 19681 9340
rect 18883 9302 18918 9303
rect 18860 9297 18918 9302
rect 18860 9277 18863 9297
rect 18883 9283 18918 9297
rect 18938 9283 18947 9303
rect 18883 9275 18947 9283
rect 18909 9274 18947 9275
rect 18910 9273 18947 9274
rect 19013 9307 19049 9308
rect 19121 9307 19157 9308
rect 19013 9302 19157 9307
rect 19013 9299 19075 9302
rect 19013 9279 19021 9299
rect 19041 9282 19075 9299
rect 19098 9299 19157 9302
rect 19098 9282 19129 9299
rect 19041 9279 19129 9282
rect 19149 9279 19157 9299
rect 19013 9273 19157 9279
rect 19223 9303 19261 9311
rect 19329 9307 19365 9308
rect 19223 9283 19232 9303
rect 19252 9283 19261 9303
rect 19223 9274 19261 9283
rect 19280 9300 19365 9307
rect 19280 9280 19287 9300
rect 19308 9299 19365 9300
rect 19308 9280 19337 9299
rect 19280 9279 19337 9280
rect 19357 9279 19365 9299
rect 19223 9273 19260 9274
rect 19280 9273 19365 9279
rect 19431 9303 19469 9311
rect 19542 9307 19578 9308
rect 19431 9283 19440 9303
rect 19460 9283 19469 9303
rect 19431 9274 19469 9283
rect 19493 9299 19578 9307
rect 19493 9279 19550 9299
rect 19570 9279 19578 9299
rect 19431 9273 19468 9274
rect 19493 9273 19578 9279
rect 19644 9303 19682 9311
rect 19644 9283 19653 9303
rect 19673 9283 19682 9303
rect 19644 9274 19682 9283
rect 19644 9273 19681 9274
rect 19067 9252 19103 9273
rect 19493 9252 19524 9273
rect 18900 9248 19000 9252
rect 18900 9244 18962 9248
rect 18900 9218 18907 9244
rect 18933 9222 18962 9244
rect 18988 9222 19000 9248
rect 18933 9218 19000 9222
rect 18900 9215 19000 9218
rect 19068 9215 19103 9252
rect 19165 9249 19524 9252
rect 19165 9244 19387 9249
rect 19165 9220 19178 9244
rect 19202 9225 19387 9244
rect 19411 9225 19524 9249
rect 19202 9220 19524 9225
rect 19165 9216 19524 9220
rect 19591 9244 19740 9252
rect 19591 9224 19602 9244
rect 19622 9224 19740 9244
rect 19591 9217 19740 9224
rect 19591 9216 19632 9217
rect 18915 9163 18952 9164
rect 19011 9163 19048 9164
rect 19067 9163 19103 9215
rect 19122 9163 19159 9164
rect 18815 9154 18953 9163
rect 18815 9134 18924 9154
rect 18944 9134 18953 9154
rect 18815 9127 18953 9134
rect 19011 9154 19159 9163
rect 19011 9134 19020 9154
rect 19040 9134 19130 9154
rect 19150 9134 19159 9154
rect 18815 9125 18911 9127
rect 19011 9124 19159 9134
rect 19218 9154 19255 9164
rect 19330 9163 19367 9164
rect 19311 9161 19367 9163
rect 19218 9134 19226 9154
rect 19246 9134 19255 9154
rect 19067 9123 19103 9124
rect 16444 9081 16554 9095
rect 16444 9078 16487 9081
rect 16444 9073 16448 9078
rect 16120 9005 16288 9007
rect 15844 8999 16288 9005
rect 15197 8941 15231 8973
rect 13649 8922 13686 8923
rect 13072 8901 13108 8922
rect 13498 8901 13529 8922
rect 14813 8920 14824 8938
rect 14842 8920 14853 8938
rect 14813 8912 14853 8920
rect 15193 8932 15231 8941
rect 15193 8914 15203 8932
rect 15221 8914 15231 8932
rect 14814 8911 14851 8912
rect 15193 8908 15231 8914
rect 15349 8910 15383 8973
rect 15505 8978 15616 8984
rect 15505 8970 15546 8978
rect 15505 8950 15513 8970
rect 15532 8950 15546 8970
rect 15505 8948 15546 8950
rect 15574 8970 15616 8978
rect 15574 8950 15590 8970
rect 15609 8950 15616 8970
rect 15574 8948 15616 8950
rect 15505 8933 15616 8948
rect 15843 8979 16288 8999
rect 15843 8910 15881 8979
rect 16120 8978 16288 8979
rect 16366 9051 16448 9073
rect 16477 9051 16487 9078
rect 16515 9054 16522 9081
rect 16551 9073 16554 9081
rect 18549 9090 18660 9105
rect 18549 9088 18591 9090
rect 16551 9054 16616 9073
rect 16515 9051 16616 9054
rect 16366 9049 16616 9051
rect 16366 8970 16403 9049
rect 16444 9036 16554 9049
rect 16518 8980 16549 8981
rect 16366 8950 16375 8970
rect 16395 8950 16403 8970
rect 16366 8940 16403 8950
rect 16462 8970 16549 8980
rect 16462 8950 16471 8970
rect 16491 8950 16549 8970
rect 16462 8941 16549 8950
rect 16462 8940 16499 8941
rect 15193 8904 15230 8908
rect 12905 8897 13005 8901
rect 12905 8893 12967 8897
rect 12905 8867 12912 8893
rect 12938 8871 12967 8893
rect 12993 8871 13005 8897
rect 12938 8867 13005 8871
rect 12905 8864 13005 8867
rect 13073 8864 13108 8901
rect 13170 8898 13529 8901
rect 13170 8893 13392 8898
rect 13170 8869 13183 8893
rect 13207 8874 13392 8893
rect 13416 8874 13529 8898
rect 13207 8869 13529 8874
rect 13170 8865 13529 8869
rect 13596 8893 13745 8901
rect 15349 8899 15881 8910
rect 13596 8873 13607 8893
rect 13627 8873 13745 8893
rect 15348 8883 15881 8899
rect 16518 8888 16549 8941
rect 16579 8970 16616 9049
rect 16787 9046 17180 9066
rect 17200 9046 17203 9066
rect 18282 9061 18323 9070
rect 16787 9041 17203 9046
rect 17877 9059 18045 9060
rect 18282 9059 18291 9061
rect 16787 9040 17128 9041
rect 16731 8980 16762 8981
rect 16579 8950 16588 8970
rect 16608 8950 16616 8970
rect 16579 8940 16616 8950
rect 16675 8973 16762 8980
rect 16675 8970 16736 8973
rect 16675 8950 16684 8970
rect 16704 8953 16736 8970
rect 16757 8953 16762 8973
rect 16704 8950 16762 8953
rect 16675 8943 16762 8950
rect 16787 8970 16824 9040
rect 17090 9039 17127 9040
rect 17877 9039 18291 9059
rect 18317 9039 18323 9061
rect 18549 9068 18556 9088
rect 18575 9068 18591 9088
rect 18549 9060 18591 9068
rect 18619 9088 18660 9090
rect 18619 9068 18633 9088
rect 18652 9068 18660 9088
rect 18619 9060 18660 9068
rect 18915 9064 18952 9065
rect 19218 9064 19255 9134
rect 19280 9154 19367 9161
rect 19280 9151 19338 9154
rect 19280 9131 19285 9151
rect 19306 9134 19338 9151
rect 19358 9134 19367 9154
rect 19306 9131 19367 9134
rect 19280 9124 19367 9131
rect 19426 9154 19463 9164
rect 19426 9134 19434 9154
rect 19454 9134 19463 9154
rect 19280 9123 19311 9124
rect 18914 9063 19255 9064
rect 18549 9054 18660 9060
rect 18839 9058 19255 9063
rect 17877 9033 18323 9039
rect 17877 9031 18045 9033
rect 16939 8980 16975 8981
rect 16787 8950 16796 8970
rect 16816 8950 16824 8970
rect 16675 8941 16731 8943
rect 16675 8940 16712 8941
rect 16787 8940 16824 8950
rect 16883 8970 17031 8980
rect 17131 8977 17227 8979
rect 16883 8950 16892 8970
rect 16912 8950 17002 8970
rect 17022 8950 17031 8970
rect 16883 8941 17031 8950
rect 17089 8970 17227 8977
rect 17089 8950 17098 8970
rect 17118 8950 17227 8970
rect 17089 8941 17227 8950
rect 16883 8940 16920 8941
rect 16939 8889 16975 8941
rect 16994 8940 17031 8941
rect 17090 8940 17127 8941
rect 16410 8887 16451 8888
rect 15348 8882 15862 8883
rect 13596 8866 13745 8873
rect 16302 8880 16451 8887
rect 14185 8870 14699 8871
rect 13596 8865 13637 8866
rect 13072 8829 13108 8864
rect 12920 8812 12957 8813
rect 13016 8812 13053 8813
rect 13072 8812 13079 8829
rect 12820 8803 12958 8812
rect 12820 8783 12929 8803
rect 12949 8783 12958 8803
rect 12820 8776 12958 8783
rect 13016 8803 13079 8812
rect 13016 8783 13025 8803
rect 13045 8788 13079 8803
rect 13100 8812 13108 8829
rect 13127 8812 13164 8813
rect 13100 8803 13164 8812
rect 13100 8788 13135 8803
rect 13045 8783 13135 8788
rect 13155 8783 13164 8803
rect 12820 8774 12916 8776
rect 13016 8773 13164 8783
rect 13223 8803 13260 8813
rect 13335 8812 13372 8813
rect 13316 8810 13372 8812
rect 13223 8783 13231 8803
rect 13251 8783 13260 8803
rect 13072 8772 13108 8773
rect 12002 8720 12170 8722
rect 11724 8714 12170 8720
rect 10792 8690 11208 8695
rect 11387 8693 11498 8699
rect 10792 8689 11133 8690
rect 10736 8629 10767 8630
rect 10584 8599 10593 8619
rect 10613 8599 10621 8619
rect 10584 8589 10621 8599
rect 10680 8622 10767 8629
rect 10680 8619 10741 8622
rect 10680 8599 10689 8619
rect 10709 8602 10741 8619
rect 10762 8602 10767 8622
rect 10709 8599 10767 8602
rect 10680 8592 10767 8599
rect 10792 8619 10829 8689
rect 11095 8688 11132 8689
rect 11387 8685 11428 8693
rect 11387 8665 11395 8685
rect 11414 8665 11428 8685
rect 11387 8663 11428 8665
rect 11456 8685 11498 8693
rect 11456 8665 11472 8685
rect 11491 8665 11498 8685
rect 11724 8692 11730 8714
rect 11756 8694 12170 8714
rect 12920 8713 12957 8714
rect 13223 8713 13260 8783
rect 13285 8803 13372 8810
rect 13285 8800 13343 8803
rect 13285 8780 13290 8800
rect 13311 8783 13343 8800
rect 13363 8783 13372 8803
rect 13311 8780 13372 8783
rect 13285 8773 13372 8780
rect 13431 8803 13468 8813
rect 13431 8783 13439 8803
rect 13459 8783 13468 8803
rect 13285 8772 13316 8773
rect 12919 8712 13260 8713
rect 11756 8692 11765 8694
rect 12002 8693 12170 8694
rect 12844 8711 13260 8712
rect 12844 8707 13220 8711
rect 11724 8683 11765 8692
rect 12844 8687 12847 8707
rect 12867 8694 13220 8707
rect 13252 8694 13260 8711
rect 12867 8687 13260 8694
rect 13431 8704 13468 8783
rect 13498 8812 13529 8865
rect 14166 8854 14699 8870
rect 16302 8860 16420 8880
rect 16440 8860 16451 8880
rect 14166 8843 14698 8854
rect 16302 8852 16451 8860
rect 16518 8884 16877 8888
rect 16518 8879 16840 8884
rect 16518 8855 16631 8879
rect 16655 8860 16840 8879
rect 16864 8860 16877 8884
rect 16655 8855 16877 8860
rect 16518 8852 16877 8855
rect 16939 8852 16974 8889
rect 17042 8886 17142 8889
rect 17042 8882 17109 8886
rect 17042 8856 17054 8882
rect 17080 8860 17109 8882
rect 17135 8860 17142 8886
rect 17080 8856 17142 8860
rect 17042 8852 17142 8856
rect 14817 8845 14854 8849
rect 13548 8812 13585 8813
rect 13498 8803 13585 8812
rect 13498 8783 13556 8803
rect 13576 8783 13585 8803
rect 13498 8773 13585 8783
rect 13644 8803 13681 8813
rect 13644 8783 13652 8803
rect 13672 8783 13681 8803
rect 13498 8772 13529 8773
rect 13493 8704 13603 8717
rect 13644 8704 13681 8783
rect 13431 8702 13681 8704
rect 13431 8699 13532 8702
rect 13431 8680 13496 8699
rect 11456 8663 11498 8665
rect 11387 8648 11498 8663
rect 13493 8672 13496 8680
rect 13525 8672 13532 8699
rect 13560 8675 13570 8702
rect 13599 8680 13681 8702
rect 13759 8774 13927 8775
rect 14166 8774 14204 8843
rect 13759 8754 14204 8774
rect 14431 8805 14542 8820
rect 14431 8803 14473 8805
rect 14431 8783 14438 8803
rect 14457 8783 14473 8803
rect 14431 8775 14473 8783
rect 14501 8803 14542 8805
rect 14501 8783 14515 8803
rect 14534 8783 14542 8803
rect 14501 8775 14542 8783
rect 14431 8769 14542 8775
rect 14664 8780 14698 8843
rect 14816 8839 14854 8845
rect 15196 8841 15233 8842
rect 14816 8821 14826 8839
rect 14844 8821 14854 8839
rect 14816 8812 14854 8821
rect 15194 8833 15234 8841
rect 15194 8815 15205 8833
rect 15223 8815 15234 8833
rect 16518 8831 16549 8852
rect 16939 8831 16975 8852
rect 16361 8830 16398 8831
rect 14816 8780 14850 8812
rect 13759 8748 14203 8754
rect 13759 8746 13927 8748
rect 13599 8675 13603 8680
rect 13560 8672 13603 8675
rect 13493 8658 13603 8672
rect 10944 8629 10980 8630
rect 10792 8599 10801 8619
rect 10821 8599 10829 8619
rect 10680 8590 10736 8592
rect 10680 8589 10717 8590
rect 10792 8589 10829 8599
rect 10888 8619 11036 8629
rect 11136 8626 11232 8628
rect 10888 8599 10897 8619
rect 10917 8599 11007 8619
rect 11027 8599 11036 8619
rect 10888 8590 11036 8599
rect 11094 8619 11232 8626
rect 11094 8599 11103 8619
rect 11123 8599 11232 8619
rect 11094 8590 11232 8599
rect 10888 8589 10925 8590
rect 10944 8538 10980 8590
rect 10999 8589 11036 8590
rect 11095 8589 11132 8590
rect 10415 8536 10456 8537
rect 10307 8529 10456 8536
rect 10307 8509 10425 8529
rect 10445 8509 10456 8529
rect 10307 8501 10456 8509
rect 10523 8533 10882 8537
rect 10523 8528 10845 8533
rect 10523 8504 10636 8528
rect 10660 8509 10845 8528
rect 10869 8509 10882 8533
rect 10660 8504 10882 8509
rect 10523 8501 10882 8504
rect 10944 8501 10979 8538
rect 11047 8535 11147 8538
rect 11047 8531 11114 8535
rect 11047 8505 11059 8531
rect 11085 8509 11114 8531
rect 11140 8509 11147 8535
rect 11085 8505 11147 8509
rect 11047 8501 11147 8505
rect 10523 8480 10554 8501
rect 10944 8480 10980 8501
rect 10366 8479 10403 8480
rect 10365 8470 10403 8479
rect 10365 8450 10374 8470
rect 10394 8450 10403 8470
rect 10365 8442 10403 8450
rect 10469 8474 10554 8480
rect 10579 8479 10616 8480
rect 10469 8454 10477 8474
rect 10497 8454 10554 8474
rect 10469 8446 10554 8454
rect 10578 8470 10616 8479
rect 10578 8450 10587 8470
rect 10607 8450 10616 8470
rect 10469 8445 10505 8446
rect 10578 8442 10616 8450
rect 10682 8474 10767 8480
rect 10787 8479 10824 8480
rect 10682 8454 10690 8474
rect 10710 8473 10767 8474
rect 10710 8454 10739 8473
rect 10682 8453 10739 8454
rect 10760 8453 10767 8473
rect 10682 8446 10767 8453
rect 10786 8470 10824 8479
rect 10786 8450 10795 8470
rect 10815 8450 10824 8470
rect 10682 8445 10718 8446
rect 10786 8442 10824 8450
rect 10890 8474 11034 8480
rect 10890 8454 10898 8474
rect 10918 8471 11006 8474
rect 10918 8454 10949 8471
rect 10890 8451 10949 8454
rect 10972 8454 11006 8471
rect 11026 8454 11034 8474
rect 10972 8451 11034 8454
rect 10890 8446 11034 8451
rect 10890 8445 10926 8446
rect 10998 8445 11034 8446
rect 11100 8479 11137 8480
rect 11100 8478 11138 8479
rect 11100 8470 11164 8478
rect 11100 8450 11109 8470
rect 11129 8456 11164 8470
rect 11184 8456 11187 8476
rect 11129 8451 11187 8456
rect 11129 8450 11164 8451
rect 10366 8413 10403 8442
rect 10367 8411 10403 8413
rect 10579 8411 10616 8442
rect 10367 8389 10616 8411
rect 10787 8410 10824 8442
rect 11100 8438 11164 8450
rect 11204 8412 11231 8590
rect 13759 8568 13786 8746
rect 13826 8708 13890 8720
rect 14166 8716 14203 8748
rect 14374 8747 14623 8769
rect 14664 8748 14850 8780
rect 14678 8747 14850 8748
rect 14374 8716 14411 8747
rect 14587 8745 14623 8747
rect 14587 8716 14624 8745
rect 14816 8719 14850 8747
rect 15194 8767 15234 8815
rect 16360 8821 16398 8830
rect 16360 8801 16369 8821
rect 16389 8801 16398 8821
rect 16360 8793 16398 8801
rect 16464 8825 16549 8831
rect 16574 8830 16611 8831
rect 16464 8805 16472 8825
rect 16492 8805 16549 8825
rect 16464 8797 16549 8805
rect 16573 8821 16611 8830
rect 16573 8801 16582 8821
rect 16602 8801 16611 8821
rect 16464 8796 16500 8797
rect 16573 8793 16611 8801
rect 16677 8825 16762 8831
rect 16782 8830 16819 8831
rect 16677 8805 16685 8825
rect 16705 8824 16762 8825
rect 16705 8805 16734 8824
rect 16677 8804 16734 8805
rect 16755 8804 16762 8824
rect 16677 8797 16762 8804
rect 16781 8821 16819 8830
rect 16781 8801 16790 8821
rect 16810 8801 16819 8821
rect 16677 8796 16713 8797
rect 16781 8793 16819 8801
rect 16885 8825 17029 8831
rect 16885 8805 16893 8825
rect 16913 8808 16949 8825
rect 16969 8808 17001 8825
rect 16913 8805 17001 8808
rect 17021 8805 17029 8825
rect 16885 8797 17029 8805
rect 16885 8796 16921 8797
rect 16993 8796 17029 8797
rect 17095 8830 17132 8831
rect 17095 8829 17133 8830
rect 17095 8821 17159 8829
rect 17095 8801 17104 8821
rect 17124 8807 17159 8821
rect 17179 8807 17182 8827
rect 17124 8802 17182 8807
rect 17124 8801 17159 8802
rect 15505 8771 15615 8785
rect 15505 8768 15548 8771
rect 15194 8760 15319 8767
rect 15505 8763 15509 8768
rect 15194 8741 15286 8760
rect 15311 8741 15319 8760
rect 15194 8731 15319 8741
rect 15427 8741 15509 8763
rect 15538 8741 15548 8768
rect 15576 8744 15583 8771
rect 15612 8763 15615 8771
rect 16361 8764 16398 8793
rect 15612 8744 15677 8763
rect 16362 8762 16398 8764
rect 16574 8762 16611 8793
rect 16782 8766 16819 8793
rect 17095 8789 17159 8801
rect 15576 8741 15677 8744
rect 15427 8739 15677 8741
rect 13826 8707 13861 8708
rect 13803 8702 13861 8707
rect 13803 8682 13806 8702
rect 13826 8688 13861 8702
rect 13881 8688 13890 8708
rect 13826 8680 13890 8688
rect 13852 8679 13890 8680
rect 13853 8678 13890 8679
rect 13956 8712 13992 8713
rect 14064 8712 14100 8713
rect 13956 8705 14100 8712
rect 13956 8704 14016 8705
rect 13956 8684 13964 8704
rect 13984 8685 14016 8704
rect 14041 8704 14100 8705
rect 14041 8685 14072 8704
rect 13984 8684 14072 8685
rect 14092 8684 14100 8704
rect 13956 8678 14100 8684
rect 14166 8708 14204 8716
rect 14272 8712 14308 8713
rect 14166 8688 14175 8708
rect 14195 8688 14204 8708
rect 14166 8679 14204 8688
rect 14223 8705 14308 8712
rect 14223 8685 14230 8705
rect 14251 8704 14308 8705
rect 14251 8685 14280 8704
rect 14223 8684 14280 8685
rect 14300 8684 14308 8704
rect 14166 8678 14203 8679
rect 14223 8678 14308 8684
rect 14374 8708 14412 8716
rect 14485 8712 14521 8713
rect 14374 8688 14383 8708
rect 14403 8688 14412 8708
rect 14374 8679 14412 8688
rect 14436 8704 14521 8712
rect 14436 8684 14493 8704
rect 14513 8684 14521 8704
rect 14374 8678 14411 8679
rect 14436 8678 14521 8684
rect 14587 8708 14625 8716
rect 14587 8688 14596 8708
rect 14616 8688 14625 8708
rect 14587 8679 14625 8688
rect 14814 8709 14851 8719
rect 15194 8711 15234 8731
rect 14814 8691 14824 8709
rect 14842 8691 14851 8709
rect 14814 8682 14851 8691
rect 15193 8702 15234 8711
rect 15193 8684 15203 8702
rect 15221 8684 15234 8702
rect 14816 8681 14850 8682
rect 14587 8678 14624 8679
rect 14010 8657 14046 8678
rect 14436 8657 14467 8678
rect 15193 8675 15234 8684
rect 15193 8674 15230 8675
rect 15427 8660 15464 8739
rect 15505 8726 15615 8739
rect 15579 8670 15610 8671
rect 13843 8653 13943 8657
rect 13843 8649 13905 8653
rect 13843 8623 13850 8649
rect 13876 8627 13905 8649
rect 13931 8627 13943 8653
rect 13876 8623 13943 8627
rect 13843 8620 13943 8623
rect 14011 8620 14046 8657
rect 14108 8654 14467 8657
rect 14108 8649 14330 8654
rect 14108 8625 14121 8649
rect 14145 8630 14330 8649
rect 14354 8630 14467 8654
rect 14145 8625 14467 8630
rect 14108 8621 14467 8625
rect 14534 8649 14683 8657
rect 14534 8629 14545 8649
rect 14565 8629 14683 8649
rect 15427 8640 15436 8660
rect 15456 8640 15464 8660
rect 15427 8630 15464 8640
rect 15523 8660 15610 8670
rect 15523 8640 15532 8660
rect 15552 8640 15610 8660
rect 15523 8631 15610 8640
rect 15523 8630 15560 8631
rect 14534 8622 14683 8629
rect 14534 8621 14575 8622
rect 13858 8568 13895 8569
rect 13954 8568 13991 8569
rect 14010 8568 14046 8620
rect 14065 8568 14102 8569
rect 13758 8559 13896 8568
rect 13353 8538 13464 8553
rect 13353 8536 13395 8538
rect 13023 8515 13128 8517
rect 12679 8507 12849 8508
rect 13023 8507 13072 8515
rect 12679 8488 13072 8507
rect 13103 8488 13128 8515
rect 13353 8516 13360 8536
rect 13379 8516 13395 8536
rect 13353 8508 13395 8516
rect 13423 8536 13464 8538
rect 13423 8516 13437 8536
rect 13456 8516 13464 8536
rect 13758 8539 13867 8559
rect 13887 8539 13896 8559
rect 13758 8532 13896 8539
rect 13954 8559 14102 8568
rect 13954 8539 13963 8559
rect 13983 8539 14073 8559
rect 14093 8539 14102 8559
rect 13758 8530 13854 8532
rect 13954 8529 14102 8539
rect 14161 8559 14198 8569
rect 14273 8568 14310 8569
rect 14254 8566 14310 8568
rect 14161 8539 14169 8559
rect 14189 8539 14198 8559
rect 14010 8528 14046 8529
rect 13423 8508 13464 8516
rect 13353 8502 13464 8508
rect 12679 8481 13128 8488
rect 12679 8479 12849 8481
rect 11529 8448 11639 8462
rect 11529 8445 11572 8448
rect 11529 8440 11533 8445
rect 11063 8410 11231 8412
rect 10787 8407 11231 8410
rect 10448 8383 10559 8389
rect 10448 8375 10489 8383
rect 10137 8320 10176 8364
rect 10448 8355 10456 8375
rect 10475 8355 10489 8375
rect 10448 8353 10489 8355
rect 10517 8375 10559 8383
rect 10517 8355 10533 8375
rect 10552 8355 10559 8375
rect 10517 8353 10559 8355
rect 10448 8338 10559 8353
rect 10785 8384 11231 8407
rect 10137 8296 10177 8320
rect 10477 8296 10524 8298
rect 10785 8296 10823 8384
rect 11063 8383 11231 8384
rect 11451 8418 11533 8440
rect 11562 8418 11572 8445
rect 11600 8421 11607 8448
rect 11636 8440 11639 8448
rect 11636 8421 11701 8440
rect 11600 8418 11701 8421
rect 11451 8416 11701 8418
rect 11451 8337 11488 8416
rect 11529 8403 11639 8416
rect 11603 8347 11634 8348
rect 11451 8317 11460 8337
rect 11480 8317 11488 8337
rect 11451 8307 11488 8317
rect 11547 8337 11634 8347
rect 11547 8317 11556 8337
rect 11576 8317 11634 8337
rect 11547 8308 11634 8317
rect 11547 8307 11584 8308
rect 10137 8263 10823 8296
rect 10137 8206 10176 8263
rect 10785 8261 10823 8263
rect 11603 8255 11634 8308
rect 11664 8337 11701 8416
rect 11872 8429 12265 8433
rect 11872 8412 11891 8429
rect 11911 8413 12265 8429
rect 12285 8413 12288 8433
rect 11911 8412 12288 8413
rect 11872 8408 12288 8412
rect 11872 8407 12213 8408
rect 11816 8347 11847 8348
rect 11664 8317 11673 8337
rect 11693 8317 11701 8337
rect 11664 8307 11701 8317
rect 11760 8340 11847 8347
rect 11760 8337 11821 8340
rect 11760 8317 11769 8337
rect 11789 8320 11821 8337
rect 11842 8320 11847 8340
rect 11789 8317 11847 8320
rect 11760 8310 11847 8317
rect 11872 8337 11909 8407
rect 12175 8406 12212 8407
rect 12024 8347 12060 8348
rect 11872 8317 11881 8337
rect 11901 8317 11909 8337
rect 11760 8308 11816 8310
rect 11760 8307 11797 8308
rect 11872 8307 11909 8317
rect 11968 8337 12116 8347
rect 12216 8344 12312 8346
rect 11968 8317 11977 8337
rect 11997 8317 12087 8337
rect 12107 8317 12116 8337
rect 11968 8308 12116 8317
rect 12174 8337 12312 8344
rect 12174 8317 12183 8337
rect 12203 8317 12312 8337
rect 12174 8308 12312 8317
rect 11968 8307 12005 8308
rect 12024 8256 12060 8308
rect 12079 8307 12116 8308
rect 12175 8307 12212 8308
rect 11495 8254 11536 8255
rect 11387 8247 11536 8254
rect 11387 8227 11505 8247
rect 11525 8227 11536 8247
rect 11387 8219 11536 8227
rect 11603 8251 11962 8255
rect 11603 8246 11925 8251
rect 11603 8222 11716 8246
rect 11740 8227 11925 8246
rect 11949 8227 11962 8251
rect 11740 8222 11962 8227
rect 11603 8219 11962 8222
rect 12024 8219 12059 8256
rect 12127 8253 12227 8256
rect 12127 8249 12194 8253
rect 12127 8223 12139 8249
rect 12165 8227 12194 8249
rect 12220 8227 12227 8253
rect 12165 8223 12227 8227
rect 12127 8219 12227 8223
rect 10137 8204 10185 8206
rect 10137 8186 10148 8204
rect 10166 8186 10185 8204
rect 11603 8198 11634 8219
rect 12024 8198 12060 8219
rect 11446 8197 11483 8198
rect 10137 8177 10185 8186
rect 10138 8176 10185 8177
rect 10451 8181 10561 8195
rect 10451 8178 10494 8181
rect 10451 8173 10455 8178
rect 10373 8151 10455 8173
rect 10484 8151 10494 8178
rect 10522 8154 10529 8181
rect 10558 8173 10561 8181
rect 11445 8188 11483 8197
rect 10558 8154 10623 8173
rect 11445 8168 11454 8188
rect 11474 8168 11483 8188
rect 10522 8151 10623 8154
rect 10373 8149 10623 8151
rect 10141 8113 10178 8114
rect 9840 8083 9850 8101
rect 9868 8083 9880 8101
rect 9840 8078 9880 8083
rect 10137 8110 10178 8113
rect 10137 8105 10179 8110
rect 10137 8087 10150 8105
rect 10168 8087 10179 8105
rect 9840 8074 9877 8078
rect 10137 8073 10179 8087
rect 10217 8073 10264 8077
rect 10137 8067 10264 8073
rect 9513 8055 9550 8056
rect 9463 8046 9550 8055
rect 9463 8026 9521 8046
rect 9541 8026 9550 8046
rect 9463 8016 9550 8026
rect 9609 8046 9646 8056
rect 9609 8026 9617 8046
rect 9637 8026 9646 8046
rect 9463 8015 9494 8016
rect 9458 7947 9568 7960
rect 9609 7947 9646 8026
rect 10137 8038 10225 8067
rect 10254 8038 10264 8067
rect 10373 8070 10410 8149
rect 10451 8136 10561 8149
rect 10525 8080 10556 8081
rect 10373 8050 10382 8070
rect 10402 8050 10410 8070
rect 10373 8040 10410 8050
rect 10469 8070 10556 8080
rect 10469 8050 10478 8070
rect 10498 8050 10556 8070
rect 10469 8041 10556 8050
rect 10469 8040 10506 8041
rect 10137 8034 10264 8038
rect 10137 8017 10176 8034
rect 10217 8033 10264 8034
rect 9843 8011 9880 8012
rect 9839 8002 9880 8011
rect 9839 7984 9852 8002
rect 9870 7984 9880 8002
rect 10137 7999 10148 8017
rect 10166 7999 10176 8017
rect 10137 7990 10176 7999
rect 10138 7989 10175 7990
rect 10525 7988 10556 8041
rect 10586 8070 10623 8149
rect 10794 8146 11187 8166
rect 11207 8146 11210 8166
rect 11445 8160 11483 8168
rect 11549 8192 11634 8198
rect 11659 8197 11696 8198
rect 11549 8172 11557 8192
rect 11577 8172 11634 8192
rect 11549 8164 11634 8172
rect 11658 8188 11696 8197
rect 11658 8168 11667 8188
rect 11687 8168 11696 8188
rect 11549 8163 11585 8164
rect 11658 8160 11696 8168
rect 11762 8192 11847 8198
rect 11867 8197 11904 8198
rect 11762 8172 11770 8192
rect 11790 8191 11847 8192
rect 11790 8172 11819 8191
rect 11762 8171 11819 8172
rect 11840 8171 11847 8191
rect 11762 8164 11847 8171
rect 11866 8188 11904 8197
rect 11866 8168 11875 8188
rect 11895 8168 11904 8188
rect 11762 8163 11798 8164
rect 11866 8160 11904 8168
rect 11970 8192 12114 8198
rect 11970 8172 11978 8192
rect 11998 8190 12086 8192
rect 11998 8172 12027 8190
rect 11970 8169 12027 8172
rect 12054 8172 12086 8190
rect 12106 8172 12114 8192
rect 12054 8169 12114 8172
rect 11970 8164 12114 8169
rect 11970 8163 12006 8164
rect 12078 8163 12114 8164
rect 12180 8197 12217 8198
rect 12180 8196 12218 8197
rect 12180 8188 12244 8196
rect 12180 8168 12189 8188
rect 12209 8174 12244 8188
rect 12264 8174 12267 8194
rect 12209 8169 12267 8174
rect 12209 8168 12244 8169
rect 10794 8141 11210 8146
rect 10794 8140 11135 8141
rect 10738 8080 10769 8081
rect 10586 8050 10595 8070
rect 10615 8050 10623 8070
rect 10586 8040 10623 8050
rect 10682 8073 10769 8080
rect 10682 8070 10743 8073
rect 10682 8050 10691 8070
rect 10711 8053 10743 8070
rect 10764 8053 10769 8073
rect 10711 8050 10769 8053
rect 10682 8043 10769 8050
rect 10794 8070 10831 8140
rect 11097 8139 11134 8140
rect 11446 8131 11483 8160
rect 11447 8129 11483 8131
rect 11659 8129 11696 8160
rect 11447 8107 11696 8129
rect 11867 8128 11904 8160
rect 12180 8156 12244 8168
rect 12284 8130 12311 8308
rect 12679 8301 12708 8479
rect 12748 8441 12812 8453
rect 13088 8449 13125 8481
rect 13296 8480 13545 8502
rect 13296 8449 13333 8480
rect 13509 8478 13545 8480
rect 13509 8449 13546 8478
rect 13858 8469 13895 8470
rect 14161 8469 14198 8539
rect 14223 8559 14310 8566
rect 14223 8556 14281 8559
rect 14223 8536 14228 8556
rect 14249 8539 14281 8556
rect 14301 8539 14310 8559
rect 14249 8536 14310 8539
rect 14223 8529 14310 8536
rect 14369 8559 14406 8569
rect 14369 8539 14377 8559
rect 14397 8539 14406 8559
rect 14223 8528 14254 8529
rect 13857 8468 14198 8469
rect 13782 8463 14198 8468
rect 12748 8440 12783 8441
rect 12725 8435 12783 8440
rect 12725 8415 12728 8435
rect 12748 8421 12783 8435
rect 12803 8421 12812 8441
rect 12748 8413 12812 8421
rect 12774 8412 12812 8413
rect 12775 8411 12812 8412
rect 12878 8445 12914 8446
rect 12986 8445 13022 8446
rect 12878 8437 13022 8445
rect 12878 8417 12886 8437
rect 12906 8417 12994 8437
rect 13014 8417 13022 8437
rect 12878 8411 13022 8417
rect 13088 8441 13126 8449
rect 13194 8445 13230 8446
rect 13088 8421 13097 8441
rect 13117 8421 13126 8441
rect 13088 8412 13126 8421
rect 13145 8438 13230 8445
rect 13145 8418 13152 8438
rect 13173 8437 13230 8438
rect 13173 8418 13202 8437
rect 13145 8417 13202 8418
rect 13222 8417 13230 8437
rect 13088 8411 13125 8412
rect 13145 8411 13230 8417
rect 13296 8441 13334 8449
rect 13407 8445 13443 8446
rect 13296 8421 13305 8441
rect 13325 8421 13334 8441
rect 13296 8412 13334 8421
rect 13358 8437 13443 8445
rect 13358 8417 13415 8437
rect 13435 8417 13443 8437
rect 13296 8411 13333 8412
rect 13358 8411 13443 8417
rect 13509 8441 13547 8449
rect 13782 8443 13785 8463
rect 13805 8443 14198 8463
rect 14369 8460 14406 8539
rect 14436 8568 14467 8621
rect 14817 8619 14854 8620
rect 14816 8610 14855 8619
rect 14816 8592 14826 8610
rect 14844 8592 14855 8610
rect 15196 8608 15233 8612
rect 14728 8575 14775 8576
rect 14816 8575 14855 8592
rect 14728 8571 14855 8575
rect 14486 8568 14523 8569
rect 14436 8559 14523 8568
rect 14436 8539 14494 8559
rect 14514 8539 14523 8559
rect 14436 8529 14523 8539
rect 14582 8559 14619 8569
rect 14582 8539 14590 8559
rect 14610 8539 14619 8559
rect 14436 8528 14467 8529
rect 14431 8460 14541 8473
rect 14582 8460 14619 8539
rect 14728 8542 14738 8571
rect 14767 8542 14855 8571
rect 14728 8536 14855 8542
rect 14728 8532 14775 8536
rect 14813 8522 14855 8536
rect 14813 8504 14824 8522
rect 14842 8504 14855 8522
rect 14813 8499 14855 8504
rect 14814 8496 14855 8499
rect 15193 8603 15233 8608
rect 15193 8585 15205 8603
rect 15223 8585 15233 8603
rect 14814 8495 14851 8496
rect 14369 8458 14619 8460
rect 14369 8455 14470 8458
rect 13509 8421 13518 8441
rect 13538 8421 13547 8441
rect 14369 8436 14434 8455
rect 13509 8412 13547 8421
rect 14431 8428 14434 8436
rect 14463 8428 14470 8455
rect 14498 8431 14508 8458
rect 14537 8436 14619 8458
rect 14537 8431 14541 8436
rect 14498 8428 14541 8431
rect 14431 8414 14541 8428
rect 14807 8432 14854 8433
rect 14807 8423 14855 8432
rect 13509 8411 13546 8412
rect 12932 8390 12968 8411
rect 13358 8390 13389 8411
rect 14807 8405 14826 8423
rect 14844 8405 14855 8423
rect 14807 8403 14855 8405
rect 12765 8386 12865 8390
rect 12765 8382 12827 8386
rect 12765 8356 12772 8382
rect 12798 8360 12827 8382
rect 12853 8360 12865 8386
rect 12798 8356 12865 8360
rect 12765 8353 12865 8356
rect 12933 8353 12968 8390
rect 13030 8387 13389 8390
rect 13030 8382 13252 8387
rect 13030 8358 13043 8382
rect 13067 8363 13252 8382
rect 13276 8363 13389 8387
rect 13067 8358 13389 8363
rect 13030 8354 13389 8358
rect 13456 8382 13605 8390
rect 13456 8362 13467 8382
rect 13487 8362 13605 8382
rect 13456 8355 13605 8362
rect 13456 8354 13497 8355
rect 12932 8314 12968 8353
rect 12780 8301 12817 8302
rect 12876 8301 12913 8302
rect 12932 8301 12939 8314
rect 12679 8292 12818 8301
rect 12679 8272 12789 8292
rect 12809 8272 12818 8292
rect 12679 8265 12818 8272
rect 12876 8292 12939 8301
rect 12876 8272 12885 8292
rect 12905 8276 12939 8292
rect 12962 8301 12968 8314
rect 12987 8301 13024 8302
rect 12962 8292 13024 8301
rect 12962 8276 12995 8292
rect 12905 8272 12995 8276
rect 13015 8272 13024 8292
rect 12679 8263 12776 8265
rect 12679 8262 12708 8263
rect 12876 8262 13024 8272
rect 13083 8292 13120 8302
rect 13195 8301 13232 8302
rect 13176 8299 13232 8301
rect 13083 8272 13091 8292
rect 13111 8272 13120 8292
rect 12932 8261 12968 8262
rect 12780 8202 12817 8203
rect 13083 8202 13120 8272
rect 13145 8292 13232 8299
rect 13145 8289 13203 8292
rect 13145 8269 13150 8289
rect 13171 8272 13203 8289
rect 13223 8272 13232 8292
rect 13171 8269 13232 8272
rect 13145 8262 13232 8269
rect 13291 8292 13328 8302
rect 13291 8272 13299 8292
rect 13319 8272 13328 8292
rect 13145 8261 13176 8262
rect 12779 8201 13120 8202
rect 12704 8197 13120 8201
rect 12704 8196 13081 8197
rect 12704 8176 12707 8196
rect 12727 8180 13081 8196
rect 13101 8180 13120 8197
rect 12727 8176 13120 8180
rect 13291 8193 13328 8272
rect 13358 8301 13389 8354
rect 14169 8346 14207 8348
rect 14816 8346 14855 8403
rect 14169 8313 14855 8346
rect 13408 8301 13445 8302
rect 13358 8292 13445 8301
rect 13358 8272 13416 8292
rect 13436 8272 13445 8292
rect 13358 8262 13445 8272
rect 13504 8292 13541 8302
rect 13504 8272 13512 8292
rect 13532 8272 13541 8292
rect 13358 8261 13389 8262
rect 13353 8193 13463 8206
rect 13504 8193 13541 8272
rect 13291 8191 13541 8193
rect 13291 8188 13392 8191
rect 13291 8169 13356 8188
rect 13353 8161 13356 8169
rect 13385 8161 13392 8188
rect 13420 8164 13430 8191
rect 13459 8169 13541 8191
rect 13761 8225 13929 8226
rect 14169 8225 14207 8313
rect 14468 8311 14515 8313
rect 14815 8289 14855 8313
rect 13761 8202 14207 8225
rect 14433 8256 14544 8271
rect 14433 8254 14475 8256
rect 14433 8234 14440 8254
rect 14459 8234 14475 8254
rect 14433 8226 14475 8234
rect 14503 8254 14544 8256
rect 14503 8234 14517 8254
rect 14536 8234 14544 8254
rect 14816 8245 14855 8289
rect 14503 8226 14544 8234
rect 14433 8220 14544 8226
rect 13761 8199 14205 8202
rect 13761 8197 13929 8199
rect 13459 8164 13463 8169
rect 13420 8161 13463 8164
rect 13353 8147 13463 8161
rect 12143 8128 12311 8130
rect 11864 8121 12311 8128
rect 11528 8101 11639 8107
rect 11528 8093 11569 8101
rect 10946 8080 10982 8081
rect 10794 8050 10803 8070
rect 10823 8050 10831 8070
rect 10682 8041 10738 8043
rect 10682 8040 10719 8041
rect 10794 8040 10831 8050
rect 10890 8070 11038 8080
rect 11138 8077 11234 8079
rect 10890 8050 10899 8070
rect 10919 8050 11009 8070
rect 11029 8050 11038 8070
rect 10890 8041 11038 8050
rect 11096 8070 11234 8077
rect 11096 8050 11105 8070
rect 11125 8050 11234 8070
rect 11528 8073 11536 8093
rect 11555 8073 11569 8093
rect 11528 8071 11569 8073
rect 11597 8093 11639 8101
rect 11597 8073 11613 8093
rect 11632 8073 11639 8093
rect 11864 8094 11889 8121
rect 11920 8102 12311 8121
rect 11920 8094 11969 8102
rect 12143 8101 12311 8102
rect 11864 8092 11969 8094
rect 11597 8071 11639 8073
rect 11528 8056 11639 8071
rect 11096 8041 11234 8050
rect 10890 8040 10927 8041
rect 10946 7989 10982 8041
rect 11001 8040 11038 8041
rect 11097 8040 11134 8041
rect 10417 7987 10458 7988
rect 9839 7975 9880 7984
rect 10309 7980 10458 7987
rect 9839 7955 9879 7975
rect 9396 7945 9646 7947
rect 9396 7942 9497 7945
rect 7914 7885 7978 7897
rect 8254 7893 8291 7920
rect 8462 7893 8499 7924
rect 8675 7922 8711 7924
rect 9396 7923 9461 7942
rect 8675 7893 8712 7922
rect 9458 7915 9461 7923
rect 9490 7915 9497 7942
rect 9525 7918 9535 7945
rect 9564 7923 9646 7945
rect 9754 7945 9879 7955
rect 10309 7960 10427 7980
rect 10447 7960 10458 7980
rect 10309 7952 10458 7960
rect 10525 7984 10884 7988
rect 10525 7979 10847 7984
rect 10525 7955 10638 7979
rect 10662 7960 10847 7979
rect 10871 7960 10884 7984
rect 10662 7955 10884 7960
rect 10525 7952 10884 7955
rect 10946 7952 10981 7989
rect 11049 7986 11149 7989
rect 11049 7982 11116 7986
rect 11049 7956 11061 7982
rect 11087 7960 11116 7982
rect 11142 7960 11149 7986
rect 11087 7956 11149 7960
rect 11049 7952 11149 7956
rect 9754 7926 9762 7945
rect 9787 7926 9879 7945
rect 10525 7931 10556 7952
rect 10946 7931 10982 7952
rect 10368 7930 10405 7931
rect 10142 7927 10176 7928
rect 9564 7918 9568 7923
rect 9754 7919 9879 7926
rect 9525 7915 9568 7918
rect 9458 7901 9568 7915
rect 7914 7884 7949 7885
rect 7891 7879 7949 7884
rect 7891 7859 7894 7879
rect 7914 7865 7949 7879
rect 7969 7865 7978 7885
rect 7914 7857 7978 7865
rect 7940 7856 7978 7857
rect 7941 7855 7978 7856
rect 8044 7889 8080 7890
rect 8152 7889 8188 7890
rect 8044 7881 8188 7889
rect 8044 7861 8052 7881
rect 8072 7878 8160 7881
rect 8072 7861 8104 7878
rect 8124 7861 8160 7878
rect 8180 7861 8188 7881
rect 8044 7855 8188 7861
rect 8254 7885 8292 7893
rect 8360 7889 8396 7890
rect 8254 7865 8263 7885
rect 8283 7865 8292 7885
rect 8254 7856 8292 7865
rect 8311 7882 8396 7889
rect 8311 7862 8318 7882
rect 8339 7881 8396 7882
rect 8339 7862 8368 7881
rect 8311 7861 8368 7862
rect 8388 7861 8396 7881
rect 8254 7855 8291 7856
rect 8311 7855 8396 7861
rect 8462 7885 8500 7893
rect 8573 7889 8609 7890
rect 8462 7865 8471 7885
rect 8491 7865 8500 7885
rect 8462 7856 8500 7865
rect 8524 7881 8609 7889
rect 8524 7861 8581 7881
rect 8601 7861 8609 7881
rect 8462 7855 8499 7856
rect 8524 7855 8609 7861
rect 8675 7885 8713 7893
rect 8675 7865 8684 7885
rect 8704 7865 8713 7885
rect 8675 7856 8713 7865
rect 9839 7871 9879 7919
rect 10141 7918 10178 7927
rect 10141 7900 10150 7918
rect 10168 7900 10178 7918
rect 10141 7890 10178 7900
rect 10367 7921 10405 7930
rect 10367 7901 10376 7921
rect 10396 7901 10405 7921
rect 10367 7893 10405 7901
rect 10471 7925 10556 7931
rect 10581 7930 10618 7931
rect 10471 7905 10479 7925
rect 10499 7905 10556 7925
rect 10471 7897 10556 7905
rect 10580 7921 10618 7930
rect 10580 7901 10589 7921
rect 10609 7901 10618 7921
rect 10471 7896 10507 7897
rect 10580 7893 10618 7901
rect 10684 7925 10769 7931
rect 10789 7930 10826 7931
rect 10684 7905 10692 7925
rect 10712 7924 10769 7925
rect 10712 7905 10741 7924
rect 10684 7904 10741 7905
rect 10762 7904 10769 7924
rect 10684 7897 10769 7904
rect 10788 7921 10826 7930
rect 10788 7901 10797 7921
rect 10817 7901 10826 7921
rect 10684 7896 10720 7897
rect 10788 7893 10826 7901
rect 10892 7925 11036 7931
rect 10892 7905 10900 7925
rect 10920 7924 11008 7925
rect 10920 7905 10951 7924
rect 10892 7904 10951 7905
rect 10976 7905 11008 7924
rect 11028 7905 11036 7925
rect 10976 7904 11036 7905
rect 10892 7897 11036 7904
rect 10892 7896 10928 7897
rect 11000 7896 11036 7897
rect 11102 7930 11139 7931
rect 11102 7929 11140 7930
rect 11102 7921 11166 7929
rect 11102 7901 11111 7921
rect 11131 7907 11166 7921
rect 11186 7907 11189 7927
rect 11131 7902 11189 7907
rect 11131 7901 11166 7902
rect 8675 7855 8712 7856
rect 8098 7834 8134 7855
rect 8524 7834 8555 7855
rect 9839 7853 9850 7871
rect 9868 7853 9879 7871
rect 9839 7845 9879 7853
rect 10142 7862 10176 7890
rect 10368 7864 10405 7893
rect 10369 7862 10405 7864
rect 10581 7862 10618 7893
rect 10142 7861 10314 7862
rect 9840 7844 9877 7845
rect 7931 7830 8031 7834
rect 7931 7826 7993 7830
rect 7931 7800 7938 7826
rect 7964 7804 7993 7826
rect 8019 7804 8031 7830
rect 7964 7800 8031 7804
rect 7931 7797 8031 7800
rect 8099 7797 8134 7834
rect 8196 7831 8555 7834
rect 8196 7826 8418 7831
rect 8196 7802 8209 7826
rect 8233 7807 8418 7826
rect 8442 7807 8555 7831
rect 8233 7802 8555 7807
rect 8196 7798 8555 7802
rect 8622 7826 8771 7834
rect 8622 7806 8633 7826
rect 8653 7806 8771 7826
rect 8622 7799 8771 7806
rect 10142 7829 10328 7861
rect 10369 7840 10618 7862
rect 10789 7861 10826 7893
rect 11102 7889 11166 7901
rect 11206 7863 11233 8041
rect 13761 8019 13788 8197
rect 13828 8159 13892 8171
rect 14168 8167 14205 8199
rect 14376 8198 14625 8220
rect 14376 8167 14413 8198
rect 14589 8196 14625 8198
rect 14589 8167 14626 8196
rect 13828 8158 13863 8159
rect 13805 8153 13863 8158
rect 13805 8133 13808 8153
rect 13828 8139 13863 8153
rect 13883 8139 13892 8159
rect 13828 8131 13892 8139
rect 13854 8130 13892 8131
rect 13855 8129 13892 8130
rect 13958 8163 13994 8164
rect 14066 8163 14102 8164
rect 13958 8158 14102 8163
rect 13958 8155 14020 8158
rect 13958 8135 13966 8155
rect 13986 8138 14020 8155
rect 14043 8155 14102 8158
rect 14043 8138 14074 8155
rect 13986 8135 14074 8138
rect 14094 8135 14102 8155
rect 13958 8129 14102 8135
rect 14168 8159 14206 8167
rect 14274 8163 14310 8164
rect 14168 8139 14177 8159
rect 14197 8139 14206 8159
rect 14168 8130 14206 8139
rect 14225 8156 14310 8163
rect 14225 8136 14232 8156
rect 14253 8155 14310 8156
rect 14253 8136 14282 8155
rect 14225 8135 14282 8136
rect 14302 8135 14310 8155
rect 14168 8129 14205 8130
rect 14225 8129 14310 8135
rect 14376 8159 14414 8167
rect 14487 8163 14523 8164
rect 14376 8139 14385 8159
rect 14405 8139 14414 8159
rect 14376 8130 14414 8139
rect 14438 8155 14523 8163
rect 14438 8135 14495 8155
rect 14515 8135 14523 8155
rect 14376 8129 14413 8130
rect 14438 8129 14523 8135
rect 14589 8159 14627 8167
rect 14589 8139 14598 8159
rect 14618 8139 14627 8159
rect 14589 8130 14627 8139
rect 14589 8129 14626 8130
rect 14012 8108 14048 8129
rect 14438 8108 14469 8129
rect 13845 8104 13945 8108
rect 13845 8100 13907 8104
rect 13845 8074 13852 8100
rect 13878 8078 13907 8100
rect 13933 8078 13945 8104
rect 13878 8074 13945 8078
rect 13845 8071 13945 8074
rect 14013 8071 14048 8108
rect 14110 8105 14469 8108
rect 14110 8100 14332 8105
rect 14110 8076 14123 8100
rect 14147 8081 14332 8100
rect 14356 8081 14469 8105
rect 14147 8076 14469 8081
rect 14110 8072 14469 8076
rect 14536 8100 14685 8108
rect 14536 8080 14547 8100
rect 14567 8080 14685 8100
rect 14536 8073 14685 8080
rect 14536 8072 14577 8073
rect 13860 8019 13897 8020
rect 13956 8019 13993 8020
rect 14012 8019 14048 8071
rect 14067 8019 14104 8020
rect 13760 8010 13898 8019
rect 13760 7990 13869 8010
rect 13889 7990 13898 8010
rect 13760 7983 13898 7990
rect 13956 8010 14104 8019
rect 13956 7990 13965 8010
rect 13985 7990 14075 8010
rect 14095 7990 14104 8010
rect 13760 7981 13856 7983
rect 13956 7980 14104 7990
rect 14163 8010 14200 8020
rect 14275 8019 14312 8020
rect 14256 8017 14312 8019
rect 14163 7990 14171 8010
rect 14191 7990 14200 8010
rect 14012 7979 14048 7980
rect 11389 7937 11499 7951
rect 11389 7934 11432 7937
rect 11389 7929 11393 7934
rect 11065 7861 11233 7863
rect 10789 7855 11233 7861
rect 9211 7803 9725 7804
rect 8622 7798 8663 7799
rect 7946 7745 7983 7746
rect 8042 7745 8079 7746
rect 8098 7745 8134 7797
rect 8153 7745 8190 7746
rect 7846 7736 7984 7745
rect 7846 7716 7955 7736
rect 7975 7716 7984 7736
rect 7846 7709 7984 7716
rect 8042 7736 8190 7745
rect 8042 7716 8051 7736
rect 8071 7716 8161 7736
rect 8181 7716 8190 7736
rect 7846 7707 7942 7709
rect 8042 7706 8190 7716
rect 8249 7736 8286 7746
rect 8361 7745 8398 7746
rect 8342 7743 8398 7745
rect 8249 7716 8257 7736
rect 8277 7716 8286 7736
rect 8098 7705 8134 7706
rect 7028 7653 7196 7655
rect 6750 7647 7196 7653
rect 5818 7623 6234 7628
rect 6413 7626 6524 7632
rect 5818 7622 6159 7623
rect 5762 7562 5793 7563
rect 5610 7532 5619 7552
rect 5639 7532 5647 7552
rect 5610 7522 5647 7532
rect 5706 7555 5793 7562
rect 5706 7552 5767 7555
rect 5706 7532 5715 7552
rect 5735 7535 5767 7552
rect 5788 7535 5793 7555
rect 5735 7532 5793 7535
rect 5706 7525 5793 7532
rect 5818 7552 5855 7622
rect 6121 7621 6158 7622
rect 6413 7618 6454 7626
rect 6413 7598 6421 7618
rect 6440 7598 6454 7618
rect 6413 7596 6454 7598
rect 6482 7618 6524 7626
rect 6482 7598 6498 7618
rect 6517 7598 6524 7618
rect 6750 7625 6756 7647
rect 6782 7627 7196 7647
rect 7946 7646 7983 7647
rect 8249 7646 8286 7716
rect 8311 7736 8398 7743
rect 8311 7733 8369 7736
rect 8311 7713 8316 7733
rect 8337 7716 8369 7733
rect 8389 7716 8398 7736
rect 8337 7713 8398 7716
rect 8311 7706 8398 7713
rect 8457 7736 8494 7746
rect 8457 7716 8465 7736
rect 8485 7716 8494 7736
rect 8311 7705 8342 7706
rect 7945 7645 8286 7646
rect 6782 7625 6791 7627
rect 7028 7626 7196 7627
rect 7870 7640 8286 7645
rect 6750 7616 6791 7625
rect 7870 7620 7873 7640
rect 7893 7620 8286 7640
rect 8457 7637 8494 7716
rect 8524 7745 8555 7798
rect 9192 7787 9725 7803
rect 10142 7797 10176 7829
rect 10138 7788 10176 7797
rect 9192 7776 9724 7787
rect 9843 7778 9880 7782
rect 8574 7745 8611 7746
rect 8524 7736 8611 7745
rect 8524 7716 8582 7736
rect 8602 7716 8611 7736
rect 8524 7706 8611 7716
rect 8670 7736 8707 7746
rect 8670 7716 8678 7736
rect 8698 7716 8707 7736
rect 8524 7705 8555 7706
rect 8519 7637 8629 7650
rect 8670 7637 8707 7716
rect 8457 7635 8707 7637
rect 8457 7632 8558 7635
rect 8457 7613 8522 7632
rect 6482 7596 6524 7598
rect 6413 7581 6524 7596
rect 8519 7605 8522 7613
rect 8551 7605 8558 7632
rect 8586 7608 8596 7635
rect 8625 7613 8707 7635
rect 8785 7707 8953 7708
rect 9192 7707 9230 7776
rect 8785 7687 9230 7707
rect 9457 7738 9568 7753
rect 9457 7736 9499 7738
rect 9457 7716 9464 7736
rect 9483 7716 9499 7736
rect 9457 7708 9499 7716
rect 9527 7736 9568 7738
rect 9527 7716 9541 7736
rect 9560 7716 9568 7736
rect 9527 7708 9568 7716
rect 9457 7702 9568 7708
rect 9690 7713 9724 7776
rect 9842 7772 9880 7778
rect 9842 7754 9852 7772
rect 9870 7754 9880 7772
rect 10138 7770 10148 7788
rect 10166 7770 10176 7788
rect 10138 7764 10176 7770
rect 10294 7766 10328 7829
rect 10450 7834 10561 7840
rect 10450 7826 10491 7834
rect 10450 7806 10458 7826
rect 10477 7806 10491 7826
rect 10450 7804 10491 7806
rect 10519 7826 10561 7834
rect 10519 7806 10535 7826
rect 10554 7806 10561 7826
rect 10519 7804 10561 7806
rect 10450 7789 10561 7804
rect 10788 7835 11233 7855
rect 10788 7766 10826 7835
rect 11065 7834 11233 7835
rect 11311 7907 11393 7929
rect 11422 7907 11432 7934
rect 11460 7910 11467 7937
rect 11496 7929 11499 7937
rect 13494 7946 13605 7961
rect 13494 7944 13536 7946
rect 11496 7910 11561 7929
rect 11460 7907 11561 7910
rect 11311 7905 11561 7907
rect 11311 7826 11348 7905
rect 11389 7892 11499 7905
rect 11463 7836 11494 7837
rect 11311 7806 11320 7826
rect 11340 7806 11348 7826
rect 11311 7796 11348 7806
rect 11407 7826 11494 7836
rect 11407 7806 11416 7826
rect 11436 7806 11494 7826
rect 11407 7797 11494 7806
rect 11407 7796 11444 7797
rect 10138 7760 10175 7764
rect 10294 7755 10826 7766
rect 9842 7745 9880 7754
rect 9842 7713 9876 7745
rect 10293 7739 10826 7755
rect 11463 7744 11494 7797
rect 11524 7826 11561 7905
rect 11732 7915 12125 7922
rect 11732 7898 11740 7915
rect 11772 7902 12125 7915
rect 12145 7902 12148 7922
rect 13227 7917 13268 7926
rect 11772 7898 12148 7902
rect 11732 7897 12148 7898
rect 12822 7915 12990 7916
rect 13227 7915 13236 7917
rect 11732 7896 12073 7897
rect 11676 7836 11707 7837
rect 11524 7806 11533 7826
rect 11553 7806 11561 7826
rect 11524 7796 11561 7806
rect 11620 7829 11707 7836
rect 11620 7826 11681 7829
rect 11620 7806 11629 7826
rect 11649 7809 11681 7826
rect 11702 7809 11707 7829
rect 11649 7806 11707 7809
rect 11620 7799 11707 7806
rect 11732 7826 11769 7896
rect 12035 7895 12072 7896
rect 12822 7895 13236 7915
rect 13262 7895 13268 7917
rect 13494 7924 13501 7944
rect 13520 7924 13536 7944
rect 13494 7916 13536 7924
rect 13564 7944 13605 7946
rect 13564 7924 13578 7944
rect 13597 7924 13605 7944
rect 13564 7916 13605 7924
rect 13860 7920 13897 7921
rect 14163 7920 14200 7990
rect 14225 8010 14312 8017
rect 14225 8007 14283 8010
rect 14225 7987 14230 8007
rect 14251 7990 14283 8007
rect 14303 7990 14312 8010
rect 14251 7987 14312 7990
rect 14225 7980 14312 7987
rect 14371 8010 14408 8020
rect 14371 7990 14379 8010
rect 14399 7990 14408 8010
rect 14225 7979 14256 7980
rect 13859 7919 14200 7920
rect 13494 7910 13605 7916
rect 13784 7914 14200 7919
rect 12822 7889 13268 7895
rect 12822 7887 12990 7889
rect 11884 7836 11920 7837
rect 11732 7806 11741 7826
rect 11761 7806 11769 7826
rect 11620 7797 11676 7799
rect 11620 7796 11657 7797
rect 11732 7796 11769 7806
rect 11828 7826 11976 7836
rect 12076 7833 12172 7835
rect 11828 7806 11837 7826
rect 11857 7821 11947 7826
rect 11857 7806 11892 7821
rect 11828 7797 11892 7806
rect 11828 7796 11865 7797
rect 11884 7780 11892 7797
rect 11913 7806 11947 7821
rect 11967 7806 11976 7826
rect 11913 7797 11976 7806
rect 12034 7826 12172 7833
rect 12034 7806 12043 7826
rect 12063 7806 12172 7826
rect 12034 7797 12172 7806
rect 11913 7780 11920 7797
rect 11939 7796 11976 7797
rect 12035 7796 12072 7797
rect 11884 7745 11920 7780
rect 11355 7743 11396 7744
rect 10293 7738 10807 7739
rect 8785 7681 9229 7687
rect 8785 7679 8953 7681
rect 8625 7608 8629 7613
rect 8586 7605 8629 7608
rect 8519 7591 8629 7605
rect 5970 7562 6006 7563
rect 5818 7532 5827 7552
rect 5847 7532 5855 7552
rect 5706 7523 5762 7525
rect 5706 7522 5743 7523
rect 5818 7522 5855 7532
rect 5914 7552 6062 7562
rect 6162 7559 6258 7561
rect 5914 7532 5923 7552
rect 5943 7532 6033 7552
rect 6053 7532 6062 7552
rect 5914 7523 6062 7532
rect 6120 7552 6258 7559
rect 6120 7532 6129 7552
rect 6149 7532 6258 7552
rect 6120 7523 6258 7532
rect 5914 7522 5951 7523
rect 5970 7471 6006 7523
rect 6025 7522 6062 7523
rect 6121 7522 6158 7523
rect 5441 7469 5482 7470
rect 5333 7462 5482 7469
rect 5333 7442 5451 7462
rect 5471 7442 5482 7462
rect 5333 7434 5482 7442
rect 5549 7466 5908 7470
rect 5549 7461 5871 7466
rect 5549 7437 5662 7461
rect 5686 7442 5871 7461
rect 5895 7442 5908 7466
rect 5686 7437 5908 7442
rect 5549 7434 5908 7437
rect 5970 7434 6005 7471
rect 6073 7468 6173 7471
rect 6073 7464 6140 7468
rect 6073 7438 6085 7464
rect 6111 7442 6140 7464
rect 6166 7442 6173 7468
rect 6111 7438 6173 7442
rect 6073 7434 6173 7438
rect 5549 7413 5580 7434
rect 5970 7413 6006 7434
rect 5392 7412 5429 7413
rect 5391 7403 5429 7412
rect 5391 7383 5400 7403
rect 5420 7383 5429 7403
rect 5391 7375 5429 7383
rect 5495 7407 5580 7413
rect 5605 7412 5642 7413
rect 5495 7387 5503 7407
rect 5523 7387 5580 7407
rect 5495 7379 5580 7387
rect 5604 7403 5642 7412
rect 5604 7383 5613 7403
rect 5633 7383 5642 7403
rect 5495 7378 5531 7379
rect 5604 7375 5642 7383
rect 5708 7407 5793 7413
rect 5813 7412 5850 7413
rect 5708 7387 5716 7407
rect 5736 7406 5793 7407
rect 5736 7387 5765 7406
rect 5708 7386 5765 7387
rect 5786 7386 5793 7406
rect 5708 7379 5793 7386
rect 5812 7403 5850 7412
rect 5812 7383 5821 7403
rect 5841 7383 5850 7403
rect 5708 7378 5744 7379
rect 5812 7375 5850 7383
rect 5916 7407 6060 7413
rect 5916 7387 5924 7407
rect 5944 7404 6032 7407
rect 5944 7387 5975 7404
rect 5916 7384 5975 7387
rect 5998 7387 6032 7404
rect 6052 7387 6060 7407
rect 5998 7384 6060 7387
rect 5916 7379 6060 7384
rect 5916 7378 5952 7379
rect 6024 7378 6060 7379
rect 6126 7412 6163 7413
rect 6126 7411 6164 7412
rect 6126 7403 6190 7411
rect 6126 7383 6135 7403
rect 6155 7389 6190 7403
rect 6210 7389 6213 7409
rect 6155 7384 6213 7389
rect 6155 7383 6190 7384
rect 5392 7346 5429 7375
rect 5393 7344 5429 7346
rect 5605 7344 5642 7375
rect 5393 7322 5642 7344
rect 5813 7343 5850 7375
rect 6126 7371 6190 7383
rect 6230 7345 6257 7523
rect 8785 7501 8812 7679
rect 8852 7641 8916 7653
rect 9192 7649 9229 7681
rect 9400 7680 9649 7702
rect 9690 7681 9876 7713
rect 11247 7736 11396 7743
rect 11247 7716 11365 7736
rect 11385 7716 11396 7736
rect 11247 7708 11396 7716
rect 11463 7740 11822 7744
rect 11463 7735 11785 7740
rect 11463 7711 11576 7735
rect 11600 7716 11785 7735
rect 11809 7716 11822 7740
rect 11600 7711 11822 7716
rect 11463 7708 11822 7711
rect 11884 7708 11919 7745
rect 11987 7742 12087 7745
rect 11987 7738 12054 7742
rect 11987 7712 11999 7738
rect 12025 7716 12054 7738
rect 12080 7716 12087 7742
rect 12025 7712 12087 7716
rect 11987 7708 12087 7712
rect 10141 7697 10178 7698
rect 9704 7680 9876 7681
rect 9400 7649 9437 7680
rect 9613 7678 9649 7680
rect 9613 7649 9650 7678
rect 9842 7652 9876 7680
rect 10139 7689 10179 7697
rect 10139 7671 10150 7689
rect 10168 7671 10179 7689
rect 11463 7687 11494 7708
rect 11884 7687 11920 7708
rect 11306 7686 11343 7687
rect 8852 7640 8887 7641
rect 8829 7635 8887 7640
rect 8829 7615 8832 7635
rect 8852 7621 8887 7635
rect 8907 7621 8916 7641
rect 8852 7613 8916 7621
rect 8878 7612 8916 7613
rect 8879 7611 8916 7612
rect 8982 7645 9018 7646
rect 9090 7645 9126 7646
rect 8982 7638 9126 7645
rect 8982 7637 9042 7638
rect 8982 7617 8990 7637
rect 9010 7618 9042 7637
rect 9067 7637 9126 7638
rect 9067 7618 9098 7637
rect 9010 7617 9098 7618
rect 9118 7617 9126 7637
rect 8982 7611 9126 7617
rect 9192 7641 9230 7649
rect 9298 7645 9334 7646
rect 9192 7621 9201 7641
rect 9221 7621 9230 7641
rect 9192 7612 9230 7621
rect 9249 7638 9334 7645
rect 9249 7618 9256 7638
rect 9277 7637 9334 7638
rect 9277 7618 9306 7637
rect 9249 7617 9306 7618
rect 9326 7617 9334 7637
rect 9192 7611 9229 7612
rect 9249 7611 9334 7617
rect 9400 7641 9438 7649
rect 9511 7645 9547 7646
rect 9400 7621 9409 7641
rect 9429 7621 9438 7641
rect 9400 7612 9438 7621
rect 9462 7637 9547 7645
rect 9462 7617 9519 7637
rect 9539 7617 9547 7637
rect 9400 7611 9437 7612
rect 9462 7611 9547 7617
rect 9613 7641 9651 7649
rect 9613 7621 9622 7641
rect 9642 7621 9651 7641
rect 9613 7612 9651 7621
rect 9840 7642 9877 7652
rect 9840 7624 9850 7642
rect 9868 7624 9877 7642
rect 9840 7615 9877 7624
rect 10139 7623 10179 7671
rect 11305 7677 11343 7686
rect 11305 7657 11314 7677
rect 11334 7657 11343 7677
rect 11305 7649 11343 7657
rect 11409 7681 11494 7687
rect 11519 7686 11556 7687
rect 11409 7661 11417 7681
rect 11437 7661 11494 7681
rect 11409 7653 11494 7661
rect 11518 7677 11556 7686
rect 11518 7657 11527 7677
rect 11547 7657 11556 7677
rect 11409 7652 11445 7653
rect 11518 7649 11556 7657
rect 11622 7681 11707 7687
rect 11727 7686 11764 7687
rect 11622 7661 11630 7681
rect 11650 7680 11707 7681
rect 11650 7661 11679 7680
rect 11622 7660 11679 7661
rect 11700 7660 11707 7680
rect 11622 7653 11707 7660
rect 11726 7677 11764 7686
rect 11726 7657 11735 7677
rect 11755 7657 11764 7677
rect 11622 7652 11658 7653
rect 11726 7649 11764 7657
rect 11830 7681 11974 7687
rect 11830 7661 11838 7681
rect 11858 7661 11946 7681
rect 11966 7661 11974 7681
rect 11830 7653 11974 7661
rect 11830 7652 11866 7653
rect 11938 7652 11974 7653
rect 12040 7686 12077 7687
rect 12040 7685 12078 7686
rect 12040 7677 12104 7685
rect 12040 7657 12049 7677
rect 12069 7663 12104 7677
rect 12124 7663 12127 7683
rect 12069 7658 12127 7663
rect 12069 7657 12104 7658
rect 10450 7627 10560 7641
rect 10450 7624 10493 7627
rect 10139 7616 10264 7623
rect 10450 7619 10454 7624
rect 9842 7614 9876 7615
rect 9613 7611 9650 7612
rect 9036 7590 9072 7611
rect 9462 7590 9493 7611
rect 10139 7597 10231 7616
rect 10256 7597 10264 7616
rect 8869 7586 8969 7590
rect 8869 7582 8931 7586
rect 8869 7556 8876 7582
rect 8902 7560 8931 7582
rect 8957 7560 8969 7586
rect 8902 7556 8969 7560
rect 8869 7553 8969 7556
rect 9037 7553 9072 7590
rect 9134 7587 9493 7590
rect 9134 7582 9356 7587
rect 9134 7558 9147 7582
rect 9171 7563 9356 7582
rect 9380 7563 9493 7587
rect 9171 7558 9493 7563
rect 9134 7554 9493 7558
rect 9560 7582 9709 7590
rect 9560 7562 9571 7582
rect 9591 7562 9709 7582
rect 10139 7587 10264 7597
rect 10372 7597 10454 7619
rect 10483 7597 10493 7624
rect 10521 7600 10528 7627
rect 10557 7619 10560 7627
rect 11306 7620 11343 7649
rect 10557 7600 10622 7619
rect 11307 7618 11343 7620
rect 11519 7618 11556 7649
rect 11727 7622 11764 7649
rect 12040 7645 12104 7657
rect 10521 7597 10622 7600
rect 10372 7595 10622 7597
rect 10139 7567 10179 7587
rect 9560 7555 9709 7562
rect 10138 7558 10179 7567
rect 9560 7554 9601 7555
rect 8884 7501 8921 7502
rect 8980 7501 9017 7502
rect 9036 7501 9072 7553
rect 9091 7501 9128 7502
rect 8784 7492 8922 7501
rect 8409 7458 8520 7473
rect 8784 7472 8893 7492
rect 8913 7472 8922 7492
rect 8784 7465 8922 7472
rect 8980 7492 9128 7501
rect 8980 7472 8989 7492
rect 9009 7472 9099 7492
rect 9119 7472 9128 7492
rect 8784 7463 8880 7465
rect 8980 7462 9128 7472
rect 9187 7492 9224 7502
rect 9299 7501 9336 7502
rect 9280 7499 9336 7501
rect 9187 7472 9195 7492
rect 9215 7472 9224 7492
rect 9036 7461 9072 7462
rect 8409 7456 8451 7458
rect 7746 7437 7816 7446
rect 7746 7428 7763 7437
rect 7737 7408 7763 7428
rect 7811 7428 7816 7437
rect 8409 7436 8416 7456
rect 8435 7436 8451 7456
rect 8409 7428 8451 7436
rect 8479 7456 8520 7458
rect 8479 7436 8493 7456
rect 8512 7436 8520 7456
rect 8479 7428 8520 7436
rect 7811 7427 7905 7428
rect 7811 7408 8181 7427
rect 8409 7422 8520 7428
rect 6524 7394 6634 7408
rect 6524 7391 6567 7394
rect 6524 7386 6528 7391
rect 6089 7343 6257 7345
rect 5813 7340 6257 7343
rect 5474 7316 5585 7322
rect 5474 7308 5515 7316
rect 5163 7253 5202 7297
rect 5474 7288 5482 7308
rect 5501 7288 5515 7308
rect 5474 7286 5515 7288
rect 5543 7308 5585 7316
rect 5543 7288 5559 7308
rect 5578 7288 5585 7308
rect 5543 7286 5585 7288
rect 5474 7272 5585 7286
rect 5811 7317 6257 7340
rect 3456 7233 3497 7234
rect 2932 7192 2968 7232
rect 2780 7180 2817 7181
rect 2876 7180 2913 7181
rect 2932 7180 2937 7192
rect 2680 7171 2818 7180
rect 2680 7151 2789 7171
rect 2809 7151 2818 7171
rect 2680 7144 2818 7151
rect 2876 7171 2937 7180
rect 2876 7151 2885 7171
rect 2905 7160 2937 7171
rect 2964 7180 2968 7192
rect 2987 7180 3024 7181
rect 2964 7171 3024 7180
rect 2964 7160 2995 7171
rect 2905 7151 2995 7160
rect 3015 7151 3024 7171
rect 2680 7142 2776 7144
rect 2876 7141 3024 7151
rect 3083 7171 3120 7181
rect 3195 7180 3232 7181
rect 3176 7178 3232 7180
rect 3083 7151 3091 7171
rect 3111 7151 3120 7171
rect 2932 7140 2968 7141
rect 2780 7081 2817 7082
rect 3083 7081 3120 7151
rect 3145 7171 3232 7178
rect 3145 7168 3203 7171
rect 3145 7148 3150 7168
rect 3171 7151 3203 7168
rect 3223 7151 3232 7171
rect 3171 7148 3232 7151
rect 3145 7141 3232 7148
rect 3291 7171 3328 7181
rect 3291 7151 3299 7171
rect 3319 7151 3328 7171
rect 3145 7140 3176 7141
rect 2779 7080 3120 7081
rect 2704 7075 3120 7080
rect 2704 7057 2707 7075
rect 2727 7073 3120 7075
rect 2727 7057 3097 7073
rect 2745 7055 3097 7057
rect 3088 7053 3097 7055
rect 3118 7053 3120 7073
rect 3088 7041 3120 7053
rect 3291 7072 3328 7151
rect 3358 7180 3389 7233
rect 4138 7205 4824 7238
rect 3408 7180 3445 7181
rect 3358 7171 3445 7180
rect 3358 7151 3416 7171
rect 3436 7151 3445 7171
rect 3358 7141 3445 7151
rect 3504 7171 3541 7181
rect 3504 7151 3512 7171
rect 3532 7151 3541 7171
rect 3358 7140 3389 7141
rect 3353 7072 3463 7085
rect 3504 7072 3541 7151
rect 3291 7070 3541 7072
rect 3291 7067 3392 7070
rect 3291 7048 3356 7067
rect 2131 7035 2250 7037
rect 2082 7033 2250 7035
rect 1467 7006 1578 7012
rect 1806 7007 2250 7033
rect 3353 7040 3356 7048
rect 3385 7040 3392 7067
rect 3420 7043 3430 7070
rect 3459 7048 3541 7070
rect 3730 7117 3898 7118
rect 4138 7117 4176 7205
rect 4437 7203 4484 7205
rect 4784 7181 4824 7205
rect 5163 7229 5203 7253
rect 5503 7229 5550 7231
rect 5811 7229 5849 7317
rect 6089 7316 6257 7317
rect 6446 7364 6528 7386
rect 6557 7364 6567 7391
rect 6595 7367 6602 7394
rect 6631 7386 6634 7394
rect 7737 7401 8181 7408
rect 7737 7399 7905 7401
rect 7737 7391 7816 7399
rect 6631 7367 6696 7386
rect 6595 7364 6696 7367
rect 6446 7362 6696 7364
rect 6446 7283 6483 7362
rect 6524 7349 6634 7362
rect 6598 7293 6629 7294
rect 6446 7263 6455 7283
rect 6475 7263 6483 7283
rect 6446 7253 6483 7263
rect 6542 7283 6629 7293
rect 6542 7263 6551 7283
rect 6571 7263 6629 7283
rect 6542 7254 6629 7263
rect 6542 7253 6579 7254
rect 5163 7196 5849 7229
rect 6598 7201 6629 7254
rect 6659 7283 6696 7362
rect 6867 7359 7260 7379
rect 7280 7359 7283 7379
rect 6867 7354 7283 7359
rect 6867 7353 7208 7354
rect 6811 7293 6842 7294
rect 6659 7263 6668 7283
rect 6688 7263 6696 7283
rect 6659 7253 6696 7263
rect 6755 7286 6842 7293
rect 6755 7283 6816 7286
rect 6755 7263 6764 7283
rect 6784 7266 6816 7283
rect 6837 7266 6842 7286
rect 6784 7263 6842 7266
rect 6755 7256 6842 7263
rect 6867 7283 6904 7353
rect 7170 7352 7207 7353
rect 7019 7293 7055 7294
rect 6867 7263 6876 7283
rect 6896 7263 6904 7283
rect 6755 7254 6811 7256
rect 6755 7253 6792 7254
rect 6867 7253 6904 7263
rect 6963 7283 7111 7293
rect 7211 7290 7307 7292
rect 6963 7263 6972 7283
rect 6992 7263 7082 7283
rect 7102 7263 7111 7283
rect 6963 7254 7111 7263
rect 7169 7283 7307 7290
rect 7169 7263 7178 7283
rect 7198 7263 7307 7283
rect 7169 7254 7307 7263
rect 6963 7253 7000 7254
rect 7019 7202 7055 7254
rect 7074 7253 7111 7254
rect 7170 7253 7207 7254
rect 6490 7200 6531 7201
rect 3730 7094 4176 7117
rect 4402 7148 4513 7162
rect 4402 7146 4444 7148
rect 4402 7126 4409 7146
rect 4428 7126 4444 7146
rect 4402 7118 4444 7126
rect 4472 7146 4513 7148
rect 4472 7126 4486 7146
rect 4505 7126 4513 7146
rect 4785 7137 4824 7181
rect 4472 7118 4513 7126
rect 4402 7112 4513 7118
rect 3730 7091 4174 7094
rect 3730 7089 3898 7091
rect 3459 7043 3463 7048
rect 3420 7040 3463 7043
rect 3353 7026 3463 7040
rect 2082 7006 2250 7007
rect 1467 6998 1508 7006
rect 1467 6978 1475 6998
rect 1494 6978 1508 6998
rect 1467 6976 1508 6978
rect 1536 6998 1578 7006
rect 2131 7005 2239 7006
rect 1536 6978 1552 6998
rect 1571 6978 1578 6998
rect 1536 6976 1578 6978
rect 915 6972 951 6973
rect 763 6942 772 6962
rect 792 6942 800 6962
rect 651 6933 707 6935
rect 651 6932 688 6933
rect 763 6932 800 6942
rect 859 6962 1007 6972
rect 1107 6969 1203 6971
rect 859 6942 868 6962
rect 888 6942 978 6962
rect 998 6942 1007 6962
rect 859 6933 1007 6942
rect 1065 6962 1203 6969
rect 1065 6942 1074 6962
rect 1094 6942 1203 6962
rect 1467 6961 1578 6976
rect 2169 7004 2239 7005
rect 1065 6933 1203 6942
rect 859 6932 896 6933
rect 915 6881 951 6933
rect 970 6932 1007 6933
rect 1066 6932 1103 6933
rect 386 6879 427 6880
rect 278 6872 427 6879
rect 278 6852 396 6872
rect 416 6852 427 6872
rect 278 6844 427 6852
rect 494 6876 853 6880
rect 494 6871 816 6876
rect 494 6847 607 6871
rect 631 6852 816 6871
rect 840 6852 853 6876
rect 631 6847 853 6852
rect 494 6844 853 6847
rect 915 6844 950 6881
rect 1018 6878 1118 6881
rect 1018 6874 1085 6878
rect 1018 6848 1030 6874
rect 1056 6852 1085 6874
rect 1111 6852 1118 6878
rect 1056 6848 1118 6852
rect 1018 6844 1118 6848
rect 494 6823 525 6844
rect 915 6823 951 6844
rect 337 6822 374 6823
rect 111 6819 145 6820
rect 110 6810 147 6819
rect 110 6792 119 6810
rect 137 6792 147 6810
rect 110 6782 147 6792
rect 336 6813 374 6822
rect 336 6793 345 6813
rect 365 6793 374 6813
rect 336 6785 374 6793
rect 440 6817 525 6823
rect 550 6822 587 6823
rect 440 6797 448 6817
rect 468 6797 525 6817
rect 440 6789 525 6797
rect 549 6813 587 6822
rect 549 6793 558 6813
rect 578 6793 587 6813
rect 440 6788 476 6789
rect 549 6785 587 6793
rect 653 6817 738 6823
rect 758 6822 795 6823
rect 653 6797 661 6817
rect 681 6816 738 6817
rect 681 6797 710 6816
rect 653 6796 710 6797
rect 731 6796 738 6816
rect 653 6789 738 6796
rect 757 6813 795 6822
rect 757 6793 766 6813
rect 786 6793 795 6813
rect 653 6788 689 6789
rect 757 6785 795 6793
rect 861 6817 1005 6823
rect 861 6797 869 6817
rect 889 6816 977 6817
rect 889 6797 920 6816
rect 861 6796 920 6797
rect 945 6797 977 6816
rect 997 6797 1005 6817
rect 945 6796 1005 6797
rect 861 6789 1005 6796
rect 861 6788 897 6789
rect 969 6788 1005 6789
rect 1071 6822 1108 6823
rect 1071 6821 1109 6822
rect 1071 6813 1135 6821
rect 1071 6793 1080 6813
rect 1100 6799 1135 6813
rect 1155 6799 1158 6819
rect 1100 6794 1158 6799
rect 1100 6793 1135 6794
rect 111 6754 145 6782
rect 337 6756 374 6785
rect 338 6754 374 6756
rect 550 6754 587 6785
rect 111 6753 283 6754
rect 111 6721 297 6753
rect 338 6732 587 6754
rect 758 6753 795 6785
rect 1071 6781 1135 6793
rect 1175 6755 1202 6933
rect 2169 6897 2230 7004
rect 3730 6911 3757 7089
rect 3797 7051 3861 7063
rect 4137 7059 4174 7091
rect 4345 7090 4594 7112
rect 4345 7059 4382 7090
rect 4558 7088 4594 7090
rect 4558 7059 4595 7088
rect 3797 7050 3832 7051
rect 3774 7045 3832 7050
rect 3774 7025 3777 7045
rect 3797 7031 3832 7045
rect 3852 7031 3861 7051
rect 3797 7023 3861 7031
rect 3823 7022 3861 7023
rect 3824 7021 3861 7022
rect 3927 7055 3963 7056
rect 4035 7055 4071 7056
rect 3927 7050 4071 7055
rect 3927 7047 3989 7050
rect 3927 7027 3935 7047
rect 3955 7030 3989 7047
rect 4012 7047 4071 7050
rect 4012 7030 4043 7047
rect 3955 7027 4043 7030
rect 4063 7027 4071 7047
rect 3927 7021 4071 7027
rect 4137 7051 4175 7059
rect 4243 7055 4279 7056
rect 4137 7031 4146 7051
rect 4166 7031 4175 7051
rect 4137 7022 4175 7031
rect 4194 7048 4279 7055
rect 4194 7028 4201 7048
rect 4222 7047 4279 7048
rect 4222 7028 4251 7047
rect 4194 7027 4251 7028
rect 4271 7027 4279 7047
rect 4137 7021 4174 7022
rect 4194 7021 4279 7027
rect 4345 7051 4383 7059
rect 4456 7055 4492 7056
rect 4345 7031 4354 7051
rect 4374 7031 4383 7051
rect 4345 7022 4383 7031
rect 4407 7047 4492 7055
rect 4407 7027 4464 7047
rect 4484 7027 4492 7047
rect 4345 7021 4382 7022
rect 4407 7021 4492 7027
rect 4558 7051 4596 7059
rect 4558 7031 4567 7051
rect 4587 7031 4596 7051
rect 4558 7022 4596 7031
rect 4558 7021 4595 7022
rect 3981 7000 4017 7021
rect 4407 7000 4438 7021
rect 3814 6996 3914 7000
rect 3814 6992 3876 6996
rect 3814 6966 3821 6992
rect 3847 6970 3876 6992
rect 3902 6970 3914 6996
rect 3847 6966 3914 6970
rect 3814 6963 3914 6966
rect 3982 6963 4017 7000
rect 4079 6997 4438 7000
rect 4079 6992 4301 6997
rect 4079 6968 4092 6992
rect 4116 6973 4301 6992
rect 4325 6973 4438 6997
rect 4116 6968 4438 6973
rect 4079 6964 4438 6968
rect 4505 6992 4654 7000
rect 4505 6972 4516 6992
rect 4536 6972 4654 6992
rect 4505 6965 4654 6972
rect 4505 6964 4546 6965
rect 3829 6911 3866 6912
rect 3925 6911 3962 6912
rect 3981 6911 4017 6963
rect 4036 6911 4073 6912
rect 3729 6902 3867 6911
rect 2169 6886 2239 6897
rect 2169 6877 2176 6886
rect 2171 6857 2176 6877
rect 2224 6857 2239 6886
rect 3729 6882 3838 6902
rect 3858 6882 3867 6902
rect 3729 6875 3867 6882
rect 3925 6902 4073 6911
rect 3925 6882 3934 6902
rect 3954 6882 4044 6902
rect 4064 6882 4073 6902
rect 3729 6873 3825 6875
rect 3925 6872 4073 6882
rect 4132 6902 4169 6912
rect 4244 6911 4281 6912
rect 4225 6909 4281 6911
rect 4132 6882 4140 6902
rect 4160 6882 4169 6902
rect 3981 6871 4017 6872
rect 2171 6848 2239 6857
rect 1358 6829 1468 6843
rect 1358 6826 1401 6829
rect 1358 6821 1362 6826
rect 1034 6753 1202 6755
rect 758 6747 1202 6753
rect 111 6689 145 6721
rect 107 6680 145 6689
rect 107 6662 117 6680
rect 135 6662 145 6680
rect 107 6656 145 6662
rect 263 6658 297 6721
rect 419 6726 530 6732
rect 419 6718 460 6726
rect 419 6698 427 6718
rect 446 6698 460 6718
rect 419 6696 460 6698
rect 488 6718 530 6726
rect 488 6698 504 6718
rect 523 6698 530 6718
rect 488 6696 530 6698
rect 419 6681 530 6696
rect 757 6727 1202 6747
rect 757 6658 795 6727
rect 1034 6726 1202 6727
rect 1280 6799 1362 6821
rect 1391 6799 1401 6826
rect 1429 6802 1436 6829
rect 1465 6821 1468 6829
rect 3463 6838 3574 6853
rect 3463 6836 3505 6838
rect 1465 6802 1530 6821
rect 1429 6799 1530 6802
rect 1280 6797 1530 6799
rect 1280 6718 1317 6797
rect 1358 6784 1468 6797
rect 1432 6728 1463 6729
rect 1280 6698 1289 6718
rect 1309 6698 1317 6718
rect 1280 6688 1317 6698
rect 1376 6718 1463 6728
rect 1376 6698 1385 6718
rect 1405 6698 1463 6718
rect 1376 6689 1463 6698
rect 1376 6688 1413 6689
rect 107 6652 144 6656
rect 263 6647 795 6658
rect 262 6631 795 6647
rect 1432 6636 1463 6689
rect 1493 6718 1530 6797
rect 1701 6794 2094 6814
rect 2114 6794 2117 6814
rect 3196 6809 3237 6818
rect 1701 6789 2117 6794
rect 2791 6807 2959 6808
rect 3196 6807 3205 6809
rect 1701 6788 2042 6789
rect 1645 6728 1676 6729
rect 1493 6698 1502 6718
rect 1522 6698 1530 6718
rect 1493 6688 1530 6698
rect 1589 6721 1676 6728
rect 1589 6718 1650 6721
rect 1589 6698 1598 6718
rect 1618 6701 1650 6718
rect 1671 6701 1676 6721
rect 1618 6698 1676 6701
rect 1589 6691 1676 6698
rect 1701 6718 1738 6788
rect 2004 6787 2041 6788
rect 2791 6787 3205 6807
rect 3231 6787 3237 6809
rect 3463 6816 3470 6836
rect 3489 6816 3505 6836
rect 3463 6808 3505 6816
rect 3533 6836 3574 6838
rect 3533 6816 3547 6836
rect 3566 6816 3574 6836
rect 3533 6808 3574 6816
rect 3829 6812 3866 6813
rect 4132 6812 4169 6882
rect 4194 6902 4281 6909
rect 4194 6899 4252 6902
rect 4194 6879 4199 6899
rect 4220 6882 4252 6899
rect 4272 6882 4281 6902
rect 4220 6879 4281 6882
rect 4194 6872 4281 6879
rect 4340 6902 4377 6912
rect 4340 6882 4348 6902
rect 4368 6882 4377 6902
rect 4194 6871 4225 6872
rect 3828 6811 4169 6812
rect 3463 6802 3574 6808
rect 3753 6806 4169 6811
rect 2791 6781 3237 6787
rect 2791 6779 2959 6781
rect 1853 6728 1889 6729
rect 1701 6698 1710 6718
rect 1730 6698 1738 6718
rect 1589 6689 1645 6691
rect 1589 6688 1626 6689
rect 1701 6688 1738 6698
rect 1797 6718 1945 6728
rect 2045 6725 2141 6727
rect 1797 6698 1806 6718
rect 1826 6698 1916 6718
rect 1936 6698 1945 6718
rect 1797 6689 1945 6698
rect 2003 6718 2141 6725
rect 2003 6698 2012 6718
rect 2032 6698 2141 6718
rect 2003 6689 2141 6698
rect 1797 6688 1834 6689
rect 1853 6637 1889 6689
rect 1908 6688 1945 6689
rect 2004 6688 2041 6689
rect 1324 6635 1365 6636
rect 262 6630 776 6631
rect 1216 6628 1365 6635
rect 1216 6608 1334 6628
rect 1354 6608 1365 6628
rect 1216 6600 1365 6608
rect 1432 6632 1791 6636
rect 1432 6627 1754 6632
rect 1432 6603 1545 6627
rect 1569 6608 1754 6627
rect 1778 6608 1791 6632
rect 1569 6603 1791 6608
rect 1432 6600 1791 6603
rect 1853 6600 1888 6637
rect 1956 6634 2056 6637
rect 1956 6630 2023 6634
rect 1956 6604 1968 6630
rect 1994 6608 2023 6630
rect 2049 6608 2056 6634
rect 1994 6604 2056 6608
rect 1956 6600 2056 6604
rect 110 6589 147 6590
rect 108 6581 148 6589
rect 108 6563 119 6581
rect 137 6563 148 6581
rect 1432 6579 1463 6600
rect 1853 6579 1889 6600
rect 1275 6578 1312 6579
rect 108 6515 148 6563
rect 1274 6569 1312 6578
rect 1274 6549 1283 6569
rect 1303 6549 1312 6569
rect 1274 6541 1312 6549
rect 1378 6573 1463 6579
rect 1488 6578 1525 6579
rect 1378 6553 1386 6573
rect 1406 6553 1463 6573
rect 1378 6545 1463 6553
rect 1487 6569 1525 6578
rect 1487 6549 1496 6569
rect 1516 6549 1525 6569
rect 1378 6544 1414 6545
rect 1487 6541 1525 6549
rect 1591 6573 1676 6579
rect 1696 6578 1733 6579
rect 1591 6553 1599 6573
rect 1619 6572 1676 6573
rect 1619 6553 1648 6572
rect 1591 6552 1648 6553
rect 1669 6552 1676 6572
rect 1591 6545 1676 6552
rect 1695 6569 1733 6578
rect 1695 6549 1704 6569
rect 1724 6549 1733 6569
rect 1591 6544 1627 6545
rect 1695 6541 1733 6549
rect 1799 6573 1943 6579
rect 1799 6553 1807 6573
rect 1827 6556 1863 6573
rect 1883 6556 1915 6573
rect 1827 6553 1915 6556
rect 1935 6553 1943 6573
rect 1799 6545 1943 6553
rect 1799 6544 1835 6545
rect 1907 6544 1943 6545
rect 2009 6578 2046 6579
rect 2009 6577 2047 6578
rect 2009 6569 2073 6577
rect 2009 6549 2018 6569
rect 2038 6555 2073 6569
rect 2093 6555 2096 6575
rect 2038 6550 2096 6555
rect 2038 6549 2073 6550
rect 419 6519 529 6533
rect 419 6516 462 6519
rect 108 6508 233 6515
rect 419 6511 423 6516
rect 108 6489 200 6508
rect 225 6489 233 6508
rect 108 6479 233 6489
rect 341 6489 423 6511
rect 452 6489 462 6516
rect 490 6492 497 6519
rect 526 6511 529 6519
rect 1275 6512 1312 6541
rect 526 6492 591 6511
rect 1276 6510 1312 6512
rect 1488 6510 1525 6541
rect 1696 6514 1733 6541
rect 2009 6537 2073 6549
rect 490 6489 591 6492
rect 341 6487 591 6489
rect 108 6459 148 6479
rect 107 6450 148 6459
rect 107 6432 117 6450
rect 135 6432 148 6450
rect 107 6423 148 6432
rect 107 6422 144 6423
rect 341 6408 378 6487
rect 419 6474 529 6487
rect 493 6418 524 6419
rect 341 6388 350 6408
rect 370 6388 378 6408
rect 341 6378 378 6388
rect 437 6408 524 6418
rect 437 6388 446 6408
rect 466 6388 524 6408
rect 437 6379 524 6388
rect 437 6378 474 6379
rect 110 6356 147 6360
rect 107 6351 147 6356
rect 107 6333 119 6351
rect 137 6333 147 6351
rect 107 6153 147 6333
rect 493 6326 524 6379
rect 554 6408 591 6487
rect 762 6484 1155 6504
rect 1175 6484 1178 6504
rect 1276 6488 1525 6510
rect 1694 6509 1735 6514
rect 2113 6511 2140 6689
rect 2791 6601 2818 6779
rect 3196 6776 3237 6781
rect 3406 6780 3655 6802
rect 3753 6786 3756 6806
rect 3776 6786 4169 6806
rect 4340 6803 4377 6882
rect 4407 6911 4438 6964
rect 4784 6957 4824 7137
rect 5162 7139 5201 7196
rect 5811 7194 5849 7196
rect 6382 7193 6531 7200
rect 6382 7173 6500 7193
rect 6520 7173 6531 7193
rect 6382 7165 6531 7173
rect 6598 7197 6957 7201
rect 6598 7192 6920 7197
rect 6598 7168 6711 7192
rect 6735 7173 6920 7192
rect 6944 7173 6957 7197
rect 6735 7168 6957 7173
rect 6598 7165 6957 7168
rect 7019 7165 7054 7202
rect 7122 7199 7222 7202
rect 7122 7195 7189 7199
rect 7122 7169 7134 7195
rect 7160 7173 7189 7195
rect 7215 7173 7222 7199
rect 7160 7169 7222 7173
rect 7122 7165 7222 7169
rect 6598 7144 6629 7165
rect 7019 7144 7055 7165
rect 6441 7143 6478 7144
rect 5162 7137 5210 7139
rect 5162 7119 5173 7137
rect 5191 7119 5210 7137
rect 6440 7134 6478 7143
rect 5162 7110 5210 7119
rect 5163 7109 5210 7110
rect 5476 7114 5586 7128
rect 5476 7111 5519 7114
rect 5476 7106 5480 7111
rect 5398 7084 5480 7106
rect 5509 7084 5519 7111
rect 5547 7087 5554 7114
rect 5583 7106 5586 7114
rect 6440 7114 6449 7134
rect 6469 7114 6478 7134
rect 6440 7106 6478 7114
rect 6544 7138 6629 7144
rect 6654 7143 6691 7144
rect 6544 7118 6552 7138
rect 6572 7118 6629 7138
rect 6544 7110 6629 7118
rect 6653 7134 6691 7143
rect 6653 7114 6662 7134
rect 6682 7114 6691 7134
rect 6544 7109 6580 7110
rect 6653 7106 6691 7114
rect 6757 7138 6842 7144
rect 6862 7143 6899 7144
rect 6757 7118 6765 7138
rect 6785 7137 6842 7138
rect 6785 7118 6814 7137
rect 6757 7117 6814 7118
rect 6835 7117 6842 7137
rect 6757 7110 6842 7117
rect 6861 7134 6899 7143
rect 6861 7114 6870 7134
rect 6890 7114 6899 7134
rect 6757 7109 6793 7110
rect 6861 7106 6899 7114
rect 6965 7138 7109 7144
rect 6965 7118 6973 7138
rect 6993 7136 7081 7138
rect 6993 7118 7022 7136
rect 6965 7117 7022 7118
rect 7051 7118 7081 7136
rect 7101 7118 7109 7138
rect 7051 7117 7109 7118
rect 6965 7110 7109 7117
rect 6965 7109 7001 7110
rect 7073 7109 7109 7110
rect 7175 7143 7212 7144
rect 7175 7142 7213 7143
rect 7175 7134 7239 7142
rect 7175 7114 7184 7134
rect 7204 7120 7239 7134
rect 7259 7120 7262 7140
rect 7204 7115 7262 7120
rect 7204 7114 7239 7115
rect 5583 7087 5648 7106
rect 5547 7084 5648 7087
rect 5398 7082 5648 7084
rect 5166 7046 5203 7047
rect 4784 6939 4794 6957
rect 4812 6939 4824 6957
rect 4784 6934 4824 6939
rect 5162 7043 5203 7046
rect 5162 7038 5204 7043
rect 5162 7020 5175 7038
rect 5193 7020 5204 7038
rect 5162 7006 5204 7020
rect 5242 7006 5289 7010
rect 5162 7000 5289 7006
rect 5162 6971 5250 7000
rect 5279 6971 5289 7000
rect 5398 7003 5435 7082
rect 5476 7069 5586 7082
rect 5550 7013 5581 7014
rect 5398 6983 5407 7003
rect 5427 6983 5435 7003
rect 5398 6973 5435 6983
rect 5494 7003 5581 7013
rect 5494 6983 5503 7003
rect 5523 6983 5581 7003
rect 5494 6974 5581 6983
rect 5494 6973 5531 6974
rect 5162 6967 5289 6971
rect 5162 6950 5201 6967
rect 5242 6966 5289 6967
rect 4784 6930 4821 6934
rect 5162 6932 5173 6950
rect 5191 6932 5201 6950
rect 5162 6923 5201 6932
rect 5163 6922 5200 6923
rect 5550 6921 5581 6974
rect 5611 7003 5648 7082
rect 5819 7079 6212 7099
rect 6232 7079 6235 7099
rect 5819 7074 6235 7079
rect 6441 7077 6478 7106
rect 6442 7075 6478 7077
rect 6654 7075 6691 7106
rect 5819 7073 6160 7074
rect 5763 7013 5794 7014
rect 5611 6983 5620 7003
rect 5640 6983 5648 7003
rect 5611 6973 5648 6983
rect 5707 7006 5794 7013
rect 5707 7003 5768 7006
rect 5707 6983 5716 7003
rect 5736 6986 5768 7003
rect 5789 6986 5794 7006
rect 5736 6983 5794 6986
rect 5707 6976 5794 6983
rect 5819 7003 5856 7073
rect 6122 7072 6159 7073
rect 6442 7053 6691 7075
rect 6862 7074 6899 7106
rect 7175 7102 7239 7114
rect 7279 7078 7306 7254
rect 7737 7221 7764 7391
rect 7804 7361 7868 7373
rect 8144 7369 8181 7401
rect 8352 7400 8601 7422
rect 8884 7402 8921 7403
rect 9187 7402 9224 7472
rect 9249 7492 9336 7499
rect 9249 7489 9307 7492
rect 9249 7469 9254 7489
rect 9275 7472 9307 7489
rect 9327 7472 9336 7492
rect 9275 7469 9336 7472
rect 9249 7462 9336 7469
rect 9395 7492 9432 7502
rect 9395 7472 9403 7492
rect 9423 7472 9432 7492
rect 9249 7461 9280 7462
rect 8883 7401 9224 7402
rect 8352 7369 8389 7400
rect 8565 7398 8601 7400
rect 8565 7369 8602 7398
rect 8808 7396 9224 7401
rect 8808 7376 8811 7396
rect 8831 7376 9224 7396
rect 9395 7393 9432 7472
rect 9462 7501 9493 7554
rect 9843 7552 9880 7553
rect 9842 7543 9881 7552
rect 9842 7525 9852 7543
rect 9870 7525 9881 7543
rect 10138 7540 10148 7558
rect 10166 7540 10179 7558
rect 10138 7531 10179 7540
rect 10138 7530 10175 7531
rect 9754 7508 9801 7509
rect 9842 7508 9881 7525
rect 9754 7504 9881 7508
rect 9512 7501 9549 7502
rect 9462 7492 9549 7501
rect 9462 7472 9520 7492
rect 9540 7472 9549 7492
rect 9462 7462 9549 7472
rect 9608 7492 9645 7502
rect 9608 7472 9616 7492
rect 9636 7472 9645 7492
rect 9462 7461 9493 7462
rect 9457 7393 9567 7406
rect 9608 7393 9645 7472
rect 9754 7475 9764 7504
rect 9793 7475 9881 7504
rect 10372 7516 10409 7595
rect 10450 7582 10560 7595
rect 10524 7526 10555 7527
rect 10372 7496 10381 7516
rect 10401 7496 10409 7516
rect 10372 7486 10409 7496
rect 10468 7516 10555 7526
rect 10468 7496 10477 7516
rect 10497 7496 10555 7516
rect 10468 7487 10555 7496
rect 10468 7486 10505 7487
rect 9754 7469 9881 7475
rect 9754 7465 9801 7469
rect 9839 7455 9881 7469
rect 10141 7464 10178 7468
rect 9839 7437 9850 7455
rect 9868 7437 9881 7455
rect 9839 7432 9881 7437
rect 9840 7429 9881 7432
rect 10138 7459 10178 7464
rect 10138 7441 10150 7459
rect 10168 7441 10178 7459
rect 9840 7428 9877 7429
rect 9395 7391 9645 7393
rect 9395 7388 9496 7391
rect 9395 7369 9460 7388
rect 7804 7360 7839 7361
rect 7781 7355 7839 7360
rect 7781 7335 7784 7355
rect 7804 7341 7839 7355
rect 7859 7341 7868 7361
rect 7804 7333 7868 7341
rect 7830 7332 7868 7333
rect 7831 7331 7868 7332
rect 7934 7365 7970 7366
rect 8042 7365 8078 7366
rect 7934 7357 8078 7365
rect 7934 7337 7942 7357
rect 7962 7337 8050 7357
rect 8070 7337 8078 7357
rect 7934 7331 8078 7337
rect 8144 7361 8182 7369
rect 8250 7365 8286 7366
rect 8144 7341 8153 7361
rect 8173 7341 8182 7361
rect 8144 7332 8182 7341
rect 8201 7358 8286 7365
rect 8201 7338 8208 7358
rect 8229 7357 8286 7358
rect 8229 7338 8258 7357
rect 8201 7337 8258 7338
rect 8278 7337 8286 7357
rect 8144 7331 8181 7332
rect 8201 7331 8286 7337
rect 8352 7361 8390 7369
rect 8463 7365 8499 7366
rect 8352 7341 8361 7361
rect 8381 7341 8390 7361
rect 8352 7332 8390 7341
rect 8414 7357 8499 7365
rect 8414 7337 8471 7357
rect 8491 7337 8499 7357
rect 8352 7331 8389 7332
rect 8414 7331 8499 7337
rect 8565 7361 8603 7369
rect 8565 7341 8574 7361
rect 8594 7341 8603 7361
rect 9457 7361 9460 7369
rect 9489 7361 9496 7388
rect 9524 7364 9534 7391
rect 9563 7369 9645 7391
rect 9563 7364 9567 7369
rect 9524 7361 9567 7364
rect 9457 7347 9567 7361
rect 9833 7365 9880 7366
rect 9833 7356 9881 7365
rect 8565 7332 8603 7341
rect 9833 7338 9852 7356
rect 9870 7338 9881 7356
rect 9833 7336 9881 7338
rect 8565 7331 8602 7332
rect 7988 7310 8024 7331
rect 8414 7310 8445 7331
rect 7821 7306 7921 7310
rect 7821 7302 7883 7306
rect 7821 7276 7828 7302
rect 7854 7280 7883 7302
rect 7909 7280 7921 7306
rect 7854 7276 7921 7280
rect 7821 7273 7921 7276
rect 7989 7273 8024 7310
rect 8086 7307 8445 7310
rect 8086 7302 8308 7307
rect 8086 7278 8099 7302
rect 8123 7283 8308 7302
rect 8332 7283 8445 7307
rect 8123 7278 8445 7283
rect 8086 7274 8445 7278
rect 8512 7302 8661 7310
rect 8512 7282 8523 7302
rect 8543 7282 8661 7302
rect 8512 7275 8661 7282
rect 9194 7279 9232 7281
rect 9842 7279 9881 7336
rect 8512 7274 8553 7275
rect 7988 7233 8024 7273
rect 7836 7221 7873 7222
rect 7932 7221 7969 7222
rect 7988 7221 7993 7233
rect 7736 7212 7874 7221
rect 7736 7192 7845 7212
rect 7865 7192 7874 7212
rect 7736 7185 7874 7192
rect 7932 7212 7993 7221
rect 7932 7192 7941 7212
rect 7961 7201 7993 7212
rect 8020 7221 8024 7233
rect 8043 7221 8080 7222
rect 8020 7212 8080 7221
rect 8020 7201 8051 7212
rect 7961 7192 8051 7201
rect 8071 7192 8080 7212
rect 7736 7183 7832 7185
rect 7932 7182 8080 7192
rect 8139 7212 8176 7222
rect 8251 7221 8288 7222
rect 8232 7219 8288 7221
rect 8139 7192 8147 7212
rect 8167 7192 8176 7212
rect 7988 7181 8024 7182
rect 7836 7122 7873 7123
rect 8139 7122 8176 7192
rect 8201 7212 8288 7219
rect 8201 7209 8259 7212
rect 8201 7189 8206 7209
rect 8227 7192 8259 7209
rect 8279 7192 8288 7212
rect 8227 7189 8288 7192
rect 8201 7182 8288 7189
rect 8347 7212 8384 7222
rect 8347 7192 8355 7212
rect 8375 7192 8384 7212
rect 8201 7181 8232 7182
rect 7835 7121 8176 7122
rect 7760 7116 8176 7121
rect 7760 7098 7763 7116
rect 7783 7114 8176 7116
rect 7783 7098 8153 7114
rect 7801 7096 8153 7098
rect 8144 7094 8153 7096
rect 8174 7094 8176 7114
rect 8144 7082 8176 7094
rect 8347 7113 8384 7192
rect 8414 7221 8445 7274
rect 9194 7246 9880 7279
rect 8464 7221 8501 7222
rect 8414 7212 8501 7221
rect 8414 7192 8472 7212
rect 8492 7192 8501 7212
rect 8414 7182 8501 7192
rect 8560 7212 8597 7222
rect 8560 7192 8568 7212
rect 8588 7192 8597 7212
rect 8414 7181 8445 7182
rect 8409 7113 8519 7126
rect 8560 7113 8597 7192
rect 8347 7111 8597 7113
rect 8347 7108 8448 7111
rect 8347 7089 8412 7108
rect 7187 7076 7306 7078
rect 7138 7074 7306 7076
rect 6523 7047 6634 7053
rect 6862 7048 7306 7074
rect 8409 7081 8412 7089
rect 8441 7081 8448 7108
rect 8476 7084 8486 7111
rect 8515 7089 8597 7111
rect 8786 7158 8954 7159
rect 9194 7158 9232 7246
rect 9493 7244 9540 7246
rect 9840 7222 9880 7246
rect 8786 7135 9232 7158
rect 9458 7189 9569 7203
rect 9458 7187 9500 7189
rect 9458 7167 9465 7187
rect 9484 7167 9500 7187
rect 9458 7159 9500 7167
rect 9528 7187 9569 7189
rect 9528 7167 9542 7187
rect 9561 7167 9569 7187
rect 9841 7178 9880 7222
rect 9528 7159 9569 7167
rect 9458 7153 9569 7159
rect 8786 7132 9230 7135
rect 8786 7130 8954 7132
rect 8515 7084 8519 7089
rect 8476 7081 8519 7084
rect 8409 7067 8519 7081
rect 7138 7047 7306 7048
rect 6523 7039 6564 7047
rect 6523 7019 6531 7039
rect 6550 7019 6564 7039
rect 6523 7017 6564 7019
rect 6592 7039 6634 7047
rect 7187 7046 7295 7047
rect 6592 7019 6608 7039
rect 6627 7019 6634 7039
rect 6592 7017 6634 7019
rect 5971 7013 6007 7014
rect 5819 6983 5828 7003
rect 5848 6983 5856 7003
rect 5707 6974 5763 6976
rect 5707 6973 5744 6974
rect 5819 6973 5856 6983
rect 5915 7003 6063 7013
rect 6163 7010 6259 7012
rect 5915 6983 5924 7003
rect 5944 6983 6034 7003
rect 6054 6983 6063 7003
rect 5915 6974 6063 6983
rect 6121 7003 6259 7010
rect 6121 6983 6130 7003
rect 6150 6983 6259 7003
rect 6523 7002 6634 7017
rect 7225 7045 7295 7046
rect 6121 6974 6259 6983
rect 5915 6973 5952 6974
rect 5971 6922 6007 6974
rect 6026 6973 6063 6974
rect 6122 6973 6159 6974
rect 5442 6920 5483 6921
rect 5334 6913 5483 6920
rect 4457 6911 4494 6912
rect 4407 6902 4494 6911
rect 4407 6882 4465 6902
rect 4485 6882 4494 6902
rect 4407 6872 4494 6882
rect 4553 6902 4590 6912
rect 4553 6882 4561 6902
rect 4581 6882 4590 6902
rect 5334 6893 5452 6913
rect 5472 6893 5483 6913
rect 5334 6885 5483 6893
rect 5550 6917 5909 6921
rect 5550 6912 5872 6917
rect 5550 6888 5663 6912
rect 5687 6893 5872 6912
rect 5896 6893 5909 6917
rect 5687 6888 5909 6893
rect 5550 6885 5909 6888
rect 5971 6885 6006 6922
rect 6074 6919 6174 6922
rect 6074 6915 6141 6919
rect 6074 6889 6086 6915
rect 6112 6893 6141 6915
rect 6167 6893 6174 6919
rect 6112 6889 6174 6893
rect 6074 6885 6174 6889
rect 4407 6871 4438 6872
rect 4402 6803 4512 6816
rect 4553 6803 4590 6882
rect 4787 6867 4824 6868
rect 4783 6858 4824 6867
rect 5550 6864 5581 6885
rect 5971 6864 6007 6885
rect 5393 6863 5430 6864
rect 5167 6860 5201 6861
rect 4783 6840 4796 6858
rect 4814 6840 4824 6858
rect 4783 6831 4824 6840
rect 5166 6851 5203 6860
rect 5166 6833 5175 6851
rect 5193 6833 5203 6851
rect 4783 6811 4823 6831
rect 5166 6823 5203 6833
rect 5392 6854 5430 6863
rect 5392 6834 5401 6854
rect 5421 6834 5430 6854
rect 5392 6826 5430 6834
rect 5496 6858 5581 6864
rect 5606 6863 5643 6864
rect 5496 6838 5504 6858
rect 5524 6838 5581 6858
rect 5496 6830 5581 6838
rect 5605 6854 5643 6863
rect 5605 6834 5614 6854
rect 5634 6834 5643 6854
rect 5496 6829 5532 6830
rect 5605 6826 5643 6834
rect 5709 6858 5794 6864
rect 5814 6863 5851 6864
rect 5709 6838 5717 6858
rect 5737 6857 5794 6858
rect 5737 6838 5766 6857
rect 5709 6837 5766 6838
rect 5787 6837 5794 6857
rect 5709 6830 5794 6837
rect 5813 6854 5851 6863
rect 5813 6834 5822 6854
rect 5842 6834 5851 6854
rect 5709 6829 5745 6830
rect 5813 6826 5851 6834
rect 5917 6858 6061 6864
rect 5917 6838 5925 6858
rect 5945 6857 6033 6858
rect 5945 6838 5976 6857
rect 5917 6837 5976 6838
rect 6001 6838 6033 6857
rect 6053 6838 6061 6858
rect 6001 6837 6061 6838
rect 5917 6830 6061 6837
rect 5917 6829 5953 6830
rect 6025 6829 6061 6830
rect 6127 6863 6164 6864
rect 6127 6862 6165 6863
rect 6127 6854 6191 6862
rect 6127 6834 6136 6854
rect 6156 6840 6191 6854
rect 6211 6840 6214 6860
rect 6156 6835 6214 6840
rect 6156 6834 6191 6835
rect 4340 6801 4590 6803
rect 4340 6798 4441 6801
rect 2858 6741 2922 6753
rect 3198 6749 3235 6776
rect 3406 6749 3443 6780
rect 3619 6778 3655 6780
rect 4340 6779 4405 6798
rect 3619 6749 3656 6778
rect 4402 6771 4405 6779
rect 4434 6771 4441 6798
rect 4469 6774 4479 6801
rect 4508 6779 4590 6801
rect 4698 6801 4823 6811
rect 4698 6782 4706 6801
rect 4731 6782 4823 6801
rect 4508 6774 4512 6779
rect 4698 6775 4823 6782
rect 4469 6771 4512 6774
rect 4402 6757 4512 6771
rect 2858 6740 2893 6741
rect 2835 6735 2893 6740
rect 2835 6715 2838 6735
rect 2858 6721 2893 6735
rect 2913 6721 2922 6741
rect 2858 6713 2922 6721
rect 2884 6712 2922 6713
rect 2885 6711 2922 6712
rect 2988 6745 3024 6746
rect 3096 6745 3132 6746
rect 2988 6737 3132 6745
rect 2988 6717 2996 6737
rect 3016 6717 3104 6737
rect 3124 6717 3132 6737
rect 2988 6711 3132 6717
rect 3198 6741 3236 6749
rect 3304 6745 3340 6746
rect 3198 6721 3207 6741
rect 3227 6721 3236 6741
rect 3198 6712 3236 6721
rect 3255 6738 3340 6745
rect 3255 6718 3262 6738
rect 3283 6737 3340 6738
rect 3283 6718 3312 6737
rect 3255 6717 3312 6718
rect 3332 6717 3340 6737
rect 3198 6711 3235 6712
rect 3255 6711 3340 6717
rect 3406 6741 3444 6749
rect 3517 6745 3553 6746
rect 3406 6721 3415 6741
rect 3435 6721 3444 6741
rect 3406 6712 3444 6721
rect 3468 6737 3553 6745
rect 3468 6717 3525 6737
rect 3545 6717 3553 6737
rect 3406 6711 3443 6712
rect 3468 6711 3553 6717
rect 3619 6741 3657 6749
rect 3619 6721 3628 6741
rect 3648 6721 3657 6741
rect 3619 6712 3657 6721
rect 4783 6727 4823 6775
rect 5167 6795 5201 6823
rect 5393 6797 5430 6826
rect 5394 6795 5430 6797
rect 5606 6795 5643 6826
rect 5167 6794 5339 6795
rect 5167 6762 5353 6794
rect 5394 6773 5643 6795
rect 5814 6794 5851 6826
rect 6127 6822 6191 6834
rect 6231 6796 6258 6974
rect 7225 6938 7286 7045
rect 8786 6952 8813 7130
rect 8853 7092 8917 7104
rect 9193 7100 9230 7132
rect 9401 7131 9650 7153
rect 9401 7100 9438 7131
rect 9614 7129 9650 7131
rect 9614 7100 9651 7129
rect 8853 7091 8888 7092
rect 8830 7086 8888 7091
rect 8830 7066 8833 7086
rect 8853 7072 8888 7086
rect 8908 7072 8917 7092
rect 8853 7064 8917 7072
rect 8879 7063 8917 7064
rect 8880 7062 8917 7063
rect 8983 7096 9019 7097
rect 9091 7096 9127 7097
rect 8983 7091 9127 7096
rect 8983 7088 9045 7091
rect 8983 7068 8991 7088
rect 9011 7071 9045 7088
rect 9068 7088 9127 7091
rect 9068 7071 9099 7088
rect 9011 7068 9099 7071
rect 9119 7068 9127 7088
rect 8983 7062 9127 7068
rect 9193 7092 9231 7100
rect 9299 7096 9335 7097
rect 9193 7072 9202 7092
rect 9222 7072 9231 7092
rect 9193 7063 9231 7072
rect 9250 7089 9335 7096
rect 9250 7069 9257 7089
rect 9278 7088 9335 7089
rect 9278 7069 9307 7088
rect 9250 7068 9307 7069
rect 9327 7068 9335 7088
rect 9193 7062 9230 7063
rect 9250 7062 9335 7068
rect 9401 7092 9439 7100
rect 9512 7096 9548 7097
rect 9401 7072 9410 7092
rect 9430 7072 9439 7092
rect 9401 7063 9439 7072
rect 9463 7088 9548 7096
rect 9463 7068 9520 7088
rect 9540 7068 9548 7088
rect 9401 7062 9438 7063
rect 9463 7062 9548 7068
rect 9614 7092 9652 7100
rect 9614 7072 9623 7092
rect 9643 7072 9652 7092
rect 9614 7063 9652 7072
rect 9614 7062 9651 7063
rect 9037 7041 9073 7062
rect 9463 7041 9494 7062
rect 8870 7037 8970 7041
rect 8870 7033 8932 7037
rect 8870 7007 8877 7033
rect 8903 7011 8932 7033
rect 8958 7011 8970 7037
rect 8903 7007 8970 7011
rect 8870 7004 8970 7007
rect 9038 7004 9073 7041
rect 9135 7038 9494 7041
rect 9135 7033 9357 7038
rect 9135 7009 9148 7033
rect 9172 7014 9357 7033
rect 9381 7014 9494 7038
rect 9172 7009 9494 7014
rect 9135 7005 9494 7009
rect 9561 7033 9710 7041
rect 9561 7013 9572 7033
rect 9592 7013 9710 7033
rect 9561 7006 9710 7013
rect 9561 7005 9602 7006
rect 8885 6952 8922 6953
rect 8981 6952 9018 6953
rect 9037 6952 9073 7004
rect 9092 6952 9129 6953
rect 8785 6943 8923 6952
rect 7225 6927 7295 6938
rect 7225 6918 7232 6927
rect 7227 6898 7232 6918
rect 7280 6898 7295 6927
rect 8785 6923 8894 6943
rect 8914 6923 8923 6943
rect 8785 6916 8923 6923
rect 8981 6943 9129 6952
rect 8981 6923 8990 6943
rect 9010 6923 9100 6943
rect 9120 6923 9129 6943
rect 8785 6914 8881 6916
rect 8981 6913 9129 6923
rect 9188 6943 9225 6953
rect 9300 6952 9337 6953
rect 9281 6950 9337 6952
rect 9188 6923 9196 6943
rect 9216 6923 9225 6943
rect 9037 6912 9073 6913
rect 7227 6889 7295 6898
rect 6414 6870 6524 6884
rect 6414 6867 6457 6870
rect 6414 6862 6418 6867
rect 6090 6794 6258 6796
rect 5814 6788 6258 6794
rect 5167 6730 5201 6762
rect 3619 6711 3656 6712
rect 3042 6690 3078 6711
rect 3468 6690 3499 6711
rect 4783 6709 4794 6727
rect 4812 6709 4823 6727
rect 4783 6701 4823 6709
rect 5163 6721 5201 6730
rect 5163 6703 5173 6721
rect 5191 6703 5201 6721
rect 4784 6700 4821 6701
rect 5163 6697 5201 6703
rect 5319 6699 5353 6762
rect 5475 6767 5586 6773
rect 5475 6759 5516 6767
rect 5475 6739 5483 6759
rect 5502 6739 5516 6759
rect 5475 6737 5516 6739
rect 5544 6759 5586 6767
rect 5544 6739 5560 6759
rect 5579 6739 5586 6759
rect 5544 6737 5586 6739
rect 5475 6722 5586 6737
rect 5813 6768 6258 6788
rect 5813 6699 5851 6768
rect 6090 6767 6258 6768
rect 6336 6840 6418 6862
rect 6447 6840 6457 6867
rect 6485 6843 6492 6870
rect 6521 6862 6524 6870
rect 8519 6879 8630 6894
rect 8519 6877 8561 6879
rect 6521 6843 6586 6862
rect 6485 6840 6586 6843
rect 6336 6838 6586 6840
rect 6336 6759 6373 6838
rect 6414 6825 6524 6838
rect 6488 6769 6519 6770
rect 6336 6739 6345 6759
rect 6365 6739 6373 6759
rect 6336 6729 6373 6739
rect 6432 6759 6519 6769
rect 6432 6739 6441 6759
rect 6461 6739 6519 6759
rect 6432 6730 6519 6739
rect 6432 6729 6469 6730
rect 5163 6693 5200 6697
rect 2875 6686 2975 6690
rect 2875 6682 2937 6686
rect 2875 6656 2882 6682
rect 2908 6660 2937 6682
rect 2963 6660 2975 6686
rect 2908 6656 2975 6660
rect 2875 6653 2975 6656
rect 3043 6653 3078 6690
rect 3140 6687 3499 6690
rect 3140 6682 3362 6687
rect 3140 6658 3153 6682
rect 3177 6663 3362 6682
rect 3386 6663 3499 6687
rect 3177 6658 3499 6663
rect 3140 6654 3499 6658
rect 3566 6682 3715 6690
rect 5319 6688 5851 6699
rect 3566 6662 3577 6682
rect 3597 6662 3715 6682
rect 5318 6672 5851 6688
rect 6488 6677 6519 6730
rect 6549 6759 6586 6838
rect 6757 6835 7150 6855
rect 7170 6835 7173 6855
rect 8252 6850 8293 6859
rect 6757 6830 7173 6835
rect 7847 6848 8015 6849
rect 8252 6848 8261 6850
rect 6757 6829 7098 6830
rect 6701 6769 6732 6770
rect 6549 6739 6558 6759
rect 6578 6739 6586 6759
rect 6549 6729 6586 6739
rect 6645 6762 6732 6769
rect 6645 6759 6706 6762
rect 6645 6739 6654 6759
rect 6674 6742 6706 6759
rect 6727 6742 6732 6762
rect 6674 6739 6732 6742
rect 6645 6732 6732 6739
rect 6757 6759 6794 6829
rect 7060 6828 7097 6829
rect 7847 6828 8261 6848
rect 8287 6828 8293 6850
rect 8519 6857 8526 6877
rect 8545 6857 8561 6877
rect 8519 6849 8561 6857
rect 8589 6877 8630 6879
rect 8589 6857 8603 6877
rect 8622 6857 8630 6877
rect 8589 6849 8630 6857
rect 8885 6853 8922 6854
rect 9188 6853 9225 6923
rect 9250 6943 9337 6950
rect 9250 6940 9308 6943
rect 9250 6920 9255 6940
rect 9276 6923 9308 6940
rect 9328 6923 9337 6943
rect 9276 6920 9337 6923
rect 9250 6913 9337 6920
rect 9396 6943 9433 6953
rect 9396 6923 9404 6943
rect 9424 6923 9433 6943
rect 9250 6912 9281 6913
rect 8884 6852 9225 6853
rect 8519 6843 8630 6849
rect 8809 6847 9225 6852
rect 7847 6822 8293 6828
rect 7847 6820 8015 6822
rect 6909 6769 6945 6770
rect 6757 6739 6766 6759
rect 6786 6739 6794 6759
rect 6645 6730 6701 6732
rect 6645 6729 6682 6730
rect 6757 6729 6794 6739
rect 6853 6759 7001 6769
rect 7101 6766 7197 6768
rect 6853 6739 6862 6759
rect 6882 6739 6972 6759
rect 6992 6739 7001 6759
rect 6853 6730 7001 6739
rect 7059 6759 7197 6766
rect 7059 6739 7068 6759
rect 7088 6739 7197 6759
rect 7059 6730 7197 6739
rect 6853 6729 6890 6730
rect 6909 6678 6945 6730
rect 6964 6729 7001 6730
rect 7060 6729 7097 6730
rect 6380 6676 6421 6677
rect 5318 6671 5832 6672
rect 3566 6655 3715 6662
rect 6272 6669 6421 6676
rect 4155 6659 4669 6660
rect 3566 6654 3607 6655
rect 3042 6618 3078 6653
rect 2890 6601 2927 6602
rect 2986 6601 3023 6602
rect 3042 6601 3049 6618
rect 2790 6592 2928 6601
rect 2790 6572 2899 6592
rect 2919 6572 2928 6592
rect 2790 6565 2928 6572
rect 2986 6592 3049 6601
rect 2986 6572 2995 6592
rect 3015 6577 3049 6592
rect 3070 6601 3078 6618
rect 3097 6601 3134 6602
rect 3070 6592 3134 6601
rect 3070 6577 3105 6592
rect 3015 6572 3105 6577
rect 3125 6572 3134 6592
rect 2790 6563 2886 6565
rect 2986 6562 3134 6572
rect 3193 6592 3230 6602
rect 3305 6601 3342 6602
rect 3286 6599 3342 6601
rect 3193 6572 3201 6592
rect 3221 6572 3230 6592
rect 3042 6561 3078 6562
rect 1972 6509 2140 6511
rect 1694 6503 2140 6509
rect 762 6479 1178 6484
rect 1357 6482 1468 6488
rect 762 6478 1103 6479
rect 706 6418 737 6419
rect 554 6388 563 6408
rect 583 6388 591 6408
rect 554 6378 591 6388
rect 650 6411 737 6418
rect 650 6408 711 6411
rect 650 6388 659 6408
rect 679 6391 711 6408
rect 732 6391 737 6411
rect 679 6388 737 6391
rect 650 6381 737 6388
rect 762 6408 799 6478
rect 1065 6477 1102 6478
rect 1357 6474 1398 6482
rect 1357 6454 1365 6474
rect 1384 6454 1398 6474
rect 1357 6452 1398 6454
rect 1426 6474 1468 6482
rect 1426 6454 1442 6474
rect 1461 6454 1468 6474
rect 1694 6481 1700 6503
rect 1726 6483 2140 6503
rect 2890 6502 2927 6503
rect 3193 6502 3230 6572
rect 3255 6592 3342 6599
rect 3255 6589 3313 6592
rect 3255 6569 3260 6589
rect 3281 6572 3313 6589
rect 3333 6572 3342 6592
rect 3281 6569 3342 6572
rect 3255 6562 3342 6569
rect 3401 6592 3438 6602
rect 3401 6572 3409 6592
rect 3429 6572 3438 6592
rect 3255 6561 3286 6562
rect 2889 6501 3230 6502
rect 1726 6481 1735 6483
rect 1972 6482 2140 6483
rect 2814 6500 3230 6501
rect 2814 6496 3190 6500
rect 1694 6472 1735 6481
rect 2814 6476 2817 6496
rect 2837 6483 3190 6496
rect 3222 6483 3230 6500
rect 2837 6476 3230 6483
rect 3401 6493 3438 6572
rect 3468 6601 3499 6654
rect 4136 6643 4669 6659
rect 6272 6649 6390 6669
rect 6410 6649 6421 6669
rect 4136 6632 4668 6643
rect 6272 6641 6421 6649
rect 6488 6673 6847 6677
rect 6488 6668 6810 6673
rect 6488 6644 6601 6668
rect 6625 6649 6810 6668
rect 6834 6649 6847 6673
rect 6625 6644 6847 6649
rect 6488 6641 6847 6644
rect 6909 6641 6944 6678
rect 7012 6675 7112 6678
rect 7012 6671 7079 6675
rect 7012 6645 7024 6671
rect 7050 6649 7079 6671
rect 7105 6649 7112 6675
rect 7050 6645 7112 6649
rect 7012 6641 7112 6645
rect 4787 6634 4824 6638
rect 3518 6601 3555 6602
rect 3468 6592 3555 6601
rect 3468 6572 3526 6592
rect 3546 6572 3555 6592
rect 3468 6562 3555 6572
rect 3614 6592 3651 6602
rect 3614 6572 3622 6592
rect 3642 6572 3651 6592
rect 3468 6561 3499 6562
rect 3463 6493 3573 6506
rect 3614 6493 3651 6572
rect 3401 6491 3651 6493
rect 3401 6488 3502 6491
rect 3401 6469 3466 6488
rect 1426 6452 1468 6454
rect 1357 6437 1468 6452
rect 3463 6461 3466 6469
rect 3495 6461 3502 6488
rect 3530 6464 3540 6491
rect 3569 6469 3651 6491
rect 3729 6563 3897 6564
rect 4136 6563 4174 6632
rect 3729 6543 4174 6563
rect 4401 6594 4512 6609
rect 4401 6592 4443 6594
rect 4401 6572 4408 6592
rect 4427 6572 4443 6592
rect 4401 6564 4443 6572
rect 4471 6592 4512 6594
rect 4471 6572 4485 6592
rect 4504 6572 4512 6592
rect 4471 6564 4512 6572
rect 4401 6558 4512 6564
rect 4634 6569 4668 6632
rect 4786 6628 4824 6634
rect 5166 6630 5203 6631
rect 4786 6610 4796 6628
rect 4814 6610 4824 6628
rect 4786 6601 4824 6610
rect 5164 6622 5204 6630
rect 5164 6604 5175 6622
rect 5193 6604 5204 6622
rect 6488 6620 6519 6641
rect 6909 6620 6945 6641
rect 6331 6619 6368 6620
rect 4786 6569 4820 6601
rect 3729 6537 4173 6543
rect 3729 6535 3897 6537
rect 3569 6464 3573 6469
rect 3530 6461 3573 6464
rect 3463 6447 3573 6461
rect 914 6418 950 6419
rect 762 6388 771 6408
rect 791 6388 799 6408
rect 650 6379 706 6381
rect 650 6378 687 6379
rect 762 6378 799 6388
rect 858 6408 1006 6418
rect 1106 6415 1202 6417
rect 858 6388 867 6408
rect 887 6388 977 6408
rect 997 6388 1006 6408
rect 858 6379 1006 6388
rect 1064 6408 1202 6415
rect 1064 6388 1073 6408
rect 1093 6388 1202 6408
rect 1064 6379 1202 6388
rect 858 6378 895 6379
rect 914 6327 950 6379
rect 969 6378 1006 6379
rect 1065 6378 1102 6379
rect 385 6325 426 6326
rect 277 6318 426 6325
rect 277 6298 395 6318
rect 415 6298 426 6318
rect 277 6290 426 6298
rect 493 6322 852 6326
rect 493 6317 815 6322
rect 493 6293 606 6317
rect 630 6298 815 6317
rect 839 6298 852 6322
rect 630 6293 852 6298
rect 493 6290 852 6293
rect 914 6290 949 6327
rect 1017 6324 1117 6327
rect 1017 6320 1084 6324
rect 1017 6294 1029 6320
rect 1055 6298 1084 6320
rect 1110 6298 1117 6324
rect 1055 6294 1117 6298
rect 1017 6290 1117 6294
rect 493 6269 524 6290
rect 914 6269 950 6290
rect 336 6268 373 6269
rect 335 6259 373 6268
rect 335 6239 344 6259
rect 364 6239 373 6259
rect 335 6231 373 6239
rect 439 6263 524 6269
rect 549 6268 586 6269
rect 439 6243 447 6263
rect 467 6243 524 6263
rect 439 6235 524 6243
rect 548 6259 586 6268
rect 548 6239 557 6259
rect 577 6239 586 6259
rect 439 6234 475 6235
rect 548 6231 586 6239
rect 652 6263 737 6269
rect 757 6268 794 6269
rect 652 6243 660 6263
rect 680 6262 737 6263
rect 680 6243 709 6262
rect 652 6242 709 6243
rect 730 6242 737 6262
rect 652 6235 737 6242
rect 756 6259 794 6268
rect 756 6239 765 6259
rect 785 6239 794 6259
rect 652 6234 688 6235
rect 756 6231 794 6239
rect 860 6263 1004 6269
rect 860 6243 868 6263
rect 888 6260 976 6263
rect 888 6243 919 6260
rect 860 6240 919 6243
rect 942 6243 976 6260
rect 996 6243 1004 6263
rect 942 6240 1004 6243
rect 860 6235 1004 6240
rect 860 6234 896 6235
rect 968 6234 1004 6235
rect 1070 6268 1107 6269
rect 1070 6267 1108 6268
rect 1070 6259 1134 6267
rect 1070 6239 1079 6259
rect 1099 6245 1134 6259
rect 1154 6245 1157 6265
rect 1099 6240 1157 6245
rect 1099 6239 1134 6240
rect 336 6202 373 6231
rect 337 6200 373 6202
rect 549 6200 586 6231
rect 337 6178 586 6200
rect 757 6199 794 6231
rect 1070 6227 1134 6239
rect 1174 6201 1201 6379
rect 3729 6357 3756 6535
rect 3796 6497 3860 6509
rect 4136 6505 4173 6537
rect 4344 6536 4593 6558
rect 4634 6537 4820 6569
rect 4648 6536 4820 6537
rect 4344 6505 4381 6536
rect 4557 6534 4593 6536
rect 4557 6505 4594 6534
rect 4786 6508 4820 6536
rect 5164 6556 5204 6604
rect 6330 6610 6368 6619
rect 6330 6590 6339 6610
rect 6359 6590 6368 6610
rect 6330 6582 6368 6590
rect 6434 6614 6519 6620
rect 6544 6619 6581 6620
rect 6434 6594 6442 6614
rect 6462 6594 6519 6614
rect 6434 6586 6519 6594
rect 6543 6610 6581 6619
rect 6543 6590 6552 6610
rect 6572 6590 6581 6610
rect 6434 6585 6470 6586
rect 6543 6582 6581 6590
rect 6647 6614 6732 6620
rect 6752 6619 6789 6620
rect 6647 6594 6655 6614
rect 6675 6613 6732 6614
rect 6675 6594 6704 6613
rect 6647 6593 6704 6594
rect 6725 6593 6732 6613
rect 6647 6586 6732 6593
rect 6751 6610 6789 6619
rect 6751 6590 6760 6610
rect 6780 6590 6789 6610
rect 6647 6585 6683 6586
rect 6751 6582 6789 6590
rect 6855 6614 6999 6620
rect 6855 6594 6863 6614
rect 6883 6597 6919 6614
rect 6939 6597 6971 6614
rect 6883 6594 6971 6597
rect 6991 6594 6999 6614
rect 6855 6586 6999 6594
rect 6855 6585 6891 6586
rect 6963 6585 6999 6586
rect 7065 6619 7102 6620
rect 7065 6618 7103 6619
rect 7065 6610 7129 6618
rect 7065 6590 7074 6610
rect 7094 6596 7129 6610
rect 7149 6596 7152 6616
rect 7094 6591 7152 6596
rect 7094 6590 7129 6591
rect 5475 6560 5585 6574
rect 5475 6557 5518 6560
rect 5164 6549 5289 6556
rect 5475 6552 5479 6557
rect 5164 6530 5256 6549
rect 5281 6530 5289 6549
rect 5164 6520 5289 6530
rect 5397 6530 5479 6552
rect 5508 6530 5518 6557
rect 5546 6533 5553 6560
rect 5582 6552 5585 6560
rect 6331 6553 6368 6582
rect 5582 6533 5647 6552
rect 6332 6551 6368 6553
rect 6544 6551 6581 6582
rect 6752 6555 6789 6582
rect 7065 6578 7129 6590
rect 5546 6530 5647 6533
rect 5397 6528 5647 6530
rect 3796 6496 3831 6497
rect 3773 6491 3831 6496
rect 3773 6471 3776 6491
rect 3796 6477 3831 6491
rect 3851 6477 3860 6497
rect 3796 6469 3860 6477
rect 3822 6468 3860 6469
rect 3823 6467 3860 6468
rect 3926 6501 3962 6502
rect 4034 6501 4070 6502
rect 3926 6494 4070 6501
rect 3926 6493 3986 6494
rect 3926 6473 3934 6493
rect 3954 6474 3986 6493
rect 4011 6493 4070 6494
rect 4011 6474 4042 6493
rect 3954 6473 4042 6474
rect 4062 6473 4070 6493
rect 3926 6467 4070 6473
rect 4136 6497 4174 6505
rect 4242 6501 4278 6502
rect 4136 6477 4145 6497
rect 4165 6477 4174 6497
rect 4136 6468 4174 6477
rect 4193 6494 4278 6501
rect 4193 6474 4200 6494
rect 4221 6493 4278 6494
rect 4221 6474 4250 6493
rect 4193 6473 4250 6474
rect 4270 6473 4278 6493
rect 4136 6467 4173 6468
rect 4193 6467 4278 6473
rect 4344 6497 4382 6505
rect 4455 6501 4491 6502
rect 4344 6477 4353 6497
rect 4373 6477 4382 6497
rect 4344 6468 4382 6477
rect 4406 6493 4491 6501
rect 4406 6473 4463 6493
rect 4483 6473 4491 6493
rect 4344 6467 4381 6468
rect 4406 6467 4491 6473
rect 4557 6497 4595 6505
rect 4557 6477 4566 6497
rect 4586 6477 4595 6497
rect 4557 6468 4595 6477
rect 4784 6498 4821 6508
rect 5164 6500 5204 6520
rect 4784 6480 4794 6498
rect 4812 6480 4821 6498
rect 4784 6471 4821 6480
rect 5163 6491 5204 6500
rect 5163 6473 5173 6491
rect 5191 6473 5204 6491
rect 4786 6470 4820 6471
rect 4557 6467 4594 6468
rect 3980 6446 4016 6467
rect 4406 6446 4437 6467
rect 5163 6464 5204 6473
rect 5163 6463 5200 6464
rect 5397 6449 5434 6528
rect 5475 6515 5585 6528
rect 5549 6459 5580 6460
rect 3813 6442 3913 6446
rect 3813 6438 3875 6442
rect 3813 6412 3820 6438
rect 3846 6416 3875 6438
rect 3901 6416 3913 6442
rect 3846 6412 3913 6416
rect 3813 6409 3913 6412
rect 3981 6409 4016 6446
rect 4078 6443 4437 6446
rect 4078 6438 4300 6443
rect 4078 6414 4091 6438
rect 4115 6419 4300 6438
rect 4324 6419 4437 6443
rect 4115 6414 4437 6419
rect 4078 6410 4437 6414
rect 4504 6438 4653 6446
rect 4504 6418 4515 6438
rect 4535 6418 4653 6438
rect 5397 6429 5406 6449
rect 5426 6429 5434 6449
rect 5397 6419 5434 6429
rect 5493 6449 5580 6459
rect 5493 6429 5502 6449
rect 5522 6429 5580 6449
rect 5493 6420 5580 6429
rect 5493 6419 5530 6420
rect 4504 6411 4653 6418
rect 4504 6410 4545 6411
rect 3828 6357 3865 6358
rect 3924 6357 3961 6358
rect 3980 6357 4016 6409
rect 4035 6357 4072 6358
rect 3728 6348 3866 6357
rect 3323 6327 3434 6342
rect 3323 6325 3365 6327
rect 2993 6304 3098 6306
rect 2651 6296 2819 6297
rect 2993 6296 3042 6304
rect 2651 6277 3042 6296
rect 3073 6277 3098 6304
rect 3323 6305 3330 6325
rect 3349 6305 3365 6325
rect 3323 6297 3365 6305
rect 3393 6325 3434 6327
rect 3393 6305 3407 6325
rect 3426 6305 3434 6325
rect 3728 6328 3837 6348
rect 3857 6328 3866 6348
rect 3728 6321 3866 6328
rect 3924 6348 4072 6357
rect 3924 6328 3933 6348
rect 3953 6328 4043 6348
rect 4063 6328 4072 6348
rect 3728 6319 3824 6321
rect 3924 6318 4072 6328
rect 4131 6348 4168 6358
rect 4243 6357 4280 6358
rect 4224 6355 4280 6357
rect 4131 6328 4139 6348
rect 4159 6328 4168 6348
rect 3980 6317 4016 6318
rect 3393 6297 3434 6305
rect 3323 6291 3434 6297
rect 2651 6270 3098 6277
rect 2651 6268 2819 6270
rect 1499 6237 1609 6251
rect 1499 6234 1542 6237
rect 1499 6229 1503 6234
rect 1033 6199 1201 6201
rect 757 6196 1201 6199
rect 418 6172 529 6178
rect 418 6164 459 6172
rect 107 6109 146 6153
rect 418 6144 426 6164
rect 445 6144 459 6164
rect 418 6142 459 6144
rect 487 6164 529 6172
rect 487 6144 503 6164
rect 522 6144 529 6164
rect 487 6142 529 6144
rect 418 6127 529 6142
rect 755 6173 1201 6196
rect 107 6085 147 6109
rect 447 6085 494 6087
rect 755 6085 793 6173
rect 1033 6172 1201 6173
rect 1421 6207 1503 6229
rect 1532 6207 1542 6234
rect 1570 6210 1577 6237
rect 1606 6229 1609 6237
rect 1606 6210 1671 6229
rect 1570 6207 1671 6210
rect 1421 6205 1671 6207
rect 1421 6126 1458 6205
rect 1499 6192 1609 6205
rect 1573 6136 1604 6137
rect 1421 6106 1430 6126
rect 1450 6106 1458 6126
rect 1421 6096 1458 6106
rect 1517 6126 1604 6136
rect 1517 6106 1526 6126
rect 1546 6106 1604 6126
rect 1517 6097 1604 6106
rect 1517 6096 1554 6097
rect 107 6052 793 6085
rect 107 5995 146 6052
rect 755 6050 793 6052
rect 1573 6044 1604 6097
rect 1634 6126 1671 6205
rect 1842 6218 2235 6222
rect 1842 6201 1861 6218
rect 1881 6202 2235 6218
rect 2255 6202 2258 6222
rect 1881 6201 2258 6202
rect 1842 6197 2258 6201
rect 1842 6196 2183 6197
rect 1786 6136 1817 6137
rect 1634 6106 1643 6126
rect 1663 6106 1671 6126
rect 1634 6096 1671 6106
rect 1730 6129 1817 6136
rect 1730 6126 1791 6129
rect 1730 6106 1739 6126
rect 1759 6109 1791 6126
rect 1812 6109 1817 6129
rect 1759 6106 1817 6109
rect 1730 6099 1817 6106
rect 1842 6126 1879 6196
rect 2145 6195 2182 6196
rect 1994 6136 2030 6137
rect 1842 6106 1851 6126
rect 1871 6106 1879 6126
rect 1730 6097 1786 6099
rect 1730 6096 1767 6097
rect 1842 6096 1879 6106
rect 1938 6126 2086 6136
rect 2254 6135 2283 6136
rect 2186 6133 2283 6135
rect 1938 6106 1947 6126
rect 1967 6122 2057 6126
rect 1967 6106 2000 6122
rect 1938 6097 2000 6106
rect 1938 6096 1975 6097
rect 1994 6084 2000 6097
rect 2023 6106 2057 6122
rect 2077 6106 2086 6126
rect 2023 6097 2086 6106
rect 2144 6126 2283 6133
rect 2144 6106 2153 6126
rect 2173 6106 2283 6126
rect 2144 6097 2283 6106
rect 2023 6084 2030 6097
rect 2049 6096 2086 6097
rect 2145 6096 2182 6097
rect 1994 6045 2030 6084
rect 1465 6043 1506 6044
rect 1357 6036 1506 6043
rect 1357 6016 1475 6036
rect 1495 6016 1506 6036
rect 1357 6008 1506 6016
rect 1573 6040 1932 6044
rect 1573 6035 1895 6040
rect 1573 6011 1686 6035
rect 1710 6016 1895 6035
rect 1919 6016 1932 6040
rect 1710 6011 1932 6016
rect 1573 6008 1932 6011
rect 1994 6008 2029 6045
rect 2097 6042 2197 6045
rect 2097 6038 2164 6042
rect 2097 6012 2109 6038
rect 2135 6016 2164 6038
rect 2190 6016 2197 6042
rect 2135 6012 2197 6016
rect 2097 6008 2197 6012
rect 107 5993 155 5995
rect 107 5975 118 5993
rect 136 5975 155 5993
rect 1573 5987 1604 6008
rect 1994 5987 2030 6008
rect 1416 5986 1453 5987
rect 107 5966 155 5975
rect 108 5965 155 5966
rect 421 5970 531 5984
rect 421 5967 464 5970
rect 421 5962 425 5967
rect 343 5940 425 5962
rect 454 5940 464 5967
rect 492 5943 499 5970
rect 528 5962 531 5970
rect 1415 5977 1453 5986
rect 528 5943 593 5962
rect 1415 5957 1424 5977
rect 1444 5957 1453 5977
rect 492 5940 593 5943
rect 343 5938 593 5940
rect 111 5902 148 5903
rect 107 5899 148 5902
rect 107 5894 149 5899
rect 107 5876 120 5894
rect 138 5876 149 5894
rect 107 5862 149 5876
rect 187 5862 234 5866
rect 107 5856 234 5862
rect 107 5827 195 5856
rect 224 5827 234 5856
rect 343 5859 380 5938
rect 421 5925 531 5938
rect 495 5869 526 5870
rect 343 5839 352 5859
rect 372 5839 380 5859
rect 343 5829 380 5839
rect 439 5859 526 5869
rect 439 5839 448 5859
rect 468 5839 526 5859
rect 439 5830 526 5839
rect 439 5829 476 5830
rect 107 5823 234 5827
rect 107 5806 146 5823
rect 187 5822 234 5823
rect 107 5788 118 5806
rect 136 5788 146 5806
rect 107 5779 146 5788
rect 108 5778 145 5779
rect 495 5777 526 5830
rect 556 5859 593 5938
rect 764 5935 1157 5955
rect 1177 5935 1180 5955
rect 1415 5949 1453 5957
rect 1519 5981 1604 5987
rect 1629 5986 1666 5987
rect 1519 5961 1527 5981
rect 1547 5961 1604 5981
rect 1519 5953 1604 5961
rect 1628 5977 1666 5986
rect 1628 5957 1637 5977
rect 1657 5957 1666 5977
rect 1519 5952 1555 5953
rect 1628 5949 1666 5957
rect 1732 5981 1817 5987
rect 1837 5986 1874 5987
rect 1732 5961 1740 5981
rect 1760 5980 1817 5981
rect 1760 5961 1789 5980
rect 1732 5960 1789 5961
rect 1810 5960 1817 5980
rect 1732 5953 1817 5960
rect 1836 5977 1874 5986
rect 1836 5957 1845 5977
rect 1865 5957 1874 5977
rect 1732 5952 1768 5953
rect 1836 5949 1874 5957
rect 1940 5981 2084 5987
rect 1940 5961 1948 5981
rect 1968 5961 2056 5981
rect 2076 5961 2084 5981
rect 1940 5953 2084 5961
rect 1940 5952 1976 5953
rect 2048 5952 2084 5953
rect 2150 5986 2187 5987
rect 2150 5985 2188 5986
rect 2150 5977 2214 5985
rect 2150 5957 2159 5977
rect 2179 5963 2214 5977
rect 2234 5963 2237 5983
rect 2179 5958 2237 5963
rect 2179 5957 2214 5958
rect 764 5930 1180 5935
rect 764 5929 1105 5930
rect 708 5869 739 5870
rect 556 5839 565 5859
rect 585 5839 593 5859
rect 556 5829 593 5839
rect 652 5862 739 5869
rect 652 5859 713 5862
rect 652 5839 661 5859
rect 681 5842 713 5859
rect 734 5842 739 5862
rect 681 5839 739 5842
rect 652 5832 739 5839
rect 764 5859 801 5929
rect 1067 5928 1104 5929
rect 1416 5920 1453 5949
rect 1417 5918 1453 5920
rect 1629 5918 1666 5949
rect 1417 5896 1666 5918
rect 1837 5917 1874 5949
rect 2150 5945 2214 5957
rect 2254 5919 2283 6097
rect 2651 6090 2678 6268
rect 2718 6230 2782 6242
rect 3058 6238 3095 6270
rect 3266 6269 3515 6291
rect 3266 6238 3303 6269
rect 3479 6267 3515 6269
rect 3479 6238 3516 6267
rect 3828 6258 3865 6259
rect 4131 6258 4168 6328
rect 4193 6348 4280 6355
rect 4193 6345 4251 6348
rect 4193 6325 4198 6345
rect 4219 6328 4251 6345
rect 4271 6328 4280 6348
rect 4219 6325 4280 6328
rect 4193 6318 4280 6325
rect 4339 6348 4376 6358
rect 4339 6328 4347 6348
rect 4367 6328 4376 6348
rect 4193 6317 4224 6318
rect 3827 6257 4168 6258
rect 3752 6252 4168 6257
rect 2718 6229 2753 6230
rect 2695 6224 2753 6229
rect 2695 6204 2698 6224
rect 2718 6210 2753 6224
rect 2773 6210 2782 6230
rect 2718 6202 2782 6210
rect 2744 6201 2782 6202
rect 2745 6200 2782 6201
rect 2848 6234 2884 6235
rect 2956 6234 2992 6235
rect 2848 6229 2992 6234
rect 2848 6226 2908 6229
rect 2848 6206 2856 6226
rect 2876 6208 2908 6226
rect 2935 6226 2992 6229
rect 2935 6208 2964 6226
rect 2876 6206 2964 6208
rect 2984 6206 2992 6226
rect 2848 6200 2992 6206
rect 3058 6230 3096 6238
rect 3164 6234 3200 6235
rect 3058 6210 3067 6230
rect 3087 6210 3096 6230
rect 3058 6201 3096 6210
rect 3115 6227 3200 6234
rect 3115 6207 3122 6227
rect 3143 6226 3200 6227
rect 3143 6207 3172 6226
rect 3115 6206 3172 6207
rect 3192 6206 3200 6226
rect 3058 6200 3095 6201
rect 3115 6200 3200 6206
rect 3266 6230 3304 6238
rect 3377 6234 3413 6235
rect 3266 6210 3275 6230
rect 3295 6210 3304 6230
rect 3266 6201 3304 6210
rect 3328 6226 3413 6234
rect 3328 6206 3385 6226
rect 3405 6206 3413 6226
rect 3266 6200 3303 6201
rect 3328 6200 3413 6206
rect 3479 6230 3517 6238
rect 3752 6232 3755 6252
rect 3775 6232 4168 6252
rect 4339 6249 4376 6328
rect 4406 6357 4437 6410
rect 4787 6408 4824 6409
rect 4786 6399 4825 6408
rect 4786 6381 4796 6399
rect 4814 6381 4825 6399
rect 5166 6397 5203 6401
rect 4698 6364 4745 6365
rect 4786 6364 4825 6381
rect 4698 6360 4825 6364
rect 4456 6357 4493 6358
rect 4406 6348 4493 6357
rect 4406 6328 4464 6348
rect 4484 6328 4493 6348
rect 4406 6318 4493 6328
rect 4552 6348 4589 6358
rect 4552 6328 4560 6348
rect 4580 6328 4589 6348
rect 4406 6317 4437 6318
rect 4401 6249 4511 6262
rect 4552 6249 4589 6328
rect 4698 6331 4708 6360
rect 4737 6331 4825 6360
rect 4698 6325 4825 6331
rect 4698 6321 4745 6325
rect 4783 6311 4825 6325
rect 4783 6293 4794 6311
rect 4812 6293 4825 6311
rect 4783 6288 4825 6293
rect 4784 6285 4825 6288
rect 5163 6392 5203 6397
rect 5163 6374 5175 6392
rect 5193 6374 5203 6392
rect 4784 6284 4821 6285
rect 4339 6247 4589 6249
rect 4339 6244 4440 6247
rect 3479 6210 3488 6230
rect 3508 6210 3517 6230
rect 4339 6225 4404 6244
rect 3479 6201 3517 6210
rect 4401 6217 4404 6225
rect 4433 6217 4440 6244
rect 4468 6220 4478 6247
rect 4507 6225 4589 6247
rect 4507 6220 4511 6225
rect 4468 6217 4511 6220
rect 4401 6203 4511 6217
rect 4777 6221 4824 6222
rect 4777 6212 4825 6221
rect 3479 6200 3516 6201
rect 2902 6179 2938 6200
rect 3328 6179 3359 6200
rect 4777 6194 4796 6212
rect 4814 6194 4825 6212
rect 4777 6192 4825 6194
rect 2735 6175 2835 6179
rect 2735 6171 2797 6175
rect 2735 6145 2742 6171
rect 2768 6149 2797 6171
rect 2823 6149 2835 6175
rect 2768 6145 2835 6149
rect 2735 6142 2835 6145
rect 2903 6142 2938 6179
rect 3000 6176 3359 6179
rect 3000 6171 3222 6176
rect 3000 6147 3013 6171
rect 3037 6152 3222 6171
rect 3246 6152 3359 6176
rect 3037 6147 3359 6152
rect 3000 6143 3359 6147
rect 3426 6171 3575 6179
rect 3426 6151 3437 6171
rect 3457 6151 3575 6171
rect 3426 6144 3575 6151
rect 3426 6143 3467 6144
rect 2750 6090 2787 6091
rect 2846 6090 2883 6091
rect 2902 6090 2938 6142
rect 2957 6090 2994 6091
rect 2650 6081 2788 6090
rect 2650 6061 2759 6081
rect 2779 6061 2788 6081
rect 2650 6054 2788 6061
rect 2846 6081 2994 6090
rect 2846 6061 2855 6081
rect 2875 6061 2965 6081
rect 2985 6061 2994 6081
rect 2650 6052 2746 6054
rect 2846 6051 2994 6061
rect 3053 6081 3090 6091
rect 3165 6090 3202 6091
rect 3146 6088 3202 6090
rect 3053 6061 3061 6081
rect 3081 6061 3090 6081
rect 2902 6050 2938 6051
rect 2750 5991 2787 5992
rect 3053 5991 3090 6061
rect 3115 6081 3202 6088
rect 3115 6078 3173 6081
rect 3115 6058 3120 6078
rect 3141 6061 3173 6078
rect 3193 6061 3202 6081
rect 3141 6058 3202 6061
rect 3115 6051 3202 6058
rect 3261 6081 3298 6091
rect 3261 6061 3269 6081
rect 3289 6061 3298 6081
rect 3115 6050 3146 6051
rect 2749 5990 3090 5991
rect 2674 5986 3090 5990
rect 2674 5985 3051 5986
rect 2674 5965 2677 5985
rect 2697 5969 3051 5985
rect 3071 5969 3090 5986
rect 2697 5965 3090 5969
rect 3261 5982 3298 6061
rect 3328 6090 3359 6143
rect 4139 6135 4177 6137
rect 4786 6135 4825 6192
rect 4139 6102 4825 6135
rect 3378 6090 3415 6091
rect 3328 6081 3415 6090
rect 3328 6061 3386 6081
rect 3406 6061 3415 6081
rect 3328 6051 3415 6061
rect 3474 6081 3511 6091
rect 3474 6061 3482 6081
rect 3502 6061 3511 6081
rect 3328 6050 3359 6051
rect 3323 5982 3433 5995
rect 3474 5982 3511 6061
rect 3261 5980 3511 5982
rect 3261 5977 3362 5980
rect 3261 5958 3326 5977
rect 3323 5950 3326 5958
rect 3355 5950 3362 5977
rect 3390 5953 3400 5980
rect 3429 5958 3511 5980
rect 3731 6014 3899 6015
rect 4139 6014 4177 6102
rect 4438 6100 4485 6102
rect 4785 6078 4825 6102
rect 3731 5991 4177 6014
rect 4403 6045 4514 6060
rect 4403 6043 4445 6045
rect 4403 6023 4410 6043
rect 4429 6023 4445 6043
rect 4403 6015 4445 6023
rect 4473 6043 4514 6045
rect 4473 6023 4487 6043
rect 4506 6023 4514 6043
rect 4786 6034 4825 6078
rect 4473 6015 4514 6023
rect 4403 6009 4514 6015
rect 3731 5988 4175 5991
rect 3731 5986 3899 5988
rect 3429 5953 3433 5958
rect 3390 5950 3433 5953
rect 3323 5936 3433 5950
rect 2113 5917 2283 5919
rect 1834 5910 2283 5917
rect 1498 5890 1609 5896
rect 1498 5882 1539 5890
rect 916 5869 952 5870
rect 764 5839 773 5859
rect 793 5839 801 5859
rect 652 5830 708 5832
rect 652 5829 689 5830
rect 764 5829 801 5839
rect 860 5859 1008 5869
rect 1108 5866 1204 5868
rect 860 5839 869 5859
rect 889 5839 979 5859
rect 999 5839 1008 5859
rect 860 5830 1008 5839
rect 1066 5859 1204 5866
rect 1066 5839 1075 5859
rect 1095 5839 1204 5859
rect 1498 5862 1506 5882
rect 1525 5862 1539 5882
rect 1498 5860 1539 5862
rect 1567 5882 1609 5890
rect 1567 5862 1583 5882
rect 1602 5862 1609 5882
rect 1834 5883 1859 5910
rect 1890 5891 2283 5910
rect 1890 5883 1939 5891
rect 2113 5890 2283 5891
rect 1834 5881 1939 5883
rect 1567 5860 1609 5862
rect 1498 5845 1609 5860
rect 1066 5830 1204 5839
rect 860 5829 897 5830
rect 916 5778 952 5830
rect 971 5829 1008 5830
rect 1067 5829 1104 5830
rect 387 5776 428 5777
rect 279 5769 428 5776
rect 279 5749 397 5769
rect 417 5749 428 5769
rect 279 5741 428 5749
rect 495 5773 854 5777
rect 495 5768 817 5773
rect 495 5744 608 5768
rect 632 5749 817 5768
rect 841 5749 854 5773
rect 632 5744 854 5749
rect 495 5741 854 5744
rect 916 5741 951 5778
rect 1019 5775 1119 5778
rect 1019 5771 1086 5775
rect 1019 5745 1031 5771
rect 1057 5749 1086 5771
rect 1112 5749 1119 5775
rect 1057 5745 1119 5749
rect 1019 5741 1119 5745
rect 495 5720 526 5741
rect 916 5720 952 5741
rect 338 5719 375 5720
rect 112 5716 146 5717
rect 111 5707 148 5716
rect 111 5689 120 5707
rect 138 5689 148 5707
rect 111 5679 148 5689
rect 337 5710 375 5719
rect 337 5690 346 5710
rect 366 5690 375 5710
rect 337 5682 375 5690
rect 441 5714 526 5720
rect 551 5719 588 5720
rect 441 5694 449 5714
rect 469 5694 526 5714
rect 441 5686 526 5694
rect 550 5710 588 5719
rect 550 5690 559 5710
rect 579 5690 588 5710
rect 441 5685 477 5686
rect 550 5682 588 5690
rect 654 5714 739 5720
rect 759 5719 796 5720
rect 654 5694 662 5714
rect 682 5713 739 5714
rect 682 5694 711 5713
rect 654 5693 711 5694
rect 732 5693 739 5713
rect 654 5686 739 5693
rect 758 5710 796 5719
rect 758 5690 767 5710
rect 787 5690 796 5710
rect 654 5685 690 5686
rect 758 5682 796 5690
rect 862 5714 1006 5720
rect 862 5694 870 5714
rect 890 5713 978 5714
rect 890 5694 921 5713
rect 862 5693 921 5694
rect 946 5694 978 5713
rect 998 5694 1006 5714
rect 946 5693 1006 5694
rect 862 5686 1006 5693
rect 862 5685 898 5686
rect 970 5685 1006 5686
rect 1072 5719 1109 5720
rect 1072 5718 1110 5719
rect 1072 5710 1136 5718
rect 1072 5690 1081 5710
rect 1101 5696 1136 5710
rect 1156 5696 1159 5716
rect 1101 5691 1159 5696
rect 1101 5690 1136 5691
rect 112 5651 146 5679
rect 338 5653 375 5682
rect 339 5651 375 5653
rect 551 5651 588 5682
rect 112 5650 284 5651
rect 112 5618 298 5650
rect 339 5629 588 5651
rect 759 5650 796 5682
rect 1072 5678 1136 5690
rect 1176 5652 1203 5830
rect 3731 5808 3758 5986
rect 3798 5948 3862 5960
rect 4138 5956 4175 5988
rect 4346 5987 4595 6009
rect 4346 5956 4383 5987
rect 4559 5985 4595 5987
rect 4559 5956 4596 5985
rect 3798 5947 3833 5948
rect 3775 5942 3833 5947
rect 3775 5922 3778 5942
rect 3798 5928 3833 5942
rect 3853 5928 3862 5948
rect 3798 5920 3862 5928
rect 3824 5919 3862 5920
rect 3825 5918 3862 5919
rect 3928 5952 3964 5953
rect 4036 5952 4072 5953
rect 3928 5947 4072 5952
rect 3928 5944 3990 5947
rect 3928 5924 3936 5944
rect 3956 5927 3990 5944
rect 4013 5944 4072 5947
rect 4013 5927 4044 5944
rect 3956 5924 4044 5927
rect 4064 5924 4072 5944
rect 3928 5918 4072 5924
rect 4138 5948 4176 5956
rect 4244 5952 4280 5953
rect 4138 5928 4147 5948
rect 4167 5928 4176 5948
rect 4138 5919 4176 5928
rect 4195 5945 4280 5952
rect 4195 5925 4202 5945
rect 4223 5944 4280 5945
rect 4223 5925 4252 5944
rect 4195 5924 4252 5925
rect 4272 5924 4280 5944
rect 4138 5918 4175 5919
rect 4195 5918 4280 5924
rect 4346 5948 4384 5956
rect 4457 5952 4493 5953
rect 4346 5928 4355 5948
rect 4375 5928 4384 5948
rect 4346 5919 4384 5928
rect 4408 5944 4493 5952
rect 4408 5924 4465 5944
rect 4485 5924 4493 5944
rect 4346 5918 4383 5919
rect 4408 5918 4493 5924
rect 4559 5948 4597 5956
rect 4559 5928 4568 5948
rect 4588 5928 4597 5948
rect 4559 5919 4597 5928
rect 4559 5918 4596 5919
rect 3982 5897 4018 5918
rect 4408 5897 4439 5918
rect 3815 5893 3915 5897
rect 3815 5889 3877 5893
rect 3815 5863 3822 5889
rect 3848 5867 3877 5889
rect 3903 5867 3915 5893
rect 3848 5863 3915 5867
rect 3815 5860 3915 5863
rect 3983 5860 4018 5897
rect 4080 5894 4439 5897
rect 4080 5889 4302 5894
rect 4080 5865 4093 5889
rect 4117 5870 4302 5889
rect 4326 5870 4439 5894
rect 4117 5865 4439 5870
rect 4080 5861 4439 5865
rect 4506 5889 4655 5897
rect 4506 5869 4517 5889
rect 4537 5869 4655 5889
rect 4506 5862 4655 5869
rect 4506 5861 4547 5862
rect 3830 5808 3867 5809
rect 3926 5808 3963 5809
rect 3982 5808 4018 5860
rect 4037 5808 4074 5809
rect 3730 5799 3868 5808
rect 3730 5779 3839 5799
rect 3859 5779 3868 5799
rect 3730 5772 3868 5779
rect 3926 5799 4074 5808
rect 3926 5779 3935 5799
rect 3955 5779 4045 5799
rect 4065 5779 4074 5799
rect 3730 5770 3826 5772
rect 3926 5769 4074 5779
rect 4133 5799 4170 5809
rect 4245 5808 4282 5809
rect 4226 5806 4282 5808
rect 4133 5779 4141 5799
rect 4161 5779 4170 5799
rect 3982 5768 4018 5769
rect 1359 5726 1469 5740
rect 1359 5723 1402 5726
rect 1359 5718 1363 5723
rect 1035 5650 1203 5652
rect 759 5644 1203 5650
rect 112 5586 146 5618
rect 108 5577 146 5586
rect 108 5559 118 5577
rect 136 5559 146 5577
rect 108 5553 146 5559
rect 264 5555 298 5618
rect 420 5623 531 5629
rect 420 5615 461 5623
rect 420 5595 428 5615
rect 447 5595 461 5615
rect 420 5593 461 5595
rect 489 5615 531 5623
rect 489 5595 505 5615
rect 524 5595 531 5615
rect 489 5593 531 5595
rect 420 5578 531 5593
rect 758 5624 1203 5644
rect 758 5555 796 5624
rect 1035 5623 1203 5624
rect 1281 5696 1363 5718
rect 1392 5696 1402 5723
rect 1430 5699 1437 5726
rect 1466 5718 1469 5726
rect 3464 5735 3575 5750
rect 3464 5733 3506 5735
rect 1466 5699 1531 5718
rect 1430 5696 1531 5699
rect 1281 5694 1531 5696
rect 1281 5615 1318 5694
rect 1359 5681 1469 5694
rect 1433 5625 1464 5626
rect 1281 5595 1290 5615
rect 1310 5595 1318 5615
rect 1281 5585 1318 5595
rect 1377 5615 1464 5625
rect 1377 5595 1386 5615
rect 1406 5595 1464 5615
rect 1377 5586 1464 5595
rect 1377 5585 1414 5586
rect 108 5549 145 5553
rect 264 5544 796 5555
rect 263 5528 796 5544
rect 1433 5533 1464 5586
rect 1494 5615 1531 5694
rect 1702 5704 2095 5711
rect 1702 5687 1710 5704
rect 1742 5691 2095 5704
rect 2115 5691 2118 5711
rect 3197 5706 3238 5715
rect 1742 5687 2118 5691
rect 1702 5686 2118 5687
rect 2792 5704 2960 5705
rect 3197 5704 3206 5706
rect 1702 5685 2043 5686
rect 1646 5625 1677 5626
rect 1494 5595 1503 5615
rect 1523 5595 1531 5615
rect 1494 5585 1531 5595
rect 1590 5618 1677 5625
rect 1590 5615 1651 5618
rect 1590 5595 1599 5615
rect 1619 5598 1651 5615
rect 1672 5598 1677 5618
rect 1619 5595 1677 5598
rect 1590 5588 1677 5595
rect 1702 5615 1739 5685
rect 2005 5684 2042 5685
rect 2792 5684 3206 5704
rect 3232 5684 3238 5706
rect 3464 5713 3471 5733
rect 3490 5713 3506 5733
rect 3464 5705 3506 5713
rect 3534 5733 3575 5735
rect 3534 5713 3548 5733
rect 3567 5713 3575 5733
rect 3534 5705 3575 5713
rect 3830 5709 3867 5710
rect 4133 5709 4170 5779
rect 4195 5799 4282 5806
rect 4195 5796 4253 5799
rect 4195 5776 4200 5796
rect 4221 5779 4253 5796
rect 4273 5779 4282 5799
rect 4221 5776 4282 5779
rect 4195 5769 4282 5776
rect 4341 5799 4378 5809
rect 4341 5779 4349 5799
rect 4369 5779 4378 5799
rect 4195 5768 4226 5769
rect 3829 5708 4170 5709
rect 3464 5699 3575 5705
rect 3754 5703 4170 5708
rect 2792 5678 3238 5684
rect 2792 5676 2960 5678
rect 1854 5625 1890 5626
rect 1702 5595 1711 5615
rect 1731 5595 1739 5615
rect 1590 5586 1646 5588
rect 1590 5585 1627 5586
rect 1702 5585 1739 5595
rect 1798 5615 1946 5625
rect 2046 5622 2142 5624
rect 1798 5595 1807 5615
rect 1827 5610 1917 5615
rect 1827 5595 1862 5610
rect 1798 5586 1862 5595
rect 1798 5585 1835 5586
rect 1854 5569 1862 5586
rect 1883 5595 1917 5610
rect 1937 5595 1946 5615
rect 1883 5586 1946 5595
rect 2004 5615 2142 5622
rect 2004 5595 2013 5615
rect 2033 5595 2142 5615
rect 2004 5586 2142 5595
rect 1883 5569 1890 5586
rect 1909 5585 1946 5586
rect 2005 5585 2042 5586
rect 1854 5534 1890 5569
rect 1325 5532 1366 5533
rect 263 5527 777 5528
rect 1217 5525 1366 5532
rect 1217 5505 1335 5525
rect 1355 5505 1366 5525
rect 1217 5497 1366 5505
rect 1433 5529 1792 5533
rect 1433 5524 1755 5529
rect 1433 5500 1546 5524
rect 1570 5505 1755 5524
rect 1779 5505 1792 5529
rect 1570 5500 1792 5505
rect 1433 5497 1792 5500
rect 1854 5497 1889 5534
rect 1957 5531 2057 5534
rect 1957 5527 2024 5531
rect 1957 5501 1969 5527
rect 1995 5505 2024 5527
rect 2050 5505 2057 5531
rect 1995 5501 2057 5505
rect 1957 5497 2057 5501
rect 111 5486 148 5487
rect 109 5478 149 5486
rect 109 5460 120 5478
rect 138 5460 149 5478
rect 1433 5476 1464 5497
rect 1854 5476 1890 5497
rect 1276 5475 1313 5476
rect 109 5412 149 5460
rect 1275 5466 1313 5475
rect 1275 5446 1284 5466
rect 1304 5446 1313 5466
rect 1275 5438 1313 5446
rect 1379 5470 1464 5476
rect 1489 5475 1526 5476
rect 1379 5450 1387 5470
rect 1407 5450 1464 5470
rect 1379 5442 1464 5450
rect 1488 5466 1526 5475
rect 1488 5446 1497 5466
rect 1517 5446 1526 5466
rect 1379 5441 1415 5442
rect 1488 5438 1526 5446
rect 1592 5470 1677 5476
rect 1697 5475 1734 5476
rect 1592 5450 1600 5470
rect 1620 5469 1677 5470
rect 1620 5450 1649 5469
rect 1592 5449 1649 5450
rect 1670 5449 1677 5469
rect 1592 5442 1677 5449
rect 1696 5466 1734 5475
rect 1696 5446 1705 5466
rect 1725 5446 1734 5466
rect 1592 5441 1628 5442
rect 1696 5438 1734 5446
rect 1800 5470 1944 5476
rect 1800 5450 1808 5470
rect 1828 5450 1916 5470
rect 1936 5450 1944 5470
rect 1800 5442 1944 5450
rect 1800 5441 1836 5442
rect 1908 5441 1944 5442
rect 2010 5475 2047 5476
rect 2010 5474 2048 5475
rect 2010 5466 2074 5474
rect 2010 5446 2019 5466
rect 2039 5452 2074 5466
rect 2094 5452 2097 5472
rect 2039 5447 2097 5452
rect 2039 5446 2074 5447
rect 420 5416 530 5430
rect 420 5413 463 5416
rect 109 5405 234 5412
rect 420 5408 424 5413
rect 109 5386 201 5405
rect 226 5386 234 5405
rect 109 5376 234 5386
rect 342 5386 424 5408
rect 453 5386 463 5413
rect 491 5389 498 5416
rect 527 5408 530 5416
rect 1276 5409 1313 5438
rect 527 5389 592 5408
rect 1277 5407 1313 5409
rect 1489 5407 1526 5438
rect 1697 5411 1734 5438
rect 2010 5434 2074 5446
rect 491 5386 592 5389
rect 342 5384 592 5386
rect 109 5356 149 5376
rect 108 5347 149 5356
rect 108 5329 118 5347
rect 136 5329 149 5347
rect 108 5320 149 5329
rect 108 5319 145 5320
rect 342 5305 379 5384
rect 420 5371 530 5384
rect 494 5315 525 5316
rect 342 5285 351 5305
rect 371 5285 379 5305
rect 342 5275 379 5285
rect 438 5305 525 5315
rect 438 5285 447 5305
rect 467 5285 525 5305
rect 438 5276 525 5285
rect 438 5275 475 5276
rect 111 5253 148 5257
rect 108 5248 148 5253
rect 108 5230 120 5248
rect 138 5230 148 5248
rect 108 5050 148 5230
rect 494 5223 525 5276
rect 555 5305 592 5384
rect 763 5381 1156 5401
rect 1176 5381 1179 5401
rect 1277 5385 1526 5407
rect 1695 5406 1736 5411
rect 2114 5408 2141 5586
rect 2792 5498 2819 5676
rect 3197 5673 3238 5678
rect 3407 5677 3656 5699
rect 3754 5683 3757 5703
rect 3777 5683 4170 5703
rect 4341 5700 4378 5779
rect 4408 5808 4439 5861
rect 4785 5854 4825 6034
rect 5163 6194 5203 6374
rect 5549 6367 5580 6420
rect 5610 6449 5647 6528
rect 5818 6525 6211 6545
rect 6231 6525 6234 6545
rect 6332 6529 6581 6551
rect 6750 6550 6791 6555
rect 7169 6552 7196 6730
rect 7847 6642 7874 6820
rect 8252 6817 8293 6822
rect 8462 6821 8711 6843
rect 8809 6827 8812 6847
rect 8832 6827 9225 6847
rect 9396 6844 9433 6923
rect 9463 6952 9494 7005
rect 9840 6998 9880 7178
rect 10138 7261 10178 7441
rect 10524 7434 10555 7487
rect 10585 7516 10622 7595
rect 10793 7592 11186 7612
rect 11206 7592 11209 7612
rect 11307 7596 11556 7618
rect 11725 7617 11766 7622
rect 12144 7619 12171 7797
rect 12822 7709 12849 7887
rect 13227 7884 13268 7889
rect 13437 7888 13686 7910
rect 13784 7894 13787 7914
rect 13807 7894 14200 7914
rect 14371 7911 14408 7990
rect 14438 8019 14469 8072
rect 14815 8065 14855 8245
rect 15193 8405 15233 8585
rect 15579 8578 15610 8631
rect 15640 8660 15677 8739
rect 15848 8736 16241 8756
rect 16261 8736 16264 8756
rect 16362 8740 16611 8762
rect 16780 8761 16821 8766
rect 17199 8763 17226 8941
rect 17877 8853 17904 9031
rect 18282 9028 18323 9033
rect 18492 9032 18741 9054
rect 18839 9038 18842 9058
rect 18862 9038 19255 9058
rect 19426 9055 19463 9134
rect 19493 9163 19524 9216
rect 19870 9209 19910 9389
rect 19870 9191 19880 9209
rect 19898 9191 19910 9209
rect 19870 9186 19910 9191
rect 19870 9182 19907 9186
rect 19543 9163 19580 9164
rect 19493 9154 19580 9163
rect 19493 9134 19551 9154
rect 19571 9134 19580 9154
rect 19493 9124 19580 9134
rect 19639 9154 19676 9164
rect 19639 9134 19647 9154
rect 19667 9134 19676 9154
rect 19493 9123 19524 9124
rect 19488 9055 19598 9068
rect 19639 9055 19676 9134
rect 19873 9119 19910 9120
rect 19869 9110 19910 9119
rect 19869 9092 19882 9110
rect 19900 9092 19910 9110
rect 19869 9083 19910 9092
rect 19869 9063 19909 9083
rect 19426 9053 19676 9055
rect 19426 9050 19527 9053
rect 17944 8993 18008 9005
rect 18284 9001 18321 9028
rect 18492 9001 18529 9032
rect 18705 9030 18741 9032
rect 19426 9031 19491 9050
rect 18705 9001 18742 9030
rect 19488 9023 19491 9031
rect 19520 9023 19527 9050
rect 19555 9026 19565 9053
rect 19594 9031 19676 9053
rect 19784 9053 19909 9063
rect 19784 9034 19792 9053
rect 19817 9034 19909 9053
rect 19594 9026 19598 9031
rect 19784 9027 19909 9034
rect 19555 9023 19598 9026
rect 19488 9009 19598 9023
rect 17944 8992 17979 8993
rect 17921 8987 17979 8992
rect 17921 8967 17924 8987
rect 17944 8973 17979 8987
rect 17999 8973 18008 8993
rect 17944 8965 18008 8973
rect 17970 8964 18008 8965
rect 17971 8963 18008 8964
rect 18074 8997 18110 8998
rect 18182 8997 18218 8998
rect 18074 8989 18218 8997
rect 18074 8969 18082 8989
rect 18102 8969 18190 8989
rect 18210 8969 18218 8989
rect 18074 8963 18218 8969
rect 18284 8993 18322 9001
rect 18390 8997 18426 8998
rect 18284 8973 18293 8993
rect 18313 8973 18322 8993
rect 18284 8964 18322 8973
rect 18341 8990 18426 8997
rect 18341 8970 18348 8990
rect 18369 8989 18426 8990
rect 18369 8970 18398 8989
rect 18341 8969 18398 8970
rect 18418 8969 18426 8989
rect 18284 8963 18321 8964
rect 18341 8963 18426 8969
rect 18492 8993 18530 9001
rect 18603 8997 18639 8998
rect 18492 8973 18501 8993
rect 18521 8973 18530 8993
rect 18492 8964 18530 8973
rect 18554 8989 18639 8997
rect 18554 8969 18611 8989
rect 18631 8969 18639 8989
rect 18492 8963 18529 8964
rect 18554 8963 18639 8969
rect 18705 8993 18743 9001
rect 18705 8973 18714 8993
rect 18734 8973 18743 8993
rect 18705 8964 18743 8973
rect 19869 8979 19909 9027
rect 18705 8963 18742 8964
rect 18128 8942 18164 8963
rect 18554 8942 18585 8963
rect 19869 8961 19880 8979
rect 19898 8961 19909 8979
rect 19869 8953 19909 8961
rect 19870 8952 19907 8953
rect 17961 8938 18061 8942
rect 17961 8934 18023 8938
rect 17961 8908 17968 8934
rect 17994 8912 18023 8934
rect 18049 8912 18061 8938
rect 17994 8908 18061 8912
rect 17961 8905 18061 8908
rect 18129 8905 18164 8942
rect 18226 8939 18585 8942
rect 18226 8934 18448 8939
rect 18226 8910 18239 8934
rect 18263 8915 18448 8934
rect 18472 8915 18585 8939
rect 18263 8910 18585 8915
rect 18226 8906 18585 8910
rect 18652 8934 18801 8942
rect 18652 8914 18663 8934
rect 18683 8914 18801 8934
rect 18652 8907 18801 8914
rect 19241 8911 19755 8912
rect 18652 8906 18693 8907
rect 18128 8870 18164 8905
rect 17976 8853 18013 8854
rect 18072 8853 18109 8854
rect 18128 8853 18135 8870
rect 17876 8844 18014 8853
rect 17876 8824 17985 8844
rect 18005 8824 18014 8844
rect 17876 8817 18014 8824
rect 18072 8844 18135 8853
rect 18072 8824 18081 8844
rect 18101 8829 18135 8844
rect 18156 8853 18164 8870
rect 18183 8853 18220 8854
rect 18156 8844 18220 8853
rect 18156 8829 18191 8844
rect 18101 8824 18191 8829
rect 18211 8824 18220 8844
rect 17876 8815 17972 8817
rect 18072 8814 18220 8824
rect 18279 8844 18316 8854
rect 18391 8853 18428 8854
rect 18372 8851 18428 8853
rect 18279 8824 18287 8844
rect 18307 8824 18316 8844
rect 18128 8813 18164 8814
rect 17058 8761 17226 8763
rect 16780 8755 17226 8761
rect 15848 8731 16264 8736
rect 16443 8734 16554 8740
rect 15848 8730 16189 8731
rect 15792 8670 15823 8671
rect 15640 8640 15649 8660
rect 15669 8640 15677 8660
rect 15640 8630 15677 8640
rect 15736 8663 15823 8670
rect 15736 8660 15797 8663
rect 15736 8640 15745 8660
rect 15765 8643 15797 8660
rect 15818 8643 15823 8663
rect 15765 8640 15823 8643
rect 15736 8633 15823 8640
rect 15848 8660 15885 8730
rect 16151 8729 16188 8730
rect 16443 8726 16484 8734
rect 16443 8706 16451 8726
rect 16470 8706 16484 8726
rect 16443 8704 16484 8706
rect 16512 8726 16554 8734
rect 16512 8706 16528 8726
rect 16547 8706 16554 8726
rect 16780 8733 16786 8755
rect 16812 8735 17226 8755
rect 17976 8754 18013 8755
rect 18279 8754 18316 8824
rect 18341 8844 18428 8851
rect 18341 8841 18399 8844
rect 18341 8821 18346 8841
rect 18367 8824 18399 8841
rect 18419 8824 18428 8844
rect 18367 8821 18428 8824
rect 18341 8814 18428 8821
rect 18487 8844 18524 8854
rect 18487 8824 18495 8844
rect 18515 8824 18524 8844
rect 18341 8813 18372 8814
rect 17975 8753 18316 8754
rect 16812 8733 16821 8735
rect 17058 8734 17226 8735
rect 17900 8752 18316 8753
rect 17900 8748 18276 8752
rect 16780 8724 16821 8733
rect 17900 8728 17903 8748
rect 17923 8735 18276 8748
rect 18308 8735 18316 8752
rect 17923 8728 18316 8735
rect 18487 8745 18524 8824
rect 18554 8853 18585 8906
rect 19222 8895 19755 8911
rect 19222 8884 19754 8895
rect 19873 8886 19910 8890
rect 18604 8853 18641 8854
rect 18554 8844 18641 8853
rect 18554 8824 18612 8844
rect 18632 8824 18641 8844
rect 18554 8814 18641 8824
rect 18700 8844 18737 8854
rect 18700 8824 18708 8844
rect 18728 8824 18737 8844
rect 18554 8813 18585 8814
rect 18549 8745 18659 8758
rect 18700 8745 18737 8824
rect 18487 8743 18737 8745
rect 18487 8740 18588 8743
rect 18487 8721 18552 8740
rect 16512 8704 16554 8706
rect 16443 8689 16554 8704
rect 18549 8713 18552 8721
rect 18581 8713 18588 8740
rect 18616 8716 18626 8743
rect 18655 8721 18737 8743
rect 18815 8815 18983 8816
rect 19222 8815 19260 8884
rect 18815 8795 19260 8815
rect 19487 8846 19598 8861
rect 19487 8844 19529 8846
rect 19487 8824 19494 8844
rect 19513 8824 19529 8844
rect 19487 8816 19529 8824
rect 19557 8844 19598 8846
rect 19557 8824 19571 8844
rect 19590 8824 19598 8844
rect 19557 8816 19598 8824
rect 19487 8810 19598 8816
rect 19720 8821 19754 8884
rect 19872 8880 19910 8886
rect 19872 8862 19882 8880
rect 19900 8862 19910 8880
rect 19872 8853 19910 8862
rect 19872 8821 19906 8853
rect 18815 8789 19259 8795
rect 18815 8787 18983 8789
rect 18655 8716 18659 8721
rect 18616 8713 18659 8716
rect 18549 8699 18659 8713
rect 16000 8670 16036 8671
rect 15848 8640 15857 8660
rect 15877 8640 15885 8660
rect 15736 8631 15792 8633
rect 15736 8630 15773 8631
rect 15848 8630 15885 8640
rect 15944 8660 16092 8670
rect 16192 8667 16288 8669
rect 15944 8640 15953 8660
rect 15973 8640 16063 8660
rect 16083 8640 16092 8660
rect 15944 8631 16092 8640
rect 16150 8660 16288 8667
rect 16150 8640 16159 8660
rect 16179 8640 16288 8660
rect 16150 8631 16288 8640
rect 15944 8630 15981 8631
rect 16000 8579 16036 8631
rect 16055 8630 16092 8631
rect 16151 8630 16188 8631
rect 15471 8577 15512 8578
rect 15363 8570 15512 8577
rect 15363 8550 15481 8570
rect 15501 8550 15512 8570
rect 15363 8542 15512 8550
rect 15579 8574 15938 8578
rect 15579 8569 15901 8574
rect 15579 8545 15692 8569
rect 15716 8550 15901 8569
rect 15925 8550 15938 8574
rect 15716 8545 15938 8550
rect 15579 8542 15938 8545
rect 16000 8542 16035 8579
rect 16103 8576 16203 8579
rect 16103 8572 16170 8576
rect 16103 8546 16115 8572
rect 16141 8550 16170 8572
rect 16196 8550 16203 8576
rect 16141 8546 16203 8550
rect 16103 8542 16203 8546
rect 15579 8521 15610 8542
rect 16000 8521 16036 8542
rect 15422 8520 15459 8521
rect 15421 8511 15459 8520
rect 15421 8491 15430 8511
rect 15450 8491 15459 8511
rect 15421 8483 15459 8491
rect 15525 8515 15610 8521
rect 15635 8520 15672 8521
rect 15525 8495 15533 8515
rect 15553 8495 15610 8515
rect 15525 8487 15610 8495
rect 15634 8511 15672 8520
rect 15634 8491 15643 8511
rect 15663 8491 15672 8511
rect 15525 8486 15561 8487
rect 15634 8483 15672 8491
rect 15738 8515 15823 8521
rect 15843 8520 15880 8521
rect 15738 8495 15746 8515
rect 15766 8514 15823 8515
rect 15766 8495 15795 8514
rect 15738 8494 15795 8495
rect 15816 8494 15823 8514
rect 15738 8487 15823 8494
rect 15842 8511 15880 8520
rect 15842 8491 15851 8511
rect 15871 8491 15880 8511
rect 15738 8486 15774 8487
rect 15842 8483 15880 8491
rect 15946 8515 16090 8521
rect 15946 8495 15954 8515
rect 15974 8512 16062 8515
rect 15974 8495 16005 8512
rect 15946 8492 16005 8495
rect 16028 8495 16062 8512
rect 16082 8495 16090 8515
rect 16028 8492 16090 8495
rect 15946 8487 16090 8492
rect 15946 8486 15982 8487
rect 16054 8486 16090 8487
rect 16156 8520 16193 8521
rect 16156 8519 16194 8520
rect 16156 8511 16220 8519
rect 16156 8491 16165 8511
rect 16185 8497 16220 8511
rect 16240 8497 16243 8517
rect 16185 8492 16243 8497
rect 16185 8491 16220 8492
rect 15422 8454 15459 8483
rect 15423 8452 15459 8454
rect 15635 8452 15672 8483
rect 15423 8430 15672 8452
rect 15843 8451 15880 8483
rect 16156 8479 16220 8491
rect 16260 8453 16287 8631
rect 18815 8609 18842 8787
rect 18882 8749 18946 8761
rect 19222 8757 19259 8789
rect 19430 8788 19679 8810
rect 19720 8789 19906 8821
rect 19734 8788 19906 8789
rect 19430 8757 19467 8788
rect 19643 8786 19679 8788
rect 19643 8757 19680 8786
rect 19872 8760 19906 8788
rect 18882 8748 18917 8749
rect 18859 8743 18917 8748
rect 18859 8723 18862 8743
rect 18882 8729 18917 8743
rect 18937 8729 18946 8749
rect 18882 8721 18946 8729
rect 18908 8720 18946 8721
rect 18909 8719 18946 8720
rect 19012 8753 19048 8754
rect 19120 8753 19156 8754
rect 19012 8746 19156 8753
rect 19012 8745 19072 8746
rect 19012 8725 19020 8745
rect 19040 8726 19072 8745
rect 19097 8745 19156 8746
rect 19097 8726 19128 8745
rect 19040 8725 19128 8726
rect 19148 8725 19156 8745
rect 19012 8719 19156 8725
rect 19222 8749 19260 8757
rect 19328 8753 19364 8754
rect 19222 8729 19231 8749
rect 19251 8729 19260 8749
rect 19222 8720 19260 8729
rect 19279 8746 19364 8753
rect 19279 8726 19286 8746
rect 19307 8745 19364 8746
rect 19307 8726 19336 8745
rect 19279 8725 19336 8726
rect 19356 8725 19364 8745
rect 19222 8719 19259 8720
rect 19279 8719 19364 8725
rect 19430 8749 19468 8757
rect 19541 8753 19577 8754
rect 19430 8729 19439 8749
rect 19459 8729 19468 8749
rect 19430 8720 19468 8729
rect 19492 8745 19577 8753
rect 19492 8725 19549 8745
rect 19569 8725 19577 8745
rect 19430 8719 19467 8720
rect 19492 8719 19577 8725
rect 19643 8749 19681 8757
rect 19643 8729 19652 8749
rect 19672 8729 19681 8749
rect 19643 8720 19681 8729
rect 19870 8750 19907 8760
rect 19870 8732 19880 8750
rect 19898 8732 19907 8750
rect 19870 8723 19907 8732
rect 19872 8722 19906 8723
rect 19643 8719 19680 8720
rect 19066 8698 19102 8719
rect 19492 8698 19523 8719
rect 18899 8694 18999 8698
rect 18899 8690 18961 8694
rect 18899 8664 18906 8690
rect 18932 8668 18961 8690
rect 18987 8668 18999 8694
rect 18932 8664 18999 8668
rect 18899 8661 18999 8664
rect 19067 8661 19102 8698
rect 19164 8695 19523 8698
rect 19164 8690 19386 8695
rect 19164 8666 19177 8690
rect 19201 8671 19386 8690
rect 19410 8671 19523 8695
rect 19201 8666 19523 8671
rect 19164 8662 19523 8666
rect 19590 8690 19739 8698
rect 19590 8670 19601 8690
rect 19621 8670 19739 8690
rect 19590 8663 19739 8670
rect 19590 8662 19631 8663
rect 18914 8609 18951 8610
rect 19010 8609 19047 8610
rect 19066 8609 19102 8661
rect 19121 8609 19158 8610
rect 18814 8600 18952 8609
rect 18409 8579 18520 8594
rect 18409 8577 18451 8579
rect 18079 8556 18184 8558
rect 17735 8548 17905 8549
rect 18079 8548 18128 8556
rect 17735 8529 18128 8548
rect 18159 8529 18184 8556
rect 18409 8557 18416 8577
rect 18435 8557 18451 8577
rect 18409 8549 18451 8557
rect 18479 8577 18520 8579
rect 18479 8557 18493 8577
rect 18512 8557 18520 8577
rect 18814 8580 18923 8600
rect 18943 8580 18952 8600
rect 18814 8573 18952 8580
rect 19010 8600 19158 8609
rect 19010 8580 19019 8600
rect 19039 8580 19129 8600
rect 19149 8580 19158 8600
rect 18814 8571 18910 8573
rect 19010 8570 19158 8580
rect 19217 8600 19254 8610
rect 19329 8609 19366 8610
rect 19310 8607 19366 8609
rect 19217 8580 19225 8600
rect 19245 8580 19254 8600
rect 19066 8569 19102 8570
rect 18479 8549 18520 8557
rect 18409 8543 18520 8549
rect 17735 8522 18184 8529
rect 17735 8520 17905 8522
rect 16585 8489 16695 8503
rect 16585 8486 16628 8489
rect 16585 8481 16589 8486
rect 16119 8451 16287 8453
rect 15843 8448 16287 8451
rect 15504 8424 15615 8430
rect 15504 8416 15545 8424
rect 15193 8361 15232 8405
rect 15504 8396 15512 8416
rect 15531 8396 15545 8416
rect 15504 8394 15545 8396
rect 15573 8416 15615 8424
rect 15573 8396 15589 8416
rect 15608 8396 15615 8416
rect 15573 8394 15615 8396
rect 15504 8379 15615 8394
rect 15841 8425 16287 8448
rect 15193 8337 15233 8361
rect 15533 8337 15580 8339
rect 15841 8337 15879 8425
rect 16119 8424 16287 8425
rect 16507 8459 16589 8481
rect 16618 8459 16628 8486
rect 16656 8462 16663 8489
rect 16692 8481 16695 8489
rect 16692 8462 16757 8481
rect 16656 8459 16757 8462
rect 16507 8457 16757 8459
rect 16507 8378 16544 8457
rect 16585 8444 16695 8457
rect 16659 8388 16690 8389
rect 16507 8358 16516 8378
rect 16536 8358 16544 8378
rect 16507 8348 16544 8358
rect 16603 8378 16690 8388
rect 16603 8358 16612 8378
rect 16632 8358 16690 8378
rect 16603 8349 16690 8358
rect 16603 8348 16640 8349
rect 15193 8304 15879 8337
rect 15193 8247 15232 8304
rect 15841 8302 15879 8304
rect 16659 8296 16690 8349
rect 16720 8378 16757 8457
rect 16928 8470 17321 8474
rect 16928 8453 16947 8470
rect 16967 8454 17321 8470
rect 17341 8454 17344 8474
rect 16967 8453 17344 8454
rect 16928 8449 17344 8453
rect 16928 8448 17269 8449
rect 16872 8388 16903 8389
rect 16720 8358 16729 8378
rect 16749 8358 16757 8378
rect 16720 8348 16757 8358
rect 16816 8381 16903 8388
rect 16816 8378 16877 8381
rect 16816 8358 16825 8378
rect 16845 8361 16877 8378
rect 16898 8361 16903 8381
rect 16845 8358 16903 8361
rect 16816 8351 16903 8358
rect 16928 8378 16965 8448
rect 17231 8447 17268 8448
rect 17080 8388 17116 8389
rect 16928 8358 16937 8378
rect 16957 8358 16965 8378
rect 16816 8349 16872 8351
rect 16816 8348 16853 8349
rect 16928 8348 16965 8358
rect 17024 8378 17172 8388
rect 17272 8385 17368 8387
rect 17024 8358 17033 8378
rect 17053 8358 17143 8378
rect 17163 8358 17172 8378
rect 17024 8349 17172 8358
rect 17230 8378 17368 8385
rect 17230 8358 17239 8378
rect 17259 8358 17368 8378
rect 17230 8349 17368 8358
rect 17024 8348 17061 8349
rect 17080 8297 17116 8349
rect 17135 8348 17172 8349
rect 17231 8348 17268 8349
rect 16551 8295 16592 8296
rect 16443 8288 16592 8295
rect 16443 8268 16561 8288
rect 16581 8268 16592 8288
rect 16443 8260 16592 8268
rect 16659 8292 17018 8296
rect 16659 8287 16981 8292
rect 16659 8263 16772 8287
rect 16796 8268 16981 8287
rect 17005 8268 17018 8292
rect 16796 8263 17018 8268
rect 16659 8260 17018 8263
rect 17080 8260 17115 8297
rect 17183 8294 17283 8297
rect 17183 8290 17250 8294
rect 17183 8264 17195 8290
rect 17221 8268 17250 8290
rect 17276 8268 17283 8294
rect 17221 8264 17283 8268
rect 17183 8260 17283 8264
rect 15193 8245 15241 8247
rect 15193 8227 15204 8245
rect 15222 8227 15241 8245
rect 16659 8239 16690 8260
rect 17080 8239 17116 8260
rect 16502 8238 16539 8239
rect 15193 8218 15241 8227
rect 15194 8217 15241 8218
rect 15507 8222 15617 8236
rect 15507 8219 15550 8222
rect 15507 8214 15511 8219
rect 15429 8192 15511 8214
rect 15540 8192 15550 8219
rect 15578 8195 15585 8222
rect 15614 8214 15617 8222
rect 16501 8229 16539 8238
rect 15614 8195 15679 8214
rect 16501 8209 16510 8229
rect 16530 8209 16539 8229
rect 15578 8192 15679 8195
rect 15429 8190 15679 8192
rect 15197 8154 15234 8155
rect 14815 8047 14825 8065
rect 14843 8047 14855 8065
rect 14815 8042 14855 8047
rect 15193 8151 15234 8154
rect 15193 8146 15235 8151
rect 15193 8128 15206 8146
rect 15224 8128 15235 8146
rect 15193 8114 15235 8128
rect 15273 8114 15320 8118
rect 15193 8108 15320 8114
rect 15193 8079 15281 8108
rect 15310 8079 15320 8108
rect 15429 8111 15466 8190
rect 15507 8177 15617 8190
rect 15581 8121 15612 8122
rect 15429 8091 15438 8111
rect 15458 8091 15466 8111
rect 15429 8081 15466 8091
rect 15525 8111 15612 8121
rect 15525 8091 15534 8111
rect 15554 8091 15612 8111
rect 15525 8082 15612 8091
rect 15525 8081 15562 8082
rect 15193 8075 15320 8079
rect 15193 8058 15232 8075
rect 15273 8074 15320 8075
rect 14815 8038 14852 8042
rect 15193 8040 15204 8058
rect 15222 8040 15232 8058
rect 15193 8031 15232 8040
rect 15194 8030 15231 8031
rect 15581 8029 15612 8082
rect 15642 8111 15679 8190
rect 15850 8187 16243 8207
rect 16263 8187 16266 8207
rect 16501 8201 16539 8209
rect 16605 8233 16690 8239
rect 16715 8238 16752 8239
rect 16605 8213 16613 8233
rect 16633 8213 16690 8233
rect 16605 8205 16690 8213
rect 16714 8229 16752 8238
rect 16714 8209 16723 8229
rect 16743 8209 16752 8229
rect 16605 8204 16641 8205
rect 16714 8201 16752 8209
rect 16818 8233 16903 8239
rect 16923 8238 16960 8239
rect 16818 8213 16826 8233
rect 16846 8232 16903 8233
rect 16846 8213 16875 8232
rect 16818 8212 16875 8213
rect 16896 8212 16903 8232
rect 16818 8205 16903 8212
rect 16922 8229 16960 8238
rect 16922 8209 16931 8229
rect 16951 8209 16960 8229
rect 16818 8204 16854 8205
rect 16922 8201 16960 8209
rect 17026 8233 17170 8239
rect 17026 8213 17034 8233
rect 17054 8231 17142 8233
rect 17054 8213 17083 8231
rect 17026 8210 17083 8213
rect 17110 8213 17142 8231
rect 17162 8213 17170 8233
rect 17110 8210 17170 8213
rect 17026 8205 17170 8210
rect 17026 8204 17062 8205
rect 17134 8204 17170 8205
rect 17236 8238 17273 8239
rect 17236 8237 17274 8238
rect 17236 8229 17300 8237
rect 17236 8209 17245 8229
rect 17265 8215 17300 8229
rect 17320 8215 17323 8235
rect 17265 8210 17323 8215
rect 17265 8209 17300 8210
rect 15850 8182 16266 8187
rect 15850 8181 16191 8182
rect 15794 8121 15825 8122
rect 15642 8091 15651 8111
rect 15671 8091 15679 8111
rect 15642 8081 15679 8091
rect 15738 8114 15825 8121
rect 15738 8111 15799 8114
rect 15738 8091 15747 8111
rect 15767 8094 15799 8111
rect 15820 8094 15825 8114
rect 15767 8091 15825 8094
rect 15738 8084 15825 8091
rect 15850 8111 15887 8181
rect 16153 8180 16190 8181
rect 16502 8172 16539 8201
rect 16503 8170 16539 8172
rect 16715 8170 16752 8201
rect 16503 8148 16752 8170
rect 16923 8169 16960 8201
rect 17236 8197 17300 8209
rect 17340 8171 17367 8349
rect 17735 8342 17764 8520
rect 17804 8482 17868 8494
rect 18144 8490 18181 8522
rect 18352 8521 18601 8543
rect 18352 8490 18389 8521
rect 18565 8519 18601 8521
rect 18565 8490 18602 8519
rect 18914 8510 18951 8511
rect 19217 8510 19254 8580
rect 19279 8600 19366 8607
rect 19279 8597 19337 8600
rect 19279 8577 19284 8597
rect 19305 8580 19337 8597
rect 19357 8580 19366 8600
rect 19305 8577 19366 8580
rect 19279 8570 19366 8577
rect 19425 8600 19462 8610
rect 19425 8580 19433 8600
rect 19453 8580 19462 8600
rect 19279 8569 19310 8570
rect 18913 8509 19254 8510
rect 18838 8504 19254 8509
rect 17804 8481 17839 8482
rect 17781 8476 17839 8481
rect 17781 8456 17784 8476
rect 17804 8462 17839 8476
rect 17859 8462 17868 8482
rect 17804 8454 17868 8462
rect 17830 8453 17868 8454
rect 17831 8452 17868 8453
rect 17934 8486 17970 8487
rect 18042 8486 18078 8487
rect 17934 8478 18078 8486
rect 17934 8458 17942 8478
rect 17962 8458 18050 8478
rect 18070 8458 18078 8478
rect 17934 8452 18078 8458
rect 18144 8482 18182 8490
rect 18250 8486 18286 8487
rect 18144 8462 18153 8482
rect 18173 8462 18182 8482
rect 18144 8453 18182 8462
rect 18201 8479 18286 8486
rect 18201 8459 18208 8479
rect 18229 8478 18286 8479
rect 18229 8459 18258 8478
rect 18201 8458 18258 8459
rect 18278 8458 18286 8478
rect 18144 8452 18181 8453
rect 18201 8452 18286 8458
rect 18352 8482 18390 8490
rect 18463 8486 18499 8487
rect 18352 8462 18361 8482
rect 18381 8462 18390 8482
rect 18352 8453 18390 8462
rect 18414 8478 18499 8486
rect 18414 8458 18471 8478
rect 18491 8458 18499 8478
rect 18352 8452 18389 8453
rect 18414 8452 18499 8458
rect 18565 8482 18603 8490
rect 18838 8484 18841 8504
rect 18861 8484 19254 8504
rect 19425 8501 19462 8580
rect 19492 8609 19523 8662
rect 19873 8660 19910 8661
rect 19872 8651 19911 8660
rect 19872 8633 19882 8651
rect 19900 8633 19911 8651
rect 19784 8616 19831 8617
rect 19872 8616 19911 8633
rect 19784 8612 19911 8616
rect 19542 8609 19579 8610
rect 19492 8600 19579 8609
rect 19492 8580 19550 8600
rect 19570 8580 19579 8600
rect 19492 8570 19579 8580
rect 19638 8600 19675 8610
rect 19638 8580 19646 8600
rect 19666 8580 19675 8600
rect 19492 8569 19523 8570
rect 19487 8501 19597 8514
rect 19638 8501 19675 8580
rect 19784 8583 19794 8612
rect 19823 8583 19911 8612
rect 19784 8577 19911 8583
rect 19784 8573 19831 8577
rect 19869 8563 19911 8577
rect 19869 8545 19880 8563
rect 19898 8545 19911 8563
rect 19869 8540 19911 8545
rect 19870 8537 19911 8540
rect 19870 8536 19907 8537
rect 19425 8499 19675 8501
rect 19425 8496 19526 8499
rect 18565 8462 18574 8482
rect 18594 8462 18603 8482
rect 19425 8477 19490 8496
rect 18565 8453 18603 8462
rect 19487 8469 19490 8477
rect 19519 8469 19526 8496
rect 19554 8472 19564 8499
rect 19593 8477 19675 8499
rect 19593 8472 19597 8477
rect 19554 8469 19597 8472
rect 19487 8455 19597 8469
rect 19863 8473 19910 8474
rect 19863 8464 19911 8473
rect 18565 8452 18602 8453
rect 17988 8431 18024 8452
rect 18414 8431 18445 8452
rect 19863 8446 19882 8464
rect 19900 8446 19911 8464
rect 19863 8444 19911 8446
rect 17821 8427 17921 8431
rect 17821 8423 17883 8427
rect 17821 8397 17828 8423
rect 17854 8401 17883 8423
rect 17909 8401 17921 8427
rect 17854 8397 17921 8401
rect 17821 8394 17921 8397
rect 17989 8394 18024 8431
rect 18086 8428 18445 8431
rect 18086 8423 18308 8428
rect 18086 8399 18099 8423
rect 18123 8404 18308 8423
rect 18332 8404 18445 8428
rect 18123 8399 18445 8404
rect 18086 8395 18445 8399
rect 18512 8423 18661 8431
rect 18512 8403 18523 8423
rect 18543 8403 18661 8423
rect 18512 8396 18661 8403
rect 18512 8395 18553 8396
rect 17988 8355 18024 8394
rect 17836 8342 17873 8343
rect 17932 8342 17969 8343
rect 17988 8342 17995 8355
rect 17735 8333 17874 8342
rect 17735 8313 17845 8333
rect 17865 8313 17874 8333
rect 17735 8306 17874 8313
rect 17932 8333 17995 8342
rect 17932 8313 17941 8333
rect 17961 8317 17995 8333
rect 18018 8342 18024 8355
rect 18043 8342 18080 8343
rect 18018 8333 18080 8342
rect 18018 8317 18051 8333
rect 17961 8313 18051 8317
rect 18071 8313 18080 8333
rect 17735 8304 17832 8306
rect 17735 8303 17764 8304
rect 17932 8303 18080 8313
rect 18139 8333 18176 8343
rect 18251 8342 18288 8343
rect 18232 8340 18288 8342
rect 18139 8313 18147 8333
rect 18167 8313 18176 8333
rect 17988 8302 18024 8303
rect 17836 8243 17873 8244
rect 18139 8243 18176 8313
rect 18201 8333 18288 8340
rect 18201 8330 18259 8333
rect 18201 8310 18206 8330
rect 18227 8313 18259 8330
rect 18279 8313 18288 8333
rect 18227 8310 18288 8313
rect 18201 8303 18288 8310
rect 18347 8333 18384 8343
rect 18347 8313 18355 8333
rect 18375 8313 18384 8333
rect 18201 8302 18232 8303
rect 17835 8242 18176 8243
rect 17760 8238 18176 8242
rect 17760 8237 18137 8238
rect 17760 8217 17763 8237
rect 17783 8221 18137 8237
rect 18157 8221 18176 8238
rect 17783 8217 18176 8221
rect 18347 8234 18384 8313
rect 18414 8342 18445 8395
rect 19225 8387 19263 8389
rect 19872 8387 19911 8444
rect 19225 8354 19911 8387
rect 18464 8342 18501 8343
rect 18414 8333 18501 8342
rect 18414 8313 18472 8333
rect 18492 8313 18501 8333
rect 18414 8303 18501 8313
rect 18560 8333 18597 8343
rect 18560 8313 18568 8333
rect 18588 8313 18597 8333
rect 18414 8302 18445 8303
rect 18409 8234 18519 8247
rect 18560 8234 18597 8313
rect 18347 8232 18597 8234
rect 18347 8229 18448 8232
rect 18347 8210 18412 8229
rect 18409 8202 18412 8210
rect 18441 8202 18448 8229
rect 18476 8205 18486 8232
rect 18515 8210 18597 8232
rect 18817 8266 18985 8267
rect 19225 8266 19263 8354
rect 19524 8352 19571 8354
rect 19871 8330 19911 8354
rect 18817 8243 19263 8266
rect 19489 8297 19600 8312
rect 19489 8295 19531 8297
rect 19489 8275 19496 8295
rect 19515 8275 19531 8295
rect 19489 8267 19531 8275
rect 19559 8295 19600 8297
rect 19559 8275 19573 8295
rect 19592 8275 19600 8295
rect 19872 8286 19911 8330
rect 19559 8267 19600 8275
rect 19489 8261 19600 8267
rect 18817 8240 19261 8243
rect 18817 8238 18985 8240
rect 18515 8205 18519 8210
rect 18476 8202 18519 8205
rect 18409 8188 18519 8202
rect 17199 8169 17367 8171
rect 16920 8162 17367 8169
rect 16584 8142 16695 8148
rect 16584 8134 16625 8142
rect 16002 8121 16038 8122
rect 15850 8091 15859 8111
rect 15879 8091 15887 8111
rect 15738 8082 15794 8084
rect 15738 8081 15775 8082
rect 15850 8081 15887 8091
rect 15946 8111 16094 8121
rect 16194 8118 16290 8120
rect 15946 8091 15955 8111
rect 15975 8091 16065 8111
rect 16085 8091 16094 8111
rect 15946 8082 16094 8091
rect 16152 8111 16290 8118
rect 16152 8091 16161 8111
rect 16181 8091 16290 8111
rect 16584 8114 16592 8134
rect 16611 8114 16625 8134
rect 16584 8112 16625 8114
rect 16653 8134 16695 8142
rect 16653 8114 16669 8134
rect 16688 8114 16695 8134
rect 16920 8135 16945 8162
rect 16976 8143 17367 8162
rect 16976 8135 17025 8143
rect 17199 8142 17367 8143
rect 16920 8133 17025 8135
rect 16653 8112 16695 8114
rect 16584 8097 16695 8112
rect 16152 8082 16290 8091
rect 15946 8081 15983 8082
rect 16002 8030 16038 8082
rect 16057 8081 16094 8082
rect 16153 8081 16190 8082
rect 15473 8028 15514 8029
rect 15365 8021 15514 8028
rect 14488 8019 14525 8020
rect 14438 8010 14525 8019
rect 14438 7990 14496 8010
rect 14516 7990 14525 8010
rect 14438 7980 14525 7990
rect 14584 8010 14621 8020
rect 14584 7990 14592 8010
rect 14612 7990 14621 8010
rect 15365 8001 15483 8021
rect 15503 8001 15514 8021
rect 15365 7993 15514 8001
rect 15581 8025 15940 8029
rect 15581 8020 15903 8025
rect 15581 7996 15694 8020
rect 15718 8001 15903 8020
rect 15927 8001 15940 8025
rect 15718 7996 15940 8001
rect 15581 7993 15940 7996
rect 16002 7993 16037 8030
rect 16105 8027 16205 8030
rect 16105 8023 16172 8027
rect 16105 7997 16117 8023
rect 16143 8001 16172 8023
rect 16198 8001 16205 8027
rect 16143 7997 16205 8001
rect 16105 7993 16205 7997
rect 14438 7979 14469 7980
rect 14433 7911 14543 7924
rect 14584 7911 14621 7990
rect 14818 7975 14855 7976
rect 14814 7966 14855 7975
rect 15581 7972 15612 7993
rect 16002 7972 16038 7993
rect 15424 7971 15461 7972
rect 15198 7968 15232 7969
rect 14814 7948 14827 7966
rect 14845 7948 14855 7966
rect 14814 7939 14855 7948
rect 15197 7959 15234 7968
rect 15197 7941 15206 7959
rect 15224 7941 15234 7959
rect 14814 7919 14854 7939
rect 15197 7931 15234 7941
rect 15423 7962 15461 7971
rect 15423 7942 15432 7962
rect 15452 7942 15461 7962
rect 15423 7934 15461 7942
rect 15527 7966 15612 7972
rect 15637 7971 15674 7972
rect 15527 7946 15535 7966
rect 15555 7946 15612 7966
rect 15527 7938 15612 7946
rect 15636 7962 15674 7971
rect 15636 7942 15645 7962
rect 15665 7942 15674 7962
rect 15527 7937 15563 7938
rect 15636 7934 15674 7942
rect 15740 7966 15825 7972
rect 15845 7971 15882 7972
rect 15740 7946 15748 7966
rect 15768 7965 15825 7966
rect 15768 7946 15797 7965
rect 15740 7945 15797 7946
rect 15818 7945 15825 7965
rect 15740 7938 15825 7945
rect 15844 7962 15882 7971
rect 15844 7942 15853 7962
rect 15873 7942 15882 7962
rect 15740 7937 15776 7938
rect 15844 7934 15882 7942
rect 15948 7966 16092 7972
rect 15948 7946 15956 7966
rect 15976 7965 16064 7966
rect 15976 7946 16007 7965
rect 15948 7945 16007 7946
rect 16032 7946 16064 7965
rect 16084 7946 16092 7966
rect 16032 7945 16092 7946
rect 15948 7938 16092 7945
rect 15948 7937 15984 7938
rect 16056 7937 16092 7938
rect 16158 7971 16195 7972
rect 16158 7970 16196 7971
rect 16158 7962 16222 7970
rect 16158 7942 16167 7962
rect 16187 7948 16222 7962
rect 16242 7948 16245 7968
rect 16187 7943 16245 7948
rect 16187 7942 16222 7943
rect 14371 7909 14621 7911
rect 14371 7906 14472 7909
rect 12889 7849 12953 7861
rect 13229 7857 13266 7884
rect 13437 7857 13474 7888
rect 13650 7886 13686 7888
rect 14371 7887 14436 7906
rect 13650 7857 13687 7886
rect 14433 7879 14436 7887
rect 14465 7879 14472 7906
rect 14500 7882 14510 7909
rect 14539 7887 14621 7909
rect 14729 7909 14854 7919
rect 14729 7890 14737 7909
rect 14762 7890 14854 7909
rect 14539 7882 14543 7887
rect 14729 7883 14854 7890
rect 14500 7879 14543 7882
rect 14433 7865 14543 7879
rect 12889 7848 12924 7849
rect 12866 7843 12924 7848
rect 12866 7823 12869 7843
rect 12889 7829 12924 7843
rect 12944 7829 12953 7849
rect 12889 7821 12953 7829
rect 12915 7820 12953 7821
rect 12916 7819 12953 7820
rect 13019 7853 13055 7854
rect 13127 7853 13163 7854
rect 13019 7845 13163 7853
rect 13019 7825 13027 7845
rect 13047 7842 13135 7845
rect 13047 7825 13079 7842
rect 13099 7825 13135 7842
rect 13155 7825 13163 7845
rect 13019 7819 13163 7825
rect 13229 7849 13267 7857
rect 13335 7853 13371 7854
rect 13229 7829 13238 7849
rect 13258 7829 13267 7849
rect 13229 7820 13267 7829
rect 13286 7846 13371 7853
rect 13286 7826 13293 7846
rect 13314 7845 13371 7846
rect 13314 7826 13343 7845
rect 13286 7825 13343 7826
rect 13363 7825 13371 7845
rect 13229 7819 13266 7820
rect 13286 7819 13371 7825
rect 13437 7849 13475 7857
rect 13548 7853 13584 7854
rect 13437 7829 13446 7849
rect 13466 7829 13475 7849
rect 13437 7820 13475 7829
rect 13499 7845 13584 7853
rect 13499 7825 13556 7845
rect 13576 7825 13584 7845
rect 13437 7819 13474 7820
rect 13499 7819 13584 7825
rect 13650 7849 13688 7857
rect 13650 7829 13659 7849
rect 13679 7829 13688 7849
rect 13650 7820 13688 7829
rect 14814 7835 14854 7883
rect 15198 7903 15232 7931
rect 15424 7905 15461 7934
rect 15425 7903 15461 7905
rect 15637 7903 15674 7934
rect 15198 7902 15370 7903
rect 15198 7870 15384 7902
rect 15425 7881 15674 7903
rect 15845 7902 15882 7934
rect 16158 7930 16222 7942
rect 16262 7904 16289 8082
rect 18817 8060 18844 8238
rect 18884 8200 18948 8212
rect 19224 8208 19261 8240
rect 19432 8239 19681 8261
rect 19432 8208 19469 8239
rect 19645 8237 19681 8239
rect 19645 8208 19682 8237
rect 18884 8199 18919 8200
rect 18861 8194 18919 8199
rect 18861 8174 18864 8194
rect 18884 8180 18919 8194
rect 18939 8180 18948 8200
rect 18884 8172 18948 8180
rect 18910 8171 18948 8172
rect 18911 8170 18948 8171
rect 19014 8204 19050 8205
rect 19122 8204 19158 8205
rect 19014 8199 19158 8204
rect 19014 8196 19076 8199
rect 19014 8176 19022 8196
rect 19042 8179 19076 8196
rect 19099 8196 19158 8199
rect 19099 8179 19130 8196
rect 19042 8176 19130 8179
rect 19150 8176 19158 8196
rect 19014 8170 19158 8176
rect 19224 8200 19262 8208
rect 19330 8204 19366 8205
rect 19224 8180 19233 8200
rect 19253 8180 19262 8200
rect 19224 8171 19262 8180
rect 19281 8197 19366 8204
rect 19281 8177 19288 8197
rect 19309 8196 19366 8197
rect 19309 8177 19338 8196
rect 19281 8176 19338 8177
rect 19358 8176 19366 8196
rect 19224 8170 19261 8171
rect 19281 8170 19366 8176
rect 19432 8200 19470 8208
rect 19543 8204 19579 8205
rect 19432 8180 19441 8200
rect 19461 8180 19470 8200
rect 19432 8171 19470 8180
rect 19494 8196 19579 8204
rect 19494 8176 19551 8196
rect 19571 8176 19579 8196
rect 19432 8170 19469 8171
rect 19494 8170 19579 8176
rect 19645 8200 19683 8208
rect 19645 8180 19654 8200
rect 19674 8180 19683 8200
rect 19645 8171 19683 8180
rect 19645 8170 19682 8171
rect 19068 8149 19104 8170
rect 19494 8149 19525 8170
rect 18901 8145 19001 8149
rect 18901 8141 18963 8145
rect 18901 8115 18908 8141
rect 18934 8119 18963 8141
rect 18989 8119 19001 8145
rect 18934 8115 19001 8119
rect 18901 8112 19001 8115
rect 19069 8112 19104 8149
rect 19166 8146 19525 8149
rect 19166 8141 19388 8146
rect 19166 8117 19179 8141
rect 19203 8122 19388 8141
rect 19412 8122 19525 8146
rect 19203 8117 19525 8122
rect 19166 8113 19525 8117
rect 19592 8141 19741 8149
rect 19592 8121 19603 8141
rect 19623 8121 19741 8141
rect 19592 8114 19741 8121
rect 19592 8113 19633 8114
rect 18916 8060 18953 8061
rect 19012 8060 19049 8061
rect 19068 8060 19104 8112
rect 19123 8060 19160 8061
rect 18816 8051 18954 8060
rect 18816 8031 18925 8051
rect 18945 8031 18954 8051
rect 18816 8024 18954 8031
rect 19012 8051 19160 8060
rect 19012 8031 19021 8051
rect 19041 8031 19131 8051
rect 19151 8031 19160 8051
rect 18816 8022 18912 8024
rect 19012 8021 19160 8031
rect 19219 8051 19256 8061
rect 19331 8060 19368 8061
rect 19312 8058 19368 8060
rect 19219 8031 19227 8051
rect 19247 8031 19256 8051
rect 19068 8020 19104 8021
rect 16445 7978 16555 7992
rect 16445 7975 16488 7978
rect 16445 7970 16449 7975
rect 16121 7902 16289 7904
rect 15845 7896 16289 7902
rect 15198 7838 15232 7870
rect 13650 7819 13687 7820
rect 13073 7798 13109 7819
rect 13499 7798 13530 7819
rect 14814 7817 14825 7835
rect 14843 7817 14854 7835
rect 14814 7809 14854 7817
rect 15194 7829 15232 7838
rect 15194 7811 15204 7829
rect 15222 7811 15232 7829
rect 14815 7808 14852 7809
rect 15194 7805 15232 7811
rect 15350 7807 15384 7870
rect 15506 7875 15617 7881
rect 15506 7867 15547 7875
rect 15506 7847 15514 7867
rect 15533 7847 15547 7867
rect 15506 7845 15547 7847
rect 15575 7867 15617 7875
rect 15575 7847 15591 7867
rect 15610 7847 15617 7867
rect 15575 7845 15617 7847
rect 15506 7830 15617 7845
rect 15844 7876 16289 7896
rect 15844 7807 15882 7876
rect 16121 7875 16289 7876
rect 16367 7948 16449 7970
rect 16478 7948 16488 7975
rect 16516 7951 16523 7978
rect 16552 7970 16555 7978
rect 18550 7987 18661 8002
rect 18550 7985 18592 7987
rect 16552 7951 16617 7970
rect 16516 7948 16617 7951
rect 16367 7946 16617 7948
rect 16367 7867 16404 7946
rect 16445 7933 16555 7946
rect 16519 7877 16550 7878
rect 16367 7847 16376 7867
rect 16396 7847 16404 7867
rect 16367 7837 16404 7847
rect 16463 7867 16550 7877
rect 16463 7847 16472 7867
rect 16492 7847 16550 7867
rect 16463 7838 16550 7847
rect 16463 7837 16500 7838
rect 15194 7801 15231 7805
rect 12906 7794 13006 7798
rect 12906 7790 12968 7794
rect 12906 7764 12913 7790
rect 12939 7768 12968 7790
rect 12994 7768 13006 7794
rect 12939 7764 13006 7768
rect 12906 7761 13006 7764
rect 13074 7761 13109 7798
rect 13171 7795 13530 7798
rect 13171 7790 13393 7795
rect 13171 7766 13184 7790
rect 13208 7771 13393 7790
rect 13417 7771 13530 7795
rect 13208 7766 13530 7771
rect 13171 7762 13530 7766
rect 13597 7790 13746 7798
rect 15350 7796 15882 7807
rect 13597 7770 13608 7790
rect 13628 7770 13746 7790
rect 15349 7780 15882 7796
rect 16519 7785 16550 7838
rect 16580 7867 16617 7946
rect 16788 7956 17181 7963
rect 16788 7939 16796 7956
rect 16828 7943 17181 7956
rect 17201 7943 17204 7963
rect 18283 7958 18324 7967
rect 16828 7939 17204 7943
rect 16788 7938 17204 7939
rect 17878 7956 18046 7957
rect 18283 7956 18292 7958
rect 16788 7937 17129 7938
rect 16732 7877 16763 7878
rect 16580 7847 16589 7867
rect 16609 7847 16617 7867
rect 16580 7837 16617 7847
rect 16676 7870 16763 7877
rect 16676 7867 16737 7870
rect 16676 7847 16685 7867
rect 16705 7850 16737 7867
rect 16758 7850 16763 7870
rect 16705 7847 16763 7850
rect 16676 7840 16763 7847
rect 16788 7867 16825 7937
rect 17091 7936 17128 7937
rect 17878 7936 18292 7956
rect 18318 7936 18324 7958
rect 18550 7965 18557 7985
rect 18576 7965 18592 7985
rect 18550 7957 18592 7965
rect 18620 7985 18661 7987
rect 18620 7965 18634 7985
rect 18653 7965 18661 7985
rect 18620 7957 18661 7965
rect 18916 7961 18953 7962
rect 19219 7961 19256 8031
rect 19281 8051 19368 8058
rect 19281 8048 19339 8051
rect 19281 8028 19286 8048
rect 19307 8031 19339 8048
rect 19359 8031 19368 8051
rect 19307 8028 19368 8031
rect 19281 8021 19368 8028
rect 19427 8051 19464 8061
rect 19427 8031 19435 8051
rect 19455 8031 19464 8051
rect 19281 8020 19312 8021
rect 18915 7960 19256 7961
rect 18550 7951 18661 7957
rect 18840 7955 19256 7960
rect 17878 7930 18324 7936
rect 17878 7928 18046 7930
rect 16940 7877 16976 7878
rect 16788 7847 16797 7867
rect 16817 7847 16825 7867
rect 16676 7838 16732 7840
rect 16676 7837 16713 7838
rect 16788 7837 16825 7847
rect 16884 7867 17032 7877
rect 17132 7874 17228 7876
rect 16884 7847 16893 7867
rect 16913 7862 17003 7867
rect 16913 7847 16948 7862
rect 16884 7838 16948 7847
rect 16884 7837 16921 7838
rect 16940 7821 16948 7838
rect 16969 7847 17003 7862
rect 17023 7847 17032 7867
rect 16969 7838 17032 7847
rect 17090 7867 17228 7874
rect 17090 7847 17099 7867
rect 17119 7847 17228 7867
rect 17090 7838 17228 7847
rect 16969 7821 16976 7838
rect 16995 7837 17032 7838
rect 17091 7837 17128 7838
rect 16940 7786 16976 7821
rect 16411 7784 16452 7785
rect 15349 7779 15863 7780
rect 13597 7763 13746 7770
rect 16303 7777 16452 7784
rect 14186 7767 14700 7768
rect 13597 7762 13638 7763
rect 12921 7709 12958 7710
rect 13017 7709 13054 7710
rect 13073 7709 13109 7761
rect 13128 7709 13165 7710
rect 12821 7700 12959 7709
rect 12821 7680 12930 7700
rect 12950 7680 12959 7700
rect 12821 7673 12959 7680
rect 13017 7700 13165 7709
rect 13017 7680 13026 7700
rect 13046 7680 13136 7700
rect 13156 7680 13165 7700
rect 12821 7671 12917 7673
rect 13017 7670 13165 7680
rect 13224 7700 13261 7710
rect 13336 7709 13373 7710
rect 13317 7707 13373 7709
rect 13224 7680 13232 7700
rect 13252 7680 13261 7700
rect 13073 7669 13109 7670
rect 12003 7617 12171 7619
rect 11725 7611 12171 7617
rect 10793 7587 11209 7592
rect 11388 7590 11499 7596
rect 10793 7586 11134 7587
rect 10737 7526 10768 7527
rect 10585 7496 10594 7516
rect 10614 7496 10622 7516
rect 10585 7486 10622 7496
rect 10681 7519 10768 7526
rect 10681 7516 10742 7519
rect 10681 7496 10690 7516
rect 10710 7499 10742 7516
rect 10763 7499 10768 7519
rect 10710 7496 10768 7499
rect 10681 7489 10768 7496
rect 10793 7516 10830 7586
rect 11096 7585 11133 7586
rect 11388 7582 11429 7590
rect 11388 7562 11396 7582
rect 11415 7562 11429 7582
rect 11388 7560 11429 7562
rect 11457 7582 11499 7590
rect 11457 7562 11473 7582
rect 11492 7562 11499 7582
rect 11725 7589 11731 7611
rect 11757 7591 12171 7611
rect 12921 7610 12958 7611
rect 13224 7610 13261 7680
rect 13286 7700 13373 7707
rect 13286 7697 13344 7700
rect 13286 7677 13291 7697
rect 13312 7680 13344 7697
rect 13364 7680 13373 7700
rect 13312 7677 13373 7680
rect 13286 7670 13373 7677
rect 13432 7700 13469 7710
rect 13432 7680 13440 7700
rect 13460 7680 13469 7700
rect 13286 7669 13317 7670
rect 12920 7609 13261 7610
rect 11757 7589 11766 7591
rect 12003 7590 12171 7591
rect 12845 7604 13261 7609
rect 11725 7580 11766 7589
rect 12845 7584 12848 7604
rect 12868 7584 13261 7604
rect 13432 7601 13469 7680
rect 13499 7709 13530 7762
rect 14167 7751 14700 7767
rect 16303 7757 16421 7777
rect 16441 7757 16452 7777
rect 14167 7740 14699 7751
rect 16303 7749 16452 7757
rect 16519 7781 16878 7785
rect 16519 7776 16841 7781
rect 16519 7752 16632 7776
rect 16656 7757 16841 7776
rect 16865 7757 16878 7781
rect 16656 7752 16878 7757
rect 16519 7749 16878 7752
rect 16940 7749 16975 7786
rect 17043 7783 17143 7786
rect 17043 7779 17110 7783
rect 17043 7753 17055 7779
rect 17081 7757 17110 7779
rect 17136 7757 17143 7783
rect 17081 7753 17143 7757
rect 17043 7749 17143 7753
rect 14818 7742 14855 7746
rect 13549 7709 13586 7710
rect 13499 7700 13586 7709
rect 13499 7680 13557 7700
rect 13577 7680 13586 7700
rect 13499 7670 13586 7680
rect 13645 7700 13682 7710
rect 13645 7680 13653 7700
rect 13673 7680 13682 7700
rect 13499 7669 13530 7670
rect 13494 7601 13604 7614
rect 13645 7601 13682 7680
rect 13432 7599 13682 7601
rect 13432 7596 13533 7599
rect 13432 7577 13497 7596
rect 11457 7560 11499 7562
rect 11388 7545 11499 7560
rect 13494 7569 13497 7577
rect 13526 7569 13533 7596
rect 13561 7572 13571 7599
rect 13600 7577 13682 7599
rect 13760 7671 13928 7672
rect 14167 7671 14205 7740
rect 13760 7651 14205 7671
rect 14432 7702 14543 7717
rect 14432 7700 14474 7702
rect 14432 7680 14439 7700
rect 14458 7680 14474 7700
rect 14432 7672 14474 7680
rect 14502 7700 14543 7702
rect 14502 7680 14516 7700
rect 14535 7680 14543 7700
rect 14502 7672 14543 7680
rect 14432 7666 14543 7672
rect 14665 7677 14699 7740
rect 14817 7736 14855 7742
rect 15197 7738 15234 7739
rect 14817 7718 14827 7736
rect 14845 7718 14855 7736
rect 14817 7709 14855 7718
rect 15195 7730 15235 7738
rect 15195 7712 15206 7730
rect 15224 7712 15235 7730
rect 16519 7728 16550 7749
rect 16940 7728 16976 7749
rect 16362 7727 16399 7728
rect 14817 7677 14851 7709
rect 13760 7645 14204 7651
rect 13760 7643 13928 7645
rect 13600 7572 13604 7577
rect 13561 7569 13604 7572
rect 13494 7555 13604 7569
rect 10945 7526 10981 7527
rect 10793 7496 10802 7516
rect 10822 7496 10830 7516
rect 10681 7487 10737 7489
rect 10681 7486 10718 7487
rect 10793 7486 10830 7496
rect 10889 7516 11037 7526
rect 11137 7523 11233 7525
rect 10889 7496 10898 7516
rect 10918 7496 11008 7516
rect 11028 7496 11037 7516
rect 10889 7487 11037 7496
rect 11095 7516 11233 7523
rect 11095 7496 11104 7516
rect 11124 7496 11233 7516
rect 11095 7487 11233 7496
rect 10889 7486 10926 7487
rect 10945 7435 10981 7487
rect 11000 7486 11037 7487
rect 11096 7486 11133 7487
rect 10416 7433 10457 7434
rect 10308 7426 10457 7433
rect 10308 7406 10426 7426
rect 10446 7406 10457 7426
rect 10308 7398 10457 7406
rect 10524 7430 10883 7434
rect 10524 7425 10846 7430
rect 10524 7401 10637 7425
rect 10661 7406 10846 7425
rect 10870 7406 10883 7430
rect 10661 7401 10883 7406
rect 10524 7398 10883 7401
rect 10945 7398 10980 7435
rect 11048 7432 11148 7435
rect 11048 7428 11115 7432
rect 11048 7402 11060 7428
rect 11086 7406 11115 7428
rect 11141 7406 11148 7432
rect 11086 7402 11148 7406
rect 11048 7398 11148 7402
rect 10524 7377 10555 7398
rect 10945 7377 10981 7398
rect 10367 7376 10404 7377
rect 10366 7367 10404 7376
rect 10366 7347 10375 7367
rect 10395 7347 10404 7367
rect 10366 7339 10404 7347
rect 10470 7371 10555 7377
rect 10580 7376 10617 7377
rect 10470 7351 10478 7371
rect 10498 7351 10555 7371
rect 10470 7343 10555 7351
rect 10579 7367 10617 7376
rect 10579 7347 10588 7367
rect 10608 7347 10617 7367
rect 10470 7342 10506 7343
rect 10579 7339 10617 7347
rect 10683 7371 10768 7377
rect 10788 7376 10825 7377
rect 10683 7351 10691 7371
rect 10711 7370 10768 7371
rect 10711 7351 10740 7370
rect 10683 7350 10740 7351
rect 10761 7350 10768 7370
rect 10683 7343 10768 7350
rect 10787 7367 10825 7376
rect 10787 7347 10796 7367
rect 10816 7347 10825 7367
rect 10683 7342 10719 7343
rect 10787 7339 10825 7347
rect 10891 7371 11035 7377
rect 10891 7351 10899 7371
rect 10919 7368 11007 7371
rect 10919 7351 10950 7368
rect 10891 7348 10950 7351
rect 10973 7351 11007 7368
rect 11027 7351 11035 7371
rect 10973 7348 11035 7351
rect 10891 7343 11035 7348
rect 10891 7342 10927 7343
rect 10999 7342 11035 7343
rect 11101 7376 11138 7377
rect 11101 7375 11139 7376
rect 11101 7367 11165 7375
rect 11101 7347 11110 7367
rect 11130 7353 11165 7367
rect 11185 7353 11188 7373
rect 11130 7348 11188 7353
rect 11130 7347 11165 7348
rect 10367 7310 10404 7339
rect 10368 7308 10404 7310
rect 10580 7308 10617 7339
rect 10368 7286 10617 7308
rect 10788 7307 10825 7339
rect 11101 7335 11165 7347
rect 11205 7309 11232 7487
rect 13760 7465 13787 7643
rect 13827 7605 13891 7617
rect 14167 7613 14204 7645
rect 14375 7644 14624 7666
rect 14665 7645 14851 7677
rect 14679 7644 14851 7645
rect 14375 7613 14412 7644
rect 14588 7642 14624 7644
rect 14588 7613 14625 7642
rect 14817 7616 14851 7644
rect 15195 7664 15235 7712
rect 16361 7718 16399 7727
rect 16361 7698 16370 7718
rect 16390 7698 16399 7718
rect 16361 7690 16399 7698
rect 16465 7722 16550 7728
rect 16575 7727 16612 7728
rect 16465 7702 16473 7722
rect 16493 7702 16550 7722
rect 16465 7694 16550 7702
rect 16574 7718 16612 7727
rect 16574 7698 16583 7718
rect 16603 7698 16612 7718
rect 16465 7693 16501 7694
rect 16574 7690 16612 7698
rect 16678 7722 16763 7728
rect 16783 7727 16820 7728
rect 16678 7702 16686 7722
rect 16706 7721 16763 7722
rect 16706 7702 16735 7721
rect 16678 7701 16735 7702
rect 16756 7701 16763 7721
rect 16678 7694 16763 7701
rect 16782 7718 16820 7727
rect 16782 7698 16791 7718
rect 16811 7698 16820 7718
rect 16678 7693 16714 7694
rect 16782 7690 16820 7698
rect 16886 7722 17030 7728
rect 16886 7702 16894 7722
rect 16914 7702 17002 7722
rect 17022 7702 17030 7722
rect 16886 7694 17030 7702
rect 16886 7693 16922 7694
rect 16994 7693 17030 7694
rect 17096 7727 17133 7728
rect 17096 7726 17134 7727
rect 17096 7718 17160 7726
rect 17096 7698 17105 7718
rect 17125 7704 17160 7718
rect 17180 7704 17183 7724
rect 17125 7699 17183 7704
rect 17125 7698 17160 7699
rect 15506 7668 15616 7682
rect 15506 7665 15549 7668
rect 15195 7657 15320 7664
rect 15506 7660 15510 7665
rect 15195 7638 15287 7657
rect 15312 7638 15320 7657
rect 15195 7628 15320 7638
rect 15428 7638 15510 7660
rect 15539 7638 15549 7665
rect 15577 7641 15584 7668
rect 15613 7660 15616 7668
rect 16362 7661 16399 7690
rect 15613 7641 15678 7660
rect 16363 7659 16399 7661
rect 16575 7659 16612 7690
rect 16783 7663 16820 7690
rect 17096 7686 17160 7698
rect 15577 7638 15678 7641
rect 15428 7636 15678 7638
rect 13827 7604 13862 7605
rect 13804 7599 13862 7604
rect 13804 7579 13807 7599
rect 13827 7585 13862 7599
rect 13882 7585 13891 7605
rect 13827 7577 13891 7585
rect 13853 7576 13891 7577
rect 13854 7575 13891 7576
rect 13957 7609 13993 7610
rect 14065 7609 14101 7610
rect 13957 7602 14101 7609
rect 13957 7601 14017 7602
rect 13957 7581 13965 7601
rect 13985 7582 14017 7601
rect 14042 7601 14101 7602
rect 14042 7582 14073 7601
rect 13985 7581 14073 7582
rect 14093 7581 14101 7601
rect 13957 7575 14101 7581
rect 14167 7605 14205 7613
rect 14273 7609 14309 7610
rect 14167 7585 14176 7605
rect 14196 7585 14205 7605
rect 14167 7576 14205 7585
rect 14224 7602 14309 7609
rect 14224 7582 14231 7602
rect 14252 7601 14309 7602
rect 14252 7582 14281 7601
rect 14224 7581 14281 7582
rect 14301 7581 14309 7601
rect 14167 7575 14204 7576
rect 14224 7575 14309 7581
rect 14375 7605 14413 7613
rect 14486 7609 14522 7610
rect 14375 7585 14384 7605
rect 14404 7585 14413 7605
rect 14375 7576 14413 7585
rect 14437 7601 14522 7609
rect 14437 7581 14494 7601
rect 14514 7581 14522 7601
rect 14375 7575 14412 7576
rect 14437 7575 14522 7581
rect 14588 7605 14626 7613
rect 14588 7585 14597 7605
rect 14617 7585 14626 7605
rect 14588 7576 14626 7585
rect 14815 7606 14852 7616
rect 15195 7608 15235 7628
rect 14815 7588 14825 7606
rect 14843 7588 14852 7606
rect 14815 7579 14852 7588
rect 15194 7599 15235 7608
rect 15194 7581 15204 7599
rect 15222 7581 15235 7599
rect 14817 7578 14851 7579
rect 14588 7575 14625 7576
rect 14011 7554 14047 7575
rect 14437 7554 14468 7575
rect 15194 7572 15235 7581
rect 15194 7571 15231 7572
rect 15428 7557 15465 7636
rect 15506 7623 15616 7636
rect 15580 7567 15611 7568
rect 13844 7550 13944 7554
rect 13844 7546 13906 7550
rect 13844 7520 13851 7546
rect 13877 7524 13906 7546
rect 13932 7524 13944 7550
rect 13877 7520 13944 7524
rect 13844 7517 13944 7520
rect 14012 7517 14047 7554
rect 14109 7551 14468 7554
rect 14109 7546 14331 7551
rect 14109 7522 14122 7546
rect 14146 7527 14331 7546
rect 14355 7527 14468 7551
rect 14146 7522 14468 7527
rect 14109 7518 14468 7522
rect 14535 7546 14684 7554
rect 14535 7526 14546 7546
rect 14566 7526 14684 7546
rect 15428 7537 15437 7557
rect 15457 7537 15465 7557
rect 15428 7527 15465 7537
rect 15524 7557 15611 7567
rect 15524 7537 15533 7557
rect 15553 7537 15611 7557
rect 15524 7528 15611 7537
rect 15524 7527 15561 7528
rect 14535 7519 14684 7526
rect 14535 7518 14576 7519
rect 13859 7465 13896 7466
rect 13955 7465 13992 7466
rect 14011 7465 14047 7517
rect 14066 7465 14103 7466
rect 13759 7456 13897 7465
rect 13384 7422 13495 7437
rect 13759 7436 13868 7456
rect 13888 7436 13897 7456
rect 13759 7429 13897 7436
rect 13955 7456 14103 7465
rect 13955 7436 13964 7456
rect 13984 7436 14074 7456
rect 14094 7436 14103 7456
rect 13759 7427 13855 7429
rect 13955 7426 14103 7436
rect 14162 7456 14199 7466
rect 14274 7465 14311 7466
rect 14255 7463 14311 7465
rect 14162 7436 14170 7456
rect 14190 7436 14199 7456
rect 14011 7425 14047 7426
rect 13384 7420 13426 7422
rect 12721 7401 12791 7410
rect 12721 7392 12738 7401
rect 12712 7372 12738 7392
rect 12786 7392 12791 7401
rect 13384 7400 13391 7420
rect 13410 7400 13426 7420
rect 13384 7392 13426 7400
rect 13454 7420 13495 7422
rect 13454 7400 13468 7420
rect 13487 7400 13495 7420
rect 13454 7392 13495 7400
rect 12786 7391 12880 7392
rect 12786 7372 13156 7391
rect 13384 7386 13495 7392
rect 11499 7358 11609 7372
rect 11499 7355 11542 7358
rect 11499 7350 11503 7355
rect 11064 7307 11232 7309
rect 10788 7304 11232 7307
rect 10449 7280 10560 7286
rect 10449 7272 10490 7280
rect 10138 7217 10177 7261
rect 10449 7252 10457 7272
rect 10476 7252 10490 7272
rect 10449 7250 10490 7252
rect 10518 7272 10560 7280
rect 10518 7252 10534 7272
rect 10553 7252 10560 7272
rect 10518 7250 10560 7252
rect 10449 7236 10560 7250
rect 10786 7281 11232 7304
rect 10138 7193 10178 7217
rect 10478 7193 10525 7195
rect 10786 7193 10824 7281
rect 11064 7280 11232 7281
rect 11421 7328 11503 7350
rect 11532 7328 11542 7355
rect 11570 7331 11577 7358
rect 11606 7350 11609 7358
rect 12712 7365 13156 7372
rect 12712 7363 12880 7365
rect 12712 7355 12791 7363
rect 11606 7331 11671 7350
rect 11570 7328 11671 7331
rect 11421 7326 11671 7328
rect 11421 7247 11458 7326
rect 11499 7313 11609 7326
rect 11573 7257 11604 7258
rect 11421 7227 11430 7247
rect 11450 7227 11458 7247
rect 11421 7217 11458 7227
rect 11517 7247 11604 7257
rect 11517 7227 11526 7247
rect 11546 7227 11604 7247
rect 11517 7218 11604 7227
rect 11517 7217 11554 7218
rect 10138 7160 10824 7193
rect 11573 7165 11604 7218
rect 11634 7247 11671 7326
rect 11842 7323 12235 7343
rect 12255 7323 12258 7343
rect 11842 7318 12258 7323
rect 11842 7317 12183 7318
rect 11786 7257 11817 7258
rect 11634 7227 11643 7247
rect 11663 7227 11671 7247
rect 11634 7217 11671 7227
rect 11730 7250 11817 7257
rect 11730 7247 11791 7250
rect 11730 7227 11739 7247
rect 11759 7230 11791 7247
rect 11812 7230 11817 7250
rect 11759 7227 11817 7230
rect 11730 7220 11817 7227
rect 11842 7247 11879 7317
rect 12145 7316 12182 7317
rect 11994 7257 12030 7258
rect 11842 7227 11851 7247
rect 11871 7227 11879 7247
rect 11730 7218 11786 7220
rect 11730 7217 11767 7218
rect 11842 7217 11879 7227
rect 11938 7247 12086 7257
rect 12186 7254 12282 7256
rect 11938 7227 11947 7247
rect 11967 7227 12057 7247
rect 12077 7227 12086 7247
rect 11938 7218 12086 7227
rect 12144 7247 12282 7254
rect 12144 7227 12153 7247
rect 12173 7227 12282 7247
rect 12144 7218 12282 7227
rect 11938 7217 11975 7218
rect 11994 7166 12030 7218
rect 12049 7217 12086 7218
rect 12145 7217 12182 7218
rect 11465 7164 11506 7165
rect 10137 7103 10176 7160
rect 10786 7158 10824 7160
rect 11357 7157 11506 7164
rect 11357 7137 11475 7157
rect 11495 7137 11506 7157
rect 11357 7129 11506 7137
rect 11573 7161 11932 7165
rect 11573 7156 11895 7161
rect 11573 7132 11686 7156
rect 11710 7137 11895 7156
rect 11919 7137 11932 7161
rect 11710 7132 11932 7137
rect 11573 7129 11932 7132
rect 11994 7129 12029 7166
rect 12097 7163 12197 7166
rect 12097 7159 12164 7163
rect 12097 7133 12109 7159
rect 12135 7137 12164 7159
rect 12190 7137 12197 7163
rect 12135 7133 12197 7137
rect 12097 7129 12197 7133
rect 11573 7108 11604 7129
rect 11994 7108 12030 7129
rect 11416 7107 11453 7108
rect 10137 7101 10185 7103
rect 10137 7083 10148 7101
rect 10166 7083 10185 7101
rect 11415 7098 11453 7107
rect 10137 7074 10185 7083
rect 10138 7073 10185 7074
rect 10451 7078 10561 7092
rect 10451 7075 10494 7078
rect 10451 7070 10455 7075
rect 10373 7048 10455 7070
rect 10484 7048 10494 7075
rect 10522 7051 10529 7078
rect 10558 7070 10561 7078
rect 11415 7078 11424 7098
rect 11444 7078 11453 7098
rect 11415 7070 11453 7078
rect 11519 7102 11604 7108
rect 11629 7107 11666 7108
rect 11519 7082 11527 7102
rect 11547 7082 11604 7102
rect 11519 7074 11604 7082
rect 11628 7098 11666 7107
rect 11628 7078 11637 7098
rect 11657 7078 11666 7098
rect 11519 7073 11555 7074
rect 11628 7070 11666 7078
rect 11732 7102 11817 7108
rect 11837 7107 11874 7108
rect 11732 7082 11740 7102
rect 11760 7101 11817 7102
rect 11760 7082 11789 7101
rect 11732 7081 11789 7082
rect 11810 7081 11817 7101
rect 11732 7074 11817 7081
rect 11836 7098 11874 7107
rect 11836 7078 11845 7098
rect 11865 7078 11874 7098
rect 11732 7073 11768 7074
rect 11836 7070 11874 7078
rect 11940 7102 12084 7108
rect 11940 7082 11948 7102
rect 11968 7100 12056 7102
rect 11968 7082 11997 7100
rect 11940 7081 11997 7082
rect 12026 7082 12056 7100
rect 12076 7082 12084 7102
rect 12026 7081 12084 7082
rect 11940 7074 12084 7081
rect 11940 7073 11976 7074
rect 12048 7073 12084 7074
rect 12150 7107 12187 7108
rect 12150 7106 12188 7107
rect 12150 7098 12214 7106
rect 12150 7078 12159 7098
rect 12179 7084 12214 7098
rect 12234 7084 12237 7104
rect 12179 7079 12237 7084
rect 12179 7078 12214 7079
rect 10558 7051 10623 7070
rect 10522 7048 10623 7051
rect 10373 7046 10623 7048
rect 10141 7010 10178 7011
rect 9840 6980 9850 6998
rect 9868 6980 9880 6998
rect 9840 6975 9880 6980
rect 10137 7007 10178 7010
rect 10137 7002 10179 7007
rect 10137 6984 10150 7002
rect 10168 6984 10179 7002
rect 9840 6971 9877 6975
rect 10137 6970 10179 6984
rect 10217 6970 10264 6974
rect 10137 6964 10264 6970
rect 9513 6952 9550 6953
rect 9463 6943 9550 6952
rect 9463 6923 9521 6943
rect 9541 6923 9550 6943
rect 9463 6913 9550 6923
rect 9609 6943 9646 6953
rect 9609 6923 9617 6943
rect 9637 6923 9646 6943
rect 9463 6912 9494 6913
rect 9458 6844 9568 6857
rect 9609 6844 9646 6923
rect 10137 6935 10225 6964
rect 10254 6935 10264 6964
rect 10373 6967 10410 7046
rect 10451 7033 10561 7046
rect 10525 6977 10556 6978
rect 10373 6947 10382 6967
rect 10402 6947 10410 6967
rect 10373 6937 10410 6947
rect 10469 6967 10556 6977
rect 10469 6947 10478 6967
rect 10498 6947 10556 6967
rect 10469 6938 10556 6947
rect 10469 6937 10506 6938
rect 10137 6931 10264 6935
rect 10137 6914 10176 6931
rect 10217 6930 10264 6931
rect 9843 6908 9880 6909
rect 9839 6899 9880 6908
rect 9839 6881 9852 6899
rect 9870 6881 9880 6899
rect 10137 6896 10148 6914
rect 10166 6896 10176 6914
rect 10137 6887 10176 6896
rect 10138 6886 10175 6887
rect 10525 6885 10556 6938
rect 10586 6967 10623 7046
rect 10794 7043 11187 7063
rect 11207 7043 11210 7063
rect 10794 7038 11210 7043
rect 11416 7041 11453 7070
rect 11417 7039 11453 7041
rect 11629 7039 11666 7070
rect 10794 7037 11135 7038
rect 10738 6977 10769 6978
rect 10586 6947 10595 6967
rect 10615 6947 10623 6967
rect 10586 6937 10623 6947
rect 10682 6970 10769 6977
rect 10682 6967 10743 6970
rect 10682 6947 10691 6967
rect 10711 6950 10743 6967
rect 10764 6950 10769 6970
rect 10711 6947 10769 6950
rect 10682 6940 10769 6947
rect 10794 6967 10831 7037
rect 11097 7036 11134 7037
rect 11417 7017 11666 7039
rect 11837 7038 11874 7070
rect 12150 7066 12214 7078
rect 12254 7042 12281 7218
rect 12712 7185 12739 7355
rect 12779 7325 12843 7337
rect 13119 7333 13156 7365
rect 13327 7364 13576 7386
rect 13859 7366 13896 7367
rect 14162 7366 14199 7436
rect 14224 7456 14311 7463
rect 14224 7453 14282 7456
rect 14224 7433 14229 7453
rect 14250 7436 14282 7453
rect 14302 7436 14311 7456
rect 14250 7433 14311 7436
rect 14224 7426 14311 7433
rect 14370 7456 14407 7466
rect 14370 7436 14378 7456
rect 14398 7436 14407 7456
rect 14224 7425 14255 7426
rect 13858 7365 14199 7366
rect 13327 7333 13364 7364
rect 13540 7362 13576 7364
rect 13540 7333 13577 7362
rect 13783 7360 14199 7365
rect 13783 7340 13786 7360
rect 13806 7340 14199 7360
rect 14370 7357 14407 7436
rect 14437 7465 14468 7518
rect 14818 7516 14855 7517
rect 14817 7507 14856 7516
rect 14817 7489 14827 7507
rect 14845 7489 14856 7507
rect 15197 7505 15234 7509
rect 14729 7472 14776 7473
rect 14817 7472 14856 7489
rect 14729 7468 14856 7472
rect 14487 7465 14524 7466
rect 14437 7456 14524 7465
rect 14437 7436 14495 7456
rect 14515 7436 14524 7456
rect 14437 7426 14524 7436
rect 14583 7456 14620 7466
rect 14583 7436 14591 7456
rect 14611 7436 14620 7456
rect 14437 7425 14468 7426
rect 14432 7357 14542 7370
rect 14583 7357 14620 7436
rect 14729 7439 14739 7468
rect 14768 7439 14856 7468
rect 14729 7433 14856 7439
rect 14729 7429 14776 7433
rect 14814 7419 14856 7433
rect 14814 7401 14825 7419
rect 14843 7401 14856 7419
rect 14814 7396 14856 7401
rect 14815 7393 14856 7396
rect 15194 7500 15234 7505
rect 15194 7482 15206 7500
rect 15224 7482 15234 7500
rect 14815 7392 14852 7393
rect 14370 7355 14620 7357
rect 14370 7352 14471 7355
rect 14370 7333 14435 7352
rect 12779 7324 12814 7325
rect 12756 7319 12814 7324
rect 12756 7299 12759 7319
rect 12779 7305 12814 7319
rect 12834 7305 12843 7325
rect 12779 7297 12843 7305
rect 12805 7296 12843 7297
rect 12806 7295 12843 7296
rect 12909 7329 12945 7330
rect 13017 7329 13053 7330
rect 12909 7321 13053 7329
rect 12909 7301 12917 7321
rect 12937 7301 13025 7321
rect 13045 7301 13053 7321
rect 12909 7295 13053 7301
rect 13119 7325 13157 7333
rect 13225 7329 13261 7330
rect 13119 7305 13128 7325
rect 13148 7305 13157 7325
rect 13119 7296 13157 7305
rect 13176 7322 13261 7329
rect 13176 7302 13183 7322
rect 13204 7321 13261 7322
rect 13204 7302 13233 7321
rect 13176 7301 13233 7302
rect 13253 7301 13261 7321
rect 13119 7295 13156 7296
rect 13176 7295 13261 7301
rect 13327 7325 13365 7333
rect 13438 7329 13474 7330
rect 13327 7305 13336 7325
rect 13356 7305 13365 7325
rect 13327 7296 13365 7305
rect 13389 7321 13474 7329
rect 13389 7301 13446 7321
rect 13466 7301 13474 7321
rect 13327 7295 13364 7296
rect 13389 7295 13474 7301
rect 13540 7325 13578 7333
rect 13540 7305 13549 7325
rect 13569 7305 13578 7325
rect 14432 7325 14435 7333
rect 14464 7325 14471 7352
rect 14499 7328 14509 7355
rect 14538 7333 14620 7355
rect 14538 7328 14542 7333
rect 14499 7325 14542 7328
rect 14432 7311 14542 7325
rect 14808 7329 14855 7330
rect 14808 7320 14856 7329
rect 13540 7296 13578 7305
rect 14808 7302 14827 7320
rect 14845 7302 14856 7320
rect 14808 7300 14856 7302
rect 13540 7295 13577 7296
rect 12963 7274 12999 7295
rect 13389 7274 13420 7295
rect 12796 7270 12896 7274
rect 12796 7266 12858 7270
rect 12796 7240 12803 7266
rect 12829 7244 12858 7266
rect 12884 7244 12896 7270
rect 12829 7240 12896 7244
rect 12796 7237 12896 7240
rect 12964 7237 12999 7274
rect 13061 7271 13420 7274
rect 13061 7266 13283 7271
rect 13061 7242 13074 7266
rect 13098 7247 13283 7266
rect 13307 7247 13420 7271
rect 13098 7242 13420 7247
rect 13061 7238 13420 7242
rect 13487 7266 13636 7274
rect 13487 7246 13498 7266
rect 13518 7246 13636 7266
rect 13487 7239 13636 7246
rect 14169 7243 14207 7245
rect 14817 7243 14856 7300
rect 15194 7302 15234 7482
rect 15580 7475 15611 7528
rect 15641 7557 15678 7636
rect 15849 7633 16242 7653
rect 16262 7633 16265 7653
rect 16363 7637 16612 7659
rect 16781 7658 16822 7663
rect 17200 7660 17227 7838
rect 17878 7750 17905 7928
rect 18283 7925 18324 7930
rect 18493 7929 18742 7951
rect 18840 7935 18843 7955
rect 18863 7935 19256 7955
rect 19427 7952 19464 8031
rect 19494 8060 19525 8113
rect 19871 8106 19911 8286
rect 19871 8088 19881 8106
rect 19899 8088 19911 8106
rect 19871 8083 19911 8088
rect 19871 8079 19908 8083
rect 19544 8060 19581 8061
rect 19494 8051 19581 8060
rect 19494 8031 19552 8051
rect 19572 8031 19581 8051
rect 19494 8021 19581 8031
rect 19640 8051 19677 8061
rect 19640 8031 19648 8051
rect 19668 8031 19677 8051
rect 19494 8020 19525 8021
rect 19489 7952 19599 7965
rect 19640 7952 19677 8031
rect 19874 8016 19911 8017
rect 19870 8007 19911 8016
rect 19870 7989 19883 8007
rect 19901 7989 19911 8007
rect 19870 7980 19911 7989
rect 19870 7960 19910 7980
rect 19427 7950 19677 7952
rect 19427 7947 19528 7950
rect 17945 7890 18009 7902
rect 18285 7898 18322 7925
rect 18493 7898 18530 7929
rect 18706 7927 18742 7929
rect 19427 7928 19492 7947
rect 18706 7898 18743 7927
rect 19489 7920 19492 7928
rect 19521 7920 19528 7947
rect 19556 7923 19566 7950
rect 19595 7928 19677 7950
rect 19785 7950 19910 7960
rect 19785 7931 19793 7950
rect 19818 7931 19910 7950
rect 19595 7923 19599 7928
rect 19785 7924 19910 7931
rect 19556 7920 19599 7923
rect 19489 7906 19599 7920
rect 17945 7889 17980 7890
rect 17922 7884 17980 7889
rect 17922 7864 17925 7884
rect 17945 7870 17980 7884
rect 18000 7870 18009 7890
rect 17945 7862 18009 7870
rect 17971 7861 18009 7862
rect 17972 7860 18009 7861
rect 18075 7894 18111 7895
rect 18183 7894 18219 7895
rect 18075 7886 18219 7894
rect 18075 7866 18083 7886
rect 18103 7883 18191 7886
rect 18103 7866 18135 7883
rect 18155 7866 18191 7883
rect 18211 7866 18219 7886
rect 18075 7860 18219 7866
rect 18285 7890 18323 7898
rect 18391 7894 18427 7895
rect 18285 7870 18294 7890
rect 18314 7870 18323 7890
rect 18285 7861 18323 7870
rect 18342 7887 18427 7894
rect 18342 7867 18349 7887
rect 18370 7886 18427 7887
rect 18370 7867 18399 7886
rect 18342 7866 18399 7867
rect 18419 7866 18427 7886
rect 18285 7860 18322 7861
rect 18342 7860 18427 7866
rect 18493 7890 18531 7898
rect 18604 7894 18640 7895
rect 18493 7870 18502 7890
rect 18522 7870 18531 7890
rect 18493 7861 18531 7870
rect 18555 7886 18640 7894
rect 18555 7866 18612 7886
rect 18632 7866 18640 7886
rect 18493 7860 18530 7861
rect 18555 7860 18640 7866
rect 18706 7890 18744 7898
rect 18706 7870 18715 7890
rect 18735 7870 18744 7890
rect 18706 7861 18744 7870
rect 19870 7876 19910 7924
rect 18706 7860 18743 7861
rect 18129 7839 18165 7860
rect 18555 7839 18586 7860
rect 19870 7858 19881 7876
rect 19899 7858 19910 7876
rect 19870 7850 19910 7858
rect 19871 7849 19908 7850
rect 17962 7835 18062 7839
rect 17962 7831 18024 7835
rect 17962 7805 17969 7831
rect 17995 7809 18024 7831
rect 18050 7809 18062 7835
rect 17995 7805 18062 7809
rect 17962 7802 18062 7805
rect 18130 7802 18165 7839
rect 18227 7836 18586 7839
rect 18227 7831 18449 7836
rect 18227 7807 18240 7831
rect 18264 7812 18449 7831
rect 18473 7812 18586 7836
rect 18264 7807 18586 7812
rect 18227 7803 18586 7807
rect 18653 7831 18802 7839
rect 18653 7811 18664 7831
rect 18684 7811 18802 7831
rect 18653 7804 18802 7811
rect 19242 7808 19756 7809
rect 18653 7803 18694 7804
rect 17977 7750 18014 7751
rect 18073 7750 18110 7751
rect 18129 7750 18165 7802
rect 18184 7750 18221 7751
rect 17877 7741 18015 7750
rect 17877 7721 17986 7741
rect 18006 7721 18015 7741
rect 17877 7714 18015 7721
rect 18073 7741 18221 7750
rect 18073 7721 18082 7741
rect 18102 7721 18192 7741
rect 18212 7721 18221 7741
rect 17877 7712 17973 7714
rect 18073 7711 18221 7721
rect 18280 7741 18317 7751
rect 18392 7750 18429 7751
rect 18373 7748 18429 7750
rect 18280 7721 18288 7741
rect 18308 7721 18317 7741
rect 18129 7710 18165 7711
rect 17059 7658 17227 7660
rect 16781 7652 17227 7658
rect 15849 7628 16265 7633
rect 16444 7631 16555 7637
rect 15849 7627 16190 7628
rect 15793 7567 15824 7568
rect 15641 7537 15650 7557
rect 15670 7537 15678 7557
rect 15641 7527 15678 7537
rect 15737 7560 15824 7567
rect 15737 7557 15798 7560
rect 15737 7537 15746 7557
rect 15766 7540 15798 7557
rect 15819 7540 15824 7560
rect 15766 7537 15824 7540
rect 15737 7530 15824 7537
rect 15849 7557 15886 7627
rect 16152 7626 16189 7627
rect 16444 7623 16485 7631
rect 16444 7603 16452 7623
rect 16471 7603 16485 7623
rect 16444 7601 16485 7603
rect 16513 7623 16555 7631
rect 16513 7603 16529 7623
rect 16548 7603 16555 7623
rect 16781 7630 16787 7652
rect 16813 7632 17227 7652
rect 17977 7651 18014 7652
rect 18280 7651 18317 7721
rect 18342 7741 18429 7748
rect 18342 7738 18400 7741
rect 18342 7718 18347 7738
rect 18368 7721 18400 7738
rect 18420 7721 18429 7741
rect 18368 7718 18429 7721
rect 18342 7711 18429 7718
rect 18488 7741 18525 7751
rect 18488 7721 18496 7741
rect 18516 7721 18525 7741
rect 18342 7710 18373 7711
rect 17976 7650 18317 7651
rect 16813 7630 16822 7632
rect 17059 7631 17227 7632
rect 17901 7645 18317 7650
rect 16781 7621 16822 7630
rect 17901 7625 17904 7645
rect 17924 7625 18317 7645
rect 18488 7642 18525 7721
rect 18555 7750 18586 7803
rect 19223 7792 19756 7808
rect 19223 7781 19755 7792
rect 19874 7783 19911 7787
rect 18605 7750 18642 7751
rect 18555 7741 18642 7750
rect 18555 7721 18613 7741
rect 18633 7721 18642 7741
rect 18555 7711 18642 7721
rect 18701 7741 18738 7751
rect 18701 7721 18709 7741
rect 18729 7721 18738 7741
rect 18555 7710 18586 7711
rect 18550 7642 18660 7655
rect 18701 7642 18738 7721
rect 18488 7640 18738 7642
rect 18488 7637 18589 7640
rect 18488 7618 18553 7637
rect 16513 7601 16555 7603
rect 16444 7586 16555 7601
rect 18550 7610 18553 7618
rect 18582 7610 18589 7637
rect 18617 7613 18627 7640
rect 18656 7618 18738 7640
rect 18816 7712 18984 7713
rect 19223 7712 19261 7781
rect 18816 7692 19261 7712
rect 19488 7743 19599 7758
rect 19488 7741 19530 7743
rect 19488 7721 19495 7741
rect 19514 7721 19530 7741
rect 19488 7713 19530 7721
rect 19558 7741 19599 7743
rect 19558 7721 19572 7741
rect 19591 7721 19599 7741
rect 19558 7713 19599 7721
rect 19488 7707 19599 7713
rect 19721 7718 19755 7781
rect 19873 7777 19911 7783
rect 19873 7759 19883 7777
rect 19901 7759 19911 7777
rect 19873 7750 19911 7759
rect 19873 7718 19907 7750
rect 18816 7686 19260 7692
rect 18816 7684 18984 7686
rect 18656 7613 18660 7618
rect 18617 7610 18660 7613
rect 18550 7596 18660 7610
rect 16001 7567 16037 7568
rect 15849 7537 15858 7557
rect 15878 7537 15886 7557
rect 15737 7528 15793 7530
rect 15737 7527 15774 7528
rect 15849 7527 15886 7537
rect 15945 7557 16093 7567
rect 16193 7564 16289 7566
rect 15945 7537 15954 7557
rect 15974 7537 16064 7557
rect 16084 7537 16093 7557
rect 15945 7528 16093 7537
rect 16151 7557 16289 7564
rect 16151 7537 16160 7557
rect 16180 7537 16289 7557
rect 16151 7528 16289 7537
rect 15945 7527 15982 7528
rect 16001 7476 16037 7528
rect 16056 7527 16093 7528
rect 16152 7527 16189 7528
rect 15472 7474 15513 7475
rect 15364 7467 15513 7474
rect 15364 7447 15482 7467
rect 15502 7447 15513 7467
rect 15364 7439 15513 7447
rect 15580 7471 15939 7475
rect 15580 7466 15902 7471
rect 15580 7442 15693 7466
rect 15717 7447 15902 7466
rect 15926 7447 15939 7471
rect 15717 7442 15939 7447
rect 15580 7439 15939 7442
rect 16001 7439 16036 7476
rect 16104 7473 16204 7476
rect 16104 7469 16171 7473
rect 16104 7443 16116 7469
rect 16142 7447 16171 7469
rect 16197 7447 16204 7473
rect 16142 7443 16204 7447
rect 16104 7439 16204 7443
rect 15580 7418 15611 7439
rect 16001 7418 16037 7439
rect 15423 7417 15460 7418
rect 15422 7408 15460 7417
rect 15422 7388 15431 7408
rect 15451 7388 15460 7408
rect 15422 7380 15460 7388
rect 15526 7412 15611 7418
rect 15636 7417 15673 7418
rect 15526 7392 15534 7412
rect 15554 7392 15611 7412
rect 15526 7384 15611 7392
rect 15635 7408 15673 7417
rect 15635 7388 15644 7408
rect 15664 7388 15673 7408
rect 15526 7383 15562 7384
rect 15635 7380 15673 7388
rect 15739 7412 15824 7418
rect 15844 7417 15881 7418
rect 15739 7392 15747 7412
rect 15767 7411 15824 7412
rect 15767 7392 15796 7411
rect 15739 7391 15796 7392
rect 15817 7391 15824 7411
rect 15739 7384 15824 7391
rect 15843 7408 15881 7417
rect 15843 7388 15852 7408
rect 15872 7388 15881 7408
rect 15739 7383 15775 7384
rect 15843 7380 15881 7388
rect 15947 7412 16091 7418
rect 15947 7392 15955 7412
rect 15975 7409 16063 7412
rect 15975 7392 16006 7409
rect 15947 7389 16006 7392
rect 16029 7392 16063 7409
rect 16083 7392 16091 7412
rect 16029 7389 16091 7392
rect 15947 7384 16091 7389
rect 15947 7383 15983 7384
rect 16055 7383 16091 7384
rect 16157 7417 16194 7418
rect 16157 7416 16195 7417
rect 16157 7408 16221 7416
rect 16157 7388 16166 7408
rect 16186 7394 16221 7408
rect 16241 7394 16244 7414
rect 16186 7389 16244 7394
rect 16186 7388 16221 7389
rect 15423 7351 15460 7380
rect 15424 7349 15460 7351
rect 15636 7349 15673 7380
rect 15424 7327 15673 7349
rect 15844 7348 15881 7380
rect 16157 7376 16221 7388
rect 16261 7350 16288 7528
rect 18816 7506 18843 7684
rect 18883 7646 18947 7658
rect 19223 7654 19260 7686
rect 19431 7685 19680 7707
rect 19721 7686 19907 7718
rect 19735 7685 19907 7686
rect 19431 7654 19468 7685
rect 19644 7683 19680 7685
rect 19644 7654 19681 7683
rect 19873 7657 19907 7685
rect 18883 7645 18918 7646
rect 18860 7640 18918 7645
rect 18860 7620 18863 7640
rect 18883 7626 18918 7640
rect 18938 7626 18947 7646
rect 18883 7618 18947 7626
rect 18909 7617 18947 7618
rect 18910 7616 18947 7617
rect 19013 7650 19049 7651
rect 19121 7650 19157 7651
rect 19013 7643 19157 7650
rect 19013 7642 19073 7643
rect 19013 7622 19021 7642
rect 19041 7623 19073 7642
rect 19098 7642 19157 7643
rect 19098 7623 19129 7642
rect 19041 7622 19129 7623
rect 19149 7622 19157 7642
rect 19013 7616 19157 7622
rect 19223 7646 19261 7654
rect 19329 7650 19365 7651
rect 19223 7626 19232 7646
rect 19252 7626 19261 7646
rect 19223 7617 19261 7626
rect 19280 7643 19365 7650
rect 19280 7623 19287 7643
rect 19308 7642 19365 7643
rect 19308 7623 19337 7642
rect 19280 7622 19337 7623
rect 19357 7622 19365 7642
rect 19223 7616 19260 7617
rect 19280 7616 19365 7622
rect 19431 7646 19469 7654
rect 19542 7650 19578 7651
rect 19431 7626 19440 7646
rect 19460 7626 19469 7646
rect 19431 7617 19469 7626
rect 19493 7642 19578 7650
rect 19493 7622 19550 7642
rect 19570 7622 19578 7642
rect 19431 7616 19468 7617
rect 19493 7616 19578 7622
rect 19644 7646 19682 7654
rect 19644 7626 19653 7646
rect 19673 7626 19682 7646
rect 19644 7617 19682 7626
rect 19871 7647 19908 7657
rect 19871 7629 19881 7647
rect 19899 7629 19908 7647
rect 19871 7620 19908 7629
rect 19873 7619 19907 7620
rect 19644 7616 19681 7617
rect 19067 7595 19103 7616
rect 19493 7595 19524 7616
rect 18900 7591 19000 7595
rect 18900 7587 18962 7591
rect 18900 7561 18907 7587
rect 18933 7565 18962 7587
rect 18988 7565 19000 7591
rect 18933 7561 19000 7565
rect 18900 7558 19000 7561
rect 19068 7558 19103 7595
rect 19165 7592 19524 7595
rect 19165 7587 19387 7592
rect 19165 7563 19178 7587
rect 19202 7568 19387 7587
rect 19411 7568 19524 7592
rect 19202 7563 19524 7568
rect 19165 7559 19524 7563
rect 19591 7587 19740 7595
rect 19591 7567 19602 7587
rect 19622 7567 19740 7587
rect 19591 7560 19740 7567
rect 19591 7559 19632 7560
rect 18915 7506 18952 7507
rect 19011 7506 19048 7507
rect 19067 7506 19103 7558
rect 19122 7506 19159 7507
rect 18815 7497 18953 7506
rect 18440 7463 18551 7478
rect 18815 7477 18924 7497
rect 18944 7477 18953 7497
rect 18815 7470 18953 7477
rect 19011 7497 19159 7506
rect 19011 7477 19020 7497
rect 19040 7477 19130 7497
rect 19150 7477 19159 7497
rect 18815 7468 18911 7470
rect 19011 7467 19159 7477
rect 19218 7497 19255 7507
rect 19330 7506 19367 7507
rect 19311 7504 19367 7506
rect 19218 7477 19226 7497
rect 19246 7477 19255 7497
rect 19067 7466 19103 7467
rect 18440 7461 18482 7463
rect 17777 7442 17847 7451
rect 17777 7433 17794 7442
rect 17768 7413 17794 7433
rect 17842 7433 17847 7442
rect 18440 7441 18447 7461
rect 18466 7441 18482 7461
rect 18440 7433 18482 7441
rect 18510 7461 18551 7463
rect 18510 7441 18524 7461
rect 18543 7441 18551 7461
rect 18510 7433 18551 7441
rect 17842 7432 17936 7433
rect 17842 7413 18212 7432
rect 18440 7427 18551 7433
rect 16555 7399 16665 7413
rect 16555 7396 16598 7399
rect 16555 7391 16559 7396
rect 16120 7348 16288 7350
rect 15844 7345 16288 7348
rect 15505 7321 15616 7327
rect 15505 7313 15546 7321
rect 15194 7258 15233 7302
rect 15505 7293 15513 7313
rect 15532 7293 15546 7313
rect 15505 7291 15546 7293
rect 15574 7313 15616 7321
rect 15574 7293 15590 7313
rect 15609 7293 15616 7313
rect 15574 7291 15616 7293
rect 15505 7277 15616 7291
rect 15842 7322 16288 7345
rect 13487 7238 13528 7239
rect 12963 7197 12999 7237
rect 12811 7185 12848 7186
rect 12907 7185 12944 7186
rect 12963 7185 12968 7197
rect 12711 7176 12849 7185
rect 12711 7156 12820 7176
rect 12840 7156 12849 7176
rect 12711 7149 12849 7156
rect 12907 7176 12968 7185
rect 12907 7156 12916 7176
rect 12936 7165 12968 7176
rect 12995 7185 12999 7197
rect 13018 7185 13055 7186
rect 12995 7176 13055 7185
rect 12995 7165 13026 7176
rect 12936 7156 13026 7165
rect 13046 7156 13055 7176
rect 12711 7147 12807 7149
rect 12907 7146 13055 7156
rect 13114 7176 13151 7186
rect 13226 7185 13263 7186
rect 13207 7183 13263 7185
rect 13114 7156 13122 7176
rect 13142 7156 13151 7176
rect 12963 7145 12999 7146
rect 12811 7086 12848 7087
rect 13114 7086 13151 7156
rect 13176 7176 13263 7183
rect 13176 7173 13234 7176
rect 13176 7153 13181 7173
rect 13202 7156 13234 7173
rect 13254 7156 13263 7176
rect 13202 7153 13263 7156
rect 13176 7146 13263 7153
rect 13322 7176 13359 7186
rect 13322 7156 13330 7176
rect 13350 7156 13359 7176
rect 13176 7145 13207 7146
rect 12810 7085 13151 7086
rect 12735 7080 13151 7085
rect 12735 7062 12738 7080
rect 12758 7078 13151 7080
rect 12758 7062 13128 7078
rect 12776 7060 13128 7062
rect 13119 7058 13128 7060
rect 13149 7058 13151 7078
rect 13119 7046 13151 7058
rect 13322 7077 13359 7156
rect 13389 7185 13420 7238
rect 14169 7210 14855 7243
rect 13439 7185 13476 7186
rect 13389 7176 13476 7185
rect 13389 7156 13447 7176
rect 13467 7156 13476 7176
rect 13389 7146 13476 7156
rect 13535 7176 13572 7186
rect 13535 7156 13543 7176
rect 13563 7156 13572 7176
rect 13389 7145 13420 7146
rect 13384 7077 13494 7090
rect 13535 7077 13572 7156
rect 13322 7075 13572 7077
rect 13322 7072 13423 7075
rect 13322 7053 13387 7072
rect 12162 7040 12281 7042
rect 12113 7038 12281 7040
rect 11498 7011 11609 7017
rect 11837 7012 12281 7038
rect 13384 7045 13387 7053
rect 13416 7045 13423 7072
rect 13451 7048 13461 7075
rect 13490 7053 13572 7075
rect 13761 7122 13929 7123
rect 14169 7122 14207 7210
rect 14468 7208 14515 7210
rect 14815 7186 14855 7210
rect 15194 7234 15234 7258
rect 15534 7234 15581 7236
rect 15842 7234 15880 7322
rect 16120 7321 16288 7322
rect 16477 7369 16559 7391
rect 16588 7369 16598 7396
rect 16626 7372 16633 7399
rect 16662 7391 16665 7399
rect 17768 7406 18212 7413
rect 17768 7404 17936 7406
rect 17768 7396 17847 7404
rect 16662 7372 16727 7391
rect 16626 7369 16727 7372
rect 16477 7367 16727 7369
rect 16477 7288 16514 7367
rect 16555 7354 16665 7367
rect 16629 7298 16660 7299
rect 16477 7268 16486 7288
rect 16506 7268 16514 7288
rect 16477 7258 16514 7268
rect 16573 7288 16660 7298
rect 16573 7268 16582 7288
rect 16602 7268 16660 7288
rect 16573 7259 16660 7268
rect 16573 7258 16610 7259
rect 15194 7201 15880 7234
rect 16629 7206 16660 7259
rect 16690 7288 16727 7367
rect 16898 7364 17291 7384
rect 17311 7364 17314 7384
rect 16898 7359 17314 7364
rect 16898 7358 17239 7359
rect 16842 7298 16873 7299
rect 16690 7268 16699 7288
rect 16719 7268 16727 7288
rect 16690 7258 16727 7268
rect 16786 7291 16873 7298
rect 16786 7288 16847 7291
rect 16786 7268 16795 7288
rect 16815 7271 16847 7288
rect 16868 7271 16873 7291
rect 16815 7268 16873 7271
rect 16786 7261 16873 7268
rect 16898 7288 16935 7358
rect 17201 7357 17238 7358
rect 17050 7298 17086 7299
rect 16898 7268 16907 7288
rect 16927 7268 16935 7288
rect 16786 7259 16842 7261
rect 16786 7258 16823 7259
rect 16898 7258 16935 7268
rect 16994 7288 17142 7298
rect 17242 7295 17338 7297
rect 16994 7268 17003 7288
rect 17023 7268 17113 7288
rect 17133 7268 17142 7288
rect 16994 7259 17142 7268
rect 17200 7288 17338 7295
rect 17200 7268 17209 7288
rect 17229 7268 17338 7288
rect 17200 7259 17338 7268
rect 16994 7258 17031 7259
rect 17050 7207 17086 7259
rect 17105 7258 17142 7259
rect 17201 7258 17238 7259
rect 16521 7205 16562 7206
rect 13761 7099 14207 7122
rect 14433 7153 14544 7167
rect 14433 7151 14475 7153
rect 14433 7131 14440 7151
rect 14459 7131 14475 7151
rect 14433 7123 14475 7131
rect 14503 7151 14544 7153
rect 14503 7131 14517 7151
rect 14536 7131 14544 7151
rect 14816 7142 14855 7186
rect 14503 7123 14544 7131
rect 14433 7117 14544 7123
rect 13761 7096 14205 7099
rect 13761 7094 13929 7096
rect 13490 7048 13494 7053
rect 13451 7045 13494 7048
rect 13384 7031 13494 7045
rect 12113 7011 12281 7012
rect 11498 7003 11539 7011
rect 11498 6983 11506 7003
rect 11525 6983 11539 7003
rect 11498 6981 11539 6983
rect 11567 7003 11609 7011
rect 12162 7010 12270 7011
rect 11567 6983 11583 7003
rect 11602 6983 11609 7003
rect 11567 6981 11609 6983
rect 10946 6977 10982 6978
rect 10794 6947 10803 6967
rect 10823 6947 10831 6967
rect 10682 6938 10738 6940
rect 10682 6937 10719 6938
rect 10794 6937 10831 6947
rect 10890 6967 11038 6977
rect 11138 6974 11234 6976
rect 10890 6947 10899 6967
rect 10919 6947 11009 6967
rect 11029 6947 11038 6967
rect 10890 6938 11038 6947
rect 11096 6967 11234 6974
rect 11096 6947 11105 6967
rect 11125 6947 11234 6967
rect 11498 6966 11609 6981
rect 12200 7009 12270 7010
rect 11096 6938 11234 6947
rect 10890 6937 10927 6938
rect 10946 6886 10982 6938
rect 11001 6937 11038 6938
rect 11097 6937 11134 6938
rect 10417 6884 10458 6885
rect 9839 6872 9880 6881
rect 10309 6877 10458 6884
rect 9839 6852 9879 6872
rect 9396 6842 9646 6844
rect 9396 6839 9497 6842
rect 7914 6782 7978 6794
rect 8254 6790 8291 6817
rect 8462 6790 8499 6821
rect 8675 6819 8711 6821
rect 9396 6820 9461 6839
rect 8675 6790 8712 6819
rect 9458 6812 9461 6820
rect 9490 6812 9497 6839
rect 9525 6815 9535 6842
rect 9564 6820 9646 6842
rect 9754 6842 9879 6852
rect 10309 6857 10427 6877
rect 10447 6857 10458 6877
rect 10309 6849 10458 6857
rect 10525 6881 10884 6885
rect 10525 6876 10847 6881
rect 10525 6852 10638 6876
rect 10662 6857 10847 6876
rect 10871 6857 10884 6881
rect 10662 6852 10884 6857
rect 10525 6849 10884 6852
rect 10946 6849 10981 6886
rect 11049 6883 11149 6886
rect 11049 6879 11116 6883
rect 11049 6853 11061 6879
rect 11087 6857 11116 6879
rect 11142 6857 11149 6883
rect 11087 6853 11149 6857
rect 11049 6849 11149 6853
rect 9754 6823 9762 6842
rect 9787 6823 9879 6842
rect 10525 6828 10556 6849
rect 10946 6828 10982 6849
rect 10368 6827 10405 6828
rect 10142 6824 10176 6825
rect 9564 6815 9568 6820
rect 9754 6816 9879 6823
rect 9525 6812 9568 6815
rect 9458 6798 9568 6812
rect 7914 6781 7949 6782
rect 7891 6776 7949 6781
rect 7891 6756 7894 6776
rect 7914 6762 7949 6776
rect 7969 6762 7978 6782
rect 7914 6754 7978 6762
rect 7940 6753 7978 6754
rect 7941 6752 7978 6753
rect 8044 6786 8080 6787
rect 8152 6786 8188 6787
rect 8044 6778 8188 6786
rect 8044 6758 8052 6778
rect 8072 6758 8160 6778
rect 8180 6758 8188 6778
rect 8044 6752 8188 6758
rect 8254 6782 8292 6790
rect 8360 6786 8396 6787
rect 8254 6762 8263 6782
rect 8283 6762 8292 6782
rect 8254 6753 8292 6762
rect 8311 6779 8396 6786
rect 8311 6759 8318 6779
rect 8339 6778 8396 6779
rect 8339 6759 8368 6778
rect 8311 6758 8368 6759
rect 8388 6758 8396 6778
rect 8254 6752 8291 6753
rect 8311 6752 8396 6758
rect 8462 6782 8500 6790
rect 8573 6786 8609 6787
rect 8462 6762 8471 6782
rect 8491 6762 8500 6782
rect 8462 6753 8500 6762
rect 8524 6778 8609 6786
rect 8524 6758 8581 6778
rect 8601 6758 8609 6778
rect 8462 6752 8499 6753
rect 8524 6752 8609 6758
rect 8675 6782 8713 6790
rect 8675 6762 8684 6782
rect 8704 6762 8713 6782
rect 8675 6753 8713 6762
rect 9839 6768 9879 6816
rect 10141 6815 10178 6824
rect 10141 6797 10150 6815
rect 10168 6797 10178 6815
rect 10141 6787 10178 6797
rect 10367 6818 10405 6827
rect 10367 6798 10376 6818
rect 10396 6798 10405 6818
rect 10367 6790 10405 6798
rect 10471 6822 10556 6828
rect 10581 6827 10618 6828
rect 10471 6802 10479 6822
rect 10499 6802 10556 6822
rect 10471 6794 10556 6802
rect 10580 6818 10618 6827
rect 10580 6798 10589 6818
rect 10609 6798 10618 6818
rect 10471 6793 10507 6794
rect 10580 6790 10618 6798
rect 10684 6822 10769 6828
rect 10789 6827 10826 6828
rect 10684 6802 10692 6822
rect 10712 6821 10769 6822
rect 10712 6802 10741 6821
rect 10684 6801 10741 6802
rect 10762 6801 10769 6821
rect 10684 6794 10769 6801
rect 10788 6818 10826 6827
rect 10788 6798 10797 6818
rect 10817 6798 10826 6818
rect 10684 6793 10720 6794
rect 10788 6790 10826 6798
rect 10892 6822 11036 6828
rect 10892 6802 10900 6822
rect 10920 6821 11008 6822
rect 10920 6802 10951 6821
rect 10892 6801 10951 6802
rect 10976 6802 11008 6821
rect 11028 6802 11036 6822
rect 10976 6801 11036 6802
rect 10892 6794 11036 6801
rect 10892 6793 10928 6794
rect 11000 6793 11036 6794
rect 11102 6827 11139 6828
rect 11102 6826 11140 6827
rect 11102 6818 11166 6826
rect 11102 6798 11111 6818
rect 11131 6804 11166 6818
rect 11186 6804 11189 6824
rect 11131 6799 11189 6804
rect 11131 6798 11166 6799
rect 8675 6752 8712 6753
rect 8098 6731 8134 6752
rect 8524 6731 8555 6752
rect 9839 6750 9850 6768
rect 9868 6750 9879 6768
rect 9839 6742 9879 6750
rect 10142 6759 10176 6787
rect 10368 6761 10405 6790
rect 10369 6759 10405 6761
rect 10581 6759 10618 6790
rect 10142 6758 10314 6759
rect 9840 6741 9877 6742
rect 7931 6727 8031 6731
rect 7931 6723 7993 6727
rect 7931 6697 7938 6723
rect 7964 6701 7993 6723
rect 8019 6701 8031 6727
rect 7964 6697 8031 6701
rect 7931 6694 8031 6697
rect 8099 6694 8134 6731
rect 8196 6728 8555 6731
rect 8196 6723 8418 6728
rect 8196 6699 8209 6723
rect 8233 6704 8418 6723
rect 8442 6704 8555 6728
rect 8233 6699 8555 6704
rect 8196 6695 8555 6699
rect 8622 6723 8771 6731
rect 8622 6703 8633 6723
rect 8653 6703 8771 6723
rect 8622 6696 8771 6703
rect 10142 6726 10328 6758
rect 10369 6737 10618 6759
rect 10789 6758 10826 6790
rect 11102 6786 11166 6798
rect 11206 6760 11233 6938
rect 12200 6902 12261 7009
rect 13761 6916 13788 7094
rect 13828 7056 13892 7068
rect 14168 7064 14205 7096
rect 14376 7095 14625 7117
rect 14376 7064 14413 7095
rect 14589 7093 14625 7095
rect 14589 7064 14626 7093
rect 13828 7055 13863 7056
rect 13805 7050 13863 7055
rect 13805 7030 13808 7050
rect 13828 7036 13863 7050
rect 13883 7036 13892 7056
rect 13828 7028 13892 7036
rect 13854 7027 13892 7028
rect 13855 7026 13892 7027
rect 13958 7060 13994 7061
rect 14066 7060 14102 7061
rect 13958 7055 14102 7060
rect 13958 7052 14020 7055
rect 13958 7032 13966 7052
rect 13986 7035 14020 7052
rect 14043 7052 14102 7055
rect 14043 7035 14074 7052
rect 13986 7032 14074 7035
rect 14094 7032 14102 7052
rect 13958 7026 14102 7032
rect 14168 7056 14206 7064
rect 14274 7060 14310 7061
rect 14168 7036 14177 7056
rect 14197 7036 14206 7056
rect 14168 7027 14206 7036
rect 14225 7053 14310 7060
rect 14225 7033 14232 7053
rect 14253 7052 14310 7053
rect 14253 7033 14282 7052
rect 14225 7032 14282 7033
rect 14302 7032 14310 7052
rect 14168 7026 14205 7027
rect 14225 7026 14310 7032
rect 14376 7056 14414 7064
rect 14487 7060 14523 7061
rect 14376 7036 14385 7056
rect 14405 7036 14414 7056
rect 14376 7027 14414 7036
rect 14438 7052 14523 7060
rect 14438 7032 14495 7052
rect 14515 7032 14523 7052
rect 14376 7026 14413 7027
rect 14438 7026 14523 7032
rect 14589 7056 14627 7064
rect 14589 7036 14598 7056
rect 14618 7036 14627 7056
rect 14589 7027 14627 7036
rect 14589 7026 14626 7027
rect 14012 7005 14048 7026
rect 14438 7005 14469 7026
rect 13845 7001 13945 7005
rect 13845 6997 13907 7001
rect 13845 6971 13852 6997
rect 13878 6975 13907 6997
rect 13933 6975 13945 7001
rect 13878 6971 13945 6975
rect 13845 6968 13945 6971
rect 14013 6968 14048 7005
rect 14110 7002 14469 7005
rect 14110 6997 14332 7002
rect 14110 6973 14123 6997
rect 14147 6978 14332 6997
rect 14356 6978 14469 7002
rect 14147 6973 14469 6978
rect 14110 6969 14469 6973
rect 14536 6997 14685 7005
rect 14536 6977 14547 6997
rect 14567 6977 14685 6997
rect 14536 6970 14685 6977
rect 14536 6969 14577 6970
rect 13860 6916 13897 6917
rect 13956 6916 13993 6917
rect 14012 6916 14048 6968
rect 14067 6916 14104 6917
rect 13760 6907 13898 6916
rect 12200 6891 12270 6902
rect 12200 6882 12207 6891
rect 12202 6862 12207 6882
rect 12255 6862 12270 6891
rect 13760 6887 13869 6907
rect 13889 6887 13898 6907
rect 13760 6880 13898 6887
rect 13956 6907 14104 6916
rect 13956 6887 13965 6907
rect 13985 6887 14075 6907
rect 14095 6887 14104 6907
rect 13760 6878 13856 6880
rect 13956 6877 14104 6887
rect 14163 6907 14200 6917
rect 14275 6916 14312 6917
rect 14256 6914 14312 6916
rect 14163 6887 14171 6907
rect 14191 6887 14200 6907
rect 14012 6876 14048 6877
rect 12202 6853 12270 6862
rect 11389 6834 11499 6848
rect 11389 6831 11432 6834
rect 11389 6826 11393 6831
rect 11065 6758 11233 6760
rect 10789 6752 11233 6758
rect 9211 6700 9725 6701
rect 8622 6695 8663 6696
rect 8098 6659 8134 6694
rect 7946 6642 7983 6643
rect 8042 6642 8079 6643
rect 8098 6642 8105 6659
rect 7846 6633 7984 6642
rect 7846 6613 7955 6633
rect 7975 6613 7984 6633
rect 7846 6606 7984 6613
rect 8042 6633 8105 6642
rect 8042 6613 8051 6633
rect 8071 6618 8105 6633
rect 8126 6642 8134 6659
rect 8153 6642 8190 6643
rect 8126 6633 8190 6642
rect 8126 6618 8161 6633
rect 8071 6613 8161 6618
rect 8181 6613 8190 6633
rect 7846 6604 7942 6606
rect 8042 6603 8190 6613
rect 8249 6633 8286 6643
rect 8361 6642 8398 6643
rect 8342 6640 8398 6642
rect 8249 6613 8257 6633
rect 8277 6613 8286 6633
rect 8098 6602 8134 6603
rect 7028 6550 7196 6552
rect 6750 6544 7196 6550
rect 5818 6520 6234 6525
rect 6413 6523 6524 6529
rect 5818 6519 6159 6520
rect 5762 6459 5793 6460
rect 5610 6429 5619 6449
rect 5639 6429 5647 6449
rect 5610 6419 5647 6429
rect 5706 6452 5793 6459
rect 5706 6449 5767 6452
rect 5706 6429 5715 6449
rect 5735 6432 5767 6449
rect 5788 6432 5793 6452
rect 5735 6429 5793 6432
rect 5706 6422 5793 6429
rect 5818 6449 5855 6519
rect 6121 6518 6158 6519
rect 6413 6515 6454 6523
rect 6413 6495 6421 6515
rect 6440 6495 6454 6515
rect 6413 6493 6454 6495
rect 6482 6515 6524 6523
rect 6482 6495 6498 6515
rect 6517 6495 6524 6515
rect 6750 6522 6756 6544
rect 6782 6524 7196 6544
rect 7946 6543 7983 6544
rect 8249 6543 8286 6613
rect 8311 6633 8398 6640
rect 8311 6630 8369 6633
rect 8311 6610 8316 6630
rect 8337 6613 8369 6630
rect 8389 6613 8398 6633
rect 8337 6610 8398 6613
rect 8311 6603 8398 6610
rect 8457 6633 8494 6643
rect 8457 6613 8465 6633
rect 8485 6613 8494 6633
rect 8311 6602 8342 6603
rect 7945 6542 8286 6543
rect 6782 6522 6791 6524
rect 7028 6523 7196 6524
rect 7870 6541 8286 6542
rect 7870 6537 8246 6541
rect 6750 6513 6791 6522
rect 7870 6517 7873 6537
rect 7893 6524 8246 6537
rect 8278 6524 8286 6541
rect 7893 6517 8286 6524
rect 8457 6534 8494 6613
rect 8524 6642 8555 6695
rect 9192 6684 9725 6700
rect 10142 6694 10176 6726
rect 10138 6685 10176 6694
rect 9192 6673 9724 6684
rect 9843 6675 9880 6679
rect 8574 6642 8611 6643
rect 8524 6633 8611 6642
rect 8524 6613 8582 6633
rect 8602 6613 8611 6633
rect 8524 6603 8611 6613
rect 8670 6633 8707 6643
rect 8670 6613 8678 6633
rect 8698 6613 8707 6633
rect 8524 6602 8555 6603
rect 8519 6534 8629 6547
rect 8670 6534 8707 6613
rect 8457 6532 8707 6534
rect 8457 6529 8558 6532
rect 8457 6510 8522 6529
rect 6482 6493 6524 6495
rect 6413 6478 6524 6493
rect 8519 6502 8522 6510
rect 8551 6502 8558 6529
rect 8586 6505 8596 6532
rect 8625 6510 8707 6532
rect 8785 6604 8953 6605
rect 9192 6604 9230 6673
rect 8785 6584 9230 6604
rect 9457 6635 9568 6650
rect 9457 6633 9499 6635
rect 9457 6613 9464 6633
rect 9483 6613 9499 6633
rect 9457 6605 9499 6613
rect 9527 6633 9568 6635
rect 9527 6613 9541 6633
rect 9560 6613 9568 6633
rect 9527 6605 9568 6613
rect 9457 6599 9568 6605
rect 9690 6610 9724 6673
rect 9842 6669 9880 6675
rect 9842 6651 9852 6669
rect 9870 6651 9880 6669
rect 10138 6667 10148 6685
rect 10166 6667 10176 6685
rect 10138 6661 10176 6667
rect 10294 6663 10328 6726
rect 10450 6731 10561 6737
rect 10450 6723 10491 6731
rect 10450 6703 10458 6723
rect 10477 6703 10491 6723
rect 10450 6701 10491 6703
rect 10519 6723 10561 6731
rect 10519 6703 10535 6723
rect 10554 6703 10561 6723
rect 10519 6701 10561 6703
rect 10450 6686 10561 6701
rect 10788 6732 11233 6752
rect 10788 6663 10826 6732
rect 11065 6731 11233 6732
rect 11311 6804 11393 6826
rect 11422 6804 11432 6831
rect 11460 6807 11467 6834
rect 11496 6826 11499 6834
rect 13494 6843 13605 6858
rect 13494 6841 13536 6843
rect 11496 6807 11561 6826
rect 11460 6804 11561 6807
rect 11311 6802 11561 6804
rect 11311 6723 11348 6802
rect 11389 6789 11499 6802
rect 11463 6733 11494 6734
rect 11311 6703 11320 6723
rect 11340 6703 11348 6723
rect 11311 6693 11348 6703
rect 11407 6723 11494 6733
rect 11407 6703 11416 6723
rect 11436 6703 11494 6723
rect 11407 6694 11494 6703
rect 11407 6693 11444 6694
rect 10138 6657 10175 6661
rect 10294 6652 10826 6663
rect 9842 6642 9880 6651
rect 9842 6610 9876 6642
rect 10293 6636 10826 6652
rect 11463 6641 11494 6694
rect 11524 6723 11561 6802
rect 11732 6799 12125 6819
rect 12145 6799 12148 6819
rect 13227 6814 13268 6823
rect 11732 6794 12148 6799
rect 12822 6812 12990 6813
rect 13227 6812 13236 6814
rect 11732 6793 12073 6794
rect 11676 6733 11707 6734
rect 11524 6703 11533 6723
rect 11553 6703 11561 6723
rect 11524 6693 11561 6703
rect 11620 6726 11707 6733
rect 11620 6723 11681 6726
rect 11620 6703 11629 6723
rect 11649 6706 11681 6723
rect 11702 6706 11707 6726
rect 11649 6703 11707 6706
rect 11620 6696 11707 6703
rect 11732 6723 11769 6793
rect 12035 6792 12072 6793
rect 12822 6792 13236 6812
rect 13262 6792 13268 6814
rect 13494 6821 13501 6841
rect 13520 6821 13536 6841
rect 13494 6813 13536 6821
rect 13564 6841 13605 6843
rect 13564 6821 13578 6841
rect 13597 6821 13605 6841
rect 13564 6813 13605 6821
rect 13860 6817 13897 6818
rect 14163 6817 14200 6887
rect 14225 6907 14312 6914
rect 14225 6904 14283 6907
rect 14225 6884 14230 6904
rect 14251 6887 14283 6904
rect 14303 6887 14312 6907
rect 14251 6884 14312 6887
rect 14225 6877 14312 6884
rect 14371 6907 14408 6917
rect 14371 6887 14379 6907
rect 14399 6887 14408 6907
rect 14225 6876 14256 6877
rect 13859 6816 14200 6817
rect 13494 6807 13605 6813
rect 13784 6811 14200 6816
rect 12822 6786 13268 6792
rect 12822 6784 12990 6786
rect 11884 6733 11920 6734
rect 11732 6703 11741 6723
rect 11761 6703 11769 6723
rect 11620 6694 11676 6696
rect 11620 6693 11657 6694
rect 11732 6693 11769 6703
rect 11828 6723 11976 6733
rect 12076 6730 12172 6732
rect 11828 6703 11837 6723
rect 11857 6703 11947 6723
rect 11967 6703 11976 6723
rect 11828 6694 11976 6703
rect 12034 6723 12172 6730
rect 12034 6703 12043 6723
rect 12063 6703 12172 6723
rect 12034 6694 12172 6703
rect 11828 6693 11865 6694
rect 11884 6642 11920 6694
rect 11939 6693 11976 6694
rect 12035 6693 12072 6694
rect 11355 6640 11396 6641
rect 10293 6635 10807 6636
rect 8785 6578 9229 6584
rect 8785 6576 8953 6578
rect 8625 6505 8629 6510
rect 8586 6502 8629 6505
rect 8519 6488 8629 6502
rect 5970 6459 6006 6460
rect 5818 6429 5827 6449
rect 5847 6429 5855 6449
rect 5706 6420 5762 6422
rect 5706 6419 5743 6420
rect 5818 6419 5855 6429
rect 5914 6449 6062 6459
rect 6162 6456 6258 6458
rect 5914 6429 5923 6449
rect 5943 6429 6033 6449
rect 6053 6429 6062 6449
rect 5914 6420 6062 6429
rect 6120 6449 6258 6456
rect 6120 6429 6129 6449
rect 6149 6429 6258 6449
rect 6120 6420 6258 6429
rect 5914 6419 5951 6420
rect 5970 6368 6006 6420
rect 6025 6419 6062 6420
rect 6121 6419 6158 6420
rect 5441 6366 5482 6367
rect 5333 6359 5482 6366
rect 5333 6339 5451 6359
rect 5471 6339 5482 6359
rect 5333 6331 5482 6339
rect 5549 6363 5908 6367
rect 5549 6358 5871 6363
rect 5549 6334 5662 6358
rect 5686 6339 5871 6358
rect 5895 6339 5908 6363
rect 5686 6334 5908 6339
rect 5549 6331 5908 6334
rect 5970 6331 6005 6368
rect 6073 6365 6173 6368
rect 6073 6361 6140 6365
rect 6073 6335 6085 6361
rect 6111 6339 6140 6361
rect 6166 6339 6173 6365
rect 6111 6335 6173 6339
rect 6073 6331 6173 6335
rect 5549 6310 5580 6331
rect 5970 6310 6006 6331
rect 5392 6309 5429 6310
rect 5391 6300 5429 6309
rect 5391 6280 5400 6300
rect 5420 6280 5429 6300
rect 5391 6272 5429 6280
rect 5495 6304 5580 6310
rect 5605 6309 5642 6310
rect 5495 6284 5503 6304
rect 5523 6284 5580 6304
rect 5495 6276 5580 6284
rect 5604 6300 5642 6309
rect 5604 6280 5613 6300
rect 5633 6280 5642 6300
rect 5495 6275 5531 6276
rect 5604 6272 5642 6280
rect 5708 6304 5793 6310
rect 5813 6309 5850 6310
rect 5708 6284 5716 6304
rect 5736 6303 5793 6304
rect 5736 6284 5765 6303
rect 5708 6283 5765 6284
rect 5786 6283 5793 6303
rect 5708 6276 5793 6283
rect 5812 6300 5850 6309
rect 5812 6280 5821 6300
rect 5841 6280 5850 6300
rect 5708 6275 5744 6276
rect 5812 6272 5850 6280
rect 5916 6304 6060 6310
rect 5916 6284 5924 6304
rect 5944 6301 6032 6304
rect 5944 6284 5975 6301
rect 5916 6281 5975 6284
rect 5998 6284 6032 6301
rect 6052 6284 6060 6304
rect 5998 6281 6060 6284
rect 5916 6276 6060 6281
rect 5916 6275 5952 6276
rect 6024 6275 6060 6276
rect 6126 6309 6163 6310
rect 6126 6308 6164 6309
rect 6126 6300 6190 6308
rect 6126 6280 6135 6300
rect 6155 6286 6190 6300
rect 6210 6286 6213 6306
rect 6155 6281 6213 6286
rect 6155 6280 6190 6281
rect 5392 6243 5429 6272
rect 5393 6241 5429 6243
rect 5605 6241 5642 6272
rect 5393 6219 5642 6241
rect 5813 6240 5850 6272
rect 6126 6268 6190 6280
rect 6230 6242 6257 6420
rect 8785 6398 8812 6576
rect 8852 6538 8916 6550
rect 9192 6546 9229 6578
rect 9400 6577 9649 6599
rect 9690 6578 9876 6610
rect 11247 6633 11396 6640
rect 11247 6613 11365 6633
rect 11385 6613 11396 6633
rect 11247 6605 11396 6613
rect 11463 6637 11822 6641
rect 11463 6632 11785 6637
rect 11463 6608 11576 6632
rect 11600 6613 11785 6632
rect 11809 6613 11822 6637
rect 11600 6608 11822 6613
rect 11463 6605 11822 6608
rect 11884 6605 11919 6642
rect 11987 6639 12087 6642
rect 11987 6635 12054 6639
rect 11987 6609 11999 6635
rect 12025 6613 12054 6635
rect 12080 6613 12087 6639
rect 12025 6609 12087 6613
rect 11987 6605 12087 6609
rect 10141 6594 10178 6595
rect 9704 6577 9876 6578
rect 9400 6546 9437 6577
rect 9613 6575 9649 6577
rect 9613 6546 9650 6575
rect 9842 6549 9876 6577
rect 10139 6586 10179 6594
rect 10139 6568 10150 6586
rect 10168 6568 10179 6586
rect 11463 6584 11494 6605
rect 11884 6584 11920 6605
rect 11306 6583 11343 6584
rect 8852 6537 8887 6538
rect 8829 6532 8887 6537
rect 8829 6512 8832 6532
rect 8852 6518 8887 6532
rect 8907 6518 8916 6538
rect 8852 6510 8916 6518
rect 8878 6509 8916 6510
rect 8879 6508 8916 6509
rect 8982 6542 9018 6543
rect 9090 6542 9126 6543
rect 8982 6535 9126 6542
rect 8982 6534 9042 6535
rect 8982 6514 8990 6534
rect 9010 6515 9042 6534
rect 9067 6534 9126 6535
rect 9067 6515 9098 6534
rect 9010 6514 9098 6515
rect 9118 6514 9126 6534
rect 8982 6508 9126 6514
rect 9192 6538 9230 6546
rect 9298 6542 9334 6543
rect 9192 6518 9201 6538
rect 9221 6518 9230 6538
rect 9192 6509 9230 6518
rect 9249 6535 9334 6542
rect 9249 6515 9256 6535
rect 9277 6534 9334 6535
rect 9277 6515 9306 6534
rect 9249 6514 9306 6515
rect 9326 6514 9334 6534
rect 9192 6508 9229 6509
rect 9249 6508 9334 6514
rect 9400 6538 9438 6546
rect 9511 6542 9547 6543
rect 9400 6518 9409 6538
rect 9429 6518 9438 6538
rect 9400 6509 9438 6518
rect 9462 6534 9547 6542
rect 9462 6514 9519 6534
rect 9539 6514 9547 6534
rect 9400 6508 9437 6509
rect 9462 6508 9547 6514
rect 9613 6538 9651 6546
rect 9613 6518 9622 6538
rect 9642 6518 9651 6538
rect 9613 6509 9651 6518
rect 9840 6539 9877 6549
rect 9840 6521 9850 6539
rect 9868 6521 9877 6539
rect 9840 6512 9877 6521
rect 10139 6520 10179 6568
rect 11305 6574 11343 6583
rect 11305 6554 11314 6574
rect 11334 6554 11343 6574
rect 11305 6546 11343 6554
rect 11409 6578 11494 6584
rect 11519 6583 11556 6584
rect 11409 6558 11417 6578
rect 11437 6558 11494 6578
rect 11409 6550 11494 6558
rect 11518 6574 11556 6583
rect 11518 6554 11527 6574
rect 11547 6554 11556 6574
rect 11409 6549 11445 6550
rect 11518 6546 11556 6554
rect 11622 6578 11707 6584
rect 11727 6583 11764 6584
rect 11622 6558 11630 6578
rect 11650 6577 11707 6578
rect 11650 6558 11679 6577
rect 11622 6557 11679 6558
rect 11700 6557 11707 6577
rect 11622 6550 11707 6557
rect 11726 6574 11764 6583
rect 11726 6554 11735 6574
rect 11755 6554 11764 6574
rect 11622 6549 11658 6550
rect 11726 6546 11764 6554
rect 11830 6578 11974 6584
rect 11830 6558 11838 6578
rect 11858 6561 11894 6578
rect 11914 6561 11946 6578
rect 11858 6558 11946 6561
rect 11966 6558 11974 6578
rect 11830 6550 11974 6558
rect 11830 6549 11866 6550
rect 11938 6549 11974 6550
rect 12040 6583 12077 6584
rect 12040 6582 12078 6583
rect 12040 6574 12104 6582
rect 12040 6554 12049 6574
rect 12069 6560 12104 6574
rect 12124 6560 12127 6580
rect 12069 6555 12127 6560
rect 12069 6554 12104 6555
rect 10450 6524 10560 6538
rect 10450 6521 10493 6524
rect 10139 6513 10264 6520
rect 10450 6516 10454 6521
rect 9842 6511 9876 6512
rect 9613 6508 9650 6509
rect 9036 6487 9072 6508
rect 9462 6487 9493 6508
rect 10139 6494 10231 6513
rect 10256 6494 10264 6513
rect 8869 6483 8969 6487
rect 8869 6479 8931 6483
rect 8869 6453 8876 6479
rect 8902 6457 8931 6479
rect 8957 6457 8969 6483
rect 8902 6453 8969 6457
rect 8869 6450 8969 6453
rect 9037 6450 9072 6487
rect 9134 6484 9493 6487
rect 9134 6479 9356 6484
rect 9134 6455 9147 6479
rect 9171 6460 9356 6479
rect 9380 6460 9493 6484
rect 9171 6455 9493 6460
rect 9134 6451 9493 6455
rect 9560 6479 9709 6487
rect 9560 6459 9571 6479
rect 9591 6459 9709 6479
rect 10139 6484 10264 6494
rect 10372 6494 10454 6516
rect 10483 6494 10493 6521
rect 10521 6497 10528 6524
rect 10557 6516 10560 6524
rect 11306 6517 11343 6546
rect 10557 6497 10622 6516
rect 11307 6515 11343 6517
rect 11519 6515 11556 6546
rect 11727 6519 11764 6546
rect 12040 6542 12104 6554
rect 10521 6494 10622 6497
rect 10372 6492 10622 6494
rect 10139 6464 10179 6484
rect 9560 6452 9709 6459
rect 10138 6455 10179 6464
rect 9560 6451 9601 6452
rect 8884 6398 8921 6399
rect 8980 6398 9017 6399
rect 9036 6398 9072 6450
rect 9091 6398 9128 6399
rect 8784 6389 8922 6398
rect 8379 6368 8490 6383
rect 8379 6366 8421 6368
rect 8049 6345 8154 6347
rect 7707 6337 7875 6338
rect 8049 6337 8098 6345
rect 7707 6318 8098 6337
rect 8129 6318 8154 6345
rect 8379 6346 8386 6366
rect 8405 6346 8421 6366
rect 8379 6338 8421 6346
rect 8449 6366 8490 6368
rect 8449 6346 8463 6366
rect 8482 6346 8490 6366
rect 8784 6369 8893 6389
rect 8913 6369 8922 6389
rect 8784 6362 8922 6369
rect 8980 6389 9128 6398
rect 8980 6369 8989 6389
rect 9009 6369 9099 6389
rect 9119 6369 9128 6389
rect 8784 6360 8880 6362
rect 8980 6359 9128 6369
rect 9187 6389 9224 6399
rect 9299 6398 9336 6399
rect 9280 6396 9336 6398
rect 9187 6369 9195 6389
rect 9215 6369 9224 6389
rect 9036 6358 9072 6359
rect 8449 6338 8490 6346
rect 8379 6332 8490 6338
rect 7707 6311 8154 6318
rect 7707 6309 7875 6311
rect 6555 6278 6665 6292
rect 6555 6275 6598 6278
rect 6555 6270 6559 6275
rect 6089 6240 6257 6242
rect 5813 6237 6257 6240
rect 5474 6213 5585 6219
rect 5474 6205 5515 6213
rect 5163 6150 5202 6194
rect 5474 6185 5482 6205
rect 5501 6185 5515 6205
rect 5474 6183 5515 6185
rect 5543 6205 5585 6213
rect 5543 6185 5559 6205
rect 5578 6185 5585 6205
rect 5543 6183 5585 6185
rect 5474 6168 5585 6183
rect 5811 6214 6257 6237
rect 5163 6126 5203 6150
rect 5503 6126 5550 6128
rect 5811 6126 5849 6214
rect 6089 6213 6257 6214
rect 6477 6248 6559 6270
rect 6588 6248 6598 6275
rect 6626 6251 6633 6278
rect 6662 6270 6665 6278
rect 6662 6251 6727 6270
rect 6626 6248 6727 6251
rect 6477 6246 6727 6248
rect 6477 6167 6514 6246
rect 6555 6233 6665 6246
rect 6629 6177 6660 6178
rect 6477 6147 6486 6167
rect 6506 6147 6514 6167
rect 6477 6137 6514 6147
rect 6573 6167 6660 6177
rect 6573 6147 6582 6167
rect 6602 6147 6660 6167
rect 6573 6138 6660 6147
rect 6573 6137 6610 6138
rect 5163 6093 5849 6126
rect 5163 6036 5202 6093
rect 5811 6091 5849 6093
rect 6629 6085 6660 6138
rect 6690 6167 6727 6246
rect 6898 6259 7291 6263
rect 6898 6242 6917 6259
rect 6937 6243 7291 6259
rect 7311 6243 7314 6263
rect 6937 6242 7314 6243
rect 6898 6238 7314 6242
rect 6898 6237 7239 6238
rect 6842 6177 6873 6178
rect 6690 6147 6699 6167
rect 6719 6147 6727 6167
rect 6690 6137 6727 6147
rect 6786 6170 6873 6177
rect 6786 6167 6847 6170
rect 6786 6147 6795 6167
rect 6815 6150 6847 6167
rect 6868 6150 6873 6170
rect 6815 6147 6873 6150
rect 6786 6140 6873 6147
rect 6898 6167 6935 6237
rect 7201 6236 7238 6237
rect 7050 6177 7086 6178
rect 6898 6147 6907 6167
rect 6927 6147 6935 6167
rect 6786 6138 6842 6140
rect 6786 6137 6823 6138
rect 6898 6137 6935 6147
rect 6994 6167 7142 6177
rect 7310 6176 7339 6177
rect 7242 6174 7339 6176
rect 6994 6147 7003 6167
rect 7023 6163 7113 6167
rect 7023 6147 7056 6163
rect 6994 6138 7056 6147
rect 6994 6137 7031 6138
rect 7050 6125 7056 6138
rect 7079 6147 7113 6163
rect 7133 6147 7142 6167
rect 7079 6138 7142 6147
rect 7200 6167 7339 6174
rect 7200 6147 7209 6167
rect 7229 6147 7339 6167
rect 7200 6138 7339 6147
rect 7079 6125 7086 6138
rect 7105 6137 7142 6138
rect 7201 6137 7238 6138
rect 7050 6086 7086 6125
rect 6521 6084 6562 6085
rect 6413 6077 6562 6084
rect 6413 6057 6531 6077
rect 6551 6057 6562 6077
rect 6413 6049 6562 6057
rect 6629 6081 6988 6085
rect 6629 6076 6951 6081
rect 6629 6052 6742 6076
rect 6766 6057 6951 6076
rect 6975 6057 6988 6081
rect 6766 6052 6988 6057
rect 6629 6049 6988 6052
rect 7050 6049 7085 6086
rect 7153 6083 7253 6086
rect 7153 6079 7220 6083
rect 7153 6053 7165 6079
rect 7191 6057 7220 6079
rect 7246 6057 7253 6083
rect 7191 6053 7253 6057
rect 7153 6049 7253 6053
rect 5163 6034 5211 6036
rect 5163 6016 5174 6034
rect 5192 6016 5211 6034
rect 6629 6028 6660 6049
rect 7050 6028 7086 6049
rect 6472 6027 6509 6028
rect 5163 6007 5211 6016
rect 5164 6006 5211 6007
rect 5477 6011 5587 6025
rect 5477 6008 5520 6011
rect 5477 6003 5481 6008
rect 5399 5981 5481 6003
rect 5510 5981 5520 6008
rect 5548 5984 5555 6011
rect 5584 6003 5587 6011
rect 6471 6018 6509 6027
rect 5584 5984 5649 6003
rect 6471 5998 6480 6018
rect 6500 5998 6509 6018
rect 5548 5981 5649 5984
rect 5399 5979 5649 5981
rect 5167 5943 5204 5944
rect 4785 5836 4795 5854
rect 4813 5836 4825 5854
rect 4785 5831 4825 5836
rect 5163 5940 5204 5943
rect 5163 5935 5205 5940
rect 5163 5917 5176 5935
rect 5194 5917 5205 5935
rect 5163 5903 5205 5917
rect 5243 5903 5290 5907
rect 5163 5897 5290 5903
rect 5163 5868 5251 5897
rect 5280 5868 5290 5897
rect 5399 5900 5436 5979
rect 5477 5966 5587 5979
rect 5551 5910 5582 5911
rect 5399 5880 5408 5900
rect 5428 5880 5436 5900
rect 5399 5870 5436 5880
rect 5495 5900 5582 5910
rect 5495 5880 5504 5900
rect 5524 5880 5582 5900
rect 5495 5871 5582 5880
rect 5495 5870 5532 5871
rect 5163 5864 5290 5868
rect 5163 5847 5202 5864
rect 5243 5863 5290 5864
rect 4785 5827 4822 5831
rect 5163 5829 5174 5847
rect 5192 5829 5202 5847
rect 5163 5820 5202 5829
rect 5164 5819 5201 5820
rect 5551 5818 5582 5871
rect 5612 5900 5649 5979
rect 5820 5976 6213 5996
rect 6233 5976 6236 5996
rect 6471 5990 6509 5998
rect 6575 6022 6660 6028
rect 6685 6027 6722 6028
rect 6575 6002 6583 6022
rect 6603 6002 6660 6022
rect 6575 5994 6660 6002
rect 6684 6018 6722 6027
rect 6684 5998 6693 6018
rect 6713 5998 6722 6018
rect 6575 5993 6611 5994
rect 6684 5990 6722 5998
rect 6788 6022 6873 6028
rect 6893 6027 6930 6028
rect 6788 6002 6796 6022
rect 6816 6021 6873 6022
rect 6816 6002 6845 6021
rect 6788 6001 6845 6002
rect 6866 6001 6873 6021
rect 6788 5994 6873 6001
rect 6892 6018 6930 6027
rect 6892 5998 6901 6018
rect 6921 5998 6930 6018
rect 6788 5993 6824 5994
rect 6892 5990 6930 5998
rect 6996 6022 7140 6028
rect 6996 6002 7004 6022
rect 7024 6002 7112 6022
rect 7132 6002 7140 6022
rect 6996 5994 7140 6002
rect 6996 5993 7032 5994
rect 7104 5993 7140 5994
rect 7206 6027 7243 6028
rect 7206 6026 7244 6027
rect 7206 6018 7270 6026
rect 7206 5998 7215 6018
rect 7235 6004 7270 6018
rect 7290 6004 7293 6024
rect 7235 5999 7293 6004
rect 7235 5998 7270 5999
rect 5820 5971 6236 5976
rect 5820 5970 6161 5971
rect 5764 5910 5795 5911
rect 5612 5880 5621 5900
rect 5641 5880 5649 5900
rect 5612 5870 5649 5880
rect 5708 5903 5795 5910
rect 5708 5900 5769 5903
rect 5708 5880 5717 5900
rect 5737 5883 5769 5900
rect 5790 5883 5795 5903
rect 5737 5880 5795 5883
rect 5708 5873 5795 5880
rect 5820 5900 5857 5970
rect 6123 5969 6160 5970
rect 6472 5961 6509 5990
rect 6473 5959 6509 5961
rect 6685 5959 6722 5990
rect 6473 5937 6722 5959
rect 6893 5958 6930 5990
rect 7206 5986 7270 5998
rect 7310 5960 7339 6138
rect 7707 6131 7734 6309
rect 7774 6271 7838 6283
rect 8114 6279 8151 6311
rect 8322 6310 8571 6332
rect 8322 6279 8359 6310
rect 8535 6308 8571 6310
rect 8535 6279 8572 6308
rect 8884 6299 8921 6300
rect 9187 6299 9224 6369
rect 9249 6389 9336 6396
rect 9249 6386 9307 6389
rect 9249 6366 9254 6386
rect 9275 6369 9307 6386
rect 9327 6369 9336 6389
rect 9275 6366 9336 6369
rect 9249 6359 9336 6366
rect 9395 6389 9432 6399
rect 9395 6369 9403 6389
rect 9423 6369 9432 6389
rect 9249 6358 9280 6359
rect 8883 6298 9224 6299
rect 8808 6293 9224 6298
rect 7774 6270 7809 6271
rect 7751 6265 7809 6270
rect 7751 6245 7754 6265
rect 7774 6251 7809 6265
rect 7829 6251 7838 6271
rect 7774 6243 7838 6251
rect 7800 6242 7838 6243
rect 7801 6241 7838 6242
rect 7904 6275 7940 6276
rect 8012 6275 8048 6276
rect 7904 6270 8048 6275
rect 7904 6267 7964 6270
rect 7904 6247 7912 6267
rect 7932 6249 7964 6267
rect 7991 6267 8048 6270
rect 7991 6249 8020 6267
rect 7932 6247 8020 6249
rect 8040 6247 8048 6267
rect 7904 6241 8048 6247
rect 8114 6271 8152 6279
rect 8220 6275 8256 6276
rect 8114 6251 8123 6271
rect 8143 6251 8152 6271
rect 8114 6242 8152 6251
rect 8171 6268 8256 6275
rect 8171 6248 8178 6268
rect 8199 6267 8256 6268
rect 8199 6248 8228 6267
rect 8171 6247 8228 6248
rect 8248 6247 8256 6267
rect 8114 6241 8151 6242
rect 8171 6241 8256 6247
rect 8322 6271 8360 6279
rect 8433 6275 8469 6276
rect 8322 6251 8331 6271
rect 8351 6251 8360 6271
rect 8322 6242 8360 6251
rect 8384 6267 8469 6275
rect 8384 6247 8441 6267
rect 8461 6247 8469 6267
rect 8322 6241 8359 6242
rect 8384 6241 8469 6247
rect 8535 6271 8573 6279
rect 8808 6273 8811 6293
rect 8831 6273 9224 6293
rect 9395 6290 9432 6369
rect 9462 6398 9493 6451
rect 9843 6449 9880 6450
rect 9842 6440 9881 6449
rect 9842 6422 9852 6440
rect 9870 6422 9881 6440
rect 10138 6437 10148 6455
rect 10166 6437 10179 6455
rect 10138 6428 10179 6437
rect 10138 6427 10175 6428
rect 9754 6405 9801 6406
rect 9842 6405 9881 6422
rect 9754 6401 9881 6405
rect 9512 6398 9549 6399
rect 9462 6389 9549 6398
rect 9462 6369 9520 6389
rect 9540 6369 9549 6389
rect 9462 6359 9549 6369
rect 9608 6389 9645 6399
rect 9608 6369 9616 6389
rect 9636 6369 9645 6389
rect 9462 6358 9493 6359
rect 9457 6290 9567 6303
rect 9608 6290 9645 6369
rect 9754 6372 9764 6401
rect 9793 6372 9881 6401
rect 10372 6413 10409 6492
rect 10450 6479 10560 6492
rect 10524 6423 10555 6424
rect 10372 6393 10381 6413
rect 10401 6393 10409 6413
rect 10372 6383 10409 6393
rect 10468 6413 10555 6423
rect 10468 6393 10477 6413
rect 10497 6393 10555 6413
rect 10468 6384 10555 6393
rect 10468 6383 10505 6384
rect 9754 6366 9881 6372
rect 9754 6362 9801 6366
rect 9839 6352 9881 6366
rect 10141 6361 10178 6365
rect 9839 6334 9850 6352
rect 9868 6334 9881 6352
rect 9839 6329 9881 6334
rect 9840 6326 9881 6329
rect 10138 6356 10178 6361
rect 10138 6338 10150 6356
rect 10168 6338 10178 6356
rect 9840 6325 9877 6326
rect 9395 6288 9645 6290
rect 9395 6285 9496 6288
rect 8535 6251 8544 6271
rect 8564 6251 8573 6271
rect 9395 6266 9460 6285
rect 8535 6242 8573 6251
rect 9457 6258 9460 6266
rect 9489 6258 9496 6285
rect 9524 6261 9534 6288
rect 9563 6266 9645 6288
rect 9563 6261 9567 6266
rect 9524 6258 9567 6261
rect 9457 6244 9567 6258
rect 9833 6262 9880 6263
rect 9833 6253 9881 6262
rect 8535 6241 8572 6242
rect 7958 6220 7994 6241
rect 8384 6220 8415 6241
rect 9833 6235 9852 6253
rect 9870 6235 9881 6253
rect 9833 6233 9881 6235
rect 7791 6216 7891 6220
rect 7791 6212 7853 6216
rect 7791 6186 7798 6212
rect 7824 6190 7853 6212
rect 7879 6190 7891 6216
rect 7824 6186 7891 6190
rect 7791 6183 7891 6186
rect 7959 6183 7994 6220
rect 8056 6217 8415 6220
rect 8056 6212 8278 6217
rect 8056 6188 8069 6212
rect 8093 6193 8278 6212
rect 8302 6193 8415 6217
rect 8093 6188 8415 6193
rect 8056 6184 8415 6188
rect 8482 6212 8631 6220
rect 8482 6192 8493 6212
rect 8513 6192 8631 6212
rect 8482 6185 8631 6192
rect 8482 6184 8523 6185
rect 7806 6131 7843 6132
rect 7902 6131 7939 6132
rect 7958 6131 7994 6183
rect 8013 6131 8050 6132
rect 7706 6122 7844 6131
rect 7706 6102 7815 6122
rect 7835 6102 7844 6122
rect 7706 6095 7844 6102
rect 7902 6122 8050 6131
rect 7902 6102 7911 6122
rect 7931 6102 8021 6122
rect 8041 6102 8050 6122
rect 7706 6093 7802 6095
rect 7902 6092 8050 6102
rect 8109 6122 8146 6132
rect 8221 6131 8258 6132
rect 8202 6129 8258 6131
rect 8109 6102 8117 6122
rect 8137 6102 8146 6122
rect 7958 6091 7994 6092
rect 7806 6032 7843 6033
rect 8109 6032 8146 6102
rect 8171 6122 8258 6129
rect 8171 6119 8229 6122
rect 8171 6099 8176 6119
rect 8197 6102 8229 6119
rect 8249 6102 8258 6122
rect 8197 6099 8258 6102
rect 8171 6092 8258 6099
rect 8317 6122 8354 6132
rect 8317 6102 8325 6122
rect 8345 6102 8354 6122
rect 8171 6091 8202 6092
rect 7805 6031 8146 6032
rect 7730 6027 8146 6031
rect 7730 6026 8107 6027
rect 7730 6006 7733 6026
rect 7753 6010 8107 6026
rect 8127 6010 8146 6027
rect 7753 6006 8146 6010
rect 8317 6023 8354 6102
rect 8384 6131 8415 6184
rect 9195 6176 9233 6178
rect 9842 6176 9881 6233
rect 9195 6143 9881 6176
rect 8434 6131 8471 6132
rect 8384 6122 8471 6131
rect 8384 6102 8442 6122
rect 8462 6102 8471 6122
rect 8384 6092 8471 6102
rect 8530 6122 8567 6132
rect 8530 6102 8538 6122
rect 8558 6102 8567 6122
rect 8384 6091 8415 6092
rect 8379 6023 8489 6036
rect 8530 6023 8567 6102
rect 8317 6021 8567 6023
rect 8317 6018 8418 6021
rect 8317 5999 8382 6018
rect 8379 5991 8382 5999
rect 8411 5991 8418 6018
rect 8446 5994 8456 6021
rect 8485 5999 8567 6021
rect 8787 6055 8955 6056
rect 9195 6055 9233 6143
rect 9494 6141 9541 6143
rect 9841 6119 9881 6143
rect 8787 6032 9233 6055
rect 9459 6086 9570 6101
rect 9459 6084 9501 6086
rect 9459 6064 9466 6084
rect 9485 6064 9501 6084
rect 9459 6056 9501 6064
rect 9529 6084 9570 6086
rect 9529 6064 9543 6084
rect 9562 6064 9570 6084
rect 9842 6075 9881 6119
rect 9529 6056 9570 6064
rect 9459 6050 9570 6056
rect 8787 6029 9231 6032
rect 8787 6027 8955 6029
rect 8485 5994 8489 5999
rect 8446 5991 8489 5994
rect 8379 5977 8489 5991
rect 7169 5958 7339 5960
rect 6890 5951 7339 5958
rect 6554 5931 6665 5937
rect 6554 5923 6595 5931
rect 5972 5910 6008 5911
rect 5820 5880 5829 5900
rect 5849 5880 5857 5900
rect 5708 5871 5764 5873
rect 5708 5870 5745 5871
rect 5820 5870 5857 5880
rect 5916 5900 6064 5910
rect 6164 5907 6260 5909
rect 5916 5880 5925 5900
rect 5945 5880 6035 5900
rect 6055 5880 6064 5900
rect 5916 5871 6064 5880
rect 6122 5900 6260 5907
rect 6122 5880 6131 5900
rect 6151 5880 6260 5900
rect 6554 5903 6562 5923
rect 6581 5903 6595 5923
rect 6554 5901 6595 5903
rect 6623 5923 6665 5931
rect 6623 5903 6639 5923
rect 6658 5903 6665 5923
rect 6890 5924 6915 5951
rect 6946 5932 7339 5951
rect 6946 5924 6995 5932
rect 7169 5931 7339 5932
rect 6890 5922 6995 5924
rect 6623 5901 6665 5903
rect 6554 5886 6665 5901
rect 6122 5871 6260 5880
rect 5916 5870 5953 5871
rect 5972 5819 6008 5871
rect 6027 5870 6064 5871
rect 6123 5870 6160 5871
rect 5443 5817 5484 5818
rect 5335 5810 5484 5817
rect 4458 5808 4495 5809
rect 4408 5799 4495 5808
rect 4408 5779 4466 5799
rect 4486 5779 4495 5799
rect 4408 5769 4495 5779
rect 4554 5799 4591 5809
rect 4554 5779 4562 5799
rect 4582 5779 4591 5799
rect 5335 5790 5453 5810
rect 5473 5790 5484 5810
rect 5335 5782 5484 5790
rect 5551 5814 5910 5818
rect 5551 5809 5873 5814
rect 5551 5785 5664 5809
rect 5688 5790 5873 5809
rect 5897 5790 5910 5814
rect 5688 5785 5910 5790
rect 5551 5782 5910 5785
rect 5972 5782 6007 5819
rect 6075 5816 6175 5819
rect 6075 5812 6142 5816
rect 6075 5786 6087 5812
rect 6113 5790 6142 5812
rect 6168 5790 6175 5816
rect 6113 5786 6175 5790
rect 6075 5782 6175 5786
rect 4408 5768 4439 5769
rect 4403 5700 4513 5713
rect 4554 5700 4591 5779
rect 4788 5764 4825 5765
rect 4784 5755 4825 5764
rect 5551 5761 5582 5782
rect 5972 5761 6008 5782
rect 5394 5760 5431 5761
rect 5168 5757 5202 5758
rect 4784 5737 4797 5755
rect 4815 5737 4825 5755
rect 4784 5728 4825 5737
rect 5167 5748 5204 5757
rect 5167 5730 5176 5748
rect 5194 5730 5204 5748
rect 4784 5708 4824 5728
rect 5167 5720 5204 5730
rect 5393 5751 5431 5760
rect 5393 5731 5402 5751
rect 5422 5731 5431 5751
rect 5393 5723 5431 5731
rect 5497 5755 5582 5761
rect 5607 5760 5644 5761
rect 5497 5735 5505 5755
rect 5525 5735 5582 5755
rect 5497 5727 5582 5735
rect 5606 5751 5644 5760
rect 5606 5731 5615 5751
rect 5635 5731 5644 5751
rect 5497 5726 5533 5727
rect 5606 5723 5644 5731
rect 5710 5755 5795 5761
rect 5815 5760 5852 5761
rect 5710 5735 5718 5755
rect 5738 5754 5795 5755
rect 5738 5735 5767 5754
rect 5710 5734 5767 5735
rect 5788 5734 5795 5754
rect 5710 5727 5795 5734
rect 5814 5751 5852 5760
rect 5814 5731 5823 5751
rect 5843 5731 5852 5751
rect 5710 5726 5746 5727
rect 5814 5723 5852 5731
rect 5918 5755 6062 5761
rect 5918 5735 5926 5755
rect 5946 5754 6034 5755
rect 5946 5735 5977 5754
rect 5918 5734 5977 5735
rect 6002 5735 6034 5754
rect 6054 5735 6062 5755
rect 6002 5734 6062 5735
rect 5918 5727 6062 5734
rect 5918 5726 5954 5727
rect 6026 5726 6062 5727
rect 6128 5760 6165 5761
rect 6128 5759 6166 5760
rect 6128 5751 6192 5759
rect 6128 5731 6137 5751
rect 6157 5737 6192 5751
rect 6212 5737 6215 5757
rect 6157 5732 6215 5737
rect 6157 5731 6192 5732
rect 4341 5698 4591 5700
rect 4341 5695 4442 5698
rect 2859 5638 2923 5650
rect 3199 5646 3236 5673
rect 3407 5646 3444 5677
rect 3620 5675 3656 5677
rect 4341 5676 4406 5695
rect 3620 5646 3657 5675
rect 4403 5668 4406 5676
rect 4435 5668 4442 5695
rect 4470 5671 4480 5698
rect 4509 5676 4591 5698
rect 4699 5698 4824 5708
rect 4699 5679 4707 5698
rect 4732 5679 4824 5698
rect 4509 5671 4513 5676
rect 4699 5672 4824 5679
rect 4470 5668 4513 5671
rect 4403 5654 4513 5668
rect 2859 5637 2894 5638
rect 2836 5632 2894 5637
rect 2836 5612 2839 5632
rect 2859 5618 2894 5632
rect 2914 5618 2923 5638
rect 2859 5610 2923 5618
rect 2885 5609 2923 5610
rect 2886 5608 2923 5609
rect 2989 5642 3025 5643
rect 3097 5642 3133 5643
rect 2989 5634 3133 5642
rect 2989 5614 2997 5634
rect 3017 5631 3105 5634
rect 3017 5614 3049 5631
rect 3069 5614 3105 5631
rect 3125 5614 3133 5634
rect 2989 5608 3133 5614
rect 3199 5638 3237 5646
rect 3305 5642 3341 5643
rect 3199 5618 3208 5638
rect 3228 5618 3237 5638
rect 3199 5609 3237 5618
rect 3256 5635 3341 5642
rect 3256 5615 3263 5635
rect 3284 5634 3341 5635
rect 3284 5615 3313 5634
rect 3256 5614 3313 5615
rect 3333 5614 3341 5634
rect 3199 5608 3236 5609
rect 3256 5608 3341 5614
rect 3407 5638 3445 5646
rect 3518 5642 3554 5643
rect 3407 5618 3416 5638
rect 3436 5618 3445 5638
rect 3407 5609 3445 5618
rect 3469 5634 3554 5642
rect 3469 5614 3526 5634
rect 3546 5614 3554 5634
rect 3407 5608 3444 5609
rect 3469 5608 3554 5614
rect 3620 5638 3658 5646
rect 3620 5618 3629 5638
rect 3649 5618 3658 5638
rect 3620 5609 3658 5618
rect 4784 5624 4824 5672
rect 5168 5692 5202 5720
rect 5394 5694 5431 5723
rect 5395 5692 5431 5694
rect 5607 5692 5644 5723
rect 5168 5691 5340 5692
rect 5168 5659 5354 5691
rect 5395 5670 5644 5692
rect 5815 5691 5852 5723
rect 6128 5719 6192 5731
rect 6232 5693 6259 5871
rect 8787 5849 8814 6027
rect 8854 5989 8918 6001
rect 9194 5997 9231 6029
rect 9402 6028 9651 6050
rect 9402 5997 9439 6028
rect 9615 6026 9651 6028
rect 9615 5997 9652 6026
rect 8854 5988 8889 5989
rect 8831 5983 8889 5988
rect 8831 5963 8834 5983
rect 8854 5969 8889 5983
rect 8909 5969 8918 5989
rect 8854 5961 8918 5969
rect 8880 5960 8918 5961
rect 8881 5959 8918 5960
rect 8984 5993 9020 5994
rect 9092 5993 9128 5994
rect 8984 5988 9128 5993
rect 8984 5985 9046 5988
rect 8984 5965 8992 5985
rect 9012 5968 9046 5985
rect 9069 5985 9128 5988
rect 9069 5968 9100 5985
rect 9012 5965 9100 5968
rect 9120 5965 9128 5985
rect 8984 5959 9128 5965
rect 9194 5989 9232 5997
rect 9300 5993 9336 5994
rect 9194 5969 9203 5989
rect 9223 5969 9232 5989
rect 9194 5960 9232 5969
rect 9251 5986 9336 5993
rect 9251 5966 9258 5986
rect 9279 5985 9336 5986
rect 9279 5966 9308 5985
rect 9251 5965 9308 5966
rect 9328 5965 9336 5985
rect 9194 5959 9231 5960
rect 9251 5959 9336 5965
rect 9402 5989 9440 5997
rect 9513 5993 9549 5994
rect 9402 5969 9411 5989
rect 9431 5969 9440 5989
rect 9402 5960 9440 5969
rect 9464 5985 9549 5993
rect 9464 5965 9521 5985
rect 9541 5965 9549 5985
rect 9402 5959 9439 5960
rect 9464 5959 9549 5965
rect 9615 5989 9653 5997
rect 9615 5969 9624 5989
rect 9644 5969 9653 5989
rect 9615 5960 9653 5969
rect 9615 5959 9652 5960
rect 9038 5938 9074 5959
rect 9464 5938 9495 5959
rect 8871 5934 8971 5938
rect 8871 5930 8933 5934
rect 8871 5904 8878 5930
rect 8904 5908 8933 5930
rect 8959 5908 8971 5934
rect 8904 5904 8971 5908
rect 8871 5901 8971 5904
rect 9039 5901 9074 5938
rect 9136 5935 9495 5938
rect 9136 5930 9358 5935
rect 9136 5906 9149 5930
rect 9173 5911 9358 5930
rect 9382 5911 9495 5935
rect 9173 5906 9495 5911
rect 9136 5902 9495 5906
rect 9562 5930 9711 5938
rect 9562 5910 9573 5930
rect 9593 5910 9711 5930
rect 9562 5903 9711 5910
rect 9562 5902 9603 5903
rect 8886 5849 8923 5850
rect 8982 5849 9019 5850
rect 9038 5849 9074 5901
rect 9093 5849 9130 5850
rect 8786 5840 8924 5849
rect 8786 5820 8895 5840
rect 8915 5820 8924 5840
rect 8786 5813 8924 5820
rect 8982 5840 9130 5849
rect 8982 5820 8991 5840
rect 9011 5820 9101 5840
rect 9121 5820 9130 5840
rect 8786 5811 8882 5813
rect 8982 5810 9130 5820
rect 9189 5840 9226 5850
rect 9301 5849 9338 5850
rect 9282 5847 9338 5849
rect 9189 5820 9197 5840
rect 9217 5820 9226 5840
rect 9038 5809 9074 5810
rect 6415 5767 6525 5781
rect 6415 5764 6458 5767
rect 6415 5759 6419 5764
rect 6091 5691 6259 5693
rect 5815 5685 6259 5691
rect 5168 5627 5202 5659
rect 3620 5608 3657 5609
rect 3043 5587 3079 5608
rect 3469 5587 3500 5608
rect 4784 5606 4795 5624
rect 4813 5606 4824 5624
rect 4784 5598 4824 5606
rect 5164 5618 5202 5627
rect 5164 5600 5174 5618
rect 5192 5600 5202 5618
rect 4785 5597 4822 5598
rect 5164 5594 5202 5600
rect 5320 5596 5354 5659
rect 5476 5664 5587 5670
rect 5476 5656 5517 5664
rect 5476 5636 5484 5656
rect 5503 5636 5517 5656
rect 5476 5634 5517 5636
rect 5545 5656 5587 5664
rect 5545 5636 5561 5656
rect 5580 5636 5587 5656
rect 5545 5634 5587 5636
rect 5476 5619 5587 5634
rect 5814 5665 6259 5685
rect 5814 5596 5852 5665
rect 6091 5664 6259 5665
rect 6337 5737 6419 5759
rect 6448 5737 6458 5764
rect 6486 5740 6493 5767
rect 6522 5759 6525 5767
rect 8520 5776 8631 5791
rect 8520 5774 8562 5776
rect 6522 5740 6587 5759
rect 6486 5737 6587 5740
rect 6337 5735 6587 5737
rect 6337 5656 6374 5735
rect 6415 5722 6525 5735
rect 6489 5666 6520 5667
rect 6337 5636 6346 5656
rect 6366 5636 6374 5656
rect 6337 5626 6374 5636
rect 6433 5656 6520 5666
rect 6433 5636 6442 5656
rect 6462 5636 6520 5656
rect 6433 5627 6520 5636
rect 6433 5626 6470 5627
rect 5164 5590 5201 5594
rect 2876 5583 2976 5587
rect 2876 5579 2938 5583
rect 2876 5553 2883 5579
rect 2909 5557 2938 5579
rect 2964 5557 2976 5583
rect 2909 5553 2976 5557
rect 2876 5550 2976 5553
rect 3044 5550 3079 5587
rect 3141 5584 3500 5587
rect 3141 5579 3363 5584
rect 3141 5555 3154 5579
rect 3178 5560 3363 5579
rect 3387 5560 3500 5584
rect 3178 5555 3500 5560
rect 3141 5551 3500 5555
rect 3567 5579 3716 5587
rect 5320 5585 5852 5596
rect 3567 5559 3578 5579
rect 3598 5559 3716 5579
rect 5319 5569 5852 5585
rect 6489 5574 6520 5627
rect 6550 5656 6587 5735
rect 6758 5745 7151 5752
rect 6758 5728 6766 5745
rect 6798 5732 7151 5745
rect 7171 5732 7174 5752
rect 8253 5747 8294 5756
rect 6798 5728 7174 5732
rect 6758 5727 7174 5728
rect 7848 5745 8016 5746
rect 8253 5745 8262 5747
rect 6758 5726 7099 5727
rect 6702 5666 6733 5667
rect 6550 5636 6559 5656
rect 6579 5636 6587 5656
rect 6550 5626 6587 5636
rect 6646 5659 6733 5666
rect 6646 5656 6707 5659
rect 6646 5636 6655 5656
rect 6675 5639 6707 5656
rect 6728 5639 6733 5659
rect 6675 5636 6733 5639
rect 6646 5629 6733 5636
rect 6758 5656 6795 5726
rect 7061 5725 7098 5726
rect 7848 5725 8262 5745
rect 8288 5725 8294 5747
rect 8520 5754 8527 5774
rect 8546 5754 8562 5774
rect 8520 5746 8562 5754
rect 8590 5774 8631 5776
rect 8590 5754 8604 5774
rect 8623 5754 8631 5774
rect 8590 5746 8631 5754
rect 8886 5750 8923 5751
rect 9189 5750 9226 5820
rect 9251 5840 9338 5847
rect 9251 5837 9309 5840
rect 9251 5817 9256 5837
rect 9277 5820 9309 5837
rect 9329 5820 9338 5840
rect 9277 5817 9338 5820
rect 9251 5810 9338 5817
rect 9397 5840 9434 5850
rect 9397 5820 9405 5840
rect 9425 5820 9434 5840
rect 9251 5809 9282 5810
rect 8885 5749 9226 5750
rect 8520 5740 8631 5746
rect 8810 5744 9226 5749
rect 7848 5719 8294 5725
rect 7848 5717 8016 5719
rect 6910 5666 6946 5667
rect 6758 5636 6767 5656
rect 6787 5636 6795 5656
rect 6646 5627 6702 5629
rect 6646 5626 6683 5627
rect 6758 5626 6795 5636
rect 6854 5656 7002 5666
rect 7102 5663 7198 5665
rect 6854 5636 6863 5656
rect 6883 5651 6973 5656
rect 6883 5636 6918 5651
rect 6854 5627 6918 5636
rect 6854 5626 6891 5627
rect 6910 5610 6918 5627
rect 6939 5636 6973 5651
rect 6993 5636 7002 5656
rect 6939 5627 7002 5636
rect 7060 5656 7198 5663
rect 7060 5636 7069 5656
rect 7089 5636 7198 5656
rect 7060 5627 7198 5636
rect 6939 5610 6946 5627
rect 6965 5626 7002 5627
rect 7061 5626 7098 5627
rect 6910 5575 6946 5610
rect 6381 5573 6422 5574
rect 5319 5568 5833 5569
rect 3567 5552 3716 5559
rect 6273 5566 6422 5573
rect 4156 5556 4670 5557
rect 3567 5551 3608 5552
rect 2891 5498 2928 5499
rect 2987 5498 3024 5499
rect 3043 5498 3079 5550
rect 3098 5498 3135 5499
rect 2791 5489 2929 5498
rect 2791 5469 2900 5489
rect 2920 5469 2929 5489
rect 2791 5462 2929 5469
rect 2987 5489 3135 5498
rect 2987 5469 2996 5489
rect 3016 5469 3106 5489
rect 3126 5469 3135 5489
rect 2791 5460 2887 5462
rect 2987 5459 3135 5469
rect 3194 5489 3231 5499
rect 3306 5498 3343 5499
rect 3287 5496 3343 5498
rect 3194 5469 3202 5489
rect 3222 5469 3231 5489
rect 3043 5458 3079 5459
rect 1973 5406 2141 5408
rect 1695 5400 2141 5406
rect 763 5376 1179 5381
rect 1358 5379 1469 5385
rect 763 5375 1104 5376
rect 707 5315 738 5316
rect 555 5285 564 5305
rect 584 5285 592 5305
rect 555 5275 592 5285
rect 651 5308 738 5315
rect 651 5305 712 5308
rect 651 5285 660 5305
rect 680 5288 712 5305
rect 733 5288 738 5308
rect 680 5285 738 5288
rect 651 5278 738 5285
rect 763 5305 800 5375
rect 1066 5374 1103 5375
rect 1358 5371 1399 5379
rect 1358 5351 1366 5371
rect 1385 5351 1399 5371
rect 1358 5349 1399 5351
rect 1427 5371 1469 5379
rect 1427 5351 1443 5371
rect 1462 5351 1469 5371
rect 1695 5378 1701 5400
rect 1727 5380 2141 5400
rect 2891 5399 2928 5400
rect 3194 5399 3231 5469
rect 3256 5489 3343 5496
rect 3256 5486 3314 5489
rect 3256 5466 3261 5486
rect 3282 5469 3314 5486
rect 3334 5469 3343 5489
rect 3282 5466 3343 5469
rect 3256 5459 3343 5466
rect 3402 5489 3439 5499
rect 3402 5469 3410 5489
rect 3430 5469 3439 5489
rect 3256 5458 3287 5459
rect 2890 5398 3231 5399
rect 1727 5378 1736 5380
rect 1973 5379 2141 5380
rect 2815 5393 3231 5398
rect 1695 5369 1736 5378
rect 2815 5373 2818 5393
rect 2838 5373 3231 5393
rect 3402 5390 3439 5469
rect 3469 5498 3500 5551
rect 4137 5540 4670 5556
rect 6273 5546 6391 5566
rect 6411 5546 6422 5566
rect 4137 5529 4669 5540
rect 6273 5538 6422 5546
rect 6489 5570 6848 5574
rect 6489 5565 6811 5570
rect 6489 5541 6602 5565
rect 6626 5546 6811 5565
rect 6835 5546 6848 5570
rect 6626 5541 6848 5546
rect 6489 5538 6848 5541
rect 6910 5538 6945 5575
rect 7013 5572 7113 5575
rect 7013 5568 7080 5572
rect 7013 5542 7025 5568
rect 7051 5546 7080 5568
rect 7106 5546 7113 5572
rect 7051 5542 7113 5546
rect 7013 5538 7113 5542
rect 4788 5531 4825 5535
rect 3519 5498 3556 5499
rect 3469 5489 3556 5498
rect 3469 5469 3527 5489
rect 3547 5469 3556 5489
rect 3469 5459 3556 5469
rect 3615 5489 3652 5499
rect 3615 5469 3623 5489
rect 3643 5469 3652 5489
rect 3469 5458 3500 5459
rect 3464 5390 3574 5403
rect 3615 5390 3652 5469
rect 3402 5388 3652 5390
rect 3402 5385 3503 5388
rect 3402 5366 3467 5385
rect 3464 5358 3467 5366
rect 3496 5358 3503 5385
rect 3531 5361 3541 5388
rect 3570 5366 3652 5388
rect 3730 5460 3898 5461
rect 4137 5460 4175 5529
rect 3730 5440 4175 5460
rect 4402 5491 4513 5506
rect 4402 5489 4444 5491
rect 4402 5469 4409 5489
rect 4428 5469 4444 5489
rect 4402 5461 4444 5469
rect 4472 5489 4513 5491
rect 4472 5469 4486 5489
rect 4505 5469 4513 5489
rect 4472 5461 4513 5469
rect 4402 5455 4513 5461
rect 4635 5466 4669 5529
rect 4787 5525 4825 5531
rect 5167 5527 5204 5528
rect 4787 5507 4797 5525
rect 4815 5507 4825 5525
rect 4787 5498 4825 5507
rect 5165 5519 5205 5527
rect 5165 5501 5176 5519
rect 5194 5501 5205 5519
rect 6489 5517 6520 5538
rect 6910 5517 6946 5538
rect 6332 5516 6369 5517
rect 4787 5466 4821 5498
rect 3730 5434 4174 5440
rect 3730 5432 3898 5434
rect 3570 5361 3574 5366
rect 3531 5358 3574 5361
rect 1427 5349 1469 5351
rect 1358 5334 1469 5349
rect 2554 5340 2602 5354
rect 3464 5344 3574 5358
rect 915 5315 951 5316
rect 763 5285 772 5305
rect 792 5285 800 5305
rect 651 5276 707 5278
rect 651 5275 688 5276
rect 763 5275 800 5285
rect 859 5305 1007 5315
rect 1107 5312 1203 5314
rect 859 5285 868 5305
rect 888 5285 978 5305
rect 998 5285 1007 5305
rect 859 5276 1007 5285
rect 1065 5305 1203 5312
rect 1065 5285 1074 5305
rect 1094 5285 1203 5305
rect 1065 5276 1203 5285
rect 2554 5300 2567 5340
rect 2594 5300 2602 5340
rect 2554 5282 2602 5300
rect 859 5275 896 5276
rect 915 5224 951 5276
rect 970 5275 1007 5276
rect 1066 5275 1103 5276
rect 386 5222 427 5223
rect 278 5215 427 5222
rect 278 5195 396 5215
rect 416 5195 427 5215
rect 278 5187 427 5195
rect 494 5219 853 5223
rect 494 5214 816 5219
rect 494 5190 607 5214
rect 631 5195 816 5214
rect 840 5195 853 5219
rect 631 5190 853 5195
rect 494 5187 853 5190
rect 915 5187 950 5224
rect 1018 5221 1118 5224
rect 1018 5217 1085 5221
rect 1018 5191 1030 5217
rect 1056 5195 1085 5217
rect 1111 5195 1118 5221
rect 1056 5191 1118 5195
rect 1018 5187 1118 5191
rect 494 5166 525 5187
rect 915 5166 951 5187
rect 337 5165 374 5166
rect 336 5156 374 5165
rect 336 5136 345 5156
rect 365 5136 374 5156
rect 336 5128 374 5136
rect 440 5160 525 5166
rect 550 5165 587 5166
rect 440 5140 448 5160
rect 468 5140 525 5160
rect 440 5132 525 5140
rect 549 5156 587 5165
rect 549 5136 558 5156
rect 578 5136 587 5156
rect 440 5131 476 5132
rect 549 5128 587 5136
rect 653 5160 738 5166
rect 758 5165 795 5166
rect 653 5140 661 5160
rect 681 5159 738 5160
rect 681 5140 710 5159
rect 653 5139 710 5140
rect 731 5139 738 5159
rect 653 5132 738 5139
rect 757 5156 795 5165
rect 757 5136 766 5156
rect 786 5136 795 5156
rect 653 5131 689 5132
rect 757 5128 795 5136
rect 861 5160 1005 5166
rect 861 5140 869 5160
rect 889 5157 977 5160
rect 889 5140 920 5157
rect 861 5137 920 5140
rect 943 5140 977 5157
rect 997 5140 1005 5160
rect 943 5137 1005 5140
rect 861 5132 1005 5137
rect 861 5131 897 5132
rect 969 5131 1005 5132
rect 1071 5165 1108 5166
rect 1071 5164 1109 5165
rect 1071 5156 1135 5164
rect 1071 5136 1080 5156
rect 1100 5142 1135 5156
rect 1155 5142 1158 5162
rect 1100 5137 1158 5142
rect 1100 5136 1135 5137
rect 337 5099 374 5128
rect 338 5097 374 5099
rect 550 5097 587 5128
rect 338 5075 587 5097
rect 758 5096 795 5128
rect 1071 5124 1135 5136
rect 1175 5098 1202 5276
rect 2549 5175 2602 5282
rect 3730 5254 3757 5432
rect 3797 5394 3861 5406
rect 4137 5402 4174 5434
rect 4345 5433 4594 5455
rect 4635 5434 4821 5466
rect 4649 5433 4821 5434
rect 4345 5402 4382 5433
rect 4558 5431 4594 5433
rect 4558 5402 4595 5431
rect 4787 5405 4821 5433
rect 5165 5453 5205 5501
rect 6331 5507 6369 5516
rect 6331 5487 6340 5507
rect 6360 5487 6369 5507
rect 6331 5479 6369 5487
rect 6435 5511 6520 5517
rect 6545 5516 6582 5517
rect 6435 5491 6443 5511
rect 6463 5491 6520 5511
rect 6435 5483 6520 5491
rect 6544 5507 6582 5516
rect 6544 5487 6553 5507
rect 6573 5487 6582 5507
rect 6435 5482 6471 5483
rect 6544 5479 6582 5487
rect 6648 5511 6733 5517
rect 6753 5516 6790 5517
rect 6648 5491 6656 5511
rect 6676 5510 6733 5511
rect 6676 5491 6705 5510
rect 6648 5490 6705 5491
rect 6726 5490 6733 5510
rect 6648 5483 6733 5490
rect 6752 5507 6790 5516
rect 6752 5487 6761 5507
rect 6781 5487 6790 5507
rect 6648 5482 6684 5483
rect 6752 5479 6790 5487
rect 6856 5511 7000 5517
rect 6856 5491 6864 5511
rect 6884 5491 6972 5511
rect 6992 5491 7000 5511
rect 6856 5483 7000 5491
rect 6856 5482 6892 5483
rect 6964 5482 7000 5483
rect 7066 5516 7103 5517
rect 7066 5515 7104 5516
rect 7066 5507 7130 5515
rect 7066 5487 7075 5507
rect 7095 5493 7130 5507
rect 7150 5493 7153 5513
rect 7095 5488 7153 5493
rect 7095 5487 7130 5488
rect 5476 5457 5586 5471
rect 5476 5454 5519 5457
rect 5165 5446 5290 5453
rect 5476 5449 5480 5454
rect 5165 5427 5257 5446
rect 5282 5427 5290 5446
rect 5165 5417 5290 5427
rect 5398 5427 5480 5449
rect 5509 5427 5519 5454
rect 5547 5430 5554 5457
rect 5583 5449 5586 5457
rect 6332 5450 6369 5479
rect 5583 5430 5648 5449
rect 6333 5448 6369 5450
rect 6545 5448 6582 5479
rect 6753 5452 6790 5479
rect 7066 5475 7130 5487
rect 5547 5427 5648 5430
rect 5398 5425 5648 5427
rect 3797 5393 3832 5394
rect 3774 5388 3832 5393
rect 3774 5368 3777 5388
rect 3797 5374 3832 5388
rect 3852 5374 3861 5394
rect 3797 5366 3861 5374
rect 3823 5365 3861 5366
rect 3824 5364 3861 5365
rect 3927 5398 3963 5399
rect 4035 5398 4071 5399
rect 3927 5391 4071 5398
rect 3927 5390 3987 5391
rect 3927 5370 3935 5390
rect 3955 5371 3987 5390
rect 4012 5390 4071 5391
rect 4012 5371 4043 5390
rect 3955 5370 4043 5371
rect 4063 5370 4071 5390
rect 3927 5364 4071 5370
rect 4137 5394 4175 5402
rect 4243 5398 4279 5399
rect 4137 5374 4146 5394
rect 4166 5374 4175 5394
rect 4137 5365 4175 5374
rect 4194 5391 4279 5398
rect 4194 5371 4201 5391
rect 4222 5390 4279 5391
rect 4222 5371 4251 5390
rect 4194 5370 4251 5371
rect 4271 5370 4279 5390
rect 4137 5364 4174 5365
rect 4194 5364 4279 5370
rect 4345 5394 4383 5402
rect 4456 5398 4492 5399
rect 4345 5374 4354 5394
rect 4374 5374 4383 5394
rect 4345 5365 4383 5374
rect 4407 5390 4492 5398
rect 4407 5370 4464 5390
rect 4484 5370 4492 5390
rect 4345 5364 4382 5365
rect 4407 5364 4492 5370
rect 4558 5394 4596 5402
rect 4558 5374 4567 5394
rect 4587 5374 4596 5394
rect 4558 5365 4596 5374
rect 4785 5395 4822 5405
rect 5165 5397 5205 5417
rect 4785 5377 4795 5395
rect 4813 5377 4822 5395
rect 4785 5368 4822 5377
rect 5164 5388 5205 5397
rect 5164 5370 5174 5388
rect 5192 5370 5205 5388
rect 4787 5367 4821 5368
rect 4558 5364 4595 5365
rect 3981 5343 4017 5364
rect 4407 5343 4438 5364
rect 5164 5361 5205 5370
rect 5164 5360 5201 5361
rect 5398 5346 5435 5425
rect 5476 5412 5586 5425
rect 5550 5356 5581 5357
rect 3814 5339 3914 5343
rect 3814 5335 3876 5339
rect 3814 5309 3821 5335
rect 3847 5313 3876 5335
rect 3902 5313 3914 5339
rect 3847 5309 3914 5313
rect 3814 5306 3914 5309
rect 3982 5306 4017 5343
rect 4079 5340 4438 5343
rect 4079 5335 4301 5340
rect 4079 5311 4092 5335
rect 4116 5316 4301 5335
rect 4325 5316 4438 5340
rect 4116 5311 4438 5316
rect 4079 5307 4438 5311
rect 4505 5335 4654 5343
rect 4505 5315 4516 5335
rect 4536 5315 4654 5335
rect 5398 5326 5407 5346
rect 5427 5326 5435 5346
rect 5398 5316 5435 5326
rect 5494 5346 5581 5356
rect 5494 5326 5503 5346
rect 5523 5326 5581 5346
rect 5494 5317 5581 5326
rect 5494 5316 5531 5317
rect 4505 5308 4654 5315
rect 4505 5307 4546 5308
rect 3829 5254 3866 5255
rect 3925 5254 3962 5255
rect 3981 5254 4017 5306
rect 4036 5254 4073 5255
rect 3729 5245 3867 5254
rect 3729 5225 3838 5245
rect 3858 5225 3867 5245
rect 3355 5205 3466 5220
rect 3729 5218 3867 5225
rect 3925 5245 4073 5254
rect 3925 5225 3934 5245
rect 3954 5225 4044 5245
rect 4064 5225 4073 5245
rect 3729 5216 3825 5218
rect 3925 5215 4073 5225
rect 4132 5245 4169 5255
rect 4244 5254 4281 5255
rect 4225 5252 4281 5254
rect 4132 5225 4140 5245
rect 4160 5225 4169 5245
rect 3981 5214 4017 5215
rect 3355 5203 3397 5205
rect 3355 5183 3362 5203
rect 3381 5183 3397 5203
rect 3355 5175 3397 5183
rect 3425 5203 3466 5205
rect 3425 5183 3439 5203
rect 3458 5183 3466 5203
rect 3425 5175 3466 5183
rect 2549 5174 2851 5175
rect 1468 5153 1578 5167
rect 1468 5150 1511 5153
rect 1468 5145 1472 5150
rect 1034 5096 1202 5098
rect 758 5093 1202 5096
rect 419 5069 530 5075
rect 419 5061 460 5069
rect 108 5006 147 5050
rect 419 5041 427 5061
rect 446 5041 460 5061
rect 419 5039 460 5041
rect 488 5061 530 5069
rect 488 5041 504 5061
rect 523 5041 530 5061
rect 488 5040 530 5041
rect 756 5070 1202 5093
rect 488 5039 531 5040
rect 419 5020 531 5039
rect 108 4982 148 5006
rect 448 4982 495 4983
rect 756 4982 794 5070
rect 1034 5069 1202 5070
rect 1390 5123 1472 5145
rect 1501 5123 1511 5150
rect 1539 5126 1546 5153
rect 1575 5145 1578 5153
rect 2549 5148 3127 5174
rect 3355 5169 3466 5175
rect 2549 5146 2851 5148
rect 2549 5145 2735 5146
rect 1575 5126 1640 5145
rect 1539 5123 1640 5126
rect 1390 5121 1640 5123
rect 1390 5042 1427 5121
rect 1468 5108 1578 5121
rect 1542 5052 1573 5053
rect 1390 5022 1399 5042
rect 1419 5022 1427 5042
rect 1390 5012 1427 5022
rect 1486 5042 1573 5052
rect 1486 5022 1495 5042
rect 1515 5022 1573 5042
rect 1486 5013 1573 5022
rect 1486 5012 1523 5013
rect 108 4972 794 4982
rect 104 4949 794 4972
rect 1542 4960 1573 5013
rect 1603 5042 1640 5121
rect 1811 5118 2204 5138
rect 2224 5118 2227 5138
rect 2549 5137 2602 5145
rect 1811 5113 2227 5118
rect 1811 5112 2152 5113
rect 1755 5052 1786 5053
rect 1603 5022 1612 5042
rect 1632 5022 1640 5042
rect 1603 5012 1640 5022
rect 1699 5045 1786 5052
rect 1699 5042 1760 5045
rect 1699 5022 1708 5042
rect 1728 5025 1760 5042
rect 1781 5025 1786 5045
rect 1728 5022 1786 5025
rect 1699 5015 1786 5022
rect 1811 5042 1848 5112
rect 2114 5111 2151 5112
rect 1963 5052 1999 5053
rect 1811 5022 1820 5042
rect 1840 5022 1848 5042
rect 1699 5013 1755 5015
rect 1699 5012 1736 5013
rect 1811 5012 1848 5022
rect 1907 5042 2055 5052
rect 2155 5049 2251 5051
rect 1907 5022 1916 5042
rect 1936 5022 2026 5042
rect 2046 5022 2055 5042
rect 1907 5013 2055 5022
rect 2113 5042 2251 5049
rect 2113 5022 2122 5042
rect 2142 5022 2251 5042
rect 2113 5013 2251 5022
rect 1907 5012 1944 5013
rect 1963 4961 1999 5013
rect 2018 5012 2055 5013
rect 2114 5012 2151 5013
rect 1434 4959 1475 4960
rect 104 4930 146 4949
rect 756 4947 794 4949
rect 1326 4952 1475 4959
rect 107 4892 146 4930
rect 1326 4932 1444 4952
rect 1464 4932 1475 4952
rect 1326 4924 1475 4932
rect 1542 4956 1901 4960
rect 1542 4951 1864 4956
rect 1542 4927 1655 4951
rect 1679 4932 1864 4951
rect 1888 4932 1901 4956
rect 1679 4927 1901 4932
rect 1542 4924 1901 4927
rect 1963 4924 1998 4961
rect 2066 4958 2166 4961
rect 2066 4954 2133 4958
rect 2066 4928 2078 4954
rect 2104 4932 2133 4954
rect 2159 4932 2166 4958
rect 2104 4928 2166 4932
rect 2066 4924 2166 4928
rect 1542 4903 1573 4924
rect 1963 4903 1999 4924
rect 1385 4902 1422 4903
rect 1384 4893 1422 4902
rect 107 4890 155 4892
rect 107 4872 118 4890
rect 136 4872 155 4890
rect 107 4863 155 4872
rect 108 4862 155 4863
rect 421 4867 531 4881
rect 421 4864 464 4867
rect 421 4859 425 4864
rect 343 4837 425 4859
rect 454 4837 464 4864
rect 492 4840 499 4867
rect 528 4859 531 4867
rect 1384 4873 1393 4893
rect 1413 4873 1422 4893
rect 1384 4865 1422 4873
rect 1488 4897 1573 4903
rect 1598 4902 1635 4903
rect 1488 4877 1496 4897
rect 1516 4877 1573 4897
rect 1488 4869 1573 4877
rect 1597 4893 1635 4902
rect 1597 4873 1606 4893
rect 1626 4873 1635 4893
rect 1488 4868 1524 4869
rect 1597 4865 1635 4873
rect 1701 4897 1786 4903
rect 1806 4902 1843 4903
rect 1701 4877 1709 4897
rect 1729 4896 1786 4897
rect 1729 4877 1758 4896
rect 1701 4876 1758 4877
rect 1779 4876 1786 4896
rect 1701 4869 1786 4876
rect 1805 4893 1843 4902
rect 1805 4873 1814 4893
rect 1834 4873 1843 4893
rect 1701 4868 1737 4869
rect 1805 4865 1843 4873
rect 1909 4899 2053 4903
rect 1909 4897 1966 4899
rect 1909 4877 1917 4897
rect 1937 4877 1966 4897
rect 1909 4875 1966 4877
rect 1992 4897 2053 4899
rect 1992 4877 2025 4897
rect 2045 4877 2053 4897
rect 1992 4875 2053 4877
rect 1909 4869 2053 4875
rect 1909 4868 1945 4869
rect 2017 4868 2053 4869
rect 2119 4902 2156 4903
rect 2119 4901 2157 4902
rect 2119 4893 2183 4901
rect 2119 4873 2128 4893
rect 2148 4879 2183 4893
rect 2203 4879 2206 4899
rect 2148 4874 2206 4879
rect 2148 4873 2183 4874
rect 528 4840 593 4859
rect 492 4837 593 4840
rect 343 4835 593 4837
rect 111 4799 148 4800
rect 107 4796 148 4799
rect 107 4791 149 4796
rect 107 4773 120 4791
rect 138 4773 149 4791
rect 107 4759 149 4773
rect 187 4759 234 4763
rect 107 4753 234 4759
rect 107 4724 195 4753
rect 224 4724 234 4753
rect 343 4756 380 4835
rect 421 4822 531 4835
rect 495 4766 526 4767
rect 343 4736 352 4756
rect 372 4736 380 4756
rect 343 4726 380 4736
rect 439 4756 526 4766
rect 439 4736 448 4756
rect 468 4736 526 4756
rect 439 4727 526 4736
rect 439 4726 476 4727
rect 107 4720 234 4724
rect 107 4703 146 4720
rect 187 4719 234 4720
rect 107 4685 118 4703
rect 136 4685 146 4703
rect 107 4676 146 4685
rect 108 4675 145 4676
rect 495 4674 526 4727
rect 556 4756 593 4835
rect 764 4832 1157 4852
rect 1177 4832 1180 4852
rect 1385 4836 1422 4865
rect 764 4827 1180 4832
rect 1386 4834 1422 4836
rect 1598 4834 1635 4865
rect 764 4826 1105 4827
rect 708 4766 739 4767
rect 556 4736 565 4756
rect 585 4736 593 4756
rect 556 4726 593 4736
rect 652 4759 739 4766
rect 652 4756 713 4759
rect 652 4736 661 4756
rect 681 4739 713 4756
rect 734 4739 739 4759
rect 681 4736 739 4739
rect 652 4729 739 4736
rect 764 4756 801 4826
rect 1067 4825 1104 4826
rect 1386 4812 1635 4834
rect 1806 4833 1843 4865
rect 2119 4861 2183 4873
rect 2223 4836 2250 5013
rect 2683 4968 2710 5145
rect 2750 5108 2814 5120
rect 3090 5116 3127 5148
rect 3298 5147 3547 5169
rect 3829 5155 3866 5156
rect 4132 5155 4169 5225
rect 4194 5245 4281 5252
rect 4194 5242 4252 5245
rect 4194 5222 4199 5242
rect 4220 5225 4252 5242
rect 4272 5225 4281 5245
rect 4220 5222 4281 5225
rect 4194 5215 4281 5222
rect 4340 5245 4377 5255
rect 4340 5225 4348 5245
rect 4368 5225 4377 5245
rect 4194 5214 4225 5215
rect 3828 5154 4169 5155
rect 3298 5116 3335 5147
rect 3511 5145 3547 5147
rect 3753 5149 4169 5154
rect 3511 5116 3548 5145
rect 3753 5129 3756 5149
rect 3776 5129 4169 5149
rect 4340 5146 4377 5225
rect 4407 5254 4438 5307
rect 4788 5305 4825 5306
rect 4787 5296 4826 5305
rect 4787 5278 4797 5296
rect 4815 5278 4826 5296
rect 5167 5294 5204 5298
rect 4699 5261 4746 5262
rect 4787 5261 4826 5278
rect 4699 5257 4826 5261
rect 4457 5254 4494 5255
rect 4407 5245 4494 5254
rect 4407 5225 4465 5245
rect 4485 5225 4494 5245
rect 4407 5215 4494 5225
rect 4553 5245 4590 5255
rect 4553 5225 4561 5245
rect 4581 5225 4590 5245
rect 4407 5214 4438 5215
rect 4402 5146 4512 5159
rect 4553 5146 4590 5225
rect 4699 5228 4709 5257
rect 4738 5228 4826 5257
rect 4699 5222 4826 5228
rect 4699 5218 4746 5222
rect 4784 5208 4826 5222
rect 4784 5190 4795 5208
rect 4813 5190 4826 5208
rect 4784 5185 4826 5190
rect 4785 5182 4826 5185
rect 5164 5289 5204 5294
rect 5164 5271 5176 5289
rect 5194 5271 5204 5289
rect 4785 5181 4822 5182
rect 4340 5144 4590 5146
rect 4340 5141 4441 5144
rect 4340 5122 4405 5141
rect 2750 5107 2785 5108
rect 2727 5102 2785 5107
rect 2727 5082 2730 5102
rect 2750 5088 2785 5102
rect 2805 5088 2814 5108
rect 2750 5080 2814 5088
rect 2776 5079 2814 5080
rect 2777 5078 2814 5079
rect 2880 5112 2916 5113
rect 2988 5112 3024 5113
rect 2880 5105 3024 5112
rect 2880 5104 2937 5105
rect 2880 5084 2888 5104
rect 2908 5085 2937 5104
rect 2962 5104 3024 5105
rect 2962 5085 2996 5104
rect 2908 5084 2996 5085
rect 3016 5084 3024 5104
rect 2880 5078 3024 5084
rect 3090 5108 3128 5116
rect 3196 5112 3232 5113
rect 3090 5088 3099 5108
rect 3119 5088 3128 5108
rect 3090 5079 3128 5088
rect 3147 5105 3232 5112
rect 3147 5085 3154 5105
rect 3175 5104 3232 5105
rect 3175 5085 3204 5104
rect 3147 5084 3204 5085
rect 3224 5084 3232 5104
rect 3090 5078 3127 5079
rect 3147 5078 3232 5084
rect 3298 5108 3336 5116
rect 3409 5112 3445 5113
rect 3298 5088 3307 5108
rect 3327 5088 3336 5108
rect 3298 5079 3336 5088
rect 3360 5104 3445 5112
rect 3360 5084 3417 5104
rect 3437 5084 3445 5104
rect 3298 5078 3335 5079
rect 3360 5078 3445 5084
rect 3511 5108 3549 5116
rect 3511 5088 3520 5108
rect 3540 5088 3549 5108
rect 4402 5114 4405 5122
rect 4434 5114 4441 5141
rect 4469 5117 4479 5144
rect 4508 5122 4590 5144
rect 4508 5117 4512 5122
rect 4469 5114 4512 5117
rect 4402 5100 4512 5114
rect 4778 5118 4825 5119
rect 4778 5109 4826 5118
rect 4778 5091 4797 5109
rect 4815 5091 4826 5109
rect 4778 5089 4826 5091
rect 3511 5079 3549 5088
rect 3511 5078 3548 5079
rect 2934 5057 2970 5078
rect 3360 5057 3391 5078
rect 2767 5053 2867 5057
rect 2767 5049 2829 5053
rect 2767 5023 2774 5049
rect 2800 5027 2829 5049
rect 2855 5027 2867 5053
rect 2800 5023 2867 5027
rect 2767 5020 2867 5023
rect 2935 5020 2970 5057
rect 3032 5054 3391 5057
rect 3032 5049 3254 5054
rect 3032 5025 3045 5049
rect 3069 5030 3254 5049
rect 3278 5030 3391 5054
rect 3069 5025 3391 5030
rect 3032 5021 3391 5025
rect 3458 5049 3607 5057
rect 3458 5029 3469 5049
rect 3489 5029 3607 5049
rect 4787 5051 4826 5089
rect 5164 5091 5204 5271
rect 5550 5264 5581 5317
rect 5611 5346 5648 5425
rect 5819 5422 6212 5442
rect 6232 5422 6235 5442
rect 6333 5426 6582 5448
rect 6751 5447 6792 5452
rect 7170 5449 7197 5627
rect 7848 5539 7875 5717
rect 8253 5714 8294 5719
rect 8463 5718 8712 5740
rect 8810 5724 8813 5744
rect 8833 5724 9226 5744
rect 9397 5741 9434 5820
rect 9464 5849 9495 5902
rect 9841 5895 9881 6075
rect 10138 6158 10178 6338
rect 10524 6331 10555 6384
rect 10585 6413 10622 6492
rect 10793 6489 11186 6509
rect 11206 6489 11209 6509
rect 11307 6493 11556 6515
rect 11725 6514 11766 6519
rect 12144 6516 12171 6694
rect 12822 6606 12849 6784
rect 13227 6781 13268 6786
rect 13437 6785 13686 6807
rect 13784 6791 13787 6811
rect 13807 6791 14200 6811
rect 14371 6808 14408 6887
rect 14438 6916 14469 6969
rect 14815 6962 14855 7142
rect 15193 7144 15232 7201
rect 15842 7199 15880 7201
rect 16413 7198 16562 7205
rect 16413 7178 16531 7198
rect 16551 7178 16562 7198
rect 16413 7170 16562 7178
rect 16629 7202 16988 7206
rect 16629 7197 16951 7202
rect 16629 7173 16742 7197
rect 16766 7178 16951 7197
rect 16975 7178 16988 7202
rect 16766 7173 16988 7178
rect 16629 7170 16988 7173
rect 17050 7170 17085 7207
rect 17153 7204 17253 7207
rect 17153 7200 17220 7204
rect 17153 7174 17165 7200
rect 17191 7178 17220 7200
rect 17246 7178 17253 7204
rect 17191 7174 17253 7178
rect 17153 7170 17253 7174
rect 16629 7149 16660 7170
rect 17050 7149 17086 7170
rect 16472 7148 16509 7149
rect 15193 7142 15241 7144
rect 15193 7124 15204 7142
rect 15222 7124 15241 7142
rect 16471 7139 16509 7148
rect 15193 7115 15241 7124
rect 15194 7114 15241 7115
rect 15507 7119 15617 7133
rect 15507 7116 15550 7119
rect 15507 7111 15511 7116
rect 15429 7089 15511 7111
rect 15540 7089 15550 7116
rect 15578 7092 15585 7119
rect 15614 7111 15617 7119
rect 16471 7119 16480 7139
rect 16500 7119 16509 7139
rect 16471 7111 16509 7119
rect 16575 7143 16660 7149
rect 16685 7148 16722 7149
rect 16575 7123 16583 7143
rect 16603 7123 16660 7143
rect 16575 7115 16660 7123
rect 16684 7139 16722 7148
rect 16684 7119 16693 7139
rect 16713 7119 16722 7139
rect 16575 7114 16611 7115
rect 16684 7111 16722 7119
rect 16788 7143 16873 7149
rect 16893 7148 16930 7149
rect 16788 7123 16796 7143
rect 16816 7142 16873 7143
rect 16816 7123 16845 7142
rect 16788 7122 16845 7123
rect 16866 7122 16873 7142
rect 16788 7115 16873 7122
rect 16892 7139 16930 7148
rect 16892 7119 16901 7139
rect 16921 7119 16930 7139
rect 16788 7114 16824 7115
rect 16892 7111 16930 7119
rect 16996 7143 17140 7149
rect 16996 7123 17004 7143
rect 17024 7141 17112 7143
rect 17024 7123 17053 7141
rect 16996 7122 17053 7123
rect 17082 7123 17112 7141
rect 17132 7123 17140 7143
rect 17082 7122 17140 7123
rect 16996 7115 17140 7122
rect 16996 7114 17032 7115
rect 17104 7114 17140 7115
rect 17206 7148 17243 7149
rect 17206 7147 17244 7148
rect 17206 7139 17270 7147
rect 17206 7119 17215 7139
rect 17235 7125 17270 7139
rect 17290 7125 17293 7145
rect 17235 7120 17293 7125
rect 17235 7119 17270 7120
rect 15614 7092 15679 7111
rect 15578 7089 15679 7092
rect 15429 7087 15679 7089
rect 15197 7051 15234 7052
rect 14815 6944 14825 6962
rect 14843 6944 14855 6962
rect 14815 6939 14855 6944
rect 15193 7048 15234 7051
rect 15193 7043 15235 7048
rect 15193 7025 15206 7043
rect 15224 7025 15235 7043
rect 15193 7011 15235 7025
rect 15273 7011 15320 7015
rect 15193 7005 15320 7011
rect 15193 6976 15281 7005
rect 15310 6976 15320 7005
rect 15429 7008 15466 7087
rect 15507 7074 15617 7087
rect 15581 7018 15612 7019
rect 15429 6988 15438 7008
rect 15458 6988 15466 7008
rect 15429 6978 15466 6988
rect 15525 7008 15612 7018
rect 15525 6988 15534 7008
rect 15554 6988 15612 7008
rect 15525 6979 15612 6988
rect 15525 6978 15562 6979
rect 15193 6972 15320 6976
rect 15193 6955 15232 6972
rect 15273 6971 15320 6972
rect 14815 6935 14852 6939
rect 15193 6937 15204 6955
rect 15222 6937 15232 6955
rect 15193 6928 15232 6937
rect 15194 6927 15231 6928
rect 15581 6926 15612 6979
rect 15642 7008 15679 7087
rect 15850 7084 16243 7104
rect 16263 7084 16266 7104
rect 15850 7079 16266 7084
rect 16472 7082 16509 7111
rect 16473 7080 16509 7082
rect 16685 7080 16722 7111
rect 15850 7078 16191 7079
rect 15794 7018 15825 7019
rect 15642 6988 15651 7008
rect 15671 6988 15679 7008
rect 15642 6978 15679 6988
rect 15738 7011 15825 7018
rect 15738 7008 15799 7011
rect 15738 6988 15747 7008
rect 15767 6991 15799 7008
rect 15820 6991 15825 7011
rect 15767 6988 15825 6991
rect 15738 6981 15825 6988
rect 15850 7008 15887 7078
rect 16153 7077 16190 7078
rect 16473 7058 16722 7080
rect 16893 7079 16930 7111
rect 17206 7107 17270 7119
rect 17310 7083 17337 7259
rect 17768 7226 17795 7396
rect 17835 7366 17899 7378
rect 18175 7374 18212 7406
rect 18383 7405 18632 7427
rect 18915 7407 18952 7408
rect 19218 7407 19255 7477
rect 19280 7497 19367 7504
rect 19280 7494 19338 7497
rect 19280 7474 19285 7494
rect 19306 7477 19338 7494
rect 19358 7477 19367 7497
rect 19306 7474 19367 7477
rect 19280 7467 19367 7474
rect 19426 7497 19463 7507
rect 19426 7477 19434 7497
rect 19454 7477 19463 7497
rect 19280 7466 19311 7467
rect 18914 7406 19255 7407
rect 18383 7374 18420 7405
rect 18596 7403 18632 7405
rect 18596 7374 18633 7403
rect 18839 7401 19255 7406
rect 18839 7381 18842 7401
rect 18862 7381 19255 7401
rect 19426 7398 19463 7477
rect 19493 7506 19524 7559
rect 19874 7557 19911 7558
rect 19873 7548 19912 7557
rect 19873 7530 19883 7548
rect 19901 7530 19912 7548
rect 19785 7513 19832 7514
rect 19873 7513 19912 7530
rect 19785 7509 19912 7513
rect 19543 7506 19580 7507
rect 19493 7497 19580 7506
rect 19493 7477 19551 7497
rect 19571 7477 19580 7497
rect 19493 7467 19580 7477
rect 19639 7497 19676 7507
rect 19639 7477 19647 7497
rect 19667 7477 19676 7497
rect 19493 7466 19524 7467
rect 19488 7398 19598 7411
rect 19639 7398 19676 7477
rect 19785 7480 19795 7509
rect 19824 7480 19912 7509
rect 19785 7474 19912 7480
rect 19785 7470 19832 7474
rect 19870 7460 19912 7474
rect 19870 7442 19881 7460
rect 19899 7442 19912 7460
rect 19870 7437 19912 7442
rect 19871 7434 19912 7437
rect 19871 7433 19908 7434
rect 19426 7396 19676 7398
rect 19426 7393 19527 7396
rect 19426 7374 19491 7393
rect 17835 7365 17870 7366
rect 17812 7360 17870 7365
rect 17812 7340 17815 7360
rect 17835 7346 17870 7360
rect 17890 7346 17899 7366
rect 17835 7338 17899 7346
rect 17861 7337 17899 7338
rect 17862 7336 17899 7337
rect 17965 7370 18001 7371
rect 18073 7370 18109 7371
rect 17965 7362 18109 7370
rect 17965 7342 17973 7362
rect 17993 7342 18081 7362
rect 18101 7342 18109 7362
rect 17965 7336 18109 7342
rect 18175 7366 18213 7374
rect 18281 7370 18317 7371
rect 18175 7346 18184 7366
rect 18204 7346 18213 7366
rect 18175 7337 18213 7346
rect 18232 7363 18317 7370
rect 18232 7343 18239 7363
rect 18260 7362 18317 7363
rect 18260 7343 18289 7362
rect 18232 7342 18289 7343
rect 18309 7342 18317 7362
rect 18175 7336 18212 7337
rect 18232 7336 18317 7342
rect 18383 7366 18421 7374
rect 18494 7370 18530 7371
rect 18383 7346 18392 7366
rect 18412 7346 18421 7366
rect 18383 7337 18421 7346
rect 18445 7362 18530 7370
rect 18445 7342 18502 7362
rect 18522 7342 18530 7362
rect 18383 7336 18420 7337
rect 18445 7336 18530 7342
rect 18596 7366 18634 7374
rect 18596 7346 18605 7366
rect 18625 7346 18634 7366
rect 19488 7366 19491 7374
rect 19520 7366 19527 7393
rect 19555 7369 19565 7396
rect 19594 7374 19676 7396
rect 19594 7369 19598 7374
rect 19555 7366 19598 7369
rect 19488 7352 19598 7366
rect 19864 7370 19911 7371
rect 19864 7361 19912 7370
rect 18596 7337 18634 7346
rect 19864 7343 19883 7361
rect 19901 7343 19912 7361
rect 19864 7341 19912 7343
rect 18596 7336 18633 7337
rect 18019 7315 18055 7336
rect 18445 7315 18476 7336
rect 17852 7311 17952 7315
rect 17852 7307 17914 7311
rect 17852 7281 17859 7307
rect 17885 7285 17914 7307
rect 17940 7285 17952 7311
rect 17885 7281 17952 7285
rect 17852 7278 17952 7281
rect 18020 7278 18055 7315
rect 18117 7312 18476 7315
rect 18117 7307 18339 7312
rect 18117 7283 18130 7307
rect 18154 7288 18339 7307
rect 18363 7288 18476 7312
rect 18154 7283 18476 7288
rect 18117 7279 18476 7283
rect 18543 7307 18692 7315
rect 18543 7287 18554 7307
rect 18574 7287 18692 7307
rect 18543 7280 18692 7287
rect 19225 7284 19263 7286
rect 19873 7284 19912 7341
rect 18543 7279 18584 7280
rect 18019 7238 18055 7278
rect 17867 7226 17904 7227
rect 17963 7226 18000 7227
rect 18019 7226 18024 7238
rect 17767 7217 17905 7226
rect 17767 7197 17876 7217
rect 17896 7197 17905 7217
rect 17767 7190 17905 7197
rect 17963 7217 18024 7226
rect 17963 7197 17972 7217
rect 17992 7206 18024 7217
rect 18051 7226 18055 7238
rect 18074 7226 18111 7227
rect 18051 7217 18111 7226
rect 18051 7206 18082 7217
rect 17992 7197 18082 7206
rect 18102 7197 18111 7217
rect 17767 7188 17863 7190
rect 17963 7187 18111 7197
rect 18170 7217 18207 7227
rect 18282 7226 18319 7227
rect 18263 7224 18319 7226
rect 18170 7197 18178 7217
rect 18198 7197 18207 7217
rect 18019 7186 18055 7187
rect 17867 7127 17904 7128
rect 18170 7127 18207 7197
rect 18232 7217 18319 7224
rect 18232 7214 18290 7217
rect 18232 7194 18237 7214
rect 18258 7197 18290 7214
rect 18310 7197 18319 7217
rect 18258 7194 18319 7197
rect 18232 7187 18319 7194
rect 18378 7217 18415 7227
rect 18378 7197 18386 7217
rect 18406 7197 18415 7217
rect 18232 7186 18263 7187
rect 17866 7126 18207 7127
rect 17791 7121 18207 7126
rect 17791 7103 17794 7121
rect 17814 7119 18207 7121
rect 17814 7103 18184 7119
rect 17832 7101 18184 7103
rect 18175 7099 18184 7101
rect 18205 7099 18207 7119
rect 18175 7087 18207 7099
rect 18378 7118 18415 7197
rect 18445 7226 18476 7279
rect 19225 7251 19911 7284
rect 18495 7226 18532 7227
rect 18445 7217 18532 7226
rect 18445 7197 18503 7217
rect 18523 7197 18532 7217
rect 18445 7187 18532 7197
rect 18591 7217 18628 7227
rect 18591 7197 18599 7217
rect 18619 7197 18628 7217
rect 18445 7186 18476 7187
rect 18440 7118 18550 7131
rect 18591 7118 18628 7197
rect 18378 7116 18628 7118
rect 18378 7113 18479 7116
rect 18378 7094 18443 7113
rect 17218 7081 17337 7083
rect 17169 7079 17337 7081
rect 16554 7052 16665 7058
rect 16893 7053 17337 7079
rect 18440 7086 18443 7094
rect 18472 7086 18479 7113
rect 18507 7089 18517 7116
rect 18546 7094 18628 7116
rect 18817 7163 18985 7164
rect 19225 7163 19263 7251
rect 19524 7249 19571 7251
rect 19871 7227 19911 7251
rect 18817 7140 19263 7163
rect 19489 7194 19600 7208
rect 19489 7192 19531 7194
rect 19489 7172 19496 7192
rect 19515 7172 19531 7192
rect 19489 7164 19531 7172
rect 19559 7192 19600 7194
rect 19559 7172 19573 7192
rect 19592 7172 19600 7192
rect 19872 7183 19911 7227
rect 19559 7164 19600 7172
rect 19489 7158 19600 7164
rect 18817 7137 19261 7140
rect 18817 7135 18985 7137
rect 18546 7089 18550 7094
rect 18507 7086 18550 7089
rect 18440 7072 18550 7086
rect 17169 7052 17337 7053
rect 16554 7044 16595 7052
rect 16554 7024 16562 7044
rect 16581 7024 16595 7044
rect 16554 7022 16595 7024
rect 16623 7044 16665 7052
rect 17218 7051 17326 7052
rect 16623 7024 16639 7044
rect 16658 7024 16665 7044
rect 16623 7022 16665 7024
rect 16002 7018 16038 7019
rect 15850 6988 15859 7008
rect 15879 6988 15887 7008
rect 15738 6979 15794 6981
rect 15738 6978 15775 6979
rect 15850 6978 15887 6988
rect 15946 7008 16094 7018
rect 16194 7015 16290 7017
rect 15946 6988 15955 7008
rect 15975 6988 16065 7008
rect 16085 6988 16094 7008
rect 15946 6979 16094 6988
rect 16152 7008 16290 7015
rect 16152 6988 16161 7008
rect 16181 6988 16290 7008
rect 16554 7007 16665 7022
rect 17256 7050 17326 7051
rect 16152 6979 16290 6988
rect 15946 6978 15983 6979
rect 16002 6927 16038 6979
rect 16057 6978 16094 6979
rect 16153 6978 16190 6979
rect 15473 6925 15514 6926
rect 15365 6918 15514 6925
rect 14488 6916 14525 6917
rect 14438 6907 14525 6916
rect 14438 6887 14496 6907
rect 14516 6887 14525 6907
rect 14438 6877 14525 6887
rect 14584 6907 14621 6917
rect 14584 6887 14592 6907
rect 14612 6887 14621 6907
rect 15365 6898 15483 6918
rect 15503 6898 15514 6918
rect 15365 6890 15514 6898
rect 15581 6922 15940 6926
rect 15581 6917 15903 6922
rect 15581 6893 15694 6917
rect 15718 6898 15903 6917
rect 15927 6898 15940 6922
rect 15718 6893 15940 6898
rect 15581 6890 15940 6893
rect 16002 6890 16037 6927
rect 16105 6924 16205 6927
rect 16105 6920 16172 6924
rect 16105 6894 16117 6920
rect 16143 6898 16172 6920
rect 16198 6898 16205 6924
rect 16143 6894 16205 6898
rect 16105 6890 16205 6894
rect 14438 6876 14469 6877
rect 14433 6808 14543 6821
rect 14584 6808 14621 6887
rect 14818 6872 14855 6873
rect 14814 6863 14855 6872
rect 15581 6869 15612 6890
rect 16002 6869 16038 6890
rect 15424 6868 15461 6869
rect 15198 6865 15232 6866
rect 14814 6845 14827 6863
rect 14845 6845 14855 6863
rect 14814 6836 14855 6845
rect 15197 6856 15234 6865
rect 15197 6838 15206 6856
rect 15224 6838 15234 6856
rect 14814 6816 14854 6836
rect 15197 6828 15234 6838
rect 15423 6859 15461 6868
rect 15423 6839 15432 6859
rect 15452 6839 15461 6859
rect 15423 6831 15461 6839
rect 15527 6863 15612 6869
rect 15637 6868 15674 6869
rect 15527 6843 15535 6863
rect 15555 6843 15612 6863
rect 15527 6835 15612 6843
rect 15636 6859 15674 6868
rect 15636 6839 15645 6859
rect 15665 6839 15674 6859
rect 15527 6834 15563 6835
rect 15636 6831 15674 6839
rect 15740 6863 15825 6869
rect 15845 6868 15882 6869
rect 15740 6843 15748 6863
rect 15768 6862 15825 6863
rect 15768 6843 15797 6862
rect 15740 6842 15797 6843
rect 15818 6842 15825 6862
rect 15740 6835 15825 6842
rect 15844 6859 15882 6868
rect 15844 6839 15853 6859
rect 15873 6839 15882 6859
rect 15740 6834 15776 6835
rect 15844 6831 15882 6839
rect 15948 6863 16092 6869
rect 15948 6843 15956 6863
rect 15976 6862 16064 6863
rect 15976 6843 16007 6862
rect 15948 6842 16007 6843
rect 16032 6843 16064 6862
rect 16084 6843 16092 6863
rect 16032 6842 16092 6843
rect 15948 6835 16092 6842
rect 15948 6834 15984 6835
rect 16056 6834 16092 6835
rect 16158 6868 16195 6869
rect 16158 6867 16196 6868
rect 16158 6859 16222 6867
rect 16158 6839 16167 6859
rect 16187 6845 16222 6859
rect 16242 6845 16245 6865
rect 16187 6840 16245 6845
rect 16187 6839 16222 6840
rect 14371 6806 14621 6808
rect 14371 6803 14472 6806
rect 12889 6746 12953 6758
rect 13229 6754 13266 6781
rect 13437 6754 13474 6785
rect 13650 6783 13686 6785
rect 14371 6784 14436 6803
rect 13650 6754 13687 6783
rect 14433 6776 14436 6784
rect 14465 6776 14472 6803
rect 14500 6779 14510 6806
rect 14539 6784 14621 6806
rect 14729 6806 14854 6816
rect 14729 6787 14737 6806
rect 14762 6787 14854 6806
rect 14539 6779 14543 6784
rect 14729 6780 14854 6787
rect 14500 6776 14543 6779
rect 14433 6762 14543 6776
rect 12889 6745 12924 6746
rect 12866 6740 12924 6745
rect 12866 6720 12869 6740
rect 12889 6726 12924 6740
rect 12944 6726 12953 6746
rect 12889 6718 12953 6726
rect 12915 6717 12953 6718
rect 12916 6716 12953 6717
rect 13019 6750 13055 6751
rect 13127 6750 13163 6751
rect 13019 6742 13163 6750
rect 13019 6722 13027 6742
rect 13047 6722 13135 6742
rect 13155 6722 13163 6742
rect 13019 6716 13163 6722
rect 13229 6746 13267 6754
rect 13335 6750 13371 6751
rect 13229 6726 13238 6746
rect 13258 6726 13267 6746
rect 13229 6717 13267 6726
rect 13286 6743 13371 6750
rect 13286 6723 13293 6743
rect 13314 6742 13371 6743
rect 13314 6723 13343 6742
rect 13286 6722 13343 6723
rect 13363 6722 13371 6742
rect 13229 6716 13266 6717
rect 13286 6716 13371 6722
rect 13437 6746 13475 6754
rect 13548 6750 13584 6751
rect 13437 6726 13446 6746
rect 13466 6726 13475 6746
rect 13437 6717 13475 6726
rect 13499 6742 13584 6750
rect 13499 6722 13556 6742
rect 13576 6722 13584 6742
rect 13437 6716 13474 6717
rect 13499 6716 13584 6722
rect 13650 6746 13688 6754
rect 13650 6726 13659 6746
rect 13679 6726 13688 6746
rect 13650 6717 13688 6726
rect 14814 6732 14854 6780
rect 15198 6800 15232 6828
rect 15424 6802 15461 6831
rect 15425 6800 15461 6802
rect 15637 6800 15674 6831
rect 15198 6799 15370 6800
rect 15198 6767 15384 6799
rect 15425 6778 15674 6800
rect 15845 6799 15882 6831
rect 16158 6827 16222 6839
rect 16262 6801 16289 6979
rect 17256 6943 17317 7050
rect 18817 6957 18844 7135
rect 18884 7097 18948 7109
rect 19224 7105 19261 7137
rect 19432 7136 19681 7158
rect 19432 7105 19469 7136
rect 19645 7134 19681 7136
rect 19645 7105 19682 7134
rect 18884 7096 18919 7097
rect 18861 7091 18919 7096
rect 18861 7071 18864 7091
rect 18884 7077 18919 7091
rect 18939 7077 18948 7097
rect 18884 7069 18948 7077
rect 18910 7068 18948 7069
rect 18911 7067 18948 7068
rect 19014 7101 19050 7102
rect 19122 7101 19158 7102
rect 19014 7096 19158 7101
rect 19014 7093 19076 7096
rect 19014 7073 19022 7093
rect 19042 7076 19076 7093
rect 19099 7093 19158 7096
rect 19099 7076 19130 7093
rect 19042 7073 19130 7076
rect 19150 7073 19158 7093
rect 19014 7067 19158 7073
rect 19224 7097 19262 7105
rect 19330 7101 19366 7102
rect 19224 7077 19233 7097
rect 19253 7077 19262 7097
rect 19224 7068 19262 7077
rect 19281 7094 19366 7101
rect 19281 7074 19288 7094
rect 19309 7093 19366 7094
rect 19309 7074 19338 7093
rect 19281 7073 19338 7074
rect 19358 7073 19366 7093
rect 19224 7067 19261 7068
rect 19281 7067 19366 7073
rect 19432 7097 19470 7105
rect 19543 7101 19579 7102
rect 19432 7077 19441 7097
rect 19461 7077 19470 7097
rect 19432 7068 19470 7077
rect 19494 7093 19579 7101
rect 19494 7073 19551 7093
rect 19571 7073 19579 7093
rect 19432 7067 19469 7068
rect 19494 7067 19579 7073
rect 19645 7097 19683 7105
rect 19645 7077 19654 7097
rect 19674 7077 19683 7097
rect 19645 7068 19683 7077
rect 19645 7067 19682 7068
rect 19068 7046 19104 7067
rect 19494 7046 19525 7067
rect 18901 7042 19001 7046
rect 18901 7038 18963 7042
rect 18901 7012 18908 7038
rect 18934 7016 18963 7038
rect 18989 7016 19001 7042
rect 18934 7012 19001 7016
rect 18901 7009 19001 7012
rect 19069 7009 19104 7046
rect 19166 7043 19525 7046
rect 19166 7038 19388 7043
rect 19166 7014 19179 7038
rect 19203 7019 19388 7038
rect 19412 7019 19525 7043
rect 19203 7014 19525 7019
rect 19166 7010 19525 7014
rect 19592 7038 19741 7046
rect 19592 7018 19603 7038
rect 19623 7018 19741 7038
rect 19592 7011 19741 7018
rect 19592 7010 19633 7011
rect 18916 6957 18953 6958
rect 19012 6957 19049 6958
rect 19068 6957 19104 7009
rect 19123 6957 19160 6958
rect 18816 6948 18954 6957
rect 17256 6932 17326 6943
rect 17256 6923 17263 6932
rect 17258 6903 17263 6923
rect 17311 6903 17326 6932
rect 18816 6928 18925 6948
rect 18945 6928 18954 6948
rect 18816 6921 18954 6928
rect 19012 6948 19160 6957
rect 19012 6928 19021 6948
rect 19041 6928 19131 6948
rect 19151 6928 19160 6948
rect 18816 6919 18912 6921
rect 19012 6918 19160 6928
rect 19219 6948 19256 6958
rect 19331 6957 19368 6958
rect 19312 6955 19368 6957
rect 19219 6928 19227 6948
rect 19247 6928 19256 6948
rect 19068 6917 19104 6918
rect 17258 6894 17326 6903
rect 16445 6875 16555 6889
rect 16445 6872 16488 6875
rect 16445 6867 16449 6872
rect 16121 6799 16289 6801
rect 15845 6793 16289 6799
rect 15198 6735 15232 6767
rect 13650 6716 13687 6717
rect 13073 6695 13109 6716
rect 13499 6695 13530 6716
rect 14814 6714 14825 6732
rect 14843 6714 14854 6732
rect 14814 6706 14854 6714
rect 15194 6726 15232 6735
rect 15194 6708 15204 6726
rect 15222 6708 15232 6726
rect 14815 6705 14852 6706
rect 15194 6702 15232 6708
rect 15350 6704 15384 6767
rect 15506 6772 15617 6778
rect 15506 6764 15547 6772
rect 15506 6744 15514 6764
rect 15533 6744 15547 6764
rect 15506 6742 15547 6744
rect 15575 6764 15617 6772
rect 15575 6744 15591 6764
rect 15610 6744 15617 6764
rect 15575 6742 15617 6744
rect 15506 6727 15617 6742
rect 15844 6773 16289 6793
rect 15844 6704 15882 6773
rect 16121 6772 16289 6773
rect 16367 6845 16449 6867
rect 16478 6845 16488 6872
rect 16516 6848 16523 6875
rect 16552 6867 16555 6875
rect 18550 6884 18661 6899
rect 18550 6882 18592 6884
rect 16552 6848 16617 6867
rect 16516 6845 16617 6848
rect 16367 6843 16617 6845
rect 16367 6764 16404 6843
rect 16445 6830 16555 6843
rect 16519 6774 16550 6775
rect 16367 6744 16376 6764
rect 16396 6744 16404 6764
rect 16367 6734 16404 6744
rect 16463 6764 16550 6774
rect 16463 6744 16472 6764
rect 16492 6744 16550 6764
rect 16463 6735 16550 6744
rect 16463 6734 16500 6735
rect 15194 6698 15231 6702
rect 12906 6691 13006 6695
rect 12906 6687 12968 6691
rect 12906 6661 12913 6687
rect 12939 6665 12968 6687
rect 12994 6665 13006 6691
rect 12939 6661 13006 6665
rect 12906 6658 13006 6661
rect 13074 6658 13109 6695
rect 13171 6692 13530 6695
rect 13171 6687 13393 6692
rect 13171 6663 13184 6687
rect 13208 6668 13393 6687
rect 13417 6668 13530 6692
rect 13208 6663 13530 6668
rect 13171 6659 13530 6663
rect 13597 6687 13746 6695
rect 15350 6693 15882 6704
rect 13597 6667 13608 6687
rect 13628 6667 13746 6687
rect 15349 6677 15882 6693
rect 16519 6682 16550 6735
rect 16580 6764 16617 6843
rect 16788 6840 17181 6860
rect 17201 6840 17204 6860
rect 18283 6855 18324 6864
rect 16788 6835 17204 6840
rect 17878 6853 18046 6854
rect 18283 6853 18292 6855
rect 16788 6834 17129 6835
rect 16732 6774 16763 6775
rect 16580 6744 16589 6764
rect 16609 6744 16617 6764
rect 16580 6734 16617 6744
rect 16676 6767 16763 6774
rect 16676 6764 16737 6767
rect 16676 6744 16685 6764
rect 16705 6747 16737 6764
rect 16758 6747 16763 6767
rect 16705 6744 16763 6747
rect 16676 6737 16763 6744
rect 16788 6764 16825 6834
rect 17091 6833 17128 6834
rect 17878 6833 18292 6853
rect 18318 6833 18324 6855
rect 18550 6862 18557 6882
rect 18576 6862 18592 6882
rect 18550 6854 18592 6862
rect 18620 6882 18661 6884
rect 18620 6862 18634 6882
rect 18653 6862 18661 6882
rect 18620 6854 18661 6862
rect 18916 6858 18953 6859
rect 19219 6858 19256 6928
rect 19281 6948 19368 6955
rect 19281 6945 19339 6948
rect 19281 6925 19286 6945
rect 19307 6928 19339 6945
rect 19359 6928 19368 6948
rect 19307 6925 19368 6928
rect 19281 6918 19368 6925
rect 19427 6948 19464 6958
rect 19427 6928 19435 6948
rect 19455 6928 19464 6948
rect 19281 6917 19312 6918
rect 18915 6857 19256 6858
rect 18550 6848 18661 6854
rect 18840 6852 19256 6857
rect 17878 6827 18324 6833
rect 17878 6825 18046 6827
rect 16940 6774 16976 6775
rect 16788 6744 16797 6764
rect 16817 6744 16825 6764
rect 16676 6735 16732 6737
rect 16676 6734 16713 6735
rect 16788 6734 16825 6744
rect 16884 6764 17032 6774
rect 17132 6771 17228 6773
rect 16884 6744 16893 6764
rect 16913 6744 17003 6764
rect 17023 6744 17032 6764
rect 16884 6735 17032 6744
rect 17090 6764 17228 6771
rect 17090 6744 17099 6764
rect 17119 6744 17228 6764
rect 17090 6735 17228 6744
rect 16884 6734 16921 6735
rect 16940 6683 16976 6735
rect 16995 6734 17032 6735
rect 17091 6734 17128 6735
rect 16411 6681 16452 6682
rect 15349 6676 15863 6677
rect 13597 6660 13746 6667
rect 16303 6674 16452 6681
rect 14186 6664 14700 6665
rect 13597 6659 13638 6660
rect 13073 6623 13109 6658
rect 12921 6606 12958 6607
rect 13017 6606 13054 6607
rect 13073 6606 13080 6623
rect 12821 6597 12959 6606
rect 12821 6577 12930 6597
rect 12950 6577 12959 6597
rect 12821 6570 12959 6577
rect 13017 6597 13080 6606
rect 13017 6577 13026 6597
rect 13046 6582 13080 6597
rect 13101 6606 13109 6623
rect 13128 6606 13165 6607
rect 13101 6597 13165 6606
rect 13101 6582 13136 6597
rect 13046 6577 13136 6582
rect 13156 6577 13165 6597
rect 12821 6568 12917 6570
rect 13017 6567 13165 6577
rect 13224 6597 13261 6607
rect 13336 6606 13373 6607
rect 13317 6604 13373 6606
rect 13224 6577 13232 6597
rect 13252 6577 13261 6597
rect 13073 6566 13109 6567
rect 12003 6514 12171 6516
rect 11725 6508 12171 6514
rect 10793 6484 11209 6489
rect 11388 6487 11499 6493
rect 10793 6483 11134 6484
rect 10737 6423 10768 6424
rect 10585 6393 10594 6413
rect 10614 6393 10622 6413
rect 10585 6383 10622 6393
rect 10681 6416 10768 6423
rect 10681 6413 10742 6416
rect 10681 6393 10690 6413
rect 10710 6396 10742 6413
rect 10763 6396 10768 6416
rect 10710 6393 10768 6396
rect 10681 6386 10768 6393
rect 10793 6413 10830 6483
rect 11096 6482 11133 6483
rect 11388 6479 11429 6487
rect 11388 6459 11396 6479
rect 11415 6459 11429 6479
rect 11388 6457 11429 6459
rect 11457 6479 11499 6487
rect 11457 6459 11473 6479
rect 11492 6459 11499 6479
rect 11725 6486 11731 6508
rect 11757 6488 12171 6508
rect 12921 6507 12958 6508
rect 13224 6507 13261 6577
rect 13286 6597 13373 6604
rect 13286 6594 13344 6597
rect 13286 6574 13291 6594
rect 13312 6577 13344 6594
rect 13364 6577 13373 6597
rect 13312 6574 13373 6577
rect 13286 6567 13373 6574
rect 13432 6597 13469 6607
rect 13432 6577 13440 6597
rect 13460 6577 13469 6597
rect 13286 6566 13317 6567
rect 12920 6506 13261 6507
rect 11757 6486 11766 6488
rect 12003 6487 12171 6488
rect 12845 6505 13261 6506
rect 12845 6501 13221 6505
rect 11725 6477 11766 6486
rect 12845 6481 12848 6501
rect 12868 6488 13221 6501
rect 13253 6488 13261 6505
rect 12868 6481 13261 6488
rect 13432 6498 13469 6577
rect 13499 6606 13530 6659
rect 14167 6648 14700 6664
rect 16303 6654 16421 6674
rect 16441 6654 16452 6674
rect 14167 6637 14699 6648
rect 16303 6646 16452 6654
rect 16519 6678 16878 6682
rect 16519 6673 16841 6678
rect 16519 6649 16632 6673
rect 16656 6654 16841 6673
rect 16865 6654 16878 6678
rect 16656 6649 16878 6654
rect 16519 6646 16878 6649
rect 16940 6646 16975 6683
rect 17043 6680 17143 6683
rect 17043 6676 17110 6680
rect 17043 6650 17055 6676
rect 17081 6654 17110 6676
rect 17136 6654 17143 6680
rect 17081 6650 17143 6654
rect 17043 6646 17143 6650
rect 14818 6639 14855 6643
rect 13549 6606 13586 6607
rect 13499 6597 13586 6606
rect 13499 6577 13557 6597
rect 13577 6577 13586 6597
rect 13499 6567 13586 6577
rect 13645 6597 13682 6607
rect 13645 6577 13653 6597
rect 13673 6577 13682 6597
rect 13499 6566 13530 6567
rect 13494 6498 13604 6511
rect 13645 6498 13682 6577
rect 13432 6496 13682 6498
rect 13432 6493 13533 6496
rect 13432 6474 13497 6493
rect 11457 6457 11499 6459
rect 11388 6442 11499 6457
rect 13494 6466 13497 6474
rect 13526 6466 13533 6493
rect 13561 6469 13571 6496
rect 13600 6474 13682 6496
rect 13760 6568 13928 6569
rect 14167 6568 14205 6637
rect 13760 6548 14205 6568
rect 14432 6599 14543 6614
rect 14432 6597 14474 6599
rect 14432 6577 14439 6597
rect 14458 6577 14474 6597
rect 14432 6569 14474 6577
rect 14502 6597 14543 6599
rect 14502 6577 14516 6597
rect 14535 6577 14543 6597
rect 14502 6569 14543 6577
rect 14432 6563 14543 6569
rect 14665 6574 14699 6637
rect 14817 6633 14855 6639
rect 15197 6635 15234 6636
rect 14817 6615 14827 6633
rect 14845 6615 14855 6633
rect 14817 6606 14855 6615
rect 15195 6627 15235 6635
rect 15195 6609 15206 6627
rect 15224 6609 15235 6627
rect 16519 6625 16550 6646
rect 16940 6625 16976 6646
rect 16362 6624 16399 6625
rect 14817 6574 14851 6606
rect 13760 6542 14204 6548
rect 13760 6540 13928 6542
rect 13600 6469 13604 6474
rect 13561 6466 13604 6469
rect 13494 6452 13604 6466
rect 10945 6423 10981 6424
rect 10793 6393 10802 6413
rect 10822 6393 10830 6413
rect 10681 6384 10737 6386
rect 10681 6383 10718 6384
rect 10793 6383 10830 6393
rect 10889 6413 11037 6423
rect 11137 6420 11233 6422
rect 10889 6393 10898 6413
rect 10918 6393 11008 6413
rect 11028 6393 11037 6413
rect 10889 6384 11037 6393
rect 11095 6413 11233 6420
rect 11095 6393 11104 6413
rect 11124 6393 11233 6413
rect 11095 6384 11233 6393
rect 10889 6383 10926 6384
rect 10945 6332 10981 6384
rect 11000 6383 11037 6384
rect 11096 6383 11133 6384
rect 10416 6330 10457 6331
rect 10308 6323 10457 6330
rect 10308 6303 10426 6323
rect 10446 6303 10457 6323
rect 10308 6295 10457 6303
rect 10524 6327 10883 6331
rect 10524 6322 10846 6327
rect 10524 6298 10637 6322
rect 10661 6303 10846 6322
rect 10870 6303 10883 6327
rect 10661 6298 10883 6303
rect 10524 6295 10883 6298
rect 10945 6295 10980 6332
rect 11048 6329 11148 6332
rect 11048 6325 11115 6329
rect 11048 6299 11060 6325
rect 11086 6303 11115 6325
rect 11141 6303 11148 6329
rect 11086 6299 11148 6303
rect 11048 6295 11148 6299
rect 10524 6274 10555 6295
rect 10945 6274 10981 6295
rect 10367 6273 10404 6274
rect 10366 6264 10404 6273
rect 10366 6244 10375 6264
rect 10395 6244 10404 6264
rect 10366 6236 10404 6244
rect 10470 6268 10555 6274
rect 10580 6273 10617 6274
rect 10470 6248 10478 6268
rect 10498 6248 10555 6268
rect 10470 6240 10555 6248
rect 10579 6264 10617 6273
rect 10579 6244 10588 6264
rect 10608 6244 10617 6264
rect 10470 6239 10506 6240
rect 10579 6236 10617 6244
rect 10683 6268 10768 6274
rect 10788 6273 10825 6274
rect 10683 6248 10691 6268
rect 10711 6267 10768 6268
rect 10711 6248 10740 6267
rect 10683 6247 10740 6248
rect 10761 6247 10768 6267
rect 10683 6240 10768 6247
rect 10787 6264 10825 6273
rect 10787 6244 10796 6264
rect 10816 6244 10825 6264
rect 10683 6239 10719 6240
rect 10787 6236 10825 6244
rect 10891 6268 11035 6274
rect 10891 6248 10899 6268
rect 10919 6265 11007 6268
rect 10919 6248 10950 6265
rect 10891 6245 10950 6248
rect 10973 6248 11007 6265
rect 11027 6248 11035 6268
rect 10973 6245 11035 6248
rect 10891 6240 11035 6245
rect 10891 6239 10927 6240
rect 10999 6239 11035 6240
rect 11101 6273 11138 6274
rect 11101 6272 11139 6273
rect 11101 6264 11165 6272
rect 11101 6244 11110 6264
rect 11130 6250 11165 6264
rect 11185 6250 11188 6270
rect 11130 6245 11188 6250
rect 11130 6244 11165 6245
rect 10367 6207 10404 6236
rect 10368 6205 10404 6207
rect 10580 6205 10617 6236
rect 10368 6183 10617 6205
rect 10788 6204 10825 6236
rect 11101 6232 11165 6244
rect 11205 6206 11232 6384
rect 13760 6362 13787 6540
rect 13827 6502 13891 6514
rect 14167 6510 14204 6542
rect 14375 6541 14624 6563
rect 14665 6542 14851 6574
rect 14679 6541 14851 6542
rect 14375 6510 14412 6541
rect 14588 6539 14624 6541
rect 14588 6510 14625 6539
rect 14817 6513 14851 6541
rect 15195 6561 15235 6609
rect 16361 6615 16399 6624
rect 16361 6595 16370 6615
rect 16390 6595 16399 6615
rect 16361 6587 16399 6595
rect 16465 6619 16550 6625
rect 16575 6624 16612 6625
rect 16465 6599 16473 6619
rect 16493 6599 16550 6619
rect 16465 6591 16550 6599
rect 16574 6615 16612 6624
rect 16574 6595 16583 6615
rect 16603 6595 16612 6615
rect 16465 6590 16501 6591
rect 16574 6587 16612 6595
rect 16678 6619 16763 6625
rect 16783 6624 16820 6625
rect 16678 6599 16686 6619
rect 16706 6618 16763 6619
rect 16706 6599 16735 6618
rect 16678 6598 16735 6599
rect 16756 6598 16763 6618
rect 16678 6591 16763 6598
rect 16782 6615 16820 6624
rect 16782 6595 16791 6615
rect 16811 6595 16820 6615
rect 16678 6590 16714 6591
rect 16782 6587 16820 6595
rect 16886 6619 17030 6625
rect 16886 6599 16894 6619
rect 16914 6602 16950 6619
rect 16970 6602 17002 6619
rect 16914 6599 17002 6602
rect 17022 6599 17030 6619
rect 16886 6591 17030 6599
rect 16886 6590 16922 6591
rect 16994 6590 17030 6591
rect 17096 6624 17133 6625
rect 17096 6623 17134 6624
rect 17096 6615 17160 6623
rect 17096 6595 17105 6615
rect 17125 6601 17160 6615
rect 17180 6601 17183 6621
rect 17125 6596 17183 6601
rect 17125 6595 17160 6596
rect 15506 6565 15616 6579
rect 15506 6562 15549 6565
rect 15195 6554 15320 6561
rect 15506 6557 15510 6562
rect 15195 6535 15287 6554
rect 15312 6535 15320 6554
rect 15195 6525 15320 6535
rect 15428 6535 15510 6557
rect 15539 6535 15549 6562
rect 15577 6538 15584 6565
rect 15613 6557 15616 6565
rect 16362 6558 16399 6587
rect 15613 6538 15678 6557
rect 16363 6556 16399 6558
rect 16575 6556 16612 6587
rect 16783 6560 16820 6587
rect 17096 6583 17160 6595
rect 15577 6535 15678 6538
rect 15428 6533 15678 6535
rect 13827 6501 13862 6502
rect 13804 6496 13862 6501
rect 13804 6476 13807 6496
rect 13827 6482 13862 6496
rect 13882 6482 13891 6502
rect 13827 6474 13891 6482
rect 13853 6473 13891 6474
rect 13854 6472 13891 6473
rect 13957 6506 13993 6507
rect 14065 6506 14101 6507
rect 13957 6499 14101 6506
rect 13957 6498 14017 6499
rect 13957 6478 13965 6498
rect 13985 6479 14017 6498
rect 14042 6498 14101 6499
rect 14042 6479 14073 6498
rect 13985 6478 14073 6479
rect 14093 6478 14101 6498
rect 13957 6472 14101 6478
rect 14167 6502 14205 6510
rect 14273 6506 14309 6507
rect 14167 6482 14176 6502
rect 14196 6482 14205 6502
rect 14167 6473 14205 6482
rect 14224 6499 14309 6506
rect 14224 6479 14231 6499
rect 14252 6498 14309 6499
rect 14252 6479 14281 6498
rect 14224 6478 14281 6479
rect 14301 6478 14309 6498
rect 14167 6472 14204 6473
rect 14224 6472 14309 6478
rect 14375 6502 14413 6510
rect 14486 6506 14522 6507
rect 14375 6482 14384 6502
rect 14404 6482 14413 6502
rect 14375 6473 14413 6482
rect 14437 6498 14522 6506
rect 14437 6478 14494 6498
rect 14514 6478 14522 6498
rect 14375 6472 14412 6473
rect 14437 6472 14522 6478
rect 14588 6502 14626 6510
rect 14588 6482 14597 6502
rect 14617 6482 14626 6502
rect 14588 6473 14626 6482
rect 14815 6503 14852 6513
rect 15195 6505 15235 6525
rect 14815 6485 14825 6503
rect 14843 6485 14852 6503
rect 14815 6476 14852 6485
rect 15194 6496 15235 6505
rect 15194 6478 15204 6496
rect 15222 6478 15235 6496
rect 14817 6475 14851 6476
rect 14588 6472 14625 6473
rect 14011 6451 14047 6472
rect 14437 6451 14468 6472
rect 15194 6469 15235 6478
rect 15194 6468 15231 6469
rect 15428 6454 15465 6533
rect 15506 6520 15616 6533
rect 15580 6464 15611 6465
rect 13844 6447 13944 6451
rect 13844 6443 13906 6447
rect 13844 6417 13851 6443
rect 13877 6421 13906 6443
rect 13932 6421 13944 6447
rect 13877 6417 13944 6421
rect 13844 6414 13944 6417
rect 14012 6414 14047 6451
rect 14109 6448 14468 6451
rect 14109 6443 14331 6448
rect 14109 6419 14122 6443
rect 14146 6424 14331 6443
rect 14355 6424 14468 6448
rect 14146 6419 14468 6424
rect 14109 6415 14468 6419
rect 14535 6443 14684 6451
rect 14535 6423 14546 6443
rect 14566 6423 14684 6443
rect 15428 6434 15437 6454
rect 15457 6434 15465 6454
rect 15428 6424 15465 6434
rect 15524 6454 15611 6464
rect 15524 6434 15533 6454
rect 15553 6434 15611 6454
rect 15524 6425 15611 6434
rect 15524 6424 15561 6425
rect 14535 6416 14684 6423
rect 14535 6415 14576 6416
rect 13859 6362 13896 6363
rect 13955 6362 13992 6363
rect 14011 6362 14047 6414
rect 14066 6362 14103 6363
rect 13759 6353 13897 6362
rect 13354 6332 13465 6347
rect 13354 6330 13396 6332
rect 13024 6309 13129 6311
rect 12682 6301 12850 6302
rect 13024 6301 13073 6309
rect 12682 6282 13073 6301
rect 13104 6282 13129 6309
rect 13354 6310 13361 6330
rect 13380 6310 13396 6330
rect 13354 6302 13396 6310
rect 13424 6330 13465 6332
rect 13424 6310 13438 6330
rect 13457 6310 13465 6330
rect 13759 6333 13868 6353
rect 13888 6333 13897 6353
rect 13759 6326 13897 6333
rect 13955 6353 14103 6362
rect 13955 6333 13964 6353
rect 13984 6333 14074 6353
rect 14094 6333 14103 6353
rect 13759 6324 13855 6326
rect 13955 6323 14103 6333
rect 14162 6353 14199 6363
rect 14274 6362 14311 6363
rect 14255 6360 14311 6362
rect 14162 6333 14170 6353
rect 14190 6333 14199 6353
rect 14011 6322 14047 6323
rect 13424 6302 13465 6310
rect 13354 6296 13465 6302
rect 12682 6275 13129 6282
rect 12682 6273 12850 6275
rect 11530 6242 11640 6256
rect 11530 6239 11573 6242
rect 11530 6234 11534 6239
rect 11064 6204 11232 6206
rect 10788 6201 11232 6204
rect 10449 6177 10560 6183
rect 10449 6169 10490 6177
rect 10138 6114 10177 6158
rect 10449 6149 10457 6169
rect 10476 6149 10490 6169
rect 10449 6147 10490 6149
rect 10518 6169 10560 6177
rect 10518 6149 10534 6169
rect 10553 6149 10560 6169
rect 10518 6147 10560 6149
rect 10449 6132 10560 6147
rect 10786 6178 11232 6201
rect 10138 6090 10178 6114
rect 10478 6090 10525 6092
rect 10786 6090 10824 6178
rect 11064 6177 11232 6178
rect 11452 6212 11534 6234
rect 11563 6212 11573 6239
rect 11601 6215 11608 6242
rect 11637 6234 11640 6242
rect 11637 6215 11702 6234
rect 11601 6212 11702 6215
rect 11452 6210 11702 6212
rect 11452 6131 11489 6210
rect 11530 6197 11640 6210
rect 11604 6141 11635 6142
rect 11452 6111 11461 6131
rect 11481 6111 11489 6131
rect 11452 6101 11489 6111
rect 11548 6131 11635 6141
rect 11548 6111 11557 6131
rect 11577 6111 11635 6131
rect 11548 6102 11635 6111
rect 11548 6101 11585 6102
rect 10138 6057 10824 6090
rect 10138 6000 10177 6057
rect 10786 6055 10824 6057
rect 11604 6049 11635 6102
rect 11665 6131 11702 6210
rect 11873 6223 12266 6227
rect 11873 6206 11892 6223
rect 11912 6207 12266 6223
rect 12286 6207 12289 6227
rect 11912 6206 12289 6207
rect 11873 6202 12289 6206
rect 11873 6201 12214 6202
rect 11817 6141 11848 6142
rect 11665 6111 11674 6131
rect 11694 6111 11702 6131
rect 11665 6101 11702 6111
rect 11761 6134 11848 6141
rect 11761 6131 11822 6134
rect 11761 6111 11770 6131
rect 11790 6114 11822 6131
rect 11843 6114 11848 6134
rect 11790 6111 11848 6114
rect 11761 6104 11848 6111
rect 11873 6131 11910 6201
rect 12176 6200 12213 6201
rect 12025 6141 12061 6142
rect 11873 6111 11882 6131
rect 11902 6111 11910 6131
rect 11761 6102 11817 6104
rect 11761 6101 11798 6102
rect 11873 6101 11910 6111
rect 11969 6131 12117 6141
rect 12285 6140 12314 6141
rect 12217 6138 12314 6140
rect 11969 6111 11978 6131
rect 11998 6127 12088 6131
rect 11998 6111 12031 6127
rect 11969 6102 12031 6111
rect 11969 6101 12006 6102
rect 12025 6089 12031 6102
rect 12054 6111 12088 6127
rect 12108 6111 12117 6131
rect 12054 6102 12117 6111
rect 12175 6131 12314 6138
rect 12175 6111 12184 6131
rect 12204 6111 12314 6131
rect 12175 6102 12314 6111
rect 12054 6089 12061 6102
rect 12080 6101 12117 6102
rect 12176 6101 12213 6102
rect 12025 6050 12061 6089
rect 11496 6048 11537 6049
rect 11388 6041 11537 6048
rect 11388 6021 11506 6041
rect 11526 6021 11537 6041
rect 11388 6013 11537 6021
rect 11604 6045 11963 6049
rect 11604 6040 11926 6045
rect 11604 6016 11717 6040
rect 11741 6021 11926 6040
rect 11950 6021 11963 6045
rect 11741 6016 11963 6021
rect 11604 6013 11963 6016
rect 12025 6013 12060 6050
rect 12128 6047 12228 6050
rect 12128 6043 12195 6047
rect 12128 6017 12140 6043
rect 12166 6021 12195 6043
rect 12221 6021 12228 6047
rect 12166 6017 12228 6021
rect 12128 6013 12228 6017
rect 10138 5998 10186 6000
rect 10138 5980 10149 5998
rect 10167 5980 10186 5998
rect 11604 5992 11635 6013
rect 12025 5992 12061 6013
rect 11447 5991 11484 5992
rect 10138 5971 10186 5980
rect 10139 5970 10186 5971
rect 10452 5975 10562 5989
rect 10452 5972 10495 5975
rect 10452 5967 10456 5972
rect 10374 5945 10456 5967
rect 10485 5945 10495 5972
rect 10523 5948 10530 5975
rect 10559 5967 10562 5975
rect 11446 5982 11484 5991
rect 10559 5948 10624 5967
rect 11446 5962 11455 5982
rect 11475 5962 11484 5982
rect 10523 5945 10624 5948
rect 10374 5943 10624 5945
rect 10142 5907 10179 5908
rect 9841 5877 9851 5895
rect 9869 5877 9881 5895
rect 9841 5872 9881 5877
rect 10138 5904 10179 5907
rect 10138 5899 10180 5904
rect 10138 5881 10151 5899
rect 10169 5881 10180 5899
rect 9841 5868 9878 5872
rect 10138 5867 10180 5881
rect 10218 5867 10265 5871
rect 10138 5861 10265 5867
rect 9514 5849 9551 5850
rect 9464 5840 9551 5849
rect 9464 5820 9522 5840
rect 9542 5820 9551 5840
rect 9464 5810 9551 5820
rect 9610 5840 9647 5850
rect 9610 5820 9618 5840
rect 9638 5820 9647 5840
rect 9464 5809 9495 5810
rect 9459 5741 9569 5754
rect 9610 5741 9647 5820
rect 10138 5832 10226 5861
rect 10255 5832 10265 5861
rect 10374 5864 10411 5943
rect 10452 5930 10562 5943
rect 10526 5874 10557 5875
rect 10374 5844 10383 5864
rect 10403 5844 10411 5864
rect 10374 5834 10411 5844
rect 10470 5864 10557 5874
rect 10470 5844 10479 5864
rect 10499 5844 10557 5864
rect 10470 5835 10557 5844
rect 10470 5834 10507 5835
rect 10138 5828 10265 5832
rect 10138 5811 10177 5828
rect 10218 5827 10265 5828
rect 9844 5805 9881 5806
rect 9840 5796 9881 5805
rect 9840 5778 9853 5796
rect 9871 5778 9881 5796
rect 10138 5793 10149 5811
rect 10167 5793 10177 5811
rect 10138 5784 10177 5793
rect 10139 5783 10176 5784
rect 10526 5782 10557 5835
rect 10587 5864 10624 5943
rect 10795 5940 11188 5960
rect 11208 5940 11211 5960
rect 11446 5954 11484 5962
rect 11550 5986 11635 5992
rect 11660 5991 11697 5992
rect 11550 5966 11558 5986
rect 11578 5966 11635 5986
rect 11550 5958 11635 5966
rect 11659 5982 11697 5991
rect 11659 5962 11668 5982
rect 11688 5962 11697 5982
rect 11550 5957 11586 5958
rect 11659 5954 11697 5962
rect 11763 5986 11848 5992
rect 11868 5991 11905 5992
rect 11763 5966 11771 5986
rect 11791 5985 11848 5986
rect 11791 5966 11820 5985
rect 11763 5965 11820 5966
rect 11841 5965 11848 5985
rect 11763 5958 11848 5965
rect 11867 5982 11905 5991
rect 11867 5962 11876 5982
rect 11896 5962 11905 5982
rect 11763 5957 11799 5958
rect 11867 5954 11905 5962
rect 11971 5986 12115 5992
rect 11971 5966 11979 5986
rect 11999 5966 12087 5986
rect 12107 5966 12115 5986
rect 11971 5958 12115 5966
rect 11971 5957 12007 5958
rect 12079 5957 12115 5958
rect 12181 5991 12218 5992
rect 12181 5990 12219 5991
rect 12181 5982 12245 5990
rect 12181 5962 12190 5982
rect 12210 5968 12245 5982
rect 12265 5968 12268 5988
rect 12210 5963 12268 5968
rect 12210 5962 12245 5963
rect 10795 5935 11211 5940
rect 10795 5934 11136 5935
rect 10739 5874 10770 5875
rect 10587 5844 10596 5864
rect 10616 5844 10624 5864
rect 10587 5834 10624 5844
rect 10683 5867 10770 5874
rect 10683 5864 10744 5867
rect 10683 5844 10692 5864
rect 10712 5847 10744 5864
rect 10765 5847 10770 5867
rect 10712 5844 10770 5847
rect 10683 5837 10770 5844
rect 10795 5864 10832 5934
rect 11098 5933 11135 5934
rect 11447 5925 11484 5954
rect 11448 5923 11484 5925
rect 11660 5923 11697 5954
rect 11448 5901 11697 5923
rect 11868 5922 11905 5954
rect 12181 5950 12245 5962
rect 12285 5924 12314 6102
rect 12682 6095 12709 6273
rect 12749 6235 12813 6247
rect 13089 6243 13126 6275
rect 13297 6274 13546 6296
rect 13297 6243 13334 6274
rect 13510 6272 13546 6274
rect 13510 6243 13547 6272
rect 13859 6263 13896 6264
rect 14162 6263 14199 6333
rect 14224 6353 14311 6360
rect 14224 6350 14282 6353
rect 14224 6330 14229 6350
rect 14250 6333 14282 6350
rect 14302 6333 14311 6353
rect 14250 6330 14311 6333
rect 14224 6323 14311 6330
rect 14370 6353 14407 6363
rect 14370 6333 14378 6353
rect 14398 6333 14407 6353
rect 14224 6322 14255 6323
rect 13858 6262 14199 6263
rect 13783 6257 14199 6262
rect 12749 6234 12784 6235
rect 12726 6229 12784 6234
rect 12726 6209 12729 6229
rect 12749 6215 12784 6229
rect 12804 6215 12813 6235
rect 12749 6207 12813 6215
rect 12775 6206 12813 6207
rect 12776 6205 12813 6206
rect 12879 6239 12915 6240
rect 12987 6239 13023 6240
rect 12879 6234 13023 6239
rect 12879 6231 12939 6234
rect 12879 6211 12887 6231
rect 12907 6213 12939 6231
rect 12966 6231 13023 6234
rect 12966 6213 12995 6231
rect 12907 6211 12995 6213
rect 13015 6211 13023 6231
rect 12879 6205 13023 6211
rect 13089 6235 13127 6243
rect 13195 6239 13231 6240
rect 13089 6215 13098 6235
rect 13118 6215 13127 6235
rect 13089 6206 13127 6215
rect 13146 6232 13231 6239
rect 13146 6212 13153 6232
rect 13174 6231 13231 6232
rect 13174 6212 13203 6231
rect 13146 6211 13203 6212
rect 13223 6211 13231 6231
rect 13089 6205 13126 6206
rect 13146 6205 13231 6211
rect 13297 6235 13335 6243
rect 13408 6239 13444 6240
rect 13297 6215 13306 6235
rect 13326 6215 13335 6235
rect 13297 6206 13335 6215
rect 13359 6231 13444 6239
rect 13359 6211 13416 6231
rect 13436 6211 13444 6231
rect 13297 6205 13334 6206
rect 13359 6205 13444 6211
rect 13510 6235 13548 6243
rect 13783 6237 13786 6257
rect 13806 6237 14199 6257
rect 14370 6254 14407 6333
rect 14437 6362 14468 6415
rect 14818 6413 14855 6414
rect 14817 6404 14856 6413
rect 14817 6386 14827 6404
rect 14845 6386 14856 6404
rect 15197 6402 15234 6406
rect 14729 6369 14776 6370
rect 14817 6369 14856 6386
rect 14729 6365 14856 6369
rect 14487 6362 14524 6363
rect 14437 6353 14524 6362
rect 14437 6333 14495 6353
rect 14515 6333 14524 6353
rect 14437 6323 14524 6333
rect 14583 6353 14620 6363
rect 14583 6333 14591 6353
rect 14611 6333 14620 6353
rect 14437 6322 14468 6323
rect 14432 6254 14542 6267
rect 14583 6254 14620 6333
rect 14729 6336 14739 6365
rect 14768 6336 14856 6365
rect 14729 6330 14856 6336
rect 14729 6326 14776 6330
rect 14814 6316 14856 6330
rect 14814 6298 14825 6316
rect 14843 6298 14856 6316
rect 14814 6293 14856 6298
rect 14815 6290 14856 6293
rect 15194 6397 15234 6402
rect 15194 6379 15206 6397
rect 15224 6379 15234 6397
rect 14815 6289 14852 6290
rect 14370 6252 14620 6254
rect 14370 6249 14471 6252
rect 13510 6215 13519 6235
rect 13539 6215 13548 6235
rect 14370 6230 14435 6249
rect 13510 6206 13548 6215
rect 14432 6222 14435 6230
rect 14464 6222 14471 6249
rect 14499 6225 14509 6252
rect 14538 6230 14620 6252
rect 14538 6225 14542 6230
rect 14499 6222 14542 6225
rect 14432 6208 14542 6222
rect 14808 6226 14855 6227
rect 14808 6217 14856 6226
rect 13510 6205 13547 6206
rect 12933 6184 12969 6205
rect 13359 6184 13390 6205
rect 14808 6199 14827 6217
rect 14845 6199 14856 6217
rect 14808 6197 14856 6199
rect 12766 6180 12866 6184
rect 12766 6176 12828 6180
rect 12766 6150 12773 6176
rect 12799 6154 12828 6176
rect 12854 6154 12866 6180
rect 12799 6150 12866 6154
rect 12766 6147 12866 6150
rect 12934 6147 12969 6184
rect 13031 6181 13390 6184
rect 13031 6176 13253 6181
rect 13031 6152 13044 6176
rect 13068 6157 13253 6176
rect 13277 6157 13390 6181
rect 13068 6152 13390 6157
rect 13031 6148 13390 6152
rect 13457 6176 13606 6184
rect 13457 6156 13468 6176
rect 13488 6156 13606 6176
rect 13457 6149 13606 6156
rect 13457 6148 13498 6149
rect 12781 6095 12818 6096
rect 12877 6095 12914 6096
rect 12933 6095 12969 6147
rect 12988 6095 13025 6096
rect 12681 6086 12819 6095
rect 12681 6066 12790 6086
rect 12810 6066 12819 6086
rect 12681 6059 12819 6066
rect 12877 6086 13025 6095
rect 12877 6066 12886 6086
rect 12906 6066 12996 6086
rect 13016 6066 13025 6086
rect 12681 6057 12777 6059
rect 12877 6056 13025 6066
rect 13084 6086 13121 6096
rect 13196 6095 13233 6096
rect 13177 6093 13233 6095
rect 13084 6066 13092 6086
rect 13112 6066 13121 6086
rect 12933 6055 12969 6056
rect 12781 5996 12818 5997
rect 13084 5996 13121 6066
rect 13146 6086 13233 6093
rect 13146 6083 13204 6086
rect 13146 6063 13151 6083
rect 13172 6066 13204 6083
rect 13224 6066 13233 6086
rect 13172 6063 13233 6066
rect 13146 6056 13233 6063
rect 13292 6086 13329 6096
rect 13292 6066 13300 6086
rect 13320 6066 13329 6086
rect 13146 6055 13177 6056
rect 12780 5995 13121 5996
rect 12705 5991 13121 5995
rect 12705 5990 13082 5991
rect 12705 5970 12708 5990
rect 12728 5974 13082 5990
rect 13102 5974 13121 5991
rect 12728 5970 13121 5974
rect 13292 5987 13329 6066
rect 13359 6095 13390 6148
rect 14170 6140 14208 6142
rect 14817 6140 14856 6197
rect 14170 6107 14856 6140
rect 13409 6095 13446 6096
rect 13359 6086 13446 6095
rect 13359 6066 13417 6086
rect 13437 6066 13446 6086
rect 13359 6056 13446 6066
rect 13505 6086 13542 6096
rect 13505 6066 13513 6086
rect 13533 6066 13542 6086
rect 13359 6055 13390 6056
rect 13354 5987 13464 6000
rect 13505 5987 13542 6066
rect 13292 5985 13542 5987
rect 13292 5982 13393 5985
rect 13292 5963 13357 5982
rect 13354 5955 13357 5963
rect 13386 5955 13393 5982
rect 13421 5958 13431 5985
rect 13460 5963 13542 5985
rect 13762 6019 13930 6020
rect 14170 6019 14208 6107
rect 14469 6105 14516 6107
rect 14816 6083 14856 6107
rect 13762 5996 14208 6019
rect 14434 6050 14545 6065
rect 14434 6048 14476 6050
rect 14434 6028 14441 6048
rect 14460 6028 14476 6048
rect 14434 6020 14476 6028
rect 14504 6048 14545 6050
rect 14504 6028 14518 6048
rect 14537 6028 14545 6048
rect 14817 6039 14856 6083
rect 14504 6020 14545 6028
rect 14434 6014 14545 6020
rect 13762 5993 14206 5996
rect 13762 5991 13930 5993
rect 13460 5958 13464 5963
rect 13421 5955 13464 5958
rect 13354 5941 13464 5955
rect 12144 5922 12314 5924
rect 11865 5915 12314 5922
rect 11529 5895 11640 5901
rect 11529 5887 11570 5895
rect 10947 5874 10983 5875
rect 10795 5844 10804 5864
rect 10824 5844 10832 5864
rect 10683 5835 10739 5837
rect 10683 5834 10720 5835
rect 10795 5834 10832 5844
rect 10891 5864 11039 5874
rect 11139 5871 11235 5873
rect 10891 5844 10900 5864
rect 10920 5844 11010 5864
rect 11030 5844 11039 5864
rect 10891 5835 11039 5844
rect 11097 5864 11235 5871
rect 11097 5844 11106 5864
rect 11126 5844 11235 5864
rect 11529 5867 11537 5887
rect 11556 5867 11570 5887
rect 11529 5865 11570 5867
rect 11598 5887 11640 5895
rect 11598 5867 11614 5887
rect 11633 5867 11640 5887
rect 11865 5888 11890 5915
rect 11921 5896 12314 5915
rect 11921 5888 11970 5896
rect 12144 5895 12314 5896
rect 11865 5886 11970 5888
rect 11598 5865 11640 5867
rect 11529 5850 11640 5865
rect 11097 5835 11235 5844
rect 10891 5834 10928 5835
rect 10947 5783 10983 5835
rect 11002 5834 11039 5835
rect 11098 5834 11135 5835
rect 10418 5781 10459 5782
rect 9840 5769 9881 5778
rect 10310 5774 10459 5781
rect 9840 5749 9880 5769
rect 9397 5739 9647 5741
rect 9397 5736 9498 5739
rect 7915 5679 7979 5691
rect 8255 5687 8292 5714
rect 8463 5687 8500 5718
rect 8676 5716 8712 5718
rect 9397 5717 9462 5736
rect 8676 5687 8713 5716
rect 9459 5709 9462 5717
rect 9491 5709 9498 5736
rect 9526 5712 9536 5739
rect 9565 5717 9647 5739
rect 9755 5739 9880 5749
rect 10310 5754 10428 5774
rect 10448 5754 10459 5774
rect 10310 5746 10459 5754
rect 10526 5778 10885 5782
rect 10526 5773 10848 5778
rect 10526 5749 10639 5773
rect 10663 5754 10848 5773
rect 10872 5754 10885 5778
rect 10663 5749 10885 5754
rect 10526 5746 10885 5749
rect 10947 5746 10982 5783
rect 11050 5780 11150 5783
rect 11050 5776 11117 5780
rect 11050 5750 11062 5776
rect 11088 5754 11117 5776
rect 11143 5754 11150 5780
rect 11088 5750 11150 5754
rect 11050 5746 11150 5750
rect 9755 5720 9763 5739
rect 9788 5720 9880 5739
rect 10526 5725 10557 5746
rect 10947 5725 10983 5746
rect 10369 5724 10406 5725
rect 10143 5721 10177 5722
rect 9565 5712 9569 5717
rect 9755 5713 9880 5720
rect 9526 5709 9569 5712
rect 9459 5695 9569 5709
rect 7915 5678 7950 5679
rect 7892 5673 7950 5678
rect 7892 5653 7895 5673
rect 7915 5659 7950 5673
rect 7970 5659 7979 5679
rect 7915 5651 7979 5659
rect 7941 5650 7979 5651
rect 7942 5649 7979 5650
rect 8045 5683 8081 5684
rect 8153 5683 8189 5684
rect 8045 5675 8189 5683
rect 8045 5655 8053 5675
rect 8073 5672 8161 5675
rect 8073 5655 8105 5672
rect 8125 5655 8161 5672
rect 8181 5655 8189 5675
rect 8045 5649 8189 5655
rect 8255 5679 8293 5687
rect 8361 5683 8397 5684
rect 8255 5659 8264 5679
rect 8284 5659 8293 5679
rect 8255 5650 8293 5659
rect 8312 5676 8397 5683
rect 8312 5656 8319 5676
rect 8340 5675 8397 5676
rect 8340 5656 8369 5675
rect 8312 5655 8369 5656
rect 8389 5655 8397 5675
rect 8255 5649 8292 5650
rect 8312 5649 8397 5655
rect 8463 5679 8501 5687
rect 8574 5683 8610 5684
rect 8463 5659 8472 5679
rect 8492 5659 8501 5679
rect 8463 5650 8501 5659
rect 8525 5675 8610 5683
rect 8525 5655 8582 5675
rect 8602 5655 8610 5675
rect 8463 5649 8500 5650
rect 8525 5649 8610 5655
rect 8676 5679 8714 5687
rect 8676 5659 8685 5679
rect 8705 5659 8714 5679
rect 8676 5650 8714 5659
rect 9840 5665 9880 5713
rect 10142 5712 10179 5721
rect 10142 5694 10151 5712
rect 10169 5694 10179 5712
rect 10142 5684 10179 5694
rect 10368 5715 10406 5724
rect 10368 5695 10377 5715
rect 10397 5695 10406 5715
rect 10368 5687 10406 5695
rect 10472 5719 10557 5725
rect 10582 5724 10619 5725
rect 10472 5699 10480 5719
rect 10500 5699 10557 5719
rect 10472 5691 10557 5699
rect 10581 5715 10619 5724
rect 10581 5695 10590 5715
rect 10610 5695 10619 5715
rect 10472 5690 10508 5691
rect 10581 5687 10619 5695
rect 10685 5719 10770 5725
rect 10790 5724 10827 5725
rect 10685 5699 10693 5719
rect 10713 5718 10770 5719
rect 10713 5699 10742 5718
rect 10685 5698 10742 5699
rect 10763 5698 10770 5718
rect 10685 5691 10770 5698
rect 10789 5715 10827 5724
rect 10789 5695 10798 5715
rect 10818 5695 10827 5715
rect 10685 5690 10721 5691
rect 10789 5687 10827 5695
rect 10893 5719 11037 5725
rect 10893 5699 10901 5719
rect 10921 5718 11009 5719
rect 10921 5699 10952 5718
rect 10893 5698 10952 5699
rect 10977 5699 11009 5718
rect 11029 5699 11037 5719
rect 10977 5698 11037 5699
rect 10893 5691 11037 5698
rect 10893 5690 10929 5691
rect 11001 5690 11037 5691
rect 11103 5724 11140 5725
rect 11103 5723 11141 5724
rect 11103 5715 11167 5723
rect 11103 5695 11112 5715
rect 11132 5701 11167 5715
rect 11187 5701 11190 5721
rect 11132 5696 11190 5701
rect 11132 5695 11167 5696
rect 8676 5649 8713 5650
rect 8099 5628 8135 5649
rect 8525 5628 8556 5649
rect 9840 5647 9851 5665
rect 9869 5647 9880 5665
rect 9840 5639 9880 5647
rect 10143 5656 10177 5684
rect 10369 5658 10406 5687
rect 10370 5656 10406 5658
rect 10582 5656 10619 5687
rect 10143 5655 10315 5656
rect 9841 5638 9878 5639
rect 7932 5624 8032 5628
rect 7932 5620 7994 5624
rect 7932 5594 7939 5620
rect 7965 5598 7994 5620
rect 8020 5598 8032 5624
rect 7965 5594 8032 5598
rect 7932 5591 8032 5594
rect 8100 5591 8135 5628
rect 8197 5625 8556 5628
rect 8197 5620 8419 5625
rect 8197 5596 8210 5620
rect 8234 5601 8419 5620
rect 8443 5601 8556 5625
rect 8234 5596 8556 5601
rect 8197 5592 8556 5596
rect 8623 5620 8772 5628
rect 8623 5600 8634 5620
rect 8654 5600 8772 5620
rect 8623 5593 8772 5600
rect 10143 5623 10329 5655
rect 10370 5634 10619 5656
rect 10790 5655 10827 5687
rect 11103 5683 11167 5695
rect 11207 5657 11234 5835
rect 13762 5813 13789 5991
rect 13829 5953 13893 5965
rect 14169 5961 14206 5993
rect 14377 5992 14626 6014
rect 14377 5961 14414 5992
rect 14590 5990 14626 5992
rect 14590 5961 14627 5990
rect 13829 5952 13864 5953
rect 13806 5947 13864 5952
rect 13806 5927 13809 5947
rect 13829 5933 13864 5947
rect 13884 5933 13893 5953
rect 13829 5925 13893 5933
rect 13855 5924 13893 5925
rect 13856 5923 13893 5924
rect 13959 5957 13995 5958
rect 14067 5957 14103 5958
rect 13959 5952 14103 5957
rect 13959 5949 14021 5952
rect 13959 5929 13967 5949
rect 13987 5932 14021 5949
rect 14044 5949 14103 5952
rect 14044 5932 14075 5949
rect 13987 5929 14075 5932
rect 14095 5929 14103 5949
rect 13959 5923 14103 5929
rect 14169 5953 14207 5961
rect 14275 5957 14311 5958
rect 14169 5933 14178 5953
rect 14198 5933 14207 5953
rect 14169 5924 14207 5933
rect 14226 5950 14311 5957
rect 14226 5930 14233 5950
rect 14254 5949 14311 5950
rect 14254 5930 14283 5949
rect 14226 5929 14283 5930
rect 14303 5929 14311 5949
rect 14169 5923 14206 5924
rect 14226 5923 14311 5929
rect 14377 5953 14415 5961
rect 14488 5957 14524 5958
rect 14377 5933 14386 5953
rect 14406 5933 14415 5953
rect 14377 5924 14415 5933
rect 14439 5949 14524 5957
rect 14439 5929 14496 5949
rect 14516 5929 14524 5949
rect 14377 5923 14414 5924
rect 14439 5923 14524 5929
rect 14590 5953 14628 5961
rect 14590 5933 14599 5953
rect 14619 5933 14628 5953
rect 14590 5924 14628 5933
rect 14590 5923 14627 5924
rect 14013 5902 14049 5923
rect 14439 5902 14470 5923
rect 13846 5898 13946 5902
rect 13846 5894 13908 5898
rect 13846 5868 13853 5894
rect 13879 5872 13908 5894
rect 13934 5872 13946 5898
rect 13879 5868 13946 5872
rect 13846 5865 13946 5868
rect 14014 5865 14049 5902
rect 14111 5899 14470 5902
rect 14111 5894 14333 5899
rect 14111 5870 14124 5894
rect 14148 5875 14333 5894
rect 14357 5875 14470 5899
rect 14148 5870 14470 5875
rect 14111 5866 14470 5870
rect 14537 5894 14686 5902
rect 14537 5874 14548 5894
rect 14568 5874 14686 5894
rect 14537 5867 14686 5874
rect 14537 5866 14578 5867
rect 13861 5813 13898 5814
rect 13957 5813 13994 5814
rect 14013 5813 14049 5865
rect 14068 5813 14105 5814
rect 13761 5804 13899 5813
rect 13761 5784 13870 5804
rect 13890 5784 13899 5804
rect 13761 5777 13899 5784
rect 13957 5804 14105 5813
rect 13957 5784 13966 5804
rect 13986 5784 14076 5804
rect 14096 5784 14105 5804
rect 13761 5775 13857 5777
rect 13957 5774 14105 5784
rect 14164 5804 14201 5814
rect 14276 5813 14313 5814
rect 14257 5811 14313 5813
rect 14164 5784 14172 5804
rect 14192 5784 14201 5804
rect 14013 5773 14049 5774
rect 11390 5731 11500 5745
rect 11390 5728 11433 5731
rect 11390 5723 11394 5728
rect 11066 5655 11234 5657
rect 10790 5649 11234 5655
rect 9212 5597 9726 5598
rect 8623 5592 8664 5593
rect 7947 5539 7984 5540
rect 8043 5539 8080 5540
rect 8099 5539 8135 5591
rect 8154 5539 8191 5540
rect 7847 5530 7985 5539
rect 7847 5510 7956 5530
rect 7976 5510 7985 5530
rect 7847 5503 7985 5510
rect 8043 5530 8191 5539
rect 8043 5510 8052 5530
rect 8072 5510 8162 5530
rect 8182 5510 8191 5530
rect 7847 5501 7943 5503
rect 8043 5500 8191 5510
rect 8250 5530 8287 5540
rect 8362 5539 8399 5540
rect 8343 5537 8399 5539
rect 8250 5510 8258 5530
rect 8278 5510 8287 5530
rect 8099 5499 8135 5500
rect 7029 5447 7197 5449
rect 6751 5441 7197 5447
rect 5819 5417 6235 5422
rect 6414 5420 6525 5426
rect 5819 5416 6160 5417
rect 5763 5356 5794 5357
rect 5611 5326 5620 5346
rect 5640 5326 5648 5346
rect 5611 5316 5648 5326
rect 5707 5349 5794 5356
rect 5707 5346 5768 5349
rect 5707 5326 5716 5346
rect 5736 5329 5768 5346
rect 5789 5329 5794 5349
rect 5736 5326 5794 5329
rect 5707 5319 5794 5326
rect 5819 5346 5856 5416
rect 6122 5415 6159 5416
rect 6414 5412 6455 5420
rect 6414 5392 6422 5412
rect 6441 5392 6455 5412
rect 6414 5390 6455 5392
rect 6483 5412 6525 5420
rect 6483 5392 6499 5412
rect 6518 5392 6525 5412
rect 6751 5419 6757 5441
rect 6783 5421 7197 5441
rect 7947 5440 7984 5441
rect 8250 5440 8287 5510
rect 8312 5530 8399 5537
rect 8312 5527 8370 5530
rect 8312 5507 8317 5527
rect 8338 5510 8370 5527
rect 8390 5510 8399 5530
rect 8338 5507 8399 5510
rect 8312 5500 8399 5507
rect 8458 5530 8495 5540
rect 8458 5510 8466 5530
rect 8486 5510 8495 5530
rect 8312 5499 8343 5500
rect 7946 5439 8287 5440
rect 6783 5419 6792 5421
rect 7029 5420 7197 5421
rect 7871 5434 8287 5439
rect 6751 5410 6792 5419
rect 7871 5414 7874 5434
rect 7894 5414 8287 5434
rect 8458 5431 8495 5510
rect 8525 5539 8556 5592
rect 9193 5581 9726 5597
rect 10143 5591 10177 5623
rect 10139 5582 10177 5591
rect 9193 5570 9725 5581
rect 9844 5572 9881 5576
rect 8575 5539 8612 5540
rect 8525 5530 8612 5539
rect 8525 5510 8583 5530
rect 8603 5510 8612 5530
rect 8525 5500 8612 5510
rect 8671 5530 8708 5540
rect 8671 5510 8679 5530
rect 8699 5510 8708 5530
rect 8525 5499 8556 5500
rect 8520 5431 8630 5444
rect 8671 5431 8708 5510
rect 8458 5429 8708 5431
rect 8458 5426 8559 5429
rect 8458 5407 8523 5426
rect 8520 5399 8523 5407
rect 8552 5399 8559 5426
rect 8587 5402 8597 5429
rect 8626 5407 8708 5429
rect 8786 5501 8954 5502
rect 9193 5501 9231 5570
rect 8786 5481 9231 5501
rect 9458 5532 9569 5547
rect 9458 5530 9500 5532
rect 9458 5510 9465 5530
rect 9484 5510 9500 5530
rect 9458 5502 9500 5510
rect 9528 5530 9569 5532
rect 9528 5510 9542 5530
rect 9561 5510 9569 5530
rect 9528 5502 9569 5510
rect 9458 5496 9569 5502
rect 9691 5507 9725 5570
rect 9843 5566 9881 5572
rect 9843 5548 9853 5566
rect 9871 5548 9881 5566
rect 10139 5564 10149 5582
rect 10167 5564 10177 5582
rect 10139 5558 10177 5564
rect 10295 5560 10329 5623
rect 10451 5628 10562 5634
rect 10451 5620 10492 5628
rect 10451 5600 10459 5620
rect 10478 5600 10492 5620
rect 10451 5598 10492 5600
rect 10520 5620 10562 5628
rect 10520 5600 10536 5620
rect 10555 5600 10562 5620
rect 10520 5598 10562 5600
rect 10451 5583 10562 5598
rect 10789 5629 11234 5649
rect 10789 5560 10827 5629
rect 11066 5628 11234 5629
rect 11312 5701 11394 5723
rect 11423 5701 11433 5728
rect 11461 5704 11468 5731
rect 11497 5723 11500 5731
rect 13495 5740 13606 5755
rect 13495 5738 13537 5740
rect 11497 5704 11562 5723
rect 11461 5701 11562 5704
rect 11312 5699 11562 5701
rect 11312 5620 11349 5699
rect 11390 5686 11500 5699
rect 11464 5630 11495 5631
rect 11312 5600 11321 5620
rect 11341 5600 11349 5620
rect 11312 5590 11349 5600
rect 11408 5620 11495 5630
rect 11408 5600 11417 5620
rect 11437 5600 11495 5620
rect 11408 5591 11495 5600
rect 11408 5590 11445 5591
rect 10139 5554 10176 5558
rect 10295 5549 10827 5560
rect 9843 5539 9881 5548
rect 9843 5507 9877 5539
rect 10294 5533 10827 5549
rect 11464 5538 11495 5591
rect 11525 5620 11562 5699
rect 11733 5709 12126 5716
rect 11733 5692 11741 5709
rect 11773 5696 12126 5709
rect 12146 5696 12149 5716
rect 13228 5711 13269 5720
rect 11773 5692 12149 5696
rect 11733 5691 12149 5692
rect 12823 5709 12991 5710
rect 13228 5709 13237 5711
rect 11733 5690 12074 5691
rect 11677 5630 11708 5631
rect 11525 5600 11534 5620
rect 11554 5600 11562 5620
rect 11525 5590 11562 5600
rect 11621 5623 11708 5630
rect 11621 5620 11682 5623
rect 11621 5600 11630 5620
rect 11650 5603 11682 5620
rect 11703 5603 11708 5623
rect 11650 5600 11708 5603
rect 11621 5593 11708 5600
rect 11733 5620 11770 5690
rect 12036 5689 12073 5690
rect 12823 5689 13237 5709
rect 13263 5689 13269 5711
rect 13495 5718 13502 5738
rect 13521 5718 13537 5738
rect 13495 5710 13537 5718
rect 13565 5738 13606 5740
rect 13565 5718 13579 5738
rect 13598 5718 13606 5738
rect 13565 5710 13606 5718
rect 13861 5714 13898 5715
rect 14164 5714 14201 5784
rect 14226 5804 14313 5811
rect 14226 5801 14284 5804
rect 14226 5781 14231 5801
rect 14252 5784 14284 5801
rect 14304 5784 14313 5804
rect 14252 5781 14313 5784
rect 14226 5774 14313 5781
rect 14372 5804 14409 5814
rect 14372 5784 14380 5804
rect 14400 5784 14409 5804
rect 14226 5773 14257 5774
rect 13860 5713 14201 5714
rect 13495 5704 13606 5710
rect 13785 5708 14201 5713
rect 12823 5683 13269 5689
rect 12823 5681 12991 5683
rect 11885 5630 11921 5631
rect 11733 5600 11742 5620
rect 11762 5600 11770 5620
rect 11621 5591 11677 5593
rect 11621 5590 11658 5591
rect 11733 5590 11770 5600
rect 11829 5620 11977 5630
rect 12077 5627 12173 5629
rect 11829 5600 11838 5620
rect 11858 5615 11948 5620
rect 11858 5600 11893 5615
rect 11829 5591 11893 5600
rect 11829 5590 11866 5591
rect 11885 5574 11893 5591
rect 11914 5600 11948 5615
rect 11968 5600 11977 5620
rect 11914 5591 11977 5600
rect 12035 5620 12173 5627
rect 12035 5600 12044 5620
rect 12064 5600 12173 5620
rect 12035 5591 12173 5600
rect 11914 5574 11921 5591
rect 11940 5590 11977 5591
rect 12036 5590 12073 5591
rect 11885 5539 11921 5574
rect 11356 5537 11397 5538
rect 10294 5532 10808 5533
rect 8786 5475 9230 5481
rect 8786 5473 8954 5475
rect 8626 5402 8630 5407
rect 8587 5399 8630 5402
rect 6483 5390 6525 5392
rect 6414 5375 6525 5390
rect 7610 5381 7658 5395
rect 8520 5385 8630 5399
rect 5971 5356 6007 5357
rect 5819 5326 5828 5346
rect 5848 5326 5856 5346
rect 5707 5317 5763 5319
rect 5707 5316 5744 5317
rect 5819 5316 5856 5326
rect 5915 5346 6063 5356
rect 6163 5353 6259 5355
rect 5915 5326 5924 5346
rect 5944 5326 6034 5346
rect 6054 5326 6063 5346
rect 5915 5317 6063 5326
rect 6121 5346 6259 5353
rect 6121 5326 6130 5346
rect 6150 5326 6259 5346
rect 6121 5317 6259 5326
rect 7610 5341 7623 5381
rect 7650 5341 7658 5381
rect 7610 5323 7658 5341
rect 5915 5316 5952 5317
rect 5971 5265 6007 5317
rect 6026 5316 6063 5317
rect 6122 5316 6159 5317
rect 5442 5263 5483 5264
rect 5334 5256 5483 5263
rect 5334 5236 5452 5256
rect 5472 5236 5483 5256
rect 5334 5228 5483 5236
rect 5550 5260 5909 5264
rect 5550 5255 5872 5260
rect 5550 5231 5663 5255
rect 5687 5236 5872 5255
rect 5896 5236 5909 5260
rect 5687 5231 5909 5236
rect 5550 5228 5909 5231
rect 5971 5228 6006 5265
rect 6074 5262 6174 5265
rect 6074 5258 6141 5262
rect 6074 5232 6086 5258
rect 6112 5236 6141 5258
rect 6167 5236 6174 5262
rect 6112 5232 6174 5236
rect 6074 5228 6174 5232
rect 5550 5207 5581 5228
rect 5971 5207 6007 5228
rect 5393 5206 5430 5207
rect 5392 5197 5430 5206
rect 5392 5177 5401 5197
rect 5421 5177 5430 5197
rect 5392 5169 5430 5177
rect 5496 5201 5581 5207
rect 5606 5206 5643 5207
rect 5496 5181 5504 5201
rect 5524 5181 5581 5201
rect 5496 5173 5581 5181
rect 5605 5197 5643 5206
rect 5605 5177 5614 5197
rect 5634 5177 5643 5197
rect 5496 5172 5532 5173
rect 5605 5169 5643 5177
rect 5709 5201 5794 5207
rect 5814 5206 5851 5207
rect 5709 5181 5717 5201
rect 5737 5200 5794 5201
rect 5737 5181 5766 5200
rect 5709 5180 5766 5181
rect 5787 5180 5794 5200
rect 5709 5173 5794 5180
rect 5813 5197 5851 5206
rect 5813 5177 5822 5197
rect 5842 5177 5851 5197
rect 5709 5172 5745 5173
rect 5813 5169 5851 5177
rect 5917 5201 6061 5207
rect 5917 5181 5925 5201
rect 5945 5198 6033 5201
rect 5945 5181 5976 5198
rect 5917 5178 5976 5181
rect 5999 5181 6033 5198
rect 6053 5181 6061 5201
rect 5999 5178 6061 5181
rect 5917 5173 6061 5178
rect 5917 5172 5953 5173
rect 6025 5172 6061 5173
rect 6127 5206 6164 5207
rect 6127 5205 6165 5206
rect 6127 5197 6191 5205
rect 6127 5177 6136 5197
rect 6156 5183 6191 5197
rect 6211 5183 6214 5203
rect 6156 5178 6214 5183
rect 6156 5177 6191 5178
rect 5393 5140 5430 5169
rect 5394 5138 5430 5140
rect 5606 5138 5643 5169
rect 5394 5116 5643 5138
rect 5814 5137 5851 5169
rect 6127 5165 6191 5177
rect 6231 5139 6258 5317
rect 7605 5216 7658 5323
rect 8786 5295 8813 5473
rect 8853 5435 8917 5447
rect 9193 5443 9230 5475
rect 9401 5474 9650 5496
rect 9691 5475 9877 5507
rect 11248 5530 11397 5537
rect 11248 5510 11366 5530
rect 11386 5510 11397 5530
rect 11248 5502 11397 5510
rect 11464 5534 11823 5538
rect 11464 5529 11786 5534
rect 11464 5505 11577 5529
rect 11601 5510 11786 5529
rect 11810 5510 11823 5534
rect 11601 5505 11823 5510
rect 11464 5502 11823 5505
rect 11885 5502 11920 5539
rect 11988 5536 12088 5539
rect 11988 5532 12055 5536
rect 11988 5506 12000 5532
rect 12026 5510 12055 5532
rect 12081 5510 12088 5536
rect 12026 5506 12088 5510
rect 11988 5502 12088 5506
rect 10142 5491 10179 5492
rect 9705 5474 9877 5475
rect 9401 5443 9438 5474
rect 9614 5472 9650 5474
rect 9614 5443 9651 5472
rect 9843 5446 9877 5474
rect 10140 5483 10180 5491
rect 10140 5465 10151 5483
rect 10169 5465 10180 5483
rect 11464 5481 11495 5502
rect 11885 5481 11921 5502
rect 11307 5480 11344 5481
rect 8853 5434 8888 5435
rect 8830 5429 8888 5434
rect 8830 5409 8833 5429
rect 8853 5415 8888 5429
rect 8908 5415 8917 5435
rect 8853 5407 8917 5415
rect 8879 5406 8917 5407
rect 8880 5405 8917 5406
rect 8983 5439 9019 5440
rect 9091 5439 9127 5440
rect 8983 5432 9127 5439
rect 8983 5431 9043 5432
rect 8983 5411 8991 5431
rect 9011 5412 9043 5431
rect 9068 5431 9127 5432
rect 9068 5412 9099 5431
rect 9011 5411 9099 5412
rect 9119 5411 9127 5431
rect 8983 5405 9127 5411
rect 9193 5435 9231 5443
rect 9299 5439 9335 5440
rect 9193 5415 9202 5435
rect 9222 5415 9231 5435
rect 9193 5406 9231 5415
rect 9250 5432 9335 5439
rect 9250 5412 9257 5432
rect 9278 5431 9335 5432
rect 9278 5412 9307 5431
rect 9250 5411 9307 5412
rect 9327 5411 9335 5431
rect 9193 5405 9230 5406
rect 9250 5405 9335 5411
rect 9401 5435 9439 5443
rect 9512 5439 9548 5440
rect 9401 5415 9410 5435
rect 9430 5415 9439 5435
rect 9401 5406 9439 5415
rect 9463 5431 9548 5439
rect 9463 5411 9520 5431
rect 9540 5411 9548 5431
rect 9401 5405 9438 5406
rect 9463 5405 9548 5411
rect 9614 5435 9652 5443
rect 9614 5415 9623 5435
rect 9643 5415 9652 5435
rect 9614 5406 9652 5415
rect 9841 5436 9878 5446
rect 9841 5418 9851 5436
rect 9869 5418 9878 5436
rect 9841 5409 9878 5418
rect 10140 5417 10180 5465
rect 11306 5471 11344 5480
rect 11306 5451 11315 5471
rect 11335 5451 11344 5471
rect 11306 5443 11344 5451
rect 11410 5475 11495 5481
rect 11520 5480 11557 5481
rect 11410 5455 11418 5475
rect 11438 5455 11495 5475
rect 11410 5447 11495 5455
rect 11519 5471 11557 5480
rect 11519 5451 11528 5471
rect 11548 5451 11557 5471
rect 11410 5446 11446 5447
rect 11519 5443 11557 5451
rect 11623 5475 11708 5481
rect 11728 5480 11765 5481
rect 11623 5455 11631 5475
rect 11651 5474 11708 5475
rect 11651 5455 11680 5474
rect 11623 5454 11680 5455
rect 11701 5454 11708 5474
rect 11623 5447 11708 5454
rect 11727 5471 11765 5480
rect 11727 5451 11736 5471
rect 11756 5451 11765 5471
rect 11623 5446 11659 5447
rect 11727 5443 11765 5451
rect 11831 5475 11975 5481
rect 11831 5455 11839 5475
rect 11859 5455 11947 5475
rect 11967 5455 11975 5475
rect 11831 5447 11975 5455
rect 11831 5446 11867 5447
rect 11939 5446 11975 5447
rect 12041 5480 12078 5481
rect 12041 5479 12079 5480
rect 12041 5471 12105 5479
rect 12041 5451 12050 5471
rect 12070 5457 12105 5471
rect 12125 5457 12128 5477
rect 12070 5452 12128 5457
rect 12070 5451 12105 5452
rect 10451 5421 10561 5435
rect 10451 5418 10494 5421
rect 10140 5410 10265 5417
rect 10451 5413 10455 5418
rect 9843 5408 9877 5409
rect 9614 5405 9651 5406
rect 9037 5384 9073 5405
rect 9463 5384 9494 5405
rect 10140 5391 10232 5410
rect 10257 5391 10265 5410
rect 8870 5380 8970 5384
rect 8870 5376 8932 5380
rect 8870 5350 8877 5376
rect 8903 5354 8932 5376
rect 8958 5354 8970 5380
rect 8903 5350 8970 5354
rect 8870 5347 8970 5350
rect 9038 5347 9073 5384
rect 9135 5381 9494 5384
rect 9135 5376 9357 5381
rect 9135 5352 9148 5376
rect 9172 5357 9357 5376
rect 9381 5357 9494 5381
rect 9172 5352 9494 5357
rect 9135 5348 9494 5352
rect 9561 5376 9710 5384
rect 9561 5356 9572 5376
rect 9592 5356 9710 5376
rect 10140 5381 10265 5391
rect 10373 5391 10455 5413
rect 10484 5391 10494 5418
rect 10522 5394 10529 5421
rect 10558 5413 10561 5421
rect 11307 5414 11344 5443
rect 10558 5394 10623 5413
rect 11308 5412 11344 5414
rect 11520 5412 11557 5443
rect 11728 5416 11765 5443
rect 12041 5439 12105 5451
rect 10522 5391 10623 5394
rect 10373 5389 10623 5391
rect 10140 5361 10180 5381
rect 9561 5349 9710 5356
rect 10139 5352 10180 5361
rect 9561 5348 9602 5349
rect 8885 5295 8922 5296
rect 8981 5295 9018 5296
rect 9037 5295 9073 5347
rect 9092 5295 9129 5296
rect 8785 5286 8923 5295
rect 8785 5266 8894 5286
rect 8914 5266 8923 5286
rect 8411 5246 8522 5261
rect 8785 5259 8923 5266
rect 8981 5286 9129 5295
rect 8981 5266 8990 5286
rect 9010 5266 9100 5286
rect 9120 5266 9129 5286
rect 8785 5257 8881 5259
rect 8981 5256 9129 5266
rect 9188 5286 9225 5296
rect 9300 5295 9337 5296
rect 9281 5293 9337 5295
rect 9188 5266 9196 5286
rect 9216 5266 9225 5286
rect 9037 5255 9073 5256
rect 8411 5244 8453 5246
rect 8411 5224 8418 5244
rect 8437 5224 8453 5244
rect 8411 5216 8453 5224
rect 8481 5244 8522 5246
rect 8481 5224 8495 5244
rect 8514 5224 8522 5244
rect 8481 5216 8522 5224
rect 7605 5215 7907 5216
rect 6524 5194 6634 5208
rect 6524 5191 6567 5194
rect 6524 5186 6528 5191
rect 6090 5137 6258 5139
rect 5814 5134 6258 5137
rect 5475 5110 5586 5116
rect 5475 5102 5516 5110
rect 3458 5022 3607 5029
rect 4139 5032 4177 5034
rect 4787 5032 4829 5051
rect 3458 5021 3499 5022
rect 2934 5016 2970 5020
rect 2934 4987 2971 5016
rect 2782 4968 2819 4969
rect 2878 4968 2915 4969
rect 2934 4968 2970 4987
rect 2989 4968 3026 4969
rect 2682 4959 2820 4968
rect 2682 4939 2791 4959
rect 2811 4939 2820 4959
rect 2682 4932 2820 4939
rect 2878 4959 3026 4968
rect 2878 4939 2887 4959
rect 2907 4939 2997 4959
rect 3017 4939 3026 4959
rect 2682 4930 2778 4932
rect 2878 4929 3026 4939
rect 3085 4959 3122 4969
rect 3197 4968 3234 4969
rect 3178 4966 3234 4968
rect 3085 4939 3093 4959
rect 3113 4939 3122 4959
rect 2934 4928 2970 4929
rect 2782 4869 2819 4870
rect 3085 4869 3122 4939
rect 3147 4959 3234 4966
rect 3147 4956 3205 4959
rect 3147 4936 3152 4956
rect 3173 4939 3205 4956
rect 3225 4939 3234 4959
rect 3173 4936 3234 4939
rect 3147 4929 3234 4936
rect 3293 4959 3330 4969
rect 3293 4939 3301 4959
rect 3321 4939 3330 4959
rect 3147 4928 3178 4929
rect 2781 4868 3122 4869
rect 2706 4863 3122 4868
rect 2331 4836 2384 4844
rect 2706 4843 2709 4863
rect 2729 4843 3122 4863
rect 3293 4860 3330 4939
rect 3360 4968 3391 5021
rect 4139 5009 4829 5032
rect 5164 5047 5203 5091
rect 5475 5082 5483 5102
rect 5502 5082 5516 5102
rect 5475 5080 5516 5082
rect 5544 5102 5586 5110
rect 5544 5082 5560 5102
rect 5579 5082 5586 5102
rect 5544 5081 5586 5082
rect 5812 5111 6258 5134
rect 5544 5080 5587 5081
rect 5475 5061 5587 5080
rect 5164 5023 5204 5047
rect 5504 5023 5551 5024
rect 5812 5023 5850 5111
rect 6090 5110 6258 5111
rect 6446 5164 6528 5186
rect 6557 5164 6567 5191
rect 6595 5167 6602 5194
rect 6631 5186 6634 5194
rect 7605 5189 8183 5215
rect 8411 5210 8522 5216
rect 7605 5187 7907 5189
rect 7605 5186 7791 5187
rect 6631 5167 6696 5186
rect 6595 5164 6696 5167
rect 6446 5162 6696 5164
rect 6446 5083 6483 5162
rect 6524 5149 6634 5162
rect 6598 5093 6629 5094
rect 6446 5063 6455 5083
rect 6475 5063 6483 5083
rect 6446 5053 6483 5063
rect 6542 5083 6629 5093
rect 6542 5063 6551 5083
rect 6571 5063 6629 5083
rect 6542 5054 6629 5063
rect 6542 5053 6579 5054
rect 5164 5013 5850 5023
rect 4139 4999 4825 5009
rect 3410 4968 3447 4969
rect 3360 4959 3447 4968
rect 3360 4939 3418 4959
rect 3438 4939 3447 4959
rect 3360 4929 3447 4939
rect 3506 4959 3543 4969
rect 3506 4939 3514 4959
rect 3534 4939 3543 4959
rect 3360 4928 3391 4929
rect 3355 4860 3465 4873
rect 3506 4860 3543 4939
rect 3293 4858 3543 4860
rect 3293 4855 3394 4858
rect 3293 4836 3358 4855
rect 2198 4835 2384 4836
rect 2082 4833 2384 4835
rect 1467 4806 1578 4812
rect 1806 4807 2384 4833
rect 3355 4828 3358 4836
rect 3387 4828 3394 4855
rect 3422 4831 3432 4858
rect 3461 4836 3543 4858
rect 3731 4911 3899 4912
rect 4139 4911 4177 4999
rect 4438 4998 4485 4999
rect 4785 4975 4825 4999
rect 4402 4942 4514 4961
rect 4402 4941 4445 4942
rect 3731 4888 4177 4911
rect 4403 4940 4445 4941
rect 4403 4920 4410 4940
rect 4429 4920 4445 4940
rect 4403 4912 4445 4920
rect 4473 4940 4514 4942
rect 4473 4920 4487 4940
rect 4506 4920 4514 4940
rect 4786 4931 4825 4975
rect 5160 4990 5850 5013
rect 6598 5001 6629 5054
rect 6659 5083 6696 5162
rect 6867 5159 7260 5179
rect 7280 5159 7283 5179
rect 7605 5178 7658 5186
rect 6867 5154 7283 5159
rect 6867 5153 7208 5154
rect 6811 5093 6842 5094
rect 6659 5063 6668 5083
rect 6688 5063 6696 5083
rect 6659 5053 6696 5063
rect 6755 5086 6842 5093
rect 6755 5083 6816 5086
rect 6755 5063 6764 5083
rect 6784 5066 6816 5083
rect 6837 5066 6842 5086
rect 6784 5063 6842 5066
rect 6755 5056 6842 5063
rect 6867 5083 6904 5153
rect 7170 5152 7207 5153
rect 7019 5093 7055 5094
rect 6867 5063 6876 5083
rect 6896 5063 6904 5083
rect 6755 5054 6811 5056
rect 6755 5053 6792 5054
rect 6867 5053 6904 5063
rect 6963 5083 7111 5093
rect 7211 5090 7307 5092
rect 6963 5063 6972 5083
rect 6992 5063 7082 5083
rect 7102 5063 7111 5083
rect 6963 5054 7111 5063
rect 7169 5083 7307 5090
rect 7169 5063 7178 5083
rect 7198 5063 7307 5083
rect 7169 5054 7307 5063
rect 6963 5053 7000 5054
rect 7019 5002 7055 5054
rect 7074 5053 7111 5054
rect 7170 5053 7207 5054
rect 6490 5000 6531 5001
rect 5160 4971 5202 4990
rect 5812 4988 5850 4990
rect 6382 4993 6531 5000
rect 4473 4912 4514 4920
rect 4403 4906 4514 4912
rect 3731 4885 4175 4888
rect 3731 4883 3899 4885
rect 3461 4831 3465 4836
rect 3422 4828 3465 4831
rect 3355 4814 3465 4828
rect 2082 4806 2384 4807
rect 1467 4798 1508 4806
rect 1467 4778 1475 4798
rect 1494 4778 1508 4798
rect 1467 4776 1508 4778
rect 1536 4798 1578 4806
rect 1536 4778 1552 4798
rect 1571 4778 1578 4798
rect 1536 4776 1578 4778
rect 916 4766 952 4767
rect 764 4736 773 4756
rect 793 4736 801 4756
rect 652 4727 708 4729
rect 652 4726 689 4727
rect 764 4726 801 4736
rect 860 4756 1008 4766
rect 1108 4763 1204 4765
rect 860 4736 869 4756
rect 889 4736 979 4756
rect 999 4736 1008 4756
rect 860 4727 1008 4736
rect 1066 4756 1204 4763
rect 1467 4761 1578 4776
rect 1066 4736 1075 4756
rect 1095 4736 1204 4756
rect 1066 4727 1204 4736
rect 860 4726 897 4727
rect 916 4675 952 4727
rect 971 4726 1008 4727
rect 1067 4726 1104 4727
rect 387 4673 428 4674
rect 279 4666 428 4673
rect 279 4646 397 4666
rect 417 4646 428 4666
rect 279 4638 428 4646
rect 495 4670 854 4674
rect 495 4665 817 4670
rect 495 4641 608 4665
rect 632 4646 817 4665
rect 841 4646 854 4670
rect 632 4641 854 4646
rect 495 4638 854 4641
rect 916 4638 951 4675
rect 1019 4672 1119 4675
rect 1019 4668 1086 4672
rect 1019 4642 1031 4668
rect 1057 4646 1086 4668
rect 1112 4646 1119 4672
rect 1057 4642 1119 4646
rect 1019 4638 1119 4642
rect 495 4617 526 4638
rect 916 4617 952 4638
rect 338 4616 375 4617
rect 112 4613 146 4614
rect 111 4604 148 4613
rect 111 4586 120 4604
rect 138 4586 148 4604
rect 111 4576 148 4586
rect 337 4607 375 4616
rect 337 4587 346 4607
rect 366 4587 375 4607
rect 337 4579 375 4587
rect 441 4611 526 4617
rect 551 4616 588 4617
rect 441 4591 449 4611
rect 469 4591 526 4611
rect 441 4583 526 4591
rect 550 4607 588 4616
rect 550 4587 559 4607
rect 579 4587 588 4607
rect 441 4582 477 4583
rect 550 4579 588 4587
rect 654 4611 739 4617
rect 759 4616 796 4617
rect 654 4591 662 4611
rect 682 4610 739 4611
rect 682 4591 711 4610
rect 654 4590 711 4591
rect 732 4590 739 4610
rect 654 4583 739 4590
rect 758 4607 796 4616
rect 758 4587 767 4607
rect 787 4587 796 4607
rect 654 4582 690 4583
rect 758 4579 796 4587
rect 862 4611 1006 4617
rect 862 4591 870 4611
rect 890 4610 978 4611
rect 890 4591 921 4610
rect 862 4590 921 4591
rect 946 4591 978 4610
rect 998 4591 1006 4611
rect 946 4590 1006 4591
rect 862 4583 1006 4590
rect 862 4582 898 4583
rect 970 4582 1006 4583
rect 1072 4616 1109 4617
rect 1072 4615 1110 4616
rect 1072 4607 1136 4615
rect 1072 4587 1081 4607
rect 1101 4593 1136 4607
rect 1156 4593 1159 4613
rect 1101 4588 1159 4593
rect 1101 4587 1136 4588
rect 112 4548 146 4576
rect 338 4550 375 4579
rect 339 4548 375 4550
rect 551 4548 588 4579
rect 112 4547 284 4548
rect 112 4515 298 4547
rect 339 4526 588 4548
rect 759 4547 796 4579
rect 1072 4575 1136 4587
rect 1176 4549 1203 4727
rect 2331 4699 2384 4806
rect 3731 4705 3758 4883
rect 3798 4845 3862 4857
rect 4138 4853 4175 4885
rect 4346 4884 4595 4906
rect 4346 4853 4383 4884
rect 4559 4882 4595 4884
rect 4559 4853 4596 4882
rect 3798 4844 3833 4845
rect 3775 4839 3833 4844
rect 3775 4819 3778 4839
rect 3798 4825 3833 4839
rect 3853 4825 3862 4845
rect 3798 4817 3862 4825
rect 3824 4816 3862 4817
rect 3825 4815 3862 4816
rect 3928 4849 3964 4850
rect 4036 4849 4072 4850
rect 3928 4844 4072 4849
rect 3928 4841 3990 4844
rect 3928 4821 3936 4841
rect 3956 4824 3990 4841
rect 4013 4841 4072 4844
rect 4013 4824 4044 4841
rect 3956 4821 4044 4824
rect 4064 4821 4072 4841
rect 3928 4815 4072 4821
rect 4138 4845 4176 4853
rect 4244 4849 4280 4850
rect 4138 4825 4147 4845
rect 4167 4825 4176 4845
rect 4138 4816 4176 4825
rect 4195 4842 4280 4849
rect 4195 4822 4202 4842
rect 4223 4841 4280 4842
rect 4223 4822 4252 4841
rect 4195 4821 4252 4822
rect 4272 4821 4280 4841
rect 4138 4815 4175 4816
rect 4195 4815 4280 4821
rect 4346 4845 4384 4853
rect 4457 4849 4493 4850
rect 4346 4825 4355 4845
rect 4375 4825 4384 4845
rect 4346 4816 4384 4825
rect 4408 4841 4493 4849
rect 4408 4821 4465 4841
rect 4485 4821 4493 4841
rect 4346 4815 4383 4816
rect 4408 4815 4493 4821
rect 4559 4845 4597 4853
rect 4559 4825 4568 4845
rect 4588 4825 4597 4845
rect 4559 4816 4597 4825
rect 4559 4815 4596 4816
rect 3982 4794 4018 4815
rect 4408 4794 4439 4815
rect 3815 4790 3915 4794
rect 3815 4786 3877 4790
rect 3815 4760 3822 4786
rect 3848 4764 3877 4786
rect 3903 4764 3915 4790
rect 3848 4760 3915 4764
rect 3815 4757 3915 4760
rect 3983 4757 4018 4794
rect 4080 4791 4439 4794
rect 4080 4786 4302 4791
rect 4080 4762 4093 4786
rect 4117 4767 4302 4786
rect 4326 4767 4439 4791
rect 4117 4762 4439 4767
rect 4080 4758 4439 4762
rect 4506 4786 4655 4794
rect 4506 4766 4517 4786
rect 4537 4766 4655 4786
rect 4506 4759 4655 4766
rect 4506 4758 4547 4759
rect 3830 4705 3867 4706
rect 3926 4705 3963 4706
rect 3982 4705 4018 4757
rect 4037 4705 4074 4706
rect 2331 4681 2379 4699
rect 2331 4641 2339 4681
rect 2366 4641 2379 4681
rect 3730 4696 3868 4705
rect 3730 4676 3839 4696
rect 3859 4676 3868 4696
rect 3730 4669 3868 4676
rect 3926 4696 4074 4705
rect 3926 4676 3935 4696
rect 3955 4676 4045 4696
rect 4065 4676 4074 4696
rect 3730 4667 3826 4669
rect 3926 4666 4074 4676
rect 4133 4696 4170 4706
rect 4245 4705 4282 4706
rect 4226 4703 4282 4705
rect 4133 4676 4141 4696
rect 4161 4676 4170 4696
rect 3982 4665 4018 4666
rect 1359 4623 1469 4637
rect 2331 4627 2379 4641
rect 3464 4632 3575 4647
rect 3464 4630 3506 4632
rect 1359 4620 1402 4623
rect 1359 4615 1363 4620
rect 1035 4547 1203 4549
rect 759 4541 1203 4547
rect 112 4483 146 4515
rect 108 4474 146 4483
rect 108 4456 118 4474
rect 136 4456 146 4474
rect 108 4450 146 4456
rect 264 4452 298 4515
rect 420 4520 531 4526
rect 420 4512 461 4520
rect 420 4492 428 4512
rect 447 4492 461 4512
rect 420 4490 461 4492
rect 489 4512 531 4520
rect 489 4492 505 4512
rect 524 4492 531 4512
rect 489 4490 531 4492
rect 420 4475 531 4490
rect 758 4521 1203 4541
rect 758 4452 796 4521
rect 1035 4520 1203 4521
rect 1281 4593 1363 4615
rect 1392 4593 1402 4620
rect 1430 4596 1437 4623
rect 1466 4615 1469 4623
rect 1466 4596 1531 4615
rect 1430 4593 1531 4596
rect 1281 4591 1531 4593
rect 1281 4512 1318 4591
rect 1359 4578 1469 4591
rect 1433 4522 1464 4523
rect 1281 4492 1290 4512
rect 1310 4492 1318 4512
rect 1281 4482 1318 4492
rect 1377 4512 1464 4522
rect 1377 4492 1386 4512
rect 1406 4492 1464 4512
rect 1377 4483 1464 4492
rect 1377 4482 1414 4483
rect 108 4446 145 4450
rect 264 4441 796 4452
rect 263 4425 796 4441
rect 1433 4430 1464 4483
rect 1494 4512 1531 4591
rect 1702 4588 2095 4608
rect 2115 4588 2118 4608
rect 3197 4603 3238 4612
rect 1702 4583 2118 4588
rect 2792 4601 2960 4602
rect 3197 4601 3206 4603
rect 1702 4582 2043 4583
rect 1646 4522 1677 4523
rect 1494 4492 1503 4512
rect 1523 4492 1531 4512
rect 1494 4482 1531 4492
rect 1590 4515 1677 4522
rect 1590 4512 1651 4515
rect 1590 4492 1599 4512
rect 1619 4495 1651 4512
rect 1672 4495 1677 4515
rect 1619 4492 1677 4495
rect 1590 4485 1677 4492
rect 1702 4512 1739 4582
rect 2005 4581 2042 4582
rect 2792 4581 3206 4601
rect 3232 4581 3238 4603
rect 3464 4610 3471 4630
rect 3490 4610 3506 4630
rect 3464 4602 3506 4610
rect 3534 4630 3575 4632
rect 3534 4610 3548 4630
rect 3567 4610 3575 4630
rect 3534 4602 3575 4610
rect 3830 4606 3867 4607
rect 4133 4606 4170 4676
rect 4195 4696 4282 4703
rect 4195 4693 4253 4696
rect 4195 4673 4200 4693
rect 4221 4676 4253 4693
rect 4273 4676 4282 4696
rect 4221 4673 4282 4676
rect 4195 4666 4282 4673
rect 4341 4696 4378 4706
rect 4341 4676 4349 4696
rect 4369 4676 4378 4696
rect 4195 4665 4226 4666
rect 3829 4605 4170 4606
rect 3464 4596 3575 4602
rect 3754 4600 4170 4605
rect 2792 4575 3238 4581
rect 2792 4573 2960 4575
rect 1854 4522 1890 4523
rect 1702 4492 1711 4512
rect 1731 4492 1739 4512
rect 1590 4483 1646 4485
rect 1590 4482 1627 4483
rect 1702 4482 1739 4492
rect 1798 4512 1946 4522
rect 2046 4519 2142 4521
rect 1798 4492 1807 4512
rect 1827 4492 1917 4512
rect 1937 4492 1946 4512
rect 1798 4483 1946 4492
rect 2004 4512 2142 4519
rect 2004 4492 2013 4512
rect 2033 4492 2142 4512
rect 2004 4483 2142 4492
rect 1798 4482 1835 4483
rect 1854 4431 1890 4483
rect 1909 4482 1946 4483
rect 2005 4482 2042 4483
rect 1325 4429 1366 4430
rect 263 4424 777 4425
rect 1217 4422 1366 4429
rect 1217 4402 1335 4422
rect 1355 4402 1366 4422
rect 1217 4394 1366 4402
rect 1433 4426 1792 4430
rect 1433 4421 1755 4426
rect 1433 4397 1546 4421
rect 1570 4402 1755 4421
rect 1779 4402 1792 4426
rect 1570 4397 1792 4402
rect 1433 4394 1792 4397
rect 1854 4394 1889 4431
rect 1957 4428 2057 4431
rect 1957 4424 2024 4428
rect 1957 4398 1969 4424
rect 1995 4402 2024 4424
rect 2050 4402 2057 4428
rect 1995 4398 2057 4402
rect 1957 4394 2057 4398
rect 111 4383 148 4384
rect 109 4375 149 4383
rect 109 4357 120 4375
rect 138 4357 149 4375
rect 1433 4373 1464 4394
rect 1854 4373 1890 4394
rect 1276 4372 1313 4373
rect 109 4309 149 4357
rect 1275 4363 1313 4372
rect 1275 4343 1284 4363
rect 1304 4343 1313 4363
rect 1275 4335 1313 4343
rect 1379 4367 1464 4373
rect 1489 4372 1526 4373
rect 1379 4347 1387 4367
rect 1407 4347 1464 4367
rect 1379 4339 1464 4347
rect 1488 4363 1526 4372
rect 1488 4343 1497 4363
rect 1517 4343 1526 4363
rect 1379 4338 1415 4339
rect 1488 4335 1526 4343
rect 1592 4367 1677 4373
rect 1697 4372 1734 4373
rect 1592 4347 1600 4367
rect 1620 4366 1677 4367
rect 1620 4347 1649 4366
rect 1592 4346 1649 4347
rect 1670 4346 1677 4366
rect 1592 4339 1677 4346
rect 1696 4363 1734 4372
rect 1696 4343 1705 4363
rect 1725 4343 1734 4363
rect 1592 4338 1628 4339
rect 1696 4335 1734 4343
rect 1800 4367 1944 4373
rect 1800 4347 1808 4367
rect 1828 4350 1864 4367
rect 1884 4350 1916 4367
rect 1828 4347 1916 4350
rect 1936 4347 1944 4367
rect 1800 4339 1944 4347
rect 1800 4338 1836 4339
rect 1908 4338 1944 4339
rect 2010 4372 2047 4373
rect 2010 4371 2048 4372
rect 2010 4363 2074 4371
rect 2010 4343 2019 4363
rect 2039 4349 2074 4363
rect 2094 4349 2097 4369
rect 2039 4344 2097 4349
rect 2039 4343 2074 4344
rect 420 4313 530 4327
rect 420 4310 463 4313
rect 109 4302 234 4309
rect 420 4305 424 4310
rect 109 4283 201 4302
rect 226 4283 234 4302
rect 109 4273 234 4283
rect 342 4283 424 4305
rect 453 4283 463 4310
rect 491 4286 498 4313
rect 527 4305 530 4313
rect 1276 4306 1313 4335
rect 527 4286 592 4305
rect 1277 4304 1313 4306
rect 1489 4304 1526 4335
rect 1697 4308 1734 4335
rect 2010 4331 2074 4343
rect 491 4283 592 4286
rect 342 4281 592 4283
rect 109 4253 149 4273
rect 108 4244 149 4253
rect 108 4226 118 4244
rect 136 4226 149 4244
rect 108 4217 149 4226
rect 108 4216 145 4217
rect 342 4202 379 4281
rect 420 4268 530 4281
rect 494 4212 525 4213
rect 342 4182 351 4202
rect 371 4182 379 4202
rect 342 4172 379 4182
rect 438 4202 525 4212
rect 438 4182 447 4202
rect 467 4182 525 4202
rect 438 4173 525 4182
rect 438 4172 475 4173
rect 111 4150 148 4154
rect 108 4145 148 4150
rect 108 4127 120 4145
rect 138 4127 148 4145
rect 108 3947 148 4127
rect 494 4120 525 4173
rect 555 4202 592 4281
rect 763 4278 1156 4298
rect 1176 4278 1179 4298
rect 1277 4282 1526 4304
rect 1695 4303 1736 4308
rect 2114 4305 2141 4483
rect 2792 4395 2819 4573
rect 3197 4570 3238 4575
rect 3407 4574 3656 4596
rect 3754 4580 3757 4600
rect 3777 4580 4170 4600
rect 4341 4597 4378 4676
rect 4408 4705 4439 4758
rect 4785 4751 4825 4931
rect 5163 4933 5202 4971
rect 6382 4973 6500 4993
rect 6520 4973 6531 4993
rect 6382 4965 6531 4973
rect 6598 4997 6957 5001
rect 6598 4992 6920 4997
rect 6598 4968 6711 4992
rect 6735 4973 6920 4992
rect 6944 4973 6957 4997
rect 6735 4968 6957 4973
rect 6598 4965 6957 4968
rect 7019 4965 7054 5002
rect 7122 4999 7222 5002
rect 7122 4995 7189 4999
rect 7122 4969 7134 4995
rect 7160 4973 7189 4995
rect 7215 4973 7222 4999
rect 7160 4969 7222 4973
rect 7122 4965 7222 4969
rect 6598 4944 6629 4965
rect 7019 4944 7055 4965
rect 6441 4943 6478 4944
rect 6440 4934 6478 4943
rect 5163 4931 5211 4933
rect 5163 4913 5174 4931
rect 5192 4913 5211 4931
rect 5163 4904 5211 4913
rect 5164 4903 5211 4904
rect 5477 4908 5587 4922
rect 5477 4905 5520 4908
rect 5477 4900 5481 4905
rect 5399 4878 5481 4900
rect 5510 4878 5520 4905
rect 5548 4881 5555 4908
rect 5584 4900 5587 4908
rect 6440 4914 6449 4934
rect 6469 4914 6478 4934
rect 6440 4906 6478 4914
rect 6544 4938 6629 4944
rect 6654 4943 6691 4944
rect 6544 4918 6552 4938
rect 6572 4918 6629 4938
rect 6544 4910 6629 4918
rect 6653 4934 6691 4943
rect 6653 4914 6662 4934
rect 6682 4914 6691 4934
rect 6544 4909 6580 4910
rect 6653 4906 6691 4914
rect 6757 4938 6842 4944
rect 6862 4943 6899 4944
rect 6757 4918 6765 4938
rect 6785 4937 6842 4938
rect 6785 4918 6814 4937
rect 6757 4917 6814 4918
rect 6835 4917 6842 4937
rect 6757 4910 6842 4917
rect 6861 4934 6899 4943
rect 6861 4914 6870 4934
rect 6890 4914 6899 4934
rect 6757 4909 6793 4910
rect 6861 4906 6899 4914
rect 6965 4940 7109 4944
rect 6965 4938 7022 4940
rect 6965 4918 6973 4938
rect 6993 4918 7022 4938
rect 6965 4916 7022 4918
rect 7048 4938 7109 4940
rect 7048 4918 7081 4938
rect 7101 4918 7109 4938
rect 7048 4916 7109 4918
rect 6965 4910 7109 4916
rect 6965 4909 7001 4910
rect 7073 4909 7109 4910
rect 7175 4943 7212 4944
rect 7175 4942 7213 4943
rect 7175 4934 7239 4942
rect 7175 4914 7184 4934
rect 7204 4920 7239 4934
rect 7259 4920 7262 4940
rect 7204 4915 7262 4920
rect 7204 4914 7239 4915
rect 5584 4881 5649 4900
rect 5548 4878 5649 4881
rect 5399 4876 5649 4878
rect 5167 4840 5204 4841
rect 4785 4733 4795 4751
rect 4813 4733 4825 4751
rect 4785 4728 4825 4733
rect 5163 4837 5204 4840
rect 5163 4832 5205 4837
rect 5163 4814 5176 4832
rect 5194 4814 5205 4832
rect 5163 4800 5205 4814
rect 5243 4800 5290 4804
rect 5163 4794 5290 4800
rect 5163 4765 5251 4794
rect 5280 4765 5290 4794
rect 5399 4797 5436 4876
rect 5477 4863 5587 4876
rect 5551 4807 5582 4808
rect 5399 4777 5408 4797
rect 5428 4777 5436 4797
rect 5399 4767 5436 4777
rect 5495 4797 5582 4807
rect 5495 4777 5504 4797
rect 5524 4777 5582 4797
rect 5495 4768 5582 4777
rect 5495 4767 5532 4768
rect 5163 4761 5290 4765
rect 5163 4744 5202 4761
rect 5243 4760 5290 4761
rect 4785 4724 4822 4728
rect 5163 4726 5174 4744
rect 5192 4726 5202 4744
rect 5163 4717 5202 4726
rect 5164 4716 5201 4717
rect 5551 4715 5582 4768
rect 5612 4797 5649 4876
rect 5820 4873 6213 4893
rect 6233 4873 6236 4893
rect 6441 4877 6478 4906
rect 5820 4868 6236 4873
rect 6442 4875 6478 4877
rect 6654 4875 6691 4906
rect 5820 4867 6161 4868
rect 5764 4807 5795 4808
rect 5612 4777 5621 4797
rect 5641 4777 5649 4797
rect 5612 4767 5649 4777
rect 5708 4800 5795 4807
rect 5708 4797 5769 4800
rect 5708 4777 5717 4797
rect 5737 4780 5769 4797
rect 5790 4780 5795 4800
rect 5737 4777 5795 4780
rect 5708 4770 5795 4777
rect 5820 4797 5857 4867
rect 6123 4866 6160 4867
rect 6442 4853 6691 4875
rect 6862 4874 6899 4906
rect 7175 4902 7239 4914
rect 7279 4877 7306 5054
rect 7739 5009 7766 5186
rect 7806 5149 7870 5161
rect 8146 5157 8183 5189
rect 8354 5188 8603 5210
rect 8885 5196 8922 5197
rect 9188 5196 9225 5266
rect 9250 5286 9337 5293
rect 9250 5283 9308 5286
rect 9250 5263 9255 5283
rect 9276 5266 9308 5283
rect 9328 5266 9337 5286
rect 9276 5263 9337 5266
rect 9250 5256 9337 5263
rect 9396 5286 9433 5296
rect 9396 5266 9404 5286
rect 9424 5266 9433 5286
rect 9250 5255 9281 5256
rect 8884 5195 9225 5196
rect 8354 5157 8391 5188
rect 8567 5186 8603 5188
rect 8809 5190 9225 5195
rect 8567 5157 8604 5186
rect 8809 5170 8812 5190
rect 8832 5170 9225 5190
rect 9396 5187 9433 5266
rect 9463 5295 9494 5348
rect 9844 5346 9881 5347
rect 9843 5337 9882 5346
rect 9843 5319 9853 5337
rect 9871 5319 9882 5337
rect 10139 5334 10149 5352
rect 10167 5334 10180 5352
rect 10139 5325 10180 5334
rect 10139 5324 10176 5325
rect 9755 5302 9802 5303
rect 9843 5302 9882 5319
rect 9755 5298 9882 5302
rect 9513 5295 9550 5296
rect 9463 5286 9550 5295
rect 9463 5266 9521 5286
rect 9541 5266 9550 5286
rect 9463 5256 9550 5266
rect 9609 5286 9646 5296
rect 9609 5266 9617 5286
rect 9637 5266 9646 5286
rect 9463 5255 9494 5256
rect 9458 5187 9568 5200
rect 9609 5187 9646 5266
rect 9755 5269 9765 5298
rect 9794 5269 9882 5298
rect 10373 5310 10410 5389
rect 10451 5376 10561 5389
rect 10525 5320 10556 5321
rect 10373 5290 10382 5310
rect 10402 5290 10410 5310
rect 10373 5280 10410 5290
rect 10469 5310 10556 5320
rect 10469 5290 10478 5310
rect 10498 5290 10556 5310
rect 10469 5281 10556 5290
rect 10469 5280 10506 5281
rect 9755 5263 9882 5269
rect 9755 5259 9802 5263
rect 9840 5249 9882 5263
rect 10142 5258 10179 5262
rect 9840 5231 9851 5249
rect 9869 5231 9882 5249
rect 9840 5226 9882 5231
rect 9841 5223 9882 5226
rect 10139 5253 10179 5258
rect 10139 5235 10151 5253
rect 10169 5235 10179 5253
rect 9841 5222 9878 5223
rect 9396 5185 9646 5187
rect 9396 5182 9497 5185
rect 9396 5163 9461 5182
rect 7806 5148 7841 5149
rect 7783 5143 7841 5148
rect 7783 5123 7786 5143
rect 7806 5129 7841 5143
rect 7861 5129 7870 5149
rect 7806 5121 7870 5129
rect 7832 5120 7870 5121
rect 7833 5119 7870 5120
rect 7936 5153 7972 5154
rect 8044 5153 8080 5154
rect 7936 5146 8080 5153
rect 7936 5145 7993 5146
rect 7936 5125 7944 5145
rect 7964 5126 7993 5145
rect 8018 5145 8080 5146
rect 8018 5126 8052 5145
rect 7964 5125 8052 5126
rect 8072 5125 8080 5145
rect 7936 5119 8080 5125
rect 8146 5149 8184 5157
rect 8252 5153 8288 5154
rect 8146 5129 8155 5149
rect 8175 5129 8184 5149
rect 8146 5120 8184 5129
rect 8203 5146 8288 5153
rect 8203 5126 8210 5146
rect 8231 5145 8288 5146
rect 8231 5126 8260 5145
rect 8203 5125 8260 5126
rect 8280 5125 8288 5145
rect 8146 5119 8183 5120
rect 8203 5119 8288 5125
rect 8354 5149 8392 5157
rect 8465 5153 8501 5154
rect 8354 5129 8363 5149
rect 8383 5129 8392 5149
rect 8354 5120 8392 5129
rect 8416 5145 8501 5153
rect 8416 5125 8473 5145
rect 8493 5125 8501 5145
rect 8354 5119 8391 5120
rect 8416 5119 8501 5125
rect 8567 5149 8605 5157
rect 8567 5129 8576 5149
rect 8596 5129 8605 5149
rect 9458 5155 9461 5163
rect 9490 5155 9497 5182
rect 9525 5158 9535 5185
rect 9564 5163 9646 5185
rect 9564 5158 9568 5163
rect 9525 5155 9568 5158
rect 9458 5141 9568 5155
rect 9834 5159 9881 5160
rect 9834 5150 9882 5159
rect 9834 5132 9853 5150
rect 9871 5132 9882 5150
rect 9834 5130 9882 5132
rect 8567 5120 8605 5129
rect 8567 5119 8604 5120
rect 7990 5098 8026 5119
rect 8416 5098 8447 5119
rect 7823 5094 7923 5098
rect 7823 5090 7885 5094
rect 7823 5064 7830 5090
rect 7856 5068 7885 5090
rect 7911 5068 7923 5094
rect 7856 5064 7923 5068
rect 7823 5061 7923 5064
rect 7991 5061 8026 5098
rect 8088 5095 8447 5098
rect 8088 5090 8310 5095
rect 8088 5066 8101 5090
rect 8125 5071 8310 5090
rect 8334 5071 8447 5095
rect 8125 5066 8447 5071
rect 8088 5062 8447 5066
rect 8514 5090 8663 5098
rect 8514 5070 8525 5090
rect 8545 5070 8663 5090
rect 9843 5092 9882 5130
rect 8514 5063 8663 5070
rect 9195 5073 9233 5075
rect 9843 5073 9885 5092
rect 8514 5062 8555 5063
rect 7990 5057 8026 5061
rect 7990 5028 8027 5057
rect 7838 5009 7875 5010
rect 7934 5009 7971 5010
rect 7990 5009 8026 5028
rect 8045 5009 8082 5010
rect 7738 5000 7876 5009
rect 7738 4980 7847 5000
rect 7867 4980 7876 5000
rect 7738 4973 7876 4980
rect 7934 5000 8082 5009
rect 7934 4980 7943 5000
rect 7963 4980 8053 5000
rect 8073 4980 8082 5000
rect 7738 4971 7834 4973
rect 7934 4970 8082 4980
rect 8141 5000 8178 5010
rect 8253 5009 8290 5010
rect 8234 5007 8290 5009
rect 8141 4980 8149 5000
rect 8169 4980 8178 5000
rect 7990 4969 8026 4970
rect 7838 4910 7875 4911
rect 8141 4910 8178 4980
rect 8203 5000 8290 5007
rect 8203 4997 8261 5000
rect 8203 4977 8208 4997
rect 8229 4980 8261 4997
rect 8281 4980 8290 5000
rect 8229 4977 8290 4980
rect 8203 4970 8290 4977
rect 8349 5000 8386 5010
rect 8349 4980 8357 5000
rect 8377 4980 8386 5000
rect 8203 4969 8234 4970
rect 7837 4909 8178 4910
rect 7762 4904 8178 4909
rect 7387 4877 7440 4885
rect 7762 4884 7765 4904
rect 7785 4884 8178 4904
rect 8349 4901 8386 4980
rect 8416 5009 8447 5062
rect 9195 5050 9885 5073
rect 10139 5055 10179 5235
rect 10525 5228 10556 5281
rect 10586 5310 10623 5389
rect 10794 5386 11187 5406
rect 11207 5386 11210 5406
rect 11308 5390 11557 5412
rect 11726 5411 11767 5416
rect 12145 5413 12172 5591
rect 12823 5503 12850 5681
rect 13228 5678 13269 5683
rect 13438 5682 13687 5704
rect 13785 5688 13788 5708
rect 13808 5688 14201 5708
rect 14372 5705 14409 5784
rect 14439 5813 14470 5866
rect 14816 5859 14856 6039
rect 15194 6199 15234 6379
rect 15580 6372 15611 6425
rect 15641 6454 15678 6533
rect 15849 6530 16242 6550
rect 16262 6530 16265 6550
rect 16363 6534 16612 6556
rect 16781 6555 16822 6560
rect 17200 6557 17227 6735
rect 17878 6647 17905 6825
rect 18283 6822 18324 6827
rect 18493 6826 18742 6848
rect 18840 6832 18843 6852
rect 18863 6832 19256 6852
rect 19427 6849 19464 6928
rect 19494 6957 19525 7010
rect 19871 7003 19911 7183
rect 19871 6985 19881 7003
rect 19899 6985 19911 7003
rect 19871 6980 19911 6985
rect 19871 6976 19908 6980
rect 19544 6957 19581 6958
rect 19494 6948 19581 6957
rect 19494 6928 19552 6948
rect 19572 6928 19581 6948
rect 19494 6918 19581 6928
rect 19640 6948 19677 6958
rect 19640 6928 19648 6948
rect 19668 6928 19677 6948
rect 19494 6917 19525 6918
rect 19489 6849 19599 6862
rect 19640 6849 19677 6928
rect 19874 6913 19911 6914
rect 19870 6904 19911 6913
rect 19870 6886 19883 6904
rect 19901 6886 19911 6904
rect 19870 6877 19911 6886
rect 19870 6857 19910 6877
rect 19427 6847 19677 6849
rect 19427 6844 19528 6847
rect 17945 6787 18009 6799
rect 18285 6795 18322 6822
rect 18493 6795 18530 6826
rect 18706 6824 18742 6826
rect 19427 6825 19492 6844
rect 18706 6795 18743 6824
rect 19489 6817 19492 6825
rect 19521 6817 19528 6844
rect 19556 6820 19566 6847
rect 19595 6825 19677 6847
rect 19785 6847 19910 6857
rect 19785 6828 19793 6847
rect 19818 6828 19910 6847
rect 19595 6820 19599 6825
rect 19785 6821 19910 6828
rect 19556 6817 19599 6820
rect 19489 6803 19599 6817
rect 17945 6786 17980 6787
rect 17922 6781 17980 6786
rect 17922 6761 17925 6781
rect 17945 6767 17980 6781
rect 18000 6767 18009 6787
rect 17945 6759 18009 6767
rect 17971 6758 18009 6759
rect 17972 6757 18009 6758
rect 18075 6791 18111 6792
rect 18183 6791 18219 6792
rect 18075 6783 18219 6791
rect 18075 6763 18083 6783
rect 18103 6763 18191 6783
rect 18211 6763 18219 6783
rect 18075 6757 18219 6763
rect 18285 6787 18323 6795
rect 18391 6791 18427 6792
rect 18285 6767 18294 6787
rect 18314 6767 18323 6787
rect 18285 6758 18323 6767
rect 18342 6784 18427 6791
rect 18342 6764 18349 6784
rect 18370 6783 18427 6784
rect 18370 6764 18399 6783
rect 18342 6763 18399 6764
rect 18419 6763 18427 6783
rect 18285 6757 18322 6758
rect 18342 6757 18427 6763
rect 18493 6787 18531 6795
rect 18604 6791 18640 6792
rect 18493 6767 18502 6787
rect 18522 6767 18531 6787
rect 18493 6758 18531 6767
rect 18555 6783 18640 6791
rect 18555 6763 18612 6783
rect 18632 6763 18640 6783
rect 18493 6757 18530 6758
rect 18555 6757 18640 6763
rect 18706 6787 18744 6795
rect 18706 6767 18715 6787
rect 18735 6767 18744 6787
rect 18706 6758 18744 6767
rect 19870 6773 19910 6821
rect 18706 6757 18743 6758
rect 18129 6736 18165 6757
rect 18555 6736 18586 6757
rect 19870 6755 19881 6773
rect 19899 6755 19910 6773
rect 19870 6747 19910 6755
rect 19871 6746 19908 6747
rect 17962 6732 18062 6736
rect 17962 6728 18024 6732
rect 17962 6702 17969 6728
rect 17995 6706 18024 6728
rect 18050 6706 18062 6732
rect 17995 6702 18062 6706
rect 17962 6699 18062 6702
rect 18130 6699 18165 6736
rect 18227 6733 18586 6736
rect 18227 6728 18449 6733
rect 18227 6704 18240 6728
rect 18264 6709 18449 6728
rect 18473 6709 18586 6733
rect 18264 6704 18586 6709
rect 18227 6700 18586 6704
rect 18653 6728 18802 6736
rect 18653 6708 18664 6728
rect 18684 6708 18802 6728
rect 18653 6701 18802 6708
rect 19242 6705 19756 6706
rect 18653 6700 18694 6701
rect 18129 6664 18165 6699
rect 17977 6647 18014 6648
rect 18073 6647 18110 6648
rect 18129 6647 18136 6664
rect 17877 6638 18015 6647
rect 17877 6618 17986 6638
rect 18006 6618 18015 6638
rect 17877 6611 18015 6618
rect 18073 6638 18136 6647
rect 18073 6618 18082 6638
rect 18102 6623 18136 6638
rect 18157 6647 18165 6664
rect 18184 6647 18221 6648
rect 18157 6638 18221 6647
rect 18157 6623 18192 6638
rect 18102 6618 18192 6623
rect 18212 6618 18221 6638
rect 17877 6609 17973 6611
rect 18073 6608 18221 6618
rect 18280 6638 18317 6648
rect 18392 6647 18429 6648
rect 18373 6645 18429 6647
rect 18280 6618 18288 6638
rect 18308 6618 18317 6638
rect 18129 6607 18165 6608
rect 17059 6555 17227 6557
rect 16781 6549 17227 6555
rect 15849 6525 16265 6530
rect 16444 6528 16555 6534
rect 15849 6524 16190 6525
rect 15793 6464 15824 6465
rect 15641 6434 15650 6454
rect 15670 6434 15678 6454
rect 15641 6424 15678 6434
rect 15737 6457 15824 6464
rect 15737 6454 15798 6457
rect 15737 6434 15746 6454
rect 15766 6437 15798 6454
rect 15819 6437 15824 6457
rect 15766 6434 15824 6437
rect 15737 6427 15824 6434
rect 15849 6454 15886 6524
rect 16152 6523 16189 6524
rect 16444 6520 16485 6528
rect 16444 6500 16452 6520
rect 16471 6500 16485 6520
rect 16444 6498 16485 6500
rect 16513 6520 16555 6528
rect 16513 6500 16529 6520
rect 16548 6500 16555 6520
rect 16781 6527 16787 6549
rect 16813 6529 17227 6549
rect 17977 6548 18014 6549
rect 18280 6548 18317 6618
rect 18342 6638 18429 6645
rect 18342 6635 18400 6638
rect 18342 6615 18347 6635
rect 18368 6618 18400 6635
rect 18420 6618 18429 6638
rect 18368 6615 18429 6618
rect 18342 6608 18429 6615
rect 18488 6638 18525 6648
rect 18488 6618 18496 6638
rect 18516 6618 18525 6638
rect 18342 6607 18373 6608
rect 17976 6547 18317 6548
rect 16813 6527 16822 6529
rect 17059 6528 17227 6529
rect 17901 6546 18317 6547
rect 17901 6542 18277 6546
rect 16781 6518 16822 6527
rect 17901 6522 17904 6542
rect 17924 6529 18277 6542
rect 18309 6529 18317 6546
rect 17924 6522 18317 6529
rect 18488 6539 18525 6618
rect 18555 6647 18586 6700
rect 19223 6689 19756 6705
rect 19223 6678 19755 6689
rect 19874 6680 19911 6684
rect 18605 6647 18642 6648
rect 18555 6638 18642 6647
rect 18555 6618 18613 6638
rect 18633 6618 18642 6638
rect 18555 6608 18642 6618
rect 18701 6638 18738 6648
rect 18701 6618 18709 6638
rect 18729 6618 18738 6638
rect 18555 6607 18586 6608
rect 18550 6539 18660 6552
rect 18701 6539 18738 6618
rect 18488 6537 18738 6539
rect 18488 6534 18589 6537
rect 18488 6515 18553 6534
rect 16513 6498 16555 6500
rect 16444 6483 16555 6498
rect 18550 6507 18553 6515
rect 18582 6507 18589 6534
rect 18617 6510 18627 6537
rect 18656 6515 18738 6537
rect 18816 6609 18984 6610
rect 19223 6609 19261 6678
rect 18816 6589 19261 6609
rect 19488 6640 19599 6655
rect 19488 6638 19530 6640
rect 19488 6618 19495 6638
rect 19514 6618 19530 6638
rect 19488 6610 19530 6618
rect 19558 6638 19599 6640
rect 19558 6618 19572 6638
rect 19591 6618 19599 6638
rect 19558 6610 19599 6618
rect 19488 6604 19599 6610
rect 19721 6615 19755 6678
rect 19873 6674 19911 6680
rect 19873 6656 19883 6674
rect 19901 6656 19911 6674
rect 19873 6647 19911 6656
rect 19873 6615 19907 6647
rect 18816 6583 19260 6589
rect 18816 6581 18984 6583
rect 18656 6510 18660 6515
rect 18617 6507 18660 6510
rect 18550 6493 18660 6507
rect 16001 6464 16037 6465
rect 15849 6434 15858 6454
rect 15878 6434 15886 6454
rect 15737 6425 15793 6427
rect 15737 6424 15774 6425
rect 15849 6424 15886 6434
rect 15945 6454 16093 6464
rect 16193 6461 16289 6463
rect 15945 6434 15954 6454
rect 15974 6434 16064 6454
rect 16084 6434 16093 6454
rect 15945 6425 16093 6434
rect 16151 6454 16289 6461
rect 16151 6434 16160 6454
rect 16180 6434 16289 6454
rect 16151 6425 16289 6434
rect 15945 6424 15982 6425
rect 16001 6373 16037 6425
rect 16056 6424 16093 6425
rect 16152 6424 16189 6425
rect 15472 6371 15513 6372
rect 15364 6364 15513 6371
rect 15364 6344 15482 6364
rect 15502 6344 15513 6364
rect 15364 6336 15513 6344
rect 15580 6368 15939 6372
rect 15580 6363 15902 6368
rect 15580 6339 15693 6363
rect 15717 6344 15902 6363
rect 15926 6344 15939 6368
rect 15717 6339 15939 6344
rect 15580 6336 15939 6339
rect 16001 6336 16036 6373
rect 16104 6370 16204 6373
rect 16104 6366 16171 6370
rect 16104 6340 16116 6366
rect 16142 6344 16171 6366
rect 16197 6344 16204 6370
rect 16142 6340 16204 6344
rect 16104 6336 16204 6340
rect 15580 6315 15611 6336
rect 16001 6315 16037 6336
rect 15423 6314 15460 6315
rect 15422 6305 15460 6314
rect 15422 6285 15431 6305
rect 15451 6285 15460 6305
rect 15422 6277 15460 6285
rect 15526 6309 15611 6315
rect 15636 6314 15673 6315
rect 15526 6289 15534 6309
rect 15554 6289 15611 6309
rect 15526 6281 15611 6289
rect 15635 6305 15673 6314
rect 15635 6285 15644 6305
rect 15664 6285 15673 6305
rect 15526 6280 15562 6281
rect 15635 6277 15673 6285
rect 15739 6309 15824 6315
rect 15844 6314 15881 6315
rect 15739 6289 15747 6309
rect 15767 6308 15824 6309
rect 15767 6289 15796 6308
rect 15739 6288 15796 6289
rect 15817 6288 15824 6308
rect 15739 6281 15824 6288
rect 15843 6305 15881 6314
rect 15843 6285 15852 6305
rect 15872 6285 15881 6305
rect 15739 6280 15775 6281
rect 15843 6277 15881 6285
rect 15947 6309 16091 6315
rect 15947 6289 15955 6309
rect 15975 6306 16063 6309
rect 15975 6289 16006 6306
rect 15947 6286 16006 6289
rect 16029 6289 16063 6306
rect 16083 6289 16091 6309
rect 16029 6286 16091 6289
rect 15947 6281 16091 6286
rect 15947 6280 15983 6281
rect 16055 6280 16091 6281
rect 16157 6314 16194 6315
rect 16157 6313 16195 6314
rect 16157 6305 16221 6313
rect 16157 6285 16166 6305
rect 16186 6291 16221 6305
rect 16241 6291 16244 6311
rect 16186 6286 16244 6291
rect 16186 6285 16221 6286
rect 15423 6248 15460 6277
rect 15424 6246 15460 6248
rect 15636 6246 15673 6277
rect 15424 6224 15673 6246
rect 15844 6245 15881 6277
rect 16157 6273 16221 6285
rect 16261 6247 16288 6425
rect 18816 6403 18843 6581
rect 18883 6543 18947 6555
rect 19223 6551 19260 6583
rect 19431 6582 19680 6604
rect 19721 6583 19907 6615
rect 19735 6582 19907 6583
rect 19431 6551 19468 6582
rect 19644 6580 19680 6582
rect 19644 6551 19681 6580
rect 19873 6554 19907 6582
rect 18883 6542 18918 6543
rect 18860 6537 18918 6542
rect 18860 6517 18863 6537
rect 18883 6523 18918 6537
rect 18938 6523 18947 6543
rect 18883 6515 18947 6523
rect 18909 6514 18947 6515
rect 18910 6513 18947 6514
rect 19013 6547 19049 6548
rect 19121 6547 19157 6548
rect 19013 6540 19157 6547
rect 19013 6539 19073 6540
rect 19013 6519 19021 6539
rect 19041 6520 19073 6539
rect 19098 6539 19157 6540
rect 19098 6520 19129 6539
rect 19041 6519 19129 6520
rect 19149 6519 19157 6539
rect 19013 6513 19157 6519
rect 19223 6543 19261 6551
rect 19329 6547 19365 6548
rect 19223 6523 19232 6543
rect 19252 6523 19261 6543
rect 19223 6514 19261 6523
rect 19280 6540 19365 6547
rect 19280 6520 19287 6540
rect 19308 6539 19365 6540
rect 19308 6520 19337 6539
rect 19280 6519 19337 6520
rect 19357 6519 19365 6539
rect 19223 6513 19260 6514
rect 19280 6513 19365 6519
rect 19431 6543 19469 6551
rect 19542 6547 19578 6548
rect 19431 6523 19440 6543
rect 19460 6523 19469 6543
rect 19431 6514 19469 6523
rect 19493 6539 19578 6547
rect 19493 6519 19550 6539
rect 19570 6519 19578 6539
rect 19431 6513 19468 6514
rect 19493 6513 19578 6519
rect 19644 6543 19682 6551
rect 19644 6523 19653 6543
rect 19673 6523 19682 6543
rect 19644 6514 19682 6523
rect 19871 6544 19908 6554
rect 19871 6526 19881 6544
rect 19899 6526 19908 6544
rect 19871 6517 19908 6526
rect 19873 6516 19907 6517
rect 19644 6513 19681 6514
rect 19067 6492 19103 6513
rect 19493 6492 19524 6513
rect 18900 6488 19000 6492
rect 18900 6484 18962 6488
rect 18900 6458 18907 6484
rect 18933 6462 18962 6484
rect 18988 6462 19000 6488
rect 18933 6458 19000 6462
rect 18900 6455 19000 6458
rect 19068 6455 19103 6492
rect 19165 6489 19524 6492
rect 19165 6484 19387 6489
rect 19165 6460 19178 6484
rect 19202 6465 19387 6484
rect 19411 6465 19524 6489
rect 19202 6460 19524 6465
rect 19165 6456 19524 6460
rect 19591 6484 19740 6492
rect 19591 6464 19602 6484
rect 19622 6464 19740 6484
rect 19591 6457 19740 6464
rect 19591 6456 19632 6457
rect 18915 6403 18952 6404
rect 19011 6403 19048 6404
rect 19067 6403 19103 6455
rect 19122 6403 19159 6404
rect 18815 6394 18953 6403
rect 18410 6373 18521 6388
rect 18410 6371 18452 6373
rect 18080 6350 18185 6352
rect 17738 6342 17906 6343
rect 18080 6342 18129 6350
rect 17738 6323 18129 6342
rect 18160 6323 18185 6350
rect 18410 6351 18417 6371
rect 18436 6351 18452 6371
rect 18410 6343 18452 6351
rect 18480 6371 18521 6373
rect 18480 6351 18494 6371
rect 18513 6351 18521 6371
rect 18815 6374 18924 6394
rect 18944 6374 18953 6394
rect 18815 6367 18953 6374
rect 19011 6394 19159 6403
rect 19011 6374 19020 6394
rect 19040 6374 19130 6394
rect 19150 6374 19159 6394
rect 18815 6365 18911 6367
rect 19011 6364 19159 6374
rect 19218 6394 19255 6404
rect 19330 6403 19367 6404
rect 19311 6401 19367 6403
rect 19218 6374 19226 6394
rect 19246 6374 19255 6394
rect 19067 6363 19103 6364
rect 18480 6343 18521 6351
rect 18410 6337 18521 6343
rect 17738 6316 18185 6323
rect 17738 6314 17906 6316
rect 16586 6283 16696 6297
rect 16586 6280 16629 6283
rect 16586 6275 16590 6280
rect 16120 6245 16288 6247
rect 15844 6242 16288 6245
rect 15505 6218 15616 6224
rect 15505 6210 15546 6218
rect 15194 6155 15233 6199
rect 15505 6190 15513 6210
rect 15532 6190 15546 6210
rect 15505 6188 15546 6190
rect 15574 6210 15616 6218
rect 15574 6190 15590 6210
rect 15609 6190 15616 6210
rect 15574 6188 15616 6190
rect 15505 6173 15616 6188
rect 15842 6219 16288 6242
rect 15194 6131 15234 6155
rect 15534 6131 15581 6133
rect 15842 6131 15880 6219
rect 16120 6218 16288 6219
rect 16508 6253 16590 6275
rect 16619 6253 16629 6280
rect 16657 6256 16664 6283
rect 16693 6275 16696 6283
rect 16693 6256 16758 6275
rect 16657 6253 16758 6256
rect 16508 6251 16758 6253
rect 16508 6172 16545 6251
rect 16586 6238 16696 6251
rect 16660 6182 16691 6183
rect 16508 6152 16517 6172
rect 16537 6152 16545 6172
rect 16508 6142 16545 6152
rect 16604 6172 16691 6182
rect 16604 6152 16613 6172
rect 16633 6152 16691 6172
rect 16604 6143 16691 6152
rect 16604 6142 16641 6143
rect 15194 6098 15880 6131
rect 15194 6041 15233 6098
rect 15842 6096 15880 6098
rect 16660 6090 16691 6143
rect 16721 6172 16758 6251
rect 16929 6264 17322 6268
rect 16929 6247 16948 6264
rect 16968 6248 17322 6264
rect 17342 6248 17345 6268
rect 16968 6247 17345 6248
rect 16929 6243 17345 6247
rect 16929 6242 17270 6243
rect 16873 6182 16904 6183
rect 16721 6152 16730 6172
rect 16750 6152 16758 6172
rect 16721 6142 16758 6152
rect 16817 6175 16904 6182
rect 16817 6172 16878 6175
rect 16817 6152 16826 6172
rect 16846 6155 16878 6172
rect 16899 6155 16904 6175
rect 16846 6152 16904 6155
rect 16817 6145 16904 6152
rect 16929 6172 16966 6242
rect 17232 6241 17269 6242
rect 17081 6182 17117 6183
rect 16929 6152 16938 6172
rect 16958 6152 16966 6172
rect 16817 6143 16873 6145
rect 16817 6142 16854 6143
rect 16929 6142 16966 6152
rect 17025 6172 17173 6182
rect 17341 6181 17370 6182
rect 17273 6179 17370 6181
rect 17025 6152 17034 6172
rect 17054 6168 17144 6172
rect 17054 6152 17087 6168
rect 17025 6143 17087 6152
rect 17025 6142 17062 6143
rect 17081 6130 17087 6143
rect 17110 6152 17144 6168
rect 17164 6152 17173 6172
rect 17110 6143 17173 6152
rect 17231 6172 17370 6179
rect 17231 6152 17240 6172
rect 17260 6152 17370 6172
rect 17231 6143 17370 6152
rect 17110 6130 17117 6143
rect 17136 6142 17173 6143
rect 17232 6142 17269 6143
rect 17081 6091 17117 6130
rect 16552 6089 16593 6090
rect 16444 6082 16593 6089
rect 16444 6062 16562 6082
rect 16582 6062 16593 6082
rect 16444 6054 16593 6062
rect 16660 6086 17019 6090
rect 16660 6081 16982 6086
rect 16660 6057 16773 6081
rect 16797 6062 16982 6081
rect 17006 6062 17019 6086
rect 16797 6057 17019 6062
rect 16660 6054 17019 6057
rect 17081 6054 17116 6091
rect 17184 6088 17284 6091
rect 17184 6084 17251 6088
rect 17184 6058 17196 6084
rect 17222 6062 17251 6084
rect 17277 6062 17284 6088
rect 17222 6058 17284 6062
rect 17184 6054 17284 6058
rect 15194 6039 15242 6041
rect 15194 6021 15205 6039
rect 15223 6021 15242 6039
rect 16660 6033 16691 6054
rect 17081 6033 17117 6054
rect 16503 6032 16540 6033
rect 15194 6012 15242 6021
rect 15195 6011 15242 6012
rect 15508 6016 15618 6030
rect 15508 6013 15551 6016
rect 15508 6008 15512 6013
rect 15430 5986 15512 6008
rect 15541 5986 15551 6013
rect 15579 5989 15586 6016
rect 15615 6008 15618 6016
rect 16502 6023 16540 6032
rect 15615 5989 15680 6008
rect 16502 6003 16511 6023
rect 16531 6003 16540 6023
rect 15579 5986 15680 5989
rect 15430 5984 15680 5986
rect 15198 5948 15235 5949
rect 14816 5841 14826 5859
rect 14844 5841 14856 5859
rect 14816 5836 14856 5841
rect 15194 5945 15235 5948
rect 15194 5940 15236 5945
rect 15194 5922 15207 5940
rect 15225 5922 15236 5940
rect 15194 5908 15236 5922
rect 15274 5908 15321 5912
rect 15194 5902 15321 5908
rect 15194 5873 15282 5902
rect 15311 5873 15321 5902
rect 15430 5905 15467 5984
rect 15508 5971 15618 5984
rect 15582 5915 15613 5916
rect 15430 5885 15439 5905
rect 15459 5885 15467 5905
rect 15430 5875 15467 5885
rect 15526 5905 15613 5915
rect 15526 5885 15535 5905
rect 15555 5885 15613 5905
rect 15526 5876 15613 5885
rect 15526 5875 15563 5876
rect 15194 5869 15321 5873
rect 15194 5852 15233 5869
rect 15274 5868 15321 5869
rect 14816 5832 14853 5836
rect 15194 5834 15205 5852
rect 15223 5834 15233 5852
rect 15194 5825 15233 5834
rect 15195 5824 15232 5825
rect 15582 5823 15613 5876
rect 15643 5905 15680 5984
rect 15851 5981 16244 6001
rect 16264 5981 16267 6001
rect 16502 5995 16540 6003
rect 16606 6027 16691 6033
rect 16716 6032 16753 6033
rect 16606 6007 16614 6027
rect 16634 6007 16691 6027
rect 16606 5999 16691 6007
rect 16715 6023 16753 6032
rect 16715 6003 16724 6023
rect 16744 6003 16753 6023
rect 16606 5998 16642 5999
rect 16715 5995 16753 6003
rect 16819 6027 16904 6033
rect 16924 6032 16961 6033
rect 16819 6007 16827 6027
rect 16847 6026 16904 6027
rect 16847 6007 16876 6026
rect 16819 6006 16876 6007
rect 16897 6006 16904 6026
rect 16819 5999 16904 6006
rect 16923 6023 16961 6032
rect 16923 6003 16932 6023
rect 16952 6003 16961 6023
rect 16819 5998 16855 5999
rect 16923 5995 16961 6003
rect 17027 6027 17171 6033
rect 17027 6007 17035 6027
rect 17055 6007 17143 6027
rect 17163 6007 17171 6027
rect 17027 5999 17171 6007
rect 17027 5998 17063 5999
rect 17135 5998 17171 5999
rect 17237 6032 17274 6033
rect 17237 6031 17275 6032
rect 17237 6023 17301 6031
rect 17237 6003 17246 6023
rect 17266 6009 17301 6023
rect 17321 6009 17324 6029
rect 17266 6004 17324 6009
rect 17266 6003 17301 6004
rect 15851 5976 16267 5981
rect 15851 5975 16192 5976
rect 15795 5915 15826 5916
rect 15643 5885 15652 5905
rect 15672 5885 15680 5905
rect 15643 5875 15680 5885
rect 15739 5908 15826 5915
rect 15739 5905 15800 5908
rect 15739 5885 15748 5905
rect 15768 5888 15800 5905
rect 15821 5888 15826 5908
rect 15768 5885 15826 5888
rect 15739 5878 15826 5885
rect 15851 5905 15888 5975
rect 16154 5974 16191 5975
rect 16503 5966 16540 5995
rect 16504 5964 16540 5966
rect 16716 5964 16753 5995
rect 16504 5942 16753 5964
rect 16924 5963 16961 5995
rect 17237 5991 17301 6003
rect 17341 5965 17370 6143
rect 17738 6136 17765 6314
rect 17805 6276 17869 6288
rect 18145 6284 18182 6316
rect 18353 6315 18602 6337
rect 18353 6284 18390 6315
rect 18566 6313 18602 6315
rect 18566 6284 18603 6313
rect 18915 6304 18952 6305
rect 19218 6304 19255 6374
rect 19280 6394 19367 6401
rect 19280 6391 19338 6394
rect 19280 6371 19285 6391
rect 19306 6374 19338 6391
rect 19358 6374 19367 6394
rect 19306 6371 19367 6374
rect 19280 6364 19367 6371
rect 19426 6394 19463 6404
rect 19426 6374 19434 6394
rect 19454 6374 19463 6394
rect 19280 6363 19311 6364
rect 18914 6303 19255 6304
rect 18839 6298 19255 6303
rect 17805 6275 17840 6276
rect 17782 6270 17840 6275
rect 17782 6250 17785 6270
rect 17805 6256 17840 6270
rect 17860 6256 17869 6276
rect 17805 6248 17869 6256
rect 17831 6247 17869 6248
rect 17832 6246 17869 6247
rect 17935 6280 17971 6281
rect 18043 6280 18079 6281
rect 17935 6275 18079 6280
rect 17935 6272 17995 6275
rect 17935 6252 17943 6272
rect 17963 6254 17995 6272
rect 18022 6272 18079 6275
rect 18022 6254 18051 6272
rect 17963 6252 18051 6254
rect 18071 6252 18079 6272
rect 17935 6246 18079 6252
rect 18145 6276 18183 6284
rect 18251 6280 18287 6281
rect 18145 6256 18154 6276
rect 18174 6256 18183 6276
rect 18145 6247 18183 6256
rect 18202 6273 18287 6280
rect 18202 6253 18209 6273
rect 18230 6272 18287 6273
rect 18230 6253 18259 6272
rect 18202 6252 18259 6253
rect 18279 6252 18287 6272
rect 18145 6246 18182 6247
rect 18202 6246 18287 6252
rect 18353 6276 18391 6284
rect 18464 6280 18500 6281
rect 18353 6256 18362 6276
rect 18382 6256 18391 6276
rect 18353 6247 18391 6256
rect 18415 6272 18500 6280
rect 18415 6252 18472 6272
rect 18492 6252 18500 6272
rect 18353 6246 18390 6247
rect 18415 6246 18500 6252
rect 18566 6276 18604 6284
rect 18839 6278 18842 6298
rect 18862 6278 19255 6298
rect 19426 6295 19463 6374
rect 19493 6403 19524 6456
rect 19874 6454 19911 6455
rect 19873 6445 19912 6454
rect 19873 6427 19883 6445
rect 19901 6427 19912 6445
rect 19785 6410 19832 6411
rect 19873 6410 19912 6427
rect 19785 6406 19912 6410
rect 19543 6403 19580 6404
rect 19493 6394 19580 6403
rect 19493 6374 19551 6394
rect 19571 6374 19580 6394
rect 19493 6364 19580 6374
rect 19639 6394 19676 6404
rect 19639 6374 19647 6394
rect 19667 6374 19676 6394
rect 19493 6363 19524 6364
rect 19488 6295 19598 6308
rect 19639 6295 19676 6374
rect 19785 6377 19795 6406
rect 19824 6377 19912 6406
rect 19785 6371 19912 6377
rect 19785 6367 19832 6371
rect 19870 6357 19912 6371
rect 19870 6339 19881 6357
rect 19899 6339 19912 6357
rect 19870 6334 19912 6339
rect 19871 6331 19912 6334
rect 19871 6330 19908 6331
rect 19426 6293 19676 6295
rect 19426 6290 19527 6293
rect 18566 6256 18575 6276
rect 18595 6256 18604 6276
rect 19426 6271 19491 6290
rect 18566 6247 18604 6256
rect 19488 6263 19491 6271
rect 19520 6263 19527 6290
rect 19555 6266 19565 6293
rect 19594 6271 19676 6293
rect 19594 6266 19598 6271
rect 19555 6263 19598 6266
rect 19488 6249 19598 6263
rect 19864 6267 19911 6268
rect 19864 6258 19912 6267
rect 18566 6246 18603 6247
rect 17989 6225 18025 6246
rect 18415 6225 18446 6246
rect 19864 6240 19883 6258
rect 19901 6240 19912 6258
rect 19864 6238 19912 6240
rect 17822 6221 17922 6225
rect 17822 6217 17884 6221
rect 17822 6191 17829 6217
rect 17855 6195 17884 6217
rect 17910 6195 17922 6221
rect 17855 6191 17922 6195
rect 17822 6188 17922 6191
rect 17990 6188 18025 6225
rect 18087 6222 18446 6225
rect 18087 6217 18309 6222
rect 18087 6193 18100 6217
rect 18124 6198 18309 6217
rect 18333 6198 18446 6222
rect 18124 6193 18446 6198
rect 18087 6189 18446 6193
rect 18513 6217 18662 6225
rect 18513 6197 18524 6217
rect 18544 6197 18662 6217
rect 18513 6190 18662 6197
rect 18513 6189 18554 6190
rect 17837 6136 17874 6137
rect 17933 6136 17970 6137
rect 17989 6136 18025 6188
rect 18044 6136 18081 6137
rect 17737 6127 17875 6136
rect 17737 6107 17846 6127
rect 17866 6107 17875 6127
rect 17737 6100 17875 6107
rect 17933 6127 18081 6136
rect 17933 6107 17942 6127
rect 17962 6107 18052 6127
rect 18072 6107 18081 6127
rect 17737 6098 17833 6100
rect 17933 6097 18081 6107
rect 18140 6127 18177 6137
rect 18252 6136 18289 6137
rect 18233 6134 18289 6136
rect 18140 6107 18148 6127
rect 18168 6107 18177 6127
rect 17989 6096 18025 6097
rect 17837 6037 17874 6038
rect 18140 6037 18177 6107
rect 18202 6127 18289 6134
rect 18202 6124 18260 6127
rect 18202 6104 18207 6124
rect 18228 6107 18260 6124
rect 18280 6107 18289 6127
rect 18228 6104 18289 6107
rect 18202 6097 18289 6104
rect 18348 6127 18385 6137
rect 18348 6107 18356 6127
rect 18376 6107 18385 6127
rect 18202 6096 18233 6097
rect 17836 6036 18177 6037
rect 17761 6032 18177 6036
rect 17761 6031 18138 6032
rect 17761 6011 17764 6031
rect 17784 6015 18138 6031
rect 18158 6015 18177 6032
rect 17784 6011 18177 6015
rect 18348 6028 18385 6107
rect 18415 6136 18446 6189
rect 19226 6181 19264 6183
rect 19873 6181 19912 6238
rect 19226 6148 19912 6181
rect 18465 6136 18502 6137
rect 18415 6127 18502 6136
rect 18415 6107 18473 6127
rect 18493 6107 18502 6127
rect 18415 6097 18502 6107
rect 18561 6127 18598 6137
rect 18561 6107 18569 6127
rect 18589 6107 18598 6127
rect 18415 6096 18446 6097
rect 18410 6028 18520 6041
rect 18561 6028 18598 6107
rect 18348 6026 18598 6028
rect 18348 6023 18449 6026
rect 18348 6004 18413 6023
rect 18410 5996 18413 6004
rect 18442 5996 18449 6023
rect 18477 5999 18487 6026
rect 18516 6004 18598 6026
rect 18818 6060 18986 6061
rect 19226 6060 19264 6148
rect 19525 6146 19572 6148
rect 19872 6124 19912 6148
rect 18818 6037 19264 6060
rect 19490 6091 19601 6106
rect 19490 6089 19532 6091
rect 19490 6069 19497 6089
rect 19516 6069 19532 6089
rect 19490 6061 19532 6069
rect 19560 6089 19601 6091
rect 19560 6069 19574 6089
rect 19593 6069 19601 6089
rect 19873 6080 19912 6124
rect 19560 6061 19601 6069
rect 19490 6055 19601 6061
rect 18818 6034 19262 6037
rect 18818 6032 18986 6034
rect 18516 5999 18520 6004
rect 18477 5996 18520 5999
rect 18410 5982 18520 5996
rect 17200 5963 17370 5965
rect 16921 5956 17370 5963
rect 16585 5936 16696 5942
rect 16585 5928 16626 5936
rect 16003 5915 16039 5916
rect 15851 5885 15860 5905
rect 15880 5885 15888 5905
rect 15739 5876 15795 5878
rect 15739 5875 15776 5876
rect 15851 5875 15888 5885
rect 15947 5905 16095 5915
rect 16195 5912 16291 5914
rect 15947 5885 15956 5905
rect 15976 5885 16066 5905
rect 16086 5885 16095 5905
rect 15947 5876 16095 5885
rect 16153 5905 16291 5912
rect 16153 5885 16162 5905
rect 16182 5885 16291 5905
rect 16585 5908 16593 5928
rect 16612 5908 16626 5928
rect 16585 5906 16626 5908
rect 16654 5928 16696 5936
rect 16654 5908 16670 5928
rect 16689 5908 16696 5928
rect 16921 5929 16946 5956
rect 16977 5937 17370 5956
rect 16977 5929 17026 5937
rect 17200 5936 17370 5937
rect 16921 5927 17026 5929
rect 16654 5906 16696 5908
rect 16585 5891 16696 5906
rect 16153 5876 16291 5885
rect 15947 5875 15984 5876
rect 16003 5824 16039 5876
rect 16058 5875 16095 5876
rect 16154 5875 16191 5876
rect 15474 5822 15515 5823
rect 15366 5815 15515 5822
rect 14489 5813 14526 5814
rect 14439 5804 14526 5813
rect 14439 5784 14497 5804
rect 14517 5784 14526 5804
rect 14439 5774 14526 5784
rect 14585 5804 14622 5814
rect 14585 5784 14593 5804
rect 14613 5784 14622 5804
rect 15366 5795 15484 5815
rect 15504 5795 15515 5815
rect 15366 5787 15515 5795
rect 15582 5819 15941 5823
rect 15582 5814 15904 5819
rect 15582 5790 15695 5814
rect 15719 5795 15904 5814
rect 15928 5795 15941 5819
rect 15719 5790 15941 5795
rect 15582 5787 15941 5790
rect 16003 5787 16038 5824
rect 16106 5821 16206 5824
rect 16106 5817 16173 5821
rect 16106 5791 16118 5817
rect 16144 5795 16173 5817
rect 16199 5795 16206 5821
rect 16144 5791 16206 5795
rect 16106 5787 16206 5791
rect 14439 5773 14470 5774
rect 14434 5705 14544 5718
rect 14585 5705 14622 5784
rect 14819 5769 14856 5770
rect 14815 5760 14856 5769
rect 15582 5766 15613 5787
rect 16003 5766 16039 5787
rect 15425 5765 15462 5766
rect 15199 5762 15233 5763
rect 14815 5742 14828 5760
rect 14846 5742 14856 5760
rect 14815 5733 14856 5742
rect 15198 5753 15235 5762
rect 15198 5735 15207 5753
rect 15225 5735 15235 5753
rect 14815 5713 14855 5733
rect 15198 5725 15235 5735
rect 15424 5756 15462 5765
rect 15424 5736 15433 5756
rect 15453 5736 15462 5756
rect 15424 5728 15462 5736
rect 15528 5760 15613 5766
rect 15638 5765 15675 5766
rect 15528 5740 15536 5760
rect 15556 5740 15613 5760
rect 15528 5732 15613 5740
rect 15637 5756 15675 5765
rect 15637 5736 15646 5756
rect 15666 5736 15675 5756
rect 15528 5731 15564 5732
rect 15637 5728 15675 5736
rect 15741 5760 15826 5766
rect 15846 5765 15883 5766
rect 15741 5740 15749 5760
rect 15769 5759 15826 5760
rect 15769 5740 15798 5759
rect 15741 5739 15798 5740
rect 15819 5739 15826 5759
rect 15741 5732 15826 5739
rect 15845 5756 15883 5765
rect 15845 5736 15854 5756
rect 15874 5736 15883 5756
rect 15741 5731 15777 5732
rect 15845 5728 15883 5736
rect 15949 5760 16093 5766
rect 15949 5740 15957 5760
rect 15977 5759 16065 5760
rect 15977 5740 16008 5759
rect 15949 5739 16008 5740
rect 16033 5740 16065 5759
rect 16085 5740 16093 5760
rect 16033 5739 16093 5740
rect 15949 5732 16093 5739
rect 15949 5731 15985 5732
rect 16057 5731 16093 5732
rect 16159 5765 16196 5766
rect 16159 5764 16197 5765
rect 16159 5756 16223 5764
rect 16159 5736 16168 5756
rect 16188 5742 16223 5756
rect 16243 5742 16246 5762
rect 16188 5737 16246 5742
rect 16188 5736 16223 5737
rect 14372 5703 14622 5705
rect 14372 5700 14473 5703
rect 12890 5643 12954 5655
rect 13230 5651 13267 5678
rect 13438 5651 13475 5682
rect 13651 5680 13687 5682
rect 14372 5681 14437 5700
rect 13651 5651 13688 5680
rect 14434 5673 14437 5681
rect 14466 5673 14473 5700
rect 14501 5676 14511 5703
rect 14540 5681 14622 5703
rect 14730 5703 14855 5713
rect 14730 5684 14738 5703
rect 14763 5684 14855 5703
rect 14540 5676 14544 5681
rect 14730 5677 14855 5684
rect 14501 5673 14544 5676
rect 14434 5659 14544 5673
rect 12890 5642 12925 5643
rect 12867 5637 12925 5642
rect 12867 5617 12870 5637
rect 12890 5623 12925 5637
rect 12945 5623 12954 5643
rect 12890 5615 12954 5623
rect 12916 5614 12954 5615
rect 12917 5613 12954 5614
rect 13020 5647 13056 5648
rect 13128 5647 13164 5648
rect 13020 5639 13164 5647
rect 13020 5619 13028 5639
rect 13048 5636 13136 5639
rect 13048 5619 13080 5636
rect 13100 5619 13136 5636
rect 13156 5619 13164 5639
rect 13020 5613 13164 5619
rect 13230 5643 13268 5651
rect 13336 5647 13372 5648
rect 13230 5623 13239 5643
rect 13259 5623 13268 5643
rect 13230 5614 13268 5623
rect 13287 5640 13372 5647
rect 13287 5620 13294 5640
rect 13315 5639 13372 5640
rect 13315 5620 13344 5639
rect 13287 5619 13344 5620
rect 13364 5619 13372 5639
rect 13230 5613 13267 5614
rect 13287 5613 13372 5619
rect 13438 5643 13476 5651
rect 13549 5647 13585 5648
rect 13438 5623 13447 5643
rect 13467 5623 13476 5643
rect 13438 5614 13476 5623
rect 13500 5639 13585 5647
rect 13500 5619 13557 5639
rect 13577 5619 13585 5639
rect 13438 5613 13475 5614
rect 13500 5613 13585 5619
rect 13651 5643 13689 5651
rect 13651 5623 13660 5643
rect 13680 5623 13689 5643
rect 13651 5614 13689 5623
rect 14815 5629 14855 5677
rect 15199 5697 15233 5725
rect 15425 5699 15462 5728
rect 15426 5697 15462 5699
rect 15638 5697 15675 5728
rect 15199 5696 15371 5697
rect 15199 5664 15385 5696
rect 15426 5675 15675 5697
rect 15846 5696 15883 5728
rect 16159 5724 16223 5736
rect 16263 5698 16290 5876
rect 18818 5854 18845 6032
rect 18885 5994 18949 6006
rect 19225 6002 19262 6034
rect 19433 6033 19682 6055
rect 19433 6002 19470 6033
rect 19646 6031 19682 6033
rect 19646 6002 19683 6031
rect 18885 5993 18920 5994
rect 18862 5988 18920 5993
rect 18862 5968 18865 5988
rect 18885 5974 18920 5988
rect 18940 5974 18949 5994
rect 18885 5966 18949 5974
rect 18911 5965 18949 5966
rect 18912 5964 18949 5965
rect 19015 5998 19051 5999
rect 19123 5998 19159 5999
rect 19015 5993 19159 5998
rect 19015 5990 19077 5993
rect 19015 5970 19023 5990
rect 19043 5973 19077 5990
rect 19100 5990 19159 5993
rect 19100 5973 19131 5990
rect 19043 5970 19131 5973
rect 19151 5970 19159 5990
rect 19015 5964 19159 5970
rect 19225 5994 19263 6002
rect 19331 5998 19367 5999
rect 19225 5974 19234 5994
rect 19254 5974 19263 5994
rect 19225 5965 19263 5974
rect 19282 5991 19367 5998
rect 19282 5971 19289 5991
rect 19310 5990 19367 5991
rect 19310 5971 19339 5990
rect 19282 5970 19339 5971
rect 19359 5970 19367 5990
rect 19225 5964 19262 5965
rect 19282 5964 19367 5970
rect 19433 5994 19471 6002
rect 19544 5998 19580 5999
rect 19433 5974 19442 5994
rect 19462 5974 19471 5994
rect 19433 5965 19471 5974
rect 19495 5990 19580 5998
rect 19495 5970 19552 5990
rect 19572 5970 19580 5990
rect 19433 5964 19470 5965
rect 19495 5964 19580 5970
rect 19646 5994 19684 6002
rect 19646 5974 19655 5994
rect 19675 5974 19684 5994
rect 19646 5965 19684 5974
rect 19646 5964 19683 5965
rect 19069 5943 19105 5964
rect 19495 5943 19526 5964
rect 18902 5939 19002 5943
rect 18902 5935 18964 5939
rect 18902 5909 18909 5935
rect 18935 5913 18964 5935
rect 18990 5913 19002 5939
rect 18935 5909 19002 5913
rect 18902 5906 19002 5909
rect 19070 5906 19105 5943
rect 19167 5940 19526 5943
rect 19167 5935 19389 5940
rect 19167 5911 19180 5935
rect 19204 5916 19389 5935
rect 19413 5916 19526 5940
rect 19204 5911 19526 5916
rect 19167 5907 19526 5911
rect 19593 5935 19742 5943
rect 19593 5915 19604 5935
rect 19624 5915 19742 5935
rect 19593 5908 19742 5915
rect 19593 5907 19634 5908
rect 18917 5854 18954 5855
rect 19013 5854 19050 5855
rect 19069 5854 19105 5906
rect 19124 5854 19161 5855
rect 18817 5845 18955 5854
rect 18817 5825 18926 5845
rect 18946 5825 18955 5845
rect 18817 5818 18955 5825
rect 19013 5845 19161 5854
rect 19013 5825 19022 5845
rect 19042 5825 19132 5845
rect 19152 5825 19161 5845
rect 18817 5816 18913 5818
rect 19013 5815 19161 5825
rect 19220 5845 19257 5855
rect 19332 5854 19369 5855
rect 19313 5852 19369 5854
rect 19220 5825 19228 5845
rect 19248 5825 19257 5845
rect 19069 5814 19105 5815
rect 16446 5772 16556 5786
rect 16446 5769 16489 5772
rect 16446 5764 16450 5769
rect 16122 5696 16290 5698
rect 15846 5690 16290 5696
rect 15199 5632 15233 5664
rect 13651 5613 13688 5614
rect 13074 5592 13110 5613
rect 13500 5592 13531 5613
rect 14815 5611 14826 5629
rect 14844 5611 14855 5629
rect 14815 5603 14855 5611
rect 15195 5623 15233 5632
rect 15195 5605 15205 5623
rect 15223 5605 15233 5623
rect 14816 5602 14853 5603
rect 15195 5599 15233 5605
rect 15351 5601 15385 5664
rect 15507 5669 15618 5675
rect 15507 5661 15548 5669
rect 15507 5641 15515 5661
rect 15534 5641 15548 5661
rect 15507 5639 15548 5641
rect 15576 5661 15618 5669
rect 15576 5641 15592 5661
rect 15611 5641 15618 5661
rect 15576 5639 15618 5641
rect 15507 5624 15618 5639
rect 15845 5670 16290 5690
rect 15845 5601 15883 5670
rect 16122 5669 16290 5670
rect 16368 5742 16450 5764
rect 16479 5742 16489 5769
rect 16517 5745 16524 5772
rect 16553 5764 16556 5772
rect 18551 5781 18662 5796
rect 18551 5779 18593 5781
rect 16553 5745 16618 5764
rect 16517 5742 16618 5745
rect 16368 5740 16618 5742
rect 16368 5661 16405 5740
rect 16446 5727 16556 5740
rect 16520 5671 16551 5672
rect 16368 5641 16377 5661
rect 16397 5641 16405 5661
rect 16368 5631 16405 5641
rect 16464 5661 16551 5671
rect 16464 5641 16473 5661
rect 16493 5641 16551 5661
rect 16464 5632 16551 5641
rect 16464 5631 16501 5632
rect 15195 5595 15232 5599
rect 12907 5588 13007 5592
rect 12907 5584 12969 5588
rect 12907 5558 12914 5584
rect 12940 5562 12969 5584
rect 12995 5562 13007 5588
rect 12940 5558 13007 5562
rect 12907 5555 13007 5558
rect 13075 5555 13110 5592
rect 13172 5589 13531 5592
rect 13172 5584 13394 5589
rect 13172 5560 13185 5584
rect 13209 5565 13394 5584
rect 13418 5565 13531 5589
rect 13209 5560 13531 5565
rect 13172 5556 13531 5560
rect 13598 5584 13747 5592
rect 15351 5590 15883 5601
rect 13598 5564 13609 5584
rect 13629 5564 13747 5584
rect 15350 5574 15883 5590
rect 16520 5579 16551 5632
rect 16581 5661 16618 5740
rect 16789 5750 17182 5757
rect 16789 5733 16797 5750
rect 16829 5737 17182 5750
rect 17202 5737 17205 5757
rect 18284 5752 18325 5761
rect 16829 5733 17205 5737
rect 16789 5732 17205 5733
rect 17879 5750 18047 5751
rect 18284 5750 18293 5752
rect 16789 5731 17130 5732
rect 16733 5671 16764 5672
rect 16581 5641 16590 5661
rect 16610 5641 16618 5661
rect 16581 5631 16618 5641
rect 16677 5664 16764 5671
rect 16677 5661 16738 5664
rect 16677 5641 16686 5661
rect 16706 5644 16738 5661
rect 16759 5644 16764 5664
rect 16706 5641 16764 5644
rect 16677 5634 16764 5641
rect 16789 5661 16826 5731
rect 17092 5730 17129 5731
rect 17879 5730 18293 5750
rect 18319 5730 18325 5752
rect 18551 5759 18558 5779
rect 18577 5759 18593 5779
rect 18551 5751 18593 5759
rect 18621 5779 18662 5781
rect 18621 5759 18635 5779
rect 18654 5759 18662 5779
rect 18621 5751 18662 5759
rect 18917 5755 18954 5756
rect 19220 5755 19257 5825
rect 19282 5845 19369 5852
rect 19282 5842 19340 5845
rect 19282 5822 19287 5842
rect 19308 5825 19340 5842
rect 19360 5825 19369 5845
rect 19308 5822 19369 5825
rect 19282 5815 19369 5822
rect 19428 5845 19465 5855
rect 19428 5825 19436 5845
rect 19456 5825 19465 5845
rect 19282 5814 19313 5815
rect 18916 5754 19257 5755
rect 18551 5745 18662 5751
rect 18841 5749 19257 5754
rect 17879 5724 18325 5730
rect 17879 5722 18047 5724
rect 16941 5671 16977 5672
rect 16789 5641 16798 5661
rect 16818 5641 16826 5661
rect 16677 5632 16733 5634
rect 16677 5631 16714 5632
rect 16789 5631 16826 5641
rect 16885 5661 17033 5671
rect 17133 5668 17229 5670
rect 16885 5641 16894 5661
rect 16914 5656 17004 5661
rect 16914 5641 16949 5656
rect 16885 5632 16949 5641
rect 16885 5631 16922 5632
rect 16941 5615 16949 5632
rect 16970 5641 17004 5656
rect 17024 5641 17033 5661
rect 16970 5632 17033 5641
rect 17091 5661 17229 5668
rect 17091 5641 17100 5661
rect 17120 5641 17229 5661
rect 17091 5632 17229 5641
rect 16970 5615 16977 5632
rect 16996 5631 17033 5632
rect 17092 5631 17129 5632
rect 16941 5580 16977 5615
rect 16412 5578 16453 5579
rect 15350 5573 15864 5574
rect 13598 5557 13747 5564
rect 16304 5571 16453 5578
rect 14187 5561 14701 5562
rect 13598 5556 13639 5557
rect 12922 5503 12959 5504
rect 13018 5503 13055 5504
rect 13074 5503 13110 5555
rect 13129 5503 13166 5504
rect 12822 5494 12960 5503
rect 12822 5474 12931 5494
rect 12951 5474 12960 5494
rect 12822 5467 12960 5474
rect 13018 5494 13166 5503
rect 13018 5474 13027 5494
rect 13047 5474 13137 5494
rect 13157 5474 13166 5494
rect 12822 5465 12918 5467
rect 13018 5464 13166 5474
rect 13225 5494 13262 5504
rect 13337 5503 13374 5504
rect 13318 5501 13374 5503
rect 13225 5474 13233 5494
rect 13253 5474 13262 5494
rect 13074 5463 13110 5464
rect 12004 5411 12172 5413
rect 11726 5405 12172 5411
rect 10794 5381 11210 5386
rect 11389 5384 11500 5390
rect 10794 5380 11135 5381
rect 10738 5320 10769 5321
rect 10586 5290 10595 5310
rect 10615 5290 10623 5310
rect 10586 5280 10623 5290
rect 10682 5313 10769 5320
rect 10682 5310 10743 5313
rect 10682 5290 10691 5310
rect 10711 5293 10743 5310
rect 10764 5293 10769 5313
rect 10711 5290 10769 5293
rect 10682 5283 10769 5290
rect 10794 5310 10831 5380
rect 11097 5379 11134 5380
rect 11389 5376 11430 5384
rect 11389 5356 11397 5376
rect 11416 5356 11430 5376
rect 11389 5354 11430 5356
rect 11458 5376 11500 5384
rect 11458 5356 11474 5376
rect 11493 5356 11500 5376
rect 11726 5383 11732 5405
rect 11758 5385 12172 5405
rect 12922 5404 12959 5405
rect 13225 5404 13262 5474
rect 13287 5494 13374 5501
rect 13287 5491 13345 5494
rect 13287 5471 13292 5491
rect 13313 5474 13345 5491
rect 13365 5474 13374 5494
rect 13313 5471 13374 5474
rect 13287 5464 13374 5471
rect 13433 5494 13470 5504
rect 13433 5474 13441 5494
rect 13461 5474 13470 5494
rect 13287 5463 13318 5464
rect 12921 5403 13262 5404
rect 11758 5383 11767 5385
rect 12004 5384 12172 5385
rect 12846 5398 13262 5403
rect 11726 5374 11767 5383
rect 12846 5378 12849 5398
rect 12869 5378 13262 5398
rect 13433 5395 13470 5474
rect 13500 5503 13531 5556
rect 14168 5545 14701 5561
rect 16304 5551 16422 5571
rect 16442 5551 16453 5571
rect 14168 5534 14700 5545
rect 16304 5543 16453 5551
rect 16520 5575 16879 5579
rect 16520 5570 16842 5575
rect 16520 5546 16633 5570
rect 16657 5551 16842 5570
rect 16866 5551 16879 5575
rect 16657 5546 16879 5551
rect 16520 5543 16879 5546
rect 16941 5543 16976 5580
rect 17044 5577 17144 5580
rect 17044 5573 17111 5577
rect 17044 5547 17056 5573
rect 17082 5551 17111 5573
rect 17137 5551 17144 5577
rect 17082 5547 17144 5551
rect 17044 5543 17144 5547
rect 14819 5536 14856 5540
rect 13550 5503 13587 5504
rect 13500 5494 13587 5503
rect 13500 5474 13558 5494
rect 13578 5474 13587 5494
rect 13500 5464 13587 5474
rect 13646 5494 13683 5504
rect 13646 5474 13654 5494
rect 13674 5474 13683 5494
rect 13500 5463 13531 5464
rect 13495 5395 13605 5408
rect 13646 5395 13683 5474
rect 13433 5393 13683 5395
rect 13433 5390 13534 5393
rect 13433 5371 13498 5390
rect 13495 5363 13498 5371
rect 13527 5363 13534 5390
rect 13562 5366 13572 5393
rect 13601 5371 13683 5393
rect 13761 5465 13929 5466
rect 14168 5465 14206 5534
rect 13761 5445 14206 5465
rect 14433 5496 14544 5511
rect 14433 5494 14475 5496
rect 14433 5474 14440 5494
rect 14459 5474 14475 5494
rect 14433 5466 14475 5474
rect 14503 5494 14544 5496
rect 14503 5474 14517 5494
rect 14536 5474 14544 5494
rect 14503 5466 14544 5474
rect 14433 5460 14544 5466
rect 14666 5471 14700 5534
rect 14818 5530 14856 5536
rect 15198 5532 15235 5533
rect 14818 5512 14828 5530
rect 14846 5512 14856 5530
rect 14818 5503 14856 5512
rect 15196 5524 15236 5532
rect 15196 5506 15207 5524
rect 15225 5506 15236 5524
rect 16520 5522 16551 5543
rect 16941 5522 16977 5543
rect 16363 5521 16400 5522
rect 14818 5471 14852 5503
rect 13761 5439 14205 5445
rect 13761 5437 13929 5439
rect 13601 5366 13605 5371
rect 13562 5363 13605 5366
rect 11458 5354 11500 5356
rect 11389 5339 11500 5354
rect 12585 5345 12633 5359
rect 13495 5349 13605 5363
rect 10946 5320 10982 5321
rect 10794 5290 10803 5310
rect 10823 5290 10831 5310
rect 10682 5281 10738 5283
rect 10682 5280 10719 5281
rect 10794 5280 10831 5290
rect 10890 5310 11038 5320
rect 11138 5317 11234 5319
rect 10890 5290 10899 5310
rect 10919 5290 11009 5310
rect 11029 5290 11038 5310
rect 10890 5281 11038 5290
rect 11096 5310 11234 5317
rect 11096 5290 11105 5310
rect 11125 5290 11234 5310
rect 11096 5281 11234 5290
rect 12585 5305 12598 5345
rect 12625 5305 12633 5345
rect 12585 5287 12633 5305
rect 10890 5280 10927 5281
rect 10946 5229 10982 5281
rect 11001 5280 11038 5281
rect 11097 5280 11134 5281
rect 10417 5227 10458 5228
rect 10309 5220 10458 5227
rect 10309 5200 10427 5220
rect 10447 5200 10458 5220
rect 10309 5192 10458 5200
rect 10525 5224 10884 5228
rect 10525 5219 10847 5224
rect 10525 5195 10638 5219
rect 10662 5200 10847 5219
rect 10871 5200 10884 5224
rect 10662 5195 10884 5200
rect 10525 5192 10884 5195
rect 10946 5192 10981 5229
rect 11049 5226 11149 5229
rect 11049 5222 11116 5226
rect 11049 5196 11061 5222
rect 11087 5200 11116 5222
rect 11142 5200 11149 5226
rect 11087 5196 11149 5200
rect 11049 5192 11149 5196
rect 10525 5171 10556 5192
rect 10946 5171 10982 5192
rect 10368 5170 10405 5171
rect 10367 5161 10405 5170
rect 10367 5141 10376 5161
rect 10396 5141 10405 5161
rect 10367 5133 10405 5141
rect 10471 5165 10556 5171
rect 10581 5170 10618 5171
rect 10471 5145 10479 5165
rect 10499 5145 10556 5165
rect 10471 5137 10556 5145
rect 10580 5161 10618 5170
rect 10580 5141 10589 5161
rect 10609 5141 10618 5161
rect 10471 5136 10507 5137
rect 10580 5133 10618 5141
rect 10684 5165 10769 5171
rect 10789 5170 10826 5171
rect 10684 5145 10692 5165
rect 10712 5164 10769 5165
rect 10712 5145 10741 5164
rect 10684 5144 10741 5145
rect 10762 5144 10769 5164
rect 10684 5137 10769 5144
rect 10788 5161 10826 5170
rect 10788 5141 10797 5161
rect 10817 5141 10826 5161
rect 10684 5136 10720 5137
rect 10788 5133 10826 5141
rect 10892 5165 11036 5171
rect 10892 5145 10900 5165
rect 10920 5162 11008 5165
rect 10920 5145 10951 5162
rect 10892 5142 10951 5145
rect 10974 5145 11008 5162
rect 11028 5145 11036 5165
rect 10974 5142 11036 5145
rect 10892 5137 11036 5142
rect 10892 5136 10928 5137
rect 11000 5136 11036 5137
rect 11102 5170 11139 5171
rect 11102 5169 11140 5170
rect 11102 5161 11166 5169
rect 11102 5141 11111 5161
rect 11131 5147 11166 5161
rect 11186 5147 11189 5167
rect 11131 5142 11189 5147
rect 11131 5141 11166 5142
rect 10368 5104 10405 5133
rect 10369 5102 10405 5104
rect 10581 5102 10618 5133
rect 10369 5080 10618 5102
rect 10789 5101 10826 5133
rect 11102 5129 11166 5141
rect 11206 5103 11233 5281
rect 12580 5180 12633 5287
rect 13761 5259 13788 5437
rect 13828 5399 13892 5411
rect 14168 5407 14205 5439
rect 14376 5438 14625 5460
rect 14666 5439 14852 5471
rect 14680 5438 14852 5439
rect 14376 5407 14413 5438
rect 14589 5436 14625 5438
rect 14589 5407 14626 5436
rect 14818 5410 14852 5438
rect 15196 5458 15236 5506
rect 16362 5512 16400 5521
rect 16362 5492 16371 5512
rect 16391 5492 16400 5512
rect 16362 5484 16400 5492
rect 16466 5516 16551 5522
rect 16576 5521 16613 5522
rect 16466 5496 16474 5516
rect 16494 5496 16551 5516
rect 16466 5488 16551 5496
rect 16575 5512 16613 5521
rect 16575 5492 16584 5512
rect 16604 5492 16613 5512
rect 16466 5487 16502 5488
rect 16575 5484 16613 5492
rect 16679 5516 16764 5522
rect 16784 5521 16821 5522
rect 16679 5496 16687 5516
rect 16707 5515 16764 5516
rect 16707 5496 16736 5515
rect 16679 5495 16736 5496
rect 16757 5495 16764 5515
rect 16679 5488 16764 5495
rect 16783 5512 16821 5521
rect 16783 5492 16792 5512
rect 16812 5492 16821 5512
rect 16679 5487 16715 5488
rect 16783 5484 16821 5492
rect 16887 5516 17031 5522
rect 16887 5496 16895 5516
rect 16915 5496 17003 5516
rect 17023 5496 17031 5516
rect 16887 5488 17031 5496
rect 16887 5487 16923 5488
rect 16995 5487 17031 5488
rect 17097 5521 17134 5522
rect 17097 5520 17135 5521
rect 17097 5512 17161 5520
rect 17097 5492 17106 5512
rect 17126 5498 17161 5512
rect 17181 5498 17184 5518
rect 17126 5493 17184 5498
rect 17126 5492 17161 5493
rect 15507 5462 15617 5476
rect 15507 5459 15550 5462
rect 15196 5451 15321 5458
rect 15507 5454 15511 5459
rect 15196 5432 15288 5451
rect 15313 5432 15321 5451
rect 15196 5422 15321 5432
rect 15429 5432 15511 5454
rect 15540 5432 15550 5459
rect 15578 5435 15585 5462
rect 15614 5454 15617 5462
rect 16363 5455 16400 5484
rect 15614 5435 15679 5454
rect 16364 5453 16400 5455
rect 16576 5453 16613 5484
rect 16784 5457 16821 5484
rect 17097 5480 17161 5492
rect 15578 5432 15679 5435
rect 15429 5430 15679 5432
rect 13828 5398 13863 5399
rect 13805 5393 13863 5398
rect 13805 5373 13808 5393
rect 13828 5379 13863 5393
rect 13883 5379 13892 5399
rect 13828 5371 13892 5379
rect 13854 5370 13892 5371
rect 13855 5369 13892 5370
rect 13958 5403 13994 5404
rect 14066 5403 14102 5404
rect 13958 5396 14102 5403
rect 13958 5395 14018 5396
rect 13958 5375 13966 5395
rect 13986 5376 14018 5395
rect 14043 5395 14102 5396
rect 14043 5376 14074 5395
rect 13986 5375 14074 5376
rect 14094 5375 14102 5395
rect 13958 5369 14102 5375
rect 14168 5399 14206 5407
rect 14274 5403 14310 5404
rect 14168 5379 14177 5399
rect 14197 5379 14206 5399
rect 14168 5370 14206 5379
rect 14225 5396 14310 5403
rect 14225 5376 14232 5396
rect 14253 5395 14310 5396
rect 14253 5376 14282 5395
rect 14225 5375 14282 5376
rect 14302 5375 14310 5395
rect 14168 5369 14205 5370
rect 14225 5369 14310 5375
rect 14376 5399 14414 5407
rect 14487 5403 14523 5404
rect 14376 5379 14385 5399
rect 14405 5379 14414 5399
rect 14376 5370 14414 5379
rect 14438 5395 14523 5403
rect 14438 5375 14495 5395
rect 14515 5375 14523 5395
rect 14376 5369 14413 5370
rect 14438 5369 14523 5375
rect 14589 5399 14627 5407
rect 14589 5379 14598 5399
rect 14618 5379 14627 5399
rect 14589 5370 14627 5379
rect 14816 5400 14853 5410
rect 15196 5402 15236 5422
rect 14816 5382 14826 5400
rect 14844 5382 14853 5400
rect 14816 5373 14853 5382
rect 15195 5393 15236 5402
rect 15195 5375 15205 5393
rect 15223 5375 15236 5393
rect 14818 5372 14852 5373
rect 14589 5369 14626 5370
rect 14012 5348 14048 5369
rect 14438 5348 14469 5369
rect 15195 5366 15236 5375
rect 15195 5365 15232 5366
rect 15429 5351 15466 5430
rect 15507 5417 15617 5430
rect 15581 5361 15612 5362
rect 13845 5344 13945 5348
rect 13845 5340 13907 5344
rect 13845 5314 13852 5340
rect 13878 5318 13907 5340
rect 13933 5318 13945 5344
rect 13878 5314 13945 5318
rect 13845 5311 13945 5314
rect 14013 5311 14048 5348
rect 14110 5345 14469 5348
rect 14110 5340 14332 5345
rect 14110 5316 14123 5340
rect 14147 5321 14332 5340
rect 14356 5321 14469 5345
rect 14147 5316 14469 5321
rect 14110 5312 14469 5316
rect 14536 5340 14685 5348
rect 14536 5320 14547 5340
rect 14567 5320 14685 5340
rect 15429 5331 15438 5351
rect 15458 5331 15466 5351
rect 15429 5321 15466 5331
rect 15525 5351 15612 5361
rect 15525 5331 15534 5351
rect 15554 5331 15612 5351
rect 15525 5322 15612 5331
rect 15525 5321 15562 5322
rect 14536 5313 14685 5320
rect 14536 5312 14577 5313
rect 13860 5259 13897 5260
rect 13956 5259 13993 5260
rect 14012 5259 14048 5311
rect 14067 5259 14104 5260
rect 13760 5250 13898 5259
rect 13760 5230 13869 5250
rect 13889 5230 13898 5250
rect 13386 5210 13497 5225
rect 13760 5223 13898 5230
rect 13956 5250 14104 5259
rect 13956 5230 13965 5250
rect 13985 5230 14075 5250
rect 14095 5230 14104 5250
rect 13760 5221 13856 5223
rect 13956 5220 14104 5230
rect 14163 5250 14200 5260
rect 14275 5259 14312 5260
rect 14256 5257 14312 5259
rect 14163 5230 14171 5250
rect 14191 5230 14200 5250
rect 14012 5219 14048 5220
rect 13386 5208 13428 5210
rect 13386 5188 13393 5208
rect 13412 5188 13428 5208
rect 13386 5180 13428 5188
rect 13456 5208 13497 5210
rect 13456 5188 13470 5208
rect 13489 5188 13497 5208
rect 13456 5180 13497 5188
rect 12580 5179 12882 5180
rect 11499 5158 11609 5172
rect 11499 5155 11542 5158
rect 11499 5150 11503 5155
rect 11065 5101 11233 5103
rect 10789 5098 11233 5101
rect 10450 5074 10561 5080
rect 10450 5066 10491 5074
rect 9195 5040 9881 5050
rect 8466 5009 8503 5010
rect 8416 5000 8503 5009
rect 8416 4980 8474 5000
rect 8494 4980 8503 5000
rect 8416 4970 8503 4980
rect 8562 5000 8599 5010
rect 8562 4980 8570 5000
rect 8590 4980 8599 5000
rect 8416 4969 8447 4970
rect 8411 4901 8521 4914
rect 8562 4901 8599 4980
rect 8349 4899 8599 4901
rect 8349 4896 8450 4899
rect 8349 4877 8414 4896
rect 7254 4876 7440 4877
rect 7138 4874 7440 4876
rect 6523 4847 6634 4853
rect 6862 4848 7440 4874
rect 8411 4869 8414 4877
rect 8443 4869 8450 4896
rect 8478 4872 8488 4899
rect 8517 4877 8599 4899
rect 8787 4952 8955 4953
rect 9195 4952 9233 5040
rect 9494 5039 9541 5040
rect 9841 5016 9881 5040
rect 9458 4983 9570 5002
rect 9458 4982 9501 4983
rect 8787 4929 9233 4952
rect 9459 4981 9501 4982
rect 9459 4961 9466 4981
rect 9485 4961 9501 4981
rect 9459 4953 9501 4961
rect 9529 4981 9570 4983
rect 9529 4961 9543 4981
rect 9562 4961 9570 4981
rect 9842 4972 9881 5016
rect 10139 5011 10178 5055
rect 10450 5046 10458 5066
rect 10477 5046 10491 5066
rect 10450 5044 10491 5046
rect 10519 5066 10561 5074
rect 10519 5046 10535 5066
rect 10554 5046 10561 5066
rect 10519 5045 10561 5046
rect 10787 5075 11233 5098
rect 10519 5044 10562 5045
rect 10450 5025 10562 5044
rect 10139 4987 10179 5011
rect 10479 4987 10526 4988
rect 10787 4987 10825 5075
rect 11065 5074 11233 5075
rect 11421 5128 11503 5150
rect 11532 5128 11542 5155
rect 11570 5131 11577 5158
rect 11606 5150 11609 5158
rect 12580 5153 13158 5179
rect 13386 5174 13497 5180
rect 12580 5151 12882 5153
rect 12580 5150 12766 5151
rect 11606 5131 11671 5150
rect 11570 5128 11671 5131
rect 11421 5126 11671 5128
rect 11421 5047 11458 5126
rect 11499 5113 11609 5126
rect 11573 5057 11604 5058
rect 11421 5027 11430 5047
rect 11450 5027 11458 5047
rect 11421 5017 11458 5027
rect 11517 5047 11604 5057
rect 11517 5027 11526 5047
rect 11546 5027 11604 5047
rect 11517 5018 11604 5027
rect 11517 5017 11554 5018
rect 10139 4977 10825 4987
rect 9529 4953 9570 4961
rect 9459 4947 9570 4953
rect 8787 4926 9231 4929
rect 8787 4924 8955 4926
rect 8517 4872 8521 4877
rect 8478 4869 8521 4872
rect 8411 4855 8521 4869
rect 7138 4847 7440 4848
rect 6523 4839 6564 4847
rect 6523 4819 6531 4839
rect 6550 4819 6564 4839
rect 6523 4817 6564 4819
rect 6592 4839 6634 4847
rect 6592 4819 6608 4839
rect 6627 4819 6634 4839
rect 6592 4817 6634 4819
rect 5972 4807 6008 4808
rect 5820 4777 5829 4797
rect 5849 4777 5857 4797
rect 5708 4768 5764 4770
rect 5708 4767 5745 4768
rect 5820 4767 5857 4777
rect 5916 4797 6064 4807
rect 6164 4804 6260 4806
rect 5916 4777 5925 4797
rect 5945 4777 6035 4797
rect 6055 4777 6064 4797
rect 5916 4768 6064 4777
rect 6122 4797 6260 4804
rect 6523 4802 6634 4817
rect 6122 4777 6131 4797
rect 6151 4777 6260 4797
rect 6122 4768 6260 4777
rect 5916 4767 5953 4768
rect 5972 4716 6008 4768
rect 6027 4767 6064 4768
rect 6123 4767 6160 4768
rect 5443 4714 5484 4715
rect 5335 4707 5484 4714
rect 4458 4705 4495 4706
rect 4408 4696 4495 4705
rect 4408 4676 4466 4696
rect 4486 4676 4495 4696
rect 4408 4666 4495 4676
rect 4554 4696 4591 4706
rect 4554 4676 4562 4696
rect 4582 4676 4591 4696
rect 5335 4687 5453 4707
rect 5473 4687 5484 4707
rect 5335 4679 5484 4687
rect 5551 4711 5910 4715
rect 5551 4706 5873 4711
rect 5551 4682 5664 4706
rect 5688 4687 5873 4706
rect 5897 4687 5910 4711
rect 5688 4682 5910 4687
rect 5551 4679 5910 4682
rect 5972 4679 6007 4716
rect 6075 4713 6175 4716
rect 6075 4709 6142 4713
rect 6075 4683 6087 4709
rect 6113 4687 6142 4709
rect 6168 4687 6175 4713
rect 6113 4683 6175 4687
rect 6075 4679 6175 4683
rect 4408 4665 4439 4666
rect 4403 4597 4513 4610
rect 4554 4597 4591 4676
rect 4788 4661 4825 4662
rect 4784 4652 4825 4661
rect 5551 4658 5582 4679
rect 5972 4658 6008 4679
rect 5394 4657 5431 4658
rect 5168 4654 5202 4655
rect 4784 4634 4797 4652
rect 4815 4634 4825 4652
rect 4784 4625 4825 4634
rect 5167 4645 5204 4654
rect 5167 4627 5176 4645
rect 5194 4627 5204 4645
rect 4784 4605 4824 4625
rect 5167 4617 5204 4627
rect 5393 4648 5431 4657
rect 5393 4628 5402 4648
rect 5422 4628 5431 4648
rect 5393 4620 5431 4628
rect 5497 4652 5582 4658
rect 5607 4657 5644 4658
rect 5497 4632 5505 4652
rect 5525 4632 5582 4652
rect 5497 4624 5582 4632
rect 5606 4648 5644 4657
rect 5606 4628 5615 4648
rect 5635 4628 5644 4648
rect 5497 4623 5533 4624
rect 5606 4620 5644 4628
rect 5710 4652 5795 4658
rect 5815 4657 5852 4658
rect 5710 4632 5718 4652
rect 5738 4651 5795 4652
rect 5738 4632 5767 4651
rect 5710 4631 5767 4632
rect 5788 4631 5795 4651
rect 5710 4624 5795 4631
rect 5814 4648 5852 4657
rect 5814 4628 5823 4648
rect 5843 4628 5852 4648
rect 5710 4623 5746 4624
rect 5814 4620 5852 4628
rect 5918 4652 6062 4658
rect 5918 4632 5926 4652
rect 5946 4651 6034 4652
rect 5946 4632 5977 4651
rect 5918 4631 5977 4632
rect 6002 4632 6034 4651
rect 6054 4632 6062 4652
rect 6002 4631 6062 4632
rect 5918 4624 6062 4631
rect 5918 4623 5954 4624
rect 6026 4623 6062 4624
rect 6128 4657 6165 4658
rect 6128 4656 6166 4657
rect 6128 4648 6192 4656
rect 6128 4628 6137 4648
rect 6157 4634 6192 4648
rect 6212 4634 6215 4654
rect 6157 4629 6215 4634
rect 6157 4628 6192 4629
rect 4341 4595 4591 4597
rect 4341 4592 4442 4595
rect 2859 4535 2923 4547
rect 3199 4543 3236 4570
rect 3407 4543 3444 4574
rect 3620 4572 3656 4574
rect 4341 4573 4406 4592
rect 3620 4543 3657 4572
rect 4403 4565 4406 4573
rect 4435 4565 4442 4592
rect 4470 4568 4480 4595
rect 4509 4573 4591 4595
rect 4699 4595 4824 4605
rect 4699 4576 4707 4595
rect 4732 4576 4824 4595
rect 4509 4568 4513 4573
rect 4699 4569 4824 4576
rect 4470 4565 4513 4568
rect 4403 4551 4513 4565
rect 2859 4534 2894 4535
rect 2836 4529 2894 4534
rect 2836 4509 2839 4529
rect 2859 4515 2894 4529
rect 2914 4515 2923 4535
rect 2859 4507 2923 4515
rect 2885 4506 2923 4507
rect 2886 4505 2923 4506
rect 2989 4539 3025 4540
rect 3097 4539 3133 4540
rect 2989 4531 3133 4539
rect 2989 4511 2997 4531
rect 3017 4511 3105 4531
rect 3125 4511 3133 4531
rect 2989 4505 3133 4511
rect 3199 4535 3237 4543
rect 3305 4539 3341 4540
rect 3199 4515 3208 4535
rect 3228 4515 3237 4535
rect 3199 4506 3237 4515
rect 3256 4532 3341 4539
rect 3256 4512 3263 4532
rect 3284 4531 3341 4532
rect 3284 4512 3313 4531
rect 3256 4511 3313 4512
rect 3333 4511 3341 4531
rect 3199 4505 3236 4506
rect 3256 4505 3341 4511
rect 3407 4535 3445 4543
rect 3518 4539 3554 4540
rect 3407 4515 3416 4535
rect 3436 4515 3445 4535
rect 3407 4506 3445 4515
rect 3469 4531 3554 4539
rect 3469 4511 3526 4531
rect 3546 4511 3554 4531
rect 3407 4505 3444 4506
rect 3469 4505 3554 4511
rect 3620 4535 3658 4543
rect 3620 4515 3629 4535
rect 3649 4515 3658 4535
rect 3620 4506 3658 4515
rect 4784 4521 4824 4569
rect 5168 4589 5202 4617
rect 5394 4591 5431 4620
rect 5395 4589 5431 4591
rect 5607 4589 5644 4620
rect 5168 4588 5340 4589
rect 5168 4556 5354 4588
rect 5395 4567 5644 4589
rect 5815 4588 5852 4620
rect 6128 4616 6192 4628
rect 6232 4590 6259 4768
rect 7387 4740 7440 4847
rect 8787 4746 8814 4924
rect 8854 4886 8918 4898
rect 9194 4894 9231 4926
rect 9402 4925 9651 4947
rect 9402 4894 9439 4925
rect 9615 4923 9651 4925
rect 9615 4894 9652 4923
rect 8854 4885 8889 4886
rect 8831 4880 8889 4885
rect 8831 4860 8834 4880
rect 8854 4866 8889 4880
rect 8909 4866 8918 4886
rect 8854 4858 8918 4866
rect 8880 4857 8918 4858
rect 8881 4856 8918 4857
rect 8984 4890 9020 4891
rect 9092 4890 9128 4891
rect 8984 4885 9128 4890
rect 8984 4882 9046 4885
rect 8984 4862 8992 4882
rect 9012 4865 9046 4882
rect 9069 4882 9128 4885
rect 9069 4865 9100 4882
rect 9012 4862 9100 4865
rect 9120 4862 9128 4882
rect 8984 4856 9128 4862
rect 9194 4886 9232 4894
rect 9300 4890 9336 4891
rect 9194 4866 9203 4886
rect 9223 4866 9232 4886
rect 9194 4857 9232 4866
rect 9251 4883 9336 4890
rect 9251 4863 9258 4883
rect 9279 4882 9336 4883
rect 9279 4863 9308 4882
rect 9251 4862 9308 4863
rect 9328 4862 9336 4882
rect 9194 4856 9231 4857
rect 9251 4856 9336 4862
rect 9402 4886 9440 4894
rect 9513 4890 9549 4891
rect 9402 4866 9411 4886
rect 9431 4866 9440 4886
rect 9402 4857 9440 4866
rect 9464 4882 9549 4890
rect 9464 4862 9521 4882
rect 9541 4862 9549 4882
rect 9402 4856 9439 4857
rect 9464 4856 9549 4862
rect 9615 4886 9653 4894
rect 9615 4866 9624 4886
rect 9644 4866 9653 4886
rect 9615 4857 9653 4866
rect 9615 4856 9652 4857
rect 9038 4835 9074 4856
rect 9464 4835 9495 4856
rect 8871 4831 8971 4835
rect 8871 4827 8933 4831
rect 8871 4801 8878 4827
rect 8904 4805 8933 4827
rect 8959 4805 8971 4831
rect 8904 4801 8971 4805
rect 8871 4798 8971 4801
rect 9039 4798 9074 4835
rect 9136 4832 9495 4835
rect 9136 4827 9358 4832
rect 9136 4803 9149 4827
rect 9173 4808 9358 4827
rect 9382 4808 9495 4832
rect 9173 4803 9495 4808
rect 9136 4799 9495 4803
rect 9562 4827 9711 4835
rect 9562 4807 9573 4827
rect 9593 4807 9711 4827
rect 9562 4800 9711 4807
rect 9562 4799 9603 4800
rect 8886 4746 8923 4747
rect 8982 4746 9019 4747
rect 9038 4746 9074 4798
rect 9093 4746 9130 4747
rect 7387 4722 7435 4740
rect 7387 4682 7395 4722
rect 7422 4682 7435 4722
rect 8786 4737 8924 4746
rect 8786 4717 8895 4737
rect 8915 4717 8924 4737
rect 8786 4710 8924 4717
rect 8982 4737 9130 4746
rect 8982 4717 8991 4737
rect 9011 4717 9101 4737
rect 9121 4717 9130 4737
rect 8786 4708 8882 4710
rect 8982 4707 9130 4717
rect 9189 4737 9226 4747
rect 9301 4746 9338 4747
rect 9282 4744 9338 4746
rect 9189 4717 9197 4737
rect 9217 4717 9226 4737
rect 9038 4706 9074 4707
rect 6415 4664 6525 4678
rect 7387 4668 7435 4682
rect 8520 4673 8631 4688
rect 8520 4671 8562 4673
rect 6415 4661 6458 4664
rect 6415 4656 6419 4661
rect 6091 4588 6259 4590
rect 5815 4582 6259 4588
rect 5168 4524 5202 4556
rect 3620 4505 3657 4506
rect 3043 4484 3079 4505
rect 3469 4484 3500 4505
rect 4784 4503 4795 4521
rect 4813 4503 4824 4521
rect 4784 4495 4824 4503
rect 5164 4515 5202 4524
rect 5164 4497 5174 4515
rect 5192 4497 5202 4515
rect 4785 4494 4822 4495
rect 5164 4491 5202 4497
rect 5320 4493 5354 4556
rect 5476 4561 5587 4567
rect 5476 4553 5517 4561
rect 5476 4533 5484 4553
rect 5503 4533 5517 4553
rect 5476 4531 5517 4533
rect 5545 4553 5587 4561
rect 5545 4533 5561 4553
rect 5580 4533 5587 4553
rect 5545 4531 5587 4533
rect 5476 4516 5587 4531
rect 5814 4562 6259 4582
rect 5814 4493 5852 4562
rect 6091 4561 6259 4562
rect 6337 4634 6419 4656
rect 6448 4634 6458 4661
rect 6486 4637 6493 4664
rect 6522 4656 6525 4664
rect 6522 4637 6587 4656
rect 6486 4634 6587 4637
rect 6337 4632 6587 4634
rect 6337 4553 6374 4632
rect 6415 4619 6525 4632
rect 6489 4563 6520 4564
rect 6337 4533 6346 4553
rect 6366 4533 6374 4553
rect 6337 4523 6374 4533
rect 6433 4553 6520 4563
rect 6433 4533 6442 4553
rect 6462 4533 6520 4553
rect 6433 4524 6520 4533
rect 6433 4523 6470 4524
rect 5164 4487 5201 4491
rect 2876 4480 2976 4484
rect 2876 4476 2938 4480
rect 2876 4450 2883 4476
rect 2909 4454 2938 4476
rect 2964 4454 2976 4480
rect 2909 4450 2976 4454
rect 2876 4447 2976 4450
rect 3044 4447 3079 4484
rect 3141 4481 3500 4484
rect 3141 4476 3363 4481
rect 3141 4452 3154 4476
rect 3178 4457 3363 4476
rect 3387 4457 3500 4481
rect 3178 4452 3500 4457
rect 3141 4448 3500 4452
rect 3567 4476 3716 4484
rect 5320 4482 5852 4493
rect 3567 4456 3578 4476
rect 3598 4456 3716 4476
rect 5319 4466 5852 4482
rect 6489 4471 6520 4524
rect 6550 4553 6587 4632
rect 6758 4629 7151 4649
rect 7171 4629 7174 4649
rect 8253 4644 8294 4653
rect 6758 4624 7174 4629
rect 7848 4642 8016 4643
rect 8253 4642 8262 4644
rect 6758 4623 7099 4624
rect 6702 4563 6733 4564
rect 6550 4533 6559 4553
rect 6579 4533 6587 4553
rect 6550 4523 6587 4533
rect 6646 4556 6733 4563
rect 6646 4553 6707 4556
rect 6646 4533 6655 4553
rect 6675 4536 6707 4553
rect 6728 4536 6733 4556
rect 6675 4533 6733 4536
rect 6646 4526 6733 4533
rect 6758 4553 6795 4623
rect 7061 4622 7098 4623
rect 7848 4622 8262 4642
rect 8288 4622 8294 4644
rect 8520 4651 8527 4671
rect 8546 4651 8562 4671
rect 8520 4643 8562 4651
rect 8590 4671 8631 4673
rect 8590 4651 8604 4671
rect 8623 4651 8631 4671
rect 8590 4643 8631 4651
rect 8886 4647 8923 4648
rect 9189 4647 9226 4717
rect 9251 4737 9338 4744
rect 9251 4734 9309 4737
rect 9251 4714 9256 4734
rect 9277 4717 9309 4734
rect 9329 4717 9338 4737
rect 9277 4714 9338 4717
rect 9251 4707 9338 4714
rect 9397 4737 9434 4747
rect 9397 4717 9405 4737
rect 9425 4717 9434 4737
rect 9251 4706 9282 4707
rect 8885 4646 9226 4647
rect 8520 4637 8631 4643
rect 8810 4641 9226 4646
rect 7848 4616 8294 4622
rect 7848 4614 8016 4616
rect 6910 4563 6946 4564
rect 6758 4533 6767 4553
rect 6787 4533 6795 4553
rect 6646 4524 6702 4526
rect 6646 4523 6683 4524
rect 6758 4523 6795 4533
rect 6854 4553 7002 4563
rect 7102 4560 7198 4562
rect 6854 4533 6863 4553
rect 6883 4533 6973 4553
rect 6993 4533 7002 4553
rect 6854 4524 7002 4533
rect 7060 4553 7198 4560
rect 7060 4533 7069 4553
rect 7089 4533 7198 4553
rect 7060 4524 7198 4533
rect 6854 4523 6891 4524
rect 6910 4472 6946 4524
rect 6965 4523 7002 4524
rect 7061 4523 7098 4524
rect 6381 4470 6422 4471
rect 5319 4465 5833 4466
rect 3567 4449 3716 4456
rect 6273 4463 6422 4470
rect 4156 4453 4670 4454
rect 3567 4448 3608 4449
rect 3043 4412 3079 4447
rect 2891 4395 2928 4396
rect 2987 4395 3024 4396
rect 3043 4395 3050 4412
rect 2791 4386 2929 4395
rect 2791 4366 2900 4386
rect 2920 4366 2929 4386
rect 2791 4359 2929 4366
rect 2987 4386 3050 4395
rect 2987 4366 2996 4386
rect 3016 4371 3050 4386
rect 3071 4395 3079 4412
rect 3098 4395 3135 4396
rect 3071 4386 3135 4395
rect 3071 4371 3106 4386
rect 3016 4366 3106 4371
rect 3126 4366 3135 4386
rect 2791 4357 2887 4359
rect 2987 4356 3135 4366
rect 3194 4386 3231 4396
rect 3306 4395 3343 4396
rect 3287 4393 3343 4395
rect 3194 4366 3202 4386
rect 3222 4366 3231 4386
rect 3043 4355 3079 4356
rect 1973 4303 2141 4305
rect 1695 4297 2141 4303
rect 763 4273 1179 4278
rect 1358 4276 1469 4282
rect 763 4272 1104 4273
rect 707 4212 738 4213
rect 555 4182 564 4202
rect 584 4182 592 4202
rect 555 4172 592 4182
rect 651 4205 738 4212
rect 651 4202 712 4205
rect 651 4182 660 4202
rect 680 4185 712 4202
rect 733 4185 738 4205
rect 680 4182 738 4185
rect 651 4175 738 4182
rect 763 4202 800 4272
rect 1066 4271 1103 4272
rect 1358 4268 1399 4276
rect 1358 4248 1366 4268
rect 1385 4248 1399 4268
rect 1358 4246 1399 4248
rect 1427 4268 1469 4276
rect 1427 4248 1443 4268
rect 1462 4248 1469 4268
rect 1695 4275 1701 4297
rect 1727 4277 2141 4297
rect 2891 4296 2928 4297
rect 3194 4296 3231 4366
rect 3256 4386 3343 4393
rect 3256 4383 3314 4386
rect 3256 4363 3261 4383
rect 3282 4366 3314 4383
rect 3334 4366 3343 4386
rect 3282 4363 3343 4366
rect 3256 4356 3343 4363
rect 3402 4386 3439 4396
rect 3402 4366 3410 4386
rect 3430 4366 3439 4386
rect 3256 4355 3287 4356
rect 2890 4295 3231 4296
rect 1727 4275 1736 4277
rect 1973 4276 2141 4277
rect 2815 4294 3231 4295
rect 2815 4290 3191 4294
rect 1695 4266 1736 4275
rect 2815 4270 2818 4290
rect 2838 4277 3191 4290
rect 3223 4277 3231 4294
rect 2838 4270 3231 4277
rect 3402 4287 3439 4366
rect 3469 4395 3500 4448
rect 4137 4437 4670 4453
rect 6273 4443 6391 4463
rect 6411 4443 6422 4463
rect 4137 4426 4669 4437
rect 6273 4435 6422 4443
rect 6489 4467 6848 4471
rect 6489 4462 6811 4467
rect 6489 4438 6602 4462
rect 6626 4443 6811 4462
rect 6835 4443 6848 4467
rect 6626 4438 6848 4443
rect 6489 4435 6848 4438
rect 6910 4435 6945 4472
rect 7013 4469 7113 4472
rect 7013 4465 7080 4469
rect 7013 4439 7025 4465
rect 7051 4443 7080 4465
rect 7106 4443 7113 4469
rect 7051 4439 7113 4443
rect 7013 4435 7113 4439
rect 4788 4428 4825 4432
rect 3519 4395 3556 4396
rect 3469 4386 3556 4395
rect 3469 4366 3527 4386
rect 3547 4366 3556 4386
rect 3469 4356 3556 4366
rect 3615 4386 3652 4396
rect 3615 4366 3623 4386
rect 3643 4366 3652 4386
rect 3469 4355 3500 4356
rect 3464 4287 3574 4300
rect 3615 4287 3652 4366
rect 3402 4285 3652 4287
rect 3402 4282 3503 4285
rect 3402 4263 3467 4282
rect 1427 4246 1469 4248
rect 1358 4231 1469 4246
rect 3464 4255 3467 4263
rect 3496 4255 3503 4282
rect 3531 4258 3541 4285
rect 3570 4263 3652 4285
rect 3730 4357 3898 4358
rect 4137 4357 4175 4426
rect 3730 4337 4175 4357
rect 4402 4388 4513 4403
rect 4402 4386 4444 4388
rect 4402 4366 4409 4386
rect 4428 4366 4444 4386
rect 4402 4358 4444 4366
rect 4472 4386 4513 4388
rect 4472 4366 4486 4386
rect 4505 4366 4513 4386
rect 4472 4358 4513 4366
rect 4402 4352 4513 4358
rect 4635 4363 4669 4426
rect 4787 4422 4825 4428
rect 5167 4424 5204 4425
rect 4787 4404 4797 4422
rect 4815 4404 4825 4422
rect 4787 4395 4825 4404
rect 5165 4416 5205 4424
rect 5165 4398 5176 4416
rect 5194 4398 5205 4416
rect 6489 4414 6520 4435
rect 6910 4414 6946 4435
rect 6332 4413 6369 4414
rect 4787 4363 4821 4395
rect 3730 4331 4174 4337
rect 3730 4329 3898 4331
rect 3570 4258 3574 4263
rect 3531 4255 3574 4258
rect 3464 4241 3574 4255
rect 915 4212 951 4213
rect 763 4182 772 4202
rect 792 4182 800 4202
rect 651 4173 707 4175
rect 651 4172 688 4173
rect 763 4172 800 4182
rect 859 4202 1007 4212
rect 1107 4209 1203 4211
rect 859 4182 868 4202
rect 888 4182 978 4202
rect 998 4182 1007 4202
rect 859 4173 1007 4182
rect 1065 4202 1203 4209
rect 1065 4182 1074 4202
rect 1094 4182 1203 4202
rect 1065 4173 1203 4182
rect 859 4172 896 4173
rect 915 4121 951 4173
rect 970 4172 1007 4173
rect 1066 4172 1103 4173
rect 386 4119 427 4120
rect 278 4112 427 4119
rect 278 4092 396 4112
rect 416 4092 427 4112
rect 278 4084 427 4092
rect 494 4116 853 4120
rect 494 4111 816 4116
rect 494 4087 607 4111
rect 631 4092 816 4111
rect 840 4092 853 4116
rect 631 4087 853 4092
rect 494 4084 853 4087
rect 915 4084 950 4121
rect 1018 4118 1118 4121
rect 1018 4114 1085 4118
rect 1018 4088 1030 4114
rect 1056 4092 1085 4114
rect 1111 4092 1118 4118
rect 1056 4088 1118 4092
rect 1018 4084 1118 4088
rect 494 4063 525 4084
rect 915 4063 951 4084
rect 337 4062 374 4063
rect 336 4053 374 4062
rect 336 4033 345 4053
rect 365 4033 374 4053
rect 336 4025 374 4033
rect 440 4057 525 4063
rect 550 4062 587 4063
rect 440 4037 448 4057
rect 468 4037 525 4057
rect 440 4029 525 4037
rect 549 4053 587 4062
rect 549 4033 558 4053
rect 578 4033 587 4053
rect 440 4028 476 4029
rect 549 4025 587 4033
rect 653 4057 738 4063
rect 758 4062 795 4063
rect 653 4037 661 4057
rect 681 4056 738 4057
rect 681 4037 710 4056
rect 653 4036 710 4037
rect 731 4036 738 4056
rect 653 4029 738 4036
rect 757 4053 795 4062
rect 757 4033 766 4053
rect 786 4033 795 4053
rect 653 4028 689 4029
rect 757 4025 795 4033
rect 861 4057 1005 4063
rect 861 4037 869 4057
rect 889 4054 977 4057
rect 889 4037 920 4054
rect 861 4034 920 4037
rect 943 4037 977 4054
rect 997 4037 1005 4057
rect 943 4034 1005 4037
rect 861 4029 1005 4034
rect 861 4028 897 4029
rect 969 4028 1005 4029
rect 1071 4062 1108 4063
rect 1071 4061 1109 4062
rect 1071 4053 1135 4061
rect 1071 4033 1080 4053
rect 1100 4039 1135 4053
rect 1155 4039 1158 4059
rect 1100 4034 1158 4039
rect 1100 4033 1135 4034
rect 337 3996 374 4025
rect 338 3994 374 3996
rect 550 3994 587 4025
rect 338 3972 587 3994
rect 758 3993 795 4025
rect 1071 4021 1135 4033
rect 1175 3995 1202 4173
rect 3730 4151 3757 4329
rect 3797 4291 3861 4303
rect 4137 4299 4174 4331
rect 4345 4330 4594 4352
rect 4635 4331 4821 4363
rect 4649 4330 4821 4331
rect 4345 4299 4382 4330
rect 4558 4328 4594 4330
rect 4558 4299 4595 4328
rect 4787 4302 4821 4330
rect 5165 4350 5205 4398
rect 6331 4404 6369 4413
rect 6331 4384 6340 4404
rect 6360 4384 6369 4404
rect 6331 4376 6369 4384
rect 6435 4408 6520 4414
rect 6545 4413 6582 4414
rect 6435 4388 6443 4408
rect 6463 4388 6520 4408
rect 6435 4380 6520 4388
rect 6544 4404 6582 4413
rect 6544 4384 6553 4404
rect 6573 4384 6582 4404
rect 6435 4379 6471 4380
rect 6544 4376 6582 4384
rect 6648 4408 6733 4414
rect 6753 4413 6790 4414
rect 6648 4388 6656 4408
rect 6676 4407 6733 4408
rect 6676 4388 6705 4407
rect 6648 4387 6705 4388
rect 6726 4387 6733 4407
rect 6648 4380 6733 4387
rect 6752 4404 6790 4413
rect 6752 4384 6761 4404
rect 6781 4384 6790 4404
rect 6648 4379 6684 4380
rect 6752 4376 6790 4384
rect 6856 4408 7000 4414
rect 6856 4388 6864 4408
rect 6884 4391 6920 4408
rect 6940 4391 6972 4408
rect 6884 4388 6972 4391
rect 6992 4388 7000 4408
rect 6856 4380 7000 4388
rect 6856 4379 6892 4380
rect 6964 4379 7000 4380
rect 7066 4413 7103 4414
rect 7066 4412 7104 4413
rect 7066 4404 7130 4412
rect 7066 4384 7075 4404
rect 7095 4390 7130 4404
rect 7150 4390 7153 4410
rect 7095 4385 7153 4390
rect 7095 4384 7130 4385
rect 5476 4354 5586 4368
rect 5476 4351 5519 4354
rect 5165 4343 5290 4350
rect 5476 4346 5480 4351
rect 5165 4324 5257 4343
rect 5282 4324 5290 4343
rect 5165 4314 5290 4324
rect 5398 4324 5480 4346
rect 5509 4324 5519 4351
rect 5547 4327 5554 4354
rect 5583 4346 5586 4354
rect 6332 4347 6369 4376
rect 5583 4327 5648 4346
rect 6333 4345 6369 4347
rect 6545 4345 6582 4376
rect 6753 4349 6790 4376
rect 7066 4372 7130 4384
rect 5547 4324 5648 4327
rect 5398 4322 5648 4324
rect 3797 4290 3832 4291
rect 3774 4285 3832 4290
rect 3774 4265 3777 4285
rect 3797 4271 3832 4285
rect 3852 4271 3861 4291
rect 3797 4263 3861 4271
rect 3823 4262 3861 4263
rect 3824 4261 3861 4262
rect 3927 4295 3963 4296
rect 4035 4295 4071 4296
rect 3927 4288 4071 4295
rect 3927 4287 3987 4288
rect 3927 4267 3935 4287
rect 3955 4268 3987 4287
rect 4012 4287 4071 4288
rect 4012 4268 4043 4287
rect 3955 4267 4043 4268
rect 4063 4267 4071 4287
rect 3927 4261 4071 4267
rect 4137 4291 4175 4299
rect 4243 4295 4279 4296
rect 4137 4271 4146 4291
rect 4166 4271 4175 4291
rect 4137 4262 4175 4271
rect 4194 4288 4279 4295
rect 4194 4268 4201 4288
rect 4222 4287 4279 4288
rect 4222 4268 4251 4287
rect 4194 4267 4251 4268
rect 4271 4267 4279 4287
rect 4137 4261 4174 4262
rect 4194 4261 4279 4267
rect 4345 4291 4383 4299
rect 4456 4295 4492 4296
rect 4345 4271 4354 4291
rect 4374 4271 4383 4291
rect 4345 4262 4383 4271
rect 4407 4287 4492 4295
rect 4407 4267 4464 4287
rect 4484 4267 4492 4287
rect 4345 4261 4382 4262
rect 4407 4261 4492 4267
rect 4558 4291 4596 4299
rect 4558 4271 4567 4291
rect 4587 4271 4596 4291
rect 4558 4262 4596 4271
rect 4785 4292 4822 4302
rect 5165 4294 5205 4314
rect 4785 4274 4795 4292
rect 4813 4274 4822 4292
rect 4785 4265 4822 4274
rect 5164 4285 5205 4294
rect 5164 4267 5174 4285
rect 5192 4267 5205 4285
rect 4787 4264 4821 4265
rect 4558 4261 4595 4262
rect 3981 4240 4017 4261
rect 4407 4240 4438 4261
rect 5164 4258 5205 4267
rect 5164 4257 5201 4258
rect 5398 4243 5435 4322
rect 5476 4309 5586 4322
rect 5550 4253 5581 4254
rect 3814 4236 3914 4240
rect 3814 4232 3876 4236
rect 3814 4206 3821 4232
rect 3847 4210 3876 4232
rect 3902 4210 3914 4236
rect 3847 4206 3914 4210
rect 3814 4203 3914 4206
rect 3982 4203 4017 4240
rect 4079 4237 4438 4240
rect 4079 4232 4301 4237
rect 4079 4208 4092 4232
rect 4116 4213 4301 4232
rect 4325 4213 4438 4237
rect 4116 4208 4438 4213
rect 4079 4204 4438 4208
rect 4505 4232 4654 4240
rect 4505 4212 4516 4232
rect 4536 4212 4654 4232
rect 5398 4223 5407 4243
rect 5427 4223 5435 4243
rect 5398 4213 5435 4223
rect 5494 4243 5581 4253
rect 5494 4223 5503 4243
rect 5523 4223 5581 4243
rect 5494 4214 5581 4223
rect 5494 4213 5531 4214
rect 4505 4205 4654 4212
rect 4505 4204 4546 4205
rect 3829 4151 3866 4152
rect 3925 4151 3962 4152
rect 3981 4151 4017 4203
rect 4036 4151 4073 4152
rect 3729 4142 3867 4151
rect 3324 4121 3435 4136
rect 3324 4119 3366 4121
rect 2994 4098 3099 4100
rect 2650 4090 2820 4091
rect 2994 4090 3043 4098
rect 2650 4071 3043 4090
rect 3074 4071 3099 4098
rect 3324 4099 3331 4119
rect 3350 4099 3366 4119
rect 3324 4091 3366 4099
rect 3394 4119 3435 4121
rect 3394 4099 3408 4119
rect 3427 4099 3435 4119
rect 3729 4122 3838 4142
rect 3858 4122 3867 4142
rect 3729 4115 3867 4122
rect 3925 4142 4073 4151
rect 3925 4122 3934 4142
rect 3954 4122 4044 4142
rect 4064 4122 4073 4142
rect 3729 4113 3825 4115
rect 3925 4112 4073 4122
rect 4132 4142 4169 4152
rect 4244 4151 4281 4152
rect 4225 4149 4281 4151
rect 4132 4122 4140 4142
rect 4160 4122 4169 4142
rect 3981 4111 4017 4112
rect 3394 4091 3435 4099
rect 3324 4085 3435 4091
rect 2650 4064 3099 4071
rect 2650 4062 2820 4064
rect 1500 4031 1610 4045
rect 1500 4028 1543 4031
rect 1500 4023 1504 4028
rect 1034 3993 1202 3995
rect 758 3990 1202 3993
rect 419 3966 530 3972
rect 419 3958 460 3966
rect 108 3903 147 3947
rect 419 3938 427 3958
rect 446 3938 460 3958
rect 419 3936 460 3938
rect 488 3958 530 3966
rect 488 3938 504 3958
rect 523 3938 530 3958
rect 488 3936 530 3938
rect 419 3921 530 3936
rect 756 3967 1202 3990
rect 108 3879 148 3903
rect 448 3879 495 3881
rect 756 3879 794 3967
rect 1034 3966 1202 3967
rect 1422 4001 1504 4023
rect 1533 4001 1543 4028
rect 1571 4004 1578 4031
rect 1607 4023 1610 4031
rect 1607 4004 1672 4023
rect 1571 4001 1672 4004
rect 1422 3999 1672 4001
rect 1422 3920 1459 3999
rect 1500 3986 1610 3999
rect 1574 3930 1605 3931
rect 1422 3900 1431 3920
rect 1451 3900 1459 3920
rect 1422 3890 1459 3900
rect 1518 3920 1605 3930
rect 1518 3900 1527 3920
rect 1547 3900 1605 3920
rect 1518 3891 1605 3900
rect 1518 3890 1555 3891
rect 108 3846 794 3879
rect 108 3789 147 3846
rect 756 3844 794 3846
rect 1574 3838 1605 3891
rect 1635 3920 1672 3999
rect 1843 4012 2236 4016
rect 1843 3995 1862 4012
rect 1882 3996 2236 4012
rect 2256 3996 2259 4016
rect 1882 3995 2259 3996
rect 1843 3991 2259 3995
rect 1843 3990 2184 3991
rect 1787 3930 1818 3931
rect 1635 3900 1644 3920
rect 1664 3900 1672 3920
rect 1635 3890 1672 3900
rect 1731 3923 1818 3930
rect 1731 3920 1792 3923
rect 1731 3900 1740 3920
rect 1760 3903 1792 3920
rect 1813 3903 1818 3923
rect 1760 3900 1818 3903
rect 1731 3893 1818 3900
rect 1843 3920 1880 3990
rect 2146 3989 2183 3990
rect 1995 3930 2031 3931
rect 1843 3900 1852 3920
rect 1872 3900 1880 3920
rect 1731 3891 1787 3893
rect 1731 3890 1768 3891
rect 1843 3890 1880 3900
rect 1939 3920 2087 3930
rect 2187 3927 2283 3929
rect 1939 3900 1948 3920
rect 1968 3900 2058 3920
rect 2078 3900 2087 3920
rect 1939 3891 2087 3900
rect 2145 3920 2283 3927
rect 2145 3900 2154 3920
rect 2174 3900 2283 3920
rect 2145 3891 2283 3900
rect 1939 3890 1976 3891
rect 1995 3839 2031 3891
rect 2050 3890 2087 3891
rect 2146 3890 2183 3891
rect 1466 3837 1507 3838
rect 1358 3830 1507 3837
rect 1358 3810 1476 3830
rect 1496 3810 1507 3830
rect 1358 3802 1507 3810
rect 1574 3834 1933 3838
rect 1574 3829 1896 3834
rect 1574 3805 1687 3829
rect 1711 3810 1896 3829
rect 1920 3810 1933 3834
rect 1711 3805 1933 3810
rect 1574 3802 1933 3805
rect 1995 3802 2030 3839
rect 2098 3836 2198 3839
rect 2098 3832 2165 3836
rect 2098 3806 2110 3832
rect 2136 3810 2165 3832
rect 2191 3810 2198 3836
rect 2136 3806 2198 3810
rect 2098 3802 2198 3806
rect 108 3787 156 3789
rect 108 3769 119 3787
rect 137 3769 156 3787
rect 1574 3781 1605 3802
rect 1995 3781 2031 3802
rect 1417 3780 1454 3781
rect 108 3760 156 3769
rect 109 3759 156 3760
rect 422 3764 532 3778
rect 422 3761 465 3764
rect 422 3756 426 3761
rect 344 3734 426 3756
rect 455 3734 465 3761
rect 493 3737 500 3764
rect 529 3756 532 3764
rect 1416 3771 1454 3780
rect 529 3737 594 3756
rect 1416 3751 1425 3771
rect 1445 3751 1454 3771
rect 493 3734 594 3737
rect 344 3732 594 3734
rect 112 3696 149 3697
rect 108 3693 149 3696
rect 108 3688 150 3693
rect 108 3670 121 3688
rect 139 3670 150 3688
rect 108 3656 150 3670
rect 188 3656 235 3660
rect 108 3650 235 3656
rect 108 3621 196 3650
rect 225 3621 235 3650
rect 344 3653 381 3732
rect 422 3719 532 3732
rect 496 3663 527 3664
rect 344 3633 353 3653
rect 373 3633 381 3653
rect 344 3623 381 3633
rect 440 3653 527 3663
rect 440 3633 449 3653
rect 469 3633 527 3653
rect 440 3624 527 3633
rect 440 3623 477 3624
rect 108 3617 235 3621
rect 108 3600 147 3617
rect 188 3616 235 3617
rect 108 3582 119 3600
rect 137 3582 147 3600
rect 108 3573 147 3582
rect 109 3572 146 3573
rect 496 3571 527 3624
rect 557 3653 594 3732
rect 765 3729 1158 3749
rect 1178 3729 1181 3749
rect 1416 3743 1454 3751
rect 1520 3775 1605 3781
rect 1630 3780 1667 3781
rect 1520 3755 1528 3775
rect 1548 3755 1605 3775
rect 1520 3747 1605 3755
rect 1629 3771 1667 3780
rect 1629 3751 1638 3771
rect 1658 3751 1667 3771
rect 1520 3746 1556 3747
rect 1629 3743 1667 3751
rect 1733 3775 1818 3781
rect 1838 3780 1875 3781
rect 1733 3755 1741 3775
rect 1761 3774 1818 3775
rect 1761 3755 1790 3774
rect 1733 3754 1790 3755
rect 1811 3754 1818 3774
rect 1733 3747 1818 3754
rect 1837 3771 1875 3780
rect 1837 3751 1846 3771
rect 1866 3751 1875 3771
rect 1733 3746 1769 3747
rect 1837 3743 1875 3751
rect 1941 3775 2085 3781
rect 1941 3755 1949 3775
rect 1969 3773 2057 3775
rect 1969 3755 1998 3773
rect 1941 3752 1998 3755
rect 2025 3755 2057 3773
rect 2077 3755 2085 3775
rect 2025 3752 2085 3755
rect 1941 3747 2085 3752
rect 1941 3746 1977 3747
rect 2049 3746 2085 3747
rect 2151 3780 2188 3781
rect 2151 3779 2189 3780
rect 2151 3771 2215 3779
rect 2151 3751 2160 3771
rect 2180 3757 2215 3771
rect 2235 3757 2238 3777
rect 2180 3752 2238 3757
rect 2180 3751 2215 3752
rect 765 3724 1181 3729
rect 765 3723 1106 3724
rect 709 3663 740 3664
rect 557 3633 566 3653
rect 586 3633 594 3653
rect 557 3623 594 3633
rect 653 3656 740 3663
rect 653 3653 714 3656
rect 653 3633 662 3653
rect 682 3636 714 3653
rect 735 3636 740 3656
rect 682 3633 740 3636
rect 653 3626 740 3633
rect 765 3653 802 3723
rect 1068 3722 1105 3723
rect 1417 3714 1454 3743
rect 1418 3712 1454 3714
rect 1630 3712 1667 3743
rect 1418 3690 1667 3712
rect 1838 3711 1875 3743
rect 2151 3739 2215 3751
rect 2255 3713 2282 3891
rect 2650 3884 2679 4062
rect 2719 4024 2783 4036
rect 3059 4032 3096 4064
rect 3267 4063 3516 4085
rect 3267 4032 3304 4063
rect 3480 4061 3516 4063
rect 3480 4032 3517 4061
rect 3829 4052 3866 4053
rect 4132 4052 4169 4122
rect 4194 4142 4281 4149
rect 4194 4139 4252 4142
rect 4194 4119 4199 4139
rect 4220 4122 4252 4139
rect 4272 4122 4281 4142
rect 4220 4119 4281 4122
rect 4194 4112 4281 4119
rect 4340 4142 4377 4152
rect 4340 4122 4348 4142
rect 4368 4122 4377 4142
rect 4194 4111 4225 4112
rect 3828 4051 4169 4052
rect 3753 4046 4169 4051
rect 2719 4023 2754 4024
rect 2696 4018 2754 4023
rect 2696 3998 2699 4018
rect 2719 4004 2754 4018
rect 2774 4004 2783 4024
rect 2719 3996 2783 4004
rect 2745 3995 2783 3996
rect 2746 3994 2783 3995
rect 2849 4028 2885 4029
rect 2957 4028 2993 4029
rect 2849 4020 2993 4028
rect 2849 4000 2857 4020
rect 2877 4000 2965 4020
rect 2985 4000 2993 4020
rect 2849 3994 2993 4000
rect 3059 4024 3097 4032
rect 3165 4028 3201 4029
rect 3059 4004 3068 4024
rect 3088 4004 3097 4024
rect 3059 3995 3097 4004
rect 3116 4021 3201 4028
rect 3116 4001 3123 4021
rect 3144 4020 3201 4021
rect 3144 4001 3173 4020
rect 3116 4000 3173 4001
rect 3193 4000 3201 4020
rect 3059 3994 3096 3995
rect 3116 3994 3201 4000
rect 3267 4024 3305 4032
rect 3378 4028 3414 4029
rect 3267 4004 3276 4024
rect 3296 4004 3305 4024
rect 3267 3995 3305 4004
rect 3329 4020 3414 4028
rect 3329 4000 3386 4020
rect 3406 4000 3414 4020
rect 3267 3994 3304 3995
rect 3329 3994 3414 4000
rect 3480 4024 3518 4032
rect 3753 4026 3756 4046
rect 3776 4026 4169 4046
rect 4340 4043 4377 4122
rect 4407 4151 4438 4204
rect 4788 4202 4825 4203
rect 4787 4193 4826 4202
rect 4787 4175 4797 4193
rect 4815 4175 4826 4193
rect 5167 4191 5204 4195
rect 4699 4158 4746 4159
rect 4787 4158 4826 4175
rect 4699 4154 4826 4158
rect 4457 4151 4494 4152
rect 4407 4142 4494 4151
rect 4407 4122 4465 4142
rect 4485 4122 4494 4142
rect 4407 4112 4494 4122
rect 4553 4142 4590 4152
rect 4553 4122 4561 4142
rect 4581 4122 4590 4142
rect 4407 4111 4438 4112
rect 4402 4043 4512 4056
rect 4553 4043 4590 4122
rect 4699 4125 4709 4154
rect 4738 4125 4826 4154
rect 4699 4119 4826 4125
rect 4699 4115 4746 4119
rect 4784 4105 4826 4119
rect 4784 4087 4795 4105
rect 4813 4087 4826 4105
rect 4784 4082 4826 4087
rect 4785 4079 4826 4082
rect 5164 4186 5204 4191
rect 5164 4168 5176 4186
rect 5194 4168 5204 4186
rect 4785 4078 4822 4079
rect 4340 4041 4590 4043
rect 4340 4038 4441 4041
rect 3480 4004 3489 4024
rect 3509 4004 3518 4024
rect 4340 4019 4405 4038
rect 3480 3995 3518 4004
rect 4402 4011 4405 4019
rect 4434 4011 4441 4038
rect 4469 4014 4479 4041
rect 4508 4019 4590 4041
rect 4508 4014 4512 4019
rect 4469 4011 4512 4014
rect 4402 3997 4512 4011
rect 4778 4015 4825 4016
rect 4778 4006 4826 4015
rect 3480 3994 3517 3995
rect 2903 3973 2939 3994
rect 3329 3973 3360 3994
rect 4778 3988 4797 4006
rect 4815 3988 4826 4006
rect 4778 3986 4826 3988
rect 2736 3969 2836 3973
rect 2736 3965 2798 3969
rect 2736 3939 2743 3965
rect 2769 3943 2798 3965
rect 2824 3943 2836 3969
rect 2769 3939 2836 3943
rect 2736 3936 2836 3939
rect 2904 3936 2939 3973
rect 3001 3970 3360 3973
rect 3001 3965 3223 3970
rect 3001 3941 3014 3965
rect 3038 3946 3223 3965
rect 3247 3946 3360 3970
rect 3038 3941 3360 3946
rect 3001 3937 3360 3941
rect 3427 3965 3576 3973
rect 3427 3945 3438 3965
rect 3458 3945 3576 3965
rect 3427 3938 3576 3945
rect 3427 3937 3468 3938
rect 2903 3897 2939 3936
rect 2751 3884 2788 3885
rect 2847 3884 2884 3885
rect 2903 3884 2910 3897
rect 2650 3875 2789 3884
rect 2650 3855 2760 3875
rect 2780 3855 2789 3875
rect 2650 3848 2789 3855
rect 2847 3875 2910 3884
rect 2847 3855 2856 3875
rect 2876 3859 2910 3875
rect 2933 3884 2939 3897
rect 2958 3884 2995 3885
rect 2933 3875 2995 3884
rect 2933 3859 2966 3875
rect 2876 3855 2966 3859
rect 2986 3855 2995 3875
rect 2650 3846 2747 3848
rect 2650 3845 2679 3846
rect 2847 3845 2995 3855
rect 3054 3875 3091 3885
rect 3166 3884 3203 3885
rect 3147 3882 3203 3884
rect 3054 3855 3062 3875
rect 3082 3855 3091 3875
rect 2903 3844 2939 3845
rect 2751 3785 2788 3786
rect 3054 3785 3091 3855
rect 3116 3875 3203 3882
rect 3116 3872 3174 3875
rect 3116 3852 3121 3872
rect 3142 3855 3174 3872
rect 3194 3855 3203 3875
rect 3142 3852 3203 3855
rect 3116 3845 3203 3852
rect 3262 3875 3299 3885
rect 3262 3855 3270 3875
rect 3290 3855 3299 3875
rect 3116 3844 3147 3845
rect 2750 3784 3091 3785
rect 2675 3780 3091 3784
rect 2675 3779 3052 3780
rect 2675 3759 2678 3779
rect 2698 3763 3052 3779
rect 3072 3763 3091 3780
rect 2698 3759 3091 3763
rect 3262 3776 3299 3855
rect 3329 3884 3360 3937
rect 4140 3929 4178 3931
rect 4787 3929 4826 3986
rect 4140 3896 4826 3929
rect 3379 3884 3416 3885
rect 3329 3875 3416 3884
rect 3329 3855 3387 3875
rect 3407 3855 3416 3875
rect 3329 3845 3416 3855
rect 3475 3875 3512 3885
rect 3475 3855 3483 3875
rect 3503 3855 3512 3875
rect 3329 3844 3360 3845
rect 3324 3776 3434 3789
rect 3475 3776 3512 3855
rect 3262 3774 3512 3776
rect 3262 3771 3363 3774
rect 3262 3752 3327 3771
rect 3324 3744 3327 3752
rect 3356 3744 3363 3771
rect 3391 3747 3401 3774
rect 3430 3752 3512 3774
rect 3732 3808 3900 3809
rect 4140 3808 4178 3896
rect 4439 3894 4486 3896
rect 4786 3872 4826 3896
rect 3732 3785 4178 3808
rect 4404 3839 4515 3854
rect 4404 3837 4446 3839
rect 4404 3817 4411 3837
rect 4430 3817 4446 3837
rect 4404 3809 4446 3817
rect 4474 3837 4515 3839
rect 4474 3817 4488 3837
rect 4507 3817 4515 3837
rect 4787 3828 4826 3872
rect 4474 3809 4515 3817
rect 4404 3803 4515 3809
rect 3732 3782 4176 3785
rect 3732 3780 3900 3782
rect 3430 3747 3434 3752
rect 3391 3744 3434 3747
rect 3324 3730 3434 3744
rect 2114 3711 2282 3713
rect 1835 3704 2282 3711
rect 1499 3684 1610 3690
rect 1499 3676 1540 3684
rect 917 3663 953 3664
rect 765 3633 774 3653
rect 794 3633 802 3653
rect 653 3624 709 3626
rect 653 3623 690 3624
rect 765 3623 802 3633
rect 861 3653 1009 3663
rect 1109 3660 1205 3662
rect 861 3633 870 3653
rect 890 3633 980 3653
rect 1000 3633 1009 3653
rect 861 3624 1009 3633
rect 1067 3653 1205 3660
rect 1067 3633 1076 3653
rect 1096 3633 1205 3653
rect 1499 3656 1507 3676
rect 1526 3656 1540 3676
rect 1499 3654 1540 3656
rect 1568 3676 1610 3684
rect 1568 3656 1584 3676
rect 1603 3656 1610 3676
rect 1835 3677 1860 3704
rect 1891 3685 2282 3704
rect 1891 3677 1940 3685
rect 2114 3684 2282 3685
rect 1835 3675 1940 3677
rect 1568 3654 1610 3656
rect 1499 3639 1610 3654
rect 1067 3624 1205 3633
rect 861 3623 898 3624
rect 917 3572 953 3624
rect 972 3623 1009 3624
rect 1068 3623 1105 3624
rect 388 3570 429 3571
rect 280 3563 429 3570
rect 280 3543 398 3563
rect 418 3543 429 3563
rect 280 3535 429 3543
rect 496 3567 855 3571
rect 496 3562 818 3567
rect 496 3538 609 3562
rect 633 3543 818 3562
rect 842 3543 855 3567
rect 633 3538 855 3543
rect 496 3535 855 3538
rect 917 3535 952 3572
rect 1020 3569 1120 3572
rect 1020 3565 1087 3569
rect 1020 3539 1032 3565
rect 1058 3543 1087 3565
rect 1113 3543 1120 3569
rect 1058 3539 1120 3543
rect 1020 3535 1120 3539
rect 496 3514 527 3535
rect 917 3514 953 3535
rect 339 3513 376 3514
rect 113 3510 147 3511
rect 112 3501 149 3510
rect 112 3483 121 3501
rect 139 3483 149 3501
rect 112 3473 149 3483
rect 338 3504 376 3513
rect 338 3484 347 3504
rect 367 3484 376 3504
rect 338 3476 376 3484
rect 442 3508 527 3514
rect 552 3513 589 3514
rect 442 3488 450 3508
rect 470 3488 527 3508
rect 442 3480 527 3488
rect 551 3504 589 3513
rect 551 3484 560 3504
rect 580 3484 589 3504
rect 442 3479 478 3480
rect 551 3476 589 3484
rect 655 3508 740 3514
rect 760 3513 797 3514
rect 655 3488 663 3508
rect 683 3507 740 3508
rect 683 3488 712 3507
rect 655 3487 712 3488
rect 733 3487 740 3507
rect 655 3480 740 3487
rect 759 3504 797 3513
rect 759 3484 768 3504
rect 788 3484 797 3504
rect 655 3479 691 3480
rect 759 3476 797 3484
rect 863 3508 1007 3514
rect 863 3488 871 3508
rect 891 3507 979 3508
rect 891 3488 922 3507
rect 863 3487 922 3488
rect 947 3488 979 3507
rect 999 3488 1007 3508
rect 947 3487 1007 3488
rect 863 3480 1007 3487
rect 863 3479 899 3480
rect 971 3479 1007 3480
rect 1073 3513 1110 3514
rect 1073 3512 1111 3513
rect 1073 3504 1137 3512
rect 1073 3484 1082 3504
rect 1102 3490 1137 3504
rect 1157 3490 1160 3510
rect 1102 3485 1160 3490
rect 1102 3484 1137 3485
rect 113 3445 147 3473
rect 339 3447 376 3476
rect 340 3445 376 3447
rect 552 3445 589 3476
rect 113 3444 285 3445
rect 113 3412 299 3444
rect 340 3423 589 3445
rect 760 3444 797 3476
rect 1073 3472 1137 3484
rect 1177 3446 1204 3624
rect 3732 3602 3759 3780
rect 3799 3742 3863 3754
rect 4139 3750 4176 3782
rect 4347 3781 4596 3803
rect 4347 3750 4384 3781
rect 4560 3779 4596 3781
rect 4560 3750 4597 3779
rect 3799 3741 3834 3742
rect 3776 3736 3834 3741
rect 3776 3716 3779 3736
rect 3799 3722 3834 3736
rect 3854 3722 3863 3742
rect 3799 3714 3863 3722
rect 3825 3713 3863 3714
rect 3826 3712 3863 3713
rect 3929 3746 3965 3747
rect 4037 3746 4073 3747
rect 3929 3741 4073 3746
rect 3929 3738 3991 3741
rect 3929 3718 3937 3738
rect 3957 3721 3991 3738
rect 4014 3738 4073 3741
rect 4014 3721 4045 3738
rect 3957 3718 4045 3721
rect 4065 3718 4073 3738
rect 3929 3712 4073 3718
rect 4139 3742 4177 3750
rect 4245 3746 4281 3747
rect 4139 3722 4148 3742
rect 4168 3722 4177 3742
rect 4139 3713 4177 3722
rect 4196 3739 4281 3746
rect 4196 3719 4203 3739
rect 4224 3738 4281 3739
rect 4224 3719 4253 3738
rect 4196 3718 4253 3719
rect 4273 3718 4281 3738
rect 4139 3712 4176 3713
rect 4196 3712 4281 3718
rect 4347 3742 4385 3750
rect 4458 3746 4494 3747
rect 4347 3722 4356 3742
rect 4376 3722 4385 3742
rect 4347 3713 4385 3722
rect 4409 3738 4494 3746
rect 4409 3718 4466 3738
rect 4486 3718 4494 3738
rect 4347 3712 4384 3713
rect 4409 3712 4494 3718
rect 4560 3742 4598 3750
rect 4560 3722 4569 3742
rect 4589 3722 4598 3742
rect 4560 3713 4598 3722
rect 4560 3712 4597 3713
rect 3983 3691 4019 3712
rect 4409 3691 4440 3712
rect 3816 3687 3916 3691
rect 3816 3683 3878 3687
rect 3816 3657 3823 3683
rect 3849 3661 3878 3683
rect 3904 3661 3916 3687
rect 3849 3657 3916 3661
rect 3816 3654 3916 3657
rect 3984 3654 4019 3691
rect 4081 3688 4440 3691
rect 4081 3683 4303 3688
rect 4081 3659 4094 3683
rect 4118 3664 4303 3683
rect 4327 3664 4440 3688
rect 4118 3659 4440 3664
rect 4081 3655 4440 3659
rect 4507 3683 4656 3691
rect 4507 3663 4518 3683
rect 4538 3663 4656 3683
rect 4507 3656 4656 3663
rect 4507 3655 4548 3656
rect 3831 3602 3868 3603
rect 3927 3602 3964 3603
rect 3983 3602 4019 3654
rect 4038 3602 4075 3603
rect 3731 3593 3869 3602
rect 3731 3573 3840 3593
rect 3860 3573 3869 3593
rect 3731 3566 3869 3573
rect 3927 3593 4075 3602
rect 3927 3573 3936 3593
rect 3956 3573 4046 3593
rect 4066 3573 4075 3593
rect 3731 3564 3827 3566
rect 3927 3563 4075 3573
rect 4134 3593 4171 3603
rect 4246 3602 4283 3603
rect 4227 3600 4283 3602
rect 4134 3573 4142 3593
rect 4162 3573 4171 3593
rect 3983 3562 4019 3563
rect 1360 3520 1470 3534
rect 1360 3517 1403 3520
rect 1360 3512 1364 3517
rect 1036 3444 1204 3446
rect 760 3438 1204 3444
rect 113 3380 147 3412
rect 109 3371 147 3380
rect 109 3353 119 3371
rect 137 3353 147 3371
rect 109 3347 147 3353
rect 265 3349 299 3412
rect 421 3417 532 3423
rect 421 3409 462 3417
rect 421 3389 429 3409
rect 448 3389 462 3409
rect 421 3387 462 3389
rect 490 3409 532 3417
rect 490 3389 506 3409
rect 525 3389 532 3409
rect 490 3387 532 3389
rect 421 3372 532 3387
rect 759 3418 1204 3438
rect 759 3349 797 3418
rect 1036 3417 1204 3418
rect 1282 3490 1364 3512
rect 1393 3490 1403 3517
rect 1431 3493 1438 3520
rect 1467 3512 1470 3520
rect 3465 3529 3576 3544
rect 3465 3527 3507 3529
rect 1467 3493 1532 3512
rect 1431 3490 1532 3493
rect 1282 3488 1532 3490
rect 1282 3409 1319 3488
rect 1360 3475 1470 3488
rect 1434 3419 1465 3420
rect 1282 3389 1291 3409
rect 1311 3389 1319 3409
rect 1282 3379 1319 3389
rect 1378 3409 1465 3419
rect 1378 3389 1387 3409
rect 1407 3389 1465 3409
rect 1378 3380 1465 3389
rect 1378 3379 1415 3380
rect 109 3343 146 3347
rect 265 3338 797 3349
rect 264 3322 797 3338
rect 1434 3327 1465 3380
rect 1495 3409 1532 3488
rect 1703 3498 2096 3505
rect 1703 3481 1711 3498
rect 1743 3485 2096 3498
rect 2116 3485 2119 3505
rect 3198 3500 3239 3509
rect 1743 3481 2119 3485
rect 1703 3480 2119 3481
rect 2793 3498 2961 3499
rect 3198 3498 3207 3500
rect 1703 3479 2044 3480
rect 1647 3419 1678 3420
rect 1495 3389 1504 3409
rect 1524 3389 1532 3409
rect 1495 3379 1532 3389
rect 1591 3412 1678 3419
rect 1591 3409 1652 3412
rect 1591 3389 1600 3409
rect 1620 3392 1652 3409
rect 1673 3392 1678 3412
rect 1620 3389 1678 3392
rect 1591 3382 1678 3389
rect 1703 3409 1740 3479
rect 2006 3478 2043 3479
rect 2793 3478 3207 3498
rect 3233 3478 3239 3500
rect 3465 3507 3472 3527
rect 3491 3507 3507 3527
rect 3465 3499 3507 3507
rect 3535 3527 3576 3529
rect 3535 3507 3549 3527
rect 3568 3507 3576 3527
rect 3535 3499 3576 3507
rect 3831 3503 3868 3504
rect 4134 3503 4171 3573
rect 4196 3593 4283 3600
rect 4196 3590 4254 3593
rect 4196 3570 4201 3590
rect 4222 3573 4254 3590
rect 4274 3573 4283 3593
rect 4222 3570 4283 3573
rect 4196 3563 4283 3570
rect 4342 3593 4379 3603
rect 4342 3573 4350 3593
rect 4370 3573 4379 3593
rect 4196 3562 4227 3563
rect 3830 3502 4171 3503
rect 3465 3493 3576 3499
rect 3755 3497 4171 3502
rect 2793 3472 3239 3478
rect 2793 3470 2961 3472
rect 1855 3419 1891 3420
rect 1703 3389 1712 3409
rect 1732 3389 1740 3409
rect 1591 3380 1647 3382
rect 1591 3379 1628 3380
rect 1703 3379 1740 3389
rect 1799 3409 1947 3419
rect 2047 3416 2143 3418
rect 1799 3389 1808 3409
rect 1828 3404 1918 3409
rect 1828 3389 1863 3404
rect 1799 3380 1863 3389
rect 1799 3379 1836 3380
rect 1855 3363 1863 3380
rect 1884 3389 1918 3404
rect 1938 3389 1947 3409
rect 1884 3380 1947 3389
rect 2005 3409 2143 3416
rect 2005 3389 2014 3409
rect 2034 3389 2143 3409
rect 2005 3380 2143 3389
rect 1884 3363 1891 3380
rect 1910 3379 1947 3380
rect 2006 3379 2043 3380
rect 1855 3328 1891 3363
rect 1326 3326 1367 3327
rect 264 3321 778 3322
rect 1218 3319 1367 3326
rect 1218 3299 1336 3319
rect 1356 3299 1367 3319
rect 1218 3291 1367 3299
rect 1434 3323 1793 3327
rect 1434 3318 1756 3323
rect 1434 3294 1547 3318
rect 1571 3299 1756 3318
rect 1780 3299 1793 3323
rect 1571 3294 1793 3299
rect 1434 3291 1793 3294
rect 1855 3291 1890 3328
rect 1958 3325 2058 3328
rect 1958 3321 2025 3325
rect 1958 3295 1970 3321
rect 1996 3299 2025 3321
rect 2051 3299 2058 3325
rect 1996 3295 2058 3299
rect 1958 3291 2058 3295
rect 112 3280 149 3281
rect 110 3272 150 3280
rect 110 3254 121 3272
rect 139 3254 150 3272
rect 1434 3270 1465 3291
rect 1855 3270 1891 3291
rect 1277 3269 1314 3270
rect 110 3206 150 3254
rect 1276 3260 1314 3269
rect 1276 3240 1285 3260
rect 1305 3240 1314 3260
rect 1276 3232 1314 3240
rect 1380 3264 1465 3270
rect 1490 3269 1527 3270
rect 1380 3244 1388 3264
rect 1408 3244 1465 3264
rect 1380 3236 1465 3244
rect 1489 3260 1527 3269
rect 1489 3240 1498 3260
rect 1518 3240 1527 3260
rect 1380 3235 1416 3236
rect 1489 3232 1527 3240
rect 1593 3264 1678 3270
rect 1698 3269 1735 3270
rect 1593 3244 1601 3264
rect 1621 3263 1678 3264
rect 1621 3244 1650 3263
rect 1593 3243 1650 3244
rect 1671 3243 1678 3263
rect 1593 3236 1678 3243
rect 1697 3260 1735 3269
rect 1697 3240 1706 3260
rect 1726 3240 1735 3260
rect 1593 3235 1629 3236
rect 1697 3232 1735 3240
rect 1801 3264 1945 3270
rect 1801 3244 1809 3264
rect 1829 3244 1917 3264
rect 1937 3244 1945 3264
rect 1801 3236 1945 3244
rect 1801 3235 1837 3236
rect 1909 3235 1945 3236
rect 2011 3269 2048 3270
rect 2011 3268 2049 3269
rect 2011 3260 2075 3268
rect 2011 3240 2020 3260
rect 2040 3246 2075 3260
rect 2095 3246 2098 3266
rect 2040 3241 2098 3246
rect 2040 3240 2075 3241
rect 421 3210 531 3224
rect 421 3207 464 3210
rect 110 3199 235 3206
rect 421 3202 425 3207
rect 110 3180 202 3199
rect 227 3180 235 3199
rect 110 3170 235 3180
rect 343 3180 425 3202
rect 454 3180 464 3207
rect 492 3183 499 3210
rect 528 3202 531 3210
rect 1277 3203 1314 3232
rect 528 3183 593 3202
rect 1278 3201 1314 3203
rect 1490 3201 1527 3232
rect 1698 3205 1735 3232
rect 2011 3228 2075 3240
rect 492 3180 593 3183
rect 343 3178 593 3180
rect 110 3150 150 3170
rect 109 3141 150 3150
rect 109 3123 119 3141
rect 137 3123 150 3141
rect 109 3114 150 3123
rect 109 3113 146 3114
rect 343 3099 380 3178
rect 421 3165 531 3178
rect 495 3109 526 3110
rect 343 3079 352 3099
rect 372 3079 380 3099
rect 343 3069 380 3079
rect 439 3099 526 3109
rect 439 3079 448 3099
rect 468 3079 526 3099
rect 439 3070 526 3079
rect 439 3069 476 3070
rect 112 3047 149 3051
rect 109 3042 149 3047
rect 109 3024 121 3042
rect 139 3024 149 3042
rect 109 2844 149 3024
rect 495 3017 526 3070
rect 556 3099 593 3178
rect 764 3175 1157 3195
rect 1177 3175 1180 3195
rect 1278 3179 1527 3201
rect 1696 3200 1737 3205
rect 2115 3202 2142 3380
rect 2793 3292 2820 3470
rect 3198 3467 3239 3472
rect 3408 3471 3657 3493
rect 3755 3477 3758 3497
rect 3778 3477 4171 3497
rect 4342 3494 4379 3573
rect 4409 3602 4440 3655
rect 4786 3648 4826 3828
rect 5164 3988 5204 4168
rect 5550 4161 5581 4214
rect 5611 4243 5648 4322
rect 5819 4319 6212 4339
rect 6232 4319 6235 4339
rect 6333 4323 6582 4345
rect 6751 4344 6792 4349
rect 7170 4346 7197 4524
rect 7848 4436 7875 4614
rect 8253 4611 8294 4616
rect 8463 4615 8712 4637
rect 8810 4621 8813 4641
rect 8833 4621 9226 4641
rect 9397 4638 9434 4717
rect 9464 4746 9495 4799
rect 9841 4792 9881 4972
rect 10135 4954 10825 4977
rect 11573 4965 11604 5018
rect 11634 5047 11671 5126
rect 11842 5123 12235 5143
rect 12255 5123 12258 5143
rect 12580 5142 12633 5150
rect 11842 5118 12258 5123
rect 11842 5117 12183 5118
rect 11786 5057 11817 5058
rect 11634 5027 11643 5047
rect 11663 5027 11671 5047
rect 11634 5017 11671 5027
rect 11730 5050 11817 5057
rect 11730 5047 11791 5050
rect 11730 5027 11739 5047
rect 11759 5030 11791 5047
rect 11812 5030 11817 5050
rect 11759 5027 11817 5030
rect 11730 5020 11817 5027
rect 11842 5047 11879 5117
rect 12145 5116 12182 5117
rect 11994 5057 12030 5058
rect 11842 5027 11851 5047
rect 11871 5027 11879 5047
rect 11730 5018 11786 5020
rect 11730 5017 11767 5018
rect 11842 5017 11879 5027
rect 11938 5047 12086 5057
rect 12186 5054 12282 5056
rect 11938 5027 11947 5047
rect 11967 5027 12057 5047
rect 12077 5027 12086 5047
rect 11938 5018 12086 5027
rect 12144 5047 12282 5054
rect 12144 5027 12153 5047
rect 12173 5027 12282 5047
rect 12144 5018 12282 5027
rect 11938 5017 11975 5018
rect 11994 4966 12030 5018
rect 12049 5017 12086 5018
rect 12145 5017 12182 5018
rect 11465 4964 11506 4965
rect 10135 4935 10177 4954
rect 10787 4952 10825 4954
rect 11357 4957 11506 4964
rect 10138 4897 10177 4935
rect 11357 4937 11475 4957
rect 11495 4937 11506 4957
rect 11357 4929 11506 4937
rect 11573 4961 11932 4965
rect 11573 4956 11895 4961
rect 11573 4932 11686 4956
rect 11710 4937 11895 4956
rect 11919 4937 11932 4961
rect 11710 4932 11932 4937
rect 11573 4929 11932 4932
rect 11994 4929 12029 4966
rect 12097 4963 12197 4966
rect 12097 4959 12164 4963
rect 12097 4933 12109 4959
rect 12135 4937 12164 4959
rect 12190 4937 12197 4963
rect 12135 4933 12197 4937
rect 12097 4929 12197 4933
rect 11573 4908 11604 4929
rect 11994 4908 12030 4929
rect 11416 4907 11453 4908
rect 11415 4898 11453 4907
rect 10138 4895 10186 4897
rect 10138 4877 10149 4895
rect 10167 4877 10186 4895
rect 10138 4868 10186 4877
rect 10139 4867 10186 4868
rect 10452 4872 10562 4886
rect 10452 4869 10495 4872
rect 10452 4864 10456 4869
rect 10374 4842 10456 4864
rect 10485 4842 10495 4869
rect 10523 4845 10530 4872
rect 10559 4864 10562 4872
rect 11415 4878 11424 4898
rect 11444 4878 11453 4898
rect 11415 4870 11453 4878
rect 11519 4902 11604 4908
rect 11629 4907 11666 4908
rect 11519 4882 11527 4902
rect 11547 4882 11604 4902
rect 11519 4874 11604 4882
rect 11628 4898 11666 4907
rect 11628 4878 11637 4898
rect 11657 4878 11666 4898
rect 11519 4873 11555 4874
rect 11628 4870 11666 4878
rect 11732 4902 11817 4908
rect 11837 4907 11874 4908
rect 11732 4882 11740 4902
rect 11760 4901 11817 4902
rect 11760 4882 11789 4901
rect 11732 4881 11789 4882
rect 11810 4881 11817 4901
rect 11732 4874 11817 4881
rect 11836 4898 11874 4907
rect 11836 4878 11845 4898
rect 11865 4878 11874 4898
rect 11732 4873 11768 4874
rect 11836 4870 11874 4878
rect 11940 4904 12084 4908
rect 11940 4902 11997 4904
rect 11940 4882 11948 4902
rect 11968 4882 11997 4902
rect 11940 4880 11997 4882
rect 12023 4902 12084 4904
rect 12023 4882 12056 4902
rect 12076 4882 12084 4902
rect 12023 4880 12084 4882
rect 11940 4874 12084 4880
rect 11940 4873 11976 4874
rect 12048 4873 12084 4874
rect 12150 4907 12187 4908
rect 12150 4906 12188 4907
rect 12150 4898 12214 4906
rect 12150 4878 12159 4898
rect 12179 4884 12214 4898
rect 12234 4884 12237 4904
rect 12179 4879 12237 4884
rect 12179 4878 12214 4879
rect 10559 4845 10624 4864
rect 10523 4842 10624 4845
rect 10374 4840 10624 4842
rect 10142 4804 10179 4805
rect 9841 4774 9851 4792
rect 9869 4774 9881 4792
rect 9841 4769 9881 4774
rect 10138 4801 10179 4804
rect 10138 4796 10180 4801
rect 10138 4778 10151 4796
rect 10169 4778 10180 4796
rect 9841 4765 9878 4769
rect 10138 4764 10180 4778
rect 10218 4764 10265 4768
rect 10138 4758 10265 4764
rect 9514 4746 9551 4747
rect 9464 4737 9551 4746
rect 9464 4717 9522 4737
rect 9542 4717 9551 4737
rect 9464 4707 9551 4717
rect 9610 4737 9647 4747
rect 9610 4717 9618 4737
rect 9638 4717 9647 4737
rect 9464 4706 9495 4707
rect 9459 4638 9569 4651
rect 9610 4638 9647 4717
rect 10138 4729 10226 4758
rect 10255 4729 10265 4758
rect 10374 4761 10411 4840
rect 10452 4827 10562 4840
rect 10526 4771 10557 4772
rect 10374 4741 10383 4761
rect 10403 4741 10411 4761
rect 10374 4731 10411 4741
rect 10470 4761 10557 4771
rect 10470 4741 10479 4761
rect 10499 4741 10557 4761
rect 10470 4732 10557 4741
rect 10470 4731 10507 4732
rect 10138 4725 10265 4729
rect 10138 4708 10177 4725
rect 10218 4724 10265 4725
rect 9844 4702 9881 4703
rect 9840 4693 9881 4702
rect 9840 4675 9853 4693
rect 9871 4675 9881 4693
rect 10138 4690 10149 4708
rect 10167 4690 10177 4708
rect 10138 4681 10177 4690
rect 10139 4680 10176 4681
rect 10526 4679 10557 4732
rect 10587 4761 10624 4840
rect 10795 4837 11188 4857
rect 11208 4837 11211 4857
rect 11416 4841 11453 4870
rect 10795 4832 11211 4837
rect 11417 4839 11453 4841
rect 11629 4839 11666 4870
rect 10795 4831 11136 4832
rect 10739 4771 10770 4772
rect 10587 4741 10596 4761
rect 10616 4741 10624 4761
rect 10587 4731 10624 4741
rect 10683 4764 10770 4771
rect 10683 4761 10744 4764
rect 10683 4741 10692 4761
rect 10712 4744 10744 4761
rect 10765 4744 10770 4764
rect 10712 4741 10770 4744
rect 10683 4734 10770 4741
rect 10795 4761 10832 4831
rect 11098 4830 11135 4831
rect 11417 4817 11666 4839
rect 11837 4838 11874 4870
rect 12150 4866 12214 4878
rect 12254 4841 12281 5018
rect 12714 4973 12741 5150
rect 12781 5113 12845 5125
rect 13121 5121 13158 5153
rect 13329 5152 13578 5174
rect 13860 5160 13897 5161
rect 14163 5160 14200 5230
rect 14225 5250 14312 5257
rect 14225 5247 14283 5250
rect 14225 5227 14230 5247
rect 14251 5230 14283 5247
rect 14303 5230 14312 5250
rect 14251 5227 14312 5230
rect 14225 5220 14312 5227
rect 14371 5250 14408 5260
rect 14371 5230 14379 5250
rect 14399 5230 14408 5250
rect 14225 5219 14256 5220
rect 13859 5159 14200 5160
rect 13329 5121 13366 5152
rect 13542 5150 13578 5152
rect 13784 5154 14200 5159
rect 13542 5121 13579 5150
rect 13784 5134 13787 5154
rect 13807 5134 14200 5154
rect 14371 5151 14408 5230
rect 14438 5259 14469 5312
rect 14819 5310 14856 5311
rect 14818 5301 14857 5310
rect 14818 5283 14828 5301
rect 14846 5283 14857 5301
rect 15198 5299 15235 5303
rect 14730 5266 14777 5267
rect 14818 5266 14857 5283
rect 14730 5262 14857 5266
rect 14488 5259 14525 5260
rect 14438 5250 14525 5259
rect 14438 5230 14496 5250
rect 14516 5230 14525 5250
rect 14438 5220 14525 5230
rect 14584 5250 14621 5260
rect 14584 5230 14592 5250
rect 14612 5230 14621 5250
rect 14438 5219 14469 5220
rect 14433 5151 14543 5164
rect 14584 5151 14621 5230
rect 14730 5233 14740 5262
rect 14769 5233 14857 5262
rect 14730 5227 14857 5233
rect 14730 5223 14777 5227
rect 14815 5213 14857 5227
rect 14815 5195 14826 5213
rect 14844 5195 14857 5213
rect 14815 5190 14857 5195
rect 14816 5187 14857 5190
rect 15195 5294 15235 5299
rect 15195 5276 15207 5294
rect 15225 5276 15235 5294
rect 14816 5186 14853 5187
rect 14371 5149 14621 5151
rect 14371 5146 14472 5149
rect 14371 5127 14436 5146
rect 12781 5112 12816 5113
rect 12758 5107 12816 5112
rect 12758 5087 12761 5107
rect 12781 5093 12816 5107
rect 12836 5093 12845 5113
rect 12781 5085 12845 5093
rect 12807 5084 12845 5085
rect 12808 5083 12845 5084
rect 12911 5117 12947 5118
rect 13019 5117 13055 5118
rect 12911 5110 13055 5117
rect 12911 5109 12968 5110
rect 12911 5089 12919 5109
rect 12939 5090 12968 5109
rect 12993 5109 13055 5110
rect 12993 5090 13027 5109
rect 12939 5089 13027 5090
rect 13047 5089 13055 5109
rect 12911 5083 13055 5089
rect 13121 5113 13159 5121
rect 13227 5117 13263 5118
rect 13121 5093 13130 5113
rect 13150 5093 13159 5113
rect 13121 5084 13159 5093
rect 13178 5110 13263 5117
rect 13178 5090 13185 5110
rect 13206 5109 13263 5110
rect 13206 5090 13235 5109
rect 13178 5089 13235 5090
rect 13255 5089 13263 5109
rect 13121 5083 13158 5084
rect 13178 5083 13263 5089
rect 13329 5113 13367 5121
rect 13440 5117 13476 5118
rect 13329 5093 13338 5113
rect 13358 5093 13367 5113
rect 13329 5084 13367 5093
rect 13391 5109 13476 5117
rect 13391 5089 13448 5109
rect 13468 5089 13476 5109
rect 13329 5083 13366 5084
rect 13391 5083 13476 5089
rect 13542 5113 13580 5121
rect 13542 5093 13551 5113
rect 13571 5093 13580 5113
rect 14433 5119 14436 5127
rect 14465 5119 14472 5146
rect 14500 5122 14510 5149
rect 14539 5127 14621 5149
rect 14539 5122 14543 5127
rect 14500 5119 14543 5122
rect 14433 5105 14543 5119
rect 14809 5123 14856 5124
rect 14809 5114 14857 5123
rect 14809 5096 14828 5114
rect 14846 5096 14857 5114
rect 14809 5094 14857 5096
rect 13542 5084 13580 5093
rect 13542 5083 13579 5084
rect 12965 5062 13001 5083
rect 13391 5062 13422 5083
rect 12798 5058 12898 5062
rect 12798 5054 12860 5058
rect 12798 5028 12805 5054
rect 12831 5032 12860 5054
rect 12886 5032 12898 5058
rect 12831 5028 12898 5032
rect 12798 5025 12898 5028
rect 12966 5025 13001 5062
rect 13063 5059 13422 5062
rect 13063 5054 13285 5059
rect 13063 5030 13076 5054
rect 13100 5035 13285 5054
rect 13309 5035 13422 5059
rect 13100 5030 13422 5035
rect 13063 5026 13422 5030
rect 13489 5054 13638 5062
rect 13489 5034 13500 5054
rect 13520 5034 13638 5054
rect 14818 5056 14857 5094
rect 15195 5096 15235 5276
rect 15581 5269 15612 5322
rect 15642 5351 15679 5430
rect 15850 5427 16243 5447
rect 16263 5427 16266 5447
rect 16364 5431 16613 5453
rect 16782 5452 16823 5457
rect 17201 5454 17228 5632
rect 17879 5544 17906 5722
rect 18284 5719 18325 5724
rect 18494 5723 18743 5745
rect 18841 5729 18844 5749
rect 18864 5729 19257 5749
rect 19428 5746 19465 5825
rect 19495 5854 19526 5907
rect 19872 5900 19912 6080
rect 19872 5882 19882 5900
rect 19900 5882 19912 5900
rect 19872 5877 19912 5882
rect 19872 5873 19909 5877
rect 19545 5854 19582 5855
rect 19495 5845 19582 5854
rect 19495 5825 19553 5845
rect 19573 5825 19582 5845
rect 19495 5815 19582 5825
rect 19641 5845 19678 5855
rect 19641 5825 19649 5845
rect 19669 5825 19678 5845
rect 19495 5814 19526 5815
rect 19490 5746 19600 5759
rect 19641 5746 19678 5825
rect 19875 5810 19912 5811
rect 19871 5801 19912 5810
rect 19871 5783 19884 5801
rect 19902 5783 19912 5801
rect 19871 5774 19912 5783
rect 19871 5754 19911 5774
rect 19428 5744 19678 5746
rect 19428 5741 19529 5744
rect 17946 5684 18010 5696
rect 18286 5692 18323 5719
rect 18494 5692 18531 5723
rect 18707 5721 18743 5723
rect 19428 5722 19493 5741
rect 18707 5692 18744 5721
rect 19490 5714 19493 5722
rect 19522 5714 19529 5741
rect 19557 5717 19567 5744
rect 19596 5722 19678 5744
rect 19786 5744 19911 5754
rect 19786 5725 19794 5744
rect 19819 5725 19911 5744
rect 19596 5717 19600 5722
rect 19786 5718 19911 5725
rect 19557 5714 19600 5717
rect 19490 5700 19600 5714
rect 17946 5683 17981 5684
rect 17923 5678 17981 5683
rect 17923 5658 17926 5678
rect 17946 5664 17981 5678
rect 18001 5664 18010 5684
rect 17946 5656 18010 5664
rect 17972 5655 18010 5656
rect 17973 5654 18010 5655
rect 18076 5688 18112 5689
rect 18184 5688 18220 5689
rect 18076 5680 18220 5688
rect 18076 5660 18084 5680
rect 18104 5677 18192 5680
rect 18104 5660 18136 5677
rect 18156 5660 18192 5677
rect 18212 5660 18220 5680
rect 18076 5654 18220 5660
rect 18286 5684 18324 5692
rect 18392 5688 18428 5689
rect 18286 5664 18295 5684
rect 18315 5664 18324 5684
rect 18286 5655 18324 5664
rect 18343 5681 18428 5688
rect 18343 5661 18350 5681
rect 18371 5680 18428 5681
rect 18371 5661 18400 5680
rect 18343 5660 18400 5661
rect 18420 5660 18428 5680
rect 18286 5654 18323 5655
rect 18343 5654 18428 5660
rect 18494 5684 18532 5692
rect 18605 5688 18641 5689
rect 18494 5664 18503 5684
rect 18523 5664 18532 5684
rect 18494 5655 18532 5664
rect 18556 5680 18641 5688
rect 18556 5660 18613 5680
rect 18633 5660 18641 5680
rect 18494 5654 18531 5655
rect 18556 5654 18641 5660
rect 18707 5684 18745 5692
rect 18707 5664 18716 5684
rect 18736 5664 18745 5684
rect 18707 5655 18745 5664
rect 19871 5670 19911 5718
rect 18707 5654 18744 5655
rect 18130 5633 18166 5654
rect 18556 5633 18587 5654
rect 19871 5652 19882 5670
rect 19900 5652 19911 5670
rect 19871 5644 19911 5652
rect 19872 5643 19909 5644
rect 17963 5629 18063 5633
rect 17963 5625 18025 5629
rect 17963 5599 17970 5625
rect 17996 5603 18025 5625
rect 18051 5603 18063 5629
rect 17996 5599 18063 5603
rect 17963 5596 18063 5599
rect 18131 5596 18166 5633
rect 18228 5630 18587 5633
rect 18228 5625 18450 5630
rect 18228 5601 18241 5625
rect 18265 5606 18450 5625
rect 18474 5606 18587 5630
rect 18265 5601 18587 5606
rect 18228 5597 18587 5601
rect 18654 5625 18803 5633
rect 18654 5605 18665 5625
rect 18685 5605 18803 5625
rect 18654 5598 18803 5605
rect 19243 5602 19757 5603
rect 18654 5597 18695 5598
rect 17978 5544 18015 5545
rect 18074 5544 18111 5545
rect 18130 5544 18166 5596
rect 18185 5544 18222 5545
rect 17878 5535 18016 5544
rect 17878 5515 17987 5535
rect 18007 5515 18016 5535
rect 17878 5508 18016 5515
rect 18074 5535 18222 5544
rect 18074 5515 18083 5535
rect 18103 5515 18193 5535
rect 18213 5515 18222 5535
rect 17878 5506 17974 5508
rect 18074 5505 18222 5515
rect 18281 5535 18318 5545
rect 18393 5544 18430 5545
rect 18374 5542 18430 5544
rect 18281 5515 18289 5535
rect 18309 5515 18318 5535
rect 18130 5504 18166 5505
rect 17060 5452 17228 5454
rect 16782 5446 17228 5452
rect 15850 5422 16266 5427
rect 16445 5425 16556 5431
rect 15850 5421 16191 5422
rect 15794 5361 15825 5362
rect 15642 5331 15651 5351
rect 15671 5331 15679 5351
rect 15642 5321 15679 5331
rect 15738 5354 15825 5361
rect 15738 5351 15799 5354
rect 15738 5331 15747 5351
rect 15767 5334 15799 5351
rect 15820 5334 15825 5354
rect 15767 5331 15825 5334
rect 15738 5324 15825 5331
rect 15850 5351 15887 5421
rect 16153 5420 16190 5421
rect 16445 5417 16486 5425
rect 16445 5397 16453 5417
rect 16472 5397 16486 5417
rect 16445 5395 16486 5397
rect 16514 5417 16556 5425
rect 16514 5397 16530 5417
rect 16549 5397 16556 5417
rect 16782 5424 16788 5446
rect 16814 5426 17228 5446
rect 17978 5445 18015 5446
rect 18281 5445 18318 5515
rect 18343 5535 18430 5542
rect 18343 5532 18401 5535
rect 18343 5512 18348 5532
rect 18369 5515 18401 5532
rect 18421 5515 18430 5535
rect 18369 5512 18430 5515
rect 18343 5505 18430 5512
rect 18489 5535 18526 5545
rect 18489 5515 18497 5535
rect 18517 5515 18526 5535
rect 18343 5504 18374 5505
rect 17977 5444 18318 5445
rect 16814 5424 16823 5426
rect 17060 5425 17228 5426
rect 17902 5439 18318 5444
rect 16782 5415 16823 5424
rect 17902 5419 17905 5439
rect 17925 5419 18318 5439
rect 18489 5436 18526 5515
rect 18556 5544 18587 5597
rect 19224 5586 19757 5602
rect 19224 5575 19756 5586
rect 19875 5577 19912 5581
rect 18606 5544 18643 5545
rect 18556 5535 18643 5544
rect 18556 5515 18614 5535
rect 18634 5515 18643 5535
rect 18556 5505 18643 5515
rect 18702 5535 18739 5545
rect 18702 5515 18710 5535
rect 18730 5515 18739 5535
rect 18556 5504 18587 5505
rect 18551 5436 18661 5449
rect 18702 5436 18739 5515
rect 18489 5434 18739 5436
rect 18489 5431 18590 5434
rect 18489 5412 18554 5431
rect 18551 5404 18554 5412
rect 18583 5404 18590 5431
rect 18618 5407 18628 5434
rect 18657 5412 18739 5434
rect 18817 5506 18985 5507
rect 19224 5506 19262 5575
rect 18817 5486 19262 5506
rect 19489 5537 19600 5552
rect 19489 5535 19531 5537
rect 19489 5515 19496 5535
rect 19515 5515 19531 5535
rect 19489 5507 19531 5515
rect 19559 5535 19600 5537
rect 19559 5515 19573 5535
rect 19592 5515 19600 5535
rect 19559 5507 19600 5515
rect 19489 5501 19600 5507
rect 19722 5512 19756 5575
rect 19874 5571 19912 5577
rect 19874 5553 19884 5571
rect 19902 5553 19912 5571
rect 19874 5544 19912 5553
rect 19874 5512 19908 5544
rect 18817 5480 19261 5486
rect 18817 5478 18985 5480
rect 18657 5407 18661 5412
rect 18618 5404 18661 5407
rect 16514 5395 16556 5397
rect 16445 5380 16556 5395
rect 17641 5386 17689 5400
rect 18551 5390 18661 5404
rect 16002 5361 16038 5362
rect 15850 5331 15859 5351
rect 15879 5331 15887 5351
rect 15738 5322 15794 5324
rect 15738 5321 15775 5322
rect 15850 5321 15887 5331
rect 15946 5351 16094 5361
rect 16194 5358 16290 5360
rect 15946 5331 15955 5351
rect 15975 5331 16065 5351
rect 16085 5331 16094 5351
rect 15946 5322 16094 5331
rect 16152 5351 16290 5358
rect 16152 5331 16161 5351
rect 16181 5331 16290 5351
rect 16152 5322 16290 5331
rect 17641 5346 17654 5386
rect 17681 5346 17689 5386
rect 17641 5328 17689 5346
rect 15946 5321 15983 5322
rect 16002 5270 16038 5322
rect 16057 5321 16094 5322
rect 16153 5321 16190 5322
rect 15473 5268 15514 5269
rect 15365 5261 15514 5268
rect 15365 5241 15483 5261
rect 15503 5241 15514 5261
rect 15365 5233 15514 5241
rect 15581 5265 15940 5269
rect 15581 5260 15903 5265
rect 15581 5236 15694 5260
rect 15718 5241 15903 5260
rect 15927 5241 15940 5265
rect 15718 5236 15940 5241
rect 15581 5233 15940 5236
rect 16002 5233 16037 5270
rect 16105 5267 16205 5270
rect 16105 5263 16172 5267
rect 16105 5237 16117 5263
rect 16143 5241 16172 5263
rect 16198 5241 16205 5267
rect 16143 5237 16205 5241
rect 16105 5233 16205 5237
rect 15581 5212 15612 5233
rect 16002 5212 16038 5233
rect 15424 5211 15461 5212
rect 15423 5202 15461 5211
rect 15423 5182 15432 5202
rect 15452 5182 15461 5202
rect 15423 5174 15461 5182
rect 15527 5206 15612 5212
rect 15637 5211 15674 5212
rect 15527 5186 15535 5206
rect 15555 5186 15612 5206
rect 15527 5178 15612 5186
rect 15636 5202 15674 5211
rect 15636 5182 15645 5202
rect 15665 5182 15674 5202
rect 15527 5177 15563 5178
rect 15636 5174 15674 5182
rect 15740 5206 15825 5212
rect 15845 5211 15882 5212
rect 15740 5186 15748 5206
rect 15768 5205 15825 5206
rect 15768 5186 15797 5205
rect 15740 5185 15797 5186
rect 15818 5185 15825 5205
rect 15740 5178 15825 5185
rect 15844 5202 15882 5211
rect 15844 5182 15853 5202
rect 15873 5182 15882 5202
rect 15740 5177 15776 5178
rect 15844 5174 15882 5182
rect 15948 5206 16092 5212
rect 15948 5186 15956 5206
rect 15976 5203 16064 5206
rect 15976 5186 16007 5203
rect 15948 5183 16007 5186
rect 16030 5186 16064 5203
rect 16084 5186 16092 5206
rect 16030 5183 16092 5186
rect 15948 5178 16092 5183
rect 15948 5177 15984 5178
rect 16056 5177 16092 5178
rect 16158 5211 16195 5212
rect 16158 5210 16196 5211
rect 16158 5202 16222 5210
rect 16158 5182 16167 5202
rect 16187 5188 16222 5202
rect 16242 5188 16245 5208
rect 16187 5183 16245 5188
rect 16187 5182 16222 5183
rect 15424 5145 15461 5174
rect 15425 5143 15461 5145
rect 15637 5143 15674 5174
rect 15425 5121 15674 5143
rect 15845 5142 15882 5174
rect 16158 5170 16222 5182
rect 16262 5144 16289 5322
rect 17636 5221 17689 5328
rect 18817 5300 18844 5478
rect 18884 5440 18948 5452
rect 19224 5448 19261 5480
rect 19432 5479 19681 5501
rect 19722 5480 19908 5512
rect 19736 5479 19908 5480
rect 19432 5448 19469 5479
rect 19645 5477 19681 5479
rect 19645 5448 19682 5477
rect 19874 5451 19908 5479
rect 18884 5439 18919 5440
rect 18861 5434 18919 5439
rect 18861 5414 18864 5434
rect 18884 5420 18919 5434
rect 18939 5420 18948 5440
rect 18884 5412 18948 5420
rect 18910 5411 18948 5412
rect 18911 5410 18948 5411
rect 19014 5444 19050 5445
rect 19122 5444 19158 5445
rect 19014 5437 19158 5444
rect 19014 5436 19074 5437
rect 19014 5416 19022 5436
rect 19042 5417 19074 5436
rect 19099 5436 19158 5437
rect 19099 5417 19130 5436
rect 19042 5416 19130 5417
rect 19150 5416 19158 5436
rect 19014 5410 19158 5416
rect 19224 5440 19262 5448
rect 19330 5444 19366 5445
rect 19224 5420 19233 5440
rect 19253 5420 19262 5440
rect 19224 5411 19262 5420
rect 19281 5437 19366 5444
rect 19281 5417 19288 5437
rect 19309 5436 19366 5437
rect 19309 5417 19338 5436
rect 19281 5416 19338 5417
rect 19358 5416 19366 5436
rect 19224 5410 19261 5411
rect 19281 5410 19366 5416
rect 19432 5440 19470 5448
rect 19543 5444 19579 5445
rect 19432 5420 19441 5440
rect 19461 5420 19470 5440
rect 19432 5411 19470 5420
rect 19494 5436 19579 5444
rect 19494 5416 19551 5436
rect 19571 5416 19579 5436
rect 19432 5410 19469 5411
rect 19494 5410 19579 5416
rect 19645 5440 19683 5448
rect 19645 5420 19654 5440
rect 19674 5420 19683 5440
rect 19645 5411 19683 5420
rect 19872 5441 19909 5451
rect 19872 5423 19882 5441
rect 19900 5423 19909 5441
rect 19872 5414 19909 5423
rect 19874 5413 19908 5414
rect 19645 5410 19682 5411
rect 19068 5389 19104 5410
rect 19494 5389 19525 5410
rect 18901 5385 19001 5389
rect 18901 5381 18963 5385
rect 18901 5355 18908 5381
rect 18934 5359 18963 5381
rect 18989 5359 19001 5385
rect 18934 5355 19001 5359
rect 18901 5352 19001 5355
rect 19069 5352 19104 5389
rect 19166 5386 19525 5389
rect 19166 5381 19388 5386
rect 19166 5357 19179 5381
rect 19203 5362 19388 5381
rect 19412 5362 19525 5386
rect 19203 5357 19525 5362
rect 19166 5353 19525 5357
rect 19592 5381 19741 5389
rect 19592 5361 19603 5381
rect 19623 5361 19741 5381
rect 19592 5354 19741 5361
rect 19592 5353 19633 5354
rect 18916 5300 18953 5301
rect 19012 5300 19049 5301
rect 19068 5300 19104 5352
rect 19123 5300 19160 5301
rect 18816 5291 18954 5300
rect 18816 5271 18925 5291
rect 18945 5271 18954 5291
rect 18442 5251 18553 5266
rect 18816 5264 18954 5271
rect 19012 5291 19160 5300
rect 19012 5271 19021 5291
rect 19041 5271 19131 5291
rect 19151 5271 19160 5291
rect 18816 5262 18912 5264
rect 19012 5261 19160 5271
rect 19219 5291 19256 5301
rect 19331 5300 19368 5301
rect 19312 5298 19368 5300
rect 19219 5271 19227 5291
rect 19247 5271 19256 5291
rect 19068 5260 19104 5261
rect 18442 5249 18484 5251
rect 18442 5229 18449 5249
rect 18468 5229 18484 5249
rect 18442 5221 18484 5229
rect 18512 5249 18553 5251
rect 18512 5229 18526 5249
rect 18545 5229 18553 5249
rect 18512 5221 18553 5229
rect 17636 5220 17938 5221
rect 16555 5199 16665 5213
rect 16555 5196 16598 5199
rect 16555 5191 16559 5196
rect 16121 5142 16289 5144
rect 15845 5139 16289 5142
rect 15506 5115 15617 5121
rect 15506 5107 15547 5115
rect 13489 5027 13638 5034
rect 14170 5037 14208 5039
rect 14818 5037 14860 5056
rect 13489 5026 13530 5027
rect 12965 5021 13001 5025
rect 12965 4992 13002 5021
rect 12813 4973 12850 4974
rect 12909 4973 12946 4974
rect 12965 4973 13001 4992
rect 13020 4973 13057 4974
rect 12713 4964 12851 4973
rect 12713 4944 12822 4964
rect 12842 4944 12851 4964
rect 12713 4937 12851 4944
rect 12909 4964 13057 4973
rect 12909 4944 12918 4964
rect 12938 4944 13028 4964
rect 13048 4944 13057 4964
rect 12713 4935 12809 4937
rect 12909 4934 13057 4944
rect 13116 4964 13153 4974
rect 13228 4973 13265 4974
rect 13209 4971 13265 4973
rect 13116 4944 13124 4964
rect 13144 4944 13153 4964
rect 12965 4933 13001 4934
rect 12813 4874 12850 4875
rect 13116 4874 13153 4944
rect 13178 4964 13265 4971
rect 13178 4961 13236 4964
rect 13178 4941 13183 4961
rect 13204 4944 13236 4961
rect 13256 4944 13265 4964
rect 13204 4941 13265 4944
rect 13178 4934 13265 4941
rect 13324 4964 13361 4974
rect 13324 4944 13332 4964
rect 13352 4944 13361 4964
rect 13178 4933 13209 4934
rect 12812 4873 13153 4874
rect 12737 4868 13153 4873
rect 12362 4841 12415 4849
rect 12737 4848 12740 4868
rect 12760 4848 13153 4868
rect 13324 4865 13361 4944
rect 13391 4973 13422 5026
rect 14170 5014 14860 5037
rect 15195 5052 15234 5096
rect 15506 5087 15514 5107
rect 15533 5087 15547 5107
rect 15506 5085 15547 5087
rect 15575 5107 15617 5115
rect 15575 5087 15591 5107
rect 15610 5087 15617 5107
rect 15575 5086 15617 5087
rect 15843 5116 16289 5139
rect 15575 5085 15618 5086
rect 15506 5066 15618 5085
rect 15195 5028 15235 5052
rect 15535 5028 15582 5029
rect 15843 5028 15881 5116
rect 16121 5115 16289 5116
rect 16477 5169 16559 5191
rect 16588 5169 16598 5196
rect 16626 5172 16633 5199
rect 16662 5191 16665 5199
rect 17636 5194 18214 5220
rect 18442 5215 18553 5221
rect 17636 5192 17938 5194
rect 17636 5191 17822 5192
rect 16662 5172 16727 5191
rect 16626 5169 16727 5172
rect 16477 5167 16727 5169
rect 16477 5088 16514 5167
rect 16555 5154 16665 5167
rect 16629 5098 16660 5099
rect 16477 5068 16486 5088
rect 16506 5068 16514 5088
rect 16477 5058 16514 5068
rect 16573 5088 16660 5098
rect 16573 5068 16582 5088
rect 16602 5068 16660 5088
rect 16573 5059 16660 5068
rect 16573 5058 16610 5059
rect 15195 5018 15881 5028
rect 14170 5004 14856 5014
rect 13441 4973 13478 4974
rect 13391 4964 13478 4973
rect 13391 4944 13449 4964
rect 13469 4944 13478 4964
rect 13391 4934 13478 4944
rect 13537 4964 13574 4974
rect 13537 4944 13545 4964
rect 13565 4944 13574 4964
rect 13391 4933 13422 4934
rect 13386 4865 13496 4878
rect 13537 4865 13574 4944
rect 13324 4863 13574 4865
rect 13324 4860 13425 4863
rect 13324 4841 13389 4860
rect 12229 4840 12415 4841
rect 12113 4838 12415 4840
rect 11498 4811 11609 4817
rect 11837 4812 12415 4838
rect 13386 4833 13389 4841
rect 13418 4833 13425 4860
rect 13453 4836 13463 4863
rect 13492 4841 13574 4863
rect 13762 4916 13930 4917
rect 14170 4916 14208 5004
rect 14469 5003 14516 5004
rect 14816 4980 14856 5004
rect 14433 4947 14545 4966
rect 14433 4946 14476 4947
rect 13762 4893 14208 4916
rect 14434 4945 14476 4946
rect 14434 4925 14441 4945
rect 14460 4925 14476 4945
rect 14434 4917 14476 4925
rect 14504 4945 14545 4947
rect 14504 4925 14518 4945
rect 14537 4925 14545 4945
rect 14817 4936 14856 4980
rect 15191 4995 15881 5018
rect 16629 5006 16660 5059
rect 16690 5088 16727 5167
rect 16898 5164 17291 5184
rect 17311 5164 17314 5184
rect 17636 5183 17689 5191
rect 16898 5159 17314 5164
rect 16898 5158 17239 5159
rect 16842 5098 16873 5099
rect 16690 5068 16699 5088
rect 16719 5068 16727 5088
rect 16690 5058 16727 5068
rect 16786 5091 16873 5098
rect 16786 5088 16847 5091
rect 16786 5068 16795 5088
rect 16815 5071 16847 5088
rect 16868 5071 16873 5091
rect 16815 5068 16873 5071
rect 16786 5061 16873 5068
rect 16898 5088 16935 5158
rect 17201 5157 17238 5158
rect 17050 5098 17086 5099
rect 16898 5068 16907 5088
rect 16927 5068 16935 5088
rect 16786 5059 16842 5061
rect 16786 5058 16823 5059
rect 16898 5058 16935 5068
rect 16994 5088 17142 5098
rect 17242 5095 17338 5097
rect 16994 5068 17003 5088
rect 17023 5068 17113 5088
rect 17133 5068 17142 5088
rect 16994 5059 17142 5068
rect 17200 5088 17338 5095
rect 17200 5068 17209 5088
rect 17229 5068 17338 5088
rect 17200 5059 17338 5068
rect 16994 5058 17031 5059
rect 17050 5007 17086 5059
rect 17105 5058 17142 5059
rect 17201 5058 17238 5059
rect 16521 5005 16562 5006
rect 15191 4976 15233 4995
rect 15843 4993 15881 4995
rect 16413 4998 16562 5005
rect 14504 4917 14545 4925
rect 14434 4911 14545 4917
rect 13762 4890 14206 4893
rect 13762 4888 13930 4890
rect 13492 4836 13496 4841
rect 13453 4833 13496 4836
rect 13386 4819 13496 4833
rect 12113 4811 12415 4812
rect 11498 4803 11539 4811
rect 11498 4783 11506 4803
rect 11525 4783 11539 4803
rect 11498 4781 11539 4783
rect 11567 4803 11609 4811
rect 11567 4783 11583 4803
rect 11602 4783 11609 4803
rect 11567 4781 11609 4783
rect 10947 4771 10983 4772
rect 10795 4741 10804 4761
rect 10824 4741 10832 4761
rect 10683 4732 10739 4734
rect 10683 4731 10720 4732
rect 10795 4731 10832 4741
rect 10891 4761 11039 4771
rect 11139 4768 11235 4770
rect 10891 4741 10900 4761
rect 10920 4741 11010 4761
rect 11030 4741 11039 4761
rect 10891 4732 11039 4741
rect 11097 4761 11235 4768
rect 11498 4766 11609 4781
rect 11097 4741 11106 4761
rect 11126 4741 11235 4761
rect 11097 4732 11235 4741
rect 10891 4731 10928 4732
rect 10947 4680 10983 4732
rect 11002 4731 11039 4732
rect 11098 4731 11135 4732
rect 10418 4678 10459 4679
rect 9840 4666 9881 4675
rect 10310 4671 10459 4678
rect 9840 4646 9880 4666
rect 9397 4636 9647 4638
rect 9397 4633 9498 4636
rect 7915 4576 7979 4588
rect 8255 4584 8292 4611
rect 8463 4584 8500 4615
rect 8676 4613 8712 4615
rect 9397 4614 9462 4633
rect 8676 4584 8713 4613
rect 9459 4606 9462 4614
rect 9491 4606 9498 4633
rect 9526 4609 9536 4636
rect 9565 4614 9647 4636
rect 9755 4636 9880 4646
rect 10310 4651 10428 4671
rect 10448 4651 10459 4671
rect 10310 4643 10459 4651
rect 10526 4675 10885 4679
rect 10526 4670 10848 4675
rect 10526 4646 10639 4670
rect 10663 4651 10848 4670
rect 10872 4651 10885 4675
rect 10663 4646 10885 4651
rect 10526 4643 10885 4646
rect 10947 4643 10982 4680
rect 11050 4677 11150 4680
rect 11050 4673 11117 4677
rect 11050 4647 11062 4673
rect 11088 4651 11117 4673
rect 11143 4651 11150 4677
rect 11088 4647 11150 4651
rect 11050 4643 11150 4647
rect 9755 4617 9763 4636
rect 9788 4617 9880 4636
rect 10526 4622 10557 4643
rect 10947 4622 10983 4643
rect 10369 4621 10406 4622
rect 10143 4618 10177 4619
rect 9565 4609 9569 4614
rect 9755 4610 9880 4617
rect 9526 4606 9569 4609
rect 9459 4592 9569 4606
rect 7915 4575 7950 4576
rect 7892 4570 7950 4575
rect 7892 4550 7895 4570
rect 7915 4556 7950 4570
rect 7970 4556 7979 4576
rect 7915 4548 7979 4556
rect 7941 4547 7979 4548
rect 7942 4546 7979 4547
rect 8045 4580 8081 4581
rect 8153 4580 8189 4581
rect 8045 4572 8189 4580
rect 8045 4552 8053 4572
rect 8073 4552 8161 4572
rect 8181 4552 8189 4572
rect 8045 4546 8189 4552
rect 8255 4576 8293 4584
rect 8361 4580 8397 4581
rect 8255 4556 8264 4576
rect 8284 4556 8293 4576
rect 8255 4547 8293 4556
rect 8312 4573 8397 4580
rect 8312 4553 8319 4573
rect 8340 4572 8397 4573
rect 8340 4553 8369 4572
rect 8312 4552 8369 4553
rect 8389 4552 8397 4572
rect 8255 4546 8292 4547
rect 8312 4546 8397 4552
rect 8463 4576 8501 4584
rect 8574 4580 8610 4581
rect 8463 4556 8472 4576
rect 8492 4556 8501 4576
rect 8463 4547 8501 4556
rect 8525 4572 8610 4580
rect 8525 4552 8582 4572
rect 8602 4552 8610 4572
rect 8463 4546 8500 4547
rect 8525 4546 8610 4552
rect 8676 4576 8714 4584
rect 8676 4556 8685 4576
rect 8705 4556 8714 4576
rect 8676 4547 8714 4556
rect 9840 4562 9880 4610
rect 10142 4609 10179 4618
rect 10142 4591 10151 4609
rect 10169 4591 10179 4609
rect 10142 4581 10179 4591
rect 10368 4612 10406 4621
rect 10368 4592 10377 4612
rect 10397 4592 10406 4612
rect 10368 4584 10406 4592
rect 10472 4616 10557 4622
rect 10582 4621 10619 4622
rect 10472 4596 10480 4616
rect 10500 4596 10557 4616
rect 10472 4588 10557 4596
rect 10581 4612 10619 4621
rect 10581 4592 10590 4612
rect 10610 4592 10619 4612
rect 10472 4587 10508 4588
rect 10581 4584 10619 4592
rect 10685 4616 10770 4622
rect 10790 4621 10827 4622
rect 10685 4596 10693 4616
rect 10713 4615 10770 4616
rect 10713 4596 10742 4615
rect 10685 4595 10742 4596
rect 10763 4595 10770 4615
rect 10685 4588 10770 4595
rect 10789 4612 10827 4621
rect 10789 4592 10798 4612
rect 10818 4592 10827 4612
rect 10685 4587 10721 4588
rect 10789 4584 10827 4592
rect 10893 4616 11037 4622
rect 10893 4596 10901 4616
rect 10921 4615 11009 4616
rect 10921 4596 10952 4615
rect 10893 4595 10952 4596
rect 10977 4596 11009 4615
rect 11029 4596 11037 4616
rect 10977 4595 11037 4596
rect 10893 4588 11037 4595
rect 10893 4587 10929 4588
rect 11001 4587 11037 4588
rect 11103 4621 11140 4622
rect 11103 4620 11141 4621
rect 11103 4612 11167 4620
rect 11103 4592 11112 4612
rect 11132 4598 11167 4612
rect 11187 4598 11190 4618
rect 11132 4593 11190 4598
rect 11132 4592 11167 4593
rect 8676 4546 8713 4547
rect 8099 4525 8135 4546
rect 8525 4525 8556 4546
rect 9840 4544 9851 4562
rect 9869 4544 9880 4562
rect 9840 4536 9880 4544
rect 10143 4553 10177 4581
rect 10369 4555 10406 4584
rect 10370 4553 10406 4555
rect 10582 4553 10619 4584
rect 10143 4552 10315 4553
rect 9841 4535 9878 4536
rect 7932 4521 8032 4525
rect 7932 4517 7994 4521
rect 7932 4491 7939 4517
rect 7965 4495 7994 4517
rect 8020 4495 8032 4521
rect 7965 4491 8032 4495
rect 7932 4488 8032 4491
rect 8100 4488 8135 4525
rect 8197 4522 8556 4525
rect 8197 4517 8419 4522
rect 8197 4493 8210 4517
rect 8234 4498 8419 4517
rect 8443 4498 8556 4522
rect 8234 4493 8556 4498
rect 8197 4489 8556 4493
rect 8623 4517 8772 4525
rect 8623 4497 8634 4517
rect 8654 4497 8772 4517
rect 8623 4490 8772 4497
rect 10143 4520 10329 4552
rect 10370 4531 10619 4553
rect 10790 4552 10827 4584
rect 11103 4580 11167 4592
rect 11207 4554 11234 4732
rect 12362 4704 12415 4811
rect 13762 4710 13789 4888
rect 13829 4850 13893 4862
rect 14169 4858 14206 4890
rect 14377 4889 14626 4911
rect 14377 4858 14414 4889
rect 14590 4887 14626 4889
rect 14590 4858 14627 4887
rect 13829 4849 13864 4850
rect 13806 4844 13864 4849
rect 13806 4824 13809 4844
rect 13829 4830 13864 4844
rect 13884 4830 13893 4850
rect 13829 4822 13893 4830
rect 13855 4821 13893 4822
rect 13856 4820 13893 4821
rect 13959 4854 13995 4855
rect 14067 4854 14103 4855
rect 13959 4849 14103 4854
rect 13959 4846 14021 4849
rect 13959 4826 13967 4846
rect 13987 4829 14021 4846
rect 14044 4846 14103 4849
rect 14044 4829 14075 4846
rect 13987 4826 14075 4829
rect 14095 4826 14103 4846
rect 13959 4820 14103 4826
rect 14169 4850 14207 4858
rect 14275 4854 14311 4855
rect 14169 4830 14178 4850
rect 14198 4830 14207 4850
rect 14169 4821 14207 4830
rect 14226 4847 14311 4854
rect 14226 4827 14233 4847
rect 14254 4846 14311 4847
rect 14254 4827 14283 4846
rect 14226 4826 14283 4827
rect 14303 4826 14311 4846
rect 14169 4820 14206 4821
rect 14226 4820 14311 4826
rect 14377 4850 14415 4858
rect 14488 4854 14524 4855
rect 14377 4830 14386 4850
rect 14406 4830 14415 4850
rect 14377 4821 14415 4830
rect 14439 4846 14524 4854
rect 14439 4826 14496 4846
rect 14516 4826 14524 4846
rect 14377 4820 14414 4821
rect 14439 4820 14524 4826
rect 14590 4850 14628 4858
rect 14590 4830 14599 4850
rect 14619 4830 14628 4850
rect 14590 4821 14628 4830
rect 14590 4820 14627 4821
rect 14013 4799 14049 4820
rect 14439 4799 14470 4820
rect 13846 4795 13946 4799
rect 13846 4791 13908 4795
rect 13846 4765 13853 4791
rect 13879 4769 13908 4791
rect 13934 4769 13946 4795
rect 13879 4765 13946 4769
rect 13846 4762 13946 4765
rect 14014 4762 14049 4799
rect 14111 4796 14470 4799
rect 14111 4791 14333 4796
rect 14111 4767 14124 4791
rect 14148 4772 14333 4791
rect 14357 4772 14470 4796
rect 14148 4767 14470 4772
rect 14111 4763 14470 4767
rect 14537 4791 14686 4799
rect 14537 4771 14548 4791
rect 14568 4771 14686 4791
rect 14537 4764 14686 4771
rect 14537 4763 14578 4764
rect 13861 4710 13898 4711
rect 13957 4710 13994 4711
rect 14013 4710 14049 4762
rect 14068 4710 14105 4711
rect 12362 4686 12410 4704
rect 12362 4646 12370 4686
rect 12397 4646 12410 4686
rect 13761 4701 13899 4710
rect 13761 4681 13870 4701
rect 13890 4681 13899 4701
rect 13761 4674 13899 4681
rect 13957 4701 14105 4710
rect 13957 4681 13966 4701
rect 13986 4681 14076 4701
rect 14096 4681 14105 4701
rect 13761 4672 13857 4674
rect 13957 4671 14105 4681
rect 14164 4701 14201 4711
rect 14276 4710 14313 4711
rect 14257 4708 14313 4710
rect 14164 4681 14172 4701
rect 14192 4681 14201 4701
rect 14013 4670 14049 4671
rect 11390 4628 11500 4642
rect 12362 4632 12410 4646
rect 13495 4637 13606 4652
rect 13495 4635 13537 4637
rect 11390 4625 11433 4628
rect 11390 4620 11394 4625
rect 11066 4552 11234 4554
rect 10790 4546 11234 4552
rect 9212 4494 9726 4495
rect 8623 4489 8664 4490
rect 8099 4453 8135 4488
rect 7947 4436 7984 4437
rect 8043 4436 8080 4437
rect 8099 4436 8106 4453
rect 7847 4427 7985 4436
rect 7847 4407 7956 4427
rect 7976 4407 7985 4427
rect 7847 4400 7985 4407
rect 8043 4427 8106 4436
rect 8043 4407 8052 4427
rect 8072 4412 8106 4427
rect 8127 4436 8135 4453
rect 8154 4436 8191 4437
rect 8127 4427 8191 4436
rect 8127 4412 8162 4427
rect 8072 4407 8162 4412
rect 8182 4407 8191 4427
rect 7847 4398 7943 4400
rect 8043 4397 8191 4407
rect 8250 4427 8287 4437
rect 8362 4436 8399 4437
rect 8343 4434 8399 4436
rect 8250 4407 8258 4427
rect 8278 4407 8287 4427
rect 8099 4396 8135 4397
rect 7029 4344 7197 4346
rect 6751 4338 7197 4344
rect 5819 4314 6235 4319
rect 6414 4317 6525 4323
rect 5819 4313 6160 4314
rect 5763 4253 5794 4254
rect 5611 4223 5620 4243
rect 5640 4223 5648 4243
rect 5611 4213 5648 4223
rect 5707 4246 5794 4253
rect 5707 4243 5768 4246
rect 5707 4223 5716 4243
rect 5736 4226 5768 4243
rect 5789 4226 5794 4246
rect 5736 4223 5794 4226
rect 5707 4216 5794 4223
rect 5819 4243 5856 4313
rect 6122 4312 6159 4313
rect 6414 4309 6455 4317
rect 6414 4289 6422 4309
rect 6441 4289 6455 4309
rect 6414 4287 6455 4289
rect 6483 4309 6525 4317
rect 6483 4289 6499 4309
rect 6518 4289 6525 4309
rect 6751 4316 6757 4338
rect 6783 4318 7197 4338
rect 7947 4337 7984 4338
rect 8250 4337 8287 4407
rect 8312 4427 8399 4434
rect 8312 4424 8370 4427
rect 8312 4404 8317 4424
rect 8338 4407 8370 4424
rect 8390 4407 8399 4427
rect 8338 4404 8399 4407
rect 8312 4397 8399 4404
rect 8458 4427 8495 4437
rect 8458 4407 8466 4427
rect 8486 4407 8495 4427
rect 8312 4396 8343 4397
rect 7946 4336 8287 4337
rect 6783 4316 6792 4318
rect 7029 4317 7197 4318
rect 7871 4335 8287 4336
rect 7871 4331 8247 4335
rect 6751 4307 6792 4316
rect 7871 4311 7874 4331
rect 7894 4318 8247 4331
rect 8279 4318 8287 4335
rect 7894 4311 8287 4318
rect 8458 4328 8495 4407
rect 8525 4436 8556 4489
rect 9193 4478 9726 4494
rect 10143 4488 10177 4520
rect 10139 4479 10177 4488
rect 9193 4467 9725 4478
rect 9844 4469 9881 4473
rect 8575 4436 8612 4437
rect 8525 4427 8612 4436
rect 8525 4407 8583 4427
rect 8603 4407 8612 4427
rect 8525 4397 8612 4407
rect 8671 4427 8708 4437
rect 8671 4407 8679 4427
rect 8699 4407 8708 4427
rect 8525 4396 8556 4397
rect 8520 4328 8630 4341
rect 8671 4328 8708 4407
rect 8458 4326 8708 4328
rect 8458 4323 8559 4326
rect 8458 4304 8523 4323
rect 6483 4287 6525 4289
rect 6414 4272 6525 4287
rect 8520 4296 8523 4304
rect 8552 4296 8559 4323
rect 8587 4299 8597 4326
rect 8626 4304 8708 4326
rect 8786 4398 8954 4399
rect 9193 4398 9231 4467
rect 8786 4378 9231 4398
rect 9458 4429 9569 4444
rect 9458 4427 9500 4429
rect 9458 4407 9465 4427
rect 9484 4407 9500 4427
rect 9458 4399 9500 4407
rect 9528 4427 9569 4429
rect 9528 4407 9542 4427
rect 9561 4407 9569 4427
rect 9528 4399 9569 4407
rect 9458 4393 9569 4399
rect 9691 4404 9725 4467
rect 9843 4463 9881 4469
rect 9843 4445 9853 4463
rect 9871 4445 9881 4463
rect 10139 4461 10149 4479
rect 10167 4461 10177 4479
rect 10139 4455 10177 4461
rect 10295 4457 10329 4520
rect 10451 4525 10562 4531
rect 10451 4517 10492 4525
rect 10451 4497 10459 4517
rect 10478 4497 10492 4517
rect 10451 4495 10492 4497
rect 10520 4517 10562 4525
rect 10520 4497 10536 4517
rect 10555 4497 10562 4517
rect 10520 4495 10562 4497
rect 10451 4480 10562 4495
rect 10789 4526 11234 4546
rect 10789 4457 10827 4526
rect 11066 4525 11234 4526
rect 11312 4598 11394 4620
rect 11423 4598 11433 4625
rect 11461 4601 11468 4628
rect 11497 4620 11500 4628
rect 11497 4601 11562 4620
rect 11461 4598 11562 4601
rect 11312 4596 11562 4598
rect 11312 4517 11349 4596
rect 11390 4583 11500 4596
rect 11464 4527 11495 4528
rect 11312 4497 11321 4517
rect 11341 4497 11349 4517
rect 11312 4487 11349 4497
rect 11408 4517 11495 4527
rect 11408 4497 11417 4517
rect 11437 4497 11495 4517
rect 11408 4488 11495 4497
rect 11408 4487 11445 4488
rect 10139 4451 10176 4455
rect 10295 4446 10827 4457
rect 9843 4436 9881 4445
rect 9843 4404 9877 4436
rect 10294 4430 10827 4446
rect 11464 4435 11495 4488
rect 11525 4517 11562 4596
rect 11733 4593 12126 4613
rect 12146 4593 12149 4613
rect 13228 4608 13269 4617
rect 11733 4588 12149 4593
rect 12823 4606 12991 4607
rect 13228 4606 13237 4608
rect 11733 4587 12074 4588
rect 11677 4527 11708 4528
rect 11525 4497 11534 4517
rect 11554 4497 11562 4517
rect 11525 4487 11562 4497
rect 11621 4520 11708 4527
rect 11621 4517 11682 4520
rect 11621 4497 11630 4517
rect 11650 4500 11682 4517
rect 11703 4500 11708 4520
rect 11650 4497 11708 4500
rect 11621 4490 11708 4497
rect 11733 4517 11770 4587
rect 12036 4586 12073 4587
rect 12823 4586 13237 4606
rect 13263 4586 13269 4608
rect 13495 4615 13502 4635
rect 13521 4615 13537 4635
rect 13495 4607 13537 4615
rect 13565 4635 13606 4637
rect 13565 4615 13579 4635
rect 13598 4615 13606 4635
rect 13565 4607 13606 4615
rect 13861 4611 13898 4612
rect 14164 4611 14201 4681
rect 14226 4701 14313 4708
rect 14226 4698 14284 4701
rect 14226 4678 14231 4698
rect 14252 4681 14284 4698
rect 14304 4681 14313 4701
rect 14252 4678 14313 4681
rect 14226 4671 14313 4678
rect 14372 4701 14409 4711
rect 14372 4681 14380 4701
rect 14400 4681 14409 4701
rect 14226 4670 14257 4671
rect 13860 4610 14201 4611
rect 13495 4601 13606 4607
rect 13785 4605 14201 4610
rect 12823 4580 13269 4586
rect 12823 4578 12991 4580
rect 11885 4527 11921 4528
rect 11733 4497 11742 4517
rect 11762 4497 11770 4517
rect 11621 4488 11677 4490
rect 11621 4487 11658 4488
rect 11733 4487 11770 4497
rect 11829 4517 11977 4527
rect 12077 4524 12173 4526
rect 11829 4497 11838 4517
rect 11858 4497 11948 4517
rect 11968 4497 11977 4517
rect 11829 4488 11977 4497
rect 12035 4517 12173 4524
rect 12035 4497 12044 4517
rect 12064 4497 12173 4517
rect 12035 4488 12173 4497
rect 11829 4487 11866 4488
rect 11885 4436 11921 4488
rect 11940 4487 11977 4488
rect 12036 4487 12073 4488
rect 11356 4434 11397 4435
rect 10294 4429 10808 4430
rect 8786 4372 9230 4378
rect 8786 4370 8954 4372
rect 8626 4299 8630 4304
rect 8587 4296 8630 4299
rect 8520 4282 8630 4296
rect 5971 4253 6007 4254
rect 5819 4223 5828 4243
rect 5848 4223 5856 4243
rect 5707 4214 5763 4216
rect 5707 4213 5744 4214
rect 5819 4213 5856 4223
rect 5915 4243 6063 4253
rect 6163 4250 6259 4252
rect 5915 4223 5924 4243
rect 5944 4223 6034 4243
rect 6054 4223 6063 4243
rect 5915 4214 6063 4223
rect 6121 4243 6259 4250
rect 6121 4223 6130 4243
rect 6150 4223 6259 4243
rect 6121 4214 6259 4223
rect 5915 4213 5952 4214
rect 5971 4162 6007 4214
rect 6026 4213 6063 4214
rect 6122 4213 6159 4214
rect 5442 4160 5483 4161
rect 5334 4153 5483 4160
rect 5334 4133 5452 4153
rect 5472 4133 5483 4153
rect 5334 4125 5483 4133
rect 5550 4157 5909 4161
rect 5550 4152 5872 4157
rect 5550 4128 5663 4152
rect 5687 4133 5872 4152
rect 5896 4133 5909 4157
rect 5687 4128 5909 4133
rect 5550 4125 5909 4128
rect 5971 4125 6006 4162
rect 6074 4159 6174 4162
rect 6074 4155 6141 4159
rect 6074 4129 6086 4155
rect 6112 4133 6141 4155
rect 6167 4133 6174 4159
rect 6112 4129 6174 4133
rect 6074 4125 6174 4129
rect 5550 4104 5581 4125
rect 5971 4104 6007 4125
rect 5393 4103 5430 4104
rect 5392 4094 5430 4103
rect 5392 4074 5401 4094
rect 5421 4074 5430 4094
rect 5392 4066 5430 4074
rect 5496 4098 5581 4104
rect 5606 4103 5643 4104
rect 5496 4078 5504 4098
rect 5524 4078 5581 4098
rect 5496 4070 5581 4078
rect 5605 4094 5643 4103
rect 5605 4074 5614 4094
rect 5634 4074 5643 4094
rect 5496 4069 5532 4070
rect 5605 4066 5643 4074
rect 5709 4098 5794 4104
rect 5814 4103 5851 4104
rect 5709 4078 5717 4098
rect 5737 4097 5794 4098
rect 5737 4078 5766 4097
rect 5709 4077 5766 4078
rect 5787 4077 5794 4097
rect 5709 4070 5794 4077
rect 5813 4094 5851 4103
rect 5813 4074 5822 4094
rect 5842 4074 5851 4094
rect 5709 4069 5745 4070
rect 5813 4066 5851 4074
rect 5917 4098 6061 4104
rect 5917 4078 5925 4098
rect 5945 4095 6033 4098
rect 5945 4078 5976 4095
rect 5917 4075 5976 4078
rect 5999 4078 6033 4095
rect 6053 4078 6061 4098
rect 5999 4075 6061 4078
rect 5917 4070 6061 4075
rect 5917 4069 5953 4070
rect 6025 4069 6061 4070
rect 6127 4103 6164 4104
rect 6127 4102 6165 4103
rect 6127 4094 6191 4102
rect 6127 4074 6136 4094
rect 6156 4080 6191 4094
rect 6211 4080 6214 4100
rect 6156 4075 6214 4080
rect 6156 4074 6191 4075
rect 5393 4037 5430 4066
rect 5394 4035 5430 4037
rect 5606 4035 5643 4066
rect 5394 4013 5643 4035
rect 5814 4034 5851 4066
rect 6127 4062 6191 4074
rect 6231 4036 6258 4214
rect 8786 4192 8813 4370
rect 8853 4332 8917 4344
rect 9193 4340 9230 4372
rect 9401 4371 9650 4393
rect 9691 4372 9877 4404
rect 11248 4427 11397 4434
rect 11248 4407 11366 4427
rect 11386 4407 11397 4427
rect 11248 4399 11397 4407
rect 11464 4431 11823 4435
rect 11464 4426 11786 4431
rect 11464 4402 11577 4426
rect 11601 4407 11786 4426
rect 11810 4407 11823 4431
rect 11601 4402 11823 4407
rect 11464 4399 11823 4402
rect 11885 4399 11920 4436
rect 11988 4433 12088 4436
rect 11988 4429 12055 4433
rect 11988 4403 12000 4429
rect 12026 4407 12055 4429
rect 12081 4407 12088 4433
rect 12026 4403 12088 4407
rect 11988 4399 12088 4403
rect 10142 4388 10179 4389
rect 9705 4371 9877 4372
rect 9401 4340 9438 4371
rect 9614 4369 9650 4371
rect 9614 4340 9651 4369
rect 9843 4343 9877 4371
rect 10140 4380 10180 4388
rect 10140 4362 10151 4380
rect 10169 4362 10180 4380
rect 11464 4378 11495 4399
rect 11885 4378 11921 4399
rect 11307 4377 11344 4378
rect 8853 4331 8888 4332
rect 8830 4326 8888 4331
rect 8830 4306 8833 4326
rect 8853 4312 8888 4326
rect 8908 4312 8917 4332
rect 8853 4304 8917 4312
rect 8879 4303 8917 4304
rect 8880 4302 8917 4303
rect 8983 4336 9019 4337
rect 9091 4336 9127 4337
rect 8983 4329 9127 4336
rect 8983 4328 9043 4329
rect 8983 4308 8991 4328
rect 9011 4309 9043 4328
rect 9068 4328 9127 4329
rect 9068 4309 9099 4328
rect 9011 4308 9099 4309
rect 9119 4308 9127 4328
rect 8983 4302 9127 4308
rect 9193 4332 9231 4340
rect 9299 4336 9335 4337
rect 9193 4312 9202 4332
rect 9222 4312 9231 4332
rect 9193 4303 9231 4312
rect 9250 4329 9335 4336
rect 9250 4309 9257 4329
rect 9278 4328 9335 4329
rect 9278 4309 9307 4328
rect 9250 4308 9307 4309
rect 9327 4308 9335 4328
rect 9193 4302 9230 4303
rect 9250 4302 9335 4308
rect 9401 4332 9439 4340
rect 9512 4336 9548 4337
rect 9401 4312 9410 4332
rect 9430 4312 9439 4332
rect 9401 4303 9439 4312
rect 9463 4328 9548 4336
rect 9463 4308 9520 4328
rect 9540 4308 9548 4328
rect 9401 4302 9438 4303
rect 9463 4302 9548 4308
rect 9614 4332 9652 4340
rect 9614 4312 9623 4332
rect 9643 4312 9652 4332
rect 9614 4303 9652 4312
rect 9841 4333 9878 4343
rect 9841 4315 9851 4333
rect 9869 4315 9878 4333
rect 9841 4306 9878 4315
rect 10140 4314 10180 4362
rect 11306 4368 11344 4377
rect 11306 4348 11315 4368
rect 11335 4348 11344 4368
rect 11306 4340 11344 4348
rect 11410 4372 11495 4378
rect 11520 4377 11557 4378
rect 11410 4352 11418 4372
rect 11438 4352 11495 4372
rect 11410 4344 11495 4352
rect 11519 4368 11557 4377
rect 11519 4348 11528 4368
rect 11548 4348 11557 4368
rect 11410 4343 11446 4344
rect 11519 4340 11557 4348
rect 11623 4372 11708 4378
rect 11728 4377 11765 4378
rect 11623 4352 11631 4372
rect 11651 4371 11708 4372
rect 11651 4352 11680 4371
rect 11623 4351 11680 4352
rect 11701 4351 11708 4371
rect 11623 4344 11708 4351
rect 11727 4368 11765 4377
rect 11727 4348 11736 4368
rect 11756 4348 11765 4368
rect 11623 4343 11659 4344
rect 11727 4340 11765 4348
rect 11831 4372 11975 4378
rect 11831 4352 11839 4372
rect 11859 4355 11895 4372
rect 11915 4355 11947 4372
rect 11859 4352 11947 4355
rect 11967 4352 11975 4372
rect 11831 4344 11975 4352
rect 11831 4343 11867 4344
rect 11939 4343 11975 4344
rect 12041 4377 12078 4378
rect 12041 4376 12079 4377
rect 12041 4368 12105 4376
rect 12041 4348 12050 4368
rect 12070 4354 12105 4368
rect 12125 4354 12128 4374
rect 12070 4349 12128 4354
rect 12070 4348 12105 4349
rect 10451 4318 10561 4332
rect 10451 4315 10494 4318
rect 10140 4307 10265 4314
rect 10451 4310 10455 4315
rect 9843 4305 9877 4306
rect 9614 4302 9651 4303
rect 9037 4281 9073 4302
rect 9463 4281 9494 4302
rect 10140 4288 10232 4307
rect 10257 4288 10265 4307
rect 8870 4277 8970 4281
rect 8870 4273 8932 4277
rect 8870 4247 8877 4273
rect 8903 4251 8932 4273
rect 8958 4251 8970 4277
rect 8903 4247 8970 4251
rect 8870 4244 8970 4247
rect 9038 4244 9073 4281
rect 9135 4278 9494 4281
rect 9135 4273 9357 4278
rect 9135 4249 9148 4273
rect 9172 4254 9357 4273
rect 9381 4254 9494 4278
rect 9172 4249 9494 4254
rect 9135 4245 9494 4249
rect 9561 4273 9710 4281
rect 9561 4253 9572 4273
rect 9592 4253 9710 4273
rect 10140 4278 10265 4288
rect 10373 4288 10455 4310
rect 10484 4288 10494 4315
rect 10522 4291 10529 4318
rect 10558 4310 10561 4318
rect 11307 4311 11344 4340
rect 10558 4291 10623 4310
rect 11308 4309 11344 4311
rect 11520 4309 11557 4340
rect 11728 4313 11765 4340
rect 12041 4336 12105 4348
rect 10522 4288 10623 4291
rect 10373 4286 10623 4288
rect 10140 4258 10180 4278
rect 9561 4246 9710 4253
rect 10139 4249 10180 4258
rect 9561 4245 9602 4246
rect 8885 4192 8922 4193
rect 8981 4192 9018 4193
rect 9037 4192 9073 4244
rect 9092 4192 9129 4193
rect 8785 4183 8923 4192
rect 8380 4162 8491 4177
rect 8380 4160 8422 4162
rect 8050 4139 8155 4141
rect 7706 4131 7876 4132
rect 8050 4131 8099 4139
rect 7706 4112 8099 4131
rect 8130 4112 8155 4139
rect 8380 4140 8387 4160
rect 8406 4140 8422 4160
rect 8380 4132 8422 4140
rect 8450 4160 8491 4162
rect 8450 4140 8464 4160
rect 8483 4140 8491 4160
rect 8785 4163 8894 4183
rect 8914 4163 8923 4183
rect 8785 4156 8923 4163
rect 8981 4183 9129 4192
rect 8981 4163 8990 4183
rect 9010 4163 9100 4183
rect 9120 4163 9129 4183
rect 8785 4154 8881 4156
rect 8981 4153 9129 4163
rect 9188 4183 9225 4193
rect 9300 4192 9337 4193
rect 9281 4190 9337 4192
rect 9188 4163 9196 4183
rect 9216 4163 9225 4183
rect 9037 4152 9073 4153
rect 8450 4132 8491 4140
rect 8380 4126 8491 4132
rect 7706 4105 8155 4112
rect 7706 4103 7876 4105
rect 6556 4072 6666 4086
rect 6556 4069 6599 4072
rect 6556 4064 6560 4069
rect 6090 4034 6258 4036
rect 5814 4031 6258 4034
rect 5475 4007 5586 4013
rect 5475 3999 5516 4007
rect 5164 3944 5203 3988
rect 5475 3979 5483 3999
rect 5502 3979 5516 3999
rect 5475 3977 5516 3979
rect 5544 3999 5586 4007
rect 5544 3979 5560 3999
rect 5579 3979 5586 3999
rect 5544 3977 5586 3979
rect 5475 3962 5586 3977
rect 5812 4008 6258 4031
rect 5164 3920 5204 3944
rect 5504 3920 5551 3922
rect 5812 3920 5850 4008
rect 6090 4007 6258 4008
rect 6478 4042 6560 4064
rect 6589 4042 6599 4069
rect 6627 4045 6634 4072
rect 6663 4064 6666 4072
rect 6663 4045 6728 4064
rect 6627 4042 6728 4045
rect 6478 4040 6728 4042
rect 6478 3961 6515 4040
rect 6556 4027 6666 4040
rect 6630 3971 6661 3972
rect 6478 3941 6487 3961
rect 6507 3941 6515 3961
rect 6478 3931 6515 3941
rect 6574 3961 6661 3971
rect 6574 3941 6583 3961
rect 6603 3941 6661 3961
rect 6574 3932 6661 3941
rect 6574 3931 6611 3932
rect 5164 3887 5850 3920
rect 5164 3830 5203 3887
rect 5812 3885 5850 3887
rect 6630 3879 6661 3932
rect 6691 3961 6728 4040
rect 6899 4053 7292 4057
rect 6899 4036 6918 4053
rect 6938 4037 7292 4053
rect 7312 4037 7315 4057
rect 6938 4036 7315 4037
rect 6899 4032 7315 4036
rect 6899 4031 7240 4032
rect 6843 3971 6874 3972
rect 6691 3941 6700 3961
rect 6720 3941 6728 3961
rect 6691 3931 6728 3941
rect 6787 3964 6874 3971
rect 6787 3961 6848 3964
rect 6787 3941 6796 3961
rect 6816 3944 6848 3961
rect 6869 3944 6874 3964
rect 6816 3941 6874 3944
rect 6787 3934 6874 3941
rect 6899 3961 6936 4031
rect 7202 4030 7239 4031
rect 7051 3971 7087 3972
rect 6899 3941 6908 3961
rect 6928 3941 6936 3961
rect 6787 3932 6843 3934
rect 6787 3931 6824 3932
rect 6899 3931 6936 3941
rect 6995 3961 7143 3971
rect 7243 3968 7339 3970
rect 6995 3941 7004 3961
rect 7024 3941 7114 3961
rect 7134 3941 7143 3961
rect 6995 3932 7143 3941
rect 7201 3961 7339 3968
rect 7201 3941 7210 3961
rect 7230 3941 7339 3961
rect 7201 3932 7339 3941
rect 6995 3931 7032 3932
rect 7051 3880 7087 3932
rect 7106 3931 7143 3932
rect 7202 3931 7239 3932
rect 6522 3878 6563 3879
rect 6414 3871 6563 3878
rect 6414 3851 6532 3871
rect 6552 3851 6563 3871
rect 6414 3843 6563 3851
rect 6630 3875 6989 3879
rect 6630 3870 6952 3875
rect 6630 3846 6743 3870
rect 6767 3851 6952 3870
rect 6976 3851 6989 3875
rect 6767 3846 6989 3851
rect 6630 3843 6989 3846
rect 7051 3843 7086 3880
rect 7154 3877 7254 3880
rect 7154 3873 7221 3877
rect 7154 3847 7166 3873
rect 7192 3851 7221 3873
rect 7247 3851 7254 3877
rect 7192 3847 7254 3851
rect 7154 3843 7254 3847
rect 5164 3828 5212 3830
rect 5164 3810 5175 3828
rect 5193 3810 5212 3828
rect 6630 3822 6661 3843
rect 7051 3822 7087 3843
rect 6473 3821 6510 3822
rect 5164 3801 5212 3810
rect 5165 3800 5212 3801
rect 5478 3805 5588 3819
rect 5478 3802 5521 3805
rect 5478 3797 5482 3802
rect 5400 3775 5482 3797
rect 5511 3775 5521 3802
rect 5549 3778 5556 3805
rect 5585 3797 5588 3805
rect 6472 3812 6510 3821
rect 5585 3778 5650 3797
rect 6472 3792 6481 3812
rect 6501 3792 6510 3812
rect 5549 3775 5650 3778
rect 5400 3773 5650 3775
rect 5168 3737 5205 3738
rect 4786 3630 4796 3648
rect 4814 3630 4826 3648
rect 4786 3625 4826 3630
rect 5164 3734 5205 3737
rect 5164 3729 5206 3734
rect 5164 3711 5177 3729
rect 5195 3711 5206 3729
rect 5164 3697 5206 3711
rect 5244 3697 5291 3701
rect 5164 3691 5291 3697
rect 5164 3662 5252 3691
rect 5281 3662 5291 3691
rect 5400 3694 5437 3773
rect 5478 3760 5588 3773
rect 5552 3704 5583 3705
rect 5400 3674 5409 3694
rect 5429 3674 5437 3694
rect 5400 3664 5437 3674
rect 5496 3694 5583 3704
rect 5496 3674 5505 3694
rect 5525 3674 5583 3694
rect 5496 3665 5583 3674
rect 5496 3664 5533 3665
rect 5164 3658 5291 3662
rect 5164 3641 5203 3658
rect 5244 3657 5291 3658
rect 4786 3621 4823 3625
rect 5164 3623 5175 3641
rect 5193 3623 5203 3641
rect 5164 3614 5203 3623
rect 5165 3613 5202 3614
rect 5552 3612 5583 3665
rect 5613 3694 5650 3773
rect 5821 3770 6214 3790
rect 6234 3770 6237 3790
rect 6472 3784 6510 3792
rect 6576 3816 6661 3822
rect 6686 3821 6723 3822
rect 6576 3796 6584 3816
rect 6604 3796 6661 3816
rect 6576 3788 6661 3796
rect 6685 3812 6723 3821
rect 6685 3792 6694 3812
rect 6714 3792 6723 3812
rect 6576 3787 6612 3788
rect 6685 3784 6723 3792
rect 6789 3816 6874 3822
rect 6894 3821 6931 3822
rect 6789 3796 6797 3816
rect 6817 3815 6874 3816
rect 6817 3796 6846 3815
rect 6789 3795 6846 3796
rect 6867 3795 6874 3815
rect 6789 3788 6874 3795
rect 6893 3812 6931 3821
rect 6893 3792 6902 3812
rect 6922 3792 6931 3812
rect 6789 3787 6825 3788
rect 6893 3784 6931 3792
rect 6997 3816 7141 3822
rect 6997 3796 7005 3816
rect 7025 3814 7113 3816
rect 7025 3796 7054 3814
rect 6997 3793 7054 3796
rect 7081 3796 7113 3814
rect 7133 3796 7141 3816
rect 7081 3793 7141 3796
rect 6997 3788 7141 3793
rect 6997 3787 7033 3788
rect 7105 3787 7141 3788
rect 7207 3821 7244 3822
rect 7207 3820 7245 3821
rect 7207 3812 7271 3820
rect 7207 3792 7216 3812
rect 7236 3798 7271 3812
rect 7291 3798 7294 3818
rect 7236 3793 7294 3798
rect 7236 3792 7271 3793
rect 5821 3765 6237 3770
rect 5821 3764 6162 3765
rect 5765 3704 5796 3705
rect 5613 3674 5622 3694
rect 5642 3674 5650 3694
rect 5613 3664 5650 3674
rect 5709 3697 5796 3704
rect 5709 3694 5770 3697
rect 5709 3674 5718 3694
rect 5738 3677 5770 3694
rect 5791 3677 5796 3697
rect 5738 3674 5796 3677
rect 5709 3667 5796 3674
rect 5821 3694 5858 3764
rect 6124 3763 6161 3764
rect 6473 3755 6510 3784
rect 6474 3753 6510 3755
rect 6686 3753 6723 3784
rect 6474 3731 6723 3753
rect 6894 3752 6931 3784
rect 7207 3780 7271 3792
rect 7311 3754 7338 3932
rect 7706 3925 7735 4103
rect 7775 4065 7839 4077
rect 8115 4073 8152 4105
rect 8323 4104 8572 4126
rect 8323 4073 8360 4104
rect 8536 4102 8572 4104
rect 8536 4073 8573 4102
rect 8885 4093 8922 4094
rect 9188 4093 9225 4163
rect 9250 4183 9337 4190
rect 9250 4180 9308 4183
rect 9250 4160 9255 4180
rect 9276 4163 9308 4180
rect 9328 4163 9337 4183
rect 9276 4160 9337 4163
rect 9250 4153 9337 4160
rect 9396 4183 9433 4193
rect 9396 4163 9404 4183
rect 9424 4163 9433 4183
rect 9250 4152 9281 4153
rect 8884 4092 9225 4093
rect 8809 4087 9225 4092
rect 7775 4064 7810 4065
rect 7752 4059 7810 4064
rect 7752 4039 7755 4059
rect 7775 4045 7810 4059
rect 7830 4045 7839 4065
rect 7775 4037 7839 4045
rect 7801 4036 7839 4037
rect 7802 4035 7839 4036
rect 7905 4069 7941 4070
rect 8013 4069 8049 4070
rect 7905 4061 8049 4069
rect 7905 4041 7913 4061
rect 7933 4041 8021 4061
rect 8041 4041 8049 4061
rect 7905 4035 8049 4041
rect 8115 4065 8153 4073
rect 8221 4069 8257 4070
rect 8115 4045 8124 4065
rect 8144 4045 8153 4065
rect 8115 4036 8153 4045
rect 8172 4062 8257 4069
rect 8172 4042 8179 4062
rect 8200 4061 8257 4062
rect 8200 4042 8229 4061
rect 8172 4041 8229 4042
rect 8249 4041 8257 4061
rect 8115 4035 8152 4036
rect 8172 4035 8257 4041
rect 8323 4065 8361 4073
rect 8434 4069 8470 4070
rect 8323 4045 8332 4065
rect 8352 4045 8361 4065
rect 8323 4036 8361 4045
rect 8385 4061 8470 4069
rect 8385 4041 8442 4061
rect 8462 4041 8470 4061
rect 8323 4035 8360 4036
rect 8385 4035 8470 4041
rect 8536 4065 8574 4073
rect 8809 4067 8812 4087
rect 8832 4067 9225 4087
rect 9396 4084 9433 4163
rect 9463 4192 9494 4245
rect 9844 4243 9881 4244
rect 9843 4234 9882 4243
rect 9843 4216 9853 4234
rect 9871 4216 9882 4234
rect 10139 4231 10149 4249
rect 10167 4231 10180 4249
rect 10139 4222 10180 4231
rect 10139 4221 10176 4222
rect 9755 4199 9802 4200
rect 9843 4199 9882 4216
rect 9755 4195 9882 4199
rect 9513 4192 9550 4193
rect 9463 4183 9550 4192
rect 9463 4163 9521 4183
rect 9541 4163 9550 4183
rect 9463 4153 9550 4163
rect 9609 4183 9646 4193
rect 9609 4163 9617 4183
rect 9637 4163 9646 4183
rect 9463 4152 9494 4153
rect 9458 4084 9568 4097
rect 9609 4084 9646 4163
rect 9755 4166 9765 4195
rect 9794 4166 9882 4195
rect 10373 4207 10410 4286
rect 10451 4273 10561 4286
rect 10525 4217 10556 4218
rect 10373 4187 10382 4207
rect 10402 4187 10410 4207
rect 10373 4177 10410 4187
rect 10469 4207 10556 4217
rect 10469 4187 10478 4207
rect 10498 4187 10556 4207
rect 10469 4178 10556 4187
rect 10469 4177 10506 4178
rect 9755 4160 9882 4166
rect 9755 4156 9802 4160
rect 9840 4146 9882 4160
rect 10142 4155 10179 4159
rect 9840 4128 9851 4146
rect 9869 4128 9882 4146
rect 9840 4123 9882 4128
rect 9841 4120 9882 4123
rect 10139 4150 10179 4155
rect 10139 4132 10151 4150
rect 10169 4132 10179 4150
rect 9841 4119 9878 4120
rect 9396 4082 9646 4084
rect 9396 4079 9497 4082
rect 8536 4045 8545 4065
rect 8565 4045 8574 4065
rect 9396 4060 9461 4079
rect 8536 4036 8574 4045
rect 9458 4052 9461 4060
rect 9490 4052 9497 4079
rect 9525 4055 9535 4082
rect 9564 4060 9646 4082
rect 9564 4055 9568 4060
rect 9525 4052 9568 4055
rect 9458 4038 9568 4052
rect 9834 4056 9881 4057
rect 9834 4047 9882 4056
rect 8536 4035 8573 4036
rect 7959 4014 7995 4035
rect 8385 4014 8416 4035
rect 9834 4029 9853 4047
rect 9871 4029 9882 4047
rect 9834 4027 9882 4029
rect 7792 4010 7892 4014
rect 7792 4006 7854 4010
rect 7792 3980 7799 4006
rect 7825 3984 7854 4006
rect 7880 3984 7892 4010
rect 7825 3980 7892 3984
rect 7792 3977 7892 3980
rect 7960 3977 7995 4014
rect 8057 4011 8416 4014
rect 8057 4006 8279 4011
rect 8057 3982 8070 4006
rect 8094 3987 8279 4006
rect 8303 3987 8416 4011
rect 8094 3982 8416 3987
rect 8057 3978 8416 3982
rect 8483 4006 8632 4014
rect 8483 3986 8494 4006
rect 8514 3986 8632 4006
rect 8483 3979 8632 3986
rect 8483 3978 8524 3979
rect 7959 3938 7995 3977
rect 7807 3925 7844 3926
rect 7903 3925 7940 3926
rect 7959 3925 7966 3938
rect 7706 3916 7845 3925
rect 7706 3896 7816 3916
rect 7836 3896 7845 3916
rect 7706 3889 7845 3896
rect 7903 3916 7966 3925
rect 7903 3896 7912 3916
rect 7932 3900 7966 3916
rect 7989 3925 7995 3938
rect 8014 3925 8051 3926
rect 7989 3916 8051 3925
rect 7989 3900 8022 3916
rect 7932 3896 8022 3900
rect 8042 3896 8051 3916
rect 7706 3887 7803 3889
rect 7706 3886 7735 3887
rect 7903 3886 8051 3896
rect 8110 3916 8147 3926
rect 8222 3925 8259 3926
rect 8203 3923 8259 3925
rect 8110 3896 8118 3916
rect 8138 3896 8147 3916
rect 7959 3885 7995 3886
rect 7807 3826 7844 3827
rect 8110 3826 8147 3896
rect 8172 3916 8259 3923
rect 8172 3913 8230 3916
rect 8172 3893 8177 3913
rect 8198 3896 8230 3913
rect 8250 3896 8259 3916
rect 8198 3893 8259 3896
rect 8172 3886 8259 3893
rect 8318 3916 8355 3926
rect 8318 3896 8326 3916
rect 8346 3896 8355 3916
rect 8172 3885 8203 3886
rect 7806 3825 8147 3826
rect 7731 3821 8147 3825
rect 7731 3820 8108 3821
rect 7731 3800 7734 3820
rect 7754 3804 8108 3820
rect 8128 3804 8147 3821
rect 7754 3800 8147 3804
rect 8318 3817 8355 3896
rect 8385 3925 8416 3978
rect 9196 3970 9234 3972
rect 9843 3970 9882 4027
rect 9196 3937 9882 3970
rect 8435 3925 8472 3926
rect 8385 3916 8472 3925
rect 8385 3896 8443 3916
rect 8463 3896 8472 3916
rect 8385 3886 8472 3896
rect 8531 3916 8568 3926
rect 8531 3896 8539 3916
rect 8559 3896 8568 3916
rect 8385 3885 8416 3886
rect 8380 3817 8490 3830
rect 8531 3817 8568 3896
rect 8318 3815 8568 3817
rect 8318 3812 8419 3815
rect 8318 3793 8383 3812
rect 8380 3785 8383 3793
rect 8412 3785 8419 3812
rect 8447 3788 8457 3815
rect 8486 3793 8568 3815
rect 8788 3849 8956 3850
rect 9196 3849 9234 3937
rect 9495 3935 9542 3937
rect 9842 3913 9882 3937
rect 8788 3826 9234 3849
rect 9460 3880 9571 3895
rect 9460 3878 9502 3880
rect 9460 3858 9467 3878
rect 9486 3858 9502 3878
rect 9460 3850 9502 3858
rect 9530 3878 9571 3880
rect 9530 3858 9544 3878
rect 9563 3858 9571 3878
rect 9843 3869 9882 3913
rect 9530 3850 9571 3858
rect 9460 3844 9571 3850
rect 8788 3823 9232 3826
rect 8788 3821 8956 3823
rect 8486 3788 8490 3793
rect 8447 3785 8490 3788
rect 8380 3771 8490 3785
rect 7170 3752 7338 3754
rect 6891 3745 7338 3752
rect 6555 3725 6666 3731
rect 6555 3717 6596 3725
rect 5973 3704 6009 3705
rect 5821 3674 5830 3694
rect 5850 3674 5858 3694
rect 5709 3665 5765 3667
rect 5709 3664 5746 3665
rect 5821 3664 5858 3674
rect 5917 3694 6065 3704
rect 6165 3701 6261 3703
rect 5917 3674 5926 3694
rect 5946 3674 6036 3694
rect 6056 3674 6065 3694
rect 5917 3665 6065 3674
rect 6123 3694 6261 3701
rect 6123 3674 6132 3694
rect 6152 3674 6261 3694
rect 6555 3697 6563 3717
rect 6582 3697 6596 3717
rect 6555 3695 6596 3697
rect 6624 3717 6666 3725
rect 6624 3697 6640 3717
rect 6659 3697 6666 3717
rect 6891 3718 6916 3745
rect 6947 3726 7338 3745
rect 6947 3718 6996 3726
rect 7170 3725 7338 3726
rect 6891 3716 6996 3718
rect 6624 3695 6666 3697
rect 6555 3680 6666 3695
rect 6123 3665 6261 3674
rect 5917 3664 5954 3665
rect 5973 3613 6009 3665
rect 6028 3664 6065 3665
rect 6124 3664 6161 3665
rect 5444 3611 5485 3612
rect 5336 3604 5485 3611
rect 4459 3602 4496 3603
rect 4409 3593 4496 3602
rect 4409 3573 4467 3593
rect 4487 3573 4496 3593
rect 4409 3563 4496 3573
rect 4555 3593 4592 3603
rect 4555 3573 4563 3593
rect 4583 3573 4592 3593
rect 5336 3584 5454 3604
rect 5474 3584 5485 3604
rect 5336 3576 5485 3584
rect 5552 3608 5911 3612
rect 5552 3603 5874 3608
rect 5552 3579 5665 3603
rect 5689 3584 5874 3603
rect 5898 3584 5911 3608
rect 5689 3579 5911 3584
rect 5552 3576 5911 3579
rect 5973 3576 6008 3613
rect 6076 3610 6176 3613
rect 6076 3606 6143 3610
rect 6076 3580 6088 3606
rect 6114 3584 6143 3606
rect 6169 3584 6176 3610
rect 6114 3580 6176 3584
rect 6076 3576 6176 3580
rect 4409 3562 4440 3563
rect 4404 3494 4514 3507
rect 4555 3494 4592 3573
rect 4789 3558 4826 3559
rect 4785 3549 4826 3558
rect 5552 3555 5583 3576
rect 5973 3555 6009 3576
rect 5395 3554 5432 3555
rect 5169 3551 5203 3552
rect 4785 3531 4798 3549
rect 4816 3531 4826 3549
rect 4785 3522 4826 3531
rect 5168 3542 5205 3551
rect 5168 3524 5177 3542
rect 5195 3524 5205 3542
rect 4785 3502 4825 3522
rect 5168 3514 5205 3524
rect 5394 3545 5432 3554
rect 5394 3525 5403 3545
rect 5423 3525 5432 3545
rect 5394 3517 5432 3525
rect 5498 3549 5583 3555
rect 5608 3554 5645 3555
rect 5498 3529 5506 3549
rect 5526 3529 5583 3549
rect 5498 3521 5583 3529
rect 5607 3545 5645 3554
rect 5607 3525 5616 3545
rect 5636 3525 5645 3545
rect 5498 3520 5534 3521
rect 5607 3517 5645 3525
rect 5711 3549 5796 3555
rect 5816 3554 5853 3555
rect 5711 3529 5719 3549
rect 5739 3548 5796 3549
rect 5739 3529 5768 3548
rect 5711 3528 5768 3529
rect 5789 3528 5796 3548
rect 5711 3521 5796 3528
rect 5815 3545 5853 3554
rect 5815 3525 5824 3545
rect 5844 3525 5853 3545
rect 5711 3520 5747 3521
rect 5815 3517 5853 3525
rect 5919 3549 6063 3555
rect 5919 3529 5927 3549
rect 5947 3548 6035 3549
rect 5947 3529 5978 3548
rect 5919 3528 5978 3529
rect 6003 3529 6035 3548
rect 6055 3529 6063 3549
rect 6003 3528 6063 3529
rect 5919 3521 6063 3528
rect 5919 3520 5955 3521
rect 6027 3520 6063 3521
rect 6129 3554 6166 3555
rect 6129 3553 6167 3554
rect 6129 3545 6193 3553
rect 6129 3525 6138 3545
rect 6158 3531 6193 3545
rect 6213 3531 6216 3551
rect 6158 3526 6216 3531
rect 6158 3525 6193 3526
rect 4342 3492 4592 3494
rect 4342 3489 4443 3492
rect 2860 3432 2924 3444
rect 3200 3440 3237 3467
rect 3408 3440 3445 3471
rect 3621 3469 3657 3471
rect 4342 3470 4407 3489
rect 3621 3440 3658 3469
rect 4404 3462 4407 3470
rect 4436 3462 4443 3489
rect 4471 3465 4481 3492
rect 4510 3470 4592 3492
rect 4700 3492 4825 3502
rect 4700 3473 4708 3492
rect 4733 3473 4825 3492
rect 4510 3465 4514 3470
rect 4700 3466 4825 3473
rect 4471 3462 4514 3465
rect 4404 3448 4514 3462
rect 2860 3431 2895 3432
rect 2837 3426 2895 3431
rect 2837 3406 2840 3426
rect 2860 3412 2895 3426
rect 2915 3412 2924 3432
rect 2860 3404 2924 3412
rect 2886 3403 2924 3404
rect 2887 3402 2924 3403
rect 2990 3436 3026 3437
rect 3098 3436 3134 3437
rect 2990 3428 3134 3436
rect 2990 3408 2998 3428
rect 3018 3425 3106 3428
rect 3018 3408 3050 3425
rect 3070 3408 3106 3425
rect 3126 3408 3134 3428
rect 2990 3402 3134 3408
rect 3200 3432 3238 3440
rect 3306 3436 3342 3437
rect 3200 3412 3209 3432
rect 3229 3412 3238 3432
rect 3200 3403 3238 3412
rect 3257 3429 3342 3436
rect 3257 3409 3264 3429
rect 3285 3428 3342 3429
rect 3285 3409 3314 3428
rect 3257 3408 3314 3409
rect 3334 3408 3342 3428
rect 3200 3402 3237 3403
rect 3257 3402 3342 3408
rect 3408 3432 3446 3440
rect 3519 3436 3555 3437
rect 3408 3412 3417 3432
rect 3437 3412 3446 3432
rect 3408 3403 3446 3412
rect 3470 3428 3555 3436
rect 3470 3408 3527 3428
rect 3547 3408 3555 3428
rect 3408 3402 3445 3403
rect 3470 3402 3555 3408
rect 3621 3432 3659 3440
rect 3621 3412 3630 3432
rect 3650 3412 3659 3432
rect 3621 3403 3659 3412
rect 4785 3418 4825 3466
rect 5169 3486 5203 3514
rect 5395 3488 5432 3517
rect 5396 3486 5432 3488
rect 5608 3486 5645 3517
rect 5169 3485 5341 3486
rect 5169 3453 5355 3485
rect 5396 3464 5645 3486
rect 5816 3485 5853 3517
rect 6129 3513 6193 3525
rect 6233 3487 6260 3665
rect 8788 3643 8815 3821
rect 8855 3783 8919 3795
rect 9195 3791 9232 3823
rect 9403 3822 9652 3844
rect 9403 3791 9440 3822
rect 9616 3820 9652 3822
rect 9616 3791 9653 3820
rect 8855 3782 8890 3783
rect 8832 3777 8890 3782
rect 8832 3757 8835 3777
rect 8855 3763 8890 3777
rect 8910 3763 8919 3783
rect 8855 3755 8919 3763
rect 8881 3754 8919 3755
rect 8882 3753 8919 3754
rect 8985 3787 9021 3788
rect 9093 3787 9129 3788
rect 8985 3782 9129 3787
rect 8985 3779 9047 3782
rect 8985 3759 8993 3779
rect 9013 3762 9047 3779
rect 9070 3779 9129 3782
rect 9070 3762 9101 3779
rect 9013 3759 9101 3762
rect 9121 3759 9129 3779
rect 8985 3753 9129 3759
rect 9195 3783 9233 3791
rect 9301 3787 9337 3788
rect 9195 3763 9204 3783
rect 9224 3763 9233 3783
rect 9195 3754 9233 3763
rect 9252 3780 9337 3787
rect 9252 3760 9259 3780
rect 9280 3779 9337 3780
rect 9280 3760 9309 3779
rect 9252 3759 9309 3760
rect 9329 3759 9337 3779
rect 9195 3753 9232 3754
rect 9252 3753 9337 3759
rect 9403 3783 9441 3791
rect 9514 3787 9550 3788
rect 9403 3763 9412 3783
rect 9432 3763 9441 3783
rect 9403 3754 9441 3763
rect 9465 3779 9550 3787
rect 9465 3759 9522 3779
rect 9542 3759 9550 3779
rect 9403 3753 9440 3754
rect 9465 3753 9550 3759
rect 9616 3783 9654 3791
rect 9616 3763 9625 3783
rect 9645 3763 9654 3783
rect 9616 3754 9654 3763
rect 9616 3753 9653 3754
rect 9039 3732 9075 3753
rect 9465 3732 9496 3753
rect 8872 3728 8972 3732
rect 8872 3724 8934 3728
rect 8872 3698 8879 3724
rect 8905 3702 8934 3724
rect 8960 3702 8972 3728
rect 8905 3698 8972 3702
rect 8872 3695 8972 3698
rect 9040 3695 9075 3732
rect 9137 3729 9496 3732
rect 9137 3724 9359 3729
rect 9137 3700 9150 3724
rect 9174 3705 9359 3724
rect 9383 3705 9496 3729
rect 9174 3700 9496 3705
rect 9137 3696 9496 3700
rect 9563 3724 9712 3732
rect 9563 3704 9574 3724
rect 9594 3704 9712 3724
rect 9563 3697 9712 3704
rect 9563 3696 9604 3697
rect 8887 3643 8924 3644
rect 8983 3643 9020 3644
rect 9039 3643 9075 3695
rect 9094 3643 9131 3644
rect 8787 3634 8925 3643
rect 8787 3614 8896 3634
rect 8916 3614 8925 3634
rect 8787 3607 8925 3614
rect 8983 3634 9131 3643
rect 8983 3614 8992 3634
rect 9012 3614 9102 3634
rect 9122 3614 9131 3634
rect 8787 3605 8883 3607
rect 8983 3604 9131 3614
rect 9190 3634 9227 3644
rect 9302 3643 9339 3644
rect 9283 3641 9339 3643
rect 9190 3614 9198 3634
rect 9218 3614 9227 3634
rect 9039 3603 9075 3604
rect 6416 3561 6526 3575
rect 6416 3558 6459 3561
rect 6416 3553 6420 3558
rect 6092 3485 6260 3487
rect 5816 3479 6260 3485
rect 5169 3421 5203 3453
rect 3621 3402 3658 3403
rect 3044 3381 3080 3402
rect 3470 3381 3501 3402
rect 4785 3400 4796 3418
rect 4814 3400 4825 3418
rect 4785 3392 4825 3400
rect 5165 3412 5203 3421
rect 5165 3394 5175 3412
rect 5193 3394 5203 3412
rect 4786 3391 4823 3392
rect 5165 3388 5203 3394
rect 5321 3390 5355 3453
rect 5477 3458 5588 3464
rect 5477 3450 5518 3458
rect 5477 3430 5485 3450
rect 5504 3430 5518 3450
rect 5477 3428 5518 3430
rect 5546 3450 5588 3458
rect 5546 3430 5562 3450
rect 5581 3430 5588 3450
rect 5546 3428 5588 3430
rect 5477 3413 5588 3428
rect 5815 3459 6260 3479
rect 5815 3390 5853 3459
rect 6092 3458 6260 3459
rect 6338 3531 6420 3553
rect 6449 3531 6459 3558
rect 6487 3534 6494 3561
rect 6523 3553 6526 3561
rect 8521 3570 8632 3585
rect 8521 3568 8563 3570
rect 6523 3534 6588 3553
rect 6487 3531 6588 3534
rect 6338 3529 6588 3531
rect 6338 3450 6375 3529
rect 6416 3516 6526 3529
rect 6490 3460 6521 3461
rect 6338 3430 6347 3450
rect 6367 3430 6375 3450
rect 6338 3420 6375 3430
rect 6434 3450 6521 3460
rect 6434 3430 6443 3450
rect 6463 3430 6521 3450
rect 6434 3421 6521 3430
rect 6434 3420 6471 3421
rect 5165 3384 5202 3388
rect 2877 3377 2977 3381
rect 2877 3373 2939 3377
rect 2877 3347 2884 3373
rect 2910 3351 2939 3373
rect 2965 3351 2977 3377
rect 2910 3347 2977 3351
rect 2877 3344 2977 3347
rect 3045 3344 3080 3381
rect 3142 3378 3501 3381
rect 3142 3373 3364 3378
rect 3142 3349 3155 3373
rect 3179 3354 3364 3373
rect 3388 3354 3501 3378
rect 3179 3349 3501 3354
rect 3142 3345 3501 3349
rect 3568 3373 3717 3381
rect 5321 3379 5853 3390
rect 3568 3353 3579 3373
rect 3599 3353 3717 3373
rect 5320 3363 5853 3379
rect 6490 3368 6521 3421
rect 6551 3450 6588 3529
rect 6759 3539 7152 3546
rect 6759 3522 6767 3539
rect 6799 3526 7152 3539
rect 7172 3526 7175 3546
rect 8254 3541 8295 3550
rect 6799 3522 7175 3526
rect 6759 3521 7175 3522
rect 7849 3539 8017 3540
rect 8254 3539 8263 3541
rect 6759 3520 7100 3521
rect 6703 3460 6734 3461
rect 6551 3430 6560 3450
rect 6580 3430 6588 3450
rect 6551 3420 6588 3430
rect 6647 3453 6734 3460
rect 6647 3450 6708 3453
rect 6647 3430 6656 3450
rect 6676 3433 6708 3450
rect 6729 3433 6734 3453
rect 6676 3430 6734 3433
rect 6647 3423 6734 3430
rect 6759 3450 6796 3520
rect 7062 3519 7099 3520
rect 7849 3519 8263 3539
rect 8289 3519 8295 3541
rect 8521 3548 8528 3568
rect 8547 3548 8563 3568
rect 8521 3540 8563 3548
rect 8591 3568 8632 3570
rect 8591 3548 8605 3568
rect 8624 3548 8632 3568
rect 8591 3540 8632 3548
rect 8887 3544 8924 3545
rect 9190 3544 9227 3614
rect 9252 3634 9339 3641
rect 9252 3631 9310 3634
rect 9252 3611 9257 3631
rect 9278 3614 9310 3631
rect 9330 3614 9339 3634
rect 9278 3611 9339 3614
rect 9252 3604 9339 3611
rect 9398 3634 9435 3644
rect 9398 3614 9406 3634
rect 9426 3614 9435 3634
rect 9252 3603 9283 3604
rect 8886 3543 9227 3544
rect 8521 3534 8632 3540
rect 8811 3538 9227 3543
rect 7849 3513 8295 3519
rect 7849 3511 8017 3513
rect 6911 3460 6947 3461
rect 6759 3430 6768 3450
rect 6788 3430 6796 3450
rect 6647 3421 6703 3423
rect 6647 3420 6684 3421
rect 6759 3420 6796 3430
rect 6855 3450 7003 3460
rect 7103 3457 7199 3459
rect 6855 3430 6864 3450
rect 6884 3445 6974 3450
rect 6884 3430 6919 3445
rect 6855 3421 6919 3430
rect 6855 3420 6892 3421
rect 6911 3404 6919 3421
rect 6940 3430 6974 3445
rect 6994 3430 7003 3450
rect 6940 3421 7003 3430
rect 7061 3450 7199 3457
rect 7061 3430 7070 3450
rect 7090 3430 7199 3450
rect 7061 3421 7199 3430
rect 6940 3404 6947 3421
rect 6966 3420 7003 3421
rect 7062 3420 7099 3421
rect 6911 3369 6947 3404
rect 6382 3367 6423 3368
rect 5320 3362 5834 3363
rect 3568 3346 3717 3353
rect 6274 3360 6423 3367
rect 4157 3350 4671 3351
rect 3568 3345 3609 3346
rect 2892 3292 2929 3293
rect 2988 3292 3025 3293
rect 3044 3292 3080 3344
rect 3099 3292 3136 3293
rect 2792 3283 2930 3292
rect 2792 3263 2901 3283
rect 2921 3263 2930 3283
rect 2792 3256 2930 3263
rect 2988 3283 3136 3292
rect 2988 3263 2997 3283
rect 3017 3263 3107 3283
rect 3127 3263 3136 3283
rect 2792 3254 2888 3256
rect 2988 3253 3136 3263
rect 3195 3283 3232 3293
rect 3307 3292 3344 3293
rect 3288 3290 3344 3292
rect 3195 3263 3203 3283
rect 3223 3263 3232 3283
rect 3044 3252 3080 3253
rect 1974 3200 2142 3202
rect 1696 3194 2142 3200
rect 764 3170 1180 3175
rect 1359 3173 1470 3179
rect 764 3169 1105 3170
rect 708 3109 739 3110
rect 556 3079 565 3099
rect 585 3079 593 3099
rect 556 3069 593 3079
rect 652 3102 739 3109
rect 652 3099 713 3102
rect 652 3079 661 3099
rect 681 3082 713 3099
rect 734 3082 739 3102
rect 681 3079 739 3082
rect 652 3072 739 3079
rect 764 3099 801 3169
rect 1067 3168 1104 3169
rect 1359 3165 1400 3173
rect 1359 3145 1367 3165
rect 1386 3145 1400 3165
rect 1359 3143 1400 3145
rect 1428 3165 1470 3173
rect 1428 3145 1444 3165
rect 1463 3145 1470 3165
rect 1696 3172 1702 3194
rect 1728 3174 2142 3194
rect 2892 3193 2929 3194
rect 3195 3193 3232 3263
rect 3257 3283 3344 3290
rect 3257 3280 3315 3283
rect 3257 3260 3262 3280
rect 3283 3263 3315 3280
rect 3335 3263 3344 3283
rect 3283 3260 3344 3263
rect 3257 3253 3344 3260
rect 3403 3283 3440 3293
rect 3403 3263 3411 3283
rect 3431 3263 3440 3283
rect 3257 3252 3288 3253
rect 2891 3192 3232 3193
rect 1728 3172 1737 3174
rect 1974 3173 2142 3174
rect 2816 3187 3232 3192
rect 1696 3163 1737 3172
rect 2816 3167 2819 3187
rect 2839 3167 3232 3187
rect 3403 3184 3440 3263
rect 3470 3292 3501 3345
rect 4138 3334 4671 3350
rect 6274 3340 6392 3360
rect 6412 3340 6423 3360
rect 4138 3323 4670 3334
rect 6274 3332 6423 3340
rect 6490 3364 6849 3368
rect 6490 3359 6812 3364
rect 6490 3335 6603 3359
rect 6627 3340 6812 3359
rect 6836 3340 6849 3364
rect 6627 3335 6849 3340
rect 6490 3332 6849 3335
rect 6911 3332 6946 3369
rect 7014 3366 7114 3369
rect 7014 3362 7081 3366
rect 7014 3336 7026 3362
rect 7052 3340 7081 3362
rect 7107 3340 7114 3366
rect 7052 3336 7114 3340
rect 7014 3332 7114 3336
rect 4789 3325 4826 3329
rect 3520 3292 3557 3293
rect 3470 3283 3557 3292
rect 3470 3263 3528 3283
rect 3548 3263 3557 3283
rect 3470 3253 3557 3263
rect 3616 3283 3653 3293
rect 3616 3263 3624 3283
rect 3644 3263 3653 3283
rect 3470 3252 3501 3253
rect 3465 3184 3575 3197
rect 3616 3184 3653 3263
rect 3403 3182 3653 3184
rect 3403 3179 3504 3182
rect 3403 3160 3468 3179
rect 1428 3143 1470 3145
rect 1359 3128 1470 3143
rect 3465 3152 3468 3160
rect 3497 3152 3504 3179
rect 3532 3155 3542 3182
rect 3571 3160 3653 3182
rect 3731 3254 3899 3255
rect 4138 3254 4176 3323
rect 3731 3234 4176 3254
rect 4403 3285 4514 3300
rect 4403 3283 4445 3285
rect 4403 3263 4410 3283
rect 4429 3263 4445 3283
rect 4403 3255 4445 3263
rect 4473 3283 4514 3285
rect 4473 3263 4487 3283
rect 4506 3263 4514 3283
rect 4473 3255 4514 3263
rect 4403 3249 4514 3255
rect 4636 3260 4670 3323
rect 4788 3319 4826 3325
rect 5168 3321 5205 3322
rect 4788 3301 4798 3319
rect 4816 3301 4826 3319
rect 4788 3292 4826 3301
rect 5166 3313 5206 3321
rect 5166 3295 5177 3313
rect 5195 3295 5206 3313
rect 6490 3311 6521 3332
rect 6911 3311 6947 3332
rect 6333 3310 6370 3311
rect 4788 3260 4822 3292
rect 3731 3228 4175 3234
rect 3731 3226 3899 3228
rect 3571 3155 3575 3160
rect 3532 3152 3575 3155
rect 3465 3138 3575 3152
rect 2694 3124 2762 3133
rect 916 3109 952 3110
rect 764 3079 773 3099
rect 793 3079 801 3099
rect 652 3070 708 3072
rect 652 3069 689 3070
rect 764 3069 801 3079
rect 860 3099 1008 3109
rect 1108 3106 1204 3108
rect 860 3079 869 3099
rect 889 3079 979 3099
rect 999 3079 1008 3099
rect 860 3070 1008 3079
rect 1066 3099 1204 3106
rect 1066 3079 1075 3099
rect 1095 3079 1204 3099
rect 2694 3095 2709 3124
rect 2757 3104 2762 3124
rect 2757 3095 2764 3104
rect 2694 3084 2764 3095
rect 1066 3070 1204 3079
rect 860 3069 897 3070
rect 916 3018 952 3070
rect 971 3069 1008 3070
rect 1067 3069 1104 3070
rect 387 3016 428 3017
rect 279 3009 428 3016
rect 279 2989 397 3009
rect 417 2989 428 3009
rect 279 2981 428 2989
rect 495 3013 854 3017
rect 495 3008 817 3013
rect 495 2984 608 3008
rect 632 2989 817 3008
rect 841 2989 854 3013
rect 632 2984 854 2989
rect 495 2981 854 2984
rect 916 2981 951 3018
rect 1019 3015 1119 3018
rect 1019 3011 1086 3015
rect 1019 2985 1031 3011
rect 1057 2989 1086 3011
rect 1112 2989 1119 3015
rect 1057 2985 1119 2989
rect 1019 2981 1119 2985
rect 495 2960 526 2981
rect 916 2960 952 2981
rect 338 2959 375 2960
rect 337 2950 375 2959
rect 337 2930 346 2950
rect 366 2930 375 2950
rect 337 2922 375 2930
rect 441 2954 526 2960
rect 551 2959 588 2960
rect 441 2934 449 2954
rect 469 2934 526 2954
rect 441 2926 526 2934
rect 550 2950 588 2959
rect 550 2930 559 2950
rect 579 2930 588 2950
rect 441 2925 477 2926
rect 550 2922 588 2930
rect 654 2954 739 2960
rect 759 2959 796 2960
rect 654 2934 662 2954
rect 682 2953 739 2954
rect 682 2934 711 2953
rect 654 2933 711 2934
rect 732 2933 739 2953
rect 654 2926 739 2933
rect 758 2950 796 2959
rect 758 2930 767 2950
rect 787 2930 796 2950
rect 654 2925 690 2926
rect 758 2922 796 2930
rect 862 2954 1006 2960
rect 862 2934 870 2954
rect 890 2951 978 2954
rect 890 2934 921 2951
rect 862 2931 921 2934
rect 944 2934 978 2951
rect 998 2934 1006 2954
rect 944 2931 1006 2934
rect 862 2926 1006 2931
rect 862 2925 898 2926
rect 970 2925 1006 2926
rect 1072 2959 1109 2960
rect 1072 2958 1110 2959
rect 1072 2950 1136 2958
rect 1072 2930 1081 2950
rect 1101 2936 1136 2950
rect 1156 2936 1159 2956
rect 1101 2931 1159 2936
rect 1101 2930 1136 2931
rect 338 2893 375 2922
rect 339 2891 375 2893
rect 551 2891 588 2922
rect 339 2869 588 2891
rect 759 2890 796 2922
rect 1072 2918 1136 2930
rect 1176 2892 1203 3070
rect 2703 2977 2764 3084
rect 3731 3048 3758 3226
rect 3798 3188 3862 3200
rect 4138 3196 4175 3228
rect 4346 3227 4595 3249
rect 4636 3228 4822 3260
rect 4650 3227 4822 3228
rect 4346 3196 4383 3227
rect 4559 3225 4595 3227
rect 4559 3196 4596 3225
rect 4788 3199 4822 3227
rect 5166 3247 5206 3295
rect 6332 3301 6370 3310
rect 6332 3281 6341 3301
rect 6361 3281 6370 3301
rect 6332 3273 6370 3281
rect 6436 3305 6521 3311
rect 6546 3310 6583 3311
rect 6436 3285 6444 3305
rect 6464 3285 6521 3305
rect 6436 3277 6521 3285
rect 6545 3301 6583 3310
rect 6545 3281 6554 3301
rect 6574 3281 6583 3301
rect 6436 3276 6472 3277
rect 6545 3273 6583 3281
rect 6649 3305 6734 3311
rect 6754 3310 6791 3311
rect 6649 3285 6657 3305
rect 6677 3304 6734 3305
rect 6677 3285 6706 3304
rect 6649 3284 6706 3285
rect 6727 3284 6734 3304
rect 6649 3277 6734 3284
rect 6753 3301 6791 3310
rect 6753 3281 6762 3301
rect 6782 3281 6791 3301
rect 6649 3276 6685 3277
rect 6753 3273 6791 3281
rect 6857 3305 7001 3311
rect 6857 3285 6865 3305
rect 6885 3285 6973 3305
rect 6993 3285 7001 3305
rect 6857 3277 7001 3285
rect 6857 3276 6893 3277
rect 6965 3276 7001 3277
rect 7067 3310 7104 3311
rect 7067 3309 7105 3310
rect 7067 3301 7131 3309
rect 7067 3281 7076 3301
rect 7096 3287 7131 3301
rect 7151 3287 7154 3307
rect 7096 3282 7154 3287
rect 7096 3281 7131 3282
rect 5477 3251 5587 3265
rect 5477 3248 5520 3251
rect 5166 3240 5291 3247
rect 5477 3243 5481 3248
rect 5166 3221 5258 3240
rect 5283 3221 5291 3240
rect 5166 3211 5291 3221
rect 5399 3221 5481 3243
rect 5510 3221 5520 3248
rect 5548 3224 5555 3251
rect 5584 3243 5587 3251
rect 6333 3244 6370 3273
rect 5584 3224 5649 3243
rect 6334 3242 6370 3244
rect 6546 3242 6583 3273
rect 6754 3246 6791 3273
rect 7067 3269 7131 3281
rect 5548 3221 5649 3224
rect 5399 3219 5649 3221
rect 3798 3187 3833 3188
rect 3775 3182 3833 3187
rect 3775 3162 3778 3182
rect 3798 3168 3833 3182
rect 3853 3168 3862 3188
rect 3798 3160 3862 3168
rect 3824 3159 3862 3160
rect 3825 3158 3862 3159
rect 3928 3192 3964 3193
rect 4036 3192 4072 3193
rect 3928 3185 4072 3192
rect 3928 3184 3988 3185
rect 3928 3164 3936 3184
rect 3956 3165 3988 3184
rect 4013 3184 4072 3185
rect 4013 3165 4044 3184
rect 3956 3164 4044 3165
rect 4064 3164 4072 3184
rect 3928 3158 4072 3164
rect 4138 3188 4176 3196
rect 4244 3192 4280 3193
rect 4138 3168 4147 3188
rect 4167 3168 4176 3188
rect 4138 3159 4176 3168
rect 4195 3185 4280 3192
rect 4195 3165 4202 3185
rect 4223 3184 4280 3185
rect 4223 3165 4252 3184
rect 4195 3164 4252 3165
rect 4272 3164 4280 3184
rect 4138 3158 4175 3159
rect 4195 3158 4280 3164
rect 4346 3188 4384 3196
rect 4457 3192 4493 3193
rect 4346 3168 4355 3188
rect 4375 3168 4384 3188
rect 4346 3159 4384 3168
rect 4408 3184 4493 3192
rect 4408 3164 4465 3184
rect 4485 3164 4493 3184
rect 4346 3158 4383 3159
rect 4408 3158 4493 3164
rect 4559 3188 4597 3196
rect 4559 3168 4568 3188
rect 4588 3168 4597 3188
rect 4559 3159 4597 3168
rect 4786 3189 4823 3199
rect 5166 3191 5206 3211
rect 4786 3171 4796 3189
rect 4814 3171 4823 3189
rect 4786 3162 4823 3171
rect 5165 3182 5206 3191
rect 5165 3164 5175 3182
rect 5193 3164 5206 3182
rect 4788 3161 4822 3162
rect 4559 3158 4596 3159
rect 3982 3137 4018 3158
rect 4408 3137 4439 3158
rect 5165 3155 5206 3164
rect 5165 3154 5202 3155
rect 5399 3140 5436 3219
rect 5477 3206 5587 3219
rect 5551 3150 5582 3151
rect 3815 3133 3915 3137
rect 3815 3129 3877 3133
rect 3815 3103 3822 3129
rect 3848 3107 3877 3129
rect 3903 3107 3915 3133
rect 3848 3103 3915 3107
rect 3815 3100 3915 3103
rect 3983 3100 4018 3137
rect 4080 3134 4439 3137
rect 4080 3129 4302 3134
rect 4080 3105 4093 3129
rect 4117 3110 4302 3129
rect 4326 3110 4439 3134
rect 4117 3105 4439 3110
rect 4080 3101 4439 3105
rect 4506 3129 4655 3137
rect 4506 3109 4517 3129
rect 4537 3109 4655 3129
rect 5399 3120 5408 3140
rect 5428 3120 5436 3140
rect 5399 3110 5436 3120
rect 5495 3140 5582 3150
rect 5495 3120 5504 3140
rect 5524 3120 5582 3140
rect 5495 3111 5582 3120
rect 5495 3110 5532 3111
rect 4506 3102 4655 3109
rect 4506 3101 4547 3102
rect 3830 3048 3867 3049
rect 3926 3048 3963 3049
rect 3982 3048 4018 3100
rect 4037 3048 4074 3049
rect 3730 3039 3868 3048
rect 2694 2976 2764 2977
rect 3355 3005 3466 3020
rect 3730 3019 3839 3039
rect 3859 3019 3868 3039
rect 3730 3012 3868 3019
rect 3926 3039 4074 3048
rect 3926 3019 3935 3039
rect 3955 3019 4045 3039
rect 4065 3019 4074 3039
rect 3730 3010 3826 3012
rect 3926 3009 4074 3019
rect 4133 3039 4170 3049
rect 4245 3048 4282 3049
rect 4226 3046 4282 3048
rect 4133 3019 4141 3039
rect 4161 3019 4170 3039
rect 3982 3008 4018 3009
rect 3355 3003 3397 3005
rect 3355 2983 3362 3003
rect 3381 2983 3397 3003
rect 2694 2975 2802 2976
rect 3355 2975 3397 2983
rect 3425 3003 3466 3005
rect 3425 2983 3439 3003
rect 3458 2983 3466 3003
rect 3425 2975 3466 2983
rect 2683 2974 2851 2975
rect 1470 2941 1580 2955
rect 1470 2938 1513 2941
rect 1470 2933 1474 2938
rect 1035 2890 1203 2892
rect 759 2887 1203 2890
rect 420 2863 531 2869
rect 420 2855 461 2863
rect 109 2800 148 2844
rect 420 2835 428 2855
rect 447 2835 461 2855
rect 420 2833 461 2835
rect 489 2855 531 2863
rect 489 2835 505 2855
rect 524 2835 531 2855
rect 489 2833 531 2835
rect 420 2819 531 2833
rect 757 2864 1203 2887
rect 109 2776 149 2800
rect 449 2776 496 2778
rect 757 2776 795 2864
rect 1035 2863 1203 2864
rect 1392 2911 1474 2933
rect 1503 2911 1513 2938
rect 1541 2914 1548 2941
rect 1577 2933 1580 2941
rect 2683 2948 3127 2974
rect 3355 2969 3466 2975
rect 2683 2946 2851 2948
rect 2683 2944 2802 2946
rect 1577 2914 1642 2933
rect 1541 2911 1642 2914
rect 1392 2909 1642 2911
rect 1392 2830 1429 2909
rect 1470 2896 1580 2909
rect 1544 2840 1575 2841
rect 1392 2810 1401 2830
rect 1421 2810 1429 2830
rect 1392 2800 1429 2810
rect 1488 2830 1575 2840
rect 1488 2810 1497 2830
rect 1517 2810 1575 2830
rect 1488 2801 1575 2810
rect 1488 2800 1525 2801
rect 109 2743 795 2776
rect 1544 2748 1575 2801
rect 1605 2830 1642 2909
rect 1813 2928 1845 2940
rect 1813 2908 1815 2928
rect 1836 2926 1845 2928
rect 1836 2924 2188 2926
rect 1836 2908 2206 2924
rect 1813 2906 2206 2908
rect 2226 2906 2229 2924
rect 1813 2901 2229 2906
rect 1813 2900 2154 2901
rect 1757 2840 1788 2841
rect 1605 2810 1614 2830
rect 1634 2810 1642 2830
rect 1605 2800 1642 2810
rect 1701 2833 1788 2840
rect 1701 2830 1762 2833
rect 1701 2810 1710 2830
rect 1730 2813 1762 2830
rect 1783 2813 1788 2833
rect 1730 2810 1788 2813
rect 1701 2803 1788 2810
rect 1813 2830 1850 2900
rect 2116 2899 2153 2900
rect 1965 2840 2001 2841
rect 1813 2810 1822 2830
rect 1842 2810 1850 2830
rect 1701 2801 1757 2803
rect 1701 2800 1738 2801
rect 1813 2800 1850 2810
rect 1909 2830 2057 2840
rect 2157 2837 2253 2839
rect 1909 2810 1918 2830
rect 1938 2821 2028 2830
rect 1938 2810 1969 2821
rect 1909 2801 1969 2810
rect 1909 2800 1946 2801
rect 1965 2789 1969 2801
rect 1996 2810 2028 2821
rect 2048 2810 2057 2830
rect 1996 2801 2057 2810
rect 2115 2830 2253 2837
rect 2115 2810 2124 2830
rect 2144 2810 2253 2830
rect 2115 2801 2253 2810
rect 1996 2789 2001 2801
rect 2020 2800 2057 2801
rect 2116 2800 2153 2801
rect 1965 2749 2001 2789
rect 1436 2747 1477 2748
rect 108 2686 147 2743
rect 757 2741 795 2743
rect 1328 2740 1477 2747
rect 1328 2720 1446 2740
rect 1466 2720 1477 2740
rect 1328 2712 1477 2720
rect 1544 2744 1903 2748
rect 1544 2739 1866 2744
rect 1544 2715 1657 2739
rect 1681 2720 1866 2739
rect 1890 2720 1903 2744
rect 1681 2715 1903 2720
rect 1544 2712 1903 2715
rect 1965 2712 2000 2749
rect 2068 2746 2168 2749
rect 2068 2742 2135 2746
rect 2068 2716 2080 2742
rect 2106 2720 2135 2742
rect 2161 2720 2168 2746
rect 2106 2716 2168 2720
rect 2068 2712 2168 2716
rect 1544 2691 1575 2712
rect 1965 2691 2001 2712
rect 1387 2690 1424 2691
rect 108 2684 156 2686
rect 108 2666 119 2684
rect 137 2666 156 2684
rect 1386 2681 1424 2690
rect 108 2657 156 2666
rect 109 2656 156 2657
rect 422 2661 532 2675
rect 422 2658 465 2661
rect 422 2653 426 2658
rect 344 2631 426 2653
rect 455 2631 465 2658
rect 493 2634 500 2661
rect 529 2653 532 2661
rect 1386 2661 1395 2681
rect 1415 2661 1424 2681
rect 1386 2653 1424 2661
rect 1490 2685 1575 2691
rect 1600 2690 1637 2691
rect 1490 2665 1498 2685
rect 1518 2665 1575 2685
rect 1490 2657 1575 2665
rect 1599 2681 1637 2690
rect 1599 2661 1608 2681
rect 1628 2661 1637 2681
rect 1490 2656 1526 2657
rect 1599 2653 1637 2661
rect 1703 2685 1788 2691
rect 1808 2690 1845 2691
rect 1703 2665 1711 2685
rect 1731 2684 1788 2685
rect 1731 2665 1760 2684
rect 1703 2664 1760 2665
rect 1781 2664 1788 2684
rect 1703 2657 1788 2664
rect 1807 2681 1845 2690
rect 1807 2661 1816 2681
rect 1836 2661 1845 2681
rect 1703 2656 1739 2657
rect 1807 2653 1845 2661
rect 1911 2685 2055 2691
rect 1911 2665 1919 2685
rect 1939 2665 2027 2685
rect 2047 2665 2055 2685
rect 1911 2657 2055 2665
rect 1911 2656 1947 2657
rect 2019 2656 2055 2657
rect 2121 2690 2158 2691
rect 2121 2689 2159 2690
rect 2121 2681 2185 2689
rect 2121 2661 2130 2681
rect 2150 2667 2185 2681
rect 2205 2667 2208 2687
rect 2150 2662 2208 2667
rect 2150 2661 2185 2662
rect 529 2634 594 2653
rect 493 2631 594 2634
rect 344 2629 594 2631
rect 112 2593 149 2594
rect 108 2590 149 2593
rect 108 2585 150 2590
rect 108 2567 121 2585
rect 139 2567 150 2585
rect 108 2553 150 2567
rect 188 2553 235 2557
rect 108 2547 235 2553
rect 108 2518 196 2547
rect 225 2518 235 2547
rect 344 2550 381 2629
rect 422 2616 532 2629
rect 496 2560 527 2561
rect 344 2530 353 2550
rect 373 2530 381 2550
rect 344 2520 381 2530
rect 440 2550 527 2560
rect 440 2530 449 2550
rect 469 2530 527 2550
rect 440 2521 527 2530
rect 440 2520 477 2521
rect 108 2514 235 2518
rect 108 2497 147 2514
rect 188 2513 235 2514
rect 108 2479 119 2497
rect 137 2479 147 2497
rect 108 2470 147 2479
rect 109 2469 146 2470
rect 496 2468 527 2521
rect 557 2550 594 2629
rect 765 2626 1158 2646
rect 1178 2626 1181 2646
rect 765 2621 1181 2626
rect 1387 2624 1424 2653
rect 1388 2622 1424 2624
rect 1600 2622 1637 2653
rect 765 2620 1106 2621
rect 709 2560 740 2561
rect 557 2530 566 2550
rect 586 2530 594 2550
rect 557 2520 594 2530
rect 653 2553 740 2560
rect 653 2550 714 2553
rect 653 2530 662 2550
rect 682 2533 714 2550
rect 735 2533 740 2553
rect 682 2530 740 2533
rect 653 2523 740 2530
rect 765 2550 802 2620
rect 1068 2619 1105 2620
rect 1388 2600 1637 2622
rect 1808 2621 1845 2653
rect 2121 2649 2185 2661
rect 2225 2631 2252 2801
rect 2683 2768 2710 2944
rect 2750 2908 2814 2920
rect 3090 2916 3127 2948
rect 3298 2947 3547 2969
rect 3830 2949 3867 2950
rect 4133 2949 4170 3019
rect 4195 3039 4282 3046
rect 4195 3036 4253 3039
rect 4195 3016 4200 3036
rect 4221 3019 4253 3036
rect 4273 3019 4282 3039
rect 4221 3016 4282 3019
rect 4195 3009 4282 3016
rect 4341 3039 4378 3049
rect 4341 3019 4349 3039
rect 4369 3019 4378 3039
rect 4195 3008 4226 3009
rect 3829 2948 4170 2949
rect 3298 2916 3335 2947
rect 3511 2945 3547 2947
rect 3511 2916 3548 2945
rect 3754 2943 4170 2948
rect 3754 2923 3757 2943
rect 3777 2923 4170 2943
rect 4341 2940 4378 3019
rect 4408 3048 4439 3101
rect 4789 3099 4826 3100
rect 4788 3090 4827 3099
rect 4788 3072 4798 3090
rect 4816 3072 4827 3090
rect 5168 3088 5205 3092
rect 4700 3055 4747 3056
rect 4788 3055 4827 3072
rect 4700 3051 4827 3055
rect 4458 3048 4495 3049
rect 4408 3039 4495 3048
rect 4408 3019 4466 3039
rect 4486 3019 4495 3039
rect 4408 3009 4495 3019
rect 4554 3039 4591 3049
rect 4554 3019 4562 3039
rect 4582 3019 4591 3039
rect 4408 3008 4439 3009
rect 4403 2940 4513 2953
rect 4554 2940 4591 3019
rect 4700 3022 4710 3051
rect 4739 3022 4827 3051
rect 4700 3016 4827 3022
rect 4700 3012 4747 3016
rect 4785 3002 4827 3016
rect 4785 2984 4796 3002
rect 4814 2984 4827 3002
rect 4785 2979 4827 2984
rect 4786 2976 4827 2979
rect 5165 3083 5205 3088
rect 5165 3065 5177 3083
rect 5195 3065 5205 3083
rect 4786 2975 4823 2976
rect 4341 2938 4591 2940
rect 4341 2935 4442 2938
rect 4341 2916 4406 2935
rect 2750 2907 2785 2908
rect 2727 2902 2785 2907
rect 2727 2882 2730 2902
rect 2750 2888 2785 2902
rect 2805 2888 2814 2908
rect 2750 2880 2814 2888
rect 2776 2879 2814 2880
rect 2777 2878 2814 2879
rect 2880 2912 2916 2913
rect 2988 2912 3024 2913
rect 2880 2905 3024 2912
rect 2880 2904 2938 2905
rect 2880 2884 2888 2904
rect 2908 2886 2938 2904
rect 2967 2904 3024 2905
rect 2967 2886 2996 2904
rect 2908 2884 2996 2886
rect 3016 2884 3024 2904
rect 2880 2878 3024 2884
rect 3090 2908 3128 2916
rect 3196 2912 3232 2913
rect 3090 2888 3099 2908
rect 3119 2888 3128 2908
rect 3090 2879 3128 2888
rect 3147 2905 3232 2912
rect 3147 2885 3154 2905
rect 3175 2904 3232 2905
rect 3175 2885 3204 2904
rect 3147 2884 3204 2885
rect 3224 2884 3232 2904
rect 3090 2878 3127 2879
rect 3147 2878 3232 2884
rect 3298 2908 3336 2916
rect 3409 2912 3445 2913
rect 3298 2888 3307 2908
rect 3327 2888 3336 2908
rect 3298 2879 3336 2888
rect 3360 2904 3445 2912
rect 3360 2884 3417 2904
rect 3437 2884 3445 2904
rect 3298 2878 3335 2879
rect 3360 2878 3445 2884
rect 3511 2908 3549 2916
rect 3511 2888 3520 2908
rect 3540 2888 3549 2908
rect 4403 2908 4406 2916
rect 4435 2908 4442 2935
rect 4470 2911 4480 2938
rect 4509 2916 4591 2938
rect 4509 2911 4513 2916
rect 4470 2908 4513 2911
rect 4403 2894 4513 2908
rect 4779 2912 4826 2913
rect 4779 2903 4827 2912
rect 3511 2879 3549 2888
rect 4779 2885 4798 2903
rect 4816 2885 4827 2903
rect 4779 2883 4827 2885
rect 3511 2878 3548 2879
rect 2934 2857 2970 2878
rect 3360 2857 3391 2878
rect 2767 2853 2867 2857
rect 2767 2849 2829 2853
rect 2767 2823 2774 2849
rect 2800 2827 2829 2849
rect 2855 2827 2867 2853
rect 2800 2823 2867 2827
rect 2767 2820 2867 2823
rect 2935 2820 2970 2857
rect 3032 2854 3391 2857
rect 3032 2849 3254 2854
rect 3032 2825 3045 2849
rect 3069 2830 3254 2849
rect 3278 2830 3391 2854
rect 3069 2825 3391 2830
rect 3032 2821 3391 2825
rect 3458 2849 3607 2857
rect 3458 2829 3469 2849
rect 3489 2829 3607 2849
rect 3458 2822 3607 2829
rect 4140 2826 4178 2828
rect 4788 2826 4827 2883
rect 5165 2885 5205 3065
rect 5551 3058 5582 3111
rect 5612 3140 5649 3219
rect 5820 3216 6213 3236
rect 6233 3216 6236 3236
rect 6334 3220 6583 3242
rect 6752 3241 6793 3246
rect 7171 3243 7198 3421
rect 7849 3333 7876 3511
rect 8254 3508 8295 3513
rect 8464 3512 8713 3534
rect 8811 3518 8814 3538
rect 8834 3518 9227 3538
rect 9398 3535 9435 3614
rect 9465 3643 9496 3696
rect 9842 3689 9882 3869
rect 10139 3952 10179 4132
rect 10525 4125 10556 4178
rect 10586 4207 10623 4286
rect 10794 4283 11187 4303
rect 11207 4283 11210 4303
rect 11308 4287 11557 4309
rect 11726 4308 11767 4313
rect 12145 4310 12172 4488
rect 12823 4400 12850 4578
rect 13228 4575 13269 4580
rect 13438 4579 13687 4601
rect 13785 4585 13788 4605
rect 13808 4585 14201 4605
rect 14372 4602 14409 4681
rect 14439 4710 14470 4763
rect 14816 4756 14856 4936
rect 15194 4938 15233 4976
rect 16413 4978 16531 4998
rect 16551 4978 16562 4998
rect 16413 4970 16562 4978
rect 16629 5002 16988 5006
rect 16629 4997 16951 5002
rect 16629 4973 16742 4997
rect 16766 4978 16951 4997
rect 16975 4978 16988 5002
rect 16766 4973 16988 4978
rect 16629 4970 16988 4973
rect 17050 4970 17085 5007
rect 17153 5004 17253 5007
rect 17153 5000 17220 5004
rect 17153 4974 17165 5000
rect 17191 4978 17220 5000
rect 17246 4978 17253 5004
rect 17191 4974 17253 4978
rect 17153 4970 17253 4974
rect 16629 4949 16660 4970
rect 17050 4949 17086 4970
rect 16472 4948 16509 4949
rect 16471 4939 16509 4948
rect 15194 4936 15242 4938
rect 15194 4918 15205 4936
rect 15223 4918 15242 4936
rect 15194 4909 15242 4918
rect 15195 4908 15242 4909
rect 15508 4913 15618 4927
rect 15508 4910 15551 4913
rect 15508 4905 15512 4910
rect 15430 4883 15512 4905
rect 15541 4883 15551 4910
rect 15579 4886 15586 4913
rect 15615 4905 15618 4913
rect 16471 4919 16480 4939
rect 16500 4919 16509 4939
rect 16471 4911 16509 4919
rect 16575 4943 16660 4949
rect 16685 4948 16722 4949
rect 16575 4923 16583 4943
rect 16603 4923 16660 4943
rect 16575 4915 16660 4923
rect 16684 4939 16722 4948
rect 16684 4919 16693 4939
rect 16713 4919 16722 4939
rect 16575 4914 16611 4915
rect 16684 4911 16722 4919
rect 16788 4943 16873 4949
rect 16893 4948 16930 4949
rect 16788 4923 16796 4943
rect 16816 4942 16873 4943
rect 16816 4923 16845 4942
rect 16788 4922 16845 4923
rect 16866 4922 16873 4942
rect 16788 4915 16873 4922
rect 16892 4939 16930 4948
rect 16892 4919 16901 4939
rect 16921 4919 16930 4939
rect 16788 4914 16824 4915
rect 16892 4911 16930 4919
rect 16996 4945 17140 4949
rect 16996 4943 17053 4945
rect 16996 4923 17004 4943
rect 17024 4923 17053 4943
rect 16996 4921 17053 4923
rect 17079 4943 17140 4945
rect 17079 4923 17112 4943
rect 17132 4923 17140 4943
rect 17079 4921 17140 4923
rect 16996 4915 17140 4921
rect 16996 4914 17032 4915
rect 17104 4914 17140 4915
rect 17206 4948 17243 4949
rect 17206 4947 17244 4948
rect 17206 4939 17270 4947
rect 17206 4919 17215 4939
rect 17235 4925 17270 4939
rect 17290 4925 17293 4945
rect 17235 4920 17293 4925
rect 17235 4919 17270 4920
rect 15615 4886 15680 4905
rect 15579 4883 15680 4886
rect 15430 4881 15680 4883
rect 15198 4845 15235 4846
rect 14816 4738 14826 4756
rect 14844 4738 14856 4756
rect 14816 4733 14856 4738
rect 15194 4842 15235 4845
rect 15194 4837 15236 4842
rect 15194 4819 15207 4837
rect 15225 4819 15236 4837
rect 15194 4805 15236 4819
rect 15274 4805 15321 4809
rect 15194 4799 15321 4805
rect 15194 4770 15282 4799
rect 15311 4770 15321 4799
rect 15430 4802 15467 4881
rect 15508 4868 15618 4881
rect 15582 4812 15613 4813
rect 15430 4782 15439 4802
rect 15459 4782 15467 4802
rect 15430 4772 15467 4782
rect 15526 4802 15613 4812
rect 15526 4782 15535 4802
rect 15555 4782 15613 4802
rect 15526 4773 15613 4782
rect 15526 4772 15563 4773
rect 15194 4766 15321 4770
rect 15194 4749 15233 4766
rect 15274 4765 15321 4766
rect 14816 4729 14853 4733
rect 15194 4731 15205 4749
rect 15223 4731 15233 4749
rect 15194 4722 15233 4731
rect 15195 4721 15232 4722
rect 15582 4720 15613 4773
rect 15643 4802 15680 4881
rect 15851 4878 16244 4898
rect 16264 4878 16267 4898
rect 16472 4882 16509 4911
rect 15851 4873 16267 4878
rect 16473 4880 16509 4882
rect 16685 4880 16722 4911
rect 15851 4872 16192 4873
rect 15795 4812 15826 4813
rect 15643 4782 15652 4802
rect 15672 4782 15680 4802
rect 15643 4772 15680 4782
rect 15739 4805 15826 4812
rect 15739 4802 15800 4805
rect 15739 4782 15748 4802
rect 15768 4785 15800 4802
rect 15821 4785 15826 4805
rect 15768 4782 15826 4785
rect 15739 4775 15826 4782
rect 15851 4802 15888 4872
rect 16154 4871 16191 4872
rect 16473 4858 16722 4880
rect 16893 4879 16930 4911
rect 17206 4907 17270 4919
rect 17310 4882 17337 5059
rect 17770 5014 17797 5191
rect 17837 5154 17901 5166
rect 18177 5162 18214 5194
rect 18385 5193 18634 5215
rect 18916 5201 18953 5202
rect 19219 5201 19256 5271
rect 19281 5291 19368 5298
rect 19281 5288 19339 5291
rect 19281 5268 19286 5288
rect 19307 5271 19339 5288
rect 19359 5271 19368 5291
rect 19307 5268 19368 5271
rect 19281 5261 19368 5268
rect 19427 5291 19464 5301
rect 19427 5271 19435 5291
rect 19455 5271 19464 5291
rect 19281 5260 19312 5261
rect 18915 5200 19256 5201
rect 18385 5162 18422 5193
rect 18598 5191 18634 5193
rect 18840 5195 19256 5200
rect 18598 5162 18635 5191
rect 18840 5175 18843 5195
rect 18863 5175 19256 5195
rect 19427 5192 19464 5271
rect 19494 5300 19525 5353
rect 19875 5351 19912 5352
rect 19874 5342 19913 5351
rect 19874 5324 19884 5342
rect 19902 5324 19913 5342
rect 19786 5307 19833 5308
rect 19874 5307 19913 5324
rect 19786 5303 19913 5307
rect 19544 5300 19581 5301
rect 19494 5291 19581 5300
rect 19494 5271 19552 5291
rect 19572 5271 19581 5291
rect 19494 5261 19581 5271
rect 19640 5291 19677 5301
rect 19640 5271 19648 5291
rect 19668 5271 19677 5291
rect 19494 5260 19525 5261
rect 19489 5192 19599 5205
rect 19640 5192 19677 5271
rect 19786 5274 19796 5303
rect 19825 5274 19913 5303
rect 19786 5268 19913 5274
rect 19786 5264 19833 5268
rect 19871 5254 19913 5268
rect 19871 5236 19882 5254
rect 19900 5236 19913 5254
rect 19871 5231 19913 5236
rect 19872 5228 19913 5231
rect 19872 5227 19909 5228
rect 19427 5190 19677 5192
rect 19427 5187 19528 5190
rect 19427 5168 19492 5187
rect 17837 5153 17872 5154
rect 17814 5148 17872 5153
rect 17814 5128 17817 5148
rect 17837 5134 17872 5148
rect 17892 5134 17901 5154
rect 17837 5126 17901 5134
rect 17863 5125 17901 5126
rect 17864 5124 17901 5125
rect 17967 5158 18003 5159
rect 18075 5158 18111 5159
rect 17967 5151 18111 5158
rect 17967 5150 18024 5151
rect 17967 5130 17975 5150
rect 17995 5131 18024 5150
rect 18049 5150 18111 5151
rect 18049 5131 18083 5150
rect 17995 5130 18083 5131
rect 18103 5130 18111 5150
rect 17967 5124 18111 5130
rect 18177 5154 18215 5162
rect 18283 5158 18319 5159
rect 18177 5134 18186 5154
rect 18206 5134 18215 5154
rect 18177 5125 18215 5134
rect 18234 5151 18319 5158
rect 18234 5131 18241 5151
rect 18262 5150 18319 5151
rect 18262 5131 18291 5150
rect 18234 5130 18291 5131
rect 18311 5130 18319 5150
rect 18177 5124 18214 5125
rect 18234 5124 18319 5130
rect 18385 5154 18423 5162
rect 18496 5158 18532 5159
rect 18385 5134 18394 5154
rect 18414 5134 18423 5154
rect 18385 5125 18423 5134
rect 18447 5150 18532 5158
rect 18447 5130 18504 5150
rect 18524 5130 18532 5150
rect 18385 5124 18422 5125
rect 18447 5124 18532 5130
rect 18598 5154 18636 5162
rect 18598 5134 18607 5154
rect 18627 5134 18636 5154
rect 19489 5160 19492 5168
rect 19521 5160 19528 5187
rect 19556 5163 19566 5190
rect 19595 5168 19677 5190
rect 19595 5163 19599 5168
rect 19556 5160 19599 5163
rect 19489 5146 19599 5160
rect 19865 5164 19912 5165
rect 19865 5155 19913 5164
rect 19865 5137 19884 5155
rect 19902 5137 19913 5155
rect 19865 5135 19913 5137
rect 18598 5125 18636 5134
rect 18598 5124 18635 5125
rect 18021 5103 18057 5124
rect 18447 5103 18478 5124
rect 17854 5099 17954 5103
rect 17854 5095 17916 5099
rect 17854 5069 17861 5095
rect 17887 5073 17916 5095
rect 17942 5073 17954 5099
rect 17887 5069 17954 5073
rect 17854 5066 17954 5069
rect 18022 5066 18057 5103
rect 18119 5100 18478 5103
rect 18119 5095 18341 5100
rect 18119 5071 18132 5095
rect 18156 5076 18341 5095
rect 18365 5076 18478 5100
rect 18156 5071 18478 5076
rect 18119 5067 18478 5071
rect 18545 5095 18694 5103
rect 18545 5075 18556 5095
rect 18576 5075 18694 5095
rect 19874 5097 19913 5135
rect 18545 5068 18694 5075
rect 19226 5078 19264 5080
rect 19874 5078 19916 5097
rect 18545 5067 18586 5068
rect 18021 5062 18057 5066
rect 18021 5033 18058 5062
rect 17869 5014 17906 5015
rect 17965 5014 18002 5015
rect 18021 5014 18057 5033
rect 18076 5014 18113 5015
rect 17769 5005 17907 5014
rect 17769 4985 17878 5005
rect 17898 4985 17907 5005
rect 17769 4978 17907 4985
rect 17965 5005 18113 5014
rect 17965 4985 17974 5005
rect 17994 4985 18084 5005
rect 18104 4985 18113 5005
rect 17769 4976 17865 4978
rect 17965 4975 18113 4985
rect 18172 5005 18209 5015
rect 18284 5014 18321 5015
rect 18265 5012 18321 5014
rect 18172 4985 18180 5005
rect 18200 4985 18209 5005
rect 18021 4974 18057 4975
rect 17869 4915 17906 4916
rect 18172 4915 18209 4985
rect 18234 5005 18321 5012
rect 18234 5002 18292 5005
rect 18234 4982 18239 5002
rect 18260 4985 18292 5002
rect 18312 4985 18321 5005
rect 18260 4982 18321 4985
rect 18234 4975 18321 4982
rect 18380 5005 18417 5015
rect 18380 4985 18388 5005
rect 18408 4985 18417 5005
rect 18234 4974 18265 4975
rect 17868 4914 18209 4915
rect 17793 4909 18209 4914
rect 17418 4882 17471 4890
rect 17793 4889 17796 4909
rect 17816 4889 18209 4909
rect 18380 4906 18417 4985
rect 18447 5014 18478 5067
rect 19226 5055 19916 5078
rect 19226 5045 19912 5055
rect 18497 5014 18534 5015
rect 18447 5005 18534 5014
rect 18447 4985 18505 5005
rect 18525 4985 18534 5005
rect 18447 4975 18534 4985
rect 18593 5005 18630 5015
rect 18593 4985 18601 5005
rect 18621 4985 18630 5005
rect 18447 4974 18478 4975
rect 18442 4906 18552 4919
rect 18593 4906 18630 4985
rect 18380 4904 18630 4906
rect 18380 4901 18481 4904
rect 18380 4882 18445 4901
rect 17285 4881 17471 4882
rect 17169 4879 17471 4881
rect 16554 4852 16665 4858
rect 16893 4853 17471 4879
rect 18442 4874 18445 4882
rect 18474 4874 18481 4901
rect 18509 4877 18519 4904
rect 18548 4882 18630 4904
rect 18818 4957 18986 4958
rect 19226 4957 19264 5045
rect 19525 5044 19572 5045
rect 19872 5021 19912 5045
rect 19489 4988 19601 5007
rect 19489 4987 19532 4988
rect 18818 4934 19264 4957
rect 19490 4986 19532 4987
rect 19490 4966 19497 4986
rect 19516 4966 19532 4986
rect 19490 4958 19532 4966
rect 19560 4986 19601 4988
rect 19560 4966 19574 4986
rect 19593 4966 19601 4986
rect 19873 4977 19912 5021
rect 19560 4958 19601 4966
rect 19490 4952 19601 4958
rect 18818 4931 19262 4934
rect 18818 4929 18986 4931
rect 18548 4877 18552 4882
rect 18509 4874 18552 4877
rect 18442 4860 18552 4874
rect 17169 4852 17471 4853
rect 16554 4844 16595 4852
rect 16554 4824 16562 4844
rect 16581 4824 16595 4844
rect 16554 4822 16595 4824
rect 16623 4844 16665 4852
rect 16623 4824 16639 4844
rect 16658 4824 16665 4844
rect 16623 4822 16665 4824
rect 16003 4812 16039 4813
rect 15851 4782 15860 4802
rect 15880 4782 15888 4802
rect 15739 4773 15795 4775
rect 15739 4772 15776 4773
rect 15851 4772 15888 4782
rect 15947 4802 16095 4812
rect 16195 4809 16291 4811
rect 15947 4782 15956 4802
rect 15976 4782 16066 4802
rect 16086 4782 16095 4802
rect 15947 4773 16095 4782
rect 16153 4802 16291 4809
rect 16554 4807 16665 4822
rect 16153 4782 16162 4802
rect 16182 4782 16291 4802
rect 16153 4773 16291 4782
rect 15947 4772 15984 4773
rect 16003 4721 16039 4773
rect 16058 4772 16095 4773
rect 16154 4772 16191 4773
rect 15474 4719 15515 4720
rect 15366 4712 15515 4719
rect 14489 4710 14526 4711
rect 14439 4701 14526 4710
rect 14439 4681 14497 4701
rect 14517 4681 14526 4701
rect 14439 4671 14526 4681
rect 14585 4701 14622 4711
rect 14585 4681 14593 4701
rect 14613 4681 14622 4701
rect 15366 4692 15484 4712
rect 15504 4692 15515 4712
rect 15366 4684 15515 4692
rect 15582 4716 15941 4720
rect 15582 4711 15904 4716
rect 15582 4687 15695 4711
rect 15719 4692 15904 4711
rect 15928 4692 15941 4716
rect 15719 4687 15941 4692
rect 15582 4684 15941 4687
rect 16003 4684 16038 4721
rect 16106 4718 16206 4721
rect 16106 4714 16173 4718
rect 16106 4688 16118 4714
rect 16144 4692 16173 4714
rect 16199 4692 16206 4718
rect 16144 4688 16206 4692
rect 16106 4684 16206 4688
rect 14439 4670 14470 4671
rect 14434 4602 14544 4615
rect 14585 4602 14622 4681
rect 14819 4666 14856 4667
rect 14815 4657 14856 4666
rect 15582 4663 15613 4684
rect 16003 4663 16039 4684
rect 15425 4662 15462 4663
rect 15199 4659 15233 4660
rect 14815 4639 14828 4657
rect 14846 4639 14856 4657
rect 14815 4630 14856 4639
rect 15198 4650 15235 4659
rect 15198 4632 15207 4650
rect 15225 4632 15235 4650
rect 14815 4610 14855 4630
rect 15198 4622 15235 4632
rect 15424 4653 15462 4662
rect 15424 4633 15433 4653
rect 15453 4633 15462 4653
rect 15424 4625 15462 4633
rect 15528 4657 15613 4663
rect 15638 4662 15675 4663
rect 15528 4637 15536 4657
rect 15556 4637 15613 4657
rect 15528 4629 15613 4637
rect 15637 4653 15675 4662
rect 15637 4633 15646 4653
rect 15666 4633 15675 4653
rect 15528 4628 15564 4629
rect 15637 4625 15675 4633
rect 15741 4657 15826 4663
rect 15846 4662 15883 4663
rect 15741 4637 15749 4657
rect 15769 4656 15826 4657
rect 15769 4637 15798 4656
rect 15741 4636 15798 4637
rect 15819 4636 15826 4656
rect 15741 4629 15826 4636
rect 15845 4653 15883 4662
rect 15845 4633 15854 4653
rect 15874 4633 15883 4653
rect 15741 4628 15777 4629
rect 15845 4625 15883 4633
rect 15949 4657 16093 4663
rect 15949 4637 15957 4657
rect 15977 4656 16065 4657
rect 15977 4637 16008 4656
rect 15949 4636 16008 4637
rect 16033 4637 16065 4656
rect 16085 4637 16093 4657
rect 16033 4636 16093 4637
rect 15949 4629 16093 4636
rect 15949 4628 15985 4629
rect 16057 4628 16093 4629
rect 16159 4662 16196 4663
rect 16159 4661 16197 4662
rect 16159 4653 16223 4661
rect 16159 4633 16168 4653
rect 16188 4639 16223 4653
rect 16243 4639 16246 4659
rect 16188 4634 16246 4639
rect 16188 4633 16223 4634
rect 14372 4600 14622 4602
rect 14372 4597 14473 4600
rect 12890 4540 12954 4552
rect 13230 4548 13267 4575
rect 13438 4548 13475 4579
rect 13651 4577 13687 4579
rect 14372 4578 14437 4597
rect 13651 4548 13688 4577
rect 14434 4570 14437 4578
rect 14466 4570 14473 4597
rect 14501 4573 14511 4600
rect 14540 4578 14622 4600
rect 14730 4600 14855 4610
rect 14730 4581 14738 4600
rect 14763 4581 14855 4600
rect 14540 4573 14544 4578
rect 14730 4574 14855 4581
rect 14501 4570 14544 4573
rect 14434 4556 14544 4570
rect 12890 4539 12925 4540
rect 12867 4534 12925 4539
rect 12867 4514 12870 4534
rect 12890 4520 12925 4534
rect 12945 4520 12954 4540
rect 12890 4512 12954 4520
rect 12916 4511 12954 4512
rect 12917 4510 12954 4511
rect 13020 4544 13056 4545
rect 13128 4544 13164 4545
rect 13020 4536 13164 4544
rect 13020 4516 13028 4536
rect 13048 4516 13136 4536
rect 13156 4516 13164 4536
rect 13020 4510 13164 4516
rect 13230 4540 13268 4548
rect 13336 4544 13372 4545
rect 13230 4520 13239 4540
rect 13259 4520 13268 4540
rect 13230 4511 13268 4520
rect 13287 4537 13372 4544
rect 13287 4517 13294 4537
rect 13315 4536 13372 4537
rect 13315 4517 13344 4536
rect 13287 4516 13344 4517
rect 13364 4516 13372 4536
rect 13230 4510 13267 4511
rect 13287 4510 13372 4516
rect 13438 4540 13476 4548
rect 13549 4544 13585 4545
rect 13438 4520 13447 4540
rect 13467 4520 13476 4540
rect 13438 4511 13476 4520
rect 13500 4536 13585 4544
rect 13500 4516 13557 4536
rect 13577 4516 13585 4536
rect 13438 4510 13475 4511
rect 13500 4510 13585 4516
rect 13651 4540 13689 4548
rect 13651 4520 13660 4540
rect 13680 4520 13689 4540
rect 13651 4511 13689 4520
rect 14815 4526 14855 4574
rect 15199 4594 15233 4622
rect 15425 4596 15462 4625
rect 15426 4594 15462 4596
rect 15638 4594 15675 4625
rect 15199 4593 15371 4594
rect 15199 4561 15385 4593
rect 15426 4572 15675 4594
rect 15846 4593 15883 4625
rect 16159 4621 16223 4633
rect 16263 4595 16290 4773
rect 17418 4745 17471 4852
rect 18818 4751 18845 4929
rect 18885 4891 18949 4903
rect 19225 4899 19262 4931
rect 19433 4930 19682 4952
rect 19433 4899 19470 4930
rect 19646 4928 19682 4930
rect 19646 4899 19683 4928
rect 18885 4890 18920 4891
rect 18862 4885 18920 4890
rect 18862 4865 18865 4885
rect 18885 4871 18920 4885
rect 18940 4871 18949 4891
rect 18885 4863 18949 4871
rect 18911 4862 18949 4863
rect 18912 4861 18949 4862
rect 19015 4895 19051 4896
rect 19123 4895 19159 4896
rect 19015 4890 19159 4895
rect 19015 4887 19077 4890
rect 19015 4867 19023 4887
rect 19043 4870 19077 4887
rect 19100 4887 19159 4890
rect 19100 4870 19131 4887
rect 19043 4867 19131 4870
rect 19151 4867 19159 4887
rect 19015 4861 19159 4867
rect 19225 4891 19263 4899
rect 19331 4895 19367 4896
rect 19225 4871 19234 4891
rect 19254 4871 19263 4891
rect 19225 4862 19263 4871
rect 19282 4888 19367 4895
rect 19282 4868 19289 4888
rect 19310 4887 19367 4888
rect 19310 4868 19339 4887
rect 19282 4867 19339 4868
rect 19359 4867 19367 4887
rect 19225 4861 19262 4862
rect 19282 4861 19367 4867
rect 19433 4891 19471 4899
rect 19544 4895 19580 4896
rect 19433 4871 19442 4891
rect 19462 4871 19471 4891
rect 19433 4862 19471 4871
rect 19495 4887 19580 4895
rect 19495 4867 19552 4887
rect 19572 4867 19580 4887
rect 19433 4861 19470 4862
rect 19495 4861 19580 4867
rect 19646 4891 19684 4899
rect 19646 4871 19655 4891
rect 19675 4871 19684 4891
rect 19646 4862 19684 4871
rect 19646 4861 19683 4862
rect 19069 4840 19105 4861
rect 19495 4840 19526 4861
rect 18902 4836 19002 4840
rect 18902 4832 18964 4836
rect 18902 4806 18909 4832
rect 18935 4810 18964 4832
rect 18990 4810 19002 4836
rect 18935 4806 19002 4810
rect 18902 4803 19002 4806
rect 19070 4803 19105 4840
rect 19167 4837 19526 4840
rect 19167 4832 19389 4837
rect 19167 4808 19180 4832
rect 19204 4813 19389 4832
rect 19413 4813 19526 4837
rect 19204 4808 19526 4813
rect 19167 4804 19526 4808
rect 19593 4832 19742 4840
rect 19593 4812 19604 4832
rect 19624 4812 19742 4832
rect 19593 4805 19742 4812
rect 19593 4804 19634 4805
rect 18917 4751 18954 4752
rect 19013 4751 19050 4752
rect 19069 4751 19105 4803
rect 19124 4751 19161 4752
rect 17418 4727 17466 4745
rect 17418 4687 17426 4727
rect 17453 4687 17466 4727
rect 18817 4742 18955 4751
rect 18817 4722 18926 4742
rect 18946 4722 18955 4742
rect 18817 4715 18955 4722
rect 19013 4742 19161 4751
rect 19013 4722 19022 4742
rect 19042 4722 19132 4742
rect 19152 4722 19161 4742
rect 18817 4713 18913 4715
rect 19013 4712 19161 4722
rect 19220 4742 19257 4752
rect 19332 4751 19369 4752
rect 19313 4749 19369 4751
rect 19220 4722 19228 4742
rect 19248 4722 19257 4742
rect 19069 4711 19105 4712
rect 16446 4669 16556 4683
rect 17418 4673 17466 4687
rect 18551 4678 18662 4693
rect 18551 4676 18593 4678
rect 16446 4666 16489 4669
rect 16446 4661 16450 4666
rect 16122 4593 16290 4595
rect 15846 4587 16290 4593
rect 15199 4529 15233 4561
rect 13651 4510 13688 4511
rect 13074 4489 13110 4510
rect 13500 4489 13531 4510
rect 14815 4508 14826 4526
rect 14844 4508 14855 4526
rect 14815 4500 14855 4508
rect 15195 4520 15233 4529
rect 15195 4502 15205 4520
rect 15223 4502 15233 4520
rect 14816 4499 14853 4500
rect 15195 4496 15233 4502
rect 15351 4498 15385 4561
rect 15507 4566 15618 4572
rect 15507 4558 15548 4566
rect 15507 4538 15515 4558
rect 15534 4538 15548 4558
rect 15507 4536 15548 4538
rect 15576 4558 15618 4566
rect 15576 4538 15592 4558
rect 15611 4538 15618 4558
rect 15576 4536 15618 4538
rect 15507 4521 15618 4536
rect 15845 4567 16290 4587
rect 15845 4498 15883 4567
rect 16122 4566 16290 4567
rect 16368 4639 16450 4661
rect 16479 4639 16489 4666
rect 16517 4642 16524 4669
rect 16553 4661 16556 4669
rect 16553 4642 16618 4661
rect 16517 4639 16618 4642
rect 16368 4637 16618 4639
rect 16368 4558 16405 4637
rect 16446 4624 16556 4637
rect 16520 4568 16551 4569
rect 16368 4538 16377 4558
rect 16397 4538 16405 4558
rect 16368 4528 16405 4538
rect 16464 4558 16551 4568
rect 16464 4538 16473 4558
rect 16493 4538 16551 4558
rect 16464 4529 16551 4538
rect 16464 4528 16501 4529
rect 15195 4492 15232 4496
rect 12907 4485 13007 4489
rect 12907 4481 12969 4485
rect 12907 4455 12914 4481
rect 12940 4459 12969 4481
rect 12995 4459 13007 4485
rect 12940 4455 13007 4459
rect 12907 4452 13007 4455
rect 13075 4452 13110 4489
rect 13172 4486 13531 4489
rect 13172 4481 13394 4486
rect 13172 4457 13185 4481
rect 13209 4462 13394 4481
rect 13418 4462 13531 4486
rect 13209 4457 13531 4462
rect 13172 4453 13531 4457
rect 13598 4481 13747 4489
rect 15351 4487 15883 4498
rect 13598 4461 13609 4481
rect 13629 4461 13747 4481
rect 15350 4471 15883 4487
rect 16520 4476 16551 4529
rect 16581 4558 16618 4637
rect 16789 4634 17182 4654
rect 17202 4634 17205 4654
rect 18284 4649 18325 4658
rect 16789 4629 17205 4634
rect 17879 4647 18047 4648
rect 18284 4647 18293 4649
rect 16789 4628 17130 4629
rect 16733 4568 16764 4569
rect 16581 4538 16590 4558
rect 16610 4538 16618 4558
rect 16581 4528 16618 4538
rect 16677 4561 16764 4568
rect 16677 4558 16738 4561
rect 16677 4538 16686 4558
rect 16706 4541 16738 4558
rect 16759 4541 16764 4561
rect 16706 4538 16764 4541
rect 16677 4531 16764 4538
rect 16789 4558 16826 4628
rect 17092 4627 17129 4628
rect 17879 4627 18293 4647
rect 18319 4627 18325 4649
rect 18551 4656 18558 4676
rect 18577 4656 18593 4676
rect 18551 4648 18593 4656
rect 18621 4676 18662 4678
rect 18621 4656 18635 4676
rect 18654 4656 18662 4676
rect 18621 4648 18662 4656
rect 18917 4652 18954 4653
rect 19220 4652 19257 4722
rect 19282 4742 19369 4749
rect 19282 4739 19340 4742
rect 19282 4719 19287 4739
rect 19308 4722 19340 4739
rect 19360 4722 19369 4742
rect 19308 4719 19369 4722
rect 19282 4712 19369 4719
rect 19428 4742 19465 4752
rect 19428 4722 19436 4742
rect 19456 4722 19465 4742
rect 19282 4711 19313 4712
rect 18916 4651 19257 4652
rect 18551 4642 18662 4648
rect 18841 4646 19257 4651
rect 17879 4621 18325 4627
rect 17879 4619 18047 4621
rect 16941 4568 16977 4569
rect 16789 4538 16798 4558
rect 16818 4538 16826 4558
rect 16677 4529 16733 4531
rect 16677 4528 16714 4529
rect 16789 4528 16826 4538
rect 16885 4558 17033 4568
rect 17133 4565 17229 4567
rect 16885 4538 16894 4558
rect 16914 4538 17004 4558
rect 17024 4538 17033 4558
rect 16885 4529 17033 4538
rect 17091 4558 17229 4565
rect 17091 4538 17100 4558
rect 17120 4538 17229 4558
rect 17091 4529 17229 4538
rect 16885 4528 16922 4529
rect 16941 4477 16977 4529
rect 16996 4528 17033 4529
rect 17092 4528 17129 4529
rect 16412 4475 16453 4476
rect 15350 4470 15864 4471
rect 13598 4454 13747 4461
rect 16304 4468 16453 4475
rect 14187 4458 14701 4459
rect 13598 4453 13639 4454
rect 13074 4417 13110 4452
rect 12922 4400 12959 4401
rect 13018 4400 13055 4401
rect 13074 4400 13081 4417
rect 12822 4391 12960 4400
rect 12822 4371 12931 4391
rect 12951 4371 12960 4391
rect 12822 4364 12960 4371
rect 13018 4391 13081 4400
rect 13018 4371 13027 4391
rect 13047 4376 13081 4391
rect 13102 4400 13110 4417
rect 13129 4400 13166 4401
rect 13102 4391 13166 4400
rect 13102 4376 13137 4391
rect 13047 4371 13137 4376
rect 13157 4371 13166 4391
rect 12822 4362 12918 4364
rect 13018 4361 13166 4371
rect 13225 4391 13262 4401
rect 13337 4400 13374 4401
rect 13318 4398 13374 4400
rect 13225 4371 13233 4391
rect 13253 4371 13262 4391
rect 13074 4360 13110 4361
rect 12004 4308 12172 4310
rect 11726 4302 12172 4308
rect 10794 4278 11210 4283
rect 11389 4281 11500 4287
rect 10794 4277 11135 4278
rect 10738 4217 10769 4218
rect 10586 4187 10595 4207
rect 10615 4187 10623 4207
rect 10586 4177 10623 4187
rect 10682 4210 10769 4217
rect 10682 4207 10743 4210
rect 10682 4187 10691 4207
rect 10711 4190 10743 4207
rect 10764 4190 10769 4210
rect 10711 4187 10769 4190
rect 10682 4180 10769 4187
rect 10794 4207 10831 4277
rect 11097 4276 11134 4277
rect 11389 4273 11430 4281
rect 11389 4253 11397 4273
rect 11416 4253 11430 4273
rect 11389 4251 11430 4253
rect 11458 4273 11500 4281
rect 11458 4253 11474 4273
rect 11493 4253 11500 4273
rect 11726 4280 11732 4302
rect 11758 4282 12172 4302
rect 12922 4301 12959 4302
rect 13225 4301 13262 4371
rect 13287 4391 13374 4398
rect 13287 4388 13345 4391
rect 13287 4368 13292 4388
rect 13313 4371 13345 4388
rect 13365 4371 13374 4391
rect 13313 4368 13374 4371
rect 13287 4361 13374 4368
rect 13433 4391 13470 4401
rect 13433 4371 13441 4391
rect 13461 4371 13470 4391
rect 13287 4360 13318 4361
rect 12921 4300 13262 4301
rect 11758 4280 11767 4282
rect 12004 4281 12172 4282
rect 12846 4299 13262 4300
rect 12846 4295 13222 4299
rect 11726 4271 11767 4280
rect 12846 4275 12849 4295
rect 12869 4282 13222 4295
rect 13254 4282 13262 4299
rect 12869 4275 13262 4282
rect 13433 4292 13470 4371
rect 13500 4400 13531 4453
rect 14168 4442 14701 4458
rect 16304 4448 16422 4468
rect 16442 4448 16453 4468
rect 14168 4431 14700 4442
rect 16304 4440 16453 4448
rect 16520 4472 16879 4476
rect 16520 4467 16842 4472
rect 16520 4443 16633 4467
rect 16657 4448 16842 4467
rect 16866 4448 16879 4472
rect 16657 4443 16879 4448
rect 16520 4440 16879 4443
rect 16941 4440 16976 4477
rect 17044 4474 17144 4477
rect 17044 4470 17111 4474
rect 17044 4444 17056 4470
rect 17082 4448 17111 4470
rect 17137 4448 17144 4474
rect 17082 4444 17144 4448
rect 17044 4440 17144 4444
rect 14819 4433 14856 4437
rect 13550 4400 13587 4401
rect 13500 4391 13587 4400
rect 13500 4371 13558 4391
rect 13578 4371 13587 4391
rect 13500 4361 13587 4371
rect 13646 4391 13683 4401
rect 13646 4371 13654 4391
rect 13674 4371 13683 4391
rect 13500 4360 13531 4361
rect 13495 4292 13605 4305
rect 13646 4292 13683 4371
rect 13433 4290 13683 4292
rect 13433 4287 13534 4290
rect 13433 4268 13498 4287
rect 11458 4251 11500 4253
rect 11389 4236 11500 4251
rect 13495 4260 13498 4268
rect 13527 4260 13534 4287
rect 13562 4263 13572 4290
rect 13601 4268 13683 4290
rect 13761 4362 13929 4363
rect 14168 4362 14206 4431
rect 13761 4342 14206 4362
rect 14433 4393 14544 4408
rect 14433 4391 14475 4393
rect 14433 4371 14440 4391
rect 14459 4371 14475 4391
rect 14433 4363 14475 4371
rect 14503 4391 14544 4393
rect 14503 4371 14517 4391
rect 14536 4371 14544 4391
rect 14503 4363 14544 4371
rect 14433 4357 14544 4363
rect 14666 4368 14700 4431
rect 14818 4427 14856 4433
rect 15198 4429 15235 4430
rect 14818 4409 14828 4427
rect 14846 4409 14856 4427
rect 14818 4400 14856 4409
rect 15196 4421 15236 4429
rect 15196 4403 15207 4421
rect 15225 4403 15236 4421
rect 16520 4419 16551 4440
rect 16941 4419 16977 4440
rect 16363 4418 16400 4419
rect 14818 4368 14852 4400
rect 13761 4336 14205 4342
rect 13761 4334 13929 4336
rect 13601 4263 13605 4268
rect 13562 4260 13605 4263
rect 13495 4246 13605 4260
rect 10946 4217 10982 4218
rect 10794 4187 10803 4207
rect 10823 4187 10831 4207
rect 10682 4178 10738 4180
rect 10682 4177 10719 4178
rect 10794 4177 10831 4187
rect 10890 4207 11038 4217
rect 11138 4214 11234 4216
rect 10890 4187 10899 4207
rect 10919 4187 11009 4207
rect 11029 4187 11038 4207
rect 10890 4178 11038 4187
rect 11096 4207 11234 4214
rect 11096 4187 11105 4207
rect 11125 4187 11234 4207
rect 11096 4178 11234 4187
rect 10890 4177 10927 4178
rect 10946 4126 10982 4178
rect 11001 4177 11038 4178
rect 11097 4177 11134 4178
rect 10417 4124 10458 4125
rect 10309 4117 10458 4124
rect 10309 4097 10427 4117
rect 10447 4097 10458 4117
rect 10309 4089 10458 4097
rect 10525 4121 10884 4125
rect 10525 4116 10847 4121
rect 10525 4092 10638 4116
rect 10662 4097 10847 4116
rect 10871 4097 10884 4121
rect 10662 4092 10884 4097
rect 10525 4089 10884 4092
rect 10946 4089 10981 4126
rect 11049 4123 11149 4126
rect 11049 4119 11116 4123
rect 11049 4093 11061 4119
rect 11087 4097 11116 4119
rect 11142 4097 11149 4123
rect 11087 4093 11149 4097
rect 11049 4089 11149 4093
rect 10525 4068 10556 4089
rect 10946 4068 10982 4089
rect 10368 4067 10405 4068
rect 10367 4058 10405 4067
rect 10367 4038 10376 4058
rect 10396 4038 10405 4058
rect 10367 4030 10405 4038
rect 10471 4062 10556 4068
rect 10581 4067 10618 4068
rect 10471 4042 10479 4062
rect 10499 4042 10556 4062
rect 10471 4034 10556 4042
rect 10580 4058 10618 4067
rect 10580 4038 10589 4058
rect 10609 4038 10618 4058
rect 10471 4033 10507 4034
rect 10580 4030 10618 4038
rect 10684 4062 10769 4068
rect 10789 4067 10826 4068
rect 10684 4042 10692 4062
rect 10712 4061 10769 4062
rect 10712 4042 10741 4061
rect 10684 4041 10741 4042
rect 10762 4041 10769 4061
rect 10684 4034 10769 4041
rect 10788 4058 10826 4067
rect 10788 4038 10797 4058
rect 10817 4038 10826 4058
rect 10684 4033 10720 4034
rect 10788 4030 10826 4038
rect 10892 4062 11036 4068
rect 10892 4042 10900 4062
rect 10920 4059 11008 4062
rect 10920 4042 10951 4059
rect 10892 4039 10951 4042
rect 10974 4042 11008 4059
rect 11028 4042 11036 4062
rect 10974 4039 11036 4042
rect 10892 4034 11036 4039
rect 10892 4033 10928 4034
rect 11000 4033 11036 4034
rect 11102 4067 11139 4068
rect 11102 4066 11140 4067
rect 11102 4058 11166 4066
rect 11102 4038 11111 4058
rect 11131 4044 11166 4058
rect 11186 4044 11189 4064
rect 11131 4039 11189 4044
rect 11131 4038 11166 4039
rect 10368 4001 10405 4030
rect 10369 3999 10405 4001
rect 10581 3999 10618 4030
rect 10369 3977 10618 3999
rect 10789 3998 10826 4030
rect 11102 4026 11166 4038
rect 11206 4000 11233 4178
rect 13761 4156 13788 4334
rect 13828 4296 13892 4308
rect 14168 4304 14205 4336
rect 14376 4335 14625 4357
rect 14666 4336 14852 4368
rect 14680 4335 14852 4336
rect 14376 4304 14413 4335
rect 14589 4333 14625 4335
rect 14589 4304 14626 4333
rect 14818 4307 14852 4335
rect 15196 4355 15236 4403
rect 16362 4409 16400 4418
rect 16362 4389 16371 4409
rect 16391 4389 16400 4409
rect 16362 4381 16400 4389
rect 16466 4413 16551 4419
rect 16576 4418 16613 4419
rect 16466 4393 16474 4413
rect 16494 4393 16551 4413
rect 16466 4385 16551 4393
rect 16575 4409 16613 4418
rect 16575 4389 16584 4409
rect 16604 4389 16613 4409
rect 16466 4384 16502 4385
rect 16575 4381 16613 4389
rect 16679 4413 16764 4419
rect 16784 4418 16821 4419
rect 16679 4393 16687 4413
rect 16707 4412 16764 4413
rect 16707 4393 16736 4412
rect 16679 4392 16736 4393
rect 16757 4392 16764 4412
rect 16679 4385 16764 4392
rect 16783 4409 16821 4418
rect 16783 4389 16792 4409
rect 16812 4389 16821 4409
rect 16679 4384 16715 4385
rect 16783 4381 16821 4389
rect 16887 4413 17031 4419
rect 16887 4393 16895 4413
rect 16915 4396 16951 4413
rect 16971 4396 17003 4413
rect 16915 4393 17003 4396
rect 17023 4393 17031 4413
rect 16887 4385 17031 4393
rect 16887 4384 16923 4385
rect 16995 4384 17031 4385
rect 17097 4418 17134 4419
rect 17097 4417 17135 4418
rect 17097 4409 17161 4417
rect 17097 4389 17106 4409
rect 17126 4395 17161 4409
rect 17181 4395 17184 4415
rect 17126 4390 17184 4395
rect 17126 4389 17161 4390
rect 15507 4359 15617 4373
rect 15507 4356 15550 4359
rect 15196 4348 15321 4355
rect 15507 4351 15511 4356
rect 15196 4329 15288 4348
rect 15313 4329 15321 4348
rect 15196 4319 15321 4329
rect 15429 4329 15511 4351
rect 15540 4329 15550 4356
rect 15578 4332 15585 4359
rect 15614 4351 15617 4359
rect 16363 4352 16400 4381
rect 15614 4332 15679 4351
rect 16364 4350 16400 4352
rect 16576 4350 16613 4381
rect 16784 4354 16821 4381
rect 17097 4377 17161 4389
rect 15578 4329 15679 4332
rect 15429 4327 15679 4329
rect 13828 4295 13863 4296
rect 13805 4290 13863 4295
rect 13805 4270 13808 4290
rect 13828 4276 13863 4290
rect 13883 4276 13892 4296
rect 13828 4268 13892 4276
rect 13854 4267 13892 4268
rect 13855 4266 13892 4267
rect 13958 4300 13994 4301
rect 14066 4300 14102 4301
rect 13958 4293 14102 4300
rect 13958 4292 14018 4293
rect 13958 4272 13966 4292
rect 13986 4273 14018 4292
rect 14043 4292 14102 4293
rect 14043 4273 14074 4292
rect 13986 4272 14074 4273
rect 14094 4272 14102 4292
rect 13958 4266 14102 4272
rect 14168 4296 14206 4304
rect 14274 4300 14310 4301
rect 14168 4276 14177 4296
rect 14197 4276 14206 4296
rect 14168 4267 14206 4276
rect 14225 4293 14310 4300
rect 14225 4273 14232 4293
rect 14253 4292 14310 4293
rect 14253 4273 14282 4292
rect 14225 4272 14282 4273
rect 14302 4272 14310 4292
rect 14168 4266 14205 4267
rect 14225 4266 14310 4272
rect 14376 4296 14414 4304
rect 14487 4300 14523 4301
rect 14376 4276 14385 4296
rect 14405 4276 14414 4296
rect 14376 4267 14414 4276
rect 14438 4292 14523 4300
rect 14438 4272 14495 4292
rect 14515 4272 14523 4292
rect 14376 4266 14413 4267
rect 14438 4266 14523 4272
rect 14589 4296 14627 4304
rect 14589 4276 14598 4296
rect 14618 4276 14627 4296
rect 14589 4267 14627 4276
rect 14816 4297 14853 4307
rect 15196 4299 15236 4319
rect 14816 4279 14826 4297
rect 14844 4279 14853 4297
rect 14816 4270 14853 4279
rect 15195 4290 15236 4299
rect 15195 4272 15205 4290
rect 15223 4272 15236 4290
rect 14818 4269 14852 4270
rect 14589 4266 14626 4267
rect 14012 4245 14048 4266
rect 14438 4245 14469 4266
rect 15195 4263 15236 4272
rect 15195 4262 15232 4263
rect 15429 4248 15466 4327
rect 15507 4314 15617 4327
rect 15581 4258 15612 4259
rect 13845 4241 13945 4245
rect 13845 4237 13907 4241
rect 13845 4211 13852 4237
rect 13878 4215 13907 4237
rect 13933 4215 13945 4241
rect 13878 4211 13945 4215
rect 13845 4208 13945 4211
rect 14013 4208 14048 4245
rect 14110 4242 14469 4245
rect 14110 4237 14332 4242
rect 14110 4213 14123 4237
rect 14147 4218 14332 4237
rect 14356 4218 14469 4242
rect 14147 4213 14469 4218
rect 14110 4209 14469 4213
rect 14536 4237 14685 4245
rect 14536 4217 14547 4237
rect 14567 4217 14685 4237
rect 15429 4228 15438 4248
rect 15458 4228 15466 4248
rect 15429 4218 15466 4228
rect 15525 4248 15612 4258
rect 15525 4228 15534 4248
rect 15554 4228 15612 4248
rect 15525 4219 15612 4228
rect 15525 4218 15562 4219
rect 14536 4210 14685 4217
rect 14536 4209 14577 4210
rect 13860 4156 13897 4157
rect 13956 4156 13993 4157
rect 14012 4156 14048 4208
rect 14067 4156 14104 4157
rect 13760 4147 13898 4156
rect 13355 4126 13466 4141
rect 13355 4124 13397 4126
rect 13025 4103 13130 4105
rect 12681 4095 12851 4096
rect 13025 4095 13074 4103
rect 12681 4076 13074 4095
rect 13105 4076 13130 4103
rect 13355 4104 13362 4124
rect 13381 4104 13397 4124
rect 13355 4096 13397 4104
rect 13425 4124 13466 4126
rect 13425 4104 13439 4124
rect 13458 4104 13466 4124
rect 13760 4127 13869 4147
rect 13889 4127 13898 4147
rect 13760 4120 13898 4127
rect 13956 4147 14104 4156
rect 13956 4127 13965 4147
rect 13985 4127 14075 4147
rect 14095 4127 14104 4147
rect 13760 4118 13856 4120
rect 13956 4117 14104 4127
rect 14163 4147 14200 4157
rect 14275 4156 14312 4157
rect 14256 4154 14312 4156
rect 14163 4127 14171 4147
rect 14191 4127 14200 4147
rect 14012 4116 14048 4117
rect 13425 4096 13466 4104
rect 13355 4090 13466 4096
rect 12681 4069 13130 4076
rect 12681 4067 12851 4069
rect 11531 4036 11641 4050
rect 11531 4033 11574 4036
rect 11531 4028 11535 4033
rect 11065 3998 11233 4000
rect 10789 3995 11233 3998
rect 10450 3971 10561 3977
rect 10450 3963 10491 3971
rect 10139 3908 10178 3952
rect 10450 3943 10458 3963
rect 10477 3943 10491 3963
rect 10450 3941 10491 3943
rect 10519 3963 10561 3971
rect 10519 3943 10535 3963
rect 10554 3943 10561 3963
rect 10519 3941 10561 3943
rect 10450 3926 10561 3941
rect 10787 3972 11233 3995
rect 10139 3884 10179 3908
rect 10479 3884 10526 3886
rect 10787 3884 10825 3972
rect 11065 3971 11233 3972
rect 11453 4006 11535 4028
rect 11564 4006 11574 4033
rect 11602 4009 11609 4036
rect 11638 4028 11641 4036
rect 11638 4009 11703 4028
rect 11602 4006 11703 4009
rect 11453 4004 11703 4006
rect 11453 3925 11490 4004
rect 11531 3991 11641 4004
rect 11605 3935 11636 3936
rect 11453 3905 11462 3925
rect 11482 3905 11490 3925
rect 11453 3895 11490 3905
rect 11549 3925 11636 3935
rect 11549 3905 11558 3925
rect 11578 3905 11636 3925
rect 11549 3896 11636 3905
rect 11549 3895 11586 3896
rect 10139 3851 10825 3884
rect 10139 3794 10178 3851
rect 10787 3849 10825 3851
rect 11605 3843 11636 3896
rect 11666 3925 11703 4004
rect 11874 4017 12267 4021
rect 11874 4000 11893 4017
rect 11913 4001 12267 4017
rect 12287 4001 12290 4021
rect 11913 4000 12290 4001
rect 11874 3996 12290 4000
rect 11874 3995 12215 3996
rect 11818 3935 11849 3936
rect 11666 3905 11675 3925
rect 11695 3905 11703 3925
rect 11666 3895 11703 3905
rect 11762 3928 11849 3935
rect 11762 3925 11823 3928
rect 11762 3905 11771 3925
rect 11791 3908 11823 3925
rect 11844 3908 11849 3928
rect 11791 3905 11849 3908
rect 11762 3898 11849 3905
rect 11874 3925 11911 3995
rect 12177 3994 12214 3995
rect 12026 3935 12062 3936
rect 11874 3905 11883 3925
rect 11903 3905 11911 3925
rect 11762 3896 11818 3898
rect 11762 3895 11799 3896
rect 11874 3895 11911 3905
rect 11970 3925 12118 3935
rect 12218 3932 12314 3934
rect 11970 3905 11979 3925
rect 11999 3905 12089 3925
rect 12109 3905 12118 3925
rect 11970 3896 12118 3905
rect 12176 3925 12314 3932
rect 12176 3905 12185 3925
rect 12205 3905 12314 3925
rect 12176 3896 12314 3905
rect 11970 3895 12007 3896
rect 12026 3844 12062 3896
rect 12081 3895 12118 3896
rect 12177 3895 12214 3896
rect 11497 3842 11538 3843
rect 11389 3835 11538 3842
rect 11389 3815 11507 3835
rect 11527 3815 11538 3835
rect 11389 3807 11538 3815
rect 11605 3839 11964 3843
rect 11605 3834 11927 3839
rect 11605 3810 11718 3834
rect 11742 3815 11927 3834
rect 11951 3815 11964 3839
rect 11742 3810 11964 3815
rect 11605 3807 11964 3810
rect 12026 3807 12061 3844
rect 12129 3841 12229 3844
rect 12129 3837 12196 3841
rect 12129 3811 12141 3837
rect 12167 3815 12196 3837
rect 12222 3815 12229 3841
rect 12167 3811 12229 3815
rect 12129 3807 12229 3811
rect 10139 3792 10187 3794
rect 10139 3774 10150 3792
rect 10168 3774 10187 3792
rect 11605 3786 11636 3807
rect 12026 3786 12062 3807
rect 11448 3785 11485 3786
rect 10139 3765 10187 3774
rect 10140 3764 10187 3765
rect 10453 3769 10563 3783
rect 10453 3766 10496 3769
rect 10453 3761 10457 3766
rect 10375 3739 10457 3761
rect 10486 3739 10496 3766
rect 10524 3742 10531 3769
rect 10560 3761 10563 3769
rect 11447 3776 11485 3785
rect 10560 3742 10625 3761
rect 11447 3756 11456 3776
rect 11476 3756 11485 3776
rect 10524 3739 10625 3742
rect 10375 3737 10625 3739
rect 10143 3701 10180 3702
rect 9842 3671 9852 3689
rect 9870 3671 9882 3689
rect 9842 3666 9882 3671
rect 10139 3698 10180 3701
rect 10139 3693 10181 3698
rect 10139 3675 10152 3693
rect 10170 3675 10181 3693
rect 9842 3662 9879 3666
rect 10139 3661 10181 3675
rect 10219 3661 10266 3665
rect 10139 3655 10266 3661
rect 9515 3643 9552 3644
rect 9465 3634 9552 3643
rect 9465 3614 9523 3634
rect 9543 3614 9552 3634
rect 9465 3604 9552 3614
rect 9611 3634 9648 3644
rect 9611 3614 9619 3634
rect 9639 3614 9648 3634
rect 9465 3603 9496 3604
rect 9460 3535 9570 3548
rect 9611 3535 9648 3614
rect 10139 3626 10227 3655
rect 10256 3626 10266 3655
rect 10375 3658 10412 3737
rect 10453 3724 10563 3737
rect 10527 3668 10558 3669
rect 10375 3638 10384 3658
rect 10404 3638 10412 3658
rect 10375 3628 10412 3638
rect 10471 3658 10558 3668
rect 10471 3638 10480 3658
rect 10500 3638 10558 3658
rect 10471 3629 10558 3638
rect 10471 3628 10508 3629
rect 10139 3622 10266 3626
rect 10139 3605 10178 3622
rect 10219 3621 10266 3622
rect 9845 3599 9882 3600
rect 9841 3590 9882 3599
rect 9841 3572 9854 3590
rect 9872 3572 9882 3590
rect 10139 3587 10150 3605
rect 10168 3587 10178 3605
rect 10139 3578 10178 3587
rect 10140 3577 10177 3578
rect 10527 3576 10558 3629
rect 10588 3658 10625 3737
rect 10796 3734 11189 3754
rect 11209 3734 11212 3754
rect 11447 3748 11485 3756
rect 11551 3780 11636 3786
rect 11661 3785 11698 3786
rect 11551 3760 11559 3780
rect 11579 3760 11636 3780
rect 11551 3752 11636 3760
rect 11660 3776 11698 3785
rect 11660 3756 11669 3776
rect 11689 3756 11698 3776
rect 11551 3751 11587 3752
rect 11660 3748 11698 3756
rect 11764 3780 11849 3786
rect 11869 3785 11906 3786
rect 11764 3760 11772 3780
rect 11792 3779 11849 3780
rect 11792 3760 11821 3779
rect 11764 3759 11821 3760
rect 11842 3759 11849 3779
rect 11764 3752 11849 3759
rect 11868 3776 11906 3785
rect 11868 3756 11877 3776
rect 11897 3756 11906 3776
rect 11764 3751 11800 3752
rect 11868 3748 11906 3756
rect 11972 3780 12116 3786
rect 11972 3760 11980 3780
rect 12000 3778 12088 3780
rect 12000 3760 12029 3778
rect 11972 3757 12029 3760
rect 12056 3760 12088 3778
rect 12108 3760 12116 3780
rect 12056 3757 12116 3760
rect 11972 3752 12116 3757
rect 11972 3751 12008 3752
rect 12080 3751 12116 3752
rect 12182 3785 12219 3786
rect 12182 3784 12220 3785
rect 12182 3776 12246 3784
rect 12182 3756 12191 3776
rect 12211 3762 12246 3776
rect 12266 3762 12269 3782
rect 12211 3757 12269 3762
rect 12211 3756 12246 3757
rect 10796 3729 11212 3734
rect 10796 3728 11137 3729
rect 10740 3668 10771 3669
rect 10588 3638 10597 3658
rect 10617 3638 10625 3658
rect 10588 3628 10625 3638
rect 10684 3661 10771 3668
rect 10684 3658 10745 3661
rect 10684 3638 10693 3658
rect 10713 3641 10745 3658
rect 10766 3641 10771 3661
rect 10713 3638 10771 3641
rect 10684 3631 10771 3638
rect 10796 3658 10833 3728
rect 11099 3727 11136 3728
rect 11448 3719 11485 3748
rect 11449 3717 11485 3719
rect 11661 3717 11698 3748
rect 11449 3695 11698 3717
rect 11869 3716 11906 3748
rect 12182 3744 12246 3756
rect 12286 3718 12313 3896
rect 12681 3889 12710 4067
rect 12750 4029 12814 4041
rect 13090 4037 13127 4069
rect 13298 4068 13547 4090
rect 13298 4037 13335 4068
rect 13511 4066 13547 4068
rect 13511 4037 13548 4066
rect 13860 4057 13897 4058
rect 14163 4057 14200 4127
rect 14225 4147 14312 4154
rect 14225 4144 14283 4147
rect 14225 4124 14230 4144
rect 14251 4127 14283 4144
rect 14303 4127 14312 4147
rect 14251 4124 14312 4127
rect 14225 4117 14312 4124
rect 14371 4147 14408 4157
rect 14371 4127 14379 4147
rect 14399 4127 14408 4147
rect 14225 4116 14256 4117
rect 13859 4056 14200 4057
rect 13784 4051 14200 4056
rect 12750 4028 12785 4029
rect 12727 4023 12785 4028
rect 12727 4003 12730 4023
rect 12750 4009 12785 4023
rect 12805 4009 12814 4029
rect 12750 4001 12814 4009
rect 12776 4000 12814 4001
rect 12777 3999 12814 4000
rect 12880 4033 12916 4034
rect 12988 4033 13024 4034
rect 12880 4025 13024 4033
rect 12880 4005 12888 4025
rect 12908 4005 12996 4025
rect 13016 4005 13024 4025
rect 12880 3999 13024 4005
rect 13090 4029 13128 4037
rect 13196 4033 13232 4034
rect 13090 4009 13099 4029
rect 13119 4009 13128 4029
rect 13090 4000 13128 4009
rect 13147 4026 13232 4033
rect 13147 4006 13154 4026
rect 13175 4025 13232 4026
rect 13175 4006 13204 4025
rect 13147 4005 13204 4006
rect 13224 4005 13232 4025
rect 13090 3999 13127 4000
rect 13147 3999 13232 4005
rect 13298 4029 13336 4037
rect 13409 4033 13445 4034
rect 13298 4009 13307 4029
rect 13327 4009 13336 4029
rect 13298 4000 13336 4009
rect 13360 4025 13445 4033
rect 13360 4005 13417 4025
rect 13437 4005 13445 4025
rect 13298 3999 13335 4000
rect 13360 3999 13445 4005
rect 13511 4029 13549 4037
rect 13784 4031 13787 4051
rect 13807 4031 14200 4051
rect 14371 4048 14408 4127
rect 14438 4156 14469 4209
rect 14819 4207 14856 4208
rect 14818 4198 14857 4207
rect 14818 4180 14828 4198
rect 14846 4180 14857 4198
rect 15198 4196 15235 4200
rect 14730 4163 14777 4164
rect 14818 4163 14857 4180
rect 14730 4159 14857 4163
rect 14488 4156 14525 4157
rect 14438 4147 14525 4156
rect 14438 4127 14496 4147
rect 14516 4127 14525 4147
rect 14438 4117 14525 4127
rect 14584 4147 14621 4157
rect 14584 4127 14592 4147
rect 14612 4127 14621 4147
rect 14438 4116 14469 4117
rect 14433 4048 14543 4061
rect 14584 4048 14621 4127
rect 14730 4130 14740 4159
rect 14769 4130 14857 4159
rect 14730 4124 14857 4130
rect 14730 4120 14777 4124
rect 14815 4110 14857 4124
rect 14815 4092 14826 4110
rect 14844 4092 14857 4110
rect 14815 4087 14857 4092
rect 14816 4084 14857 4087
rect 15195 4191 15235 4196
rect 15195 4173 15207 4191
rect 15225 4173 15235 4191
rect 14816 4083 14853 4084
rect 14371 4046 14621 4048
rect 14371 4043 14472 4046
rect 13511 4009 13520 4029
rect 13540 4009 13549 4029
rect 14371 4024 14436 4043
rect 13511 4000 13549 4009
rect 14433 4016 14436 4024
rect 14465 4016 14472 4043
rect 14500 4019 14510 4046
rect 14539 4024 14621 4046
rect 14539 4019 14543 4024
rect 14500 4016 14543 4019
rect 14433 4002 14543 4016
rect 14809 4020 14856 4021
rect 14809 4011 14857 4020
rect 13511 3999 13548 4000
rect 12934 3978 12970 3999
rect 13360 3978 13391 3999
rect 14809 3993 14828 4011
rect 14846 3993 14857 4011
rect 14809 3991 14857 3993
rect 12767 3974 12867 3978
rect 12767 3970 12829 3974
rect 12767 3944 12774 3970
rect 12800 3948 12829 3970
rect 12855 3948 12867 3974
rect 12800 3944 12867 3948
rect 12767 3941 12867 3944
rect 12935 3941 12970 3978
rect 13032 3975 13391 3978
rect 13032 3970 13254 3975
rect 13032 3946 13045 3970
rect 13069 3951 13254 3970
rect 13278 3951 13391 3975
rect 13069 3946 13391 3951
rect 13032 3942 13391 3946
rect 13458 3970 13607 3978
rect 13458 3950 13469 3970
rect 13489 3950 13607 3970
rect 13458 3943 13607 3950
rect 13458 3942 13499 3943
rect 12934 3902 12970 3941
rect 12782 3889 12819 3890
rect 12878 3889 12915 3890
rect 12934 3889 12941 3902
rect 12681 3880 12820 3889
rect 12681 3860 12791 3880
rect 12811 3860 12820 3880
rect 12681 3853 12820 3860
rect 12878 3880 12941 3889
rect 12878 3860 12887 3880
rect 12907 3864 12941 3880
rect 12964 3889 12970 3902
rect 12989 3889 13026 3890
rect 12964 3880 13026 3889
rect 12964 3864 12997 3880
rect 12907 3860 12997 3864
rect 13017 3860 13026 3880
rect 12681 3851 12778 3853
rect 12681 3850 12710 3851
rect 12878 3850 13026 3860
rect 13085 3880 13122 3890
rect 13197 3889 13234 3890
rect 13178 3887 13234 3889
rect 13085 3860 13093 3880
rect 13113 3860 13122 3880
rect 12934 3849 12970 3850
rect 12782 3790 12819 3791
rect 13085 3790 13122 3860
rect 13147 3880 13234 3887
rect 13147 3877 13205 3880
rect 13147 3857 13152 3877
rect 13173 3860 13205 3877
rect 13225 3860 13234 3880
rect 13173 3857 13234 3860
rect 13147 3850 13234 3857
rect 13293 3880 13330 3890
rect 13293 3860 13301 3880
rect 13321 3860 13330 3880
rect 13147 3849 13178 3850
rect 12781 3789 13122 3790
rect 12706 3785 13122 3789
rect 12706 3784 13083 3785
rect 12706 3764 12709 3784
rect 12729 3768 13083 3784
rect 13103 3768 13122 3785
rect 12729 3764 13122 3768
rect 13293 3781 13330 3860
rect 13360 3889 13391 3942
rect 14171 3934 14209 3936
rect 14818 3934 14857 3991
rect 14171 3901 14857 3934
rect 13410 3889 13447 3890
rect 13360 3880 13447 3889
rect 13360 3860 13418 3880
rect 13438 3860 13447 3880
rect 13360 3850 13447 3860
rect 13506 3880 13543 3890
rect 13506 3860 13514 3880
rect 13534 3860 13543 3880
rect 13360 3849 13391 3850
rect 13355 3781 13465 3794
rect 13506 3781 13543 3860
rect 13293 3779 13543 3781
rect 13293 3776 13394 3779
rect 13293 3757 13358 3776
rect 13355 3749 13358 3757
rect 13387 3749 13394 3776
rect 13422 3752 13432 3779
rect 13461 3757 13543 3779
rect 13763 3813 13931 3814
rect 14171 3813 14209 3901
rect 14470 3899 14517 3901
rect 14817 3877 14857 3901
rect 13763 3790 14209 3813
rect 14435 3844 14546 3859
rect 14435 3842 14477 3844
rect 14435 3822 14442 3842
rect 14461 3822 14477 3842
rect 14435 3814 14477 3822
rect 14505 3842 14546 3844
rect 14505 3822 14519 3842
rect 14538 3822 14546 3842
rect 14818 3833 14857 3877
rect 14505 3814 14546 3822
rect 14435 3808 14546 3814
rect 13763 3787 14207 3790
rect 13763 3785 13931 3787
rect 13461 3752 13465 3757
rect 13422 3749 13465 3752
rect 13355 3735 13465 3749
rect 12145 3716 12313 3718
rect 11866 3709 12313 3716
rect 11530 3689 11641 3695
rect 11530 3681 11571 3689
rect 10948 3668 10984 3669
rect 10796 3638 10805 3658
rect 10825 3638 10833 3658
rect 10684 3629 10740 3631
rect 10684 3628 10721 3629
rect 10796 3628 10833 3638
rect 10892 3658 11040 3668
rect 11140 3665 11236 3667
rect 10892 3638 10901 3658
rect 10921 3638 11011 3658
rect 11031 3638 11040 3658
rect 10892 3629 11040 3638
rect 11098 3658 11236 3665
rect 11098 3638 11107 3658
rect 11127 3638 11236 3658
rect 11530 3661 11538 3681
rect 11557 3661 11571 3681
rect 11530 3659 11571 3661
rect 11599 3681 11641 3689
rect 11599 3661 11615 3681
rect 11634 3661 11641 3681
rect 11866 3682 11891 3709
rect 11922 3690 12313 3709
rect 11922 3682 11971 3690
rect 12145 3689 12313 3690
rect 11866 3680 11971 3682
rect 11599 3659 11641 3661
rect 11530 3644 11641 3659
rect 11098 3629 11236 3638
rect 10892 3628 10929 3629
rect 10948 3577 10984 3629
rect 11003 3628 11040 3629
rect 11099 3628 11136 3629
rect 10419 3575 10460 3576
rect 9841 3563 9882 3572
rect 10311 3568 10460 3575
rect 9841 3543 9881 3563
rect 9398 3533 9648 3535
rect 9398 3530 9499 3533
rect 7916 3473 7980 3485
rect 8256 3481 8293 3508
rect 8464 3481 8501 3512
rect 8677 3510 8713 3512
rect 9398 3511 9463 3530
rect 8677 3481 8714 3510
rect 9460 3503 9463 3511
rect 9492 3503 9499 3530
rect 9527 3506 9537 3533
rect 9566 3511 9648 3533
rect 9756 3533 9881 3543
rect 10311 3548 10429 3568
rect 10449 3548 10460 3568
rect 10311 3540 10460 3548
rect 10527 3572 10886 3576
rect 10527 3567 10849 3572
rect 10527 3543 10640 3567
rect 10664 3548 10849 3567
rect 10873 3548 10886 3572
rect 10664 3543 10886 3548
rect 10527 3540 10886 3543
rect 10948 3540 10983 3577
rect 11051 3574 11151 3577
rect 11051 3570 11118 3574
rect 11051 3544 11063 3570
rect 11089 3548 11118 3570
rect 11144 3548 11151 3574
rect 11089 3544 11151 3548
rect 11051 3540 11151 3544
rect 9756 3514 9764 3533
rect 9789 3514 9881 3533
rect 10527 3519 10558 3540
rect 10948 3519 10984 3540
rect 10370 3518 10407 3519
rect 10144 3515 10178 3516
rect 9566 3506 9570 3511
rect 9756 3507 9881 3514
rect 9527 3503 9570 3506
rect 9460 3489 9570 3503
rect 7916 3472 7951 3473
rect 7893 3467 7951 3472
rect 7893 3447 7896 3467
rect 7916 3453 7951 3467
rect 7971 3453 7980 3473
rect 7916 3445 7980 3453
rect 7942 3444 7980 3445
rect 7943 3443 7980 3444
rect 8046 3477 8082 3478
rect 8154 3477 8190 3478
rect 8046 3469 8190 3477
rect 8046 3449 8054 3469
rect 8074 3466 8162 3469
rect 8074 3449 8106 3466
rect 8126 3449 8162 3466
rect 8182 3449 8190 3469
rect 8046 3443 8190 3449
rect 8256 3473 8294 3481
rect 8362 3477 8398 3478
rect 8256 3453 8265 3473
rect 8285 3453 8294 3473
rect 8256 3444 8294 3453
rect 8313 3470 8398 3477
rect 8313 3450 8320 3470
rect 8341 3469 8398 3470
rect 8341 3450 8370 3469
rect 8313 3449 8370 3450
rect 8390 3449 8398 3469
rect 8256 3443 8293 3444
rect 8313 3443 8398 3449
rect 8464 3473 8502 3481
rect 8575 3477 8611 3478
rect 8464 3453 8473 3473
rect 8493 3453 8502 3473
rect 8464 3444 8502 3453
rect 8526 3469 8611 3477
rect 8526 3449 8583 3469
rect 8603 3449 8611 3469
rect 8464 3443 8501 3444
rect 8526 3443 8611 3449
rect 8677 3473 8715 3481
rect 8677 3453 8686 3473
rect 8706 3453 8715 3473
rect 8677 3444 8715 3453
rect 9841 3459 9881 3507
rect 10143 3506 10180 3515
rect 10143 3488 10152 3506
rect 10170 3488 10180 3506
rect 10143 3478 10180 3488
rect 10369 3509 10407 3518
rect 10369 3489 10378 3509
rect 10398 3489 10407 3509
rect 10369 3481 10407 3489
rect 10473 3513 10558 3519
rect 10583 3518 10620 3519
rect 10473 3493 10481 3513
rect 10501 3493 10558 3513
rect 10473 3485 10558 3493
rect 10582 3509 10620 3518
rect 10582 3489 10591 3509
rect 10611 3489 10620 3509
rect 10473 3484 10509 3485
rect 10582 3481 10620 3489
rect 10686 3513 10771 3519
rect 10791 3518 10828 3519
rect 10686 3493 10694 3513
rect 10714 3512 10771 3513
rect 10714 3493 10743 3512
rect 10686 3492 10743 3493
rect 10764 3492 10771 3512
rect 10686 3485 10771 3492
rect 10790 3509 10828 3518
rect 10790 3489 10799 3509
rect 10819 3489 10828 3509
rect 10686 3484 10722 3485
rect 10790 3481 10828 3489
rect 10894 3513 11038 3519
rect 10894 3493 10902 3513
rect 10922 3512 11010 3513
rect 10922 3493 10953 3512
rect 10894 3492 10953 3493
rect 10978 3493 11010 3512
rect 11030 3493 11038 3513
rect 10978 3492 11038 3493
rect 10894 3485 11038 3492
rect 10894 3484 10930 3485
rect 11002 3484 11038 3485
rect 11104 3518 11141 3519
rect 11104 3517 11142 3518
rect 11104 3509 11168 3517
rect 11104 3489 11113 3509
rect 11133 3495 11168 3509
rect 11188 3495 11191 3515
rect 11133 3490 11191 3495
rect 11133 3489 11168 3490
rect 8677 3443 8714 3444
rect 8100 3422 8136 3443
rect 8526 3422 8557 3443
rect 9841 3441 9852 3459
rect 9870 3441 9881 3459
rect 9841 3433 9881 3441
rect 10144 3450 10178 3478
rect 10370 3452 10407 3481
rect 10371 3450 10407 3452
rect 10583 3450 10620 3481
rect 10144 3449 10316 3450
rect 9842 3432 9879 3433
rect 7933 3418 8033 3422
rect 7933 3414 7995 3418
rect 7933 3388 7940 3414
rect 7966 3392 7995 3414
rect 8021 3392 8033 3418
rect 7966 3388 8033 3392
rect 7933 3385 8033 3388
rect 8101 3385 8136 3422
rect 8198 3419 8557 3422
rect 8198 3414 8420 3419
rect 8198 3390 8211 3414
rect 8235 3395 8420 3414
rect 8444 3395 8557 3419
rect 8235 3390 8557 3395
rect 8198 3386 8557 3390
rect 8624 3414 8773 3422
rect 8624 3394 8635 3414
rect 8655 3394 8773 3414
rect 8624 3387 8773 3394
rect 10144 3417 10330 3449
rect 10371 3428 10620 3450
rect 10791 3449 10828 3481
rect 11104 3477 11168 3489
rect 11208 3451 11235 3629
rect 13763 3607 13790 3785
rect 13830 3747 13894 3759
rect 14170 3755 14207 3787
rect 14378 3786 14627 3808
rect 14378 3755 14415 3786
rect 14591 3784 14627 3786
rect 14591 3755 14628 3784
rect 13830 3746 13865 3747
rect 13807 3741 13865 3746
rect 13807 3721 13810 3741
rect 13830 3727 13865 3741
rect 13885 3727 13894 3747
rect 13830 3719 13894 3727
rect 13856 3718 13894 3719
rect 13857 3717 13894 3718
rect 13960 3751 13996 3752
rect 14068 3751 14104 3752
rect 13960 3746 14104 3751
rect 13960 3743 14022 3746
rect 13960 3723 13968 3743
rect 13988 3726 14022 3743
rect 14045 3743 14104 3746
rect 14045 3726 14076 3743
rect 13988 3723 14076 3726
rect 14096 3723 14104 3743
rect 13960 3717 14104 3723
rect 14170 3747 14208 3755
rect 14276 3751 14312 3752
rect 14170 3727 14179 3747
rect 14199 3727 14208 3747
rect 14170 3718 14208 3727
rect 14227 3744 14312 3751
rect 14227 3724 14234 3744
rect 14255 3743 14312 3744
rect 14255 3724 14284 3743
rect 14227 3723 14284 3724
rect 14304 3723 14312 3743
rect 14170 3717 14207 3718
rect 14227 3717 14312 3723
rect 14378 3747 14416 3755
rect 14489 3751 14525 3752
rect 14378 3727 14387 3747
rect 14407 3727 14416 3747
rect 14378 3718 14416 3727
rect 14440 3743 14525 3751
rect 14440 3723 14497 3743
rect 14517 3723 14525 3743
rect 14378 3717 14415 3718
rect 14440 3717 14525 3723
rect 14591 3747 14629 3755
rect 14591 3727 14600 3747
rect 14620 3727 14629 3747
rect 14591 3718 14629 3727
rect 14591 3717 14628 3718
rect 14014 3696 14050 3717
rect 14440 3696 14471 3717
rect 13847 3692 13947 3696
rect 13847 3688 13909 3692
rect 13847 3662 13854 3688
rect 13880 3666 13909 3688
rect 13935 3666 13947 3692
rect 13880 3662 13947 3666
rect 13847 3659 13947 3662
rect 14015 3659 14050 3696
rect 14112 3693 14471 3696
rect 14112 3688 14334 3693
rect 14112 3664 14125 3688
rect 14149 3669 14334 3688
rect 14358 3669 14471 3693
rect 14149 3664 14471 3669
rect 14112 3660 14471 3664
rect 14538 3688 14687 3696
rect 14538 3668 14549 3688
rect 14569 3668 14687 3688
rect 14538 3661 14687 3668
rect 14538 3660 14579 3661
rect 13862 3607 13899 3608
rect 13958 3607 13995 3608
rect 14014 3607 14050 3659
rect 14069 3607 14106 3608
rect 13762 3598 13900 3607
rect 13762 3578 13871 3598
rect 13891 3578 13900 3598
rect 13762 3571 13900 3578
rect 13958 3598 14106 3607
rect 13958 3578 13967 3598
rect 13987 3578 14077 3598
rect 14097 3578 14106 3598
rect 13762 3569 13858 3571
rect 13958 3568 14106 3578
rect 14165 3598 14202 3608
rect 14277 3607 14314 3608
rect 14258 3605 14314 3607
rect 14165 3578 14173 3598
rect 14193 3578 14202 3598
rect 14014 3567 14050 3568
rect 11391 3525 11501 3539
rect 11391 3522 11434 3525
rect 11391 3517 11395 3522
rect 11067 3449 11235 3451
rect 10791 3443 11235 3449
rect 9213 3391 9727 3392
rect 8624 3386 8665 3387
rect 7948 3333 7985 3334
rect 8044 3333 8081 3334
rect 8100 3333 8136 3385
rect 8155 3333 8192 3334
rect 7848 3324 7986 3333
rect 7848 3304 7957 3324
rect 7977 3304 7986 3324
rect 7848 3297 7986 3304
rect 8044 3324 8192 3333
rect 8044 3304 8053 3324
rect 8073 3304 8163 3324
rect 8183 3304 8192 3324
rect 7848 3295 7944 3297
rect 8044 3294 8192 3304
rect 8251 3324 8288 3334
rect 8363 3333 8400 3334
rect 8344 3331 8400 3333
rect 8251 3304 8259 3324
rect 8279 3304 8288 3324
rect 8100 3293 8136 3294
rect 7030 3241 7198 3243
rect 6752 3235 7198 3241
rect 5820 3211 6236 3216
rect 6415 3214 6526 3220
rect 5820 3210 6161 3211
rect 5764 3150 5795 3151
rect 5612 3120 5621 3140
rect 5641 3120 5649 3140
rect 5612 3110 5649 3120
rect 5708 3143 5795 3150
rect 5708 3140 5769 3143
rect 5708 3120 5717 3140
rect 5737 3123 5769 3140
rect 5790 3123 5795 3143
rect 5737 3120 5795 3123
rect 5708 3113 5795 3120
rect 5820 3140 5857 3210
rect 6123 3209 6160 3210
rect 6415 3206 6456 3214
rect 6415 3186 6423 3206
rect 6442 3186 6456 3206
rect 6415 3184 6456 3186
rect 6484 3206 6526 3214
rect 6484 3186 6500 3206
rect 6519 3186 6526 3206
rect 6752 3213 6758 3235
rect 6784 3215 7198 3235
rect 7948 3234 7985 3235
rect 8251 3234 8288 3304
rect 8313 3324 8400 3331
rect 8313 3321 8371 3324
rect 8313 3301 8318 3321
rect 8339 3304 8371 3321
rect 8391 3304 8400 3324
rect 8339 3301 8400 3304
rect 8313 3294 8400 3301
rect 8459 3324 8496 3334
rect 8459 3304 8467 3324
rect 8487 3304 8496 3324
rect 8313 3293 8344 3294
rect 7947 3233 8288 3234
rect 6784 3213 6793 3215
rect 7030 3214 7198 3215
rect 7872 3228 8288 3233
rect 6752 3204 6793 3213
rect 7872 3208 7875 3228
rect 7895 3208 8288 3228
rect 8459 3225 8496 3304
rect 8526 3333 8557 3386
rect 9194 3375 9727 3391
rect 10144 3385 10178 3417
rect 10140 3376 10178 3385
rect 9194 3364 9726 3375
rect 9845 3366 9882 3370
rect 8576 3333 8613 3334
rect 8526 3324 8613 3333
rect 8526 3304 8584 3324
rect 8604 3304 8613 3324
rect 8526 3294 8613 3304
rect 8672 3324 8709 3334
rect 8672 3304 8680 3324
rect 8700 3304 8709 3324
rect 8526 3293 8557 3294
rect 8521 3225 8631 3238
rect 8672 3225 8709 3304
rect 8459 3223 8709 3225
rect 8459 3220 8560 3223
rect 8459 3201 8524 3220
rect 6484 3184 6526 3186
rect 6415 3169 6526 3184
rect 8521 3193 8524 3201
rect 8553 3193 8560 3220
rect 8588 3196 8598 3223
rect 8627 3201 8709 3223
rect 8787 3295 8955 3296
rect 9194 3295 9232 3364
rect 8787 3275 9232 3295
rect 9459 3326 9570 3341
rect 9459 3324 9501 3326
rect 9459 3304 9466 3324
rect 9485 3304 9501 3324
rect 9459 3296 9501 3304
rect 9529 3324 9570 3326
rect 9529 3304 9543 3324
rect 9562 3304 9570 3324
rect 9529 3296 9570 3304
rect 9459 3290 9570 3296
rect 9692 3301 9726 3364
rect 9844 3360 9882 3366
rect 9844 3342 9854 3360
rect 9872 3342 9882 3360
rect 10140 3358 10150 3376
rect 10168 3358 10178 3376
rect 10140 3352 10178 3358
rect 10296 3354 10330 3417
rect 10452 3422 10563 3428
rect 10452 3414 10493 3422
rect 10452 3394 10460 3414
rect 10479 3394 10493 3414
rect 10452 3392 10493 3394
rect 10521 3414 10563 3422
rect 10521 3394 10537 3414
rect 10556 3394 10563 3414
rect 10521 3392 10563 3394
rect 10452 3377 10563 3392
rect 10790 3423 11235 3443
rect 10790 3354 10828 3423
rect 11067 3422 11235 3423
rect 11313 3495 11395 3517
rect 11424 3495 11434 3522
rect 11462 3498 11469 3525
rect 11498 3517 11501 3525
rect 13496 3534 13607 3549
rect 13496 3532 13538 3534
rect 11498 3498 11563 3517
rect 11462 3495 11563 3498
rect 11313 3493 11563 3495
rect 11313 3414 11350 3493
rect 11391 3480 11501 3493
rect 11465 3424 11496 3425
rect 11313 3394 11322 3414
rect 11342 3394 11350 3414
rect 11313 3384 11350 3394
rect 11409 3414 11496 3424
rect 11409 3394 11418 3414
rect 11438 3394 11496 3414
rect 11409 3385 11496 3394
rect 11409 3384 11446 3385
rect 10140 3348 10177 3352
rect 10296 3343 10828 3354
rect 9844 3333 9882 3342
rect 9844 3301 9878 3333
rect 10295 3327 10828 3343
rect 11465 3332 11496 3385
rect 11526 3414 11563 3493
rect 11734 3503 12127 3510
rect 11734 3486 11742 3503
rect 11774 3490 12127 3503
rect 12147 3490 12150 3510
rect 13229 3505 13270 3514
rect 11774 3486 12150 3490
rect 11734 3485 12150 3486
rect 12824 3503 12992 3504
rect 13229 3503 13238 3505
rect 11734 3484 12075 3485
rect 11678 3424 11709 3425
rect 11526 3394 11535 3414
rect 11555 3394 11563 3414
rect 11526 3384 11563 3394
rect 11622 3417 11709 3424
rect 11622 3414 11683 3417
rect 11622 3394 11631 3414
rect 11651 3397 11683 3414
rect 11704 3397 11709 3417
rect 11651 3394 11709 3397
rect 11622 3387 11709 3394
rect 11734 3414 11771 3484
rect 12037 3483 12074 3484
rect 12824 3483 13238 3503
rect 13264 3483 13270 3505
rect 13496 3512 13503 3532
rect 13522 3512 13538 3532
rect 13496 3504 13538 3512
rect 13566 3532 13607 3534
rect 13566 3512 13580 3532
rect 13599 3512 13607 3532
rect 13566 3504 13607 3512
rect 13862 3508 13899 3509
rect 14165 3508 14202 3578
rect 14227 3598 14314 3605
rect 14227 3595 14285 3598
rect 14227 3575 14232 3595
rect 14253 3578 14285 3595
rect 14305 3578 14314 3598
rect 14253 3575 14314 3578
rect 14227 3568 14314 3575
rect 14373 3598 14410 3608
rect 14373 3578 14381 3598
rect 14401 3578 14410 3598
rect 14227 3567 14258 3568
rect 13861 3507 14202 3508
rect 13496 3498 13607 3504
rect 13786 3502 14202 3507
rect 12824 3477 13270 3483
rect 12824 3475 12992 3477
rect 11886 3424 11922 3425
rect 11734 3394 11743 3414
rect 11763 3394 11771 3414
rect 11622 3385 11678 3387
rect 11622 3384 11659 3385
rect 11734 3384 11771 3394
rect 11830 3414 11978 3424
rect 12078 3421 12174 3423
rect 11830 3394 11839 3414
rect 11859 3409 11949 3414
rect 11859 3394 11894 3409
rect 11830 3385 11894 3394
rect 11830 3384 11867 3385
rect 11886 3368 11894 3385
rect 11915 3394 11949 3409
rect 11969 3394 11978 3414
rect 11915 3385 11978 3394
rect 12036 3414 12174 3421
rect 12036 3394 12045 3414
rect 12065 3394 12174 3414
rect 12036 3385 12174 3394
rect 11915 3368 11922 3385
rect 11941 3384 11978 3385
rect 12037 3384 12074 3385
rect 11886 3333 11922 3368
rect 11357 3331 11398 3332
rect 10295 3326 10809 3327
rect 8787 3269 9231 3275
rect 8787 3267 8955 3269
rect 8627 3196 8631 3201
rect 8588 3193 8631 3196
rect 8521 3179 8631 3193
rect 7750 3165 7818 3174
rect 5972 3150 6008 3151
rect 5820 3120 5829 3140
rect 5849 3120 5857 3140
rect 5708 3111 5764 3113
rect 5708 3110 5745 3111
rect 5820 3110 5857 3120
rect 5916 3140 6064 3150
rect 6164 3147 6260 3149
rect 5916 3120 5925 3140
rect 5945 3120 6035 3140
rect 6055 3120 6064 3140
rect 5916 3111 6064 3120
rect 6122 3140 6260 3147
rect 6122 3120 6131 3140
rect 6151 3120 6260 3140
rect 7750 3136 7765 3165
rect 7813 3145 7818 3165
rect 7813 3136 7820 3145
rect 7750 3125 7820 3136
rect 6122 3111 6260 3120
rect 5916 3110 5953 3111
rect 5972 3059 6008 3111
rect 6027 3110 6064 3111
rect 6123 3110 6160 3111
rect 5443 3057 5484 3058
rect 5335 3050 5484 3057
rect 5335 3030 5453 3050
rect 5473 3030 5484 3050
rect 5335 3022 5484 3030
rect 5551 3054 5910 3058
rect 5551 3049 5873 3054
rect 5551 3025 5664 3049
rect 5688 3030 5873 3049
rect 5897 3030 5910 3054
rect 5688 3025 5910 3030
rect 5551 3022 5910 3025
rect 5972 3022 6007 3059
rect 6075 3056 6175 3059
rect 6075 3052 6142 3056
rect 6075 3026 6087 3052
rect 6113 3030 6142 3052
rect 6168 3030 6175 3056
rect 6113 3026 6175 3030
rect 6075 3022 6175 3026
rect 5551 3001 5582 3022
rect 5972 3001 6008 3022
rect 5394 3000 5431 3001
rect 5393 2991 5431 3000
rect 5393 2971 5402 2991
rect 5422 2971 5431 2991
rect 5393 2963 5431 2971
rect 5497 2995 5582 3001
rect 5607 3000 5644 3001
rect 5497 2975 5505 2995
rect 5525 2975 5582 2995
rect 5497 2967 5582 2975
rect 5606 2991 5644 3000
rect 5606 2971 5615 2991
rect 5635 2971 5644 2991
rect 5497 2966 5533 2967
rect 5606 2963 5644 2971
rect 5710 2995 5795 3001
rect 5815 3000 5852 3001
rect 5710 2975 5718 2995
rect 5738 2994 5795 2995
rect 5738 2975 5767 2994
rect 5710 2974 5767 2975
rect 5788 2974 5795 2994
rect 5710 2967 5795 2974
rect 5814 2991 5852 3000
rect 5814 2971 5823 2991
rect 5843 2971 5852 2991
rect 5710 2966 5746 2967
rect 5814 2963 5852 2971
rect 5918 2995 6062 3001
rect 5918 2975 5926 2995
rect 5946 2992 6034 2995
rect 5946 2975 5977 2992
rect 5918 2972 5977 2975
rect 6000 2975 6034 2992
rect 6054 2975 6062 2995
rect 6000 2972 6062 2975
rect 5918 2967 6062 2972
rect 5918 2966 5954 2967
rect 6026 2966 6062 2967
rect 6128 3000 6165 3001
rect 6128 2999 6166 3000
rect 6128 2991 6192 2999
rect 6128 2971 6137 2991
rect 6157 2977 6192 2991
rect 6212 2977 6215 2997
rect 6157 2972 6215 2977
rect 6157 2971 6192 2972
rect 5394 2934 5431 2963
rect 5395 2932 5431 2934
rect 5607 2932 5644 2963
rect 5395 2910 5644 2932
rect 5815 2931 5852 2963
rect 6128 2959 6192 2971
rect 6232 2933 6259 3111
rect 7759 3018 7820 3125
rect 8787 3089 8814 3267
rect 8854 3229 8918 3241
rect 9194 3237 9231 3269
rect 9402 3268 9651 3290
rect 9692 3269 9878 3301
rect 11249 3324 11398 3331
rect 11249 3304 11367 3324
rect 11387 3304 11398 3324
rect 11249 3296 11398 3304
rect 11465 3328 11824 3332
rect 11465 3323 11787 3328
rect 11465 3299 11578 3323
rect 11602 3304 11787 3323
rect 11811 3304 11824 3328
rect 11602 3299 11824 3304
rect 11465 3296 11824 3299
rect 11886 3296 11921 3333
rect 11989 3330 12089 3333
rect 11989 3326 12056 3330
rect 11989 3300 12001 3326
rect 12027 3304 12056 3326
rect 12082 3304 12089 3330
rect 12027 3300 12089 3304
rect 11989 3296 12089 3300
rect 10143 3285 10180 3286
rect 9706 3268 9878 3269
rect 9402 3237 9439 3268
rect 9615 3266 9651 3268
rect 9615 3237 9652 3266
rect 9844 3240 9878 3268
rect 10141 3277 10181 3285
rect 10141 3259 10152 3277
rect 10170 3259 10181 3277
rect 11465 3275 11496 3296
rect 11886 3275 11922 3296
rect 11308 3274 11345 3275
rect 8854 3228 8889 3229
rect 8831 3223 8889 3228
rect 8831 3203 8834 3223
rect 8854 3209 8889 3223
rect 8909 3209 8918 3229
rect 8854 3201 8918 3209
rect 8880 3200 8918 3201
rect 8881 3199 8918 3200
rect 8984 3233 9020 3234
rect 9092 3233 9128 3234
rect 8984 3226 9128 3233
rect 8984 3225 9044 3226
rect 8984 3205 8992 3225
rect 9012 3206 9044 3225
rect 9069 3225 9128 3226
rect 9069 3206 9100 3225
rect 9012 3205 9100 3206
rect 9120 3205 9128 3225
rect 8984 3199 9128 3205
rect 9194 3229 9232 3237
rect 9300 3233 9336 3234
rect 9194 3209 9203 3229
rect 9223 3209 9232 3229
rect 9194 3200 9232 3209
rect 9251 3226 9336 3233
rect 9251 3206 9258 3226
rect 9279 3225 9336 3226
rect 9279 3206 9308 3225
rect 9251 3205 9308 3206
rect 9328 3205 9336 3225
rect 9194 3199 9231 3200
rect 9251 3199 9336 3205
rect 9402 3229 9440 3237
rect 9513 3233 9549 3234
rect 9402 3209 9411 3229
rect 9431 3209 9440 3229
rect 9402 3200 9440 3209
rect 9464 3225 9549 3233
rect 9464 3205 9521 3225
rect 9541 3205 9549 3225
rect 9402 3199 9439 3200
rect 9464 3199 9549 3205
rect 9615 3229 9653 3237
rect 9615 3209 9624 3229
rect 9644 3209 9653 3229
rect 9615 3200 9653 3209
rect 9842 3230 9879 3240
rect 9842 3212 9852 3230
rect 9870 3212 9879 3230
rect 9842 3203 9879 3212
rect 10141 3211 10181 3259
rect 11307 3265 11345 3274
rect 11307 3245 11316 3265
rect 11336 3245 11345 3265
rect 11307 3237 11345 3245
rect 11411 3269 11496 3275
rect 11521 3274 11558 3275
rect 11411 3249 11419 3269
rect 11439 3249 11496 3269
rect 11411 3241 11496 3249
rect 11520 3265 11558 3274
rect 11520 3245 11529 3265
rect 11549 3245 11558 3265
rect 11411 3240 11447 3241
rect 11520 3237 11558 3245
rect 11624 3269 11709 3275
rect 11729 3274 11766 3275
rect 11624 3249 11632 3269
rect 11652 3268 11709 3269
rect 11652 3249 11681 3268
rect 11624 3248 11681 3249
rect 11702 3248 11709 3268
rect 11624 3241 11709 3248
rect 11728 3265 11766 3274
rect 11728 3245 11737 3265
rect 11757 3245 11766 3265
rect 11624 3240 11660 3241
rect 11728 3237 11766 3245
rect 11832 3269 11976 3275
rect 11832 3249 11840 3269
rect 11860 3249 11948 3269
rect 11968 3249 11976 3269
rect 11832 3241 11976 3249
rect 11832 3240 11868 3241
rect 11940 3240 11976 3241
rect 12042 3274 12079 3275
rect 12042 3273 12080 3274
rect 12042 3265 12106 3273
rect 12042 3245 12051 3265
rect 12071 3251 12106 3265
rect 12126 3251 12129 3271
rect 12071 3246 12129 3251
rect 12071 3245 12106 3246
rect 10452 3215 10562 3229
rect 10452 3212 10495 3215
rect 10141 3204 10266 3211
rect 10452 3207 10456 3212
rect 9844 3202 9878 3203
rect 9615 3199 9652 3200
rect 9038 3178 9074 3199
rect 9464 3178 9495 3199
rect 10141 3185 10233 3204
rect 10258 3185 10266 3204
rect 8871 3174 8971 3178
rect 8871 3170 8933 3174
rect 8871 3144 8878 3170
rect 8904 3148 8933 3170
rect 8959 3148 8971 3174
rect 8904 3144 8971 3148
rect 8871 3141 8971 3144
rect 9039 3141 9074 3178
rect 9136 3175 9495 3178
rect 9136 3170 9358 3175
rect 9136 3146 9149 3170
rect 9173 3151 9358 3170
rect 9382 3151 9495 3175
rect 9173 3146 9495 3151
rect 9136 3142 9495 3146
rect 9562 3170 9711 3178
rect 9562 3150 9573 3170
rect 9593 3150 9711 3170
rect 10141 3175 10266 3185
rect 10374 3185 10456 3207
rect 10485 3185 10495 3212
rect 10523 3188 10530 3215
rect 10559 3207 10562 3215
rect 11308 3208 11345 3237
rect 10559 3188 10624 3207
rect 11309 3206 11345 3208
rect 11521 3206 11558 3237
rect 11729 3210 11766 3237
rect 12042 3233 12106 3245
rect 10523 3185 10624 3188
rect 10374 3183 10624 3185
rect 10141 3155 10181 3175
rect 9562 3143 9711 3150
rect 10140 3146 10181 3155
rect 9562 3142 9603 3143
rect 8886 3089 8923 3090
rect 8982 3089 9019 3090
rect 9038 3089 9074 3141
rect 9093 3089 9130 3090
rect 8786 3080 8924 3089
rect 7750 3017 7820 3018
rect 8411 3046 8522 3061
rect 8786 3060 8895 3080
rect 8915 3060 8924 3080
rect 8786 3053 8924 3060
rect 8982 3080 9130 3089
rect 8982 3060 8991 3080
rect 9011 3060 9101 3080
rect 9121 3060 9130 3080
rect 8786 3051 8882 3053
rect 8982 3050 9130 3060
rect 9189 3080 9226 3090
rect 9301 3089 9338 3090
rect 9282 3087 9338 3089
rect 9189 3060 9197 3080
rect 9217 3060 9226 3080
rect 9038 3049 9074 3050
rect 8411 3044 8453 3046
rect 8411 3024 8418 3044
rect 8437 3024 8453 3044
rect 7750 3016 7858 3017
rect 8411 3016 8453 3024
rect 8481 3044 8522 3046
rect 8481 3024 8495 3044
rect 8514 3024 8522 3044
rect 8481 3016 8522 3024
rect 7739 3015 7907 3016
rect 6526 2982 6636 2996
rect 6526 2979 6569 2982
rect 6526 2974 6530 2979
rect 6091 2931 6259 2933
rect 5815 2928 6259 2931
rect 5476 2904 5587 2910
rect 5476 2896 5517 2904
rect 5165 2841 5204 2885
rect 5476 2876 5484 2896
rect 5503 2876 5517 2896
rect 5476 2874 5517 2876
rect 5545 2896 5587 2904
rect 5545 2876 5561 2896
rect 5580 2876 5587 2896
rect 5545 2874 5587 2876
rect 5476 2860 5587 2874
rect 5813 2905 6259 2928
rect 3458 2821 3499 2822
rect 2782 2768 2819 2769
rect 2878 2768 2915 2769
rect 2934 2768 2970 2820
rect 2989 2768 3026 2769
rect 2682 2759 2820 2768
rect 2682 2739 2791 2759
rect 2811 2739 2820 2759
rect 2682 2732 2820 2739
rect 2878 2759 3026 2768
rect 2878 2739 2887 2759
rect 2907 2739 2997 2759
rect 3017 2739 3026 2759
rect 2682 2730 2778 2732
rect 2878 2729 3026 2739
rect 3085 2759 3122 2769
rect 3197 2768 3234 2769
rect 3178 2766 3234 2768
rect 3085 2739 3093 2759
rect 3113 2739 3122 2759
rect 2934 2728 2970 2729
rect 2782 2669 2819 2670
rect 3085 2669 3122 2739
rect 3147 2759 3234 2766
rect 3147 2756 3205 2759
rect 3147 2736 3152 2756
rect 3173 2739 3205 2756
rect 3225 2739 3234 2759
rect 3173 2736 3234 2739
rect 3147 2729 3234 2736
rect 3293 2759 3330 2769
rect 3293 2739 3301 2759
rect 3321 2739 3330 2759
rect 3147 2728 3178 2729
rect 2781 2668 3122 2669
rect 2706 2663 3122 2668
rect 2706 2643 2709 2663
rect 2729 2643 3122 2663
rect 3293 2660 3330 2739
rect 3360 2768 3391 2821
rect 4140 2793 4826 2826
rect 3410 2768 3447 2769
rect 3360 2759 3447 2768
rect 3360 2739 3418 2759
rect 3438 2739 3447 2759
rect 3360 2729 3447 2739
rect 3506 2759 3543 2769
rect 3506 2739 3514 2759
rect 3534 2739 3543 2759
rect 3360 2728 3391 2729
rect 3355 2660 3465 2673
rect 3506 2660 3543 2739
rect 3293 2658 3543 2660
rect 3293 2655 3394 2658
rect 3293 2636 3358 2655
rect 2173 2623 2252 2631
rect 2084 2621 2252 2623
rect 1808 2614 2252 2621
rect 3355 2628 3358 2636
rect 3387 2628 3394 2655
rect 3422 2631 3432 2658
rect 3461 2636 3543 2658
rect 3732 2705 3900 2706
rect 4140 2705 4178 2793
rect 4439 2791 4486 2793
rect 4786 2769 4826 2793
rect 5165 2817 5205 2841
rect 5505 2817 5552 2819
rect 5813 2817 5851 2905
rect 6091 2904 6259 2905
rect 6448 2952 6530 2974
rect 6559 2952 6569 2979
rect 6597 2955 6604 2982
rect 6633 2974 6636 2982
rect 7739 2989 8183 3015
rect 8411 3010 8522 3016
rect 7739 2987 7907 2989
rect 7739 2985 7858 2987
rect 6633 2955 6698 2974
rect 6597 2952 6698 2955
rect 6448 2950 6698 2952
rect 6448 2871 6485 2950
rect 6526 2937 6636 2950
rect 6600 2881 6631 2882
rect 6448 2851 6457 2871
rect 6477 2851 6485 2871
rect 6448 2841 6485 2851
rect 6544 2871 6631 2881
rect 6544 2851 6553 2871
rect 6573 2851 6631 2871
rect 6544 2842 6631 2851
rect 6544 2841 6581 2842
rect 5165 2784 5851 2817
rect 6600 2789 6631 2842
rect 6661 2871 6698 2950
rect 6869 2969 6901 2981
rect 6869 2949 6871 2969
rect 6892 2967 6901 2969
rect 6892 2965 7244 2967
rect 6892 2949 7262 2965
rect 6869 2947 7262 2949
rect 7282 2947 7285 2965
rect 6869 2942 7285 2947
rect 6869 2941 7210 2942
rect 6813 2881 6844 2882
rect 6661 2851 6670 2871
rect 6690 2851 6698 2871
rect 6661 2841 6698 2851
rect 6757 2874 6844 2881
rect 6757 2871 6818 2874
rect 6757 2851 6766 2871
rect 6786 2854 6818 2871
rect 6839 2854 6844 2874
rect 6786 2851 6844 2854
rect 6757 2844 6844 2851
rect 6869 2871 6906 2941
rect 7172 2940 7209 2941
rect 7021 2881 7057 2882
rect 6869 2851 6878 2871
rect 6898 2851 6906 2871
rect 6757 2842 6813 2844
rect 6757 2841 6794 2842
rect 6869 2841 6906 2851
rect 6965 2871 7113 2881
rect 7213 2878 7309 2880
rect 6965 2851 6974 2871
rect 6994 2862 7084 2871
rect 6994 2851 7025 2862
rect 6965 2842 7025 2851
rect 6965 2841 7002 2842
rect 7021 2830 7025 2842
rect 7052 2851 7084 2862
rect 7104 2851 7113 2871
rect 7052 2842 7113 2851
rect 7171 2871 7309 2878
rect 7171 2851 7180 2871
rect 7200 2851 7309 2871
rect 7171 2842 7309 2851
rect 7052 2830 7057 2842
rect 7076 2841 7113 2842
rect 7172 2841 7209 2842
rect 7021 2790 7057 2830
rect 6492 2788 6533 2789
rect 3732 2682 4178 2705
rect 4404 2736 4515 2750
rect 4404 2734 4446 2736
rect 4404 2714 4411 2734
rect 4430 2714 4446 2734
rect 4404 2706 4446 2714
rect 4474 2734 4515 2736
rect 4474 2714 4488 2734
rect 4507 2714 4515 2734
rect 4787 2725 4826 2769
rect 4474 2706 4515 2714
rect 4404 2700 4515 2706
rect 3732 2679 4176 2682
rect 3732 2677 3900 2679
rect 3461 2631 3465 2636
rect 3422 2628 3465 2631
rect 3355 2614 3465 2628
rect 1469 2594 1580 2600
rect 1808 2595 2178 2614
rect 2084 2594 2178 2595
rect 1469 2586 1510 2594
rect 1469 2566 1477 2586
rect 1496 2566 1510 2586
rect 1469 2564 1510 2566
rect 1538 2586 1580 2594
rect 1538 2566 1554 2586
rect 1573 2566 1580 2586
rect 2173 2585 2178 2594
rect 2226 2594 2252 2614
rect 2226 2585 2243 2594
rect 2173 2576 2243 2585
rect 1538 2564 1580 2566
rect 917 2560 953 2561
rect 765 2530 774 2550
rect 794 2530 802 2550
rect 653 2521 709 2523
rect 653 2520 690 2521
rect 765 2520 802 2530
rect 861 2550 1009 2560
rect 1109 2557 1205 2559
rect 861 2530 870 2550
rect 890 2530 980 2550
rect 1000 2530 1009 2550
rect 861 2521 1009 2530
rect 1067 2550 1205 2557
rect 1067 2530 1076 2550
rect 1096 2530 1205 2550
rect 1469 2549 1580 2564
rect 1067 2521 1205 2530
rect 861 2520 898 2521
rect 917 2469 953 2521
rect 972 2520 1009 2521
rect 1068 2520 1105 2521
rect 388 2467 429 2468
rect 280 2460 429 2467
rect 280 2440 398 2460
rect 418 2440 429 2460
rect 280 2432 429 2440
rect 496 2464 855 2468
rect 496 2459 818 2464
rect 496 2435 609 2459
rect 633 2440 818 2459
rect 842 2440 855 2464
rect 633 2435 855 2440
rect 496 2432 855 2435
rect 917 2432 952 2469
rect 1020 2466 1120 2469
rect 1020 2462 1087 2466
rect 1020 2436 1032 2462
rect 1058 2440 1087 2462
rect 1113 2440 1120 2466
rect 1058 2436 1120 2440
rect 1020 2432 1120 2436
rect 496 2411 527 2432
rect 917 2411 953 2432
rect 339 2410 376 2411
rect 113 2407 147 2408
rect 112 2398 149 2407
rect 112 2380 121 2398
rect 139 2380 149 2398
rect 112 2370 149 2380
rect 338 2401 376 2410
rect 338 2381 347 2401
rect 367 2381 376 2401
rect 338 2373 376 2381
rect 442 2405 527 2411
rect 552 2410 589 2411
rect 442 2385 450 2405
rect 470 2385 527 2405
rect 442 2377 527 2385
rect 551 2401 589 2410
rect 551 2381 560 2401
rect 580 2381 589 2401
rect 442 2376 478 2377
rect 551 2373 589 2381
rect 655 2405 740 2411
rect 760 2410 797 2411
rect 655 2385 663 2405
rect 683 2404 740 2405
rect 683 2385 712 2404
rect 655 2384 712 2385
rect 733 2384 740 2404
rect 655 2377 740 2384
rect 759 2401 797 2410
rect 759 2381 768 2401
rect 788 2381 797 2401
rect 655 2376 691 2377
rect 759 2373 797 2381
rect 863 2405 1007 2411
rect 863 2385 871 2405
rect 891 2404 979 2405
rect 891 2385 922 2404
rect 863 2384 922 2385
rect 947 2385 979 2404
rect 999 2385 1007 2405
rect 947 2384 1007 2385
rect 863 2377 1007 2384
rect 863 2376 899 2377
rect 971 2376 1007 2377
rect 1073 2410 1110 2411
rect 1073 2409 1111 2410
rect 1073 2401 1137 2409
rect 1073 2381 1082 2401
rect 1102 2387 1137 2401
rect 1157 2387 1160 2407
rect 1102 2382 1160 2387
rect 1102 2381 1137 2382
rect 113 2342 147 2370
rect 339 2344 376 2373
rect 340 2342 376 2344
rect 552 2342 589 2373
rect 113 2341 285 2342
rect 113 2309 299 2341
rect 340 2320 589 2342
rect 760 2341 797 2373
rect 1073 2369 1137 2381
rect 1177 2343 1204 2521
rect 3732 2499 3759 2677
rect 3799 2639 3863 2651
rect 4139 2647 4176 2679
rect 4347 2678 4596 2700
rect 4347 2647 4384 2678
rect 4560 2676 4596 2678
rect 4560 2647 4597 2676
rect 3799 2638 3834 2639
rect 3776 2633 3834 2638
rect 3776 2613 3779 2633
rect 3799 2619 3834 2633
rect 3854 2619 3863 2639
rect 3799 2611 3863 2619
rect 3825 2610 3863 2611
rect 3826 2609 3863 2610
rect 3929 2643 3965 2644
rect 4037 2643 4073 2644
rect 3929 2638 4073 2643
rect 3929 2635 3991 2638
rect 3929 2615 3937 2635
rect 3957 2618 3991 2635
rect 4014 2635 4073 2638
rect 4014 2618 4045 2635
rect 3957 2615 4045 2618
rect 4065 2615 4073 2635
rect 3929 2609 4073 2615
rect 4139 2639 4177 2647
rect 4245 2643 4281 2644
rect 4139 2619 4148 2639
rect 4168 2619 4177 2639
rect 4139 2610 4177 2619
rect 4196 2636 4281 2643
rect 4196 2616 4203 2636
rect 4224 2635 4281 2636
rect 4224 2616 4253 2635
rect 4196 2615 4253 2616
rect 4273 2615 4281 2635
rect 4139 2609 4176 2610
rect 4196 2609 4281 2615
rect 4347 2639 4385 2647
rect 4458 2643 4494 2644
rect 4347 2619 4356 2639
rect 4376 2619 4385 2639
rect 4347 2610 4385 2619
rect 4409 2635 4494 2643
rect 4409 2615 4466 2635
rect 4486 2615 4494 2635
rect 4347 2609 4384 2610
rect 4409 2609 4494 2615
rect 4560 2639 4598 2647
rect 4560 2619 4569 2639
rect 4589 2619 4598 2639
rect 4560 2610 4598 2619
rect 4560 2609 4597 2610
rect 3983 2588 4019 2609
rect 4409 2588 4440 2609
rect 3816 2584 3916 2588
rect 3816 2580 3878 2584
rect 3816 2554 3823 2580
rect 3849 2558 3878 2580
rect 3904 2558 3916 2584
rect 3849 2554 3916 2558
rect 3816 2551 3916 2554
rect 3984 2551 4019 2588
rect 4081 2585 4440 2588
rect 4081 2580 4303 2585
rect 4081 2556 4094 2580
rect 4118 2561 4303 2580
rect 4327 2561 4440 2585
rect 4118 2556 4440 2561
rect 4081 2552 4440 2556
rect 4507 2580 4656 2588
rect 4507 2560 4518 2580
rect 4538 2560 4656 2580
rect 4507 2553 4656 2560
rect 4507 2552 4548 2553
rect 3831 2499 3868 2500
rect 3927 2499 3964 2500
rect 3983 2499 4019 2551
rect 4038 2499 4075 2500
rect 3731 2490 3869 2499
rect 3731 2470 3840 2490
rect 3860 2470 3869 2490
rect 3731 2463 3869 2470
rect 3927 2490 4075 2499
rect 3927 2470 3936 2490
rect 3956 2470 4046 2490
rect 4066 2470 4075 2490
rect 3731 2461 3827 2463
rect 3927 2460 4075 2470
rect 4134 2490 4171 2500
rect 4246 2499 4283 2500
rect 4227 2497 4283 2499
rect 4134 2470 4142 2490
rect 4162 2470 4171 2490
rect 3983 2459 4019 2460
rect 1360 2417 1470 2431
rect 1360 2414 1403 2417
rect 1360 2409 1364 2414
rect 1036 2341 1204 2343
rect 760 2335 1204 2341
rect 113 2277 147 2309
rect 109 2268 147 2277
rect 109 2250 119 2268
rect 137 2250 147 2268
rect 109 2244 147 2250
rect 265 2246 299 2309
rect 421 2314 532 2320
rect 421 2306 462 2314
rect 421 2286 429 2306
rect 448 2286 462 2306
rect 421 2284 462 2286
rect 490 2306 532 2314
rect 490 2286 506 2306
rect 525 2286 532 2306
rect 490 2284 532 2286
rect 421 2269 532 2284
rect 759 2315 1204 2335
rect 759 2246 797 2315
rect 1036 2314 1204 2315
rect 1282 2387 1364 2409
rect 1393 2387 1403 2414
rect 1431 2390 1438 2417
rect 1467 2409 1470 2417
rect 3465 2426 3576 2441
rect 3465 2424 3507 2426
rect 1467 2390 1532 2409
rect 1431 2387 1532 2390
rect 1282 2385 1532 2387
rect 1282 2306 1319 2385
rect 1360 2372 1470 2385
rect 1434 2316 1465 2317
rect 1282 2286 1291 2306
rect 1311 2286 1319 2306
rect 1282 2276 1319 2286
rect 1378 2306 1465 2316
rect 1378 2286 1387 2306
rect 1407 2286 1465 2306
rect 1378 2277 1465 2286
rect 1378 2276 1415 2277
rect 109 2240 146 2244
rect 265 2235 797 2246
rect 264 2219 797 2235
rect 1434 2224 1465 2277
rect 1495 2306 1532 2385
rect 1703 2382 2096 2402
rect 2116 2382 2119 2402
rect 3198 2397 3239 2406
rect 1703 2377 2119 2382
rect 2793 2395 2961 2396
rect 3198 2395 3207 2397
rect 1703 2376 2044 2377
rect 1647 2316 1678 2317
rect 1495 2286 1504 2306
rect 1524 2286 1532 2306
rect 1495 2276 1532 2286
rect 1591 2309 1678 2316
rect 1591 2306 1652 2309
rect 1591 2286 1600 2306
rect 1620 2289 1652 2306
rect 1673 2289 1678 2309
rect 1620 2286 1678 2289
rect 1591 2279 1678 2286
rect 1703 2306 1740 2376
rect 2006 2375 2043 2376
rect 2793 2375 3207 2395
rect 3233 2375 3239 2397
rect 3465 2404 3472 2424
rect 3491 2404 3507 2424
rect 3465 2396 3507 2404
rect 3535 2424 3576 2426
rect 3535 2404 3549 2424
rect 3568 2404 3576 2424
rect 3535 2396 3576 2404
rect 3831 2400 3868 2401
rect 4134 2400 4171 2470
rect 4196 2490 4283 2497
rect 4196 2487 4254 2490
rect 4196 2467 4201 2487
rect 4222 2470 4254 2487
rect 4274 2470 4283 2490
rect 4222 2467 4283 2470
rect 4196 2460 4283 2467
rect 4342 2490 4379 2500
rect 4342 2470 4350 2490
rect 4370 2470 4379 2490
rect 4196 2459 4227 2460
rect 3830 2399 4171 2400
rect 3465 2390 3576 2396
rect 3755 2394 4171 2399
rect 2793 2369 3239 2375
rect 2793 2367 2961 2369
rect 1855 2316 1891 2317
rect 1703 2286 1712 2306
rect 1732 2286 1740 2306
rect 1591 2277 1647 2279
rect 1591 2276 1628 2277
rect 1703 2276 1740 2286
rect 1799 2306 1947 2316
rect 2047 2313 2143 2315
rect 1799 2286 1808 2306
rect 1828 2286 1918 2306
rect 1938 2286 1947 2306
rect 1799 2277 1947 2286
rect 2005 2306 2143 2313
rect 2005 2286 2014 2306
rect 2034 2286 2143 2306
rect 2005 2277 2143 2286
rect 1799 2276 1836 2277
rect 1855 2225 1891 2277
rect 1910 2276 1947 2277
rect 2006 2276 2043 2277
rect 1326 2223 1367 2224
rect 264 2218 778 2219
rect 1218 2216 1367 2223
rect 1218 2196 1336 2216
rect 1356 2196 1367 2216
rect 1218 2188 1367 2196
rect 1434 2220 1793 2224
rect 1434 2215 1756 2220
rect 1434 2191 1547 2215
rect 1571 2196 1756 2215
rect 1780 2196 1793 2220
rect 1571 2191 1793 2196
rect 1434 2188 1793 2191
rect 1855 2188 1890 2225
rect 1958 2222 2058 2225
rect 1958 2218 2025 2222
rect 1958 2192 1970 2218
rect 1996 2196 2025 2218
rect 2051 2196 2058 2222
rect 1996 2192 2058 2196
rect 1958 2188 2058 2192
rect 112 2177 149 2178
rect 110 2169 150 2177
rect 110 2151 121 2169
rect 139 2151 150 2169
rect 1434 2167 1465 2188
rect 1855 2167 1891 2188
rect 1277 2166 1314 2167
rect 110 2103 150 2151
rect 1276 2157 1314 2166
rect 1276 2137 1285 2157
rect 1305 2137 1314 2157
rect 1276 2129 1314 2137
rect 1380 2161 1465 2167
rect 1490 2166 1527 2167
rect 1380 2141 1388 2161
rect 1408 2141 1465 2161
rect 1380 2133 1465 2141
rect 1489 2157 1527 2166
rect 1489 2137 1498 2157
rect 1518 2137 1527 2157
rect 1380 2132 1416 2133
rect 1489 2129 1527 2137
rect 1593 2161 1678 2167
rect 1698 2166 1735 2167
rect 1593 2141 1601 2161
rect 1621 2160 1678 2161
rect 1621 2141 1650 2160
rect 1593 2140 1650 2141
rect 1671 2140 1678 2160
rect 1593 2133 1678 2140
rect 1697 2157 1735 2166
rect 1697 2137 1706 2157
rect 1726 2137 1735 2157
rect 1593 2132 1629 2133
rect 1697 2129 1735 2137
rect 1801 2161 1945 2167
rect 1801 2141 1809 2161
rect 1829 2144 1865 2161
rect 1885 2144 1917 2161
rect 1829 2141 1917 2144
rect 1937 2141 1945 2161
rect 1801 2133 1945 2141
rect 1801 2132 1837 2133
rect 1909 2132 1945 2133
rect 2011 2166 2048 2167
rect 2011 2165 2049 2166
rect 2011 2157 2075 2165
rect 2011 2137 2020 2157
rect 2040 2143 2075 2157
rect 2095 2143 2098 2163
rect 2040 2138 2098 2143
rect 2040 2137 2075 2138
rect 421 2107 531 2121
rect 421 2104 464 2107
rect 110 2096 235 2103
rect 421 2099 425 2104
rect 110 2077 202 2096
rect 227 2077 235 2096
rect 110 2067 235 2077
rect 343 2077 425 2099
rect 454 2077 464 2104
rect 492 2080 499 2107
rect 528 2099 531 2107
rect 1277 2100 1314 2129
rect 528 2080 593 2099
rect 1278 2098 1314 2100
rect 1490 2098 1527 2129
rect 1698 2102 1735 2129
rect 2011 2125 2075 2137
rect 492 2077 593 2080
rect 343 2075 593 2077
rect 110 2047 150 2067
rect 109 2038 150 2047
rect 109 2020 119 2038
rect 137 2020 150 2038
rect 109 2011 150 2020
rect 109 2010 146 2011
rect 343 1996 380 2075
rect 421 2062 531 2075
rect 495 2006 526 2007
rect 343 1976 352 1996
rect 372 1976 380 1996
rect 343 1966 380 1976
rect 439 1996 526 2006
rect 439 1976 448 1996
rect 468 1976 526 1996
rect 439 1967 526 1976
rect 439 1966 476 1967
rect 112 1944 149 1948
rect 109 1939 149 1944
rect 109 1921 121 1939
rect 139 1921 149 1939
rect 109 1741 149 1921
rect 495 1914 526 1967
rect 556 1996 593 2075
rect 764 2072 1157 2092
rect 1177 2072 1180 2092
rect 1278 2076 1527 2098
rect 1696 2097 1737 2102
rect 2115 2099 2142 2277
rect 2793 2189 2820 2367
rect 3198 2364 3239 2369
rect 3408 2368 3657 2390
rect 3755 2374 3758 2394
rect 3778 2374 4171 2394
rect 4342 2391 4379 2470
rect 4409 2499 4440 2552
rect 4786 2545 4826 2725
rect 5164 2727 5203 2784
rect 5813 2782 5851 2784
rect 6384 2781 6533 2788
rect 6384 2761 6502 2781
rect 6522 2761 6533 2781
rect 6384 2753 6533 2761
rect 6600 2785 6959 2789
rect 6600 2780 6922 2785
rect 6600 2756 6713 2780
rect 6737 2761 6922 2780
rect 6946 2761 6959 2785
rect 6737 2756 6959 2761
rect 6600 2753 6959 2756
rect 7021 2753 7056 2790
rect 7124 2787 7224 2790
rect 7124 2783 7191 2787
rect 7124 2757 7136 2783
rect 7162 2761 7191 2783
rect 7217 2761 7224 2787
rect 7162 2757 7224 2761
rect 7124 2753 7224 2757
rect 6600 2732 6631 2753
rect 7021 2732 7057 2753
rect 6443 2731 6480 2732
rect 5164 2725 5212 2727
rect 5164 2707 5175 2725
rect 5193 2707 5212 2725
rect 6442 2722 6480 2731
rect 5164 2698 5212 2707
rect 5165 2697 5212 2698
rect 5478 2702 5588 2716
rect 5478 2699 5521 2702
rect 5478 2694 5482 2699
rect 5400 2672 5482 2694
rect 5511 2672 5521 2699
rect 5549 2675 5556 2702
rect 5585 2694 5588 2702
rect 6442 2702 6451 2722
rect 6471 2702 6480 2722
rect 6442 2694 6480 2702
rect 6546 2726 6631 2732
rect 6656 2731 6693 2732
rect 6546 2706 6554 2726
rect 6574 2706 6631 2726
rect 6546 2698 6631 2706
rect 6655 2722 6693 2731
rect 6655 2702 6664 2722
rect 6684 2702 6693 2722
rect 6546 2697 6582 2698
rect 6655 2694 6693 2702
rect 6759 2726 6844 2732
rect 6864 2731 6901 2732
rect 6759 2706 6767 2726
rect 6787 2725 6844 2726
rect 6787 2706 6816 2725
rect 6759 2705 6816 2706
rect 6837 2705 6844 2725
rect 6759 2698 6844 2705
rect 6863 2722 6901 2731
rect 6863 2702 6872 2722
rect 6892 2702 6901 2722
rect 6759 2697 6795 2698
rect 6863 2694 6901 2702
rect 6967 2726 7111 2732
rect 6967 2706 6975 2726
rect 6995 2706 7083 2726
rect 7103 2706 7111 2726
rect 6967 2698 7111 2706
rect 6967 2697 7003 2698
rect 7075 2697 7111 2698
rect 7177 2731 7214 2732
rect 7177 2730 7215 2731
rect 7177 2722 7241 2730
rect 7177 2702 7186 2722
rect 7206 2708 7241 2722
rect 7261 2708 7264 2728
rect 7206 2703 7264 2708
rect 7206 2702 7241 2703
rect 5585 2675 5650 2694
rect 5549 2672 5650 2675
rect 5400 2670 5650 2672
rect 5168 2634 5205 2635
rect 4786 2527 4796 2545
rect 4814 2527 4826 2545
rect 4786 2522 4826 2527
rect 5164 2631 5205 2634
rect 5164 2626 5206 2631
rect 5164 2608 5177 2626
rect 5195 2608 5206 2626
rect 5164 2594 5206 2608
rect 5244 2594 5291 2598
rect 5164 2588 5291 2594
rect 5164 2559 5252 2588
rect 5281 2559 5291 2588
rect 5400 2591 5437 2670
rect 5478 2657 5588 2670
rect 5552 2601 5583 2602
rect 5400 2571 5409 2591
rect 5429 2571 5437 2591
rect 5400 2561 5437 2571
rect 5496 2591 5583 2601
rect 5496 2571 5505 2591
rect 5525 2571 5583 2591
rect 5496 2562 5583 2571
rect 5496 2561 5533 2562
rect 5164 2555 5291 2559
rect 5164 2538 5203 2555
rect 5244 2554 5291 2555
rect 4786 2518 4823 2522
rect 5164 2520 5175 2538
rect 5193 2520 5203 2538
rect 5164 2511 5203 2520
rect 5165 2510 5202 2511
rect 5552 2509 5583 2562
rect 5613 2591 5650 2670
rect 5821 2667 6214 2687
rect 6234 2667 6237 2687
rect 5821 2662 6237 2667
rect 6443 2665 6480 2694
rect 6444 2663 6480 2665
rect 6656 2663 6693 2694
rect 5821 2661 6162 2662
rect 5765 2601 5796 2602
rect 5613 2571 5622 2591
rect 5642 2571 5650 2591
rect 5613 2561 5650 2571
rect 5709 2594 5796 2601
rect 5709 2591 5770 2594
rect 5709 2571 5718 2591
rect 5738 2574 5770 2591
rect 5791 2574 5796 2594
rect 5738 2571 5796 2574
rect 5709 2564 5796 2571
rect 5821 2591 5858 2661
rect 6124 2660 6161 2661
rect 6444 2641 6693 2663
rect 6864 2662 6901 2694
rect 7177 2690 7241 2702
rect 7281 2672 7308 2842
rect 7739 2809 7766 2985
rect 7806 2949 7870 2961
rect 8146 2957 8183 2989
rect 8354 2988 8603 3010
rect 8886 2990 8923 2991
rect 9189 2990 9226 3060
rect 9251 3080 9338 3087
rect 9251 3077 9309 3080
rect 9251 3057 9256 3077
rect 9277 3060 9309 3077
rect 9329 3060 9338 3080
rect 9277 3057 9338 3060
rect 9251 3050 9338 3057
rect 9397 3080 9434 3090
rect 9397 3060 9405 3080
rect 9425 3060 9434 3080
rect 9251 3049 9282 3050
rect 8885 2989 9226 2990
rect 8354 2957 8391 2988
rect 8567 2986 8603 2988
rect 8567 2957 8604 2986
rect 8810 2984 9226 2989
rect 8810 2964 8813 2984
rect 8833 2964 9226 2984
rect 9397 2981 9434 3060
rect 9464 3089 9495 3142
rect 9845 3140 9882 3141
rect 9844 3131 9883 3140
rect 9844 3113 9854 3131
rect 9872 3113 9883 3131
rect 10140 3128 10150 3146
rect 10168 3128 10181 3146
rect 10140 3119 10181 3128
rect 10140 3118 10177 3119
rect 9756 3096 9803 3097
rect 9844 3096 9883 3113
rect 9756 3092 9883 3096
rect 9514 3089 9551 3090
rect 9464 3080 9551 3089
rect 9464 3060 9522 3080
rect 9542 3060 9551 3080
rect 9464 3050 9551 3060
rect 9610 3080 9647 3090
rect 9610 3060 9618 3080
rect 9638 3060 9647 3080
rect 9464 3049 9495 3050
rect 9459 2981 9569 2994
rect 9610 2981 9647 3060
rect 9756 3063 9766 3092
rect 9795 3063 9883 3092
rect 10374 3104 10411 3183
rect 10452 3170 10562 3183
rect 10526 3114 10557 3115
rect 10374 3084 10383 3104
rect 10403 3084 10411 3104
rect 10374 3074 10411 3084
rect 10470 3104 10557 3114
rect 10470 3084 10479 3104
rect 10499 3084 10557 3104
rect 10470 3075 10557 3084
rect 10470 3074 10507 3075
rect 9756 3057 9883 3063
rect 9756 3053 9803 3057
rect 9841 3043 9883 3057
rect 10143 3052 10180 3056
rect 9841 3025 9852 3043
rect 9870 3025 9883 3043
rect 9841 3020 9883 3025
rect 9842 3017 9883 3020
rect 10140 3047 10180 3052
rect 10140 3029 10152 3047
rect 10170 3029 10180 3047
rect 9842 3016 9879 3017
rect 9397 2979 9647 2981
rect 9397 2976 9498 2979
rect 9397 2957 9462 2976
rect 7806 2948 7841 2949
rect 7783 2943 7841 2948
rect 7783 2923 7786 2943
rect 7806 2929 7841 2943
rect 7861 2929 7870 2949
rect 7806 2921 7870 2929
rect 7832 2920 7870 2921
rect 7833 2919 7870 2920
rect 7936 2953 7972 2954
rect 8044 2953 8080 2954
rect 7936 2946 8080 2953
rect 7936 2945 7994 2946
rect 7936 2925 7944 2945
rect 7964 2927 7994 2945
rect 8023 2945 8080 2946
rect 8023 2927 8052 2945
rect 7964 2925 8052 2927
rect 8072 2925 8080 2945
rect 7936 2919 8080 2925
rect 8146 2949 8184 2957
rect 8252 2953 8288 2954
rect 8146 2929 8155 2949
rect 8175 2929 8184 2949
rect 8146 2920 8184 2929
rect 8203 2946 8288 2953
rect 8203 2926 8210 2946
rect 8231 2945 8288 2946
rect 8231 2926 8260 2945
rect 8203 2925 8260 2926
rect 8280 2925 8288 2945
rect 8146 2919 8183 2920
rect 8203 2919 8288 2925
rect 8354 2949 8392 2957
rect 8465 2953 8501 2954
rect 8354 2929 8363 2949
rect 8383 2929 8392 2949
rect 8354 2920 8392 2929
rect 8416 2945 8501 2953
rect 8416 2925 8473 2945
rect 8493 2925 8501 2945
rect 8354 2919 8391 2920
rect 8416 2919 8501 2925
rect 8567 2949 8605 2957
rect 8567 2929 8576 2949
rect 8596 2929 8605 2949
rect 9459 2949 9462 2957
rect 9491 2949 9498 2976
rect 9526 2952 9536 2979
rect 9565 2957 9647 2979
rect 9565 2952 9569 2957
rect 9526 2949 9569 2952
rect 9459 2935 9569 2949
rect 9835 2953 9882 2954
rect 9835 2944 9883 2953
rect 8567 2920 8605 2929
rect 9835 2926 9854 2944
rect 9872 2926 9883 2944
rect 9835 2924 9883 2926
rect 8567 2919 8604 2920
rect 7990 2898 8026 2919
rect 8416 2898 8447 2919
rect 7823 2894 7923 2898
rect 7823 2890 7885 2894
rect 7823 2864 7830 2890
rect 7856 2868 7885 2890
rect 7911 2868 7923 2894
rect 7856 2864 7923 2868
rect 7823 2861 7923 2864
rect 7991 2861 8026 2898
rect 8088 2895 8447 2898
rect 8088 2890 8310 2895
rect 8088 2866 8101 2890
rect 8125 2871 8310 2890
rect 8334 2871 8447 2895
rect 8125 2866 8447 2871
rect 8088 2862 8447 2866
rect 8514 2890 8663 2898
rect 8514 2870 8525 2890
rect 8545 2870 8663 2890
rect 8514 2863 8663 2870
rect 9196 2867 9234 2869
rect 9844 2867 9883 2924
rect 8514 2862 8555 2863
rect 7838 2809 7875 2810
rect 7934 2809 7971 2810
rect 7990 2809 8026 2861
rect 8045 2809 8082 2810
rect 7738 2800 7876 2809
rect 7738 2780 7847 2800
rect 7867 2780 7876 2800
rect 7738 2773 7876 2780
rect 7934 2800 8082 2809
rect 7934 2780 7943 2800
rect 7963 2780 8053 2800
rect 8073 2780 8082 2800
rect 7738 2771 7834 2773
rect 7934 2770 8082 2780
rect 8141 2800 8178 2810
rect 8253 2809 8290 2810
rect 8234 2807 8290 2809
rect 8141 2780 8149 2800
rect 8169 2780 8178 2800
rect 7990 2769 8026 2770
rect 7838 2710 7875 2711
rect 8141 2710 8178 2780
rect 8203 2800 8290 2807
rect 8203 2797 8261 2800
rect 8203 2777 8208 2797
rect 8229 2780 8261 2797
rect 8281 2780 8290 2800
rect 8229 2777 8290 2780
rect 8203 2770 8290 2777
rect 8349 2800 8386 2810
rect 8349 2780 8357 2800
rect 8377 2780 8386 2800
rect 8203 2769 8234 2770
rect 7837 2709 8178 2710
rect 7762 2704 8178 2709
rect 7762 2684 7765 2704
rect 7785 2684 8178 2704
rect 8349 2701 8386 2780
rect 8416 2809 8447 2862
rect 9196 2834 9882 2867
rect 8466 2809 8503 2810
rect 8416 2800 8503 2809
rect 8416 2780 8474 2800
rect 8494 2780 8503 2800
rect 8416 2770 8503 2780
rect 8562 2800 8599 2810
rect 8562 2780 8570 2800
rect 8590 2780 8599 2800
rect 8416 2769 8447 2770
rect 8411 2701 8521 2714
rect 8562 2701 8599 2780
rect 8349 2699 8599 2701
rect 8349 2696 8450 2699
rect 8349 2677 8414 2696
rect 7229 2664 7308 2672
rect 7140 2662 7308 2664
rect 6864 2655 7308 2662
rect 8411 2669 8414 2677
rect 8443 2669 8450 2696
rect 8478 2672 8488 2699
rect 8517 2677 8599 2699
rect 8788 2746 8956 2747
rect 9196 2746 9234 2834
rect 9495 2832 9542 2834
rect 9842 2810 9882 2834
rect 8788 2723 9234 2746
rect 9460 2777 9571 2791
rect 9460 2775 9502 2777
rect 9460 2755 9467 2775
rect 9486 2755 9502 2775
rect 9460 2747 9502 2755
rect 9530 2775 9571 2777
rect 9530 2755 9544 2775
rect 9563 2755 9571 2775
rect 9843 2766 9882 2810
rect 9530 2747 9571 2755
rect 9460 2741 9571 2747
rect 8788 2720 9232 2723
rect 8788 2718 8956 2720
rect 8517 2672 8521 2677
rect 8478 2669 8521 2672
rect 8411 2655 8521 2669
rect 6525 2635 6636 2641
rect 6864 2636 7234 2655
rect 7140 2635 7234 2636
rect 6525 2627 6566 2635
rect 6525 2607 6533 2627
rect 6552 2607 6566 2627
rect 6525 2605 6566 2607
rect 6594 2627 6636 2635
rect 6594 2607 6610 2627
rect 6629 2607 6636 2627
rect 7229 2626 7234 2635
rect 7282 2635 7308 2655
rect 7282 2626 7299 2635
rect 7229 2617 7299 2626
rect 6594 2605 6636 2607
rect 5973 2601 6009 2602
rect 5821 2571 5830 2591
rect 5850 2571 5858 2591
rect 5709 2562 5765 2564
rect 5709 2561 5746 2562
rect 5821 2561 5858 2571
rect 5917 2591 6065 2601
rect 6165 2598 6261 2600
rect 5917 2571 5926 2591
rect 5946 2571 6036 2591
rect 6056 2571 6065 2591
rect 5917 2562 6065 2571
rect 6123 2591 6261 2598
rect 6123 2571 6132 2591
rect 6152 2571 6261 2591
rect 6525 2590 6636 2605
rect 6123 2562 6261 2571
rect 5917 2561 5954 2562
rect 5973 2510 6009 2562
rect 6028 2561 6065 2562
rect 6124 2561 6161 2562
rect 5444 2508 5485 2509
rect 5336 2501 5485 2508
rect 4459 2499 4496 2500
rect 4409 2490 4496 2499
rect 4409 2470 4467 2490
rect 4487 2470 4496 2490
rect 4409 2460 4496 2470
rect 4555 2490 4592 2500
rect 4555 2470 4563 2490
rect 4583 2470 4592 2490
rect 5336 2481 5454 2501
rect 5474 2481 5485 2501
rect 5336 2473 5485 2481
rect 5552 2505 5911 2509
rect 5552 2500 5874 2505
rect 5552 2476 5665 2500
rect 5689 2481 5874 2500
rect 5898 2481 5911 2505
rect 5689 2476 5911 2481
rect 5552 2473 5911 2476
rect 5973 2473 6008 2510
rect 6076 2507 6176 2510
rect 6076 2503 6143 2507
rect 6076 2477 6088 2503
rect 6114 2481 6143 2503
rect 6169 2481 6176 2507
rect 6114 2477 6176 2481
rect 6076 2473 6176 2477
rect 4409 2459 4440 2460
rect 4404 2391 4514 2404
rect 4555 2391 4592 2470
rect 4789 2455 4826 2456
rect 4785 2446 4826 2455
rect 5552 2452 5583 2473
rect 5973 2452 6009 2473
rect 5395 2451 5432 2452
rect 5169 2448 5203 2449
rect 4785 2428 4798 2446
rect 4816 2428 4826 2446
rect 4785 2419 4826 2428
rect 5168 2439 5205 2448
rect 5168 2421 5177 2439
rect 5195 2421 5205 2439
rect 4785 2399 4825 2419
rect 5168 2411 5205 2421
rect 5394 2442 5432 2451
rect 5394 2422 5403 2442
rect 5423 2422 5432 2442
rect 5394 2414 5432 2422
rect 5498 2446 5583 2452
rect 5608 2451 5645 2452
rect 5498 2426 5506 2446
rect 5526 2426 5583 2446
rect 5498 2418 5583 2426
rect 5607 2442 5645 2451
rect 5607 2422 5616 2442
rect 5636 2422 5645 2442
rect 5498 2417 5534 2418
rect 5607 2414 5645 2422
rect 5711 2446 5796 2452
rect 5816 2451 5853 2452
rect 5711 2426 5719 2446
rect 5739 2445 5796 2446
rect 5739 2426 5768 2445
rect 5711 2425 5768 2426
rect 5789 2425 5796 2445
rect 5711 2418 5796 2425
rect 5815 2442 5853 2451
rect 5815 2422 5824 2442
rect 5844 2422 5853 2442
rect 5711 2417 5747 2418
rect 5815 2414 5853 2422
rect 5919 2446 6063 2452
rect 5919 2426 5927 2446
rect 5947 2445 6035 2446
rect 5947 2426 5978 2445
rect 5919 2425 5978 2426
rect 6003 2426 6035 2445
rect 6055 2426 6063 2446
rect 6003 2425 6063 2426
rect 5919 2418 6063 2425
rect 5919 2417 5955 2418
rect 6027 2417 6063 2418
rect 6129 2451 6166 2452
rect 6129 2450 6167 2451
rect 6129 2442 6193 2450
rect 6129 2422 6138 2442
rect 6158 2428 6193 2442
rect 6213 2428 6216 2448
rect 6158 2423 6216 2428
rect 6158 2422 6193 2423
rect 4342 2389 4592 2391
rect 4342 2386 4443 2389
rect 2860 2329 2924 2341
rect 3200 2337 3237 2364
rect 3408 2337 3445 2368
rect 3621 2366 3657 2368
rect 4342 2367 4407 2386
rect 3621 2337 3658 2366
rect 4404 2359 4407 2367
rect 4436 2359 4443 2386
rect 4471 2362 4481 2389
rect 4510 2367 4592 2389
rect 4700 2389 4825 2399
rect 4700 2370 4708 2389
rect 4733 2370 4825 2389
rect 4510 2362 4514 2367
rect 4700 2363 4825 2370
rect 4471 2359 4514 2362
rect 4404 2345 4514 2359
rect 2860 2328 2895 2329
rect 2837 2323 2895 2328
rect 2837 2303 2840 2323
rect 2860 2309 2895 2323
rect 2915 2309 2924 2329
rect 2860 2301 2924 2309
rect 2886 2300 2924 2301
rect 2887 2299 2924 2300
rect 2990 2333 3026 2334
rect 3098 2333 3134 2334
rect 2990 2325 3134 2333
rect 2990 2305 2998 2325
rect 3018 2305 3106 2325
rect 3126 2305 3134 2325
rect 2990 2299 3134 2305
rect 3200 2329 3238 2337
rect 3306 2333 3342 2334
rect 3200 2309 3209 2329
rect 3229 2309 3238 2329
rect 3200 2300 3238 2309
rect 3257 2326 3342 2333
rect 3257 2306 3264 2326
rect 3285 2325 3342 2326
rect 3285 2306 3314 2325
rect 3257 2305 3314 2306
rect 3334 2305 3342 2325
rect 3200 2299 3237 2300
rect 3257 2299 3342 2305
rect 3408 2329 3446 2337
rect 3519 2333 3555 2334
rect 3408 2309 3417 2329
rect 3437 2309 3446 2329
rect 3408 2300 3446 2309
rect 3470 2325 3555 2333
rect 3470 2305 3527 2325
rect 3547 2305 3555 2325
rect 3408 2299 3445 2300
rect 3470 2299 3555 2305
rect 3621 2329 3659 2337
rect 3621 2309 3630 2329
rect 3650 2309 3659 2329
rect 3621 2300 3659 2309
rect 4785 2315 4825 2363
rect 5169 2383 5203 2411
rect 5395 2385 5432 2414
rect 5396 2383 5432 2385
rect 5608 2383 5645 2414
rect 5169 2382 5341 2383
rect 5169 2350 5355 2382
rect 5396 2361 5645 2383
rect 5816 2382 5853 2414
rect 6129 2410 6193 2422
rect 6233 2384 6260 2562
rect 8788 2540 8815 2718
rect 8855 2680 8919 2692
rect 9195 2688 9232 2720
rect 9403 2719 9652 2741
rect 9403 2688 9440 2719
rect 9616 2717 9652 2719
rect 9616 2688 9653 2717
rect 8855 2679 8890 2680
rect 8832 2674 8890 2679
rect 8832 2654 8835 2674
rect 8855 2660 8890 2674
rect 8910 2660 8919 2680
rect 8855 2652 8919 2660
rect 8881 2651 8919 2652
rect 8882 2650 8919 2651
rect 8985 2684 9021 2685
rect 9093 2684 9129 2685
rect 8985 2679 9129 2684
rect 8985 2676 9047 2679
rect 8985 2656 8993 2676
rect 9013 2659 9047 2676
rect 9070 2676 9129 2679
rect 9070 2659 9101 2676
rect 9013 2656 9101 2659
rect 9121 2656 9129 2676
rect 8985 2650 9129 2656
rect 9195 2680 9233 2688
rect 9301 2684 9337 2685
rect 9195 2660 9204 2680
rect 9224 2660 9233 2680
rect 9195 2651 9233 2660
rect 9252 2677 9337 2684
rect 9252 2657 9259 2677
rect 9280 2676 9337 2677
rect 9280 2657 9309 2676
rect 9252 2656 9309 2657
rect 9329 2656 9337 2676
rect 9195 2650 9232 2651
rect 9252 2650 9337 2656
rect 9403 2680 9441 2688
rect 9514 2684 9550 2685
rect 9403 2660 9412 2680
rect 9432 2660 9441 2680
rect 9403 2651 9441 2660
rect 9465 2676 9550 2684
rect 9465 2656 9522 2676
rect 9542 2656 9550 2676
rect 9403 2650 9440 2651
rect 9465 2650 9550 2656
rect 9616 2680 9654 2688
rect 9616 2660 9625 2680
rect 9645 2660 9654 2680
rect 9616 2651 9654 2660
rect 9616 2650 9653 2651
rect 9039 2629 9075 2650
rect 9465 2629 9496 2650
rect 8872 2625 8972 2629
rect 8872 2621 8934 2625
rect 8872 2595 8879 2621
rect 8905 2599 8934 2621
rect 8960 2599 8972 2625
rect 8905 2595 8972 2599
rect 8872 2592 8972 2595
rect 9040 2592 9075 2629
rect 9137 2626 9496 2629
rect 9137 2621 9359 2626
rect 9137 2597 9150 2621
rect 9174 2602 9359 2621
rect 9383 2602 9496 2626
rect 9174 2597 9496 2602
rect 9137 2593 9496 2597
rect 9563 2621 9712 2629
rect 9563 2601 9574 2621
rect 9594 2601 9712 2621
rect 9563 2594 9712 2601
rect 9563 2593 9604 2594
rect 8887 2540 8924 2541
rect 8983 2540 9020 2541
rect 9039 2540 9075 2592
rect 9094 2540 9131 2541
rect 8787 2531 8925 2540
rect 8787 2511 8896 2531
rect 8916 2511 8925 2531
rect 8787 2504 8925 2511
rect 8983 2531 9131 2540
rect 8983 2511 8992 2531
rect 9012 2511 9102 2531
rect 9122 2511 9131 2531
rect 8787 2502 8883 2504
rect 8983 2501 9131 2511
rect 9190 2531 9227 2541
rect 9302 2540 9339 2541
rect 9283 2538 9339 2540
rect 9190 2511 9198 2531
rect 9218 2511 9227 2531
rect 9039 2500 9075 2501
rect 6416 2458 6526 2472
rect 6416 2455 6459 2458
rect 6416 2450 6420 2455
rect 6092 2382 6260 2384
rect 5816 2376 6260 2382
rect 5169 2318 5203 2350
rect 3621 2299 3658 2300
rect 3044 2278 3080 2299
rect 3470 2278 3501 2299
rect 4785 2297 4796 2315
rect 4814 2297 4825 2315
rect 4785 2289 4825 2297
rect 5165 2309 5203 2318
rect 5165 2291 5175 2309
rect 5193 2291 5203 2309
rect 4786 2288 4823 2289
rect 5165 2285 5203 2291
rect 5321 2287 5355 2350
rect 5477 2355 5588 2361
rect 5477 2347 5518 2355
rect 5477 2327 5485 2347
rect 5504 2327 5518 2347
rect 5477 2325 5518 2327
rect 5546 2347 5588 2355
rect 5546 2327 5562 2347
rect 5581 2327 5588 2347
rect 5546 2325 5588 2327
rect 5477 2310 5588 2325
rect 5815 2356 6260 2376
rect 5815 2287 5853 2356
rect 6092 2355 6260 2356
rect 6338 2428 6420 2450
rect 6449 2428 6459 2455
rect 6487 2431 6494 2458
rect 6523 2450 6526 2458
rect 8521 2467 8632 2482
rect 8521 2465 8563 2467
rect 6523 2431 6588 2450
rect 6487 2428 6588 2431
rect 6338 2426 6588 2428
rect 6338 2347 6375 2426
rect 6416 2413 6526 2426
rect 6490 2357 6521 2358
rect 6338 2327 6347 2347
rect 6367 2327 6375 2347
rect 6338 2317 6375 2327
rect 6434 2347 6521 2357
rect 6434 2327 6443 2347
rect 6463 2327 6521 2347
rect 6434 2318 6521 2327
rect 6434 2317 6471 2318
rect 5165 2281 5202 2285
rect 2877 2274 2977 2278
rect 2877 2270 2939 2274
rect 2877 2244 2884 2270
rect 2910 2248 2939 2270
rect 2965 2248 2977 2274
rect 2910 2244 2977 2248
rect 2877 2241 2977 2244
rect 3045 2241 3080 2278
rect 3142 2275 3501 2278
rect 3142 2270 3364 2275
rect 3142 2246 3155 2270
rect 3179 2251 3364 2270
rect 3388 2251 3501 2275
rect 3179 2246 3501 2251
rect 3142 2242 3501 2246
rect 3568 2270 3717 2278
rect 5321 2276 5853 2287
rect 3568 2250 3579 2270
rect 3599 2250 3717 2270
rect 5320 2260 5853 2276
rect 6490 2265 6521 2318
rect 6551 2347 6588 2426
rect 6759 2423 7152 2443
rect 7172 2423 7175 2443
rect 8254 2438 8295 2447
rect 6759 2418 7175 2423
rect 7849 2436 8017 2437
rect 8254 2436 8263 2438
rect 6759 2417 7100 2418
rect 6703 2357 6734 2358
rect 6551 2327 6560 2347
rect 6580 2327 6588 2347
rect 6551 2317 6588 2327
rect 6647 2350 6734 2357
rect 6647 2347 6708 2350
rect 6647 2327 6656 2347
rect 6676 2330 6708 2347
rect 6729 2330 6734 2350
rect 6676 2327 6734 2330
rect 6647 2320 6734 2327
rect 6759 2347 6796 2417
rect 7062 2416 7099 2417
rect 7849 2416 8263 2436
rect 8289 2416 8295 2438
rect 8521 2445 8528 2465
rect 8547 2445 8563 2465
rect 8521 2437 8563 2445
rect 8591 2465 8632 2467
rect 8591 2445 8605 2465
rect 8624 2445 8632 2465
rect 8591 2437 8632 2445
rect 8887 2441 8924 2442
rect 9190 2441 9227 2511
rect 9252 2531 9339 2538
rect 9252 2528 9310 2531
rect 9252 2508 9257 2528
rect 9278 2511 9310 2528
rect 9330 2511 9339 2531
rect 9278 2508 9339 2511
rect 9252 2501 9339 2508
rect 9398 2531 9435 2541
rect 9398 2511 9406 2531
rect 9426 2511 9435 2531
rect 9252 2500 9283 2501
rect 8886 2440 9227 2441
rect 8521 2431 8632 2437
rect 8811 2435 9227 2440
rect 7849 2410 8295 2416
rect 7849 2408 8017 2410
rect 6911 2357 6947 2358
rect 6759 2327 6768 2347
rect 6788 2327 6796 2347
rect 6647 2318 6703 2320
rect 6647 2317 6684 2318
rect 6759 2317 6796 2327
rect 6855 2347 7003 2357
rect 7103 2354 7199 2356
rect 6855 2327 6864 2347
rect 6884 2327 6974 2347
rect 6994 2327 7003 2347
rect 6855 2318 7003 2327
rect 7061 2347 7199 2354
rect 7061 2327 7070 2347
rect 7090 2327 7199 2347
rect 7061 2318 7199 2327
rect 6855 2317 6892 2318
rect 6911 2266 6947 2318
rect 6966 2317 7003 2318
rect 7062 2317 7099 2318
rect 6382 2264 6423 2265
rect 5320 2259 5834 2260
rect 3568 2243 3717 2250
rect 6274 2257 6423 2264
rect 4157 2247 4671 2248
rect 3568 2242 3609 2243
rect 3044 2206 3080 2241
rect 2892 2189 2929 2190
rect 2988 2189 3025 2190
rect 3044 2189 3051 2206
rect 2792 2180 2930 2189
rect 2792 2160 2901 2180
rect 2921 2160 2930 2180
rect 2792 2153 2930 2160
rect 2988 2180 3051 2189
rect 2988 2160 2997 2180
rect 3017 2165 3051 2180
rect 3072 2189 3080 2206
rect 3099 2189 3136 2190
rect 3072 2180 3136 2189
rect 3072 2165 3107 2180
rect 3017 2160 3107 2165
rect 3127 2160 3136 2180
rect 2792 2151 2888 2153
rect 2988 2150 3136 2160
rect 3195 2180 3232 2190
rect 3307 2189 3344 2190
rect 3288 2187 3344 2189
rect 3195 2160 3203 2180
rect 3223 2160 3232 2180
rect 3044 2149 3080 2150
rect 1974 2097 2142 2099
rect 1696 2091 2142 2097
rect 764 2067 1180 2072
rect 1359 2070 1470 2076
rect 764 2066 1105 2067
rect 708 2006 739 2007
rect 556 1976 565 1996
rect 585 1976 593 1996
rect 556 1966 593 1976
rect 652 1999 739 2006
rect 652 1996 713 1999
rect 652 1976 661 1996
rect 681 1979 713 1996
rect 734 1979 739 1999
rect 681 1976 739 1979
rect 652 1969 739 1976
rect 764 1996 801 2066
rect 1067 2065 1104 2066
rect 1359 2062 1400 2070
rect 1359 2042 1367 2062
rect 1386 2042 1400 2062
rect 1359 2040 1400 2042
rect 1428 2062 1470 2070
rect 1428 2042 1444 2062
rect 1463 2042 1470 2062
rect 1696 2069 1702 2091
rect 1728 2071 2142 2091
rect 2892 2090 2929 2091
rect 3195 2090 3232 2160
rect 3257 2180 3344 2187
rect 3257 2177 3315 2180
rect 3257 2157 3262 2177
rect 3283 2160 3315 2177
rect 3335 2160 3344 2180
rect 3283 2157 3344 2160
rect 3257 2150 3344 2157
rect 3403 2180 3440 2190
rect 3403 2160 3411 2180
rect 3431 2160 3440 2180
rect 3257 2149 3288 2150
rect 2891 2089 3232 2090
rect 1728 2069 1737 2071
rect 1974 2070 2142 2071
rect 2816 2088 3232 2089
rect 2816 2084 3192 2088
rect 1696 2060 1737 2069
rect 2816 2064 2819 2084
rect 2839 2071 3192 2084
rect 3224 2071 3232 2088
rect 2839 2064 3232 2071
rect 3403 2081 3440 2160
rect 3470 2189 3501 2242
rect 4138 2231 4671 2247
rect 6274 2237 6392 2257
rect 6412 2237 6423 2257
rect 4138 2220 4670 2231
rect 6274 2229 6423 2237
rect 6490 2261 6849 2265
rect 6490 2256 6812 2261
rect 6490 2232 6603 2256
rect 6627 2237 6812 2256
rect 6836 2237 6849 2261
rect 6627 2232 6849 2237
rect 6490 2229 6849 2232
rect 6911 2229 6946 2266
rect 7014 2263 7114 2266
rect 7014 2259 7081 2263
rect 7014 2233 7026 2259
rect 7052 2237 7081 2259
rect 7107 2237 7114 2263
rect 7052 2233 7114 2237
rect 7014 2229 7114 2233
rect 4789 2222 4826 2226
rect 3520 2189 3557 2190
rect 3470 2180 3557 2189
rect 3470 2160 3528 2180
rect 3548 2160 3557 2180
rect 3470 2150 3557 2160
rect 3616 2180 3653 2190
rect 3616 2160 3624 2180
rect 3644 2160 3653 2180
rect 3470 2149 3501 2150
rect 3465 2081 3575 2094
rect 3616 2081 3653 2160
rect 3403 2079 3653 2081
rect 3403 2076 3504 2079
rect 3403 2057 3468 2076
rect 1428 2040 1470 2042
rect 1359 2025 1470 2040
rect 3465 2049 3468 2057
rect 3497 2049 3504 2076
rect 3532 2052 3542 2079
rect 3571 2057 3653 2079
rect 3731 2151 3899 2152
rect 4138 2151 4176 2220
rect 3731 2131 4176 2151
rect 4403 2182 4514 2197
rect 4403 2180 4445 2182
rect 4403 2160 4410 2180
rect 4429 2160 4445 2180
rect 4403 2152 4445 2160
rect 4473 2180 4514 2182
rect 4473 2160 4487 2180
rect 4506 2160 4514 2180
rect 4473 2152 4514 2160
rect 4403 2146 4514 2152
rect 4636 2157 4670 2220
rect 4788 2216 4826 2222
rect 5168 2218 5205 2219
rect 4788 2198 4798 2216
rect 4816 2198 4826 2216
rect 4788 2189 4826 2198
rect 5166 2210 5206 2218
rect 5166 2192 5177 2210
rect 5195 2192 5206 2210
rect 6490 2208 6521 2229
rect 6911 2208 6947 2229
rect 6333 2207 6370 2208
rect 4788 2157 4822 2189
rect 3731 2125 4175 2131
rect 3731 2123 3899 2125
rect 3571 2052 3575 2057
rect 3532 2049 3575 2052
rect 3465 2035 3575 2049
rect 916 2006 952 2007
rect 764 1976 773 1996
rect 793 1976 801 1996
rect 652 1967 708 1969
rect 652 1966 689 1967
rect 764 1966 801 1976
rect 860 1996 1008 2006
rect 1108 2003 1204 2005
rect 860 1976 869 1996
rect 889 1976 979 1996
rect 999 1976 1008 1996
rect 860 1967 1008 1976
rect 1066 1996 1204 2003
rect 1066 1976 1075 1996
rect 1095 1976 1204 1996
rect 1066 1967 1204 1976
rect 860 1966 897 1967
rect 916 1915 952 1967
rect 971 1966 1008 1967
rect 1067 1966 1104 1967
rect 387 1913 428 1914
rect 279 1906 428 1913
rect 279 1886 397 1906
rect 417 1886 428 1906
rect 279 1878 428 1886
rect 495 1910 854 1914
rect 495 1905 817 1910
rect 495 1881 608 1905
rect 632 1886 817 1905
rect 841 1886 854 1910
rect 632 1881 854 1886
rect 495 1878 854 1881
rect 916 1878 951 1915
rect 1019 1912 1119 1915
rect 1019 1908 1086 1912
rect 1019 1882 1031 1908
rect 1057 1886 1086 1908
rect 1112 1886 1119 1912
rect 1057 1882 1119 1886
rect 1019 1878 1119 1882
rect 495 1857 526 1878
rect 916 1857 952 1878
rect 338 1856 375 1857
rect 337 1847 375 1856
rect 337 1827 346 1847
rect 366 1827 375 1847
rect 337 1819 375 1827
rect 441 1851 526 1857
rect 551 1856 588 1857
rect 441 1831 449 1851
rect 469 1831 526 1851
rect 441 1823 526 1831
rect 550 1847 588 1856
rect 550 1827 559 1847
rect 579 1827 588 1847
rect 441 1822 477 1823
rect 550 1819 588 1827
rect 654 1851 739 1857
rect 759 1856 796 1857
rect 654 1831 662 1851
rect 682 1850 739 1851
rect 682 1831 711 1850
rect 654 1830 711 1831
rect 732 1830 739 1850
rect 654 1823 739 1830
rect 758 1847 796 1856
rect 758 1827 767 1847
rect 787 1827 796 1847
rect 654 1822 690 1823
rect 758 1819 796 1827
rect 862 1851 1006 1857
rect 862 1831 870 1851
rect 890 1848 978 1851
rect 890 1831 921 1848
rect 862 1828 921 1831
rect 944 1831 978 1848
rect 998 1831 1006 1851
rect 944 1828 1006 1831
rect 862 1823 1006 1828
rect 862 1822 898 1823
rect 970 1822 1006 1823
rect 1072 1856 1109 1857
rect 1072 1855 1110 1856
rect 1072 1847 1136 1855
rect 1072 1827 1081 1847
rect 1101 1833 1136 1847
rect 1156 1833 1159 1853
rect 1101 1828 1159 1833
rect 1101 1827 1136 1828
rect 338 1790 375 1819
rect 339 1788 375 1790
rect 551 1788 588 1819
rect 339 1766 588 1788
rect 759 1787 796 1819
rect 1072 1815 1136 1827
rect 1176 1789 1203 1967
rect 3731 1945 3758 2123
rect 3798 2085 3862 2097
rect 4138 2093 4175 2125
rect 4346 2124 4595 2146
rect 4636 2125 4822 2157
rect 4650 2124 4822 2125
rect 4346 2093 4383 2124
rect 4559 2122 4595 2124
rect 4559 2093 4596 2122
rect 4788 2096 4822 2124
rect 5166 2144 5206 2192
rect 6332 2198 6370 2207
rect 6332 2178 6341 2198
rect 6361 2178 6370 2198
rect 6332 2170 6370 2178
rect 6436 2202 6521 2208
rect 6546 2207 6583 2208
rect 6436 2182 6444 2202
rect 6464 2182 6521 2202
rect 6436 2174 6521 2182
rect 6545 2198 6583 2207
rect 6545 2178 6554 2198
rect 6574 2178 6583 2198
rect 6436 2173 6472 2174
rect 6545 2170 6583 2178
rect 6649 2202 6734 2208
rect 6754 2207 6791 2208
rect 6649 2182 6657 2202
rect 6677 2201 6734 2202
rect 6677 2182 6706 2201
rect 6649 2181 6706 2182
rect 6727 2181 6734 2201
rect 6649 2174 6734 2181
rect 6753 2198 6791 2207
rect 6753 2178 6762 2198
rect 6782 2178 6791 2198
rect 6649 2173 6685 2174
rect 6753 2170 6791 2178
rect 6857 2202 7001 2208
rect 6857 2182 6865 2202
rect 6885 2185 6921 2202
rect 6941 2185 6973 2202
rect 6885 2182 6973 2185
rect 6993 2182 7001 2202
rect 6857 2174 7001 2182
rect 6857 2173 6893 2174
rect 6965 2173 7001 2174
rect 7067 2207 7104 2208
rect 7067 2206 7105 2207
rect 7067 2198 7131 2206
rect 7067 2178 7076 2198
rect 7096 2184 7131 2198
rect 7151 2184 7154 2204
rect 7096 2179 7154 2184
rect 7096 2178 7131 2179
rect 5477 2148 5587 2162
rect 5477 2145 5520 2148
rect 5166 2137 5291 2144
rect 5477 2140 5481 2145
rect 5166 2118 5258 2137
rect 5283 2118 5291 2137
rect 5166 2108 5291 2118
rect 5399 2118 5481 2140
rect 5510 2118 5520 2145
rect 5548 2121 5555 2148
rect 5584 2140 5587 2148
rect 6333 2141 6370 2170
rect 5584 2121 5649 2140
rect 6334 2139 6370 2141
rect 6546 2139 6583 2170
rect 6754 2143 6791 2170
rect 7067 2166 7131 2178
rect 5548 2118 5649 2121
rect 5399 2116 5649 2118
rect 3798 2084 3833 2085
rect 3775 2079 3833 2084
rect 3775 2059 3778 2079
rect 3798 2065 3833 2079
rect 3853 2065 3862 2085
rect 3798 2057 3862 2065
rect 3824 2056 3862 2057
rect 3825 2055 3862 2056
rect 3928 2089 3964 2090
rect 4036 2089 4072 2090
rect 3928 2082 4072 2089
rect 3928 2081 3988 2082
rect 3928 2061 3936 2081
rect 3956 2062 3988 2081
rect 4013 2081 4072 2082
rect 4013 2062 4044 2081
rect 3956 2061 4044 2062
rect 4064 2061 4072 2081
rect 3928 2055 4072 2061
rect 4138 2085 4176 2093
rect 4244 2089 4280 2090
rect 4138 2065 4147 2085
rect 4167 2065 4176 2085
rect 4138 2056 4176 2065
rect 4195 2082 4280 2089
rect 4195 2062 4202 2082
rect 4223 2081 4280 2082
rect 4223 2062 4252 2081
rect 4195 2061 4252 2062
rect 4272 2061 4280 2081
rect 4138 2055 4175 2056
rect 4195 2055 4280 2061
rect 4346 2085 4384 2093
rect 4457 2089 4493 2090
rect 4346 2065 4355 2085
rect 4375 2065 4384 2085
rect 4346 2056 4384 2065
rect 4408 2081 4493 2089
rect 4408 2061 4465 2081
rect 4485 2061 4493 2081
rect 4346 2055 4383 2056
rect 4408 2055 4493 2061
rect 4559 2085 4597 2093
rect 4559 2065 4568 2085
rect 4588 2065 4597 2085
rect 4559 2056 4597 2065
rect 4786 2086 4823 2096
rect 5166 2088 5206 2108
rect 4786 2068 4796 2086
rect 4814 2068 4823 2086
rect 4786 2059 4823 2068
rect 5165 2079 5206 2088
rect 5165 2061 5175 2079
rect 5193 2061 5206 2079
rect 4788 2058 4822 2059
rect 4559 2055 4596 2056
rect 3982 2034 4018 2055
rect 4408 2034 4439 2055
rect 5165 2052 5206 2061
rect 5165 2051 5202 2052
rect 5399 2037 5436 2116
rect 5477 2103 5587 2116
rect 5551 2047 5582 2048
rect 3815 2030 3915 2034
rect 3815 2026 3877 2030
rect 3815 2000 3822 2026
rect 3848 2004 3877 2026
rect 3903 2004 3915 2030
rect 3848 2000 3915 2004
rect 3815 1997 3915 2000
rect 3983 1997 4018 2034
rect 4080 2031 4439 2034
rect 4080 2026 4302 2031
rect 4080 2002 4093 2026
rect 4117 2007 4302 2026
rect 4326 2007 4439 2031
rect 4117 2002 4439 2007
rect 4080 1998 4439 2002
rect 4506 2026 4655 2034
rect 4506 2006 4517 2026
rect 4537 2006 4655 2026
rect 5399 2017 5408 2037
rect 5428 2017 5436 2037
rect 5399 2007 5436 2017
rect 5495 2037 5582 2047
rect 5495 2017 5504 2037
rect 5524 2017 5582 2037
rect 5495 2008 5582 2017
rect 5495 2007 5532 2008
rect 4506 1999 4655 2006
rect 4506 1998 4547 1999
rect 3830 1945 3867 1946
rect 3926 1945 3963 1946
rect 3982 1945 4018 1997
rect 4037 1945 4074 1946
rect 3730 1936 3868 1945
rect 3325 1915 3436 1930
rect 3325 1913 3367 1915
rect 2995 1892 3100 1894
rect 2653 1884 2821 1885
rect 2995 1884 3044 1892
rect 2653 1865 3044 1884
rect 3075 1865 3100 1892
rect 3325 1893 3332 1913
rect 3351 1893 3367 1913
rect 3325 1885 3367 1893
rect 3395 1913 3436 1915
rect 3395 1893 3409 1913
rect 3428 1893 3436 1913
rect 3730 1916 3839 1936
rect 3859 1916 3868 1936
rect 3730 1909 3868 1916
rect 3926 1936 4074 1945
rect 3926 1916 3935 1936
rect 3955 1916 4045 1936
rect 4065 1916 4074 1936
rect 3730 1907 3826 1909
rect 3926 1906 4074 1916
rect 4133 1936 4170 1946
rect 4245 1945 4282 1946
rect 4226 1943 4282 1945
rect 4133 1916 4141 1936
rect 4161 1916 4170 1936
rect 3982 1905 4018 1906
rect 3395 1885 3436 1893
rect 3325 1879 3436 1885
rect 2653 1858 3100 1865
rect 2653 1856 2821 1858
rect 1501 1825 1611 1839
rect 1501 1822 1544 1825
rect 1501 1817 1505 1822
rect 1035 1787 1203 1789
rect 759 1784 1203 1787
rect 420 1760 531 1766
rect 420 1752 461 1760
rect 109 1697 148 1741
rect 420 1732 428 1752
rect 447 1732 461 1752
rect 420 1730 461 1732
rect 489 1752 531 1760
rect 489 1732 505 1752
rect 524 1732 531 1752
rect 489 1730 531 1732
rect 420 1715 531 1730
rect 757 1761 1203 1784
rect 109 1673 149 1697
rect 449 1673 496 1675
rect 757 1673 795 1761
rect 1035 1760 1203 1761
rect 1423 1795 1505 1817
rect 1534 1795 1544 1822
rect 1572 1798 1579 1825
rect 1608 1817 1611 1825
rect 1608 1798 1673 1817
rect 1572 1795 1673 1798
rect 1423 1793 1673 1795
rect 1423 1714 1460 1793
rect 1501 1780 1611 1793
rect 1575 1724 1606 1725
rect 1423 1694 1432 1714
rect 1452 1694 1460 1714
rect 1423 1684 1460 1694
rect 1519 1714 1606 1724
rect 1519 1694 1528 1714
rect 1548 1694 1606 1714
rect 1519 1685 1606 1694
rect 1519 1684 1556 1685
rect 109 1640 795 1673
rect 109 1583 148 1640
rect 757 1638 795 1640
rect 1575 1632 1606 1685
rect 1636 1714 1673 1793
rect 1844 1806 2237 1810
rect 1844 1789 1863 1806
rect 1883 1790 2237 1806
rect 2257 1790 2260 1810
rect 1883 1789 2260 1790
rect 1844 1785 2260 1789
rect 1844 1784 2185 1785
rect 1788 1724 1819 1725
rect 1636 1694 1645 1714
rect 1665 1694 1673 1714
rect 1636 1684 1673 1694
rect 1732 1717 1819 1724
rect 1732 1714 1793 1717
rect 1732 1694 1741 1714
rect 1761 1697 1793 1714
rect 1814 1697 1819 1717
rect 1761 1694 1819 1697
rect 1732 1687 1819 1694
rect 1844 1714 1881 1784
rect 2147 1783 2184 1784
rect 1996 1724 2032 1725
rect 1844 1694 1853 1714
rect 1873 1694 1881 1714
rect 1732 1685 1788 1687
rect 1732 1684 1769 1685
rect 1844 1684 1881 1694
rect 1940 1714 2088 1724
rect 2256 1723 2285 1724
rect 2188 1721 2285 1723
rect 1940 1694 1949 1714
rect 1969 1710 2059 1714
rect 1969 1694 2002 1710
rect 1940 1685 2002 1694
rect 1940 1684 1977 1685
rect 1996 1672 2002 1685
rect 2025 1694 2059 1710
rect 2079 1694 2088 1714
rect 2025 1685 2088 1694
rect 2146 1714 2285 1721
rect 2146 1694 2155 1714
rect 2175 1694 2285 1714
rect 2146 1685 2285 1694
rect 2025 1672 2032 1685
rect 2051 1684 2088 1685
rect 2147 1684 2184 1685
rect 1996 1633 2032 1672
rect 1467 1631 1508 1632
rect 1359 1624 1508 1631
rect 1359 1604 1477 1624
rect 1497 1604 1508 1624
rect 1359 1596 1508 1604
rect 1575 1628 1934 1632
rect 1575 1623 1897 1628
rect 1575 1599 1688 1623
rect 1712 1604 1897 1623
rect 1921 1604 1934 1628
rect 1712 1599 1934 1604
rect 1575 1596 1934 1599
rect 1996 1596 2031 1633
rect 2099 1630 2199 1633
rect 2099 1626 2166 1630
rect 2099 1600 2111 1626
rect 2137 1604 2166 1626
rect 2192 1604 2199 1630
rect 2137 1600 2199 1604
rect 2099 1596 2199 1600
rect 109 1581 157 1583
rect 109 1563 120 1581
rect 138 1563 157 1581
rect 1575 1575 1606 1596
rect 1996 1575 2032 1596
rect 1418 1574 1455 1575
rect 109 1554 157 1563
rect 110 1553 157 1554
rect 423 1558 533 1572
rect 423 1555 466 1558
rect 423 1550 427 1555
rect 345 1528 427 1550
rect 456 1528 466 1555
rect 494 1531 501 1558
rect 530 1550 533 1558
rect 1417 1565 1455 1574
rect 530 1531 595 1550
rect 1417 1545 1426 1565
rect 1446 1545 1455 1565
rect 494 1528 595 1531
rect 345 1526 595 1528
rect 113 1490 150 1491
rect 109 1487 150 1490
rect 109 1482 151 1487
rect 109 1464 122 1482
rect 140 1464 151 1482
rect 109 1450 151 1464
rect 189 1450 236 1454
rect 109 1444 236 1450
rect 109 1415 197 1444
rect 226 1415 236 1444
rect 345 1447 382 1526
rect 423 1513 533 1526
rect 497 1457 528 1458
rect 345 1427 354 1447
rect 374 1427 382 1447
rect 345 1417 382 1427
rect 441 1447 528 1457
rect 441 1427 450 1447
rect 470 1427 528 1447
rect 441 1418 528 1427
rect 441 1417 478 1418
rect 109 1411 236 1415
rect 109 1394 148 1411
rect 189 1410 236 1411
rect 109 1376 120 1394
rect 138 1376 148 1394
rect 109 1367 148 1376
rect 110 1366 147 1367
rect 497 1365 528 1418
rect 558 1447 595 1526
rect 766 1523 1159 1543
rect 1179 1523 1182 1543
rect 1417 1537 1455 1545
rect 1521 1569 1606 1575
rect 1631 1574 1668 1575
rect 1521 1549 1529 1569
rect 1549 1549 1606 1569
rect 1521 1541 1606 1549
rect 1630 1565 1668 1574
rect 1630 1545 1639 1565
rect 1659 1545 1668 1565
rect 1521 1540 1557 1541
rect 1630 1537 1668 1545
rect 1734 1569 1819 1575
rect 1839 1574 1876 1575
rect 1734 1549 1742 1569
rect 1762 1568 1819 1569
rect 1762 1549 1791 1568
rect 1734 1548 1791 1549
rect 1812 1548 1819 1568
rect 1734 1541 1819 1548
rect 1838 1565 1876 1574
rect 1838 1545 1847 1565
rect 1867 1545 1876 1565
rect 1734 1540 1770 1541
rect 1838 1537 1876 1545
rect 1942 1569 2086 1575
rect 1942 1549 1950 1569
rect 1970 1549 2058 1569
rect 2078 1549 2086 1569
rect 1942 1541 2086 1549
rect 1942 1540 1978 1541
rect 2050 1540 2086 1541
rect 2152 1574 2189 1575
rect 2152 1573 2190 1574
rect 2152 1565 2216 1573
rect 2152 1545 2161 1565
rect 2181 1551 2216 1565
rect 2236 1551 2239 1571
rect 2181 1546 2239 1551
rect 2181 1545 2216 1546
rect 766 1518 1182 1523
rect 766 1517 1107 1518
rect 710 1457 741 1458
rect 558 1427 567 1447
rect 587 1427 595 1447
rect 558 1417 595 1427
rect 654 1450 741 1457
rect 654 1447 715 1450
rect 654 1427 663 1447
rect 683 1430 715 1447
rect 736 1430 741 1450
rect 683 1427 741 1430
rect 654 1420 741 1427
rect 766 1447 803 1517
rect 1069 1516 1106 1517
rect 1418 1508 1455 1537
rect 1419 1506 1455 1508
rect 1631 1506 1668 1537
rect 1419 1484 1668 1506
rect 1839 1505 1876 1537
rect 2152 1533 2216 1545
rect 2256 1507 2285 1685
rect 2653 1678 2680 1856
rect 2720 1818 2784 1830
rect 3060 1826 3097 1858
rect 3268 1857 3517 1879
rect 3268 1826 3305 1857
rect 3481 1855 3517 1857
rect 3481 1826 3518 1855
rect 3830 1846 3867 1847
rect 4133 1846 4170 1916
rect 4195 1936 4282 1943
rect 4195 1933 4253 1936
rect 4195 1913 4200 1933
rect 4221 1916 4253 1933
rect 4273 1916 4282 1936
rect 4221 1913 4282 1916
rect 4195 1906 4282 1913
rect 4341 1936 4378 1946
rect 4341 1916 4349 1936
rect 4369 1916 4378 1936
rect 4195 1905 4226 1906
rect 3829 1845 4170 1846
rect 3754 1840 4170 1845
rect 2720 1817 2755 1818
rect 2697 1812 2755 1817
rect 2697 1792 2700 1812
rect 2720 1798 2755 1812
rect 2775 1798 2784 1818
rect 2720 1790 2784 1798
rect 2746 1789 2784 1790
rect 2747 1788 2784 1789
rect 2850 1822 2886 1823
rect 2958 1822 2994 1823
rect 2850 1817 2994 1822
rect 2850 1814 2910 1817
rect 2850 1794 2858 1814
rect 2878 1796 2910 1814
rect 2937 1814 2994 1817
rect 2937 1796 2966 1814
rect 2878 1794 2966 1796
rect 2986 1794 2994 1814
rect 2850 1788 2994 1794
rect 3060 1818 3098 1826
rect 3166 1822 3202 1823
rect 3060 1798 3069 1818
rect 3089 1798 3098 1818
rect 3060 1789 3098 1798
rect 3117 1815 3202 1822
rect 3117 1795 3124 1815
rect 3145 1814 3202 1815
rect 3145 1795 3174 1814
rect 3117 1794 3174 1795
rect 3194 1794 3202 1814
rect 3060 1788 3097 1789
rect 3117 1788 3202 1794
rect 3268 1818 3306 1826
rect 3379 1822 3415 1823
rect 3268 1798 3277 1818
rect 3297 1798 3306 1818
rect 3268 1789 3306 1798
rect 3330 1814 3415 1822
rect 3330 1794 3387 1814
rect 3407 1794 3415 1814
rect 3268 1788 3305 1789
rect 3330 1788 3415 1794
rect 3481 1818 3519 1826
rect 3754 1820 3757 1840
rect 3777 1820 4170 1840
rect 4341 1837 4378 1916
rect 4408 1945 4439 1998
rect 4789 1996 4826 1997
rect 4788 1987 4827 1996
rect 4788 1969 4798 1987
rect 4816 1969 4827 1987
rect 5168 1985 5205 1989
rect 4700 1952 4747 1953
rect 4788 1952 4827 1969
rect 4700 1948 4827 1952
rect 4458 1945 4495 1946
rect 4408 1936 4495 1945
rect 4408 1916 4466 1936
rect 4486 1916 4495 1936
rect 4408 1906 4495 1916
rect 4554 1936 4591 1946
rect 4554 1916 4562 1936
rect 4582 1916 4591 1936
rect 4408 1905 4439 1906
rect 4403 1837 4513 1850
rect 4554 1837 4591 1916
rect 4700 1919 4710 1948
rect 4739 1919 4827 1948
rect 4700 1913 4827 1919
rect 4700 1909 4747 1913
rect 4785 1899 4827 1913
rect 4785 1881 4796 1899
rect 4814 1881 4827 1899
rect 4785 1876 4827 1881
rect 4786 1873 4827 1876
rect 5165 1980 5205 1985
rect 5165 1962 5177 1980
rect 5195 1962 5205 1980
rect 4786 1872 4823 1873
rect 4341 1835 4591 1837
rect 4341 1832 4442 1835
rect 3481 1798 3490 1818
rect 3510 1798 3519 1818
rect 4341 1813 4406 1832
rect 3481 1789 3519 1798
rect 4403 1805 4406 1813
rect 4435 1805 4442 1832
rect 4470 1808 4480 1835
rect 4509 1813 4591 1835
rect 4509 1808 4513 1813
rect 4470 1805 4513 1808
rect 4403 1791 4513 1805
rect 4779 1809 4826 1810
rect 4779 1800 4827 1809
rect 3481 1788 3518 1789
rect 2904 1767 2940 1788
rect 3330 1767 3361 1788
rect 4779 1782 4798 1800
rect 4816 1782 4827 1800
rect 4779 1780 4827 1782
rect 2737 1763 2837 1767
rect 2737 1759 2799 1763
rect 2737 1733 2744 1759
rect 2770 1737 2799 1759
rect 2825 1737 2837 1763
rect 2770 1733 2837 1737
rect 2737 1730 2837 1733
rect 2905 1730 2940 1767
rect 3002 1764 3361 1767
rect 3002 1759 3224 1764
rect 3002 1735 3015 1759
rect 3039 1740 3224 1759
rect 3248 1740 3361 1764
rect 3039 1735 3361 1740
rect 3002 1731 3361 1735
rect 3428 1759 3577 1767
rect 3428 1739 3439 1759
rect 3459 1739 3577 1759
rect 3428 1732 3577 1739
rect 3428 1731 3469 1732
rect 2752 1678 2789 1679
rect 2848 1678 2885 1679
rect 2904 1678 2940 1730
rect 2959 1678 2996 1679
rect 2652 1669 2790 1678
rect 2652 1649 2761 1669
rect 2781 1649 2790 1669
rect 2652 1642 2790 1649
rect 2848 1669 2996 1678
rect 2848 1649 2857 1669
rect 2877 1649 2967 1669
rect 2987 1649 2996 1669
rect 2652 1640 2748 1642
rect 2848 1639 2996 1649
rect 3055 1669 3092 1679
rect 3167 1678 3204 1679
rect 3148 1676 3204 1678
rect 3055 1649 3063 1669
rect 3083 1649 3092 1669
rect 2904 1638 2940 1639
rect 2752 1579 2789 1580
rect 3055 1579 3092 1649
rect 3117 1669 3204 1676
rect 3117 1666 3175 1669
rect 3117 1646 3122 1666
rect 3143 1649 3175 1666
rect 3195 1649 3204 1669
rect 3143 1646 3204 1649
rect 3117 1639 3204 1646
rect 3263 1669 3300 1679
rect 3263 1649 3271 1669
rect 3291 1649 3300 1669
rect 3117 1638 3148 1639
rect 2751 1578 3092 1579
rect 2676 1574 3092 1578
rect 2676 1573 3053 1574
rect 2676 1553 2679 1573
rect 2699 1557 3053 1573
rect 3073 1557 3092 1574
rect 2699 1553 3092 1557
rect 3263 1570 3300 1649
rect 3330 1678 3361 1731
rect 4141 1723 4179 1725
rect 4788 1723 4827 1780
rect 4141 1690 4827 1723
rect 3380 1678 3417 1679
rect 3330 1669 3417 1678
rect 3330 1649 3388 1669
rect 3408 1649 3417 1669
rect 3330 1639 3417 1649
rect 3476 1669 3513 1679
rect 3476 1649 3484 1669
rect 3504 1649 3513 1669
rect 3330 1638 3361 1639
rect 3325 1570 3435 1583
rect 3476 1570 3513 1649
rect 3263 1568 3513 1570
rect 3263 1565 3364 1568
rect 3263 1546 3328 1565
rect 3325 1538 3328 1546
rect 3357 1538 3364 1565
rect 3392 1541 3402 1568
rect 3431 1546 3513 1568
rect 3733 1602 3901 1603
rect 4141 1602 4179 1690
rect 4440 1688 4487 1690
rect 4787 1666 4827 1690
rect 3733 1579 4179 1602
rect 4405 1633 4516 1648
rect 4405 1631 4447 1633
rect 4405 1611 4412 1631
rect 4431 1611 4447 1631
rect 4405 1603 4447 1611
rect 4475 1631 4516 1633
rect 4475 1611 4489 1631
rect 4508 1611 4516 1631
rect 4788 1622 4827 1666
rect 4475 1603 4516 1611
rect 4405 1597 4516 1603
rect 3733 1576 4177 1579
rect 3733 1574 3901 1576
rect 3431 1541 3435 1546
rect 3392 1538 3435 1541
rect 3325 1524 3435 1538
rect 2115 1505 2285 1507
rect 1836 1498 2285 1505
rect 1500 1478 1611 1484
rect 1500 1470 1541 1478
rect 918 1457 954 1458
rect 766 1427 775 1447
rect 795 1427 803 1447
rect 654 1418 710 1420
rect 654 1417 691 1418
rect 766 1417 803 1427
rect 862 1447 1010 1457
rect 1110 1454 1206 1456
rect 862 1427 871 1447
rect 891 1427 981 1447
rect 1001 1427 1010 1447
rect 862 1418 1010 1427
rect 1068 1447 1206 1454
rect 1068 1427 1077 1447
rect 1097 1427 1206 1447
rect 1500 1450 1508 1470
rect 1527 1450 1541 1470
rect 1500 1448 1541 1450
rect 1569 1470 1611 1478
rect 1569 1450 1585 1470
rect 1604 1450 1611 1470
rect 1836 1471 1861 1498
rect 1892 1479 2285 1498
rect 1892 1471 1941 1479
rect 2115 1478 2285 1479
rect 1836 1469 1941 1471
rect 1569 1448 1611 1450
rect 1500 1433 1611 1448
rect 1068 1418 1206 1427
rect 862 1417 899 1418
rect 918 1366 954 1418
rect 973 1417 1010 1418
rect 1069 1417 1106 1418
rect 389 1364 430 1365
rect 281 1357 430 1364
rect 281 1337 399 1357
rect 419 1337 430 1357
rect 281 1329 430 1337
rect 497 1361 856 1365
rect 497 1356 819 1361
rect 497 1332 610 1356
rect 634 1337 819 1356
rect 843 1337 856 1361
rect 634 1332 856 1337
rect 497 1329 856 1332
rect 918 1329 953 1366
rect 1021 1363 1121 1366
rect 1021 1359 1088 1363
rect 1021 1333 1033 1359
rect 1059 1337 1088 1359
rect 1114 1337 1121 1363
rect 1059 1333 1121 1337
rect 1021 1329 1121 1333
rect 497 1308 528 1329
rect 918 1308 954 1329
rect 340 1307 377 1308
rect 114 1304 148 1305
rect 113 1295 150 1304
rect 113 1277 122 1295
rect 140 1277 150 1295
rect 113 1267 150 1277
rect 339 1298 377 1307
rect 339 1278 348 1298
rect 368 1278 377 1298
rect 339 1270 377 1278
rect 443 1302 528 1308
rect 553 1307 590 1308
rect 443 1282 451 1302
rect 471 1282 528 1302
rect 443 1274 528 1282
rect 552 1298 590 1307
rect 552 1278 561 1298
rect 581 1278 590 1298
rect 443 1273 479 1274
rect 552 1270 590 1278
rect 656 1302 741 1308
rect 761 1307 798 1308
rect 656 1282 664 1302
rect 684 1301 741 1302
rect 684 1282 713 1301
rect 656 1281 713 1282
rect 734 1281 741 1301
rect 656 1274 741 1281
rect 760 1298 798 1307
rect 760 1278 769 1298
rect 789 1278 798 1298
rect 656 1273 692 1274
rect 760 1270 798 1278
rect 864 1302 1008 1308
rect 864 1282 872 1302
rect 892 1301 980 1302
rect 892 1282 923 1301
rect 864 1281 923 1282
rect 948 1282 980 1301
rect 1000 1282 1008 1302
rect 948 1281 1008 1282
rect 864 1274 1008 1281
rect 864 1273 900 1274
rect 972 1273 1008 1274
rect 1074 1307 1111 1308
rect 1074 1306 1112 1307
rect 1074 1298 1138 1306
rect 1074 1278 1083 1298
rect 1103 1284 1138 1298
rect 1158 1284 1161 1304
rect 1103 1279 1161 1284
rect 1103 1278 1138 1279
rect 114 1239 148 1267
rect 340 1241 377 1270
rect 341 1239 377 1241
rect 553 1239 590 1270
rect 114 1238 286 1239
rect 114 1206 300 1238
rect 341 1217 590 1239
rect 761 1238 798 1270
rect 1074 1266 1138 1278
rect 1178 1240 1205 1418
rect 3733 1396 3760 1574
rect 3800 1536 3864 1548
rect 4140 1544 4177 1576
rect 4348 1575 4597 1597
rect 4348 1544 4385 1575
rect 4561 1573 4597 1575
rect 4561 1544 4598 1573
rect 3800 1535 3835 1536
rect 3777 1530 3835 1535
rect 3777 1510 3780 1530
rect 3800 1516 3835 1530
rect 3855 1516 3864 1536
rect 3800 1508 3864 1516
rect 3826 1507 3864 1508
rect 3827 1506 3864 1507
rect 3930 1540 3966 1541
rect 4038 1540 4074 1541
rect 3930 1535 4074 1540
rect 3930 1532 3992 1535
rect 3930 1512 3938 1532
rect 3958 1515 3992 1532
rect 4015 1532 4074 1535
rect 4015 1515 4046 1532
rect 3958 1512 4046 1515
rect 4066 1512 4074 1532
rect 3930 1506 4074 1512
rect 4140 1536 4178 1544
rect 4246 1540 4282 1541
rect 4140 1516 4149 1536
rect 4169 1516 4178 1536
rect 4140 1507 4178 1516
rect 4197 1533 4282 1540
rect 4197 1513 4204 1533
rect 4225 1532 4282 1533
rect 4225 1513 4254 1532
rect 4197 1512 4254 1513
rect 4274 1512 4282 1532
rect 4140 1506 4177 1507
rect 4197 1506 4282 1512
rect 4348 1536 4386 1544
rect 4459 1540 4495 1541
rect 4348 1516 4357 1536
rect 4377 1516 4386 1536
rect 4348 1507 4386 1516
rect 4410 1532 4495 1540
rect 4410 1512 4467 1532
rect 4487 1512 4495 1532
rect 4348 1506 4385 1507
rect 4410 1506 4495 1512
rect 4561 1536 4599 1544
rect 4561 1516 4570 1536
rect 4590 1516 4599 1536
rect 4561 1507 4599 1516
rect 4561 1506 4598 1507
rect 3984 1485 4020 1506
rect 4410 1485 4441 1506
rect 3817 1481 3917 1485
rect 3817 1477 3879 1481
rect 3817 1451 3824 1477
rect 3850 1455 3879 1477
rect 3905 1455 3917 1481
rect 3850 1451 3917 1455
rect 3817 1448 3917 1451
rect 3985 1448 4020 1485
rect 4082 1482 4441 1485
rect 4082 1477 4304 1482
rect 4082 1453 4095 1477
rect 4119 1458 4304 1477
rect 4328 1458 4441 1482
rect 4119 1453 4441 1458
rect 4082 1449 4441 1453
rect 4508 1477 4657 1485
rect 4508 1457 4519 1477
rect 4539 1457 4657 1477
rect 4508 1450 4657 1457
rect 4508 1449 4549 1450
rect 3832 1396 3869 1397
rect 3928 1396 3965 1397
rect 3984 1396 4020 1448
rect 4039 1396 4076 1397
rect 3732 1387 3870 1396
rect 3732 1367 3841 1387
rect 3861 1367 3870 1387
rect 3732 1360 3870 1367
rect 3928 1387 4076 1396
rect 3928 1367 3937 1387
rect 3957 1367 4047 1387
rect 4067 1367 4076 1387
rect 3732 1358 3828 1360
rect 3928 1357 4076 1367
rect 4135 1387 4172 1397
rect 4247 1396 4284 1397
rect 4228 1394 4284 1396
rect 4135 1367 4143 1387
rect 4163 1367 4172 1387
rect 3984 1356 4020 1357
rect 1361 1314 1471 1328
rect 1361 1311 1404 1314
rect 1361 1306 1365 1311
rect 1037 1238 1205 1240
rect 761 1232 1205 1238
rect 114 1174 148 1206
rect 110 1165 148 1174
rect 110 1147 120 1165
rect 138 1147 148 1165
rect 110 1141 148 1147
rect 266 1143 300 1206
rect 422 1211 533 1217
rect 422 1203 463 1211
rect 422 1183 430 1203
rect 449 1183 463 1203
rect 422 1181 463 1183
rect 491 1203 533 1211
rect 491 1183 507 1203
rect 526 1183 533 1203
rect 491 1181 533 1183
rect 422 1166 533 1181
rect 760 1212 1205 1232
rect 760 1143 798 1212
rect 1037 1211 1205 1212
rect 1283 1284 1365 1306
rect 1394 1284 1404 1311
rect 1432 1287 1439 1314
rect 1468 1306 1471 1314
rect 3466 1323 3577 1338
rect 3466 1321 3508 1323
rect 1468 1287 1533 1306
rect 1432 1284 1533 1287
rect 1283 1282 1533 1284
rect 1283 1203 1320 1282
rect 1361 1269 1471 1282
rect 1435 1213 1466 1214
rect 1283 1183 1292 1203
rect 1312 1183 1320 1203
rect 1283 1173 1320 1183
rect 1379 1203 1466 1213
rect 1379 1183 1388 1203
rect 1408 1183 1466 1203
rect 1379 1174 1466 1183
rect 1379 1173 1416 1174
rect 110 1137 147 1141
rect 266 1132 798 1143
rect 265 1116 798 1132
rect 1435 1121 1466 1174
rect 1496 1203 1533 1282
rect 1704 1292 2097 1299
rect 1704 1275 1712 1292
rect 1744 1279 2097 1292
rect 2117 1279 2120 1299
rect 3199 1294 3240 1303
rect 1744 1275 2120 1279
rect 1704 1274 2120 1275
rect 2794 1292 2962 1293
rect 3199 1292 3208 1294
rect 1704 1273 2045 1274
rect 1648 1213 1679 1214
rect 1496 1183 1505 1203
rect 1525 1183 1533 1203
rect 1496 1173 1533 1183
rect 1592 1206 1679 1213
rect 1592 1203 1653 1206
rect 1592 1183 1601 1203
rect 1621 1186 1653 1203
rect 1674 1186 1679 1206
rect 1621 1183 1679 1186
rect 1592 1176 1679 1183
rect 1704 1203 1741 1273
rect 2007 1272 2044 1273
rect 2794 1272 3208 1292
rect 3234 1272 3240 1294
rect 3466 1301 3473 1321
rect 3492 1301 3508 1321
rect 3466 1293 3508 1301
rect 3536 1321 3577 1323
rect 3536 1301 3550 1321
rect 3569 1301 3577 1321
rect 3536 1293 3577 1301
rect 3832 1297 3869 1298
rect 4135 1297 4172 1367
rect 4197 1387 4284 1394
rect 4197 1384 4255 1387
rect 4197 1364 4202 1384
rect 4223 1367 4255 1384
rect 4275 1367 4284 1387
rect 4223 1364 4284 1367
rect 4197 1357 4284 1364
rect 4343 1387 4380 1397
rect 4343 1367 4351 1387
rect 4371 1367 4380 1387
rect 4197 1356 4228 1357
rect 3831 1296 4172 1297
rect 3466 1287 3577 1293
rect 3756 1291 4172 1296
rect 2794 1266 3240 1272
rect 2794 1264 2962 1266
rect 1856 1213 1892 1214
rect 1704 1183 1713 1203
rect 1733 1183 1741 1203
rect 1592 1174 1648 1176
rect 1592 1173 1629 1174
rect 1704 1173 1741 1183
rect 1800 1203 1948 1213
rect 2048 1210 2144 1212
rect 1800 1183 1809 1203
rect 1829 1198 1919 1203
rect 1829 1183 1864 1198
rect 1800 1174 1864 1183
rect 1800 1173 1837 1174
rect 1856 1157 1864 1174
rect 1885 1183 1919 1198
rect 1939 1183 1948 1203
rect 1885 1174 1948 1183
rect 2006 1203 2144 1210
rect 2006 1183 2015 1203
rect 2035 1183 2144 1203
rect 2006 1174 2144 1183
rect 1885 1157 1892 1174
rect 1911 1173 1948 1174
rect 2007 1173 2044 1174
rect 1856 1122 1892 1157
rect 1327 1120 1368 1121
rect 265 1115 779 1116
rect 1219 1113 1368 1120
rect 1219 1093 1337 1113
rect 1357 1093 1368 1113
rect 1219 1085 1368 1093
rect 1435 1117 1794 1121
rect 1435 1112 1757 1117
rect 1435 1088 1548 1112
rect 1572 1093 1757 1112
rect 1781 1093 1794 1117
rect 1572 1088 1794 1093
rect 1435 1085 1794 1088
rect 1856 1085 1891 1122
rect 1959 1119 2059 1122
rect 1959 1115 2026 1119
rect 1959 1089 1971 1115
rect 1997 1093 2026 1115
rect 2052 1093 2059 1119
rect 1997 1089 2059 1093
rect 1959 1085 2059 1089
rect 113 1074 150 1075
rect 111 1066 151 1074
rect 111 1048 122 1066
rect 140 1048 151 1066
rect 1435 1064 1466 1085
rect 1856 1064 1892 1085
rect 1278 1063 1315 1064
rect 111 1000 151 1048
rect 1277 1054 1315 1063
rect 1277 1034 1286 1054
rect 1306 1034 1315 1054
rect 1277 1026 1315 1034
rect 1381 1058 1466 1064
rect 1491 1063 1528 1064
rect 1381 1038 1389 1058
rect 1409 1038 1466 1058
rect 1381 1030 1466 1038
rect 1490 1054 1528 1063
rect 1490 1034 1499 1054
rect 1519 1034 1528 1054
rect 1381 1029 1417 1030
rect 1490 1026 1528 1034
rect 1594 1058 1679 1064
rect 1699 1063 1736 1064
rect 1594 1038 1602 1058
rect 1622 1057 1679 1058
rect 1622 1038 1651 1057
rect 1594 1037 1651 1038
rect 1672 1037 1679 1057
rect 1594 1030 1679 1037
rect 1698 1054 1736 1063
rect 1698 1034 1707 1054
rect 1727 1034 1736 1054
rect 1594 1029 1630 1030
rect 1698 1026 1736 1034
rect 1802 1058 1946 1064
rect 1802 1038 1810 1058
rect 1830 1038 1918 1058
rect 1938 1038 1946 1058
rect 1802 1030 1946 1038
rect 1802 1029 1838 1030
rect 1910 1029 1946 1030
rect 2012 1063 2049 1064
rect 2012 1062 2050 1063
rect 2012 1054 2076 1062
rect 2012 1034 2021 1054
rect 2041 1040 2076 1054
rect 2096 1040 2099 1060
rect 2041 1035 2099 1040
rect 2041 1034 2076 1035
rect 422 1004 532 1018
rect 422 1001 465 1004
rect 111 993 236 1000
rect 422 996 426 1001
rect 111 974 203 993
rect 228 974 236 993
rect 111 964 236 974
rect 344 974 426 996
rect 455 974 465 1001
rect 493 977 500 1004
rect 529 996 532 1004
rect 1278 997 1315 1026
rect 529 977 594 996
rect 1279 995 1315 997
rect 1491 995 1528 1026
rect 1699 999 1736 1026
rect 2012 1022 2076 1034
rect 493 974 594 977
rect 344 972 594 974
rect 111 944 151 964
rect 110 935 151 944
rect 110 917 120 935
rect 138 917 151 935
rect 110 908 151 917
rect 110 907 147 908
rect 344 893 381 972
rect 422 959 532 972
rect 496 903 527 904
rect 344 873 353 893
rect 373 873 381 893
rect 344 863 381 873
rect 440 893 527 903
rect 440 873 449 893
rect 469 873 527 893
rect 440 864 527 873
rect 440 863 477 864
rect 113 841 150 845
rect 110 836 150 841
rect 110 818 122 836
rect 140 818 150 836
rect 110 638 150 818
rect 496 811 527 864
rect 557 893 594 972
rect 765 969 1158 989
rect 1178 969 1181 989
rect 1279 973 1528 995
rect 1697 994 1738 999
rect 2116 996 2143 1174
rect 2794 1086 2821 1264
rect 3199 1261 3240 1266
rect 3409 1265 3658 1287
rect 3756 1271 3759 1291
rect 3779 1271 4172 1291
rect 4343 1288 4380 1367
rect 4410 1396 4441 1449
rect 4787 1442 4827 1622
rect 5165 1782 5205 1962
rect 5551 1955 5582 2008
rect 5612 2037 5649 2116
rect 5820 2113 6213 2133
rect 6233 2113 6236 2133
rect 6334 2117 6583 2139
rect 6752 2138 6793 2143
rect 7171 2140 7198 2318
rect 7849 2230 7876 2408
rect 8254 2405 8295 2410
rect 8464 2409 8713 2431
rect 8811 2415 8814 2435
rect 8834 2415 9227 2435
rect 9398 2432 9435 2511
rect 9465 2540 9496 2593
rect 9842 2586 9882 2766
rect 10140 2849 10180 3029
rect 10526 3022 10557 3075
rect 10587 3104 10624 3183
rect 10795 3180 11188 3200
rect 11208 3180 11211 3200
rect 11309 3184 11558 3206
rect 11727 3205 11768 3210
rect 12146 3207 12173 3385
rect 12824 3297 12851 3475
rect 13229 3472 13270 3477
rect 13439 3476 13688 3498
rect 13786 3482 13789 3502
rect 13809 3482 14202 3502
rect 14373 3499 14410 3578
rect 14440 3607 14471 3660
rect 14817 3653 14857 3833
rect 15195 3993 15235 4173
rect 15581 4166 15612 4219
rect 15642 4248 15679 4327
rect 15850 4324 16243 4344
rect 16263 4324 16266 4344
rect 16364 4328 16613 4350
rect 16782 4349 16823 4354
rect 17201 4351 17228 4529
rect 17879 4441 17906 4619
rect 18284 4616 18325 4621
rect 18494 4620 18743 4642
rect 18841 4626 18844 4646
rect 18864 4626 19257 4646
rect 19428 4643 19465 4722
rect 19495 4751 19526 4804
rect 19872 4797 19912 4977
rect 19872 4779 19882 4797
rect 19900 4779 19912 4797
rect 19872 4774 19912 4779
rect 19872 4770 19909 4774
rect 19545 4751 19582 4752
rect 19495 4742 19582 4751
rect 19495 4722 19553 4742
rect 19573 4722 19582 4742
rect 19495 4712 19582 4722
rect 19641 4742 19678 4752
rect 19641 4722 19649 4742
rect 19669 4722 19678 4742
rect 19495 4711 19526 4712
rect 19490 4643 19600 4656
rect 19641 4643 19678 4722
rect 19875 4707 19912 4708
rect 19871 4698 19912 4707
rect 19871 4680 19884 4698
rect 19902 4680 19912 4698
rect 19871 4671 19912 4680
rect 19871 4651 19911 4671
rect 19428 4641 19678 4643
rect 19428 4638 19529 4641
rect 17946 4581 18010 4593
rect 18286 4589 18323 4616
rect 18494 4589 18531 4620
rect 18707 4618 18743 4620
rect 19428 4619 19493 4638
rect 18707 4589 18744 4618
rect 19490 4611 19493 4619
rect 19522 4611 19529 4638
rect 19557 4614 19567 4641
rect 19596 4619 19678 4641
rect 19786 4641 19911 4651
rect 19786 4622 19794 4641
rect 19819 4622 19911 4641
rect 19596 4614 19600 4619
rect 19786 4615 19911 4622
rect 19557 4611 19600 4614
rect 19490 4597 19600 4611
rect 17946 4580 17981 4581
rect 17923 4575 17981 4580
rect 17923 4555 17926 4575
rect 17946 4561 17981 4575
rect 18001 4561 18010 4581
rect 17946 4553 18010 4561
rect 17972 4552 18010 4553
rect 17973 4551 18010 4552
rect 18076 4585 18112 4586
rect 18184 4585 18220 4586
rect 18076 4577 18220 4585
rect 18076 4557 18084 4577
rect 18104 4557 18192 4577
rect 18212 4557 18220 4577
rect 18076 4551 18220 4557
rect 18286 4581 18324 4589
rect 18392 4585 18428 4586
rect 18286 4561 18295 4581
rect 18315 4561 18324 4581
rect 18286 4552 18324 4561
rect 18343 4578 18428 4585
rect 18343 4558 18350 4578
rect 18371 4577 18428 4578
rect 18371 4558 18400 4577
rect 18343 4557 18400 4558
rect 18420 4557 18428 4577
rect 18286 4551 18323 4552
rect 18343 4551 18428 4557
rect 18494 4581 18532 4589
rect 18605 4585 18641 4586
rect 18494 4561 18503 4581
rect 18523 4561 18532 4581
rect 18494 4552 18532 4561
rect 18556 4577 18641 4585
rect 18556 4557 18613 4577
rect 18633 4557 18641 4577
rect 18494 4551 18531 4552
rect 18556 4551 18641 4557
rect 18707 4581 18745 4589
rect 18707 4561 18716 4581
rect 18736 4561 18745 4581
rect 18707 4552 18745 4561
rect 19871 4567 19911 4615
rect 18707 4551 18744 4552
rect 18130 4530 18166 4551
rect 18556 4530 18587 4551
rect 19871 4549 19882 4567
rect 19900 4549 19911 4567
rect 19871 4541 19911 4549
rect 19872 4540 19909 4541
rect 17963 4526 18063 4530
rect 17963 4522 18025 4526
rect 17963 4496 17970 4522
rect 17996 4500 18025 4522
rect 18051 4500 18063 4526
rect 17996 4496 18063 4500
rect 17963 4493 18063 4496
rect 18131 4493 18166 4530
rect 18228 4527 18587 4530
rect 18228 4522 18450 4527
rect 18228 4498 18241 4522
rect 18265 4503 18450 4522
rect 18474 4503 18587 4527
rect 18265 4498 18587 4503
rect 18228 4494 18587 4498
rect 18654 4522 18803 4530
rect 18654 4502 18665 4522
rect 18685 4502 18803 4522
rect 18654 4495 18803 4502
rect 19243 4499 19757 4500
rect 18654 4494 18695 4495
rect 18130 4458 18166 4493
rect 17978 4441 18015 4442
rect 18074 4441 18111 4442
rect 18130 4441 18137 4458
rect 17878 4432 18016 4441
rect 17878 4412 17987 4432
rect 18007 4412 18016 4432
rect 17878 4405 18016 4412
rect 18074 4432 18137 4441
rect 18074 4412 18083 4432
rect 18103 4417 18137 4432
rect 18158 4441 18166 4458
rect 18185 4441 18222 4442
rect 18158 4432 18222 4441
rect 18158 4417 18193 4432
rect 18103 4412 18193 4417
rect 18213 4412 18222 4432
rect 17878 4403 17974 4405
rect 18074 4402 18222 4412
rect 18281 4432 18318 4442
rect 18393 4441 18430 4442
rect 18374 4439 18430 4441
rect 18281 4412 18289 4432
rect 18309 4412 18318 4432
rect 18130 4401 18166 4402
rect 17060 4349 17228 4351
rect 16782 4343 17228 4349
rect 15850 4319 16266 4324
rect 16445 4322 16556 4328
rect 15850 4318 16191 4319
rect 15794 4258 15825 4259
rect 15642 4228 15651 4248
rect 15671 4228 15679 4248
rect 15642 4218 15679 4228
rect 15738 4251 15825 4258
rect 15738 4248 15799 4251
rect 15738 4228 15747 4248
rect 15767 4231 15799 4248
rect 15820 4231 15825 4251
rect 15767 4228 15825 4231
rect 15738 4221 15825 4228
rect 15850 4248 15887 4318
rect 16153 4317 16190 4318
rect 16445 4314 16486 4322
rect 16445 4294 16453 4314
rect 16472 4294 16486 4314
rect 16445 4292 16486 4294
rect 16514 4314 16556 4322
rect 16514 4294 16530 4314
rect 16549 4294 16556 4314
rect 16782 4321 16788 4343
rect 16814 4323 17228 4343
rect 17978 4342 18015 4343
rect 18281 4342 18318 4412
rect 18343 4432 18430 4439
rect 18343 4429 18401 4432
rect 18343 4409 18348 4429
rect 18369 4412 18401 4429
rect 18421 4412 18430 4432
rect 18369 4409 18430 4412
rect 18343 4402 18430 4409
rect 18489 4432 18526 4442
rect 18489 4412 18497 4432
rect 18517 4412 18526 4432
rect 18343 4401 18374 4402
rect 17977 4341 18318 4342
rect 16814 4321 16823 4323
rect 17060 4322 17228 4323
rect 17902 4340 18318 4341
rect 17902 4336 18278 4340
rect 16782 4312 16823 4321
rect 17902 4316 17905 4336
rect 17925 4323 18278 4336
rect 18310 4323 18318 4340
rect 17925 4316 18318 4323
rect 18489 4333 18526 4412
rect 18556 4441 18587 4494
rect 19224 4483 19757 4499
rect 19224 4472 19756 4483
rect 19875 4474 19912 4478
rect 18606 4441 18643 4442
rect 18556 4432 18643 4441
rect 18556 4412 18614 4432
rect 18634 4412 18643 4432
rect 18556 4402 18643 4412
rect 18702 4432 18739 4442
rect 18702 4412 18710 4432
rect 18730 4412 18739 4432
rect 18556 4401 18587 4402
rect 18551 4333 18661 4346
rect 18702 4333 18739 4412
rect 18489 4331 18739 4333
rect 18489 4328 18590 4331
rect 18489 4309 18554 4328
rect 16514 4292 16556 4294
rect 16445 4277 16556 4292
rect 18551 4301 18554 4309
rect 18583 4301 18590 4328
rect 18618 4304 18628 4331
rect 18657 4309 18739 4331
rect 18817 4403 18985 4404
rect 19224 4403 19262 4472
rect 18817 4383 19262 4403
rect 19489 4434 19600 4449
rect 19489 4432 19531 4434
rect 19489 4412 19496 4432
rect 19515 4412 19531 4432
rect 19489 4404 19531 4412
rect 19559 4432 19600 4434
rect 19559 4412 19573 4432
rect 19592 4412 19600 4432
rect 19559 4404 19600 4412
rect 19489 4398 19600 4404
rect 19722 4409 19756 4472
rect 19874 4468 19912 4474
rect 19874 4450 19884 4468
rect 19902 4450 19912 4468
rect 19874 4441 19912 4450
rect 19874 4409 19908 4441
rect 18817 4377 19261 4383
rect 18817 4375 18985 4377
rect 18657 4304 18661 4309
rect 18618 4301 18661 4304
rect 18551 4287 18661 4301
rect 16002 4258 16038 4259
rect 15850 4228 15859 4248
rect 15879 4228 15887 4248
rect 15738 4219 15794 4221
rect 15738 4218 15775 4219
rect 15850 4218 15887 4228
rect 15946 4248 16094 4258
rect 16194 4255 16290 4257
rect 15946 4228 15955 4248
rect 15975 4228 16065 4248
rect 16085 4228 16094 4248
rect 15946 4219 16094 4228
rect 16152 4248 16290 4255
rect 16152 4228 16161 4248
rect 16181 4228 16290 4248
rect 16152 4219 16290 4228
rect 15946 4218 15983 4219
rect 16002 4167 16038 4219
rect 16057 4218 16094 4219
rect 16153 4218 16190 4219
rect 15473 4165 15514 4166
rect 15365 4158 15514 4165
rect 15365 4138 15483 4158
rect 15503 4138 15514 4158
rect 15365 4130 15514 4138
rect 15581 4162 15940 4166
rect 15581 4157 15903 4162
rect 15581 4133 15694 4157
rect 15718 4138 15903 4157
rect 15927 4138 15940 4162
rect 15718 4133 15940 4138
rect 15581 4130 15940 4133
rect 16002 4130 16037 4167
rect 16105 4164 16205 4167
rect 16105 4160 16172 4164
rect 16105 4134 16117 4160
rect 16143 4138 16172 4160
rect 16198 4138 16205 4164
rect 16143 4134 16205 4138
rect 16105 4130 16205 4134
rect 15581 4109 15612 4130
rect 16002 4109 16038 4130
rect 15424 4108 15461 4109
rect 15423 4099 15461 4108
rect 15423 4079 15432 4099
rect 15452 4079 15461 4099
rect 15423 4071 15461 4079
rect 15527 4103 15612 4109
rect 15637 4108 15674 4109
rect 15527 4083 15535 4103
rect 15555 4083 15612 4103
rect 15527 4075 15612 4083
rect 15636 4099 15674 4108
rect 15636 4079 15645 4099
rect 15665 4079 15674 4099
rect 15527 4074 15563 4075
rect 15636 4071 15674 4079
rect 15740 4103 15825 4109
rect 15845 4108 15882 4109
rect 15740 4083 15748 4103
rect 15768 4102 15825 4103
rect 15768 4083 15797 4102
rect 15740 4082 15797 4083
rect 15818 4082 15825 4102
rect 15740 4075 15825 4082
rect 15844 4099 15882 4108
rect 15844 4079 15853 4099
rect 15873 4079 15882 4099
rect 15740 4074 15776 4075
rect 15844 4071 15882 4079
rect 15948 4103 16092 4109
rect 15948 4083 15956 4103
rect 15976 4100 16064 4103
rect 15976 4083 16007 4100
rect 15948 4080 16007 4083
rect 16030 4083 16064 4100
rect 16084 4083 16092 4103
rect 16030 4080 16092 4083
rect 15948 4075 16092 4080
rect 15948 4074 15984 4075
rect 16056 4074 16092 4075
rect 16158 4108 16195 4109
rect 16158 4107 16196 4108
rect 16158 4099 16222 4107
rect 16158 4079 16167 4099
rect 16187 4085 16222 4099
rect 16242 4085 16245 4105
rect 16187 4080 16245 4085
rect 16187 4079 16222 4080
rect 15424 4042 15461 4071
rect 15425 4040 15461 4042
rect 15637 4040 15674 4071
rect 15425 4018 15674 4040
rect 15845 4039 15882 4071
rect 16158 4067 16222 4079
rect 16262 4041 16289 4219
rect 18817 4197 18844 4375
rect 18884 4337 18948 4349
rect 19224 4345 19261 4377
rect 19432 4376 19681 4398
rect 19722 4377 19908 4409
rect 19736 4376 19908 4377
rect 19432 4345 19469 4376
rect 19645 4374 19681 4376
rect 19645 4345 19682 4374
rect 19874 4348 19908 4376
rect 18884 4336 18919 4337
rect 18861 4331 18919 4336
rect 18861 4311 18864 4331
rect 18884 4317 18919 4331
rect 18939 4317 18948 4337
rect 18884 4309 18948 4317
rect 18910 4308 18948 4309
rect 18911 4307 18948 4308
rect 19014 4341 19050 4342
rect 19122 4341 19158 4342
rect 19014 4334 19158 4341
rect 19014 4333 19074 4334
rect 19014 4313 19022 4333
rect 19042 4314 19074 4333
rect 19099 4333 19158 4334
rect 19099 4314 19130 4333
rect 19042 4313 19130 4314
rect 19150 4313 19158 4333
rect 19014 4307 19158 4313
rect 19224 4337 19262 4345
rect 19330 4341 19366 4342
rect 19224 4317 19233 4337
rect 19253 4317 19262 4337
rect 19224 4308 19262 4317
rect 19281 4334 19366 4341
rect 19281 4314 19288 4334
rect 19309 4333 19366 4334
rect 19309 4314 19338 4333
rect 19281 4313 19338 4314
rect 19358 4313 19366 4333
rect 19224 4307 19261 4308
rect 19281 4307 19366 4313
rect 19432 4337 19470 4345
rect 19543 4341 19579 4342
rect 19432 4317 19441 4337
rect 19461 4317 19470 4337
rect 19432 4308 19470 4317
rect 19494 4333 19579 4341
rect 19494 4313 19551 4333
rect 19571 4313 19579 4333
rect 19432 4307 19469 4308
rect 19494 4307 19579 4313
rect 19645 4337 19683 4345
rect 19645 4317 19654 4337
rect 19674 4317 19683 4337
rect 19645 4308 19683 4317
rect 19872 4338 19909 4348
rect 19872 4320 19882 4338
rect 19900 4320 19909 4338
rect 19872 4311 19909 4320
rect 19874 4310 19908 4311
rect 19645 4307 19682 4308
rect 19068 4286 19104 4307
rect 19494 4286 19525 4307
rect 18901 4282 19001 4286
rect 18901 4278 18963 4282
rect 18901 4252 18908 4278
rect 18934 4256 18963 4278
rect 18989 4256 19001 4282
rect 18934 4252 19001 4256
rect 18901 4249 19001 4252
rect 19069 4249 19104 4286
rect 19166 4283 19525 4286
rect 19166 4278 19388 4283
rect 19166 4254 19179 4278
rect 19203 4259 19388 4278
rect 19412 4259 19525 4283
rect 19203 4254 19525 4259
rect 19166 4250 19525 4254
rect 19592 4278 19741 4286
rect 19592 4258 19603 4278
rect 19623 4258 19741 4278
rect 19592 4251 19741 4258
rect 19592 4250 19633 4251
rect 18916 4197 18953 4198
rect 19012 4197 19049 4198
rect 19068 4197 19104 4249
rect 19123 4197 19160 4198
rect 18816 4188 18954 4197
rect 18411 4167 18522 4182
rect 18411 4165 18453 4167
rect 18081 4144 18186 4146
rect 17737 4136 17907 4137
rect 18081 4136 18130 4144
rect 17737 4117 18130 4136
rect 18161 4117 18186 4144
rect 18411 4145 18418 4165
rect 18437 4145 18453 4165
rect 18411 4137 18453 4145
rect 18481 4165 18522 4167
rect 18481 4145 18495 4165
rect 18514 4145 18522 4165
rect 18816 4168 18925 4188
rect 18945 4168 18954 4188
rect 18816 4161 18954 4168
rect 19012 4188 19160 4197
rect 19012 4168 19021 4188
rect 19041 4168 19131 4188
rect 19151 4168 19160 4188
rect 18816 4159 18912 4161
rect 19012 4158 19160 4168
rect 19219 4188 19256 4198
rect 19331 4197 19368 4198
rect 19312 4195 19368 4197
rect 19219 4168 19227 4188
rect 19247 4168 19256 4188
rect 19068 4157 19104 4158
rect 18481 4137 18522 4145
rect 18411 4131 18522 4137
rect 17737 4110 18186 4117
rect 17737 4108 17907 4110
rect 16587 4077 16697 4091
rect 16587 4074 16630 4077
rect 16587 4069 16591 4074
rect 16121 4039 16289 4041
rect 15845 4036 16289 4039
rect 15506 4012 15617 4018
rect 15506 4004 15547 4012
rect 15195 3949 15234 3993
rect 15506 3984 15514 4004
rect 15533 3984 15547 4004
rect 15506 3982 15547 3984
rect 15575 4004 15617 4012
rect 15575 3984 15591 4004
rect 15610 3984 15617 4004
rect 15575 3982 15617 3984
rect 15506 3967 15617 3982
rect 15843 4013 16289 4036
rect 15195 3925 15235 3949
rect 15535 3925 15582 3927
rect 15843 3925 15881 4013
rect 16121 4012 16289 4013
rect 16509 4047 16591 4069
rect 16620 4047 16630 4074
rect 16658 4050 16665 4077
rect 16694 4069 16697 4077
rect 16694 4050 16759 4069
rect 16658 4047 16759 4050
rect 16509 4045 16759 4047
rect 16509 3966 16546 4045
rect 16587 4032 16697 4045
rect 16661 3976 16692 3977
rect 16509 3946 16518 3966
rect 16538 3946 16546 3966
rect 16509 3936 16546 3946
rect 16605 3966 16692 3976
rect 16605 3946 16614 3966
rect 16634 3946 16692 3966
rect 16605 3937 16692 3946
rect 16605 3936 16642 3937
rect 15195 3892 15881 3925
rect 15195 3835 15234 3892
rect 15843 3890 15881 3892
rect 16661 3884 16692 3937
rect 16722 3966 16759 4045
rect 16930 4058 17323 4062
rect 16930 4041 16949 4058
rect 16969 4042 17323 4058
rect 17343 4042 17346 4062
rect 16969 4041 17346 4042
rect 16930 4037 17346 4041
rect 16930 4036 17271 4037
rect 16874 3976 16905 3977
rect 16722 3946 16731 3966
rect 16751 3946 16759 3966
rect 16722 3936 16759 3946
rect 16818 3969 16905 3976
rect 16818 3966 16879 3969
rect 16818 3946 16827 3966
rect 16847 3949 16879 3966
rect 16900 3949 16905 3969
rect 16847 3946 16905 3949
rect 16818 3939 16905 3946
rect 16930 3966 16967 4036
rect 17233 4035 17270 4036
rect 17082 3976 17118 3977
rect 16930 3946 16939 3966
rect 16959 3946 16967 3966
rect 16818 3937 16874 3939
rect 16818 3936 16855 3937
rect 16930 3936 16967 3946
rect 17026 3966 17174 3976
rect 17274 3973 17370 3975
rect 17026 3946 17035 3966
rect 17055 3946 17145 3966
rect 17165 3946 17174 3966
rect 17026 3937 17174 3946
rect 17232 3966 17370 3973
rect 17232 3946 17241 3966
rect 17261 3946 17370 3966
rect 17232 3937 17370 3946
rect 17026 3936 17063 3937
rect 17082 3885 17118 3937
rect 17137 3936 17174 3937
rect 17233 3936 17270 3937
rect 16553 3883 16594 3884
rect 16445 3876 16594 3883
rect 16445 3856 16563 3876
rect 16583 3856 16594 3876
rect 16445 3848 16594 3856
rect 16661 3880 17020 3884
rect 16661 3875 16983 3880
rect 16661 3851 16774 3875
rect 16798 3856 16983 3875
rect 17007 3856 17020 3880
rect 16798 3851 17020 3856
rect 16661 3848 17020 3851
rect 17082 3848 17117 3885
rect 17185 3882 17285 3885
rect 17185 3878 17252 3882
rect 17185 3852 17197 3878
rect 17223 3856 17252 3878
rect 17278 3856 17285 3882
rect 17223 3852 17285 3856
rect 17185 3848 17285 3852
rect 15195 3833 15243 3835
rect 15195 3815 15206 3833
rect 15224 3815 15243 3833
rect 16661 3827 16692 3848
rect 17082 3827 17118 3848
rect 16504 3826 16541 3827
rect 15195 3806 15243 3815
rect 15196 3805 15243 3806
rect 15509 3810 15619 3824
rect 15509 3807 15552 3810
rect 15509 3802 15513 3807
rect 15431 3780 15513 3802
rect 15542 3780 15552 3807
rect 15580 3783 15587 3810
rect 15616 3802 15619 3810
rect 16503 3817 16541 3826
rect 15616 3783 15681 3802
rect 16503 3797 16512 3817
rect 16532 3797 16541 3817
rect 15580 3780 15681 3783
rect 15431 3778 15681 3780
rect 15199 3742 15236 3743
rect 14817 3635 14827 3653
rect 14845 3635 14857 3653
rect 14817 3630 14857 3635
rect 15195 3739 15236 3742
rect 15195 3734 15237 3739
rect 15195 3716 15208 3734
rect 15226 3716 15237 3734
rect 15195 3702 15237 3716
rect 15275 3702 15322 3706
rect 15195 3696 15322 3702
rect 15195 3667 15283 3696
rect 15312 3667 15322 3696
rect 15431 3699 15468 3778
rect 15509 3765 15619 3778
rect 15583 3709 15614 3710
rect 15431 3679 15440 3699
rect 15460 3679 15468 3699
rect 15431 3669 15468 3679
rect 15527 3699 15614 3709
rect 15527 3679 15536 3699
rect 15556 3679 15614 3699
rect 15527 3670 15614 3679
rect 15527 3669 15564 3670
rect 15195 3663 15322 3667
rect 15195 3646 15234 3663
rect 15275 3662 15322 3663
rect 14817 3626 14854 3630
rect 15195 3628 15206 3646
rect 15224 3628 15234 3646
rect 15195 3619 15234 3628
rect 15196 3618 15233 3619
rect 15583 3617 15614 3670
rect 15644 3699 15681 3778
rect 15852 3775 16245 3795
rect 16265 3775 16268 3795
rect 16503 3789 16541 3797
rect 16607 3821 16692 3827
rect 16717 3826 16754 3827
rect 16607 3801 16615 3821
rect 16635 3801 16692 3821
rect 16607 3793 16692 3801
rect 16716 3817 16754 3826
rect 16716 3797 16725 3817
rect 16745 3797 16754 3817
rect 16607 3792 16643 3793
rect 16716 3789 16754 3797
rect 16820 3821 16905 3827
rect 16925 3826 16962 3827
rect 16820 3801 16828 3821
rect 16848 3820 16905 3821
rect 16848 3801 16877 3820
rect 16820 3800 16877 3801
rect 16898 3800 16905 3820
rect 16820 3793 16905 3800
rect 16924 3817 16962 3826
rect 16924 3797 16933 3817
rect 16953 3797 16962 3817
rect 16820 3792 16856 3793
rect 16924 3789 16962 3797
rect 17028 3821 17172 3827
rect 17028 3801 17036 3821
rect 17056 3819 17144 3821
rect 17056 3801 17085 3819
rect 17028 3798 17085 3801
rect 17112 3801 17144 3819
rect 17164 3801 17172 3821
rect 17112 3798 17172 3801
rect 17028 3793 17172 3798
rect 17028 3792 17064 3793
rect 17136 3792 17172 3793
rect 17238 3826 17275 3827
rect 17238 3825 17276 3826
rect 17238 3817 17302 3825
rect 17238 3797 17247 3817
rect 17267 3803 17302 3817
rect 17322 3803 17325 3823
rect 17267 3798 17325 3803
rect 17267 3797 17302 3798
rect 15852 3770 16268 3775
rect 15852 3769 16193 3770
rect 15796 3709 15827 3710
rect 15644 3679 15653 3699
rect 15673 3679 15681 3699
rect 15644 3669 15681 3679
rect 15740 3702 15827 3709
rect 15740 3699 15801 3702
rect 15740 3679 15749 3699
rect 15769 3682 15801 3699
rect 15822 3682 15827 3702
rect 15769 3679 15827 3682
rect 15740 3672 15827 3679
rect 15852 3699 15889 3769
rect 16155 3768 16192 3769
rect 16504 3760 16541 3789
rect 16505 3758 16541 3760
rect 16717 3758 16754 3789
rect 16505 3736 16754 3758
rect 16925 3757 16962 3789
rect 17238 3785 17302 3797
rect 17342 3759 17369 3937
rect 17737 3930 17766 4108
rect 17806 4070 17870 4082
rect 18146 4078 18183 4110
rect 18354 4109 18603 4131
rect 18354 4078 18391 4109
rect 18567 4107 18603 4109
rect 18567 4078 18604 4107
rect 18916 4098 18953 4099
rect 19219 4098 19256 4168
rect 19281 4188 19368 4195
rect 19281 4185 19339 4188
rect 19281 4165 19286 4185
rect 19307 4168 19339 4185
rect 19359 4168 19368 4188
rect 19307 4165 19368 4168
rect 19281 4158 19368 4165
rect 19427 4188 19464 4198
rect 19427 4168 19435 4188
rect 19455 4168 19464 4188
rect 19281 4157 19312 4158
rect 18915 4097 19256 4098
rect 18840 4092 19256 4097
rect 17806 4069 17841 4070
rect 17783 4064 17841 4069
rect 17783 4044 17786 4064
rect 17806 4050 17841 4064
rect 17861 4050 17870 4070
rect 17806 4042 17870 4050
rect 17832 4041 17870 4042
rect 17833 4040 17870 4041
rect 17936 4074 17972 4075
rect 18044 4074 18080 4075
rect 17936 4066 18080 4074
rect 17936 4046 17944 4066
rect 17964 4046 18052 4066
rect 18072 4046 18080 4066
rect 17936 4040 18080 4046
rect 18146 4070 18184 4078
rect 18252 4074 18288 4075
rect 18146 4050 18155 4070
rect 18175 4050 18184 4070
rect 18146 4041 18184 4050
rect 18203 4067 18288 4074
rect 18203 4047 18210 4067
rect 18231 4066 18288 4067
rect 18231 4047 18260 4066
rect 18203 4046 18260 4047
rect 18280 4046 18288 4066
rect 18146 4040 18183 4041
rect 18203 4040 18288 4046
rect 18354 4070 18392 4078
rect 18465 4074 18501 4075
rect 18354 4050 18363 4070
rect 18383 4050 18392 4070
rect 18354 4041 18392 4050
rect 18416 4066 18501 4074
rect 18416 4046 18473 4066
rect 18493 4046 18501 4066
rect 18354 4040 18391 4041
rect 18416 4040 18501 4046
rect 18567 4070 18605 4078
rect 18840 4072 18843 4092
rect 18863 4072 19256 4092
rect 19427 4089 19464 4168
rect 19494 4197 19525 4250
rect 19875 4248 19912 4249
rect 19874 4239 19913 4248
rect 19874 4221 19884 4239
rect 19902 4221 19913 4239
rect 19786 4204 19833 4205
rect 19874 4204 19913 4221
rect 19786 4200 19913 4204
rect 19544 4197 19581 4198
rect 19494 4188 19581 4197
rect 19494 4168 19552 4188
rect 19572 4168 19581 4188
rect 19494 4158 19581 4168
rect 19640 4188 19677 4198
rect 19640 4168 19648 4188
rect 19668 4168 19677 4188
rect 19494 4157 19525 4158
rect 19489 4089 19599 4102
rect 19640 4089 19677 4168
rect 19786 4171 19796 4200
rect 19825 4171 19913 4200
rect 19786 4165 19913 4171
rect 19786 4161 19833 4165
rect 19871 4151 19913 4165
rect 19871 4133 19882 4151
rect 19900 4133 19913 4151
rect 19871 4128 19913 4133
rect 19872 4125 19913 4128
rect 19872 4124 19909 4125
rect 19427 4087 19677 4089
rect 19427 4084 19528 4087
rect 18567 4050 18576 4070
rect 18596 4050 18605 4070
rect 19427 4065 19492 4084
rect 18567 4041 18605 4050
rect 19489 4057 19492 4065
rect 19521 4057 19528 4084
rect 19556 4060 19566 4087
rect 19595 4065 19677 4087
rect 19595 4060 19599 4065
rect 19556 4057 19599 4060
rect 19489 4043 19599 4057
rect 19865 4061 19912 4062
rect 19865 4052 19913 4061
rect 18567 4040 18604 4041
rect 17990 4019 18026 4040
rect 18416 4019 18447 4040
rect 19865 4034 19884 4052
rect 19902 4034 19913 4052
rect 19865 4032 19913 4034
rect 17823 4015 17923 4019
rect 17823 4011 17885 4015
rect 17823 3985 17830 4011
rect 17856 3989 17885 4011
rect 17911 3989 17923 4015
rect 17856 3985 17923 3989
rect 17823 3982 17923 3985
rect 17991 3982 18026 4019
rect 18088 4016 18447 4019
rect 18088 4011 18310 4016
rect 18088 3987 18101 4011
rect 18125 3992 18310 4011
rect 18334 3992 18447 4016
rect 18125 3987 18447 3992
rect 18088 3983 18447 3987
rect 18514 4011 18663 4019
rect 18514 3991 18525 4011
rect 18545 3991 18663 4011
rect 18514 3984 18663 3991
rect 18514 3983 18555 3984
rect 17990 3943 18026 3982
rect 17838 3930 17875 3931
rect 17934 3930 17971 3931
rect 17990 3930 17997 3943
rect 17737 3921 17876 3930
rect 17737 3901 17847 3921
rect 17867 3901 17876 3921
rect 17737 3894 17876 3901
rect 17934 3921 17997 3930
rect 17934 3901 17943 3921
rect 17963 3905 17997 3921
rect 18020 3930 18026 3943
rect 18045 3930 18082 3931
rect 18020 3921 18082 3930
rect 18020 3905 18053 3921
rect 17963 3901 18053 3905
rect 18073 3901 18082 3921
rect 17737 3892 17834 3894
rect 17737 3891 17766 3892
rect 17934 3891 18082 3901
rect 18141 3921 18178 3931
rect 18253 3930 18290 3931
rect 18234 3928 18290 3930
rect 18141 3901 18149 3921
rect 18169 3901 18178 3921
rect 17990 3890 18026 3891
rect 17838 3831 17875 3832
rect 18141 3831 18178 3901
rect 18203 3921 18290 3928
rect 18203 3918 18261 3921
rect 18203 3898 18208 3918
rect 18229 3901 18261 3918
rect 18281 3901 18290 3921
rect 18229 3898 18290 3901
rect 18203 3891 18290 3898
rect 18349 3921 18386 3931
rect 18349 3901 18357 3921
rect 18377 3901 18386 3921
rect 18203 3890 18234 3891
rect 17837 3830 18178 3831
rect 17762 3826 18178 3830
rect 17762 3825 18139 3826
rect 17762 3805 17765 3825
rect 17785 3809 18139 3825
rect 18159 3809 18178 3826
rect 17785 3805 18178 3809
rect 18349 3822 18386 3901
rect 18416 3930 18447 3983
rect 19227 3975 19265 3977
rect 19874 3975 19913 4032
rect 19227 3942 19913 3975
rect 18466 3930 18503 3931
rect 18416 3921 18503 3930
rect 18416 3901 18474 3921
rect 18494 3901 18503 3921
rect 18416 3891 18503 3901
rect 18562 3921 18599 3931
rect 18562 3901 18570 3921
rect 18590 3901 18599 3921
rect 18416 3890 18447 3891
rect 18411 3822 18521 3835
rect 18562 3822 18599 3901
rect 18349 3820 18599 3822
rect 18349 3817 18450 3820
rect 18349 3798 18414 3817
rect 18411 3790 18414 3798
rect 18443 3790 18450 3817
rect 18478 3793 18488 3820
rect 18517 3798 18599 3820
rect 18819 3854 18987 3855
rect 19227 3854 19265 3942
rect 19526 3940 19573 3942
rect 19873 3918 19913 3942
rect 18819 3831 19265 3854
rect 19491 3885 19602 3900
rect 19491 3883 19533 3885
rect 19491 3863 19498 3883
rect 19517 3863 19533 3883
rect 19491 3855 19533 3863
rect 19561 3883 19602 3885
rect 19561 3863 19575 3883
rect 19594 3863 19602 3883
rect 19874 3874 19913 3918
rect 19561 3855 19602 3863
rect 19491 3849 19602 3855
rect 18819 3828 19263 3831
rect 18819 3826 18987 3828
rect 18517 3793 18521 3798
rect 18478 3790 18521 3793
rect 18411 3776 18521 3790
rect 17201 3757 17369 3759
rect 16922 3750 17369 3757
rect 16586 3730 16697 3736
rect 16586 3722 16627 3730
rect 16004 3709 16040 3710
rect 15852 3679 15861 3699
rect 15881 3679 15889 3699
rect 15740 3670 15796 3672
rect 15740 3669 15777 3670
rect 15852 3669 15889 3679
rect 15948 3699 16096 3709
rect 16196 3706 16292 3708
rect 15948 3679 15957 3699
rect 15977 3679 16067 3699
rect 16087 3679 16096 3699
rect 15948 3670 16096 3679
rect 16154 3699 16292 3706
rect 16154 3679 16163 3699
rect 16183 3679 16292 3699
rect 16586 3702 16594 3722
rect 16613 3702 16627 3722
rect 16586 3700 16627 3702
rect 16655 3722 16697 3730
rect 16655 3702 16671 3722
rect 16690 3702 16697 3722
rect 16922 3723 16947 3750
rect 16978 3731 17369 3750
rect 16978 3723 17027 3731
rect 17201 3730 17369 3731
rect 16922 3721 17027 3723
rect 16655 3700 16697 3702
rect 16586 3685 16697 3700
rect 16154 3670 16292 3679
rect 15948 3669 15985 3670
rect 16004 3618 16040 3670
rect 16059 3669 16096 3670
rect 16155 3669 16192 3670
rect 15475 3616 15516 3617
rect 15367 3609 15516 3616
rect 14490 3607 14527 3608
rect 14440 3598 14527 3607
rect 14440 3578 14498 3598
rect 14518 3578 14527 3598
rect 14440 3568 14527 3578
rect 14586 3598 14623 3608
rect 14586 3578 14594 3598
rect 14614 3578 14623 3598
rect 15367 3589 15485 3609
rect 15505 3589 15516 3609
rect 15367 3581 15516 3589
rect 15583 3613 15942 3617
rect 15583 3608 15905 3613
rect 15583 3584 15696 3608
rect 15720 3589 15905 3608
rect 15929 3589 15942 3613
rect 15720 3584 15942 3589
rect 15583 3581 15942 3584
rect 16004 3581 16039 3618
rect 16107 3615 16207 3618
rect 16107 3611 16174 3615
rect 16107 3585 16119 3611
rect 16145 3589 16174 3611
rect 16200 3589 16207 3615
rect 16145 3585 16207 3589
rect 16107 3581 16207 3585
rect 14440 3567 14471 3568
rect 14435 3499 14545 3512
rect 14586 3499 14623 3578
rect 14820 3563 14857 3564
rect 14816 3554 14857 3563
rect 15583 3560 15614 3581
rect 16004 3560 16040 3581
rect 15426 3559 15463 3560
rect 15200 3556 15234 3557
rect 14816 3536 14829 3554
rect 14847 3536 14857 3554
rect 14816 3527 14857 3536
rect 15199 3547 15236 3556
rect 15199 3529 15208 3547
rect 15226 3529 15236 3547
rect 14816 3507 14856 3527
rect 15199 3519 15236 3529
rect 15425 3550 15463 3559
rect 15425 3530 15434 3550
rect 15454 3530 15463 3550
rect 15425 3522 15463 3530
rect 15529 3554 15614 3560
rect 15639 3559 15676 3560
rect 15529 3534 15537 3554
rect 15557 3534 15614 3554
rect 15529 3526 15614 3534
rect 15638 3550 15676 3559
rect 15638 3530 15647 3550
rect 15667 3530 15676 3550
rect 15529 3525 15565 3526
rect 15638 3522 15676 3530
rect 15742 3554 15827 3560
rect 15847 3559 15884 3560
rect 15742 3534 15750 3554
rect 15770 3553 15827 3554
rect 15770 3534 15799 3553
rect 15742 3533 15799 3534
rect 15820 3533 15827 3553
rect 15742 3526 15827 3533
rect 15846 3550 15884 3559
rect 15846 3530 15855 3550
rect 15875 3530 15884 3550
rect 15742 3525 15778 3526
rect 15846 3522 15884 3530
rect 15950 3554 16094 3560
rect 15950 3534 15958 3554
rect 15978 3553 16066 3554
rect 15978 3534 16009 3553
rect 15950 3533 16009 3534
rect 16034 3534 16066 3553
rect 16086 3534 16094 3554
rect 16034 3533 16094 3534
rect 15950 3526 16094 3533
rect 15950 3525 15986 3526
rect 16058 3525 16094 3526
rect 16160 3559 16197 3560
rect 16160 3558 16198 3559
rect 16160 3550 16224 3558
rect 16160 3530 16169 3550
rect 16189 3536 16224 3550
rect 16244 3536 16247 3556
rect 16189 3531 16247 3536
rect 16189 3530 16224 3531
rect 14373 3497 14623 3499
rect 14373 3494 14474 3497
rect 12891 3437 12955 3449
rect 13231 3445 13268 3472
rect 13439 3445 13476 3476
rect 13652 3474 13688 3476
rect 14373 3475 14438 3494
rect 13652 3445 13689 3474
rect 14435 3467 14438 3475
rect 14467 3467 14474 3494
rect 14502 3470 14512 3497
rect 14541 3475 14623 3497
rect 14731 3497 14856 3507
rect 14731 3478 14739 3497
rect 14764 3478 14856 3497
rect 14541 3470 14545 3475
rect 14731 3471 14856 3478
rect 14502 3467 14545 3470
rect 14435 3453 14545 3467
rect 12891 3436 12926 3437
rect 12868 3431 12926 3436
rect 12868 3411 12871 3431
rect 12891 3417 12926 3431
rect 12946 3417 12955 3437
rect 12891 3409 12955 3417
rect 12917 3408 12955 3409
rect 12918 3407 12955 3408
rect 13021 3441 13057 3442
rect 13129 3441 13165 3442
rect 13021 3433 13165 3441
rect 13021 3413 13029 3433
rect 13049 3430 13137 3433
rect 13049 3413 13081 3430
rect 13101 3413 13137 3430
rect 13157 3413 13165 3433
rect 13021 3407 13165 3413
rect 13231 3437 13269 3445
rect 13337 3441 13373 3442
rect 13231 3417 13240 3437
rect 13260 3417 13269 3437
rect 13231 3408 13269 3417
rect 13288 3434 13373 3441
rect 13288 3414 13295 3434
rect 13316 3433 13373 3434
rect 13316 3414 13345 3433
rect 13288 3413 13345 3414
rect 13365 3413 13373 3433
rect 13231 3407 13268 3408
rect 13288 3407 13373 3413
rect 13439 3437 13477 3445
rect 13550 3441 13586 3442
rect 13439 3417 13448 3437
rect 13468 3417 13477 3437
rect 13439 3408 13477 3417
rect 13501 3433 13586 3441
rect 13501 3413 13558 3433
rect 13578 3413 13586 3433
rect 13439 3407 13476 3408
rect 13501 3407 13586 3413
rect 13652 3437 13690 3445
rect 13652 3417 13661 3437
rect 13681 3417 13690 3437
rect 13652 3408 13690 3417
rect 14816 3423 14856 3471
rect 15200 3491 15234 3519
rect 15426 3493 15463 3522
rect 15427 3491 15463 3493
rect 15639 3491 15676 3522
rect 15200 3490 15372 3491
rect 15200 3458 15386 3490
rect 15427 3469 15676 3491
rect 15847 3490 15884 3522
rect 16160 3518 16224 3530
rect 16264 3492 16291 3670
rect 18819 3648 18846 3826
rect 18886 3788 18950 3800
rect 19226 3796 19263 3828
rect 19434 3827 19683 3849
rect 19434 3796 19471 3827
rect 19647 3825 19683 3827
rect 19647 3796 19684 3825
rect 18886 3787 18921 3788
rect 18863 3782 18921 3787
rect 18863 3762 18866 3782
rect 18886 3768 18921 3782
rect 18941 3768 18950 3788
rect 18886 3760 18950 3768
rect 18912 3759 18950 3760
rect 18913 3758 18950 3759
rect 19016 3792 19052 3793
rect 19124 3792 19160 3793
rect 19016 3787 19160 3792
rect 19016 3784 19078 3787
rect 19016 3764 19024 3784
rect 19044 3767 19078 3784
rect 19101 3784 19160 3787
rect 19101 3767 19132 3784
rect 19044 3764 19132 3767
rect 19152 3764 19160 3784
rect 19016 3758 19160 3764
rect 19226 3788 19264 3796
rect 19332 3792 19368 3793
rect 19226 3768 19235 3788
rect 19255 3768 19264 3788
rect 19226 3759 19264 3768
rect 19283 3785 19368 3792
rect 19283 3765 19290 3785
rect 19311 3784 19368 3785
rect 19311 3765 19340 3784
rect 19283 3764 19340 3765
rect 19360 3764 19368 3784
rect 19226 3758 19263 3759
rect 19283 3758 19368 3764
rect 19434 3788 19472 3796
rect 19545 3792 19581 3793
rect 19434 3768 19443 3788
rect 19463 3768 19472 3788
rect 19434 3759 19472 3768
rect 19496 3784 19581 3792
rect 19496 3764 19553 3784
rect 19573 3764 19581 3784
rect 19434 3758 19471 3759
rect 19496 3758 19581 3764
rect 19647 3788 19685 3796
rect 19647 3768 19656 3788
rect 19676 3768 19685 3788
rect 19647 3759 19685 3768
rect 19647 3758 19684 3759
rect 19070 3737 19106 3758
rect 19496 3737 19527 3758
rect 18903 3733 19003 3737
rect 18903 3729 18965 3733
rect 18903 3703 18910 3729
rect 18936 3707 18965 3729
rect 18991 3707 19003 3733
rect 18936 3703 19003 3707
rect 18903 3700 19003 3703
rect 19071 3700 19106 3737
rect 19168 3734 19527 3737
rect 19168 3729 19390 3734
rect 19168 3705 19181 3729
rect 19205 3710 19390 3729
rect 19414 3710 19527 3734
rect 19205 3705 19527 3710
rect 19168 3701 19527 3705
rect 19594 3729 19743 3737
rect 19594 3709 19605 3729
rect 19625 3709 19743 3729
rect 19594 3702 19743 3709
rect 19594 3701 19635 3702
rect 18918 3648 18955 3649
rect 19014 3648 19051 3649
rect 19070 3648 19106 3700
rect 19125 3648 19162 3649
rect 18818 3639 18956 3648
rect 18818 3619 18927 3639
rect 18947 3619 18956 3639
rect 18818 3612 18956 3619
rect 19014 3639 19162 3648
rect 19014 3619 19023 3639
rect 19043 3619 19133 3639
rect 19153 3619 19162 3639
rect 18818 3610 18914 3612
rect 19014 3609 19162 3619
rect 19221 3639 19258 3649
rect 19333 3648 19370 3649
rect 19314 3646 19370 3648
rect 19221 3619 19229 3639
rect 19249 3619 19258 3639
rect 19070 3608 19106 3609
rect 16447 3566 16557 3580
rect 16447 3563 16490 3566
rect 16447 3558 16451 3563
rect 16123 3490 16291 3492
rect 15847 3484 16291 3490
rect 15200 3426 15234 3458
rect 13652 3407 13689 3408
rect 13075 3386 13111 3407
rect 13501 3386 13532 3407
rect 14816 3405 14827 3423
rect 14845 3405 14856 3423
rect 14816 3397 14856 3405
rect 15196 3417 15234 3426
rect 15196 3399 15206 3417
rect 15224 3399 15234 3417
rect 14817 3396 14854 3397
rect 15196 3393 15234 3399
rect 15352 3395 15386 3458
rect 15508 3463 15619 3469
rect 15508 3455 15549 3463
rect 15508 3435 15516 3455
rect 15535 3435 15549 3455
rect 15508 3433 15549 3435
rect 15577 3455 15619 3463
rect 15577 3435 15593 3455
rect 15612 3435 15619 3455
rect 15577 3433 15619 3435
rect 15508 3418 15619 3433
rect 15846 3464 16291 3484
rect 15846 3395 15884 3464
rect 16123 3463 16291 3464
rect 16369 3536 16451 3558
rect 16480 3536 16490 3563
rect 16518 3539 16525 3566
rect 16554 3558 16557 3566
rect 18552 3575 18663 3590
rect 18552 3573 18594 3575
rect 16554 3539 16619 3558
rect 16518 3536 16619 3539
rect 16369 3534 16619 3536
rect 16369 3455 16406 3534
rect 16447 3521 16557 3534
rect 16521 3465 16552 3466
rect 16369 3435 16378 3455
rect 16398 3435 16406 3455
rect 16369 3425 16406 3435
rect 16465 3455 16552 3465
rect 16465 3435 16474 3455
rect 16494 3435 16552 3455
rect 16465 3426 16552 3435
rect 16465 3425 16502 3426
rect 15196 3389 15233 3393
rect 12908 3382 13008 3386
rect 12908 3378 12970 3382
rect 12908 3352 12915 3378
rect 12941 3356 12970 3378
rect 12996 3356 13008 3382
rect 12941 3352 13008 3356
rect 12908 3349 13008 3352
rect 13076 3349 13111 3386
rect 13173 3383 13532 3386
rect 13173 3378 13395 3383
rect 13173 3354 13186 3378
rect 13210 3359 13395 3378
rect 13419 3359 13532 3383
rect 13210 3354 13532 3359
rect 13173 3350 13532 3354
rect 13599 3378 13748 3386
rect 15352 3384 15884 3395
rect 13599 3358 13610 3378
rect 13630 3358 13748 3378
rect 15351 3368 15884 3384
rect 16521 3373 16552 3426
rect 16582 3455 16619 3534
rect 16790 3544 17183 3551
rect 16790 3527 16798 3544
rect 16830 3531 17183 3544
rect 17203 3531 17206 3551
rect 18285 3546 18326 3555
rect 16830 3527 17206 3531
rect 16790 3526 17206 3527
rect 17880 3544 18048 3545
rect 18285 3544 18294 3546
rect 16790 3525 17131 3526
rect 16734 3465 16765 3466
rect 16582 3435 16591 3455
rect 16611 3435 16619 3455
rect 16582 3425 16619 3435
rect 16678 3458 16765 3465
rect 16678 3455 16739 3458
rect 16678 3435 16687 3455
rect 16707 3438 16739 3455
rect 16760 3438 16765 3458
rect 16707 3435 16765 3438
rect 16678 3428 16765 3435
rect 16790 3455 16827 3525
rect 17093 3524 17130 3525
rect 17880 3524 18294 3544
rect 18320 3524 18326 3546
rect 18552 3553 18559 3573
rect 18578 3553 18594 3573
rect 18552 3545 18594 3553
rect 18622 3573 18663 3575
rect 18622 3553 18636 3573
rect 18655 3553 18663 3573
rect 18622 3545 18663 3553
rect 18918 3549 18955 3550
rect 19221 3549 19258 3619
rect 19283 3639 19370 3646
rect 19283 3636 19341 3639
rect 19283 3616 19288 3636
rect 19309 3619 19341 3636
rect 19361 3619 19370 3639
rect 19309 3616 19370 3619
rect 19283 3609 19370 3616
rect 19429 3639 19466 3649
rect 19429 3619 19437 3639
rect 19457 3619 19466 3639
rect 19283 3608 19314 3609
rect 18917 3548 19258 3549
rect 18552 3539 18663 3545
rect 18842 3543 19258 3548
rect 17880 3518 18326 3524
rect 17880 3516 18048 3518
rect 16942 3465 16978 3466
rect 16790 3435 16799 3455
rect 16819 3435 16827 3455
rect 16678 3426 16734 3428
rect 16678 3425 16715 3426
rect 16790 3425 16827 3435
rect 16886 3455 17034 3465
rect 17134 3462 17230 3464
rect 16886 3435 16895 3455
rect 16915 3450 17005 3455
rect 16915 3435 16950 3450
rect 16886 3426 16950 3435
rect 16886 3425 16923 3426
rect 16942 3409 16950 3426
rect 16971 3435 17005 3450
rect 17025 3435 17034 3455
rect 16971 3426 17034 3435
rect 17092 3455 17230 3462
rect 17092 3435 17101 3455
rect 17121 3435 17230 3455
rect 17092 3426 17230 3435
rect 16971 3409 16978 3426
rect 16997 3425 17034 3426
rect 17093 3425 17130 3426
rect 16942 3374 16978 3409
rect 16413 3372 16454 3373
rect 15351 3367 15865 3368
rect 13599 3351 13748 3358
rect 16305 3365 16454 3372
rect 14188 3355 14702 3356
rect 13599 3350 13640 3351
rect 12923 3297 12960 3298
rect 13019 3297 13056 3298
rect 13075 3297 13111 3349
rect 13130 3297 13167 3298
rect 12823 3288 12961 3297
rect 12823 3268 12932 3288
rect 12952 3268 12961 3288
rect 12823 3261 12961 3268
rect 13019 3288 13167 3297
rect 13019 3268 13028 3288
rect 13048 3268 13138 3288
rect 13158 3268 13167 3288
rect 12823 3259 12919 3261
rect 13019 3258 13167 3268
rect 13226 3288 13263 3298
rect 13338 3297 13375 3298
rect 13319 3295 13375 3297
rect 13226 3268 13234 3288
rect 13254 3268 13263 3288
rect 13075 3257 13111 3258
rect 12005 3205 12173 3207
rect 11727 3199 12173 3205
rect 10795 3175 11211 3180
rect 11390 3178 11501 3184
rect 10795 3174 11136 3175
rect 10739 3114 10770 3115
rect 10587 3084 10596 3104
rect 10616 3084 10624 3104
rect 10587 3074 10624 3084
rect 10683 3107 10770 3114
rect 10683 3104 10744 3107
rect 10683 3084 10692 3104
rect 10712 3087 10744 3104
rect 10765 3087 10770 3107
rect 10712 3084 10770 3087
rect 10683 3077 10770 3084
rect 10795 3104 10832 3174
rect 11098 3173 11135 3174
rect 11390 3170 11431 3178
rect 11390 3150 11398 3170
rect 11417 3150 11431 3170
rect 11390 3148 11431 3150
rect 11459 3170 11501 3178
rect 11459 3150 11475 3170
rect 11494 3150 11501 3170
rect 11727 3177 11733 3199
rect 11759 3179 12173 3199
rect 12923 3198 12960 3199
rect 13226 3198 13263 3268
rect 13288 3288 13375 3295
rect 13288 3285 13346 3288
rect 13288 3265 13293 3285
rect 13314 3268 13346 3285
rect 13366 3268 13375 3288
rect 13314 3265 13375 3268
rect 13288 3258 13375 3265
rect 13434 3288 13471 3298
rect 13434 3268 13442 3288
rect 13462 3268 13471 3288
rect 13288 3257 13319 3258
rect 12922 3197 13263 3198
rect 11759 3177 11768 3179
rect 12005 3178 12173 3179
rect 12847 3192 13263 3197
rect 11727 3168 11768 3177
rect 12847 3172 12850 3192
rect 12870 3172 13263 3192
rect 13434 3189 13471 3268
rect 13501 3297 13532 3350
rect 14169 3339 14702 3355
rect 16305 3345 16423 3365
rect 16443 3345 16454 3365
rect 14169 3328 14701 3339
rect 16305 3337 16454 3345
rect 16521 3369 16880 3373
rect 16521 3364 16843 3369
rect 16521 3340 16634 3364
rect 16658 3345 16843 3364
rect 16867 3345 16880 3369
rect 16658 3340 16880 3345
rect 16521 3337 16880 3340
rect 16942 3337 16977 3374
rect 17045 3371 17145 3374
rect 17045 3367 17112 3371
rect 17045 3341 17057 3367
rect 17083 3345 17112 3367
rect 17138 3345 17145 3371
rect 17083 3341 17145 3345
rect 17045 3337 17145 3341
rect 14820 3330 14857 3334
rect 13551 3297 13588 3298
rect 13501 3288 13588 3297
rect 13501 3268 13559 3288
rect 13579 3268 13588 3288
rect 13501 3258 13588 3268
rect 13647 3288 13684 3298
rect 13647 3268 13655 3288
rect 13675 3268 13684 3288
rect 13501 3257 13532 3258
rect 13496 3189 13606 3202
rect 13647 3189 13684 3268
rect 13434 3187 13684 3189
rect 13434 3184 13535 3187
rect 13434 3165 13499 3184
rect 11459 3148 11501 3150
rect 11390 3133 11501 3148
rect 13496 3157 13499 3165
rect 13528 3157 13535 3184
rect 13563 3160 13573 3187
rect 13602 3165 13684 3187
rect 13762 3259 13930 3260
rect 14169 3259 14207 3328
rect 13762 3239 14207 3259
rect 14434 3290 14545 3305
rect 14434 3288 14476 3290
rect 14434 3268 14441 3288
rect 14460 3268 14476 3288
rect 14434 3260 14476 3268
rect 14504 3288 14545 3290
rect 14504 3268 14518 3288
rect 14537 3268 14545 3288
rect 14504 3260 14545 3268
rect 14434 3254 14545 3260
rect 14667 3265 14701 3328
rect 14819 3324 14857 3330
rect 15199 3326 15236 3327
rect 14819 3306 14829 3324
rect 14847 3306 14857 3324
rect 14819 3297 14857 3306
rect 15197 3318 15237 3326
rect 15197 3300 15208 3318
rect 15226 3300 15237 3318
rect 16521 3316 16552 3337
rect 16942 3316 16978 3337
rect 16364 3315 16401 3316
rect 14819 3265 14853 3297
rect 13762 3233 14206 3239
rect 13762 3231 13930 3233
rect 13602 3160 13606 3165
rect 13563 3157 13606 3160
rect 13496 3143 13606 3157
rect 12725 3129 12793 3138
rect 10947 3114 10983 3115
rect 10795 3084 10804 3104
rect 10824 3084 10832 3104
rect 10683 3075 10739 3077
rect 10683 3074 10720 3075
rect 10795 3074 10832 3084
rect 10891 3104 11039 3114
rect 11139 3111 11235 3113
rect 10891 3084 10900 3104
rect 10920 3084 11010 3104
rect 11030 3084 11039 3104
rect 10891 3075 11039 3084
rect 11097 3104 11235 3111
rect 11097 3084 11106 3104
rect 11126 3084 11235 3104
rect 12725 3100 12740 3129
rect 12788 3109 12793 3129
rect 12788 3100 12795 3109
rect 12725 3089 12795 3100
rect 11097 3075 11235 3084
rect 10891 3074 10928 3075
rect 10947 3023 10983 3075
rect 11002 3074 11039 3075
rect 11098 3074 11135 3075
rect 10418 3021 10459 3022
rect 10310 3014 10459 3021
rect 10310 2994 10428 3014
rect 10448 2994 10459 3014
rect 10310 2986 10459 2994
rect 10526 3018 10885 3022
rect 10526 3013 10848 3018
rect 10526 2989 10639 3013
rect 10663 2994 10848 3013
rect 10872 2994 10885 3018
rect 10663 2989 10885 2994
rect 10526 2986 10885 2989
rect 10947 2986 10982 3023
rect 11050 3020 11150 3023
rect 11050 3016 11117 3020
rect 11050 2990 11062 3016
rect 11088 2994 11117 3016
rect 11143 2994 11150 3020
rect 11088 2990 11150 2994
rect 11050 2986 11150 2990
rect 10526 2965 10557 2986
rect 10947 2965 10983 2986
rect 10369 2964 10406 2965
rect 10368 2955 10406 2964
rect 10368 2935 10377 2955
rect 10397 2935 10406 2955
rect 10368 2927 10406 2935
rect 10472 2959 10557 2965
rect 10582 2964 10619 2965
rect 10472 2939 10480 2959
rect 10500 2939 10557 2959
rect 10472 2931 10557 2939
rect 10581 2955 10619 2964
rect 10581 2935 10590 2955
rect 10610 2935 10619 2955
rect 10472 2930 10508 2931
rect 10581 2927 10619 2935
rect 10685 2959 10770 2965
rect 10790 2964 10827 2965
rect 10685 2939 10693 2959
rect 10713 2958 10770 2959
rect 10713 2939 10742 2958
rect 10685 2938 10742 2939
rect 10763 2938 10770 2958
rect 10685 2931 10770 2938
rect 10789 2955 10827 2964
rect 10789 2935 10798 2955
rect 10818 2935 10827 2955
rect 10685 2930 10721 2931
rect 10789 2927 10827 2935
rect 10893 2959 11037 2965
rect 10893 2939 10901 2959
rect 10921 2956 11009 2959
rect 10921 2939 10952 2956
rect 10893 2936 10952 2939
rect 10975 2939 11009 2956
rect 11029 2939 11037 2959
rect 10975 2936 11037 2939
rect 10893 2931 11037 2936
rect 10893 2930 10929 2931
rect 11001 2930 11037 2931
rect 11103 2964 11140 2965
rect 11103 2963 11141 2964
rect 11103 2955 11167 2963
rect 11103 2935 11112 2955
rect 11132 2941 11167 2955
rect 11187 2941 11190 2961
rect 11132 2936 11190 2941
rect 11132 2935 11167 2936
rect 10369 2898 10406 2927
rect 10370 2896 10406 2898
rect 10582 2896 10619 2927
rect 10370 2874 10619 2896
rect 10790 2895 10827 2927
rect 11103 2923 11167 2935
rect 11207 2897 11234 3075
rect 12734 2982 12795 3089
rect 13762 3053 13789 3231
rect 13829 3193 13893 3205
rect 14169 3201 14206 3233
rect 14377 3232 14626 3254
rect 14667 3233 14853 3265
rect 14681 3232 14853 3233
rect 14377 3201 14414 3232
rect 14590 3230 14626 3232
rect 14590 3201 14627 3230
rect 14819 3204 14853 3232
rect 15197 3252 15237 3300
rect 16363 3306 16401 3315
rect 16363 3286 16372 3306
rect 16392 3286 16401 3306
rect 16363 3278 16401 3286
rect 16467 3310 16552 3316
rect 16577 3315 16614 3316
rect 16467 3290 16475 3310
rect 16495 3290 16552 3310
rect 16467 3282 16552 3290
rect 16576 3306 16614 3315
rect 16576 3286 16585 3306
rect 16605 3286 16614 3306
rect 16467 3281 16503 3282
rect 16576 3278 16614 3286
rect 16680 3310 16765 3316
rect 16785 3315 16822 3316
rect 16680 3290 16688 3310
rect 16708 3309 16765 3310
rect 16708 3290 16737 3309
rect 16680 3289 16737 3290
rect 16758 3289 16765 3309
rect 16680 3282 16765 3289
rect 16784 3306 16822 3315
rect 16784 3286 16793 3306
rect 16813 3286 16822 3306
rect 16680 3281 16716 3282
rect 16784 3278 16822 3286
rect 16888 3310 17032 3316
rect 16888 3290 16896 3310
rect 16916 3290 17004 3310
rect 17024 3290 17032 3310
rect 16888 3282 17032 3290
rect 16888 3281 16924 3282
rect 16996 3281 17032 3282
rect 17098 3315 17135 3316
rect 17098 3314 17136 3315
rect 17098 3306 17162 3314
rect 17098 3286 17107 3306
rect 17127 3292 17162 3306
rect 17182 3292 17185 3312
rect 17127 3287 17185 3292
rect 17127 3286 17162 3287
rect 15508 3256 15618 3270
rect 15508 3253 15551 3256
rect 15197 3245 15322 3252
rect 15508 3248 15512 3253
rect 15197 3226 15289 3245
rect 15314 3226 15322 3245
rect 15197 3216 15322 3226
rect 15430 3226 15512 3248
rect 15541 3226 15551 3253
rect 15579 3229 15586 3256
rect 15615 3248 15618 3256
rect 16364 3249 16401 3278
rect 15615 3229 15680 3248
rect 16365 3247 16401 3249
rect 16577 3247 16614 3278
rect 16785 3251 16822 3278
rect 17098 3274 17162 3286
rect 15579 3226 15680 3229
rect 15430 3224 15680 3226
rect 13829 3192 13864 3193
rect 13806 3187 13864 3192
rect 13806 3167 13809 3187
rect 13829 3173 13864 3187
rect 13884 3173 13893 3193
rect 13829 3165 13893 3173
rect 13855 3164 13893 3165
rect 13856 3163 13893 3164
rect 13959 3197 13995 3198
rect 14067 3197 14103 3198
rect 13959 3190 14103 3197
rect 13959 3189 14019 3190
rect 13959 3169 13967 3189
rect 13987 3170 14019 3189
rect 14044 3189 14103 3190
rect 14044 3170 14075 3189
rect 13987 3169 14075 3170
rect 14095 3169 14103 3189
rect 13959 3163 14103 3169
rect 14169 3193 14207 3201
rect 14275 3197 14311 3198
rect 14169 3173 14178 3193
rect 14198 3173 14207 3193
rect 14169 3164 14207 3173
rect 14226 3190 14311 3197
rect 14226 3170 14233 3190
rect 14254 3189 14311 3190
rect 14254 3170 14283 3189
rect 14226 3169 14283 3170
rect 14303 3169 14311 3189
rect 14169 3163 14206 3164
rect 14226 3163 14311 3169
rect 14377 3193 14415 3201
rect 14488 3197 14524 3198
rect 14377 3173 14386 3193
rect 14406 3173 14415 3193
rect 14377 3164 14415 3173
rect 14439 3189 14524 3197
rect 14439 3169 14496 3189
rect 14516 3169 14524 3189
rect 14377 3163 14414 3164
rect 14439 3163 14524 3169
rect 14590 3193 14628 3201
rect 14590 3173 14599 3193
rect 14619 3173 14628 3193
rect 14590 3164 14628 3173
rect 14817 3194 14854 3204
rect 15197 3196 15237 3216
rect 14817 3176 14827 3194
rect 14845 3176 14854 3194
rect 14817 3167 14854 3176
rect 15196 3187 15237 3196
rect 15196 3169 15206 3187
rect 15224 3169 15237 3187
rect 14819 3166 14853 3167
rect 14590 3163 14627 3164
rect 14013 3142 14049 3163
rect 14439 3142 14470 3163
rect 15196 3160 15237 3169
rect 15196 3159 15233 3160
rect 15430 3145 15467 3224
rect 15508 3211 15618 3224
rect 15582 3155 15613 3156
rect 13846 3138 13946 3142
rect 13846 3134 13908 3138
rect 13846 3108 13853 3134
rect 13879 3112 13908 3134
rect 13934 3112 13946 3138
rect 13879 3108 13946 3112
rect 13846 3105 13946 3108
rect 14014 3105 14049 3142
rect 14111 3139 14470 3142
rect 14111 3134 14333 3139
rect 14111 3110 14124 3134
rect 14148 3115 14333 3134
rect 14357 3115 14470 3139
rect 14148 3110 14470 3115
rect 14111 3106 14470 3110
rect 14537 3134 14686 3142
rect 14537 3114 14548 3134
rect 14568 3114 14686 3134
rect 15430 3125 15439 3145
rect 15459 3125 15467 3145
rect 15430 3115 15467 3125
rect 15526 3145 15613 3155
rect 15526 3125 15535 3145
rect 15555 3125 15613 3145
rect 15526 3116 15613 3125
rect 15526 3115 15563 3116
rect 14537 3107 14686 3114
rect 14537 3106 14578 3107
rect 13861 3053 13898 3054
rect 13957 3053 13994 3054
rect 14013 3053 14049 3105
rect 14068 3053 14105 3054
rect 13761 3044 13899 3053
rect 12725 2981 12795 2982
rect 13386 3010 13497 3025
rect 13761 3024 13870 3044
rect 13890 3024 13899 3044
rect 13761 3017 13899 3024
rect 13957 3044 14105 3053
rect 13957 3024 13966 3044
rect 13986 3024 14076 3044
rect 14096 3024 14105 3044
rect 13761 3015 13857 3017
rect 13957 3014 14105 3024
rect 14164 3044 14201 3054
rect 14276 3053 14313 3054
rect 14257 3051 14313 3053
rect 14164 3024 14172 3044
rect 14192 3024 14201 3044
rect 14013 3013 14049 3014
rect 13386 3008 13428 3010
rect 13386 2988 13393 3008
rect 13412 2988 13428 3008
rect 12725 2980 12833 2981
rect 13386 2980 13428 2988
rect 13456 3008 13497 3010
rect 13456 2988 13470 3008
rect 13489 2988 13497 3008
rect 13456 2980 13497 2988
rect 12714 2979 12882 2980
rect 11501 2946 11611 2960
rect 11501 2943 11544 2946
rect 11501 2938 11505 2943
rect 11066 2895 11234 2897
rect 10790 2892 11234 2895
rect 10451 2868 10562 2874
rect 10451 2860 10492 2868
rect 10140 2805 10179 2849
rect 10451 2840 10459 2860
rect 10478 2840 10492 2860
rect 10451 2838 10492 2840
rect 10520 2860 10562 2868
rect 10520 2840 10536 2860
rect 10555 2840 10562 2860
rect 10520 2838 10562 2840
rect 10451 2824 10562 2838
rect 10788 2869 11234 2892
rect 10140 2781 10180 2805
rect 10480 2781 10527 2783
rect 10788 2781 10826 2869
rect 11066 2868 11234 2869
rect 11423 2916 11505 2938
rect 11534 2916 11544 2943
rect 11572 2919 11579 2946
rect 11608 2938 11611 2946
rect 12714 2953 13158 2979
rect 13386 2974 13497 2980
rect 12714 2951 12882 2953
rect 12714 2949 12833 2951
rect 11608 2919 11673 2938
rect 11572 2916 11673 2919
rect 11423 2914 11673 2916
rect 11423 2835 11460 2914
rect 11501 2901 11611 2914
rect 11575 2845 11606 2846
rect 11423 2815 11432 2835
rect 11452 2815 11460 2835
rect 11423 2805 11460 2815
rect 11519 2835 11606 2845
rect 11519 2815 11528 2835
rect 11548 2815 11606 2835
rect 11519 2806 11606 2815
rect 11519 2805 11556 2806
rect 10140 2748 10826 2781
rect 11575 2753 11606 2806
rect 11636 2835 11673 2914
rect 11844 2933 11876 2945
rect 11844 2913 11846 2933
rect 11867 2931 11876 2933
rect 11867 2929 12219 2931
rect 11867 2913 12237 2929
rect 11844 2911 12237 2913
rect 12257 2911 12260 2929
rect 11844 2906 12260 2911
rect 11844 2905 12185 2906
rect 11788 2845 11819 2846
rect 11636 2815 11645 2835
rect 11665 2815 11673 2835
rect 11636 2805 11673 2815
rect 11732 2838 11819 2845
rect 11732 2835 11793 2838
rect 11732 2815 11741 2835
rect 11761 2818 11793 2835
rect 11814 2818 11819 2838
rect 11761 2815 11819 2818
rect 11732 2808 11819 2815
rect 11844 2835 11881 2905
rect 12147 2904 12184 2905
rect 11996 2845 12032 2846
rect 11844 2815 11853 2835
rect 11873 2815 11881 2835
rect 11732 2806 11788 2808
rect 11732 2805 11769 2806
rect 11844 2805 11881 2815
rect 11940 2835 12088 2845
rect 12188 2842 12284 2844
rect 11940 2815 11949 2835
rect 11969 2826 12059 2835
rect 11969 2815 12000 2826
rect 11940 2806 12000 2815
rect 11940 2805 11977 2806
rect 11996 2794 12000 2806
rect 12027 2815 12059 2826
rect 12079 2815 12088 2835
rect 12027 2806 12088 2815
rect 12146 2835 12284 2842
rect 12146 2815 12155 2835
rect 12175 2815 12284 2835
rect 12146 2806 12284 2815
rect 12027 2794 12032 2806
rect 12051 2805 12088 2806
rect 12147 2805 12184 2806
rect 11996 2754 12032 2794
rect 11467 2752 11508 2753
rect 10139 2691 10178 2748
rect 10788 2746 10826 2748
rect 11359 2745 11508 2752
rect 11359 2725 11477 2745
rect 11497 2725 11508 2745
rect 11359 2717 11508 2725
rect 11575 2749 11934 2753
rect 11575 2744 11897 2749
rect 11575 2720 11688 2744
rect 11712 2725 11897 2744
rect 11921 2725 11934 2749
rect 11712 2720 11934 2725
rect 11575 2717 11934 2720
rect 11996 2717 12031 2754
rect 12099 2751 12199 2754
rect 12099 2747 12166 2751
rect 12099 2721 12111 2747
rect 12137 2725 12166 2747
rect 12192 2725 12199 2751
rect 12137 2721 12199 2725
rect 12099 2717 12199 2721
rect 11575 2696 11606 2717
rect 11996 2696 12032 2717
rect 11418 2695 11455 2696
rect 10139 2689 10187 2691
rect 10139 2671 10150 2689
rect 10168 2671 10187 2689
rect 11417 2686 11455 2695
rect 10139 2662 10187 2671
rect 10140 2661 10187 2662
rect 10453 2666 10563 2680
rect 10453 2663 10496 2666
rect 10453 2658 10457 2663
rect 10375 2636 10457 2658
rect 10486 2636 10496 2663
rect 10524 2639 10531 2666
rect 10560 2658 10563 2666
rect 11417 2666 11426 2686
rect 11446 2666 11455 2686
rect 11417 2658 11455 2666
rect 11521 2690 11606 2696
rect 11631 2695 11668 2696
rect 11521 2670 11529 2690
rect 11549 2670 11606 2690
rect 11521 2662 11606 2670
rect 11630 2686 11668 2695
rect 11630 2666 11639 2686
rect 11659 2666 11668 2686
rect 11521 2661 11557 2662
rect 11630 2658 11668 2666
rect 11734 2690 11819 2696
rect 11839 2695 11876 2696
rect 11734 2670 11742 2690
rect 11762 2689 11819 2690
rect 11762 2670 11791 2689
rect 11734 2669 11791 2670
rect 11812 2669 11819 2689
rect 11734 2662 11819 2669
rect 11838 2686 11876 2695
rect 11838 2666 11847 2686
rect 11867 2666 11876 2686
rect 11734 2661 11770 2662
rect 11838 2658 11876 2666
rect 11942 2690 12086 2696
rect 11942 2670 11950 2690
rect 11970 2670 12058 2690
rect 12078 2670 12086 2690
rect 11942 2662 12086 2670
rect 11942 2661 11978 2662
rect 12050 2661 12086 2662
rect 12152 2695 12189 2696
rect 12152 2694 12190 2695
rect 12152 2686 12216 2694
rect 12152 2666 12161 2686
rect 12181 2672 12216 2686
rect 12236 2672 12239 2692
rect 12181 2667 12239 2672
rect 12181 2666 12216 2667
rect 10560 2639 10625 2658
rect 10524 2636 10625 2639
rect 10375 2634 10625 2636
rect 10143 2598 10180 2599
rect 9842 2568 9852 2586
rect 9870 2568 9882 2586
rect 9842 2563 9882 2568
rect 10139 2595 10180 2598
rect 10139 2590 10181 2595
rect 10139 2572 10152 2590
rect 10170 2572 10181 2590
rect 9842 2559 9879 2563
rect 10139 2558 10181 2572
rect 10219 2558 10266 2562
rect 10139 2552 10266 2558
rect 9515 2540 9552 2541
rect 9465 2531 9552 2540
rect 9465 2511 9523 2531
rect 9543 2511 9552 2531
rect 9465 2501 9552 2511
rect 9611 2531 9648 2541
rect 9611 2511 9619 2531
rect 9639 2511 9648 2531
rect 9465 2500 9496 2501
rect 9460 2432 9570 2445
rect 9611 2432 9648 2511
rect 10139 2523 10227 2552
rect 10256 2523 10266 2552
rect 10375 2555 10412 2634
rect 10453 2621 10563 2634
rect 10527 2565 10558 2566
rect 10375 2535 10384 2555
rect 10404 2535 10412 2555
rect 10375 2525 10412 2535
rect 10471 2555 10558 2565
rect 10471 2535 10480 2555
rect 10500 2535 10558 2555
rect 10471 2526 10558 2535
rect 10471 2525 10508 2526
rect 10139 2519 10266 2523
rect 10139 2502 10178 2519
rect 10219 2518 10266 2519
rect 9845 2496 9882 2497
rect 9841 2487 9882 2496
rect 9841 2469 9854 2487
rect 9872 2469 9882 2487
rect 10139 2484 10150 2502
rect 10168 2484 10178 2502
rect 10139 2475 10178 2484
rect 10140 2474 10177 2475
rect 10527 2473 10558 2526
rect 10588 2555 10625 2634
rect 10796 2631 11189 2651
rect 11209 2631 11212 2651
rect 10796 2626 11212 2631
rect 11418 2629 11455 2658
rect 11419 2627 11455 2629
rect 11631 2627 11668 2658
rect 10796 2625 11137 2626
rect 10740 2565 10771 2566
rect 10588 2535 10597 2555
rect 10617 2535 10625 2555
rect 10588 2525 10625 2535
rect 10684 2558 10771 2565
rect 10684 2555 10745 2558
rect 10684 2535 10693 2555
rect 10713 2538 10745 2555
rect 10766 2538 10771 2558
rect 10713 2535 10771 2538
rect 10684 2528 10771 2535
rect 10796 2555 10833 2625
rect 11099 2624 11136 2625
rect 11419 2605 11668 2627
rect 11839 2626 11876 2658
rect 12152 2654 12216 2666
rect 12256 2636 12283 2806
rect 12714 2773 12741 2949
rect 12781 2913 12845 2925
rect 13121 2921 13158 2953
rect 13329 2952 13578 2974
rect 13861 2954 13898 2955
rect 14164 2954 14201 3024
rect 14226 3044 14313 3051
rect 14226 3041 14284 3044
rect 14226 3021 14231 3041
rect 14252 3024 14284 3041
rect 14304 3024 14313 3044
rect 14252 3021 14313 3024
rect 14226 3014 14313 3021
rect 14372 3044 14409 3054
rect 14372 3024 14380 3044
rect 14400 3024 14409 3044
rect 14226 3013 14257 3014
rect 13860 2953 14201 2954
rect 13329 2921 13366 2952
rect 13542 2950 13578 2952
rect 13542 2921 13579 2950
rect 13785 2948 14201 2953
rect 13785 2928 13788 2948
rect 13808 2928 14201 2948
rect 14372 2945 14409 3024
rect 14439 3053 14470 3106
rect 14820 3104 14857 3105
rect 14819 3095 14858 3104
rect 14819 3077 14829 3095
rect 14847 3077 14858 3095
rect 15199 3093 15236 3097
rect 14731 3060 14778 3061
rect 14819 3060 14858 3077
rect 14731 3056 14858 3060
rect 14489 3053 14526 3054
rect 14439 3044 14526 3053
rect 14439 3024 14497 3044
rect 14517 3024 14526 3044
rect 14439 3014 14526 3024
rect 14585 3044 14622 3054
rect 14585 3024 14593 3044
rect 14613 3024 14622 3044
rect 14439 3013 14470 3014
rect 14434 2945 14544 2958
rect 14585 2945 14622 3024
rect 14731 3027 14741 3056
rect 14770 3027 14858 3056
rect 14731 3021 14858 3027
rect 14731 3017 14778 3021
rect 14816 3007 14858 3021
rect 14816 2989 14827 3007
rect 14845 2989 14858 3007
rect 14816 2984 14858 2989
rect 14817 2981 14858 2984
rect 15196 3088 15236 3093
rect 15196 3070 15208 3088
rect 15226 3070 15236 3088
rect 14817 2980 14854 2981
rect 14372 2943 14622 2945
rect 14372 2940 14473 2943
rect 14372 2921 14437 2940
rect 12781 2912 12816 2913
rect 12758 2907 12816 2912
rect 12758 2887 12761 2907
rect 12781 2893 12816 2907
rect 12836 2893 12845 2913
rect 12781 2885 12845 2893
rect 12807 2884 12845 2885
rect 12808 2883 12845 2884
rect 12911 2917 12947 2918
rect 13019 2917 13055 2918
rect 12911 2910 13055 2917
rect 12911 2909 12969 2910
rect 12911 2889 12919 2909
rect 12939 2891 12969 2909
rect 12998 2909 13055 2910
rect 12998 2891 13027 2909
rect 12939 2889 13027 2891
rect 13047 2889 13055 2909
rect 12911 2883 13055 2889
rect 13121 2913 13159 2921
rect 13227 2917 13263 2918
rect 13121 2893 13130 2913
rect 13150 2893 13159 2913
rect 13121 2884 13159 2893
rect 13178 2910 13263 2917
rect 13178 2890 13185 2910
rect 13206 2909 13263 2910
rect 13206 2890 13235 2909
rect 13178 2889 13235 2890
rect 13255 2889 13263 2909
rect 13121 2883 13158 2884
rect 13178 2883 13263 2889
rect 13329 2913 13367 2921
rect 13440 2917 13476 2918
rect 13329 2893 13338 2913
rect 13358 2893 13367 2913
rect 13329 2884 13367 2893
rect 13391 2909 13476 2917
rect 13391 2889 13448 2909
rect 13468 2889 13476 2909
rect 13329 2883 13366 2884
rect 13391 2883 13476 2889
rect 13542 2913 13580 2921
rect 13542 2893 13551 2913
rect 13571 2893 13580 2913
rect 14434 2913 14437 2921
rect 14466 2913 14473 2940
rect 14501 2916 14511 2943
rect 14540 2921 14622 2943
rect 14540 2916 14544 2921
rect 14501 2913 14544 2916
rect 14434 2899 14544 2913
rect 14810 2917 14857 2918
rect 14810 2908 14858 2917
rect 13542 2884 13580 2893
rect 14810 2890 14829 2908
rect 14847 2890 14858 2908
rect 14810 2888 14858 2890
rect 13542 2883 13579 2884
rect 12965 2862 13001 2883
rect 13391 2862 13422 2883
rect 12798 2858 12898 2862
rect 12798 2854 12860 2858
rect 12798 2828 12805 2854
rect 12831 2832 12860 2854
rect 12886 2832 12898 2858
rect 12831 2828 12898 2832
rect 12798 2825 12898 2828
rect 12966 2825 13001 2862
rect 13063 2859 13422 2862
rect 13063 2854 13285 2859
rect 13063 2830 13076 2854
rect 13100 2835 13285 2854
rect 13309 2835 13422 2859
rect 13100 2830 13422 2835
rect 13063 2826 13422 2830
rect 13489 2854 13638 2862
rect 13489 2834 13500 2854
rect 13520 2834 13638 2854
rect 13489 2827 13638 2834
rect 14171 2831 14209 2833
rect 14819 2831 14858 2888
rect 15196 2890 15236 3070
rect 15582 3063 15613 3116
rect 15643 3145 15680 3224
rect 15851 3221 16244 3241
rect 16264 3221 16267 3241
rect 16365 3225 16614 3247
rect 16783 3246 16824 3251
rect 17202 3248 17229 3426
rect 17880 3338 17907 3516
rect 18285 3513 18326 3518
rect 18495 3517 18744 3539
rect 18842 3523 18845 3543
rect 18865 3523 19258 3543
rect 19429 3540 19466 3619
rect 19496 3648 19527 3701
rect 19873 3694 19913 3874
rect 19873 3676 19883 3694
rect 19901 3676 19913 3694
rect 19873 3671 19913 3676
rect 19873 3667 19910 3671
rect 19546 3648 19583 3649
rect 19496 3639 19583 3648
rect 19496 3619 19554 3639
rect 19574 3619 19583 3639
rect 19496 3609 19583 3619
rect 19642 3639 19679 3649
rect 19642 3619 19650 3639
rect 19670 3619 19679 3639
rect 19496 3608 19527 3609
rect 19491 3540 19601 3553
rect 19642 3540 19679 3619
rect 19876 3604 19913 3605
rect 19872 3595 19913 3604
rect 19872 3577 19885 3595
rect 19903 3577 19913 3595
rect 19872 3568 19913 3577
rect 19872 3548 19912 3568
rect 19429 3538 19679 3540
rect 19429 3535 19530 3538
rect 17947 3478 18011 3490
rect 18287 3486 18324 3513
rect 18495 3486 18532 3517
rect 18708 3515 18744 3517
rect 19429 3516 19494 3535
rect 18708 3486 18745 3515
rect 19491 3508 19494 3516
rect 19523 3508 19530 3535
rect 19558 3511 19568 3538
rect 19597 3516 19679 3538
rect 19787 3538 19912 3548
rect 19787 3519 19795 3538
rect 19820 3519 19912 3538
rect 19597 3511 19601 3516
rect 19787 3512 19912 3519
rect 19558 3508 19601 3511
rect 19491 3494 19601 3508
rect 17947 3477 17982 3478
rect 17924 3472 17982 3477
rect 17924 3452 17927 3472
rect 17947 3458 17982 3472
rect 18002 3458 18011 3478
rect 17947 3450 18011 3458
rect 17973 3449 18011 3450
rect 17974 3448 18011 3449
rect 18077 3482 18113 3483
rect 18185 3482 18221 3483
rect 18077 3474 18221 3482
rect 18077 3454 18085 3474
rect 18105 3471 18193 3474
rect 18105 3454 18137 3471
rect 18157 3454 18193 3471
rect 18213 3454 18221 3474
rect 18077 3448 18221 3454
rect 18287 3478 18325 3486
rect 18393 3482 18429 3483
rect 18287 3458 18296 3478
rect 18316 3458 18325 3478
rect 18287 3449 18325 3458
rect 18344 3475 18429 3482
rect 18344 3455 18351 3475
rect 18372 3474 18429 3475
rect 18372 3455 18401 3474
rect 18344 3454 18401 3455
rect 18421 3454 18429 3474
rect 18287 3448 18324 3449
rect 18344 3448 18429 3454
rect 18495 3478 18533 3486
rect 18606 3482 18642 3483
rect 18495 3458 18504 3478
rect 18524 3458 18533 3478
rect 18495 3449 18533 3458
rect 18557 3474 18642 3482
rect 18557 3454 18614 3474
rect 18634 3454 18642 3474
rect 18495 3448 18532 3449
rect 18557 3448 18642 3454
rect 18708 3478 18746 3486
rect 18708 3458 18717 3478
rect 18737 3458 18746 3478
rect 18708 3449 18746 3458
rect 19872 3464 19912 3512
rect 18708 3448 18745 3449
rect 18131 3427 18167 3448
rect 18557 3427 18588 3448
rect 19872 3446 19883 3464
rect 19901 3446 19912 3464
rect 19872 3438 19912 3446
rect 19873 3437 19910 3438
rect 17964 3423 18064 3427
rect 17964 3419 18026 3423
rect 17964 3393 17971 3419
rect 17997 3397 18026 3419
rect 18052 3397 18064 3423
rect 17997 3393 18064 3397
rect 17964 3390 18064 3393
rect 18132 3390 18167 3427
rect 18229 3424 18588 3427
rect 18229 3419 18451 3424
rect 18229 3395 18242 3419
rect 18266 3400 18451 3419
rect 18475 3400 18588 3424
rect 18266 3395 18588 3400
rect 18229 3391 18588 3395
rect 18655 3419 18804 3427
rect 18655 3399 18666 3419
rect 18686 3399 18804 3419
rect 18655 3392 18804 3399
rect 19244 3396 19758 3397
rect 18655 3391 18696 3392
rect 17979 3338 18016 3339
rect 18075 3338 18112 3339
rect 18131 3338 18167 3390
rect 18186 3338 18223 3339
rect 17879 3329 18017 3338
rect 17879 3309 17988 3329
rect 18008 3309 18017 3329
rect 17879 3302 18017 3309
rect 18075 3329 18223 3338
rect 18075 3309 18084 3329
rect 18104 3309 18194 3329
rect 18214 3309 18223 3329
rect 17879 3300 17975 3302
rect 18075 3299 18223 3309
rect 18282 3329 18319 3339
rect 18394 3338 18431 3339
rect 18375 3336 18431 3338
rect 18282 3309 18290 3329
rect 18310 3309 18319 3329
rect 18131 3298 18167 3299
rect 17061 3246 17229 3248
rect 16783 3240 17229 3246
rect 15851 3216 16267 3221
rect 16446 3219 16557 3225
rect 15851 3215 16192 3216
rect 15795 3155 15826 3156
rect 15643 3125 15652 3145
rect 15672 3125 15680 3145
rect 15643 3115 15680 3125
rect 15739 3148 15826 3155
rect 15739 3145 15800 3148
rect 15739 3125 15748 3145
rect 15768 3128 15800 3145
rect 15821 3128 15826 3148
rect 15768 3125 15826 3128
rect 15739 3118 15826 3125
rect 15851 3145 15888 3215
rect 16154 3214 16191 3215
rect 16446 3211 16487 3219
rect 16446 3191 16454 3211
rect 16473 3191 16487 3211
rect 16446 3189 16487 3191
rect 16515 3211 16557 3219
rect 16515 3191 16531 3211
rect 16550 3191 16557 3211
rect 16783 3218 16789 3240
rect 16815 3220 17229 3240
rect 17979 3239 18016 3240
rect 18282 3239 18319 3309
rect 18344 3329 18431 3336
rect 18344 3326 18402 3329
rect 18344 3306 18349 3326
rect 18370 3309 18402 3326
rect 18422 3309 18431 3329
rect 18370 3306 18431 3309
rect 18344 3299 18431 3306
rect 18490 3329 18527 3339
rect 18490 3309 18498 3329
rect 18518 3309 18527 3329
rect 18344 3298 18375 3299
rect 17978 3238 18319 3239
rect 16815 3218 16824 3220
rect 17061 3219 17229 3220
rect 17903 3233 18319 3238
rect 16783 3209 16824 3218
rect 17903 3213 17906 3233
rect 17926 3213 18319 3233
rect 18490 3230 18527 3309
rect 18557 3338 18588 3391
rect 19225 3380 19758 3396
rect 19225 3369 19757 3380
rect 19876 3371 19913 3375
rect 18607 3338 18644 3339
rect 18557 3329 18644 3338
rect 18557 3309 18615 3329
rect 18635 3309 18644 3329
rect 18557 3299 18644 3309
rect 18703 3329 18740 3339
rect 18703 3309 18711 3329
rect 18731 3309 18740 3329
rect 18557 3298 18588 3299
rect 18552 3230 18662 3243
rect 18703 3230 18740 3309
rect 18490 3228 18740 3230
rect 18490 3225 18591 3228
rect 18490 3206 18555 3225
rect 16515 3189 16557 3191
rect 16446 3174 16557 3189
rect 18552 3198 18555 3206
rect 18584 3198 18591 3225
rect 18619 3201 18629 3228
rect 18658 3206 18740 3228
rect 18818 3300 18986 3301
rect 19225 3300 19263 3369
rect 18818 3280 19263 3300
rect 19490 3331 19601 3346
rect 19490 3329 19532 3331
rect 19490 3309 19497 3329
rect 19516 3309 19532 3329
rect 19490 3301 19532 3309
rect 19560 3329 19601 3331
rect 19560 3309 19574 3329
rect 19593 3309 19601 3329
rect 19560 3301 19601 3309
rect 19490 3295 19601 3301
rect 19723 3306 19757 3369
rect 19875 3365 19913 3371
rect 19875 3347 19885 3365
rect 19903 3347 19913 3365
rect 19875 3338 19913 3347
rect 19875 3306 19909 3338
rect 18818 3274 19262 3280
rect 18818 3272 18986 3274
rect 18658 3201 18662 3206
rect 18619 3198 18662 3201
rect 18552 3184 18662 3198
rect 17781 3170 17849 3179
rect 16003 3155 16039 3156
rect 15851 3125 15860 3145
rect 15880 3125 15888 3145
rect 15739 3116 15795 3118
rect 15739 3115 15776 3116
rect 15851 3115 15888 3125
rect 15947 3145 16095 3155
rect 16195 3152 16291 3154
rect 15947 3125 15956 3145
rect 15976 3125 16066 3145
rect 16086 3125 16095 3145
rect 15947 3116 16095 3125
rect 16153 3145 16291 3152
rect 16153 3125 16162 3145
rect 16182 3125 16291 3145
rect 17781 3141 17796 3170
rect 17844 3150 17849 3170
rect 17844 3141 17851 3150
rect 17781 3130 17851 3141
rect 16153 3116 16291 3125
rect 15947 3115 15984 3116
rect 16003 3064 16039 3116
rect 16058 3115 16095 3116
rect 16154 3115 16191 3116
rect 15474 3062 15515 3063
rect 15366 3055 15515 3062
rect 15366 3035 15484 3055
rect 15504 3035 15515 3055
rect 15366 3027 15515 3035
rect 15582 3059 15941 3063
rect 15582 3054 15904 3059
rect 15582 3030 15695 3054
rect 15719 3035 15904 3054
rect 15928 3035 15941 3059
rect 15719 3030 15941 3035
rect 15582 3027 15941 3030
rect 16003 3027 16038 3064
rect 16106 3061 16206 3064
rect 16106 3057 16173 3061
rect 16106 3031 16118 3057
rect 16144 3035 16173 3057
rect 16199 3035 16206 3061
rect 16144 3031 16206 3035
rect 16106 3027 16206 3031
rect 15582 3006 15613 3027
rect 16003 3006 16039 3027
rect 15425 3005 15462 3006
rect 15424 2996 15462 3005
rect 15424 2976 15433 2996
rect 15453 2976 15462 2996
rect 15424 2968 15462 2976
rect 15528 3000 15613 3006
rect 15638 3005 15675 3006
rect 15528 2980 15536 3000
rect 15556 2980 15613 3000
rect 15528 2972 15613 2980
rect 15637 2996 15675 3005
rect 15637 2976 15646 2996
rect 15666 2976 15675 2996
rect 15528 2971 15564 2972
rect 15637 2968 15675 2976
rect 15741 3000 15826 3006
rect 15846 3005 15883 3006
rect 15741 2980 15749 3000
rect 15769 2999 15826 3000
rect 15769 2980 15798 2999
rect 15741 2979 15798 2980
rect 15819 2979 15826 2999
rect 15741 2972 15826 2979
rect 15845 2996 15883 3005
rect 15845 2976 15854 2996
rect 15874 2976 15883 2996
rect 15741 2971 15777 2972
rect 15845 2968 15883 2976
rect 15949 3000 16093 3006
rect 15949 2980 15957 3000
rect 15977 2997 16065 3000
rect 15977 2980 16008 2997
rect 15949 2977 16008 2980
rect 16031 2980 16065 2997
rect 16085 2980 16093 3000
rect 16031 2977 16093 2980
rect 15949 2972 16093 2977
rect 15949 2971 15985 2972
rect 16057 2971 16093 2972
rect 16159 3005 16196 3006
rect 16159 3004 16197 3005
rect 16159 2996 16223 3004
rect 16159 2976 16168 2996
rect 16188 2982 16223 2996
rect 16243 2982 16246 3002
rect 16188 2977 16246 2982
rect 16188 2976 16223 2977
rect 15425 2939 15462 2968
rect 15426 2937 15462 2939
rect 15638 2937 15675 2968
rect 15426 2915 15675 2937
rect 15846 2936 15883 2968
rect 16159 2964 16223 2976
rect 16263 2938 16290 3116
rect 17790 3023 17851 3130
rect 18818 3094 18845 3272
rect 18885 3234 18949 3246
rect 19225 3242 19262 3274
rect 19433 3273 19682 3295
rect 19723 3274 19909 3306
rect 19737 3273 19909 3274
rect 19433 3242 19470 3273
rect 19646 3271 19682 3273
rect 19646 3242 19683 3271
rect 19875 3245 19909 3273
rect 18885 3233 18920 3234
rect 18862 3228 18920 3233
rect 18862 3208 18865 3228
rect 18885 3214 18920 3228
rect 18940 3214 18949 3234
rect 18885 3206 18949 3214
rect 18911 3205 18949 3206
rect 18912 3204 18949 3205
rect 19015 3238 19051 3239
rect 19123 3238 19159 3239
rect 19015 3231 19159 3238
rect 19015 3230 19075 3231
rect 19015 3210 19023 3230
rect 19043 3211 19075 3230
rect 19100 3230 19159 3231
rect 19100 3211 19131 3230
rect 19043 3210 19131 3211
rect 19151 3210 19159 3230
rect 19015 3204 19159 3210
rect 19225 3234 19263 3242
rect 19331 3238 19367 3239
rect 19225 3214 19234 3234
rect 19254 3214 19263 3234
rect 19225 3205 19263 3214
rect 19282 3231 19367 3238
rect 19282 3211 19289 3231
rect 19310 3230 19367 3231
rect 19310 3211 19339 3230
rect 19282 3210 19339 3211
rect 19359 3210 19367 3230
rect 19225 3204 19262 3205
rect 19282 3204 19367 3210
rect 19433 3234 19471 3242
rect 19544 3238 19580 3239
rect 19433 3214 19442 3234
rect 19462 3214 19471 3234
rect 19433 3205 19471 3214
rect 19495 3230 19580 3238
rect 19495 3210 19552 3230
rect 19572 3210 19580 3230
rect 19433 3204 19470 3205
rect 19495 3204 19580 3210
rect 19646 3234 19684 3242
rect 19646 3214 19655 3234
rect 19675 3214 19684 3234
rect 19646 3205 19684 3214
rect 19873 3235 19910 3245
rect 19873 3217 19883 3235
rect 19901 3217 19910 3235
rect 19873 3208 19910 3217
rect 19875 3207 19909 3208
rect 19646 3204 19683 3205
rect 19069 3183 19105 3204
rect 19495 3183 19526 3204
rect 18902 3179 19002 3183
rect 18902 3175 18964 3179
rect 18902 3149 18909 3175
rect 18935 3153 18964 3175
rect 18990 3153 19002 3179
rect 18935 3149 19002 3153
rect 18902 3146 19002 3149
rect 19070 3146 19105 3183
rect 19167 3180 19526 3183
rect 19167 3175 19389 3180
rect 19167 3151 19180 3175
rect 19204 3156 19389 3175
rect 19413 3156 19526 3180
rect 19204 3151 19526 3156
rect 19167 3147 19526 3151
rect 19593 3175 19742 3183
rect 19593 3155 19604 3175
rect 19624 3155 19742 3175
rect 19593 3148 19742 3155
rect 19593 3147 19634 3148
rect 18917 3094 18954 3095
rect 19013 3094 19050 3095
rect 19069 3094 19105 3146
rect 19124 3094 19161 3095
rect 18817 3085 18955 3094
rect 17781 3022 17851 3023
rect 18442 3051 18553 3066
rect 18817 3065 18926 3085
rect 18946 3065 18955 3085
rect 18817 3058 18955 3065
rect 19013 3085 19161 3094
rect 19013 3065 19022 3085
rect 19042 3065 19132 3085
rect 19152 3065 19161 3085
rect 18817 3056 18913 3058
rect 19013 3055 19161 3065
rect 19220 3085 19257 3095
rect 19332 3094 19369 3095
rect 19313 3092 19369 3094
rect 19220 3065 19228 3085
rect 19248 3065 19257 3085
rect 19069 3054 19105 3055
rect 18442 3049 18484 3051
rect 18442 3029 18449 3049
rect 18468 3029 18484 3049
rect 17781 3021 17889 3022
rect 18442 3021 18484 3029
rect 18512 3049 18553 3051
rect 18512 3029 18526 3049
rect 18545 3029 18553 3049
rect 18512 3021 18553 3029
rect 17770 3020 17938 3021
rect 16557 2987 16667 3001
rect 16557 2984 16600 2987
rect 16557 2979 16561 2984
rect 16122 2936 16290 2938
rect 15846 2933 16290 2936
rect 15507 2909 15618 2915
rect 15507 2901 15548 2909
rect 15196 2846 15235 2890
rect 15507 2881 15515 2901
rect 15534 2881 15548 2901
rect 15507 2879 15548 2881
rect 15576 2901 15618 2909
rect 15576 2881 15592 2901
rect 15611 2881 15618 2901
rect 15576 2879 15618 2881
rect 15507 2865 15618 2879
rect 15844 2910 16290 2933
rect 13489 2826 13530 2827
rect 12813 2773 12850 2774
rect 12909 2773 12946 2774
rect 12965 2773 13001 2825
rect 13020 2773 13057 2774
rect 12713 2764 12851 2773
rect 12713 2744 12822 2764
rect 12842 2744 12851 2764
rect 12713 2737 12851 2744
rect 12909 2764 13057 2773
rect 12909 2744 12918 2764
rect 12938 2744 13028 2764
rect 13048 2744 13057 2764
rect 12713 2735 12809 2737
rect 12909 2734 13057 2744
rect 13116 2764 13153 2774
rect 13228 2773 13265 2774
rect 13209 2771 13265 2773
rect 13116 2744 13124 2764
rect 13144 2744 13153 2764
rect 12965 2733 13001 2734
rect 12813 2674 12850 2675
rect 13116 2674 13153 2744
rect 13178 2764 13265 2771
rect 13178 2761 13236 2764
rect 13178 2741 13183 2761
rect 13204 2744 13236 2761
rect 13256 2744 13265 2764
rect 13204 2741 13265 2744
rect 13178 2734 13265 2741
rect 13324 2764 13361 2774
rect 13324 2744 13332 2764
rect 13352 2744 13361 2764
rect 13178 2733 13209 2734
rect 12812 2673 13153 2674
rect 12737 2668 13153 2673
rect 12737 2648 12740 2668
rect 12760 2648 13153 2668
rect 13324 2665 13361 2744
rect 13391 2773 13422 2826
rect 14171 2798 14857 2831
rect 13441 2773 13478 2774
rect 13391 2764 13478 2773
rect 13391 2744 13449 2764
rect 13469 2744 13478 2764
rect 13391 2734 13478 2744
rect 13537 2764 13574 2774
rect 13537 2744 13545 2764
rect 13565 2744 13574 2764
rect 13391 2733 13422 2734
rect 13386 2665 13496 2678
rect 13537 2665 13574 2744
rect 13324 2663 13574 2665
rect 13324 2660 13425 2663
rect 13324 2641 13389 2660
rect 12204 2628 12283 2636
rect 12115 2626 12283 2628
rect 11839 2619 12283 2626
rect 13386 2633 13389 2641
rect 13418 2633 13425 2660
rect 13453 2636 13463 2663
rect 13492 2641 13574 2663
rect 13763 2710 13931 2711
rect 14171 2710 14209 2798
rect 14470 2796 14517 2798
rect 14817 2774 14857 2798
rect 15196 2822 15236 2846
rect 15536 2822 15583 2824
rect 15844 2822 15882 2910
rect 16122 2909 16290 2910
rect 16479 2957 16561 2979
rect 16590 2957 16600 2984
rect 16628 2960 16635 2987
rect 16664 2979 16667 2987
rect 17770 2994 18214 3020
rect 18442 3015 18553 3021
rect 17770 2992 17938 2994
rect 17770 2990 17889 2992
rect 16664 2960 16729 2979
rect 16628 2957 16729 2960
rect 16479 2955 16729 2957
rect 16479 2876 16516 2955
rect 16557 2942 16667 2955
rect 16631 2886 16662 2887
rect 16479 2856 16488 2876
rect 16508 2856 16516 2876
rect 16479 2846 16516 2856
rect 16575 2876 16662 2886
rect 16575 2856 16584 2876
rect 16604 2856 16662 2876
rect 16575 2847 16662 2856
rect 16575 2846 16612 2847
rect 15196 2789 15882 2822
rect 16631 2794 16662 2847
rect 16692 2876 16729 2955
rect 16900 2974 16932 2986
rect 16900 2954 16902 2974
rect 16923 2972 16932 2974
rect 16923 2970 17275 2972
rect 16923 2954 17293 2970
rect 16900 2952 17293 2954
rect 17313 2952 17316 2970
rect 16900 2947 17316 2952
rect 16900 2946 17241 2947
rect 16844 2886 16875 2887
rect 16692 2856 16701 2876
rect 16721 2856 16729 2876
rect 16692 2846 16729 2856
rect 16788 2879 16875 2886
rect 16788 2876 16849 2879
rect 16788 2856 16797 2876
rect 16817 2859 16849 2876
rect 16870 2859 16875 2879
rect 16817 2856 16875 2859
rect 16788 2849 16875 2856
rect 16900 2876 16937 2946
rect 17203 2945 17240 2946
rect 17052 2886 17088 2887
rect 16900 2856 16909 2876
rect 16929 2856 16937 2876
rect 16788 2847 16844 2849
rect 16788 2846 16825 2847
rect 16900 2846 16937 2856
rect 16996 2876 17144 2886
rect 17244 2883 17340 2885
rect 16996 2856 17005 2876
rect 17025 2867 17115 2876
rect 17025 2856 17056 2867
rect 16996 2847 17056 2856
rect 16996 2846 17033 2847
rect 17052 2835 17056 2847
rect 17083 2856 17115 2867
rect 17135 2856 17144 2876
rect 17083 2847 17144 2856
rect 17202 2876 17340 2883
rect 17202 2856 17211 2876
rect 17231 2856 17340 2876
rect 17202 2847 17340 2856
rect 17083 2835 17088 2847
rect 17107 2846 17144 2847
rect 17203 2846 17240 2847
rect 17052 2795 17088 2835
rect 16523 2793 16564 2794
rect 13763 2687 14209 2710
rect 14435 2741 14546 2755
rect 14435 2739 14477 2741
rect 14435 2719 14442 2739
rect 14461 2719 14477 2739
rect 14435 2711 14477 2719
rect 14505 2739 14546 2741
rect 14505 2719 14519 2739
rect 14538 2719 14546 2739
rect 14818 2730 14857 2774
rect 14505 2711 14546 2719
rect 14435 2705 14546 2711
rect 13763 2684 14207 2687
rect 13763 2682 13931 2684
rect 13492 2636 13496 2641
rect 13453 2633 13496 2636
rect 13386 2619 13496 2633
rect 11500 2599 11611 2605
rect 11839 2600 12209 2619
rect 12115 2599 12209 2600
rect 11500 2591 11541 2599
rect 11500 2571 11508 2591
rect 11527 2571 11541 2591
rect 11500 2569 11541 2571
rect 11569 2591 11611 2599
rect 11569 2571 11585 2591
rect 11604 2571 11611 2591
rect 12204 2590 12209 2599
rect 12257 2599 12283 2619
rect 12257 2590 12274 2599
rect 12204 2581 12274 2590
rect 11569 2569 11611 2571
rect 10948 2565 10984 2566
rect 10796 2535 10805 2555
rect 10825 2535 10833 2555
rect 10684 2526 10740 2528
rect 10684 2525 10721 2526
rect 10796 2525 10833 2535
rect 10892 2555 11040 2565
rect 11140 2562 11236 2564
rect 10892 2535 10901 2555
rect 10921 2535 11011 2555
rect 11031 2535 11040 2555
rect 10892 2526 11040 2535
rect 11098 2555 11236 2562
rect 11098 2535 11107 2555
rect 11127 2535 11236 2555
rect 11500 2554 11611 2569
rect 11098 2526 11236 2535
rect 10892 2525 10929 2526
rect 10948 2474 10984 2526
rect 11003 2525 11040 2526
rect 11099 2525 11136 2526
rect 10419 2472 10460 2473
rect 9841 2460 9882 2469
rect 10311 2465 10460 2472
rect 9841 2440 9881 2460
rect 9398 2430 9648 2432
rect 9398 2427 9499 2430
rect 7916 2370 7980 2382
rect 8256 2378 8293 2405
rect 8464 2378 8501 2409
rect 8677 2407 8713 2409
rect 9398 2408 9463 2427
rect 8677 2378 8714 2407
rect 9460 2400 9463 2408
rect 9492 2400 9499 2427
rect 9527 2403 9537 2430
rect 9566 2408 9648 2430
rect 9756 2430 9881 2440
rect 10311 2445 10429 2465
rect 10449 2445 10460 2465
rect 10311 2437 10460 2445
rect 10527 2469 10886 2473
rect 10527 2464 10849 2469
rect 10527 2440 10640 2464
rect 10664 2445 10849 2464
rect 10873 2445 10886 2469
rect 10664 2440 10886 2445
rect 10527 2437 10886 2440
rect 10948 2437 10983 2474
rect 11051 2471 11151 2474
rect 11051 2467 11118 2471
rect 11051 2441 11063 2467
rect 11089 2445 11118 2467
rect 11144 2445 11151 2471
rect 11089 2441 11151 2445
rect 11051 2437 11151 2441
rect 9756 2411 9764 2430
rect 9789 2411 9881 2430
rect 10527 2416 10558 2437
rect 10948 2416 10984 2437
rect 10370 2415 10407 2416
rect 10144 2412 10178 2413
rect 9566 2403 9570 2408
rect 9756 2404 9881 2411
rect 9527 2400 9570 2403
rect 9460 2386 9570 2400
rect 7916 2369 7951 2370
rect 7893 2364 7951 2369
rect 7893 2344 7896 2364
rect 7916 2350 7951 2364
rect 7971 2350 7980 2370
rect 7916 2342 7980 2350
rect 7942 2341 7980 2342
rect 7943 2340 7980 2341
rect 8046 2374 8082 2375
rect 8154 2374 8190 2375
rect 8046 2366 8190 2374
rect 8046 2346 8054 2366
rect 8074 2346 8162 2366
rect 8182 2346 8190 2366
rect 8046 2340 8190 2346
rect 8256 2370 8294 2378
rect 8362 2374 8398 2375
rect 8256 2350 8265 2370
rect 8285 2350 8294 2370
rect 8256 2341 8294 2350
rect 8313 2367 8398 2374
rect 8313 2347 8320 2367
rect 8341 2366 8398 2367
rect 8341 2347 8370 2366
rect 8313 2346 8370 2347
rect 8390 2346 8398 2366
rect 8256 2340 8293 2341
rect 8313 2340 8398 2346
rect 8464 2370 8502 2378
rect 8575 2374 8611 2375
rect 8464 2350 8473 2370
rect 8493 2350 8502 2370
rect 8464 2341 8502 2350
rect 8526 2366 8611 2374
rect 8526 2346 8583 2366
rect 8603 2346 8611 2366
rect 8464 2340 8501 2341
rect 8526 2340 8611 2346
rect 8677 2370 8715 2378
rect 8677 2350 8686 2370
rect 8706 2350 8715 2370
rect 8677 2341 8715 2350
rect 9841 2356 9881 2404
rect 10143 2403 10180 2412
rect 10143 2385 10152 2403
rect 10170 2385 10180 2403
rect 10143 2375 10180 2385
rect 10369 2406 10407 2415
rect 10369 2386 10378 2406
rect 10398 2386 10407 2406
rect 10369 2378 10407 2386
rect 10473 2410 10558 2416
rect 10583 2415 10620 2416
rect 10473 2390 10481 2410
rect 10501 2390 10558 2410
rect 10473 2382 10558 2390
rect 10582 2406 10620 2415
rect 10582 2386 10591 2406
rect 10611 2386 10620 2406
rect 10473 2381 10509 2382
rect 10582 2378 10620 2386
rect 10686 2410 10771 2416
rect 10791 2415 10828 2416
rect 10686 2390 10694 2410
rect 10714 2409 10771 2410
rect 10714 2390 10743 2409
rect 10686 2389 10743 2390
rect 10764 2389 10771 2409
rect 10686 2382 10771 2389
rect 10790 2406 10828 2415
rect 10790 2386 10799 2406
rect 10819 2386 10828 2406
rect 10686 2381 10722 2382
rect 10790 2378 10828 2386
rect 10894 2410 11038 2416
rect 10894 2390 10902 2410
rect 10922 2409 11010 2410
rect 10922 2390 10953 2409
rect 10894 2389 10953 2390
rect 10978 2390 11010 2409
rect 11030 2390 11038 2410
rect 10978 2389 11038 2390
rect 10894 2382 11038 2389
rect 10894 2381 10930 2382
rect 11002 2381 11038 2382
rect 11104 2415 11141 2416
rect 11104 2414 11142 2415
rect 11104 2406 11168 2414
rect 11104 2386 11113 2406
rect 11133 2392 11168 2406
rect 11188 2392 11191 2412
rect 11133 2387 11191 2392
rect 11133 2386 11168 2387
rect 8677 2340 8714 2341
rect 8100 2319 8136 2340
rect 8526 2319 8557 2340
rect 9841 2338 9852 2356
rect 9870 2338 9881 2356
rect 9841 2330 9881 2338
rect 10144 2347 10178 2375
rect 10370 2349 10407 2378
rect 10371 2347 10407 2349
rect 10583 2347 10620 2378
rect 10144 2346 10316 2347
rect 9842 2329 9879 2330
rect 7933 2315 8033 2319
rect 7933 2311 7995 2315
rect 7933 2285 7940 2311
rect 7966 2289 7995 2311
rect 8021 2289 8033 2315
rect 7966 2285 8033 2289
rect 7933 2282 8033 2285
rect 8101 2282 8136 2319
rect 8198 2316 8557 2319
rect 8198 2311 8420 2316
rect 8198 2287 8211 2311
rect 8235 2292 8420 2311
rect 8444 2292 8557 2316
rect 8235 2287 8557 2292
rect 8198 2283 8557 2287
rect 8624 2311 8773 2319
rect 8624 2291 8635 2311
rect 8655 2291 8773 2311
rect 8624 2284 8773 2291
rect 10144 2314 10330 2346
rect 10371 2325 10620 2347
rect 10791 2346 10828 2378
rect 11104 2374 11168 2386
rect 11208 2348 11235 2526
rect 13763 2504 13790 2682
rect 13830 2644 13894 2656
rect 14170 2652 14207 2684
rect 14378 2683 14627 2705
rect 14378 2652 14415 2683
rect 14591 2681 14627 2683
rect 14591 2652 14628 2681
rect 13830 2643 13865 2644
rect 13807 2638 13865 2643
rect 13807 2618 13810 2638
rect 13830 2624 13865 2638
rect 13885 2624 13894 2644
rect 13830 2616 13894 2624
rect 13856 2615 13894 2616
rect 13857 2614 13894 2615
rect 13960 2648 13996 2649
rect 14068 2648 14104 2649
rect 13960 2643 14104 2648
rect 13960 2640 14022 2643
rect 13960 2620 13968 2640
rect 13988 2623 14022 2640
rect 14045 2640 14104 2643
rect 14045 2623 14076 2640
rect 13988 2620 14076 2623
rect 14096 2620 14104 2640
rect 13960 2614 14104 2620
rect 14170 2644 14208 2652
rect 14276 2648 14312 2649
rect 14170 2624 14179 2644
rect 14199 2624 14208 2644
rect 14170 2615 14208 2624
rect 14227 2641 14312 2648
rect 14227 2621 14234 2641
rect 14255 2640 14312 2641
rect 14255 2621 14284 2640
rect 14227 2620 14284 2621
rect 14304 2620 14312 2640
rect 14170 2614 14207 2615
rect 14227 2614 14312 2620
rect 14378 2644 14416 2652
rect 14489 2648 14525 2649
rect 14378 2624 14387 2644
rect 14407 2624 14416 2644
rect 14378 2615 14416 2624
rect 14440 2640 14525 2648
rect 14440 2620 14497 2640
rect 14517 2620 14525 2640
rect 14378 2614 14415 2615
rect 14440 2614 14525 2620
rect 14591 2644 14629 2652
rect 14591 2624 14600 2644
rect 14620 2624 14629 2644
rect 14591 2615 14629 2624
rect 14591 2614 14628 2615
rect 14014 2593 14050 2614
rect 14440 2593 14471 2614
rect 13847 2589 13947 2593
rect 13847 2585 13909 2589
rect 13847 2559 13854 2585
rect 13880 2563 13909 2585
rect 13935 2563 13947 2589
rect 13880 2559 13947 2563
rect 13847 2556 13947 2559
rect 14015 2556 14050 2593
rect 14112 2590 14471 2593
rect 14112 2585 14334 2590
rect 14112 2561 14125 2585
rect 14149 2566 14334 2585
rect 14358 2566 14471 2590
rect 14149 2561 14471 2566
rect 14112 2557 14471 2561
rect 14538 2585 14687 2593
rect 14538 2565 14549 2585
rect 14569 2565 14687 2585
rect 14538 2558 14687 2565
rect 14538 2557 14579 2558
rect 13862 2504 13899 2505
rect 13958 2504 13995 2505
rect 14014 2504 14050 2556
rect 14069 2504 14106 2505
rect 13762 2495 13900 2504
rect 13762 2475 13871 2495
rect 13891 2475 13900 2495
rect 13762 2468 13900 2475
rect 13958 2495 14106 2504
rect 13958 2475 13967 2495
rect 13987 2475 14077 2495
rect 14097 2475 14106 2495
rect 13762 2466 13858 2468
rect 13958 2465 14106 2475
rect 14165 2495 14202 2505
rect 14277 2504 14314 2505
rect 14258 2502 14314 2504
rect 14165 2475 14173 2495
rect 14193 2475 14202 2495
rect 14014 2464 14050 2465
rect 11391 2422 11501 2436
rect 11391 2419 11434 2422
rect 11391 2414 11395 2419
rect 11067 2346 11235 2348
rect 10791 2340 11235 2346
rect 9213 2288 9727 2289
rect 8624 2283 8665 2284
rect 8100 2247 8136 2282
rect 7948 2230 7985 2231
rect 8044 2230 8081 2231
rect 8100 2230 8107 2247
rect 7848 2221 7986 2230
rect 7848 2201 7957 2221
rect 7977 2201 7986 2221
rect 7848 2194 7986 2201
rect 8044 2221 8107 2230
rect 8044 2201 8053 2221
rect 8073 2206 8107 2221
rect 8128 2230 8136 2247
rect 8155 2230 8192 2231
rect 8128 2221 8192 2230
rect 8128 2206 8163 2221
rect 8073 2201 8163 2206
rect 8183 2201 8192 2221
rect 7848 2192 7944 2194
rect 8044 2191 8192 2201
rect 8251 2221 8288 2231
rect 8363 2230 8400 2231
rect 8344 2228 8400 2230
rect 8251 2201 8259 2221
rect 8279 2201 8288 2221
rect 8100 2190 8136 2191
rect 7030 2138 7198 2140
rect 6752 2132 7198 2138
rect 5820 2108 6236 2113
rect 6415 2111 6526 2117
rect 5820 2107 6161 2108
rect 5764 2047 5795 2048
rect 5612 2017 5621 2037
rect 5641 2017 5649 2037
rect 5612 2007 5649 2017
rect 5708 2040 5795 2047
rect 5708 2037 5769 2040
rect 5708 2017 5717 2037
rect 5737 2020 5769 2037
rect 5790 2020 5795 2040
rect 5737 2017 5795 2020
rect 5708 2010 5795 2017
rect 5820 2037 5857 2107
rect 6123 2106 6160 2107
rect 6415 2103 6456 2111
rect 6415 2083 6423 2103
rect 6442 2083 6456 2103
rect 6415 2081 6456 2083
rect 6484 2103 6526 2111
rect 6484 2083 6500 2103
rect 6519 2083 6526 2103
rect 6752 2110 6758 2132
rect 6784 2112 7198 2132
rect 7948 2131 7985 2132
rect 8251 2131 8288 2201
rect 8313 2221 8400 2228
rect 8313 2218 8371 2221
rect 8313 2198 8318 2218
rect 8339 2201 8371 2218
rect 8391 2201 8400 2221
rect 8339 2198 8400 2201
rect 8313 2191 8400 2198
rect 8459 2221 8496 2231
rect 8459 2201 8467 2221
rect 8487 2201 8496 2221
rect 8313 2190 8344 2191
rect 7947 2130 8288 2131
rect 6784 2110 6793 2112
rect 7030 2111 7198 2112
rect 7872 2129 8288 2130
rect 7872 2125 8248 2129
rect 6752 2101 6793 2110
rect 7872 2105 7875 2125
rect 7895 2112 8248 2125
rect 8280 2112 8288 2129
rect 7895 2105 8288 2112
rect 8459 2122 8496 2201
rect 8526 2230 8557 2283
rect 9194 2272 9727 2288
rect 10144 2282 10178 2314
rect 10140 2273 10178 2282
rect 9194 2261 9726 2272
rect 9845 2263 9882 2267
rect 8576 2230 8613 2231
rect 8526 2221 8613 2230
rect 8526 2201 8584 2221
rect 8604 2201 8613 2221
rect 8526 2191 8613 2201
rect 8672 2221 8709 2231
rect 8672 2201 8680 2221
rect 8700 2201 8709 2221
rect 8526 2190 8557 2191
rect 8521 2122 8631 2135
rect 8672 2122 8709 2201
rect 8459 2120 8709 2122
rect 8459 2117 8560 2120
rect 8459 2098 8524 2117
rect 6484 2081 6526 2083
rect 6415 2066 6526 2081
rect 8521 2090 8524 2098
rect 8553 2090 8560 2117
rect 8588 2093 8598 2120
rect 8627 2098 8709 2120
rect 8787 2192 8955 2193
rect 9194 2192 9232 2261
rect 8787 2172 9232 2192
rect 9459 2223 9570 2238
rect 9459 2221 9501 2223
rect 9459 2201 9466 2221
rect 9485 2201 9501 2221
rect 9459 2193 9501 2201
rect 9529 2221 9570 2223
rect 9529 2201 9543 2221
rect 9562 2201 9570 2221
rect 9529 2193 9570 2201
rect 9459 2187 9570 2193
rect 9692 2198 9726 2261
rect 9844 2257 9882 2263
rect 9844 2239 9854 2257
rect 9872 2239 9882 2257
rect 10140 2255 10150 2273
rect 10168 2255 10178 2273
rect 10140 2249 10178 2255
rect 10296 2251 10330 2314
rect 10452 2319 10563 2325
rect 10452 2311 10493 2319
rect 10452 2291 10460 2311
rect 10479 2291 10493 2311
rect 10452 2289 10493 2291
rect 10521 2311 10563 2319
rect 10521 2291 10537 2311
rect 10556 2291 10563 2311
rect 10521 2289 10563 2291
rect 10452 2274 10563 2289
rect 10790 2320 11235 2340
rect 10790 2251 10828 2320
rect 11067 2319 11235 2320
rect 11313 2392 11395 2414
rect 11424 2392 11434 2419
rect 11462 2395 11469 2422
rect 11498 2414 11501 2422
rect 13496 2431 13607 2446
rect 13496 2429 13538 2431
rect 11498 2395 11563 2414
rect 11462 2392 11563 2395
rect 11313 2390 11563 2392
rect 11313 2311 11350 2390
rect 11391 2377 11501 2390
rect 11465 2321 11496 2322
rect 11313 2291 11322 2311
rect 11342 2291 11350 2311
rect 11313 2281 11350 2291
rect 11409 2311 11496 2321
rect 11409 2291 11418 2311
rect 11438 2291 11496 2311
rect 11409 2282 11496 2291
rect 11409 2281 11446 2282
rect 10140 2245 10177 2249
rect 10296 2240 10828 2251
rect 9844 2230 9882 2239
rect 9844 2198 9878 2230
rect 10295 2224 10828 2240
rect 11465 2229 11496 2282
rect 11526 2311 11563 2390
rect 11734 2387 12127 2407
rect 12147 2387 12150 2407
rect 13229 2402 13270 2411
rect 11734 2382 12150 2387
rect 12824 2400 12992 2401
rect 13229 2400 13238 2402
rect 11734 2381 12075 2382
rect 11678 2321 11709 2322
rect 11526 2291 11535 2311
rect 11555 2291 11563 2311
rect 11526 2281 11563 2291
rect 11622 2314 11709 2321
rect 11622 2311 11683 2314
rect 11622 2291 11631 2311
rect 11651 2294 11683 2311
rect 11704 2294 11709 2314
rect 11651 2291 11709 2294
rect 11622 2284 11709 2291
rect 11734 2311 11771 2381
rect 12037 2380 12074 2381
rect 12824 2380 13238 2400
rect 13264 2380 13270 2402
rect 13496 2409 13503 2429
rect 13522 2409 13538 2429
rect 13496 2401 13538 2409
rect 13566 2429 13607 2431
rect 13566 2409 13580 2429
rect 13599 2409 13607 2429
rect 13566 2401 13607 2409
rect 13862 2405 13899 2406
rect 14165 2405 14202 2475
rect 14227 2495 14314 2502
rect 14227 2492 14285 2495
rect 14227 2472 14232 2492
rect 14253 2475 14285 2492
rect 14305 2475 14314 2495
rect 14253 2472 14314 2475
rect 14227 2465 14314 2472
rect 14373 2495 14410 2505
rect 14373 2475 14381 2495
rect 14401 2475 14410 2495
rect 14227 2464 14258 2465
rect 13861 2404 14202 2405
rect 13496 2395 13607 2401
rect 13786 2399 14202 2404
rect 12824 2374 13270 2380
rect 12824 2372 12992 2374
rect 11886 2321 11922 2322
rect 11734 2291 11743 2311
rect 11763 2291 11771 2311
rect 11622 2282 11678 2284
rect 11622 2281 11659 2282
rect 11734 2281 11771 2291
rect 11830 2311 11978 2321
rect 12078 2318 12174 2320
rect 11830 2291 11839 2311
rect 11859 2291 11949 2311
rect 11969 2291 11978 2311
rect 11830 2282 11978 2291
rect 12036 2311 12174 2318
rect 12036 2291 12045 2311
rect 12065 2291 12174 2311
rect 12036 2282 12174 2291
rect 11830 2281 11867 2282
rect 11886 2230 11922 2282
rect 11941 2281 11978 2282
rect 12037 2281 12074 2282
rect 11357 2228 11398 2229
rect 10295 2223 10809 2224
rect 8787 2166 9231 2172
rect 8787 2164 8955 2166
rect 8627 2093 8631 2098
rect 8588 2090 8631 2093
rect 8521 2076 8631 2090
rect 5972 2047 6008 2048
rect 5820 2017 5829 2037
rect 5849 2017 5857 2037
rect 5708 2008 5764 2010
rect 5708 2007 5745 2008
rect 5820 2007 5857 2017
rect 5916 2037 6064 2047
rect 6164 2044 6260 2046
rect 5916 2017 5925 2037
rect 5945 2017 6035 2037
rect 6055 2017 6064 2037
rect 5916 2008 6064 2017
rect 6122 2037 6260 2044
rect 6122 2017 6131 2037
rect 6151 2017 6260 2037
rect 6122 2008 6260 2017
rect 5916 2007 5953 2008
rect 5972 1956 6008 2008
rect 6027 2007 6064 2008
rect 6123 2007 6160 2008
rect 5443 1954 5484 1955
rect 5335 1947 5484 1954
rect 5335 1927 5453 1947
rect 5473 1927 5484 1947
rect 5335 1919 5484 1927
rect 5551 1951 5910 1955
rect 5551 1946 5873 1951
rect 5551 1922 5664 1946
rect 5688 1927 5873 1946
rect 5897 1927 5910 1951
rect 5688 1922 5910 1927
rect 5551 1919 5910 1922
rect 5972 1919 6007 1956
rect 6075 1953 6175 1956
rect 6075 1949 6142 1953
rect 6075 1923 6087 1949
rect 6113 1927 6142 1949
rect 6168 1927 6175 1953
rect 6113 1923 6175 1927
rect 6075 1919 6175 1923
rect 5551 1898 5582 1919
rect 5972 1898 6008 1919
rect 5394 1897 5431 1898
rect 5393 1888 5431 1897
rect 5393 1868 5402 1888
rect 5422 1868 5431 1888
rect 5393 1860 5431 1868
rect 5497 1892 5582 1898
rect 5607 1897 5644 1898
rect 5497 1872 5505 1892
rect 5525 1872 5582 1892
rect 5497 1864 5582 1872
rect 5606 1888 5644 1897
rect 5606 1868 5615 1888
rect 5635 1868 5644 1888
rect 5497 1863 5533 1864
rect 5606 1860 5644 1868
rect 5710 1892 5795 1898
rect 5815 1897 5852 1898
rect 5710 1872 5718 1892
rect 5738 1891 5795 1892
rect 5738 1872 5767 1891
rect 5710 1871 5767 1872
rect 5788 1871 5795 1891
rect 5710 1864 5795 1871
rect 5814 1888 5852 1897
rect 5814 1868 5823 1888
rect 5843 1868 5852 1888
rect 5710 1863 5746 1864
rect 5814 1860 5852 1868
rect 5918 1892 6062 1898
rect 5918 1872 5926 1892
rect 5946 1889 6034 1892
rect 5946 1872 5977 1889
rect 5918 1869 5977 1872
rect 6000 1872 6034 1889
rect 6054 1872 6062 1892
rect 6000 1869 6062 1872
rect 5918 1864 6062 1869
rect 5918 1863 5954 1864
rect 6026 1863 6062 1864
rect 6128 1897 6165 1898
rect 6128 1896 6166 1897
rect 6128 1888 6192 1896
rect 6128 1868 6137 1888
rect 6157 1874 6192 1888
rect 6212 1874 6215 1894
rect 6157 1869 6215 1874
rect 6157 1868 6192 1869
rect 5394 1831 5431 1860
rect 5395 1829 5431 1831
rect 5607 1829 5644 1860
rect 5395 1807 5644 1829
rect 5815 1828 5852 1860
rect 6128 1856 6192 1868
rect 6232 1830 6259 2008
rect 8787 1986 8814 2164
rect 8854 2126 8918 2138
rect 9194 2134 9231 2166
rect 9402 2165 9651 2187
rect 9692 2166 9878 2198
rect 11249 2221 11398 2228
rect 11249 2201 11367 2221
rect 11387 2201 11398 2221
rect 11249 2193 11398 2201
rect 11465 2225 11824 2229
rect 11465 2220 11787 2225
rect 11465 2196 11578 2220
rect 11602 2201 11787 2220
rect 11811 2201 11824 2225
rect 11602 2196 11824 2201
rect 11465 2193 11824 2196
rect 11886 2193 11921 2230
rect 11989 2227 12089 2230
rect 11989 2223 12056 2227
rect 11989 2197 12001 2223
rect 12027 2201 12056 2223
rect 12082 2201 12089 2227
rect 12027 2197 12089 2201
rect 11989 2193 12089 2197
rect 10143 2182 10180 2183
rect 9706 2165 9878 2166
rect 9402 2134 9439 2165
rect 9615 2163 9651 2165
rect 9615 2134 9652 2163
rect 9844 2137 9878 2165
rect 10141 2174 10181 2182
rect 10141 2156 10152 2174
rect 10170 2156 10181 2174
rect 11465 2172 11496 2193
rect 11886 2172 11922 2193
rect 11308 2171 11345 2172
rect 8854 2125 8889 2126
rect 8831 2120 8889 2125
rect 8831 2100 8834 2120
rect 8854 2106 8889 2120
rect 8909 2106 8918 2126
rect 8854 2098 8918 2106
rect 8880 2097 8918 2098
rect 8881 2096 8918 2097
rect 8984 2130 9020 2131
rect 9092 2130 9128 2131
rect 8984 2123 9128 2130
rect 8984 2122 9044 2123
rect 8984 2102 8992 2122
rect 9012 2103 9044 2122
rect 9069 2122 9128 2123
rect 9069 2103 9100 2122
rect 9012 2102 9100 2103
rect 9120 2102 9128 2122
rect 8984 2096 9128 2102
rect 9194 2126 9232 2134
rect 9300 2130 9336 2131
rect 9194 2106 9203 2126
rect 9223 2106 9232 2126
rect 9194 2097 9232 2106
rect 9251 2123 9336 2130
rect 9251 2103 9258 2123
rect 9279 2122 9336 2123
rect 9279 2103 9308 2122
rect 9251 2102 9308 2103
rect 9328 2102 9336 2122
rect 9194 2096 9231 2097
rect 9251 2096 9336 2102
rect 9402 2126 9440 2134
rect 9513 2130 9549 2131
rect 9402 2106 9411 2126
rect 9431 2106 9440 2126
rect 9402 2097 9440 2106
rect 9464 2122 9549 2130
rect 9464 2102 9521 2122
rect 9541 2102 9549 2122
rect 9402 2096 9439 2097
rect 9464 2096 9549 2102
rect 9615 2126 9653 2134
rect 9615 2106 9624 2126
rect 9644 2106 9653 2126
rect 9615 2097 9653 2106
rect 9842 2127 9879 2137
rect 9842 2109 9852 2127
rect 9870 2109 9879 2127
rect 9842 2100 9879 2109
rect 10141 2108 10181 2156
rect 11307 2162 11345 2171
rect 11307 2142 11316 2162
rect 11336 2142 11345 2162
rect 11307 2134 11345 2142
rect 11411 2166 11496 2172
rect 11521 2171 11558 2172
rect 11411 2146 11419 2166
rect 11439 2146 11496 2166
rect 11411 2138 11496 2146
rect 11520 2162 11558 2171
rect 11520 2142 11529 2162
rect 11549 2142 11558 2162
rect 11411 2137 11447 2138
rect 11520 2134 11558 2142
rect 11624 2166 11709 2172
rect 11729 2171 11766 2172
rect 11624 2146 11632 2166
rect 11652 2165 11709 2166
rect 11652 2146 11681 2165
rect 11624 2145 11681 2146
rect 11702 2145 11709 2165
rect 11624 2138 11709 2145
rect 11728 2162 11766 2171
rect 11728 2142 11737 2162
rect 11757 2142 11766 2162
rect 11624 2137 11660 2138
rect 11728 2134 11766 2142
rect 11832 2166 11976 2172
rect 11832 2146 11840 2166
rect 11860 2149 11896 2166
rect 11916 2149 11948 2166
rect 11860 2146 11948 2149
rect 11968 2146 11976 2166
rect 11832 2138 11976 2146
rect 11832 2137 11868 2138
rect 11940 2137 11976 2138
rect 12042 2171 12079 2172
rect 12042 2170 12080 2171
rect 12042 2162 12106 2170
rect 12042 2142 12051 2162
rect 12071 2148 12106 2162
rect 12126 2148 12129 2168
rect 12071 2143 12129 2148
rect 12071 2142 12106 2143
rect 10452 2112 10562 2126
rect 10452 2109 10495 2112
rect 10141 2101 10266 2108
rect 10452 2104 10456 2109
rect 9844 2099 9878 2100
rect 9615 2096 9652 2097
rect 9038 2075 9074 2096
rect 9464 2075 9495 2096
rect 10141 2082 10233 2101
rect 10258 2082 10266 2101
rect 8871 2071 8971 2075
rect 8871 2067 8933 2071
rect 8871 2041 8878 2067
rect 8904 2045 8933 2067
rect 8959 2045 8971 2071
rect 8904 2041 8971 2045
rect 8871 2038 8971 2041
rect 9039 2038 9074 2075
rect 9136 2072 9495 2075
rect 9136 2067 9358 2072
rect 9136 2043 9149 2067
rect 9173 2048 9358 2067
rect 9382 2048 9495 2072
rect 9173 2043 9495 2048
rect 9136 2039 9495 2043
rect 9562 2067 9711 2075
rect 9562 2047 9573 2067
rect 9593 2047 9711 2067
rect 10141 2072 10266 2082
rect 10374 2082 10456 2104
rect 10485 2082 10495 2109
rect 10523 2085 10530 2112
rect 10559 2104 10562 2112
rect 11308 2105 11345 2134
rect 10559 2085 10624 2104
rect 11309 2103 11345 2105
rect 11521 2103 11558 2134
rect 11729 2107 11766 2134
rect 12042 2130 12106 2142
rect 10523 2082 10624 2085
rect 10374 2080 10624 2082
rect 10141 2052 10181 2072
rect 9562 2040 9711 2047
rect 10140 2043 10181 2052
rect 9562 2039 9603 2040
rect 8886 1986 8923 1987
rect 8982 1986 9019 1987
rect 9038 1986 9074 2038
rect 9093 1986 9130 1987
rect 8786 1977 8924 1986
rect 8381 1956 8492 1971
rect 8381 1954 8423 1956
rect 8051 1933 8156 1935
rect 7709 1925 7877 1926
rect 8051 1925 8100 1933
rect 7709 1906 8100 1925
rect 8131 1906 8156 1933
rect 8381 1934 8388 1954
rect 8407 1934 8423 1954
rect 8381 1926 8423 1934
rect 8451 1954 8492 1956
rect 8451 1934 8465 1954
rect 8484 1934 8492 1954
rect 8786 1957 8895 1977
rect 8915 1957 8924 1977
rect 8786 1950 8924 1957
rect 8982 1977 9130 1986
rect 8982 1957 8991 1977
rect 9011 1957 9101 1977
rect 9121 1957 9130 1977
rect 8786 1948 8882 1950
rect 8982 1947 9130 1957
rect 9189 1977 9226 1987
rect 9301 1986 9338 1987
rect 9282 1984 9338 1986
rect 9189 1957 9197 1977
rect 9217 1957 9226 1977
rect 9038 1946 9074 1947
rect 8451 1926 8492 1934
rect 8381 1920 8492 1926
rect 7709 1899 8156 1906
rect 7709 1897 7877 1899
rect 6557 1866 6667 1880
rect 6557 1863 6600 1866
rect 6557 1858 6561 1863
rect 6091 1828 6259 1830
rect 5815 1825 6259 1828
rect 5476 1801 5587 1807
rect 5476 1793 5517 1801
rect 5165 1738 5204 1782
rect 5476 1773 5484 1793
rect 5503 1773 5517 1793
rect 5476 1771 5517 1773
rect 5545 1793 5587 1801
rect 5545 1773 5561 1793
rect 5580 1773 5587 1793
rect 5545 1771 5587 1773
rect 5476 1756 5587 1771
rect 5813 1802 6259 1825
rect 5165 1714 5205 1738
rect 5505 1714 5552 1716
rect 5813 1714 5851 1802
rect 6091 1801 6259 1802
rect 6479 1836 6561 1858
rect 6590 1836 6600 1863
rect 6628 1839 6635 1866
rect 6664 1858 6667 1866
rect 6664 1839 6729 1858
rect 6628 1836 6729 1839
rect 6479 1834 6729 1836
rect 6479 1755 6516 1834
rect 6557 1821 6667 1834
rect 6631 1765 6662 1766
rect 6479 1735 6488 1755
rect 6508 1735 6516 1755
rect 6479 1725 6516 1735
rect 6575 1755 6662 1765
rect 6575 1735 6584 1755
rect 6604 1735 6662 1755
rect 6575 1726 6662 1735
rect 6575 1725 6612 1726
rect 5165 1681 5851 1714
rect 5165 1624 5204 1681
rect 5813 1679 5851 1681
rect 6631 1673 6662 1726
rect 6692 1755 6729 1834
rect 6900 1847 7293 1851
rect 6900 1830 6919 1847
rect 6939 1831 7293 1847
rect 7313 1831 7316 1851
rect 6939 1830 7316 1831
rect 6900 1826 7316 1830
rect 6900 1825 7241 1826
rect 6844 1765 6875 1766
rect 6692 1735 6701 1755
rect 6721 1735 6729 1755
rect 6692 1725 6729 1735
rect 6788 1758 6875 1765
rect 6788 1755 6849 1758
rect 6788 1735 6797 1755
rect 6817 1738 6849 1755
rect 6870 1738 6875 1758
rect 6817 1735 6875 1738
rect 6788 1728 6875 1735
rect 6900 1755 6937 1825
rect 7203 1824 7240 1825
rect 7052 1765 7088 1766
rect 6900 1735 6909 1755
rect 6929 1735 6937 1755
rect 6788 1726 6844 1728
rect 6788 1725 6825 1726
rect 6900 1725 6937 1735
rect 6996 1755 7144 1765
rect 7312 1764 7341 1765
rect 7244 1762 7341 1764
rect 6996 1735 7005 1755
rect 7025 1751 7115 1755
rect 7025 1735 7058 1751
rect 6996 1726 7058 1735
rect 6996 1725 7033 1726
rect 7052 1713 7058 1726
rect 7081 1735 7115 1751
rect 7135 1735 7144 1755
rect 7081 1726 7144 1735
rect 7202 1755 7341 1762
rect 7202 1735 7211 1755
rect 7231 1735 7341 1755
rect 7202 1726 7341 1735
rect 7081 1713 7088 1726
rect 7107 1725 7144 1726
rect 7203 1725 7240 1726
rect 7052 1674 7088 1713
rect 6523 1672 6564 1673
rect 6415 1665 6564 1672
rect 6415 1645 6533 1665
rect 6553 1645 6564 1665
rect 6415 1637 6564 1645
rect 6631 1669 6990 1673
rect 6631 1664 6953 1669
rect 6631 1640 6744 1664
rect 6768 1645 6953 1664
rect 6977 1645 6990 1669
rect 6768 1640 6990 1645
rect 6631 1637 6990 1640
rect 7052 1637 7087 1674
rect 7155 1671 7255 1674
rect 7155 1667 7222 1671
rect 7155 1641 7167 1667
rect 7193 1645 7222 1667
rect 7248 1645 7255 1671
rect 7193 1641 7255 1645
rect 7155 1637 7255 1641
rect 5165 1622 5213 1624
rect 5165 1604 5176 1622
rect 5194 1604 5213 1622
rect 6631 1616 6662 1637
rect 7052 1616 7088 1637
rect 6474 1615 6511 1616
rect 5165 1595 5213 1604
rect 5166 1594 5213 1595
rect 5479 1599 5589 1613
rect 5479 1596 5522 1599
rect 5479 1591 5483 1596
rect 5401 1569 5483 1591
rect 5512 1569 5522 1596
rect 5550 1572 5557 1599
rect 5586 1591 5589 1599
rect 6473 1606 6511 1615
rect 5586 1572 5651 1591
rect 6473 1586 6482 1606
rect 6502 1586 6511 1606
rect 5550 1569 5651 1572
rect 5401 1567 5651 1569
rect 5169 1531 5206 1532
rect 4787 1424 4797 1442
rect 4815 1424 4827 1442
rect 4787 1419 4827 1424
rect 5165 1528 5206 1531
rect 5165 1523 5207 1528
rect 5165 1505 5178 1523
rect 5196 1505 5207 1523
rect 5165 1491 5207 1505
rect 5245 1491 5292 1495
rect 5165 1485 5292 1491
rect 5165 1456 5253 1485
rect 5282 1456 5292 1485
rect 5401 1488 5438 1567
rect 5479 1554 5589 1567
rect 5553 1498 5584 1499
rect 5401 1468 5410 1488
rect 5430 1468 5438 1488
rect 5401 1458 5438 1468
rect 5497 1488 5584 1498
rect 5497 1468 5506 1488
rect 5526 1468 5584 1488
rect 5497 1459 5584 1468
rect 5497 1458 5534 1459
rect 5165 1452 5292 1456
rect 5165 1435 5204 1452
rect 5245 1451 5292 1452
rect 4787 1415 4824 1419
rect 5165 1417 5176 1435
rect 5194 1417 5204 1435
rect 5165 1408 5204 1417
rect 5166 1407 5203 1408
rect 5553 1406 5584 1459
rect 5614 1488 5651 1567
rect 5822 1564 6215 1584
rect 6235 1564 6238 1584
rect 6473 1578 6511 1586
rect 6577 1610 6662 1616
rect 6687 1615 6724 1616
rect 6577 1590 6585 1610
rect 6605 1590 6662 1610
rect 6577 1582 6662 1590
rect 6686 1606 6724 1615
rect 6686 1586 6695 1606
rect 6715 1586 6724 1606
rect 6577 1581 6613 1582
rect 6686 1578 6724 1586
rect 6790 1610 6875 1616
rect 6895 1615 6932 1616
rect 6790 1590 6798 1610
rect 6818 1609 6875 1610
rect 6818 1590 6847 1609
rect 6790 1589 6847 1590
rect 6868 1589 6875 1609
rect 6790 1582 6875 1589
rect 6894 1606 6932 1615
rect 6894 1586 6903 1606
rect 6923 1586 6932 1606
rect 6790 1581 6826 1582
rect 6894 1578 6932 1586
rect 6998 1610 7142 1616
rect 6998 1590 7006 1610
rect 7026 1590 7114 1610
rect 7134 1590 7142 1610
rect 6998 1582 7142 1590
rect 6998 1581 7034 1582
rect 7106 1581 7142 1582
rect 7208 1615 7245 1616
rect 7208 1614 7246 1615
rect 7208 1606 7272 1614
rect 7208 1586 7217 1606
rect 7237 1592 7272 1606
rect 7292 1592 7295 1612
rect 7237 1587 7295 1592
rect 7237 1586 7272 1587
rect 5822 1559 6238 1564
rect 5822 1558 6163 1559
rect 5766 1498 5797 1499
rect 5614 1468 5623 1488
rect 5643 1468 5651 1488
rect 5614 1458 5651 1468
rect 5710 1491 5797 1498
rect 5710 1488 5771 1491
rect 5710 1468 5719 1488
rect 5739 1471 5771 1488
rect 5792 1471 5797 1491
rect 5739 1468 5797 1471
rect 5710 1461 5797 1468
rect 5822 1488 5859 1558
rect 6125 1557 6162 1558
rect 6474 1549 6511 1578
rect 6475 1547 6511 1549
rect 6687 1547 6724 1578
rect 6475 1525 6724 1547
rect 6895 1546 6932 1578
rect 7208 1574 7272 1586
rect 7312 1548 7341 1726
rect 7709 1719 7736 1897
rect 7776 1859 7840 1871
rect 8116 1867 8153 1899
rect 8324 1898 8573 1920
rect 8324 1867 8361 1898
rect 8537 1896 8573 1898
rect 8537 1867 8574 1896
rect 8886 1887 8923 1888
rect 9189 1887 9226 1957
rect 9251 1977 9338 1984
rect 9251 1974 9309 1977
rect 9251 1954 9256 1974
rect 9277 1957 9309 1974
rect 9329 1957 9338 1977
rect 9277 1954 9338 1957
rect 9251 1947 9338 1954
rect 9397 1977 9434 1987
rect 9397 1957 9405 1977
rect 9425 1957 9434 1977
rect 9251 1946 9282 1947
rect 8885 1886 9226 1887
rect 8810 1881 9226 1886
rect 7776 1858 7811 1859
rect 7753 1853 7811 1858
rect 7753 1833 7756 1853
rect 7776 1839 7811 1853
rect 7831 1839 7840 1859
rect 7776 1831 7840 1839
rect 7802 1830 7840 1831
rect 7803 1829 7840 1830
rect 7906 1863 7942 1864
rect 8014 1863 8050 1864
rect 7906 1858 8050 1863
rect 7906 1855 7966 1858
rect 7906 1835 7914 1855
rect 7934 1837 7966 1855
rect 7993 1855 8050 1858
rect 7993 1837 8022 1855
rect 7934 1835 8022 1837
rect 8042 1835 8050 1855
rect 7906 1829 8050 1835
rect 8116 1859 8154 1867
rect 8222 1863 8258 1864
rect 8116 1839 8125 1859
rect 8145 1839 8154 1859
rect 8116 1830 8154 1839
rect 8173 1856 8258 1863
rect 8173 1836 8180 1856
rect 8201 1855 8258 1856
rect 8201 1836 8230 1855
rect 8173 1835 8230 1836
rect 8250 1835 8258 1855
rect 8116 1829 8153 1830
rect 8173 1829 8258 1835
rect 8324 1859 8362 1867
rect 8435 1863 8471 1864
rect 8324 1839 8333 1859
rect 8353 1839 8362 1859
rect 8324 1830 8362 1839
rect 8386 1855 8471 1863
rect 8386 1835 8443 1855
rect 8463 1835 8471 1855
rect 8324 1829 8361 1830
rect 8386 1829 8471 1835
rect 8537 1859 8575 1867
rect 8810 1861 8813 1881
rect 8833 1861 9226 1881
rect 9397 1878 9434 1957
rect 9464 1986 9495 2039
rect 9845 2037 9882 2038
rect 9844 2028 9883 2037
rect 9844 2010 9854 2028
rect 9872 2010 9883 2028
rect 10140 2025 10150 2043
rect 10168 2025 10181 2043
rect 10140 2016 10181 2025
rect 10140 2015 10177 2016
rect 9756 1993 9803 1994
rect 9844 1993 9883 2010
rect 9756 1989 9883 1993
rect 9514 1986 9551 1987
rect 9464 1977 9551 1986
rect 9464 1957 9522 1977
rect 9542 1957 9551 1977
rect 9464 1947 9551 1957
rect 9610 1977 9647 1987
rect 9610 1957 9618 1977
rect 9638 1957 9647 1977
rect 9464 1946 9495 1947
rect 9459 1878 9569 1891
rect 9610 1878 9647 1957
rect 9756 1960 9766 1989
rect 9795 1960 9883 1989
rect 10374 2001 10411 2080
rect 10452 2067 10562 2080
rect 10526 2011 10557 2012
rect 10374 1981 10383 2001
rect 10403 1981 10411 2001
rect 10374 1971 10411 1981
rect 10470 2001 10557 2011
rect 10470 1981 10479 2001
rect 10499 1981 10557 2001
rect 10470 1972 10557 1981
rect 10470 1971 10507 1972
rect 9756 1954 9883 1960
rect 9756 1950 9803 1954
rect 9841 1940 9883 1954
rect 10143 1949 10180 1953
rect 9841 1922 9852 1940
rect 9870 1922 9883 1940
rect 9841 1917 9883 1922
rect 9842 1914 9883 1917
rect 10140 1944 10180 1949
rect 10140 1926 10152 1944
rect 10170 1926 10180 1944
rect 9842 1913 9879 1914
rect 9397 1876 9647 1878
rect 9397 1873 9498 1876
rect 8537 1839 8546 1859
rect 8566 1839 8575 1859
rect 9397 1854 9462 1873
rect 8537 1830 8575 1839
rect 9459 1846 9462 1854
rect 9491 1846 9498 1873
rect 9526 1849 9536 1876
rect 9565 1854 9647 1876
rect 9565 1849 9569 1854
rect 9526 1846 9569 1849
rect 9459 1832 9569 1846
rect 9835 1850 9882 1851
rect 9835 1841 9883 1850
rect 8537 1829 8574 1830
rect 7960 1808 7996 1829
rect 8386 1808 8417 1829
rect 9835 1823 9854 1841
rect 9872 1823 9883 1841
rect 9835 1821 9883 1823
rect 7793 1804 7893 1808
rect 7793 1800 7855 1804
rect 7793 1774 7800 1800
rect 7826 1778 7855 1800
rect 7881 1778 7893 1804
rect 7826 1774 7893 1778
rect 7793 1771 7893 1774
rect 7961 1771 7996 1808
rect 8058 1805 8417 1808
rect 8058 1800 8280 1805
rect 8058 1776 8071 1800
rect 8095 1781 8280 1800
rect 8304 1781 8417 1805
rect 8095 1776 8417 1781
rect 8058 1772 8417 1776
rect 8484 1800 8633 1808
rect 8484 1780 8495 1800
rect 8515 1780 8633 1800
rect 8484 1773 8633 1780
rect 8484 1772 8525 1773
rect 7808 1719 7845 1720
rect 7904 1719 7941 1720
rect 7960 1719 7996 1771
rect 8015 1719 8052 1720
rect 7708 1710 7846 1719
rect 7708 1690 7817 1710
rect 7837 1690 7846 1710
rect 7708 1683 7846 1690
rect 7904 1710 8052 1719
rect 7904 1690 7913 1710
rect 7933 1690 8023 1710
rect 8043 1690 8052 1710
rect 7708 1681 7804 1683
rect 7904 1680 8052 1690
rect 8111 1710 8148 1720
rect 8223 1719 8260 1720
rect 8204 1717 8260 1719
rect 8111 1690 8119 1710
rect 8139 1690 8148 1710
rect 7960 1679 7996 1680
rect 7808 1620 7845 1621
rect 8111 1620 8148 1690
rect 8173 1710 8260 1717
rect 8173 1707 8231 1710
rect 8173 1687 8178 1707
rect 8199 1690 8231 1707
rect 8251 1690 8260 1710
rect 8199 1687 8260 1690
rect 8173 1680 8260 1687
rect 8319 1710 8356 1720
rect 8319 1690 8327 1710
rect 8347 1690 8356 1710
rect 8173 1679 8204 1680
rect 7807 1619 8148 1620
rect 7732 1615 8148 1619
rect 7732 1614 8109 1615
rect 7732 1594 7735 1614
rect 7755 1598 8109 1614
rect 8129 1598 8148 1615
rect 7755 1594 8148 1598
rect 8319 1611 8356 1690
rect 8386 1719 8417 1772
rect 9197 1764 9235 1766
rect 9844 1764 9883 1821
rect 9197 1731 9883 1764
rect 8436 1719 8473 1720
rect 8386 1710 8473 1719
rect 8386 1690 8444 1710
rect 8464 1690 8473 1710
rect 8386 1680 8473 1690
rect 8532 1710 8569 1720
rect 8532 1690 8540 1710
rect 8560 1690 8569 1710
rect 8386 1679 8417 1680
rect 8381 1611 8491 1624
rect 8532 1611 8569 1690
rect 8319 1609 8569 1611
rect 8319 1606 8420 1609
rect 8319 1587 8384 1606
rect 8381 1579 8384 1587
rect 8413 1579 8420 1606
rect 8448 1582 8458 1609
rect 8487 1587 8569 1609
rect 8789 1643 8957 1644
rect 9197 1643 9235 1731
rect 9496 1729 9543 1731
rect 9843 1707 9883 1731
rect 8789 1620 9235 1643
rect 9461 1674 9572 1689
rect 9461 1672 9503 1674
rect 9461 1652 9468 1672
rect 9487 1652 9503 1672
rect 9461 1644 9503 1652
rect 9531 1672 9572 1674
rect 9531 1652 9545 1672
rect 9564 1652 9572 1672
rect 9844 1663 9883 1707
rect 9531 1644 9572 1652
rect 9461 1638 9572 1644
rect 8789 1617 9233 1620
rect 8789 1615 8957 1617
rect 8487 1582 8491 1587
rect 8448 1579 8491 1582
rect 8381 1565 8491 1579
rect 7171 1546 7341 1548
rect 6892 1539 7341 1546
rect 6556 1519 6667 1525
rect 6556 1511 6597 1519
rect 5974 1498 6010 1499
rect 5822 1468 5831 1488
rect 5851 1468 5859 1488
rect 5710 1459 5766 1461
rect 5710 1458 5747 1459
rect 5822 1458 5859 1468
rect 5918 1488 6066 1498
rect 6166 1495 6262 1497
rect 5918 1468 5927 1488
rect 5947 1468 6037 1488
rect 6057 1468 6066 1488
rect 5918 1459 6066 1468
rect 6124 1488 6262 1495
rect 6124 1468 6133 1488
rect 6153 1468 6262 1488
rect 6556 1491 6564 1511
rect 6583 1491 6597 1511
rect 6556 1489 6597 1491
rect 6625 1511 6667 1519
rect 6625 1491 6641 1511
rect 6660 1491 6667 1511
rect 6892 1512 6917 1539
rect 6948 1520 7341 1539
rect 6948 1512 6997 1520
rect 7171 1519 7341 1520
rect 6892 1510 6997 1512
rect 6625 1489 6667 1491
rect 6556 1474 6667 1489
rect 6124 1459 6262 1468
rect 5918 1458 5955 1459
rect 5974 1407 6010 1459
rect 6029 1458 6066 1459
rect 6125 1458 6162 1459
rect 5445 1405 5486 1406
rect 5337 1398 5486 1405
rect 4460 1396 4497 1397
rect 4410 1387 4497 1396
rect 4410 1367 4468 1387
rect 4488 1367 4497 1387
rect 4410 1357 4497 1367
rect 4556 1387 4593 1397
rect 4556 1367 4564 1387
rect 4584 1367 4593 1387
rect 5337 1378 5455 1398
rect 5475 1378 5486 1398
rect 5337 1370 5486 1378
rect 5553 1402 5912 1406
rect 5553 1397 5875 1402
rect 5553 1373 5666 1397
rect 5690 1378 5875 1397
rect 5899 1378 5912 1402
rect 5690 1373 5912 1378
rect 5553 1370 5912 1373
rect 5974 1370 6009 1407
rect 6077 1404 6177 1407
rect 6077 1400 6144 1404
rect 6077 1374 6089 1400
rect 6115 1378 6144 1400
rect 6170 1378 6177 1404
rect 6115 1374 6177 1378
rect 6077 1370 6177 1374
rect 4410 1356 4441 1357
rect 4405 1288 4515 1301
rect 4556 1288 4593 1367
rect 4790 1352 4827 1353
rect 4786 1343 4827 1352
rect 5553 1349 5584 1370
rect 5974 1349 6010 1370
rect 5396 1348 5433 1349
rect 5170 1345 5204 1346
rect 4786 1325 4799 1343
rect 4817 1325 4827 1343
rect 4786 1316 4827 1325
rect 5169 1336 5206 1345
rect 5169 1318 5178 1336
rect 5196 1318 5206 1336
rect 4786 1296 4826 1316
rect 5169 1308 5206 1318
rect 5395 1339 5433 1348
rect 5395 1319 5404 1339
rect 5424 1319 5433 1339
rect 5395 1311 5433 1319
rect 5499 1343 5584 1349
rect 5609 1348 5646 1349
rect 5499 1323 5507 1343
rect 5527 1323 5584 1343
rect 5499 1315 5584 1323
rect 5608 1339 5646 1348
rect 5608 1319 5617 1339
rect 5637 1319 5646 1339
rect 5499 1314 5535 1315
rect 5608 1311 5646 1319
rect 5712 1343 5797 1349
rect 5817 1348 5854 1349
rect 5712 1323 5720 1343
rect 5740 1342 5797 1343
rect 5740 1323 5769 1342
rect 5712 1322 5769 1323
rect 5790 1322 5797 1342
rect 5712 1315 5797 1322
rect 5816 1339 5854 1348
rect 5816 1319 5825 1339
rect 5845 1319 5854 1339
rect 5712 1314 5748 1315
rect 5816 1311 5854 1319
rect 5920 1343 6064 1349
rect 5920 1323 5928 1343
rect 5948 1342 6036 1343
rect 5948 1323 5979 1342
rect 5920 1322 5979 1323
rect 6004 1323 6036 1342
rect 6056 1323 6064 1343
rect 6004 1322 6064 1323
rect 5920 1315 6064 1322
rect 5920 1314 5956 1315
rect 6028 1314 6064 1315
rect 6130 1348 6167 1349
rect 6130 1347 6168 1348
rect 6130 1339 6194 1347
rect 6130 1319 6139 1339
rect 6159 1325 6194 1339
rect 6214 1325 6217 1345
rect 6159 1320 6217 1325
rect 6159 1319 6194 1320
rect 4343 1286 4593 1288
rect 4343 1283 4444 1286
rect 2861 1226 2925 1238
rect 3201 1234 3238 1261
rect 3409 1234 3446 1265
rect 3622 1263 3658 1265
rect 4343 1264 4408 1283
rect 3622 1234 3659 1263
rect 4405 1256 4408 1264
rect 4437 1256 4444 1283
rect 4472 1259 4482 1286
rect 4511 1264 4593 1286
rect 4701 1286 4826 1296
rect 4701 1267 4709 1286
rect 4734 1267 4826 1286
rect 4511 1259 4515 1264
rect 4701 1260 4826 1267
rect 4472 1256 4515 1259
rect 4405 1242 4515 1256
rect 2861 1225 2896 1226
rect 2838 1220 2896 1225
rect 2838 1200 2841 1220
rect 2861 1206 2896 1220
rect 2916 1206 2925 1226
rect 2861 1198 2925 1206
rect 2887 1197 2925 1198
rect 2888 1196 2925 1197
rect 2991 1230 3027 1231
rect 3099 1230 3135 1231
rect 2991 1222 3135 1230
rect 2991 1202 2999 1222
rect 3019 1219 3107 1222
rect 3019 1202 3051 1219
rect 3071 1202 3107 1219
rect 3127 1202 3135 1222
rect 2991 1196 3135 1202
rect 3201 1226 3239 1234
rect 3307 1230 3343 1231
rect 3201 1206 3210 1226
rect 3230 1206 3239 1226
rect 3201 1197 3239 1206
rect 3258 1223 3343 1230
rect 3258 1203 3265 1223
rect 3286 1222 3343 1223
rect 3286 1203 3315 1222
rect 3258 1202 3315 1203
rect 3335 1202 3343 1222
rect 3201 1196 3238 1197
rect 3258 1196 3343 1202
rect 3409 1226 3447 1234
rect 3520 1230 3556 1231
rect 3409 1206 3418 1226
rect 3438 1206 3447 1226
rect 3409 1197 3447 1206
rect 3471 1222 3556 1230
rect 3471 1202 3528 1222
rect 3548 1202 3556 1222
rect 3409 1196 3446 1197
rect 3471 1196 3556 1202
rect 3622 1226 3660 1234
rect 3622 1206 3631 1226
rect 3651 1206 3660 1226
rect 3622 1197 3660 1206
rect 4786 1212 4826 1260
rect 5170 1280 5204 1308
rect 5396 1282 5433 1311
rect 5397 1280 5433 1282
rect 5609 1280 5646 1311
rect 5170 1279 5342 1280
rect 5170 1247 5356 1279
rect 5397 1258 5646 1280
rect 5817 1279 5854 1311
rect 6130 1307 6194 1319
rect 6234 1281 6261 1459
rect 8789 1437 8816 1615
rect 8856 1577 8920 1589
rect 9196 1585 9233 1617
rect 9404 1616 9653 1638
rect 9404 1585 9441 1616
rect 9617 1614 9653 1616
rect 9617 1585 9654 1614
rect 8856 1576 8891 1577
rect 8833 1571 8891 1576
rect 8833 1551 8836 1571
rect 8856 1557 8891 1571
rect 8911 1557 8920 1577
rect 8856 1549 8920 1557
rect 8882 1548 8920 1549
rect 8883 1547 8920 1548
rect 8986 1581 9022 1582
rect 9094 1581 9130 1582
rect 8986 1576 9130 1581
rect 8986 1573 9048 1576
rect 8986 1553 8994 1573
rect 9014 1556 9048 1573
rect 9071 1573 9130 1576
rect 9071 1556 9102 1573
rect 9014 1553 9102 1556
rect 9122 1553 9130 1573
rect 8986 1547 9130 1553
rect 9196 1577 9234 1585
rect 9302 1581 9338 1582
rect 9196 1557 9205 1577
rect 9225 1557 9234 1577
rect 9196 1548 9234 1557
rect 9253 1574 9338 1581
rect 9253 1554 9260 1574
rect 9281 1573 9338 1574
rect 9281 1554 9310 1573
rect 9253 1553 9310 1554
rect 9330 1553 9338 1573
rect 9196 1547 9233 1548
rect 9253 1547 9338 1553
rect 9404 1577 9442 1585
rect 9515 1581 9551 1582
rect 9404 1557 9413 1577
rect 9433 1557 9442 1577
rect 9404 1548 9442 1557
rect 9466 1573 9551 1581
rect 9466 1553 9523 1573
rect 9543 1553 9551 1573
rect 9404 1547 9441 1548
rect 9466 1547 9551 1553
rect 9617 1577 9655 1585
rect 9617 1557 9626 1577
rect 9646 1557 9655 1577
rect 9617 1548 9655 1557
rect 9617 1547 9654 1548
rect 9040 1526 9076 1547
rect 9466 1526 9497 1547
rect 8873 1522 8973 1526
rect 8873 1518 8935 1522
rect 8873 1492 8880 1518
rect 8906 1496 8935 1518
rect 8961 1496 8973 1522
rect 8906 1492 8973 1496
rect 8873 1489 8973 1492
rect 9041 1489 9076 1526
rect 9138 1523 9497 1526
rect 9138 1518 9360 1523
rect 9138 1494 9151 1518
rect 9175 1499 9360 1518
rect 9384 1499 9497 1523
rect 9175 1494 9497 1499
rect 9138 1490 9497 1494
rect 9564 1518 9713 1526
rect 9564 1498 9575 1518
rect 9595 1498 9713 1518
rect 9564 1491 9713 1498
rect 9564 1490 9605 1491
rect 8888 1437 8925 1438
rect 8984 1437 9021 1438
rect 9040 1437 9076 1489
rect 9095 1437 9132 1438
rect 8788 1428 8926 1437
rect 8788 1408 8897 1428
rect 8917 1408 8926 1428
rect 8788 1401 8926 1408
rect 8984 1428 9132 1437
rect 8984 1408 8993 1428
rect 9013 1408 9103 1428
rect 9123 1408 9132 1428
rect 8788 1399 8884 1401
rect 8984 1398 9132 1408
rect 9191 1428 9228 1438
rect 9303 1437 9340 1438
rect 9284 1435 9340 1437
rect 9191 1408 9199 1428
rect 9219 1408 9228 1428
rect 9040 1397 9076 1398
rect 6417 1355 6527 1369
rect 6417 1352 6460 1355
rect 6417 1347 6421 1352
rect 6093 1279 6261 1281
rect 5817 1273 6261 1279
rect 5170 1215 5204 1247
rect 3622 1196 3659 1197
rect 3045 1175 3081 1196
rect 3471 1175 3502 1196
rect 4786 1194 4797 1212
rect 4815 1194 4826 1212
rect 4786 1186 4826 1194
rect 5166 1206 5204 1215
rect 5166 1188 5176 1206
rect 5194 1188 5204 1206
rect 4787 1185 4824 1186
rect 5166 1182 5204 1188
rect 5322 1184 5356 1247
rect 5478 1252 5589 1258
rect 5478 1244 5519 1252
rect 5478 1224 5486 1244
rect 5505 1224 5519 1244
rect 5478 1222 5519 1224
rect 5547 1244 5589 1252
rect 5547 1224 5563 1244
rect 5582 1224 5589 1244
rect 5547 1222 5589 1224
rect 5478 1207 5589 1222
rect 5816 1253 6261 1273
rect 5816 1184 5854 1253
rect 6093 1252 6261 1253
rect 6339 1325 6421 1347
rect 6450 1325 6460 1352
rect 6488 1328 6495 1355
rect 6524 1347 6527 1355
rect 8522 1364 8633 1379
rect 8522 1362 8564 1364
rect 6524 1328 6589 1347
rect 6488 1325 6589 1328
rect 6339 1323 6589 1325
rect 6339 1244 6376 1323
rect 6417 1310 6527 1323
rect 6491 1254 6522 1255
rect 6339 1224 6348 1244
rect 6368 1224 6376 1244
rect 6339 1214 6376 1224
rect 6435 1244 6522 1254
rect 6435 1224 6444 1244
rect 6464 1224 6522 1244
rect 6435 1215 6522 1224
rect 6435 1214 6472 1215
rect 5166 1178 5203 1182
rect 2878 1171 2978 1175
rect 2878 1167 2940 1171
rect 2878 1141 2885 1167
rect 2911 1145 2940 1167
rect 2966 1145 2978 1171
rect 2911 1141 2978 1145
rect 2878 1138 2978 1141
rect 3046 1138 3081 1175
rect 3143 1172 3502 1175
rect 3143 1167 3365 1172
rect 3143 1143 3156 1167
rect 3180 1148 3365 1167
rect 3389 1148 3502 1172
rect 3180 1143 3502 1148
rect 3143 1139 3502 1143
rect 3569 1167 3718 1175
rect 5322 1173 5854 1184
rect 3569 1147 3580 1167
rect 3600 1147 3718 1167
rect 5321 1157 5854 1173
rect 6491 1162 6522 1215
rect 6552 1244 6589 1323
rect 6760 1333 7153 1340
rect 6760 1316 6768 1333
rect 6800 1320 7153 1333
rect 7173 1320 7176 1340
rect 8255 1335 8296 1344
rect 6800 1316 7176 1320
rect 6760 1315 7176 1316
rect 7850 1333 8018 1334
rect 8255 1333 8264 1335
rect 6760 1314 7101 1315
rect 6704 1254 6735 1255
rect 6552 1224 6561 1244
rect 6581 1224 6589 1244
rect 6552 1214 6589 1224
rect 6648 1247 6735 1254
rect 6648 1244 6709 1247
rect 6648 1224 6657 1244
rect 6677 1227 6709 1244
rect 6730 1227 6735 1247
rect 6677 1224 6735 1227
rect 6648 1217 6735 1224
rect 6760 1244 6797 1314
rect 7063 1313 7100 1314
rect 7850 1313 8264 1333
rect 8290 1313 8296 1335
rect 8522 1342 8529 1362
rect 8548 1342 8564 1362
rect 8522 1334 8564 1342
rect 8592 1362 8633 1364
rect 8592 1342 8606 1362
rect 8625 1342 8633 1362
rect 8592 1334 8633 1342
rect 8888 1338 8925 1339
rect 9191 1338 9228 1408
rect 9253 1428 9340 1435
rect 9253 1425 9311 1428
rect 9253 1405 9258 1425
rect 9279 1408 9311 1425
rect 9331 1408 9340 1428
rect 9279 1405 9340 1408
rect 9253 1398 9340 1405
rect 9399 1428 9436 1438
rect 9399 1408 9407 1428
rect 9427 1408 9436 1428
rect 9253 1397 9284 1398
rect 8887 1337 9228 1338
rect 8522 1328 8633 1334
rect 8812 1332 9228 1337
rect 7850 1307 8296 1313
rect 7850 1305 8018 1307
rect 6912 1254 6948 1255
rect 6760 1224 6769 1244
rect 6789 1224 6797 1244
rect 6648 1215 6704 1217
rect 6648 1214 6685 1215
rect 6760 1214 6797 1224
rect 6856 1244 7004 1254
rect 7104 1251 7200 1253
rect 6856 1224 6865 1244
rect 6885 1239 6975 1244
rect 6885 1224 6920 1239
rect 6856 1215 6920 1224
rect 6856 1214 6893 1215
rect 6912 1198 6920 1215
rect 6941 1224 6975 1239
rect 6995 1224 7004 1244
rect 6941 1215 7004 1224
rect 7062 1244 7200 1251
rect 7062 1224 7071 1244
rect 7091 1224 7200 1244
rect 7062 1215 7200 1224
rect 6941 1198 6948 1215
rect 6967 1214 7004 1215
rect 7063 1214 7100 1215
rect 6912 1163 6948 1198
rect 6383 1161 6424 1162
rect 5321 1156 5835 1157
rect 3569 1140 3718 1147
rect 6275 1154 6424 1161
rect 4158 1144 4672 1145
rect 3569 1139 3610 1140
rect 2893 1086 2930 1087
rect 2989 1086 3026 1087
rect 3045 1086 3081 1138
rect 3100 1086 3137 1087
rect 2793 1077 2931 1086
rect 2793 1057 2902 1077
rect 2922 1057 2931 1077
rect 2793 1050 2931 1057
rect 2989 1077 3137 1086
rect 2989 1057 2998 1077
rect 3018 1057 3108 1077
rect 3128 1057 3137 1077
rect 2793 1048 2889 1050
rect 2989 1047 3137 1057
rect 3196 1077 3233 1087
rect 3308 1086 3345 1087
rect 3289 1084 3345 1086
rect 3196 1057 3204 1077
rect 3224 1057 3233 1077
rect 3045 1046 3081 1047
rect 1975 994 2143 996
rect 1697 988 2143 994
rect 765 964 1181 969
rect 1360 967 1471 973
rect 765 963 1106 964
rect 709 903 740 904
rect 557 873 566 893
rect 586 873 594 893
rect 557 863 594 873
rect 653 896 740 903
rect 653 893 714 896
rect 653 873 662 893
rect 682 876 714 893
rect 735 876 740 896
rect 682 873 740 876
rect 653 866 740 873
rect 765 893 802 963
rect 1068 962 1105 963
rect 1360 959 1401 967
rect 1360 939 1368 959
rect 1387 939 1401 959
rect 1360 937 1401 939
rect 1429 959 1471 967
rect 1429 939 1445 959
rect 1464 939 1471 959
rect 1697 966 1703 988
rect 1729 968 2143 988
rect 2893 987 2930 988
rect 3196 987 3233 1057
rect 3258 1077 3345 1084
rect 3258 1074 3316 1077
rect 3258 1054 3263 1074
rect 3284 1057 3316 1074
rect 3336 1057 3345 1077
rect 3284 1054 3345 1057
rect 3258 1047 3345 1054
rect 3404 1077 3441 1087
rect 3404 1057 3412 1077
rect 3432 1057 3441 1077
rect 3258 1046 3289 1047
rect 2892 986 3233 987
rect 1729 966 1738 968
rect 1975 967 2143 968
rect 2817 981 3233 986
rect 1697 957 1738 966
rect 2817 961 2820 981
rect 2840 961 3233 981
rect 3404 978 3441 1057
rect 3471 1086 3502 1139
rect 4139 1128 4672 1144
rect 6275 1134 6393 1154
rect 6413 1134 6424 1154
rect 4139 1117 4671 1128
rect 6275 1126 6424 1134
rect 6491 1158 6850 1162
rect 6491 1153 6813 1158
rect 6491 1129 6604 1153
rect 6628 1134 6813 1153
rect 6837 1134 6850 1158
rect 6628 1129 6850 1134
rect 6491 1126 6850 1129
rect 6912 1126 6947 1163
rect 7015 1160 7115 1163
rect 7015 1156 7082 1160
rect 7015 1130 7027 1156
rect 7053 1134 7082 1156
rect 7108 1134 7115 1160
rect 7053 1130 7115 1134
rect 7015 1126 7115 1130
rect 4790 1119 4827 1123
rect 3521 1086 3558 1087
rect 3471 1077 3558 1086
rect 3471 1057 3529 1077
rect 3549 1057 3558 1077
rect 3471 1047 3558 1057
rect 3617 1077 3654 1087
rect 3617 1057 3625 1077
rect 3645 1057 3654 1077
rect 3471 1046 3502 1047
rect 3466 978 3576 991
rect 3617 978 3654 1057
rect 3404 976 3654 978
rect 3404 973 3505 976
rect 3404 954 3469 973
rect 1429 937 1471 939
rect 1360 922 1471 937
rect 3466 946 3469 954
rect 3498 946 3505 973
rect 3533 949 3543 976
rect 3572 954 3654 976
rect 3732 1048 3900 1049
rect 4139 1048 4177 1117
rect 3732 1028 4177 1048
rect 4404 1079 4515 1094
rect 4404 1077 4446 1079
rect 4404 1057 4411 1077
rect 4430 1057 4446 1077
rect 4404 1049 4446 1057
rect 4474 1077 4515 1079
rect 4474 1057 4488 1077
rect 4507 1057 4515 1077
rect 4474 1049 4515 1057
rect 4404 1043 4515 1049
rect 4637 1054 4671 1117
rect 4789 1113 4827 1119
rect 5169 1115 5206 1116
rect 4789 1095 4799 1113
rect 4817 1095 4827 1113
rect 4789 1086 4827 1095
rect 5167 1107 5207 1115
rect 5167 1089 5178 1107
rect 5196 1089 5207 1107
rect 6491 1105 6522 1126
rect 6912 1105 6948 1126
rect 6334 1104 6371 1105
rect 4789 1054 4823 1086
rect 3732 1022 4176 1028
rect 3732 1020 3900 1022
rect 3572 949 3576 954
rect 3533 946 3576 949
rect 3466 932 3576 946
rect 917 903 953 904
rect 765 873 774 893
rect 794 873 802 893
rect 653 864 709 866
rect 653 863 690 864
rect 765 863 802 873
rect 861 893 1009 903
rect 1109 900 1205 902
rect 861 873 870 893
rect 890 873 980 893
rect 1000 873 1009 893
rect 861 864 1009 873
rect 1067 893 1205 900
rect 1067 873 1076 893
rect 1096 873 1205 893
rect 1067 864 1205 873
rect 861 863 898 864
rect 917 812 953 864
rect 972 863 1009 864
rect 1068 863 1105 864
rect 388 810 429 811
rect 280 803 429 810
rect 280 783 398 803
rect 418 783 429 803
rect 280 775 429 783
rect 496 807 855 811
rect 496 802 818 807
rect 496 778 609 802
rect 633 783 818 802
rect 842 783 855 807
rect 633 778 855 783
rect 496 775 855 778
rect 917 775 952 812
rect 1020 809 1120 812
rect 1020 805 1087 809
rect 1020 779 1032 805
rect 1058 783 1087 805
rect 1113 783 1120 809
rect 1058 779 1120 783
rect 1020 775 1120 779
rect 496 754 527 775
rect 917 754 953 775
rect 339 753 376 754
rect 338 744 376 753
rect 338 724 347 744
rect 367 724 376 744
rect 338 716 376 724
rect 442 748 527 754
rect 552 753 589 754
rect 442 728 450 748
rect 470 728 527 748
rect 442 720 527 728
rect 551 744 589 753
rect 551 724 560 744
rect 580 724 589 744
rect 442 719 478 720
rect 551 716 589 724
rect 655 748 740 754
rect 760 753 797 754
rect 655 728 663 748
rect 683 747 740 748
rect 683 728 712 747
rect 655 727 712 728
rect 733 727 740 747
rect 655 720 740 727
rect 759 744 797 753
rect 759 724 768 744
rect 788 724 797 744
rect 655 719 691 720
rect 759 716 797 724
rect 863 748 1007 754
rect 863 728 871 748
rect 891 745 979 748
rect 891 728 922 745
rect 863 725 922 728
rect 945 728 979 745
rect 999 728 1007 748
rect 945 725 1007 728
rect 863 720 1007 725
rect 863 719 899 720
rect 971 719 1007 720
rect 1073 753 1110 754
rect 1073 752 1111 753
rect 1073 744 1137 752
rect 1073 724 1082 744
rect 1102 730 1137 744
rect 1157 730 1160 750
rect 1102 725 1160 730
rect 1102 724 1137 725
rect 339 687 376 716
rect 340 685 376 687
rect 552 685 589 716
rect 340 663 589 685
rect 760 684 797 716
rect 1073 712 1137 724
rect 1177 686 1204 864
rect 3732 842 3759 1020
rect 3799 982 3863 994
rect 4139 990 4176 1022
rect 4347 1021 4596 1043
rect 4637 1022 4823 1054
rect 4651 1021 4823 1022
rect 4347 990 4384 1021
rect 4560 1019 4596 1021
rect 4560 990 4597 1019
rect 4789 993 4823 1021
rect 5167 1041 5207 1089
rect 6333 1095 6371 1104
rect 6333 1075 6342 1095
rect 6362 1075 6371 1095
rect 6333 1067 6371 1075
rect 6437 1099 6522 1105
rect 6547 1104 6584 1105
rect 6437 1079 6445 1099
rect 6465 1079 6522 1099
rect 6437 1071 6522 1079
rect 6546 1095 6584 1104
rect 6546 1075 6555 1095
rect 6575 1075 6584 1095
rect 6437 1070 6473 1071
rect 6546 1067 6584 1075
rect 6650 1099 6735 1105
rect 6755 1104 6792 1105
rect 6650 1079 6658 1099
rect 6678 1098 6735 1099
rect 6678 1079 6707 1098
rect 6650 1078 6707 1079
rect 6728 1078 6735 1098
rect 6650 1071 6735 1078
rect 6754 1095 6792 1104
rect 6754 1075 6763 1095
rect 6783 1075 6792 1095
rect 6650 1070 6686 1071
rect 6754 1067 6792 1075
rect 6858 1099 7002 1105
rect 6858 1079 6866 1099
rect 6886 1079 6974 1099
rect 6994 1079 7002 1099
rect 6858 1071 7002 1079
rect 6858 1070 6894 1071
rect 6966 1070 7002 1071
rect 7068 1104 7105 1105
rect 7068 1103 7106 1104
rect 7068 1095 7132 1103
rect 7068 1075 7077 1095
rect 7097 1081 7132 1095
rect 7152 1081 7155 1101
rect 7097 1076 7155 1081
rect 7097 1075 7132 1076
rect 5478 1045 5588 1059
rect 5478 1042 5521 1045
rect 5167 1034 5292 1041
rect 5478 1037 5482 1042
rect 5167 1015 5259 1034
rect 5284 1015 5292 1034
rect 5167 1005 5292 1015
rect 5400 1015 5482 1037
rect 5511 1015 5521 1042
rect 5549 1018 5556 1045
rect 5585 1037 5588 1045
rect 6334 1038 6371 1067
rect 5585 1018 5650 1037
rect 6335 1036 6371 1038
rect 6547 1036 6584 1067
rect 6755 1040 6792 1067
rect 7068 1063 7132 1075
rect 5549 1015 5650 1018
rect 5400 1013 5650 1015
rect 3799 981 3834 982
rect 3776 976 3834 981
rect 3776 956 3779 976
rect 3799 962 3834 976
rect 3854 962 3863 982
rect 3799 954 3863 962
rect 3825 953 3863 954
rect 3826 952 3863 953
rect 3929 986 3965 987
rect 4037 986 4073 987
rect 3929 979 4073 986
rect 3929 978 3989 979
rect 3929 958 3937 978
rect 3957 959 3989 978
rect 4014 978 4073 979
rect 4014 959 4045 978
rect 3957 958 4045 959
rect 4065 958 4073 978
rect 3929 952 4073 958
rect 4139 982 4177 990
rect 4245 986 4281 987
rect 4139 962 4148 982
rect 4168 962 4177 982
rect 4139 953 4177 962
rect 4196 979 4281 986
rect 4196 959 4203 979
rect 4224 978 4281 979
rect 4224 959 4253 978
rect 4196 958 4253 959
rect 4273 958 4281 978
rect 4139 952 4176 953
rect 4196 952 4281 958
rect 4347 982 4385 990
rect 4458 986 4494 987
rect 4347 962 4356 982
rect 4376 962 4385 982
rect 4347 953 4385 962
rect 4409 978 4494 986
rect 4409 958 4466 978
rect 4486 958 4494 978
rect 4347 952 4384 953
rect 4409 952 4494 958
rect 4560 982 4598 990
rect 4560 962 4569 982
rect 4589 962 4598 982
rect 4560 953 4598 962
rect 4787 983 4824 993
rect 5167 985 5207 1005
rect 4787 965 4797 983
rect 4815 965 4824 983
rect 4787 956 4824 965
rect 5166 976 5207 985
rect 5166 958 5176 976
rect 5194 958 5207 976
rect 4789 955 4823 956
rect 4560 952 4597 953
rect 3983 931 4019 952
rect 4409 931 4440 952
rect 5166 949 5207 958
rect 5166 948 5203 949
rect 5400 934 5437 1013
rect 5478 1000 5588 1013
rect 5552 944 5583 945
rect 3816 927 3916 931
rect 3816 923 3878 927
rect 3816 897 3823 923
rect 3849 901 3878 923
rect 3904 901 3916 927
rect 3849 897 3916 901
rect 3816 894 3916 897
rect 3984 894 4019 931
rect 4081 928 4440 931
rect 4081 923 4303 928
rect 4081 899 4094 923
rect 4118 904 4303 923
rect 4327 904 4440 928
rect 4118 899 4440 904
rect 4081 895 4440 899
rect 4507 923 4656 931
rect 4507 903 4518 923
rect 4538 903 4656 923
rect 5400 914 5409 934
rect 5429 914 5437 934
rect 5400 904 5437 914
rect 5496 934 5583 944
rect 5496 914 5505 934
rect 5525 914 5583 934
rect 5496 905 5583 914
rect 5496 904 5533 905
rect 4507 896 4656 903
rect 4507 895 4548 896
rect 3831 842 3868 843
rect 3927 842 3964 843
rect 3983 842 4019 894
rect 4038 842 4075 843
rect 3731 833 3869 842
rect 3731 813 3840 833
rect 3860 813 3869 833
rect 3731 806 3869 813
rect 3927 833 4075 842
rect 3927 813 3936 833
rect 3956 813 4046 833
rect 4066 813 4075 833
rect 3731 804 3827 806
rect 3927 803 4075 813
rect 4134 833 4171 843
rect 4246 842 4283 843
rect 4227 840 4283 842
rect 4134 813 4142 833
rect 4162 813 4171 833
rect 3983 802 4019 803
rect 3831 743 3868 744
rect 4134 743 4171 813
rect 4196 833 4283 840
rect 4196 830 4254 833
rect 4196 810 4201 830
rect 4222 813 4254 830
rect 4274 813 4283 833
rect 4222 810 4283 813
rect 4196 803 4283 810
rect 4342 833 4379 843
rect 4342 813 4350 833
rect 4370 813 4379 833
rect 4196 802 4227 803
rect 3830 742 4171 743
rect 3755 737 4171 742
rect 3755 717 3758 737
rect 3778 717 4171 737
rect 4342 734 4379 813
rect 4409 842 4440 895
rect 4790 893 4827 894
rect 4789 884 4828 893
rect 4789 866 4799 884
rect 4817 866 4828 884
rect 5169 882 5206 886
rect 4701 849 4748 850
rect 4789 849 4828 866
rect 4701 845 4828 849
rect 4459 842 4496 843
rect 4409 833 4496 842
rect 4409 813 4467 833
rect 4487 813 4496 833
rect 4409 803 4496 813
rect 4555 833 4592 843
rect 4555 813 4563 833
rect 4583 813 4592 833
rect 4409 802 4440 803
rect 4404 734 4514 747
rect 4555 734 4592 813
rect 4701 816 4711 845
rect 4740 816 4828 845
rect 4701 810 4828 816
rect 4701 806 4748 810
rect 4786 796 4828 810
rect 4786 778 4797 796
rect 4815 778 4828 796
rect 4786 773 4828 778
rect 4787 770 4828 773
rect 5166 877 5206 882
rect 5166 859 5178 877
rect 5196 859 5206 877
rect 4787 769 4824 770
rect 4342 732 4592 734
rect 4342 729 4443 732
rect 4342 710 4407 729
rect 4404 702 4407 710
rect 4436 702 4443 729
rect 4471 705 4481 732
rect 4510 710 4592 732
rect 4510 705 4514 710
rect 4471 702 4514 705
rect 4404 688 4514 702
rect 4780 706 4827 707
rect 4780 697 4828 706
rect 1036 684 1204 686
rect 760 681 1204 684
rect 421 657 532 663
rect 421 649 462 657
rect 110 594 149 638
rect 421 629 429 649
rect 448 629 462 649
rect 421 627 462 629
rect 490 651 532 657
rect 758 658 1204 681
rect 4780 679 4799 697
rect 4817 679 4828 697
rect 4780 677 4828 679
rect 4789 658 4828 677
rect 5166 679 5206 859
rect 5552 852 5583 905
rect 5613 934 5650 1013
rect 5821 1010 6214 1030
rect 6234 1010 6237 1030
rect 6335 1014 6584 1036
rect 6753 1035 6794 1040
rect 7172 1037 7199 1215
rect 7850 1127 7877 1305
rect 8255 1302 8296 1307
rect 8465 1306 8714 1328
rect 8812 1312 8815 1332
rect 8835 1312 9228 1332
rect 9399 1329 9436 1408
rect 9466 1437 9497 1490
rect 9843 1483 9883 1663
rect 10140 1746 10180 1926
rect 10526 1919 10557 1972
rect 10587 2001 10624 2080
rect 10795 2077 11188 2097
rect 11208 2077 11211 2097
rect 11309 2081 11558 2103
rect 11727 2102 11768 2107
rect 12146 2104 12173 2282
rect 12824 2194 12851 2372
rect 13229 2369 13270 2374
rect 13439 2373 13688 2395
rect 13786 2379 13789 2399
rect 13809 2379 14202 2399
rect 14373 2396 14410 2475
rect 14440 2504 14471 2557
rect 14817 2550 14857 2730
rect 15195 2732 15234 2789
rect 15844 2787 15882 2789
rect 16415 2786 16564 2793
rect 16415 2766 16533 2786
rect 16553 2766 16564 2786
rect 16415 2758 16564 2766
rect 16631 2790 16990 2794
rect 16631 2785 16953 2790
rect 16631 2761 16744 2785
rect 16768 2766 16953 2785
rect 16977 2766 16990 2790
rect 16768 2761 16990 2766
rect 16631 2758 16990 2761
rect 17052 2758 17087 2795
rect 17155 2792 17255 2795
rect 17155 2788 17222 2792
rect 17155 2762 17167 2788
rect 17193 2766 17222 2788
rect 17248 2766 17255 2792
rect 17193 2762 17255 2766
rect 17155 2758 17255 2762
rect 16631 2737 16662 2758
rect 17052 2737 17088 2758
rect 16474 2736 16511 2737
rect 15195 2730 15243 2732
rect 15195 2712 15206 2730
rect 15224 2712 15243 2730
rect 16473 2727 16511 2736
rect 15195 2703 15243 2712
rect 15196 2702 15243 2703
rect 15509 2707 15619 2721
rect 15509 2704 15552 2707
rect 15509 2699 15513 2704
rect 15431 2677 15513 2699
rect 15542 2677 15552 2704
rect 15580 2680 15587 2707
rect 15616 2699 15619 2707
rect 16473 2707 16482 2727
rect 16502 2707 16511 2727
rect 16473 2699 16511 2707
rect 16577 2731 16662 2737
rect 16687 2736 16724 2737
rect 16577 2711 16585 2731
rect 16605 2711 16662 2731
rect 16577 2703 16662 2711
rect 16686 2727 16724 2736
rect 16686 2707 16695 2727
rect 16715 2707 16724 2727
rect 16577 2702 16613 2703
rect 16686 2699 16724 2707
rect 16790 2731 16875 2737
rect 16895 2736 16932 2737
rect 16790 2711 16798 2731
rect 16818 2730 16875 2731
rect 16818 2711 16847 2730
rect 16790 2710 16847 2711
rect 16868 2710 16875 2730
rect 16790 2703 16875 2710
rect 16894 2727 16932 2736
rect 16894 2707 16903 2727
rect 16923 2707 16932 2727
rect 16790 2702 16826 2703
rect 16894 2699 16932 2707
rect 16998 2731 17142 2737
rect 16998 2711 17006 2731
rect 17026 2711 17114 2731
rect 17134 2711 17142 2731
rect 16998 2703 17142 2711
rect 16998 2702 17034 2703
rect 17106 2702 17142 2703
rect 17208 2736 17245 2737
rect 17208 2735 17246 2736
rect 17208 2727 17272 2735
rect 17208 2707 17217 2727
rect 17237 2713 17272 2727
rect 17292 2713 17295 2733
rect 17237 2708 17295 2713
rect 17237 2707 17272 2708
rect 15616 2680 15681 2699
rect 15580 2677 15681 2680
rect 15431 2675 15681 2677
rect 15199 2639 15236 2640
rect 14817 2532 14827 2550
rect 14845 2532 14857 2550
rect 14817 2527 14857 2532
rect 15195 2636 15236 2639
rect 15195 2631 15237 2636
rect 15195 2613 15208 2631
rect 15226 2613 15237 2631
rect 15195 2599 15237 2613
rect 15275 2599 15322 2603
rect 15195 2593 15322 2599
rect 15195 2564 15283 2593
rect 15312 2564 15322 2593
rect 15431 2596 15468 2675
rect 15509 2662 15619 2675
rect 15583 2606 15614 2607
rect 15431 2576 15440 2596
rect 15460 2576 15468 2596
rect 15431 2566 15468 2576
rect 15527 2596 15614 2606
rect 15527 2576 15536 2596
rect 15556 2576 15614 2596
rect 15527 2567 15614 2576
rect 15527 2566 15564 2567
rect 15195 2560 15322 2564
rect 15195 2543 15234 2560
rect 15275 2559 15322 2560
rect 14817 2523 14854 2527
rect 15195 2525 15206 2543
rect 15224 2525 15234 2543
rect 15195 2516 15234 2525
rect 15196 2515 15233 2516
rect 15583 2514 15614 2567
rect 15644 2596 15681 2675
rect 15852 2672 16245 2692
rect 16265 2672 16268 2692
rect 15852 2667 16268 2672
rect 16474 2670 16511 2699
rect 16475 2668 16511 2670
rect 16687 2668 16724 2699
rect 15852 2666 16193 2667
rect 15796 2606 15827 2607
rect 15644 2576 15653 2596
rect 15673 2576 15681 2596
rect 15644 2566 15681 2576
rect 15740 2599 15827 2606
rect 15740 2596 15801 2599
rect 15740 2576 15749 2596
rect 15769 2579 15801 2596
rect 15822 2579 15827 2599
rect 15769 2576 15827 2579
rect 15740 2569 15827 2576
rect 15852 2596 15889 2666
rect 16155 2665 16192 2666
rect 16475 2646 16724 2668
rect 16895 2667 16932 2699
rect 17208 2695 17272 2707
rect 17312 2677 17339 2847
rect 17770 2814 17797 2990
rect 17837 2954 17901 2966
rect 18177 2962 18214 2994
rect 18385 2993 18634 3015
rect 18917 2995 18954 2996
rect 19220 2995 19257 3065
rect 19282 3085 19369 3092
rect 19282 3082 19340 3085
rect 19282 3062 19287 3082
rect 19308 3065 19340 3082
rect 19360 3065 19369 3085
rect 19308 3062 19369 3065
rect 19282 3055 19369 3062
rect 19428 3085 19465 3095
rect 19428 3065 19436 3085
rect 19456 3065 19465 3085
rect 19282 3054 19313 3055
rect 18916 2994 19257 2995
rect 18385 2962 18422 2993
rect 18598 2991 18634 2993
rect 18598 2962 18635 2991
rect 18841 2989 19257 2994
rect 18841 2969 18844 2989
rect 18864 2969 19257 2989
rect 19428 2986 19465 3065
rect 19495 3094 19526 3147
rect 19876 3145 19913 3146
rect 19875 3136 19914 3145
rect 19875 3118 19885 3136
rect 19903 3118 19914 3136
rect 19787 3101 19834 3102
rect 19875 3101 19914 3118
rect 19787 3097 19914 3101
rect 19545 3094 19582 3095
rect 19495 3085 19582 3094
rect 19495 3065 19553 3085
rect 19573 3065 19582 3085
rect 19495 3055 19582 3065
rect 19641 3085 19678 3095
rect 19641 3065 19649 3085
rect 19669 3065 19678 3085
rect 19495 3054 19526 3055
rect 19490 2986 19600 2999
rect 19641 2986 19678 3065
rect 19787 3068 19797 3097
rect 19826 3068 19914 3097
rect 19787 3062 19914 3068
rect 19787 3058 19834 3062
rect 19872 3048 19914 3062
rect 19872 3030 19883 3048
rect 19901 3030 19914 3048
rect 19872 3025 19914 3030
rect 19873 3022 19914 3025
rect 19873 3021 19910 3022
rect 19428 2984 19678 2986
rect 19428 2981 19529 2984
rect 19428 2962 19493 2981
rect 17837 2953 17872 2954
rect 17814 2948 17872 2953
rect 17814 2928 17817 2948
rect 17837 2934 17872 2948
rect 17892 2934 17901 2954
rect 17837 2926 17901 2934
rect 17863 2925 17901 2926
rect 17864 2924 17901 2925
rect 17967 2958 18003 2959
rect 18075 2958 18111 2959
rect 17967 2951 18111 2958
rect 17967 2950 18025 2951
rect 17967 2930 17975 2950
rect 17995 2932 18025 2950
rect 18054 2950 18111 2951
rect 18054 2932 18083 2950
rect 17995 2930 18083 2932
rect 18103 2930 18111 2950
rect 17967 2924 18111 2930
rect 18177 2954 18215 2962
rect 18283 2958 18319 2959
rect 18177 2934 18186 2954
rect 18206 2934 18215 2954
rect 18177 2925 18215 2934
rect 18234 2951 18319 2958
rect 18234 2931 18241 2951
rect 18262 2950 18319 2951
rect 18262 2931 18291 2950
rect 18234 2930 18291 2931
rect 18311 2930 18319 2950
rect 18177 2924 18214 2925
rect 18234 2924 18319 2930
rect 18385 2954 18423 2962
rect 18496 2958 18532 2959
rect 18385 2934 18394 2954
rect 18414 2934 18423 2954
rect 18385 2925 18423 2934
rect 18447 2950 18532 2958
rect 18447 2930 18504 2950
rect 18524 2930 18532 2950
rect 18385 2924 18422 2925
rect 18447 2924 18532 2930
rect 18598 2954 18636 2962
rect 18598 2934 18607 2954
rect 18627 2934 18636 2954
rect 19490 2954 19493 2962
rect 19522 2954 19529 2981
rect 19557 2957 19567 2984
rect 19596 2962 19678 2984
rect 19596 2957 19600 2962
rect 19557 2954 19600 2957
rect 19490 2940 19600 2954
rect 19866 2958 19913 2959
rect 19866 2949 19914 2958
rect 18598 2925 18636 2934
rect 19866 2931 19885 2949
rect 19903 2931 19914 2949
rect 19866 2929 19914 2931
rect 18598 2924 18635 2925
rect 18021 2903 18057 2924
rect 18447 2903 18478 2924
rect 17854 2899 17954 2903
rect 17854 2895 17916 2899
rect 17854 2869 17861 2895
rect 17887 2873 17916 2895
rect 17942 2873 17954 2899
rect 17887 2869 17954 2873
rect 17854 2866 17954 2869
rect 18022 2866 18057 2903
rect 18119 2900 18478 2903
rect 18119 2895 18341 2900
rect 18119 2871 18132 2895
rect 18156 2876 18341 2895
rect 18365 2876 18478 2900
rect 18156 2871 18478 2876
rect 18119 2867 18478 2871
rect 18545 2895 18694 2903
rect 18545 2875 18556 2895
rect 18576 2875 18694 2895
rect 18545 2868 18694 2875
rect 19227 2872 19265 2874
rect 19875 2872 19914 2929
rect 18545 2867 18586 2868
rect 17869 2814 17906 2815
rect 17965 2814 18002 2815
rect 18021 2814 18057 2866
rect 18076 2814 18113 2815
rect 17769 2805 17907 2814
rect 17769 2785 17878 2805
rect 17898 2785 17907 2805
rect 17769 2778 17907 2785
rect 17965 2805 18113 2814
rect 17965 2785 17974 2805
rect 17994 2785 18084 2805
rect 18104 2785 18113 2805
rect 17769 2776 17865 2778
rect 17965 2775 18113 2785
rect 18172 2805 18209 2815
rect 18284 2814 18321 2815
rect 18265 2812 18321 2814
rect 18172 2785 18180 2805
rect 18200 2785 18209 2805
rect 18021 2774 18057 2775
rect 17869 2715 17906 2716
rect 18172 2715 18209 2785
rect 18234 2805 18321 2812
rect 18234 2802 18292 2805
rect 18234 2782 18239 2802
rect 18260 2785 18292 2802
rect 18312 2785 18321 2805
rect 18260 2782 18321 2785
rect 18234 2775 18321 2782
rect 18380 2805 18417 2815
rect 18380 2785 18388 2805
rect 18408 2785 18417 2805
rect 18234 2774 18265 2775
rect 17868 2714 18209 2715
rect 17793 2709 18209 2714
rect 17793 2689 17796 2709
rect 17816 2689 18209 2709
rect 18380 2706 18417 2785
rect 18447 2814 18478 2867
rect 19227 2839 19913 2872
rect 18497 2814 18534 2815
rect 18447 2805 18534 2814
rect 18447 2785 18505 2805
rect 18525 2785 18534 2805
rect 18447 2775 18534 2785
rect 18593 2805 18630 2815
rect 18593 2785 18601 2805
rect 18621 2785 18630 2805
rect 18447 2774 18478 2775
rect 18442 2706 18552 2719
rect 18593 2706 18630 2785
rect 18380 2704 18630 2706
rect 18380 2701 18481 2704
rect 18380 2682 18445 2701
rect 17260 2669 17339 2677
rect 17171 2667 17339 2669
rect 16895 2660 17339 2667
rect 18442 2674 18445 2682
rect 18474 2674 18481 2701
rect 18509 2677 18519 2704
rect 18548 2682 18630 2704
rect 18819 2751 18987 2752
rect 19227 2751 19265 2839
rect 19526 2837 19573 2839
rect 19873 2815 19913 2839
rect 18819 2728 19265 2751
rect 19491 2782 19602 2796
rect 19491 2780 19533 2782
rect 19491 2760 19498 2780
rect 19517 2760 19533 2780
rect 19491 2752 19533 2760
rect 19561 2780 19602 2782
rect 19561 2760 19575 2780
rect 19594 2760 19602 2780
rect 19874 2771 19913 2815
rect 19561 2752 19602 2760
rect 19491 2746 19602 2752
rect 18819 2725 19263 2728
rect 18819 2723 18987 2725
rect 18548 2677 18552 2682
rect 18509 2674 18552 2677
rect 18442 2660 18552 2674
rect 16556 2640 16667 2646
rect 16895 2641 17265 2660
rect 17171 2640 17265 2641
rect 16556 2632 16597 2640
rect 16556 2612 16564 2632
rect 16583 2612 16597 2632
rect 16556 2610 16597 2612
rect 16625 2632 16667 2640
rect 16625 2612 16641 2632
rect 16660 2612 16667 2632
rect 17260 2631 17265 2640
rect 17313 2640 17339 2660
rect 17313 2631 17330 2640
rect 17260 2622 17330 2631
rect 16625 2610 16667 2612
rect 16004 2606 16040 2607
rect 15852 2576 15861 2596
rect 15881 2576 15889 2596
rect 15740 2567 15796 2569
rect 15740 2566 15777 2567
rect 15852 2566 15889 2576
rect 15948 2596 16096 2606
rect 16196 2603 16292 2605
rect 15948 2576 15957 2596
rect 15977 2576 16067 2596
rect 16087 2576 16096 2596
rect 15948 2567 16096 2576
rect 16154 2596 16292 2603
rect 16154 2576 16163 2596
rect 16183 2576 16292 2596
rect 16556 2595 16667 2610
rect 16154 2567 16292 2576
rect 15948 2566 15985 2567
rect 16004 2515 16040 2567
rect 16059 2566 16096 2567
rect 16155 2566 16192 2567
rect 15475 2513 15516 2514
rect 15367 2506 15516 2513
rect 14490 2504 14527 2505
rect 14440 2495 14527 2504
rect 14440 2475 14498 2495
rect 14518 2475 14527 2495
rect 14440 2465 14527 2475
rect 14586 2495 14623 2505
rect 14586 2475 14594 2495
rect 14614 2475 14623 2495
rect 15367 2486 15485 2506
rect 15505 2486 15516 2506
rect 15367 2478 15516 2486
rect 15583 2510 15942 2514
rect 15583 2505 15905 2510
rect 15583 2481 15696 2505
rect 15720 2486 15905 2505
rect 15929 2486 15942 2510
rect 15720 2481 15942 2486
rect 15583 2478 15942 2481
rect 16004 2478 16039 2515
rect 16107 2512 16207 2515
rect 16107 2508 16174 2512
rect 16107 2482 16119 2508
rect 16145 2486 16174 2508
rect 16200 2486 16207 2512
rect 16145 2482 16207 2486
rect 16107 2478 16207 2482
rect 14440 2464 14471 2465
rect 14435 2396 14545 2409
rect 14586 2396 14623 2475
rect 14820 2460 14857 2461
rect 14816 2451 14857 2460
rect 15583 2457 15614 2478
rect 16004 2457 16040 2478
rect 15426 2456 15463 2457
rect 15200 2453 15234 2454
rect 14816 2433 14829 2451
rect 14847 2433 14857 2451
rect 14816 2424 14857 2433
rect 15199 2444 15236 2453
rect 15199 2426 15208 2444
rect 15226 2426 15236 2444
rect 14816 2404 14856 2424
rect 15199 2416 15236 2426
rect 15425 2447 15463 2456
rect 15425 2427 15434 2447
rect 15454 2427 15463 2447
rect 15425 2419 15463 2427
rect 15529 2451 15614 2457
rect 15639 2456 15676 2457
rect 15529 2431 15537 2451
rect 15557 2431 15614 2451
rect 15529 2423 15614 2431
rect 15638 2447 15676 2456
rect 15638 2427 15647 2447
rect 15667 2427 15676 2447
rect 15529 2422 15565 2423
rect 15638 2419 15676 2427
rect 15742 2451 15827 2457
rect 15847 2456 15884 2457
rect 15742 2431 15750 2451
rect 15770 2450 15827 2451
rect 15770 2431 15799 2450
rect 15742 2430 15799 2431
rect 15820 2430 15827 2450
rect 15742 2423 15827 2430
rect 15846 2447 15884 2456
rect 15846 2427 15855 2447
rect 15875 2427 15884 2447
rect 15742 2422 15778 2423
rect 15846 2419 15884 2427
rect 15950 2451 16094 2457
rect 15950 2431 15958 2451
rect 15978 2450 16066 2451
rect 15978 2431 16009 2450
rect 15950 2430 16009 2431
rect 16034 2431 16066 2450
rect 16086 2431 16094 2451
rect 16034 2430 16094 2431
rect 15950 2423 16094 2430
rect 15950 2422 15986 2423
rect 16058 2422 16094 2423
rect 16160 2456 16197 2457
rect 16160 2455 16198 2456
rect 16160 2447 16224 2455
rect 16160 2427 16169 2447
rect 16189 2433 16224 2447
rect 16244 2433 16247 2453
rect 16189 2428 16247 2433
rect 16189 2427 16224 2428
rect 14373 2394 14623 2396
rect 14373 2391 14474 2394
rect 12891 2334 12955 2346
rect 13231 2342 13268 2369
rect 13439 2342 13476 2373
rect 13652 2371 13688 2373
rect 14373 2372 14438 2391
rect 13652 2342 13689 2371
rect 14435 2364 14438 2372
rect 14467 2364 14474 2391
rect 14502 2367 14512 2394
rect 14541 2372 14623 2394
rect 14731 2394 14856 2404
rect 14731 2375 14739 2394
rect 14764 2375 14856 2394
rect 14541 2367 14545 2372
rect 14731 2368 14856 2375
rect 14502 2364 14545 2367
rect 14435 2350 14545 2364
rect 12891 2333 12926 2334
rect 12868 2328 12926 2333
rect 12868 2308 12871 2328
rect 12891 2314 12926 2328
rect 12946 2314 12955 2334
rect 12891 2306 12955 2314
rect 12917 2305 12955 2306
rect 12918 2304 12955 2305
rect 13021 2338 13057 2339
rect 13129 2338 13165 2339
rect 13021 2330 13165 2338
rect 13021 2310 13029 2330
rect 13049 2310 13137 2330
rect 13157 2310 13165 2330
rect 13021 2304 13165 2310
rect 13231 2334 13269 2342
rect 13337 2338 13373 2339
rect 13231 2314 13240 2334
rect 13260 2314 13269 2334
rect 13231 2305 13269 2314
rect 13288 2331 13373 2338
rect 13288 2311 13295 2331
rect 13316 2330 13373 2331
rect 13316 2311 13345 2330
rect 13288 2310 13345 2311
rect 13365 2310 13373 2330
rect 13231 2304 13268 2305
rect 13288 2304 13373 2310
rect 13439 2334 13477 2342
rect 13550 2338 13586 2339
rect 13439 2314 13448 2334
rect 13468 2314 13477 2334
rect 13439 2305 13477 2314
rect 13501 2330 13586 2338
rect 13501 2310 13558 2330
rect 13578 2310 13586 2330
rect 13439 2304 13476 2305
rect 13501 2304 13586 2310
rect 13652 2334 13690 2342
rect 13652 2314 13661 2334
rect 13681 2314 13690 2334
rect 13652 2305 13690 2314
rect 14816 2320 14856 2368
rect 15200 2388 15234 2416
rect 15426 2390 15463 2419
rect 15427 2388 15463 2390
rect 15639 2388 15676 2419
rect 15200 2387 15372 2388
rect 15200 2355 15386 2387
rect 15427 2366 15676 2388
rect 15847 2387 15884 2419
rect 16160 2415 16224 2427
rect 16264 2389 16291 2567
rect 18819 2545 18846 2723
rect 18886 2685 18950 2697
rect 19226 2693 19263 2725
rect 19434 2724 19683 2746
rect 19434 2693 19471 2724
rect 19647 2722 19683 2724
rect 19647 2693 19684 2722
rect 18886 2684 18921 2685
rect 18863 2679 18921 2684
rect 18863 2659 18866 2679
rect 18886 2665 18921 2679
rect 18941 2665 18950 2685
rect 18886 2657 18950 2665
rect 18912 2656 18950 2657
rect 18913 2655 18950 2656
rect 19016 2689 19052 2690
rect 19124 2689 19160 2690
rect 19016 2684 19160 2689
rect 19016 2681 19078 2684
rect 19016 2661 19024 2681
rect 19044 2664 19078 2681
rect 19101 2681 19160 2684
rect 19101 2664 19132 2681
rect 19044 2661 19132 2664
rect 19152 2661 19160 2681
rect 19016 2655 19160 2661
rect 19226 2685 19264 2693
rect 19332 2689 19368 2690
rect 19226 2665 19235 2685
rect 19255 2665 19264 2685
rect 19226 2656 19264 2665
rect 19283 2682 19368 2689
rect 19283 2662 19290 2682
rect 19311 2681 19368 2682
rect 19311 2662 19340 2681
rect 19283 2661 19340 2662
rect 19360 2661 19368 2681
rect 19226 2655 19263 2656
rect 19283 2655 19368 2661
rect 19434 2685 19472 2693
rect 19545 2689 19581 2690
rect 19434 2665 19443 2685
rect 19463 2665 19472 2685
rect 19434 2656 19472 2665
rect 19496 2681 19581 2689
rect 19496 2661 19553 2681
rect 19573 2661 19581 2681
rect 19434 2655 19471 2656
rect 19496 2655 19581 2661
rect 19647 2685 19685 2693
rect 19647 2665 19656 2685
rect 19676 2665 19685 2685
rect 19647 2656 19685 2665
rect 19647 2655 19684 2656
rect 19070 2634 19106 2655
rect 19496 2634 19527 2655
rect 18903 2630 19003 2634
rect 18903 2626 18965 2630
rect 18903 2600 18910 2626
rect 18936 2604 18965 2626
rect 18991 2604 19003 2630
rect 18936 2600 19003 2604
rect 18903 2597 19003 2600
rect 19071 2597 19106 2634
rect 19168 2631 19527 2634
rect 19168 2626 19390 2631
rect 19168 2602 19181 2626
rect 19205 2607 19390 2626
rect 19414 2607 19527 2631
rect 19205 2602 19527 2607
rect 19168 2598 19527 2602
rect 19594 2626 19743 2634
rect 19594 2606 19605 2626
rect 19625 2606 19743 2626
rect 19594 2599 19743 2606
rect 19594 2598 19635 2599
rect 18918 2545 18955 2546
rect 19014 2545 19051 2546
rect 19070 2545 19106 2597
rect 19125 2545 19162 2546
rect 18818 2536 18956 2545
rect 18818 2516 18927 2536
rect 18947 2516 18956 2536
rect 18818 2509 18956 2516
rect 19014 2536 19162 2545
rect 19014 2516 19023 2536
rect 19043 2516 19133 2536
rect 19153 2516 19162 2536
rect 18818 2507 18914 2509
rect 19014 2506 19162 2516
rect 19221 2536 19258 2546
rect 19333 2545 19370 2546
rect 19314 2543 19370 2545
rect 19221 2516 19229 2536
rect 19249 2516 19258 2536
rect 19070 2505 19106 2506
rect 16447 2463 16557 2477
rect 16447 2460 16490 2463
rect 16447 2455 16451 2460
rect 16123 2387 16291 2389
rect 15847 2381 16291 2387
rect 15200 2323 15234 2355
rect 13652 2304 13689 2305
rect 13075 2283 13111 2304
rect 13501 2283 13532 2304
rect 14816 2302 14827 2320
rect 14845 2302 14856 2320
rect 14816 2294 14856 2302
rect 15196 2314 15234 2323
rect 15196 2296 15206 2314
rect 15224 2296 15234 2314
rect 14817 2293 14854 2294
rect 15196 2290 15234 2296
rect 15352 2292 15386 2355
rect 15508 2360 15619 2366
rect 15508 2352 15549 2360
rect 15508 2332 15516 2352
rect 15535 2332 15549 2352
rect 15508 2330 15549 2332
rect 15577 2352 15619 2360
rect 15577 2332 15593 2352
rect 15612 2332 15619 2352
rect 15577 2330 15619 2332
rect 15508 2315 15619 2330
rect 15846 2361 16291 2381
rect 15846 2292 15884 2361
rect 16123 2360 16291 2361
rect 16369 2433 16451 2455
rect 16480 2433 16490 2460
rect 16518 2436 16525 2463
rect 16554 2455 16557 2463
rect 18552 2472 18663 2487
rect 18552 2470 18594 2472
rect 16554 2436 16619 2455
rect 16518 2433 16619 2436
rect 16369 2431 16619 2433
rect 16369 2352 16406 2431
rect 16447 2418 16557 2431
rect 16521 2362 16552 2363
rect 16369 2332 16378 2352
rect 16398 2332 16406 2352
rect 16369 2322 16406 2332
rect 16465 2352 16552 2362
rect 16465 2332 16474 2352
rect 16494 2332 16552 2352
rect 16465 2323 16552 2332
rect 16465 2322 16502 2323
rect 15196 2286 15233 2290
rect 12908 2279 13008 2283
rect 12908 2275 12970 2279
rect 12908 2249 12915 2275
rect 12941 2253 12970 2275
rect 12996 2253 13008 2279
rect 12941 2249 13008 2253
rect 12908 2246 13008 2249
rect 13076 2246 13111 2283
rect 13173 2280 13532 2283
rect 13173 2275 13395 2280
rect 13173 2251 13186 2275
rect 13210 2256 13395 2275
rect 13419 2256 13532 2280
rect 13210 2251 13532 2256
rect 13173 2247 13532 2251
rect 13599 2275 13748 2283
rect 15352 2281 15884 2292
rect 13599 2255 13610 2275
rect 13630 2255 13748 2275
rect 15351 2265 15884 2281
rect 16521 2270 16552 2323
rect 16582 2352 16619 2431
rect 16790 2428 17183 2448
rect 17203 2428 17206 2448
rect 18285 2443 18326 2452
rect 16790 2423 17206 2428
rect 17880 2441 18048 2442
rect 18285 2441 18294 2443
rect 16790 2422 17131 2423
rect 16734 2362 16765 2363
rect 16582 2332 16591 2352
rect 16611 2332 16619 2352
rect 16582 2322 16619 2332
rect 16678 2355 16765 2362
rect 16678 2352 16739 2355
rect 16678 2332 16687 2352
rect 16707 2335 16739 2352
rect 16760 2335 16765 2355
rect 16707 2332 16765 2335
rect 16678 2325 16765 2332
rect 16790 2352 16827 2422
rect 17093 2421 17130 2422
rect 17880 2421 18294 2441
rect 18320 2421 18326 2443
rect 18552 2450 18559 2470
rect 18578 2450 18594 2470
rect 18552 2442 18594 2450
rect 18622 2470 18663 2472
rect 18622 2450 18636 2470
rect 18655 2450 18663 2470
rect 18622 2442 18663 2450
rect 18918 2446 18955 2447
rect 19221 2446 19258 2516
rect 19283 2536 19370 2543
rect 19283 2533 19341 2536
rect 19283 2513 19288 2533
rect 19309 2516 19341 2533
rect 19361 2516 19370 2536
rect 19309 2513 19370 2516
rect 19283 2506 19370 2513
rect 19429 2536 19466 2546
rect 19429 2516 19437 2536
rect 19457 2516 19466 2536
rect 19283 2505 19314 2506
rect 18917 2445 19258 2446
rect 18552 2436 18663 2442
rect 18842 2440 19258 2445
rect 17880 2415 18326 2421
rect 17880 2413 18048 2415
rect 16942 2362 16978 2363
rect 16790 2332 16799 2352
rect 16819 2332 16827 2352
rect 16678 2323 16734 2325
rect 16678 2322 16715 2323
rect 16790 2322 16827 2332
rect 16886 2352 17034 2362
rect 17134 2359 17230 2361
rect 16886 2332 16895 2352
rect 16915 2332 17005 2352
rect 17025 2332 17034 2352
rect 16886 2323 17034 2332
rect 17092 2352 17230 2359
rect 17092 2332 17101 2352
rect 17121 2332 17230 2352
rect 17092 2323 17230 2332
rect 16886 2322 16923 2323
rect 16942 2271 16978 2323
rect 16997 2322 17034 2323
rect 17093 2322 17130 2323
rect 16413 2269 16454 2270
rect 15351 2264 15865 2265
rect 13599 2248 13748 2255
rect 16305 2262 16454 2269
rect 14188 2252 14702 2253
rect 13599 2247 13640 2248
rect 13075 2211 13111 2246
rect 12923 2194 12960 2195
rect 13019 2194 13056 2195
rect 13075 2194 13082 2211
rect 12823 2185 12961 2194
rect 12823 2165 12932 2185
rect 12952 2165 12961 2185
rect 12823 2158 12961 2165
rect 13019 2185 13082 2194
rect 13019 2165 13028 2185
rect 13048 2170 13082 2185
rect 13103 2194 13111 2211
rect 13130 2194 13167 2195
rect 13103 2185 13167 2194
rect 13103 2170 13138 2185
rect 13048 2165 13138 2170
rect 13158 2165 13167 2185
rect 12823 2156 12919 2158
rect 13019 2155 13167 2165
rect 13226 2185 13263 2195
rect 13338 2194 13375 2195
rect 13319 2192 13375 2194
rect 13226 2165 13234 2185
rect 13254 2165 13263 2185
rect 13075 2154 13111 2155
rect 12005 2102 12173 2104
rect 11727 2096 12173 2102
rect 10795 2072 11211 2077
rect 11390 2075 11501 2081
rect 10795 2071 11136 2072
rect 10739 2011 10770 2012
rect 10587 1981 10596 2001
rect 10616 1981 10624 2001
rect 10587 1971 10624 1981
rect 10683 2004 10770 2011
rect 10683 2001 10744 2004
rect 10683 1981 10692 2001
rect 10712 1984 10744 2001
rect 10765 1984 10770 2004
rect 10712 1981 10770 1984
rect 10683 1974 10770 1981
rect 10795 2001 10832 2071
rect 11098 2070 11135 2071
rect 11390 2067 11431 2075
rect 11390 2047 11398 2067
rect 11417 2047 11431 2067
rect 11390 2045 11431 2047
rect 11459 2067 11501 2075
rect 11459 2047 11475 2067
rect 11494 2047 11501 2067
rect 11727 2074 11733 2096
rect 11759 2076 12173 2096
rect 12923 2095 12960 2096
rect 13226 2095 13263 2165
rect 13288 2185 13375 2192
rect 13288 2182 13346 2185
rect 13288 2162 13293 2182
rect 13314 2165 13346 2182
rect 13366 2165 13375 2185
rect 13314 2162 13375 2165
rect 13288 2155 13375 2162
rect 13434 2185 13471 2195
rect 13434 2165 13442 2185
rect 13462 2165 13471 2185
rect 13288 2154 13319 2155
rect 12922 2094 13263 2095
rect 11759 2074 11768 2076
rect 12005 2075 12173 2076
rect 12847 2093 13263 2094
rect 12847 2089 13223 2093
rect 11727 2065 11768 2074
rect 12847 2069 12850 2089
rect 12870 2076 13223 2089
rect 13255 2076 13263 2093
rect 12870 2069 13263 2076
rect 13434 2086 13471 2165
rect 13501 2194 13532 2247
rect 14169 2236 14702 2252
rect 16305 2242 16423 2262
rect 16443 2242 16454 2262
rect 14169 2225 14701 2236
rect 16305 2234 16454 2242
rect 16521 2266 16880 2270
rect 16521 2261 16843 2266
rect 16521 2237 16634 2261
rect 16658 2242 16843 2261
rect 16867 2242 16880 2266
rect 16658 2237 16880 2242
rect 16521 2234 16880 2237
rect 16942 2234 16977 2271
rect 17045 2268 17145 2271
rect 17045 2264 17112 2268
rect 17045 2238 17057 2264
rect 17083 2242 17112 2264
rect 17138 2242 17145 2268
rect 17083 2238 17145 2242
rect 17045 2234 17145 2238
rect 14820 2227 14857 2231
rect 13551 2194 13588 2195
rect 13501 2185 13588 2194
rect 13501 2165 13559 2185
rect 13579 2165 13588 2185
rect 13501 2155 13588 2165
rect 13647 2185 13684 2195
rect 13647 2165 13655 2185
rect 13675 2165 13684 2185
rect 13501 2154 13532 2155
rect 13496 2086 13606 2099
rect 13647 2086 13684 2165
rect 13434 2084 13684 2086
rect 13434 2081 13535 2084
rect 13434 2062 13499 2081
rect 11459 2045 11501 2047
rect 11390 2030 11501 2045
rect 13496 2054 13499 2062
rect 13528 2054 13535 2081
rect 13563 2057 13573 2084
rect 13602 2062 13684 2084
rect 13762 2156 13930 2157
rect 14169 2156 14207 2225
rect 13762 2136 14207 2156
rect 14434 2187 14545 2202
rect 14434 2185 14476 2187
rect 14434 2165 14441 2185
rect 14460 2165 14476 2185
rect 14434 2157 14476 2165
rect 14504 2185 14545 2187
rect 14504 2165 14518 2185
rect 14537 2165 14545 2185
rect 14504 2157 14545 2165
rect 14434 2151 14545 2157
rect 14667 2162 14701 2225
rect 14819 2221 14857 2227
rect 15199 2223 15236 2224
rect 14819 2203 14829 2221
rect 14847 2203 14857 2221
rect 14819 2194 14857 2203
rect 15197 2215 15237 2223
rect 15197 2197 15208 2215
rect 15226 2197 15237 2215
rect 16521 2213 16552 2234
rect 16942 2213 16978 2234
rect 16364 2212 16401 2213
rect 14819 2162 14853 2194
rect 13762 2130 14206 2136
rect 13762 2128 13930 2130
rect 13602 2057 13606 2062
rect 13563 2054 13606 2057
rect 13496 2040 13606 2054
rect 10947 2011 10983 2012
rect 10795 1981 10804 2001
rect 10824 1981 10832 2001
rect 10683 1972 10739 1974
rect 10683 1971 10720 1972
rect 10795 1971 10832 1981
rect 10891 2001 11039 2011
rect 11139 2008 11235 2010
rect 10891 1981 10900 2001
rect 10920 1981 11010 2001
rect 11030 1981 11039 2001
rect 10891 1972 11039 1981
rect 11097 2001 11235 2008
rect 11097 1981 11106 2001
rect 11126 1981 11235 2001
rect 11097 1972 11235 1981
rect 10891 1971 10928 1972
rect 10947 1920 10983 1972
rect 11002 1971 11039 1972
rect 11098 1971 11135 1972
rect 10418 1918 10459 1919
rect 10310 1911 10459 1918
rect 10310 1891 10428 1911
rect 10448 1891 10459 1911
rect 10310 1883 10459 1891
rect 10526 1915 10885 1919
rect 10526 1910 10848 1915
rect 10526 1886 10639 1910
rect 10663 1891 10848 1910
rect 10872 1891 10885 1915
rect 10663 1886 10885 1891
rect 10526 1883 10885 1886
rect 10947 1883 10982 1920
rect 11050 1917 11150 1920
rect 11050 1913 11117 1917
rect 11050 1887 11062 1913
rect 11088 1891 11117 1913
rect 11143 1891 11150 1917
rect 11088 1887 11150 1891
rect 11050 1883 11150 1887
rect 10526 1862 10557 1883
rect 10947 1862 10983 1883
rect 10369 1861 10406 1862
rect 10368 1852 10406 1861
rect 10368 1832 10377 1852
rect 10397 1832 10406 1852
rect 10368 1824 10406 1832
rect 10472 1856 10557 1862
rect 10582 1861 10619 1862
rect 10472 1836 10480 1856
rect 10500 1836 10557 1856
rect 10472 1828 10557 1836
rect 10581 1852 10619 1861
rect 10581 1832 10590 1852
rect 10610 1832 10619 1852
rect 10472 1827 10508 1828
rect 10581 1824 10619 1832
rect 10685 1856 10770 1862
rect 10790 1861 10827 1862
rect 10685 1836 10693 1856
rect 10713 1855 10770 1856
rect 10713 1836 10742 1855
rect 10685 1835 10742 1836
rect 10763 1835 10770 1855
rect 10685 1828 10770 1835
rect 10789 1852 10827 1861
rect 10789 1832 10798 1852
rect 10818 1832 10827 1852
rect 10685 1827 10721 1828
rect 10789 1824 10827 1832
rect 10893 1856 11037 1862
rect 10893 1836 10901 1856
rect 10921 1853 11009 1856
rect 10921 1836 10952 1853
rect 10893 1833 10952 1836
rect 10975 1836 11009 1853
rect 11029 1836 11037 1856
rect 10975 1833 11037 1836
rect 10893 1828 11037 1833
rect 10893 1827 10929 1828
rect 11001 1827 11037 1828
rect 11103 1861 11140 1862
rect 11103 1860 11141 1861
rect 11103 1852 11167 1860
rect 11103 1832 11112 1852
rect 11132 1838 11167 1852
rect 11187 1838 11190 1858
rect 11132 1833 11190 1838
rect 11132 1832 11167 1833
rect 10369 1795 10406 1824
rect 10370 1793 10406 1795
rect 10582 1793 10619 1824
rect 10370 1771 10619 1793
rect 10790 1792 10827 1824
rect 11103 1820 11167 1832
rect 11207 1794 11234 1972
rect 13762 1950 13789 2128
rect 13829 2090 13893 2102
rect 14169 2098 14206 2130
rect 14377 2129 14626 2151
rect 14667 2130 14853 2162
rect 14681 2129 14853 2130
rect 14377 2098 14414 2129
rect 14590 2127 14626 2129
rect 14590 2098 14627 2127
rect 14819 2101 14853 2129
rect 15197 2149 15237 2197
rect 16363 2203 16401 2212
rect 16363 2183 16372 2203
rect 16392 2183 16401 2203
rect 16363 2175 16401 2183
rect 16467 2207 16552 2213
rect 16577 2212 16614 2213
rect 16467 2187 16475 2207
rect 16495 2187 16552 2207
rect 16467 2179 16552 2187
rect 16576 2203 16614 2212
rect 16576 2183 16585 2203
rect 16605 2183 16614 2203
rect 16467 2178 16503 2179
rect 16576 2175 16614 2183
rect 16680 2207 16765 2213
rect 16785 2212 16822 2213
rect 16680 2187 16688 2207
rect 16708 2206 16765 2207
rect 16708 2187 16737 2206
rect 16680 2186 16737 2187
rect 16758 2186 16765 2206
rect 16680 2179 16765 2186
rect 16784 2203 16822 2212
rect 16784 2183 16793 2203
rect 16813 2183 16822 2203
rect 16680 2178 16716 2179
rect 16784 2175 16822 2183
rect 16888 2207 17032 2213
rect 16888 2187 16896 2207
rect 16916 2190 16952 2207
rect 16972 2190 17004 2207
rect 16916 2187 17004 2190
rect 17024 2187 17032 2207
rect 16888 2179 17032 2187
rect 16888 2178 16924 2179
rect 16996 2178 17032 2179
rect 17098 2212 17135 2213
rect 17098 2211 17136 2212
rect 17098 2203 17162 2211
rect 17098 2183 17107 2203
rect 17127 2189 17162 2203
rect 17182 2189 17185 2209
rect 17127 2184 17185 2189
rect 17127 2183 17162 2184
rect 15508 2153 15618 2167
rect 15508 2150 15551 2153
rect 15197 2142 15322 2149
rect 15508 2145 15512 2150
rect 15197 2123 15289 2142
rect 15314 2123 15322 2142
rect 15197 2113 15322 2123
rect 15430 2123 15512 2145
rect 15541 2123 15551 2150
rect 15579 2126 15586 2153
rect 15615 2145 15618 2153
rect 16364 2146 16401 2175
rect 15615 2126 15680 2145
rect 16365 2144 16401 2146
rect 16577 2144 16614 2175
rect 16785 2148 16822 2175
rect 17098 2171 17162 2183
rect 15579 2123 15680 2126
rect 15430 2121 15680 2123
rect 13829 2089 13864 2090
rect 13806 2084 13864 2089
rect 13806 2064 13809 2084
rect 13829 2070 13864 2084
rect 13884 2070 13893 2090
rect 13829 2062 13893 2070
rect 13855 2061 13893 2062
rect 13856 2060 13893 2061
rect 13959 2094 13995 2095
rect 14067 2094 14103 2095
rect 13959 2087 14103 2094
rect 13959 2086 14019 2087
rect 13959 2066 13967 2086
rect 13987 2067 14019 2086
rect 14044 2086 14103 2087
rect 14044 2067 14075 2086
rect 13987 2066 14075 2067
rect 14095 2066 14103 2086
rect 13959 2060 14103 2066
rect 14169 2090 14207 2098
rect 14275 2094 14311 2095
rect 14169 2070 14178 2090
rect 14198 2070 14207 2090
rect 14169 2061 14207 2070
rect 14226 2087 14311 2094
rect 14226 2067 14233 2087
rect 14254 2086 14311 2087
rect 14254 2067 14283 2086
rect 14226 2066 14283 2067
rect 14303 2066 14311 2086
rect 14169 2060 14206 2061
rect 14226 2060 14311 2066
rect 14377 2090 14415 2098
rect 14488 2094 14524 2095
rect 14377 2070 14386 2090
rect 14406 2070 14415 2090
rect 14377 2061 14415 2070
rect 14439 2086 14524 2094
rect 14439 2066 14496 2086
rect 14516 2066 14524 2086
rect 14377 2060 14414 2061
rect 14439 2060 14524 2066
rect 14590 2090 14628 2098
rect 14590 2070 14599 2090
rect 14619 2070 14628 2090
rect 14590 2061 14628 2070
rect 14817 2091 14854 2101
rect 15197 2093 15237 2113
rect 14817 2073 14827 2091
rect 14845 2073 14854 2091
rect 14817 2064 14854 2073
rect 15196 2084 15237 2093
rect 15196 2066 15206 2084
rect 15224 2066 15237 2084
rect 14819 2063 14853 2064
rect 14590 2060 14627 2061
rect 14013 2039 14049 2060
rect 14439 2039 14470 2060
rect 15196 2057 15237 2066
rect 15196 2056 15233 2057
rect 15430 2042 15467 2121
rect 15508 2108 15618 2121
rect 15582 2052 15613 2053
rect 13846 2035 13946 2039
rect 13846 2031 13908 2035
rect 13846 2005 13853 2031
rect 13879 2009 13908 2031
rect 13934 2009 13946 2035
rect 13879 2005 13946 2009
rect 13846 2002 13946 2005
rect 14014 2002 14049 2039
rect 14111 2036 14470 2039
rect 14111 2031 14333 2036
rect 14111 2007 14124 2031
rect 14148 2012 14333 2031
rect 14357 2012 14470 2036
rect 14148 2007 14470 2012
rect 14111 2003 14470 2007
rect 14537 2031 14686 2039
rect 14537 2011 14548 2031
rect 14568 2011 14686 2031
rect 15430 2022 15439 2042
rect 15459 2022 15467 2042
rect 15430 2012 15467 2022
rect 15526 2042 15613 2052
rect 15526 2022 15535 2042
rect 15555 2022 15613 2042
rect 15526 2013 15613 2022
rect 15526 2012 15563 2013
rect 14537 2004 14686 2011
rect 14537 2003 14578 2004
rect 13861 1950 13898 1951
rect 13957 1950 13994 1951
rect 14013 1950 14049 2002
rect 14068 1950 14105 1951
rect 13761 1941 13899 1950
rect 13356 1920 13467 1935
rect 13356 1918 13398 1920
rect 13026 1897 13131 1899
rect 12684 1889 12852 1890
rect 13026 1889 13075 1897
rect 12684 1870 13075 1889
rect 13106 1870 13131 1897
rect 13356 1898 13363 1918
rect 13382 1898 13398 1918
rect 13356 1890 13398 1898
rect 13426 1918 13467 1920
rect 13426 1898 13440 1918
rect 13459 1898 13467 1918
rect 13761 1921 13870 1941
rect 13890 1921 13899 1941
rect 13761 1914 13899 1921
rect 13957 1941 14105 1950
rect 13957 1921 13966 1941
rect 13986 1921 14076 1941
rect 14096 1921 14105 1941
rect 13761 1912 13857 1914
rect 13957 1911 14105 1921
rect 14164 1941 14201 1951
rect 14276 1950 14313 1951
rect 14257 1948 14313 1950
rect 14164 1921 14172 1941
rect 14192 1921 14201 1941
rect 14013 1910 14049 1911
rect 13426 1890 13467 1898
rect 13356 1884 13467 1890
rect 12684 1863 13131 1870
rect 12684 1861 12852 1863
rect 11532 1830 11642 1844
rect 11532 1827 11575 1830
rect 11532 1822 11536 1827
rect 11066 1792 11234 1794
rect 10790 1789 11234 1792
rect 10451 1765 10562 1771
rect 10451 1757 10492 1765
rect 10140 1702 10179 1746
rect 10451 1737 10459 1757
rect 10478 1737 10492 1757
rect 10451 1735 10492 1737
rect 10520 1757 10562 1765
rect 10520 1737 10536 1757
rect 10555 1737 10562 1757
rect 10520 1735 10562 1737
rect 10451 1720 10562 1735
rect 10788 1766 11234 1789
rect 10140 1678 10180 1702
rect 10480 1678 10527 1680
rect 10788 1678 10826 1766
rect 11066 1765 11234 1766
rect 11454 1800 11536 1822
rect 11565 1800 11575 1827
rect 11603 1803 11610 1830
rect 11639 1822 11642 1830
rect 11639 1803 11704 1822
rect 11603 1800 11704 1803
rect 11454 1798 11704 1800
rect 11454 1719 11491 1798
rect 11532 1785 11642 1798
rect 11606 1729 11637 1730
rect 11454 1699 11463 1719
rect 11483 1699 11491 1719
rect 11454 1689 11491 1699
rect 11550 1719 11637 1729
rect 11550 1699 11559 1719
rect 11579 1699 11637 1719
rect 11550 1690 11637 1699
rect 11550 1689 11587 1690
rect 10140 1645 10826 1678
rect 10140 1588 10179 1645
rect 10788 1643 10826 1645
rect 11606 1637 11637 1690
rect 11667 1719 11704 1798
rect 11875 1811 12268 1815
rect 11875 1794 11894 1811
rect 11914 1795 12268 1811
rect 12288 1795 12291 1815
rect 11914 1794 12291 1795
rect 11875 1790 12291 1794
rect 11875 1789 12216 1790
rect 11819 1729 11850 1730
rect 11667 1699 11676 1719
rect 11696 1699 11704 1719
rect 11667 1689 11704 1699
rect 11763 1722 11850 1729
rect 11763 1719 11824 1722
rect 11763 1699 11772 1719
rect 11792 1702 11824 1719
rect 11845 1702 11850 1722
rect 11792 1699 11850 1702
rect 11763 1692 11850 1699
rect 11875 1719 11912 1789
rect 12178 1788 12215 1789
rect 12027 1729 12063 1730
rect 11875 1699 11884 1719
rect 11904 1699 11912 1719
rect 11763 1690 11819 1692
rect 11763 1689 11800 1690
rect 11875 1689 11912 1699
rect 11971 1719 12119 1729
rect 12287 1728 12316 1729
rect 12219 1726 12316 1728
rect 11971 1699 11980 1719
rect 12000 1715 12090 1719
rect 12000 1699 12033 1715
rect 11971 1690 12033 1699
rect 11971 1689 12008 1690
rect 12027 1677 12033 1690
rect 12056 1699 12090 1715
rect 12110 1699 12119 1719
rect 12056 1690 12119 1699
rect 12177 1719 12316 1726
rect 12177 1699 12186 1719
rect 12206 1699 12316 1719
rect 12177 1690 12316 1699
rect 12056 1677 12063 1690
rect 12082 1689 12119 1690
rect 12178 1689 12215 1690
rect 12027 1638 12063 1677
rect 11498 1636 11539 1637
rect 11390 1629 11539 1636
rect 11390 1609 11508 1629
rect 11528 1609 11539 1629
rect 11390 1601 11539 1609
rect 11606 1633 11965 1637
rect 11606 1628 11928 1633
rect 11606 1604 11719 1628
rect 11743 1609 11928 1628
rect 11952 1609 11965 1633
rect 11743 1604 11965 1609
rect 11606 1601 11965 1604
rect 12027 1601 12062 1638
rect 12130 1635 12230 1638
rect 12130 1631 12197 1635
rect 12130 1605 12142 1631
rect 12168 1609 12197 1631
rect 12223 1609 12230 1635
rect 12168 1605 12230 1609
rect 12130 1601 12230 1605
rect 10140 1586 10188 1588
rect 10140 1568 10151 1586
rect 10169 1568 10188 1586
rect 11606 1580 11637 1601
rect 12027 1580 12063 1601
rect 11449 1579 11486 1580
rect 10140 1559 10188 1568
rect 10141 1558 10188 1559
rect 10454 1563 10564 1577
rect 10454 1560 10497 1563
rect 10454 1555 10458 1560
rect 10376 1533 10458 1555
rect 10487 1533 10497 1560
rect 10525 1536 10532 1563
rect 10561 1555 10564 1563
rect 11448 1570 11486 1579
rect 10561 1536 10626 1555
rect 11448 1550 11457 1570
rect 11477 1550 11486 1570
rect 10525 1533 10626 1536
rect 10376 1531 10626 1533
rect 10144 1495 10181 1496
rect 9843 1465 9853 1483
rect 9871 1465 9883 1483
rect 9843 1460 9883 1465
rect 10140 1492 10181 1495
rect 10140 1487 10182 1492
rect 10140 1469 10153 1487
rect 10171 1469 10182 1487
rect 9843 1456 9880 1460
rect 10140 1455 10182 1469
rect 10220 1455 10267 1459
rect 10140 1449 10267 1455
rect 9516 1437 9553 1438
rect 9466 1428 9553 1437
rect 9466 1408 9524 1428
rect 9544 1408 9553 1428
rect 9466 1398 9553 1408
rect 9612 1428 9649 1438
rect 9612 1408 9620 1428
rect 9640 1408 9649 1428
rect 9466 1397 9497 1398
rect 9461 1329 9571 1342
rect 9612 1329 9649 1408
rect 10140 1420 10228 1449
rect 10257 1420 10267 1449
rect 10376 1452 10413 1531
rect 10454 1518 10564 1531
rect 10528 1462 10559 1463
rect 10376 1432 10385 1452
rect 10405 1432 10413 1452
rect 10376 1422 10413 1432
rect 10472 1452 10559 1462
rect 10472 1432 10481 1452
rect 10501 1432 10559 1452
rect 10472 1423 10559 1432
rect 10472 1422 10509 1423
rect 10140 1416 10267 1420
rect 10140 1399 10179 1416
rect 10220 1415 10267 1416
rect 9846 1393 9883 1394
rect 9842 1384 9883 1393
rect 9842 1366 9855 1384
rect 9873 1366 9883 1384
rect 10140 1381 10151 1399
rect 10169 1381 10179 1399
rect 10140 1372 10179 1381
rect 10141 1371 10178 1372
rect 10528 1370 10559 1423
rect 10589 1452 10626 1531
rect 10797 1528 11190 1548
rect 11210 1528 11213 1548
rect 11448 1542 11486 1550
rect 11552 1574 11637 1580
rect 11662 1579 11699 1580
rect 11552 1554 11560 1574
rect 11580 1554 11637 1574
rect 11552 1546 11637 1554
rect 11661 1570 11699 1579
rect 11661 1550 11670 1570
rect 11690 1550 11699 1570
rect 11552 1545 11588 1546
rect 11661 1542 11699 1550
rect 11765 1574 11850 1580
rect 11870 1579 11907 1580
rect 11765 1554 11773 1574
rect 11793 1573 11850 1574
rect 11793 1554 11822 1573
rect 11765 1553 11822 1554
rect 11843 1553 11850 1573
rect 11765 1546 11850 1553
rect 11869 1570 11907 1579
rect 11869 1550 11878 1570
rect 11898 1550 11907 1570
rect 11765 1545 11801 1546
rect 11869 1542 11907 1550
rect 11973 1574 12117 1580
rect 11973 1554 11981 1574
rect 12001 1554 12089 1574
rect 12109 1554 12117 1574
rect 11973 1546 12117 1554
rect 11973 1545 12009 1546
rect 12081 1545 12117 1546
rect 12183 1579 12220 1580
rect 12183 1578 12221 1579
rect 12183 1570 12247 1578
rect 12183 1550 12192 1570
rect 12212 1556 12247 1570
rect 12267 1556 12270 1576
rect 12212 1551 12270 1556
rect 12212 1550 12247 1551
rect 10797 1523 11213 1528
rect 10797 1522 11138 1523
rect 10741 1462 10772 1463
rect 10589 1432 10598 1452
rect 10618 1432 10626 1452
rect 10589 1422 10626 1432
rect 10685 1455 10772 1462
rect 10685 1452 10746 1455
rect 10685 1432 10694 1452
rect 10714 1435 10746 1452
rect 10767 1435 10772 1455
rect 10714 1432 10772 1435
rect 10685 1425 10772 1432
rect 10797 1452 10834 1522
rect 11100 1521 11137 1522
rect 11449 1513 11486 1542
rect 11450 1511 11486 1513
rect 11662 1511 11699 1542
rect 11450 1489 11699 1511
rect 11870 1510 11907 1542
rect 12183 1538 12247 1550
rect 12287 1512 12316 1690
rect 12684 1683 12711 1861
rect 12751 1823 12815 1835
rect 13091 1831 13128 1863
rect 13299 1862 13548 1884
rect 13299 1831 13336 1862
rect 13512 1860 13548 1862
rect 13512 1831 13549 1860
rect 13861 1851 13898 1852
rect 14164 1851 14201 1921
rect 14226 1941 14313 1948
rect 14226 1938 14284 1941
rect 14226 1918 14231 1938
rect 14252 1921 14284 1938
rect 14304 1921 14313 1941
rect 14252 1918 14313 1921
rect 14226 1911 14313 1918
rect 14372 1941 14409 1951
rect 14372 1921 14380 1941
rect 14400 1921 14409 1941
rect 14226 1910 14257 1911
rect 13860 1850 14201 1851
rect 13785 1845 14201 1850
rect 12751 1822 12786 1823
rect 12728 1817 12786 1822
rect 12728 1797 12731 1817
rect 12751 1803 12786 1817
rect 12806 1803 12815 1823
rect 12751 1795 12815 1803
rect 12777 1794 12815 1795
rect 12778 1793 12815 1794
rect 12881 1827 12917 1828
rect 12989 1827 13025 1828
rect 12881 1822 13025 1827
rect 12881 1819 12941 1822
rect 12881 1799 12889 1819
rect 12909 1801 12941 1819
rect 12968 1819 13025 1822
rect 12968 1801 12997 1819
rect 12909 1799 12997 1801
rect 13017 1799 13025 1819
rect 12881 1793 13025 1799
rect 13091 1823 13129 1831
rect 13197 1827 13233 1828
rect 13091 1803 13100 1823
rect 13120 1803 13129 1823
rect 13091 1794 13129 1803
rect 13148 1820 13233 1827
rect 13148 1800 13155 1820
rect 13176 1819 13233 1820
rect 13176 1800 13205 1819
rect 13148 1799 13205 1800
rect 13225 1799 13233 1819
rect 13091 1793 13128 1794
rect 13148 1793 13233 1799
rect 13299 1823 13337 1831
rect 13410 1827 13446 1828
rect 13299 1803 13308 1823
rect 13328 1803 13337 1823
rect 13299 1794 13337 1803
rect 13361 1819 13446 1827
rect 13361 1799 13418 1819
rect 13438 1799 13446 1819
rect 13299 1793 13336 1794
rect 13361 1793 13446 1799
rect 13512 1823 13550 1831
rect 13785 1825 13788 1845
rect 13808 1825 14201 1845
rect 14372 1842 14409 1921
rect 14439 1950 14470 2003
rect 14820 2001 14857 2002
rect 14819 1992 14858 2001
rect 14819 1974 14829 1992
rect 14847 1974 14858 1992
rect 15199 1990 15236 1994
rect 14731 1957 14778 1958
rect 14819 1957 14858 1974
rect 14731 1953 14858 1957
rect 14489 1950 14526 1951
rect 14439 1941 14526 1950
rect 14439 1921 14497 1941
rect 14517 1921 14526 1941
rect 14439 1911 14526 1921
rect 14585 1941 14622 1951
rect 14585 1921 14593 1941
rect 14613 1921 14622 1941
rect 14439 1910 14470 1911
rect 14434 1842 14544 1855
rect 14585 1842 14622 1921
rect 14731 1924 14741 1953
rect 14770 1924 14858 1953
rect 14731 1918 14858 1924
rect 14731 1914 14778 1918
rect 14816 1904 14858 1918
rect 14816 1886 14827 1904
rect 14845 1886 14858 1904
rect 14816 1881 14858 1886
rect 14817 1878 14858 1881
rect 15196 1985 15236 1990
rect 15196 1967 15208 1985
rect 15226 1967 15236 1985
rect 14817 1877 14854 1878
rect 14372 1840 14622 1842
rect 14372 1837 14473 1840
rect 13512 1803 13521 1823
rect 13541 1803 13550 1823
rect 14372 1818 14437 1837
rect 13512 1794 13550 1803
rect 14434 1810 14437 1818
rect 14466 1810 14473 1837
rect 14501 1813 14511 1840
rect 14540 1818 14622 1840
rect 14540 1813 14544 1818
rect 14501 1810 14544 1813
rect 14434 1796 14544 1810
rect 14810 1814 14857 1815
rect 14810 1805 14858 1814
rect 13512 1793 13549 1794
rect 12935 1772 12971 1793
rect 13361 1772 13392 1793
rect 14810 1787 14829 1805
rect 14847 1787 14858 1805
rect 14810 1785 14858 1787
rect 12768 1768 12868 1772
rect 12768 1764 12830 1768
rect 12768 1738 12775 1764
rect 12801 1742 12830 1764
rect 12856 1742 12868 1768
rect 12801 1738 12868 1742
rect 12768 1735 12868 1738
rect 12936 1735 12971 1772
rect 13033 1769 13392 1772
rect 13033 1764 13255 1769
rect 13033 1740 13046 1764
rect 13070 1745 13255 1764
rect 13279 1745 13392 1769
rect 13070 1740 13392 1745
rect 13033 1736 13392 1740
rect 13459 1764 13608 1772
rect 13459 1744 13470 1764
rect 13490 1744 13608 1764
rect 13459 1737 13608 1744
rect 13459 1736 13500 1737
rect 12783 1683 12820 1684
rect 12879 1683 12916 1684
rect 12935 1683 12971 1735
rect 12990 1683 13027 1684
rect 12683 1674 12821 1683
rect 12683 1654 12792 1674
rect 12812 1654 12821 1674
rect 12683 1647 12821 1654
rect 12879 1674 13027 1683
rect 12879 1654 12888 1674
rect 12908 1654 12998 1674
rect 13018 1654 13027 1674
rect 12683 1645 12779 1647
rect 12879 1644 13027 1654
rect 13086 1674 13123 1684
rect 13198 1683 13235 1684
rect 13179 1681 13235 1683
rect 13086 1654 13094 1674
rect 13114 1654 13123 1674
rect 12935 1643 12971 1644
rect 12783 1584 12820 1585
rect 13086 1584 13123 1654
rect 13148 1674 13235 1681
rect 13148 1671 13206 1674
rect 13148 1651 13153 1671
rect 13174 1654 13206 1671
rect 13226 1654 13235 1674
rect 13174 1651 13235 1654
rect 13148 1644 13235 1651
rect 13294 1674 13331 1684
rect 13294 1654 13302 1674
rect 13322 1654 13331 1674
rect 13148 1643 13179 1644
rect 12782 1583 13123 1584
rect 12707 1579 13123 1583
rect 12707 1578 13084 1579
rect 12707 1558 12710 1578
rect 12730 1562 13084 1578
rect 13104 1562 13123 1579
rect 12730 1558 13123 1562
rect 13294 1575 13331 1654
rect 13361 1683 13392 1736
rect 14172 1728 14210 1730
rect 14819 1728 14858 1785
rect 14172 1695 14858 1728
rect 13411 1683 13448 1684
rect 13361 1674 13448 1683
rect 13361 1654 13419 1674
rect 13439 1654 13448 1674
rect 13361 1644 13448 1654
rect 13507 1674 13544 1684
rect 13507 1654 13515 1674
rect 13535 1654 13544 1674
rect 13361 1643 13392 1644
rect 13356 1575 13466 1588
rect 13507 1575 13544 1654
rect 13294 1573 13544 1575
rect 13294 1570 13395 1573
rect 13294 1551 13359 1570
rect 13356 1543 13359 1551
rect 13388 1543 13395 1570
rect 13423 1546 13433 1573
rect 13462 1551 13544 1573
rect 13764 1607 13932 1608
rect 14172 1607 14210 1695
rect 14471 1693 14518 1695
rect 14818 1671 14858 1695
rect 13764 1584 14210 1607
rect 14436 1638 14547 1653
rect 14436 1636 14478 1638
rect 14436 1616 14443 1636
rect 14462 1616 14478 1636
rect 14436 1608 14478 1616
rect 14506 1636 14547 1638
rect 14506 1616 14520 1636
rect 14539 1616 14547 1636
rect 14819 1627 14858 1671
rect 14506 1608 14547 1616
rect 14436 1602 14547 1608
rect 13764 1581 14208 1584
rect 13764 1579 13932 1581
rect 13462 1546 13466 1551
rect 13423 1543 13466 1546
rect 13356 1529 13466 1543
rect 12146 1510 12316 1512
rect 11867 1503 12316 1510
rect 11531 1483 11642 1489
rect 11531 1475 11572 1483
rect 10949 1462 10985 1463
rect 10797 1432 10806 1452
rect 10826 1432 10834 1452
rect 10685 1423 10741 1425
rect 10685 1422 10722 1423
rect 10797 1422 10834 1432
rect 10893 1452 11041 1462
rect 11141 1459 11237 1461
rect 10893 1432 10902 1452
rect 10922 1432 11012 1452
rect 11032 1432 11041 1452
rect 10893 1423 11041 1432
rect 11099 1452 11237 1459
rect 11099 1432 11108 1452
rect 11128 1432 11237 1452
rect 11531 1455 11539 1475
rect 11558 1455 11572 1475
rect 11531 1453 11572 1455
rect 11600 1475 11642 1483
rect 11600 1455 11616 1475
rect 11635 1455 11642 1475
rect 11867 1476 11892 1503
rect 11923 1484 12316 1503
rect 11923 1476 11972 1484
rect 12146 1483 12316 1484
rect 11867 1474 11972 1476
rect 11600 1453 11642 1455
rect 11531 1438 11642 1453
rect 11099 1423 11237 1432
rect 10893 1422 10930 1423
rect 10949 1371 10985 1423
rect 11004 1422 11041 1423
rect 11100 1422 11137 1423
rect 10420 1369 10461 1370
rect 9842 1357 9883 1366
rect 10312 1362 10461 1369
rect 9842 1337 9882 1357
rect 9399 1327 9649 1329
rect 9399 1324 9500 1327
rect 7917 1267 7981 1279
rect 8257 1275 8294 1302
rect 8465 1275 8502 1306
rect 8678 1304 8714 1306
rect 9399 1305 9464 1324
rect 8678 1275 8715 1304
rect 9461 1297 9464 1305
rect 9493 1297 9500 1324
rect 9528 1300 9538 1327
rect 9567 1305 9649 1327
rect 9757 1327 9882 1337
rect 10312 1342 10430 1362
rect 10450 1342 10461 1362
rect 10312 1334 10461 1342
rect 10528 1366 10887 1370
rect 10528 1361 10850 1366
rect 10528 1337 10641 1361
rect 10665 1342 10850 1361
rect 10874 1342 10887 1366
rect 10665 1337 10887 1342
rect 10528 1334 10887 1337
rect 10949 1334 10984 1371
rect 11052 1368 11152 1371
rect 11052 1364 11119 1368
rect 11052 1338 11064 1364
rect 11090 1342 11119 1364
rect 11145 1342 11152 1368
rect 11090 1338 11152 1342
rect 11052 1334 11152 1338
rect 9757 1308 9765 1327
rect 9790 1308 9882 1327
rect 10528 1313 10559 1334
rect 10949 1313 10985 1334
rect 10371 1312 10408 1313
rect 10145 1309 10179 1310
rect 9567 1300 9571 1305
rect 9757 1301 9882 1308
rect 9528 1297 9571 1300
rect 9461 1283 9571 1297
rect 7917 1266 7952 1267
rect 7894 1261 7952 1266
rect 7894 1241 7897 1261
rect 7917 1247 7952 1261
rect 7972 1247 7981 1267
rect 7917 1239 7981 1247
rect 7943 1238 7981 1239
rect 7944 1237 7981 1238
rect 8047 1271 8083 1272
rect 8155 1271 8191 1272
rect 8047 1263 8191 1271
rect 8047 1243 8055 1263
rect 8075 1260 8163 1263
rect 8075 1243 8107 1260
rect 8127 1243 8163 1260
rect 8183 1243 8191 1263
rect 8047 1237 8191 1243
rect 8257 1267 8295 1275
rect 8363 1271 8399 1272
rect 8257 1247 8266 1267
rect 8286 1247 8295 1267
rect 8257 1238 8295 1247
rect 8314 1264 8399 1271
rect 8314 1244 8321 1264
rect 8342 1263 8399 1264
rect 8342 1244 8371 1263
rect 8314 1243 8371 1244
rect 8391 1243 8399 1263
rect 8257 1237 8294 1238
rect 8314 1237 8399 1243
rect 8465 1267 8503 1275
rect 8576 1271 8612 1272
rect 8465 1247 8474 1267
rect 8494 1247 8503 1267
rect 8465 1238 8503 1247
rect 8527 1263 8612 1271
rect 8527 1243 8584 1263
rect 8604 1243 8612 1263
rect 8465 1237 8502 1238
rect 8527 1237 8612 1243
rect 8678 1267 8716 1275
rect 8678 1247 8687 1267
rect 8707 1247 8716 1267
rect 8678 1238 8716 1247
rect 9842 1253 9882 1301
rect 10144 1300 10181 1309
rect 10144 1282 10153 1300
rect 10171 1282 10181 1300
rect 10144 1272 10181 1282
rect 10370 1303 10408 1312
rect 10370 1283 10379 1303
rect 10399 1283 10408 1303
rect 10370 1275 10408 1283
rect 10474 1307 10559 1313
rect 10584 1312 10621 1313
rect 10474 1287 10482 1307
rect 10502 1287 10559 1307
rect 10474 1279 10559 1287
rect 10583 1303 10621 1312
rect 10583 1283 10592 1303
rect 10612 1283 10621 1303
rect 10474 1278 10510 1279
rect 10583 1275 10621 1283
rect 10687 1307 10772 1313
rect 10792 1312 10829 1313
rect 10687 1287 10695 1307
rect 10715 1306 10772 1307
rect 10715 1287 10744 1306
rect 10687 1286 10744 1287
rect 10765 1286 10772 1306
rect 10687 1279 10772 1286
rect 10791 1303 10829 1312
rect 10791 1283 10800 1303
rect 10820 1283 10829 1303
rect 10687 1278 10723 1279
rect 10791 1275 10829 1283
rect 10895 1307 11039 1313
rect 10895 1287 10903 1307
rect 10923 1306 11011 1307
rect 10923 1287 10954 1306
rect 10895 1286 10954 1287
rect 10979 1287 11011 1306
rect 11031 1287 11039 1307
rect 10979 1286 11039 1287
rect 10895 1279 11039 1286
rect 10895 1278 10931 1279
rect 11003 1278 11039 1279
rect 11105 1312 11142 1313
rect 11105 1311 11143 1312
rect 11105 1303 11169 1311
rect 11105 1283 11114 1303
rect 11134 1289 11169 1303
rect 11189 1289 11192 1309
rect 11134 1284 11192 1289
rect 11134 1283 11169 1284
rect 8678 1237 8715 1238
rect 8101 1216 8137 1237
rect 8527 1216 8558 1237
rect 9842 1235 9853 1253
rect 9871 1235 9882 1253
rect 9842 1227 9882 1235
rect 10145 1244 10179 1272
rect 10371 1246 10408 1275
rect 10372 1244 10408 1246
rect 10584 1244 10621 1275
rect 10145 1243 10317 1244
rect 9843 1226 9880 1227
rect 7934 1212 8034 1216
rect 7934 1208 7996 1212
rect 7934 1182 7941 1208
rect 7967 1186 7996 1208
rect 8022 1186 8034 1212
rect 7967 1182 8034 1186
rect 7934 1179 8034 1182
rect 8102 1179 8137 1216
rect 8199 1213 8558 1216
rect 8199 1208 8421 1213
rect 8199 1184 8212 1208
rect 8236 1189 8421 1208
rect 8445 1189 8558 1213
rect 8236 1184 8558 1189
rect 8199 1180 8558 1184
rect 8625 1208 8774 1216
rect 8625 1188 8636 1208
rect 8656 1188 8774 1208
rect 8625 1181 8774 1188
rect 10145 1211 10331 1243
rect 10372 1222 10621 1244
rect 10792 1243 10829 1275
rect 11105 1271 11169 1283
rect 11209 1245 11236 1423
rect 13764 1401 13791 1579
rect 13831 1541 13895 1553
rect 14171 1549 14208 1581
rect 14379 1580 14628 1602
rect 14379 1549 14416 1580
rect 14592 1578 14628 1580
rect 14592 1549 14629 1578
rect 13831 1540 13866 1541
rect 13808 1535 13866 1540
rect 13808 1515 13811 1535
rect 13831 1521 13866 1535
rect 13886 1521 13895 1541
rect 13831 1513 13895 1521
rect 13857 1512 13895 1513
rect 13858 1511 13895 1512
rect 13961 1545 13997 1546
rect 14069 1545 14105 1546
rect 13961 1540 14105 1545
rect 13961 1537 14023 1540
rect 13961 1517 13969 1537
rect 13989 1520 14023 1537
rect 14046 1537 14105 1540
rect 14046 1520 14077 1537
rect 13989 1517 14077 1520
rect 14097 1517 14105 1537
rect 13961 1511 14105 1517
rect 14171 1541 14209 1549
rect 14277 1545 14313 1546
rect 14171 1521 14180 1541
rect 14200 1521 14209 1541
rect 14171 1512 14209 1521
rect 14228 1538 14313 1545
rect 14228 1518 14235 1538
rect 14256 1537 14313 1538
rect 14256 1518 14285 1537
rect 14228 1517 14285 1518
rect 14305 1517 14313 1537
rect 14171 1511 14208 1512
rect 14228 1511 14313 1517
rect 14379 1541 14417 1549
rect 14490 1545 14526 1546
rect 14379 1521 14388 1541
rect 14408 1521 14417 1541
rect 14379 1512 14417 1521
rect 14441 1537 14526 1545
rect 14441 1517 14498 1537
rect 14518 1517 14526 1537
rect 14379 1511 14416 1512
rect 14441 1511 14526 1517
rect 14592 1541 14630 1549
rect 14592 1521 14601 1541
rect 14621 1521 14630 1541
rect 14592 1512 14630 1521
rect 14592 1511 14629 1512
rect 14015 1490 14051 1511
rect 14441 1490 14472 1511
rect 13848 1486 13948 1490
rect 13848 1482 13910 1486
rect 13848 1456 13855 1482
rect 13881 1460 13910 1482
rect 13936 1460 13948 1486
rect 13881 1456 13948 1460
rect 13848 1453 13948 1456
rect 14016 1453 14051 1490
rect 14113 1487 14472 1490
rect 14113 1482 14335 1487
rect 14113 1458 14126 1482
rect 14150 1463 14335 1482
rect 14359 1463 14472 1487
rect 14150 1458 14472 1463
rect 14113 1454 14472 1458
rect 14539 1482 14688 1490
rect 14539 1462 14550 1482
rect 14570 1462 14688 1482
rect 14539 1455 14688 1462
rect 14539 1454 14580 1455
rect 13863 1401 13900 1402
rect 13959 1401 13996 1402
rect 14015 1401 14051 1453
rect 14070 1401 14107 1402
rect 13763 1392 13901 1401
rect 13763 1372 13872 1392
rect 13892 1372 13901 1392
rect 13763 1365 13901 1372
rect 13959 1392 14107 1401
rect 13959 1372 13968 1392
rect 13988 1372 14078 1392
rect 14098 1372 14107 1392
rect 13763 1363 13859 1365
rect 13959 1362 14107 1372
rect 14166 1392 14203 1402
rect 14278 1401 14315 1402
rect 14259 1399 14315 1401
rect 14166 1372 14174 1392
rect 14194 1372 14203 1392
rect 14015 1361 14051 1362
rect 11392 1319 11502 1333
rect 11392 1316 11435 1319
rect 11392 1311 11396 1316
rect 11068 1243 11236 1245
rect 10792 1237 11236 1243
rect 9214 1185 9728 1186
rect 8625 1180 8666 1181
rect 7949 1127 7986 1128
rect 8045 1127 8082 1128
rect 8101 1127 8137 1179
rect 8156 1127 8193 1128
rect 7849 1118 7987 1127
rect 7849 1098 7958 1118
rect 7978 1098 7987 1118
rect 7849 1091 7987 1098
rect 8045 1118 8193 1127
rect 8045 1098 8054 1118
rect 8074 1098 8164 1118
rect 8184 1098 8193 1118
rect 7849 1089 7945 1091
rect 8045 1088 8193 1098
rect 8252 1118 8289 1128
rect 8364 1127 8401 1128
rect 8345 1125 8401 1127
rect 8252 1098 8260 1118
rect 8280 1098 8289 1118
rect 8101 1087 8137 1088
rect 7031 1035 7199 1037
rect 6753 1029 7199 1035
rect 5821 1005 6237 1010
rect 6416 1008 6527 1014
rect 5821 1004 6162 1005
rect 5765 944 5796 945
rect 5613 914 5622 934
rect 5642 914 5650 934
rect 5613 904 5650 914
rect 5709 937 5796 944
rect 5709 934 5770 937
rect 5709 914 5718 934
rect 5738 917 5770 934
rect 5791 917 5796 937
rect 5738 914 5796 917
rect 5709 907 5796 914
rect 5821 934 5858 1004
rect 6124 1003 6161 1004
rect 6416 1000 6457 1008
rect 6416 980 6424 1000
rect 6443 980 6457 1000
rect 6416 978 6457 980
rect 6485 1000 6527 1008
rect 6485 980 6501 1000
rect 6520 980 6527 1000
rect 6753 1007 6759 1029
rect 6785 1009 7199 1029
rect 7949 1028 7986 1029
rect 8252 1028 8289 1098
rect 8314 1118 8401 1125
rect 8314 1115 8372 1118
rect 8314 1095 8319 1115
rect 8340 1098 8372 1115
rect 8392 1098 8401 1118
rect 8340 1095 8401 1098
rect 8314 1088 8401 1095
rect 8460 1118 8497 1128
rect 8460 1098 8468 1118
rect 8488 1098 8497 1118
rect 8314 1087 8345 1088
rect 7948 1027 8289 1028
rect 6785 1007 6794 1009
rect 7031 1008 7199 1009
rect 7873 1022 8289 1027
rect 6753 998 6794 1007
rect 7873 1002 7876 1022
rect 7896 1002 8289 1022
rect 8460 1019 8497 1098
rect 8527 1127 8558 1180
rect 9195 1169 9728 1185
rect 10145 1179 10179 1211
rect 10141 1170 10179 1179
rect 9195 1158 9727 1169
rect 9846 1160 9883 1164
rect 8577 1127 8614 1128
rect 8527 1118 8614 1127
rect 8527 1098 8585 1118
rect 8605 1098 8614 1118
rect 8527 1088 8614 1098
rect 8673 1118 8710 1128
rect 8673 1098 8681 1118
rect 8701 1098 8710 1118
rect 8527 1087 8558 1088
rect 8522 1019 8632 1032
rect 8673 1019 8710 1098
rect 8460 1017 8710 1019
rect 8460 1014 8561 1017
rect 8460 995 8525 1014
rect 6485 978 6527 980
rect 6416 963 6527 978
rect 8522 987 8525 995
rect 8554 987 8561 1014
rect 8589 990 8599 1017
rect 8628 995 8710 1017
rect 8788 1089 8956 1090
rect 9195 1089 9233 1158
rect 8788 1069 9233 1089
rect 9460 1120 9571 1135
rect 9460 1118 9502 1120
rect 9460 1098 9467 1118
rect 9486 1098 9502 1118
rect 9460 1090 9502 1098
rect 9530 1118 9571 1120
rect 9530 1098 9544 1118
rect 9563 1098 9571 1118
rect 9530 1090 9571 1098
rect 9460 1084 9571 1090
rect 9693 1095 9727 1158
rect 9845 1154 9883 1160
rect 9845 1136 9855 1154
rect 9873 1136 9883 1154
rect 10141 1152 10151 1170
rect 10169 1152 10179 1170
rect 10141 1146 10179 1152
rect 10297 1148 10331 1211
rect 10453 1216 10564 1222
rect 10453 1208 10494 1216
rect 10453 1188 10461 1208
rect 10480 1188 10494 1208
rect 10453 1186 10494 1188
rect 10522 1208 10564 1216
rect 10522 1188 10538 1208
rect 10557 1188 10564 1208
rect 10522 1186 10564 1188
rect 10453 1171 10564 1186
rect 10791 1217 11236 1237
rect 10791 1148 10829 1217
rect 11068 1216 11236 1217
rect 11314 1289 11396 1311
rect 11425 1289 11435 1316
rect 11463 1292 11470 1319
rect 11499 1311 11502 1319
rect 13497 1328 13608 1343
rect 13497 1326 13539 1328
rect 11499 1292 11564 1311
rect 11463 1289 11564 1292
rect 11314 1287 11564 1289
rect 11314 1208 11351 1287
rect 11392 1274 11502 1287
rect 11466 1218 11497 1219
rect 11314 1188 11323 1208
rect 11343 1188 11351 1208
rect 11314 1178 11351 1188
rect 11410 1208 11497 1218
rect 11410 1188 11419 1208
rect 11439 1188 11497 1208
rect 11410 1179 11497 1188
rect 11410 1178 11447 1179
rect 10141 1142 10178 1146
rect 10297 1137 10829 1148
rect 9845 1127 9883 1136
rect 9845 1095 9879 1127
rect 10296 1121 10829 1137
rect 11466 1126 11497 1179
rect 11527 1208 11564 1287
rect 11735 1297 12128 1304
rect 11735 1280 11743 1297
rect 11775 1284 12128 1297
rect 12148 1284 12151 1304
rect 13230 1299 13271 1308
rect 11775 1280 12151 1284
rect 11735 1279 12151 1280
rect 12825 1297 12993 1298
rect 13230 1297 13239 1299
rect 11735 1278 12076 1279
rect 11679 1218 11710 1219
rect 11527 1188 11536 1208
rect 11556 1188 11564 1208
rect 11527 1178 11564 1188
rect 11623 1211 11710 1218
rect 11623 1208 11684 1211
rect 11623 1188 11632 1208
rect 11652 1191 11684 1208
rect 11705 1191 11710 1211
rect 11652 1188 11710 1191
rect 11623 1181 11710 1188
rect 11735 1208 11772 1278
rect 12038 1277 12075 1278
rect 12825 1277 13239 1297
rect 13265 1277 13271 1299
rect 13497 1306 13504 1326
rect 13523 1306 13539 1326
rect 13497 1298 13539 1306
rect 13567 1326 13608 1328
rect 13567 1306 13581 1326
rect 13600 1306 13608 1326
rect 13567 1298 13608 1306
rect 13863 1302 13900 1303
rect 14166 1302 14203 1372
rect 14228 1392 14315 1399
rect 14228 1389 14286 1392
rect 14228 1369 14233 1389
rect 14254 1372 14286 1389
rect 14306 1372 14315 1392
rect 14254 1369 14315 1372
rect 14228 1362 14315 1369
rect 14374 1392 14411 1402
rect 14374 1372 14382 1392
rect 14402 1372 14411 1392
rect 14228 1361 14259 1362
rect 13862 1301 14203 1302
rect 13497 1292 13608 1298
rect 13787 1296 14203 1301
rect 12825 1271 13271 1277
rect 12825 1269 12993 1271
rect 11887 1218 11923 1219
rect 11735 1188 11744 1208
rect 11764 1188 11772 1208
rect 11623 1179 11679 1181
rect 11623 1178 11660 1179
rect 11735 1178 11772 1188
rect 11831 1208 11979 1218
rect 12079 1215 12175 1217
rect 11831 1188 11840 1208
rect 11860 1203 11950 1208
rect 11860 1188 11895 1203
rect 11831 1179 11895 1188
rect 11831 1178 11868 1179
rect 11887 1162 11895 1179
rect 11916 1188 11950 1203
rect 11970 1188 11979 1208
rect 11916 1179 11979 1188
rect 12037 1208 12175 1215
rect 12037 1188 12046 1208
rect 12066 1188 12175 1208
rect 12037 1179 12175 1188
rect 11916 1162 11923 1179
rect 11942 1178 11979 1179
rect 12038 1178 12075 1179
rect 11887 1127 11923 1162
rect 11358 1125 11399 1126
rect 10296 1120 10810 1121
rect 8788 1063 9232 1069
rect 8788 1061 8956 1063
rect 8628 990 8632 995
rect 8589 987 8632 990
rect 8522 973 8632 987
rect 5973 944 6009 945
rect 5821 914 5830 934
rect 5850 914 5858 934
rect 5709 905 5765 907
rect 5709 904 5746 905
rect 5821 904 5858 914
rect 5917 934 6065 944
rect 6165 941 6261 943
rect 5917 914 5926 934
rect 5946 914 6036 934
rect 6056 914 6065 934
rect 5917 905 6065 914
rect 6123 934 6261 941
rect 6123 914 6132 934
rect 6152 914 6261 934
rect 6123 905 6261 914
rect 5917 904 5954 905
rect 5973 853 6009 905
rect 6028 904 6065 905
rect 6124 904 6161 905
rect 5444 851 5485 852
rect 5336 844 5485 851
rect 5336 824 5454 844
rect 5474 824 5485 844
rect 5336 816 5485 824
rect 5552 848 5911 852
rect 5552 843 5874 848
rect 5552 819 5665 843
rect 5689 824 5874 843
rect 5898 824 5911 848
rect 5689 819 5911 824
rect 5552 816 5911 819
rect 5973 816 6008 853
rect 6076 850 6176 853
rect 6076 846 6143 850
rect 6076 820 6088 846
rect 6114 824 6143 846
rect 6169 824 6176 850
rect 6114 820 6176 824
rect 6076 816 6176 820
rect 5552 795 5583 816
rect 5973 795 6009 816
rect 5395 794 5432 795
rect 5394 785 5432 794
rect 5394 765 5403 785
rect 5423 765 5432 785
rect 5394 757 5432 765
rect 5498 789 5583 795
rect 5608 794 5645 795
rect 5498 769 5506 789
rect 5526 769 5583 789
rect 5498 761 5583 769
rect 5607 785 5645 794
rect 5607 765 5616 785
rect 5636 765 5645 785
rect 5498 760 5534 761
rect 5607 757 5645 765
rect 5711 789 5796 795
rect 5816 794 5853 795
rect 5711 769 5719 789
rect 5739 788 5796 789
rect 5739 769 5768 788
rect 5711 768 5768 769
rect 5789 768 5796 788
rect 5711 761 5796 768
rect 5815 785 5853 794
rect 5815 765 5824 785
rect 5844 765 5853 785
rect 5711 760 5747 761
rect 5815 757 5853 765
rect 5919 789 6063 795
rect 5919 769 5927 789
rect 5947 786 6035 789
rect 5947 769 5978 786
rect 5919 766 5978 769
rect 6001 769 6035 786
rect 6055 769 6063 789
rect 6001 766 6063 769
rect 5919 761 6063 766
rect 5919 760 5955 761
rect 6027 760 6063 761
rect 6129 794 6166 795
rect 6129 793 6167 794
rect 6129 785 6193 793
rect 6129 765 6138 785
rect 6158 771 6193 785
rect 6213 771 6216 791
rect 6158 766 6216 771
rect 6158 765 6193 766
rect 5395 728 5432 757
rect 5396 726 5432 728
rect 5608 726 5645 757
rect 5396 704 5645 726
rect 5816 725 5853 757
rect 6129 753 6193 765
rect 6233 727 6260 905
rect 8788 883 8815 1061
rect 8855 1023 8919 1035
rect 9195 1031 9232 1063
rect 9403 1062 9652 1084
rect 9693 1063 9879 1095
rect 11250 1118 11399 1125
rect 11250 1098 11368 1118
rect 11388 1098 11399 1118
rect 11250 1090 11399 1098
rect 11466 1122 11825 1126
rect 11466 1117 11788 1122
rect 11466 1093 11579 1117
rect 11603 1098 11788 1117
rect 11812 1098 11825 1122
rect 11603 1093 11825 1098
rect 11466 1090 11825 1093
rect 11887 1090 11922 1127
rect 11990 1124 12090 1127
rect 11990 1120 12057 1124
rect 11990 1094 12002 1120
rect 12028 1098 12057 1120
rect 12083 1098 12090 1124
rect 12028 1094 12090 1098
rect 11990 1090 12090 1094
rect 10144 1079 10181 1080
rect 9707 1062 9879 1063
rect 9403 1031 9440 1062
rect 9616 1060 9652 1062
rect 9616 1031 9653 1060
rect 9845 1034 9879 1062
rect 10142 1071 10182 1079
rect 10142 1053 10153 1071
rect 10171 1053 10182 1071
rect 11466 1069 11497 1090
rect 11887 1069 11923 1090
rect 11309 1068 11346 1069
rect 8855 1022 8890 1023
rect 8832 1017 8890 1022
rect 8832 997 8835 1017
rect 8855 1003 8890 1017
rect 8910 1003 8919 1023
rect 8855 995 8919 1003
rect 8881 994 8919 995
rect 8882 993 8919 994
rect 8985 1027 9021 1028
rect 9093 1027 9129 1028
rect 8985 1020 9129 1027
rect 8985 1019 9045 1020
rect 8985 999 8993 1019
rect 9013 1000 9045 1019
rect 9070 1019 9129 1020
rect 9070 1000 9101 1019
rect 9013 999 9101 1000
rect 9121 999 9129 1019
rect 8985 993 9129 999
rect 9195 1023 9233 1031
rect 9301 1027 9337 1028
rect 9195 1003 9204 1023
rect 9224 1003 9233 1023
rect 9195 994 9233 1003
rect 9252 1020 9337 1027
rect 9252 1000 9259 1020
rect 9280 1019 9337 1020
rect 9280 1000 9309 1019
rect 9252 999 9309 1000
rect 9329 999 9337 1019
rect 9195 993 9232 994
rect 9252 993 9337 999
rect 9403 1023 9441 1031
rect 9514 1027 9550 1028
rect 9403 1003 9412 1023
rect 9432 1003 9441 1023
rect 9403 994 9441 1003
rect 9465 1019 9550 1027
rect 9465 999 9522 1019
rect 9542 999 9550 1019
rect 9403 993 9440 994
rect 9465 993 9550 999
rect 9616 1023 9654 1031
rect 9616 1003 9625 1023
rect 9645 1003 9654 1023
rect 9616 994 9654 1003
rect 9843 1024 9880 1034
rect 9843 1006 9853 1024
rect 9871 1006 9880 1024
rect 9843 997 9880 1006
rect 10142 1005 10182 1053
rect 11308 1059 11346 1068
rect 11308 1039 11317 1059
rect 11337 1039 11346 1059
rect 11308 1031 11346 1039
rect 11412 1063 11497 1069
rect 11522 1068 11559 1069
rect 11412 1043 11420 1063
rect 11440 1043 11497 1063
rect 11412 1035 11497 1043
rect 11521 1059 11559 1068
rect 11521 1039 11530 1059
rect 11550 1039 11559 1059
rect 11412 1034 11448 1035
rect 11521 1031 11559 1039
rect 11625 1063 11710 1069
rect 11730 1068 11767 1069
rect 11625 1043 11633 1063
rect 11653 1062 11710 1063
rect 11653 1043 11682 1062
rect 11625 1042 11682 1043
rect 11703 1042 11710 1062
rect 11625 1035 11710 1042
rect 11729 1059 11767 1068
rect 11729 1039 11738 1059
rect 11758 1039 11767 1059
rect 11625 1034 11661 1035
rect 11729 1031 11767 1039
rect 11833 1063 11977 1069
rect 11833 1043 11841 1063
rect 11861 1043 11949 1063
rect 11969 1043 11977 1063
rect 11833 1035 11977 1043
rect 11833 1034 11869 1035
rect 11941 1034 11977 1035
rect 12043 1068 12080 1069
rect 12043 1067 12081 1068
rect 12043 1059 12107 1067
rect 12043 1039 12052 1059
rect 12072 1045 12107 1059
rect 12127 1045 12130 1065
rect 12072 1040 12130 1045
rect 12072 1039 12107 1040
rect 10453 1009 10563 1023
rect 10453 1006 10496 1009
rect 10142 998 10267 1005
rect 10453 1001 10457 1006
rect 9845 996 9879 997
rect 9616 993 9653 994
rect 9039 972 9075 993
rect 9465 972 9496 993
rect 10142 979 10234 998
rect 10259 979 10267 998
rect 8872 968 8972 972
rect 8872 964 8934 968
rect 8872 938 8879 964
rect 8905 942 8934 964
rect 8960 942 8972 968
rect 8905 938 8972 942
rect 8872 935 8972 938
rect 9040 935 9075 972
rect 9137 969 9496 972
rect 9137 964 9359 969
rect 9137 940 9150 964
rect 9174 945 9359 964
rect 9383 945 9496 969
rect 9174 940 9496 945
rect 9137 936 9496 940
rect 9563 964 9712 972
rect 9563 944 9574 964
rect 9594 944 9712 964
rect 10142 969 10267 979
rect 10375 979 10457 1001
rect 10486 979 10496 1006
rect 10524 982 10531 1009
rect 10560 1001 10563 1009
rect 11309 1002 11346 1031
rect 10560 982 10625 1001
rect 11310 1000 11346 1002
rect 11522 1000 11559 1031
rect 11730 1004 11767 1031
rect 12043 1027 12107 1039
rect 10524 979 10625 982
rect 10375 977 10625 979
rect 10142 949 10182 969
rect 9563 937 9712 944
rect 10141 940 10182 949
rect 9563 936 9604 937
rect 8887 883 8924 884
rect 8983 883 9020 884
rect 9039 883 9075 935
rect 9094 883 9131 884
rect 8787 874 8925 883
rect 8787 854 8896 874
rect 8916 854 8925 874
rect 8787 847 8925 854
rect 8983 874 9131 883
rect 8983 854 8992 874
rect 9012 854 9102 874
rect 9122 854 9131 874
rect 8787 845 8883 847
rect 8983 844 9131 854
rect 9190 874 9227 884
rect 9302 883 9339 884
rect 9283 881 9339 883
rect 9190 854 9198 874
rect 9218 854 9227 874
rect 9039 843 9075 844
rect 8887 784 8924 785
rect 9190 784 9227 854
rect 9252 874 9339 881
rect 9252 871 9310 874
rect 9252 851 9257 871
rect 9278 854 9310 871
rect 9330 854 9339 874
rect 9278 851 9339 854
rect 9252 844 9339 851
rect 9398 874 9435 884
rect 9398 854 9406 874
rect 9426 854 9435 874
rect 9252 843 9283 844
rect 8886 783 9227 784
rect 8811 778 9227 783
rect 8811 758 8814 778
rect 8834 758 9227 778
rect 9398 775 9435 854
rect 9465 883 9496 936
rect 9846 934 9883 935
rect 9845 925 9884 934
rect 9845 907 9855 925
rect 9873 907 9884 925
rect 10141 922 10151 940
rect 10169 922 10182 940
rect 10141 913 10182 922
rect 10141 912 10178 913
rect 9757 890 9804 891
rect 9845 890 9884 907
rect 9757 886 9884 890
rect 9515 883 9552 884
rect 9465 874 9552 883
rect 9465 854 9523 874
rect 9543 854 9552 874
rect 9465 844 9552 854
rect 9611 874 9648 884
rect 9611 854 9619 874
rect 9639 854 9648 874
rect 9465 843 9496 844
rect 9460 775 9570 788
rect 9611 775 9648 854
rect 9757 857 9767 886
rect 9796 857 9884 886
rect 10375 898 10412 977
rect 10453 964 10563 977
rect 10527 908 10558 909
rect 10375 878 10384 898
rect 10404 878 10412 898
rect 10375 868 10412 878
rect 10471 898 10558 908
rect 10471 878 10480 898
rect 10500 878 10558 898
rect 10471 869 10558 878
rect 10471 868 10508 869
rect 9757 851 9884 857
rect 9757 847 9804 851
rect 9842 837 9884 851
rect 10144 846 10181 850
rect 9842 819 9853 837
rect 9871 819 9884 837
rect 9842 814 9884 819
rect 9843 811 9884 814
rect 10141 841 10181 846
rect 10141 823 10153 841
rect 10171 823 10181 841
rect 9843 810 9880 811
rect 9398 773 9648 775
rect 9398 770 9499 773
rect 9398 751 9463 770
rect 9460 743 9463 751
rect 9492 743 9499 770
rect 9527 746 9537 773
rect 9566 751 9648 773
rect 9566 746 9570 751
rect 9527 743 9570 746
rect 9460 729 9570 743
rect 9836 747 9883 748
rect 9836 738 9884 747
rect 6092 725 6260 727
rect 5816 722 6260 725
rect 5477 698 5588 704
rect 5477 690 5518 698
rect 490 649 531 651
rect 490 629 506 649
rect 525 629 531 649
rect 490 627 531 629
rect 421 612 531 627
rect 110 570 150 594
rect 758 584 796 658
rect 1036 657 1204 658
rect 718 570 797 584
rect 110 569 400 570
rect 566 569 797 570
rect 110 567 797 569
rect 110 546 757 567
rect 786 546 797 567
rect 110 537 797 546
rect 4787 571 4831 658
rect 5166 635 5205 679
rect 5477 670 5485 690
rect 5504 670 5518 690
rect 5477 668 5518 670
rect 5546 692 5588 698
rect 5814 699 6260 722
rect 9836 720 9855 738
rect 9873 720 9884 738
rect 9836 718 9884 720
rect 9845 699 9884 718
rect 5546 690 5587 692
rect 5546 670 5562 690
rect 5581 670 5587 690
rect 5546 668 5587 670
rect 5477 653 5587 668
rect 5166 611 5206 635
rect 5814 625 5852 699
rect 6092 698 6260 699
rect 5774 611 5853 625
rect 5166 610 5456 611
rect 5622 610 5853 611
rect 5166 608 5853 610
rect 5166 587 5813 608
rect 5842 587 5853 608
rect 5166 578 5853 587
rect 9843 612 9887 699
rect 9843 591 9848 612
rect 9877 591 9887 612
rect 9843 578 9887 591
rect 10141 643 10181 823
rect 10527 816 10558 869
rect 10588 898 10625 977
rect 10796 974 11189 994
rect 11209 974 11212 994
rect 11310 978 11559 1000
rect 11728 999 11769 1004
rect 12147 1001 12174 1179
rect 12825 1091 12852 1269
rect 13230 1266 13271 1271
rect 13440 1270 13689 1292
rect 13787 1276 13790 1296
rect 13810 1276 14203 1296
rect 14374 1293 14411 1372
rect 14441 1401 14472 1454
rect 14818 1447 14858 1627
rect 15196 1787 15236 1967
rect 15582 1960 15613 2013
rect 15643 2042 15680 2121
rect 15851 2118 16244 2138
rect 16264 2118 16267 2138
rect 16365 2122 16614 2144
rect 16783 2143 16824 2148
rect 17202 2145 17229 2323
rect 17880 2235 17907 2413
rect 18285 2410 18326 2415
rect 18495 2414 18744 2436
rect 18842 2420 18845 2440
rect 18865 2420 19258 2440
rect 19429 2437 19466 2516
rect 19496 2545 19527 2598
rect 19873 2591 19913 2771
rect 19873 2573 19883 2591
rect 19901 2573 19913 2591
rect 19873 2568 19913 2573
rect 19873 2564 19910 2568
rect 19546 2545 19583 2546
rect 19496 2536 19583 2545
rect 19496 2516 19554 2536
rect 19574 2516 19583 2536
rect 19496 2506 19583 2516
rect 19642 2536 19679 2546
rect 19642 2516 19650 2536
rect 19670 2516 19679 2536
rect 19496 2505 19527 2506
rect 19491 2437 19601 2450
rect 19642 2437 19679 2516
rect 19876 2501 19913 2502
rect 19872 2492 19913 2501
rect 19872 2474 19885 2492
rect 19903 2474 19913 2492
rect 19872 2465 19913 2474
rect 19872 2445 19912 2465
rect 19429 2435 19679 2437
rect 19429 2432 19530 2435
rect 17947 2375 18011 2387
rect 18287 2383 18324 2410
rect 18495 2383 18532 2414
rect 18708 2412 18744 2414
rect 19429 2413 19494 2432
rect 18708 2383 18745 2412
rect 19491 2405 19494 2413
rect 19523 2405 19530 2432
rect 19558 2408 19568 2435
rect 19597 2413 19679 2435
rect 19787 2435 19912 2445
rect 19787 2416 19795 2435
rect 19820 2416 19912 2435
rect 19597 2408 19601 2413
rect 19787 2409 19912 2416
rect 19558 2405 19601 2408
rect 19491 2391 19601 2405
rect 17947 2374 17982 2375
rect 17924 2369 17982 2374
rect 17924 2349 17927 2369
rect 17947 2355 17982 2369
rect 18002 2355 18011 2375
rect 17947 2347 18011 2355
rect 17973 2346 18011 2347
rect 17974 2345 18011 2346
rect 18077 2379 18113 2380
rect 18185 2379 18221 2380
rect 18077 2371 18221 2379
rect 18077 2351 18085 2371
rect 18105 2351 18193 2371
rect 18213 2351 18221 2371
rect 18077 2345 18221 2351
rect 18287 2375 18325 2383
rect 18393 2379 18429 2380
rect 18287 2355 18296 2375
rect 18316 2355 18325 2375
rect 18287 2346 18325 2355
rect 18344 2372 18429 2379
rect 18344 2352 18351 2372
rect 18372 2371 18429 2372
rect 18372 2352 18401 2371
rect 18344 2351 18401 2352
rect 18421 2351 18429 2371
rect 18287 2345 18324 2346
rect 18344 2345 18429 2351
rect 18495 2375 18533 2383
rect 18606 2379 18642 2380
rect 18495 2355 18504 2375
rect 18524 2355 18533 2375
rect 18495 2346 18533 2355
rect 18557 2371 18642 2379
rect 18557 2351 18614 2371
rect 18634 2351 18642 2371
rect 18495 2345 18532 2346
rect 18557 2345 18642 2351
rect 18708 2375 18746 2383
rect 18708 2355 18717 2375
rect 18737 2355 18746 2375
rect 18708 2346 18746 2355
rect 19872 2361 19912 2409
rect 18708 2345 18745 2346
rect 18131 2324 18167 2345
rect 18557 2324 18588 2345
rect 19872 2343 19883 2361
rect 19901 2343 19912 2361
rect 19872 2335 19912 2343
rect 19873 2334 19910 2335
rect 17964 2320 18064 2324
rect 17964 2316 18026 2320
rect 17964 2290 17971 2316
rect 17997 2294 18026 2316
rect 18052 2294 18064 2320
rect 17997 2290 18064 2294
rect 17964 2287 18064 2290
rect 18132 2287 18167 2324
rect 18229 2321 18588 2324
rect 18229 2316 18451 2321
rect 18229 2292 18242 2316
rect 18266 2297 18451 2316
rect 18475 2297 18588 2321
rect 18266 2292 18588 2297
rect 18229 2288 18588 2292
rect 18655 2316 18804 2324
rect 18655 2296 18666 2316
rect 18686 2296 18804 2316
rect 18655 2289 18804 2296
rect 19244 2293 19758 2294
rect 18655 2288 18696 2289
rect 18131 2252 18167 2287
rect 17979 2235 18016 2236
rect 18075 2235 18112 2236
rect 18131 2235 18138 2252
rect 17879 2226 18017 2235
rect 17879 2206 17988 2226
rect 18008 2206 18017 2226
rect 17879 2199 18017 2206
rect 18075 2226 18138 2235
rect 18075 2206 18084 2226
rect 18104 2211 18138 2226
rect 18159 2235 18167 2252
rect 18186 2235 18223 2236
rect 18159 2226 18223 2235
rect 18159 2211 18194 2226
rect 18104 2206 18194 2211
rect 18214 2206 18223 2226
rect 17879 2197 17975 2199
rect 18075 2196 18223 2206
rect 18282 2226 18319 2236
rect 18394 2235 18431 2236
rect 18375 2233 18431 2235
rect 18282 2206 18290 2226
rect 18310 2206 18319 2226
rect 18131 2195 18167 2196
rect 17061 2143 17229 2145
rect 16783 2137 17229 2143
rect 15851 2113 16267 2118
rect 16446 2116 16557 2122
rect 15851 2112 16192 2113
rect 15795 2052 15826 2053
rect 15643 2022 15652 2042
rect 15672 2022 15680 2042
rect 15643 2012 15680 2022
rect 15739 2045 15826 2052
rect 15739 2042 15800 2045
rect 15739 2022 15748 2042
rect 15768 2025 15800 2042
rect 15821 2025 15826 2045
rect 15768 2022 15826 2025
rect 15739 2015 15826 2022
rect 15851 2042 15888 2112
rect 16154 2111 16191 2112
rect 16446 2108 16487 2116
rect 16446 2088 16454 2108
rect 16473 2088 16487 2108
rect 16446 2086 16487 2088
rect 16515 2108 16557 2116
rect 16515 2088 16531 2108
rect 16550 2088 16557 2108
rect 16783 2115 16789 2137
rect 16815 2117 17229 2137
rect 17979 2136 18016 2137
rect 18282 2136 18319 2206
rect 18344 2226 18431 2233
rect 18344 2223 18402 2226
rect 18344 2203 18349 2223
rect 18370 2206 18402 2223
rect 18422 2206 18431 2226
rect 18370 2203 18431 2206
rect 18344 2196 18431 2203
rect 18490 2226 18527 2236
rect 18490 2206 18498 2226
rect 18518 2206 18527 2226
rect 18344 2195 18375 2196
rect 17978 2135 18319 2136
rect 16815 2115 16824 2117
rect 17061 2116 17229 2117
rect 17903 2134 18319 2135
rect 17903 2130 18279 2134
rect 16783 2106 16824 2115
rect 17903 2110 17906 2130
rect 17926 2117 18279 2130
rect 18311 2117 18319 2134
rect 17926 2110 18319 2117
rect 18490 2127 18527 2206
rect 18557 2235 18588 2288
rect 19225 2277 19758 2293
rect 19225 2266 19757 2277
rect 19876 2268 19913 2272
rect 18607 2235 18644 2236
rect 18557 2226 18644 2235
rect 18557 2206 18615 2226
rect 18635 2206 18644 2226
rect 18557 2196 18644 2206
rect 18703 2226 18740 2236
rect 18703 2206 18711 2226
rect 18731 2206 18740 2226
rect 18557 2195 18588 2196
rect 18552 2127 18662 2140
rect 18703 2127 18740 2206
rect 18490 2125 18740 2127
rect 18490 2122 18591 2125
rect 18490 2103 18555 2122
rect 16515 2086 16557 2088
rect 16446 2071 16557 2086
rect 18552 2095 18555 2103
rect 18584 2095 18591 2122
rect 18619 2098 18629 2125
rect 18658 2103 18740 2125
rect 18818 2197 18986 2198
rect 19225 2197 19263 2266
rect 18818 2177 19263 2197
rect 19490 2228 19601 2243
rect 19490 2226 19532 2228
rect 19490 2206 19497 2226
rect 19516 2206 19532 2226
rect 19490 2198 19532 2206
rect 19560 2226 19601 2228
rect 19560 2206 19574 2226
rect 19593 2206 19601 2226
rect 19560 2198 19601 2206
rect 19490 2192 19601 2198
rect 19723 2203 19757 2266
rect 19875 2262 19913 2268
rect 19875 2244 19885 2262
rect 19903 2244 19913 2262
rect 19875 2235 19913 2244
rect 19875 2203 19909 2235
rect 18818 2171 19262 2177
rect 18818 2169 18986 2171
rect 18658 2098 18662 2103
rect 18619 2095 18662 2098
rect 18552 2081 18662 2095
rect 16003 2052 16039 2053
rect 15851 2022 15860 2042
rect 15880 2022 15888 2042
rect 15739 2013 15795 2015
rect 15739 2012 15776 2013
rect 15851 2012 15888 2022
rect 15947 2042 16095 2052
rect 16195 2049 16291 2051
rect 15947 2022 15956 2042
rect 15976 2022 16066 2042
rect 16086 2022 16095 2042
rect 15947 2013 16095 2022
rect 16153 2042 16291 2049
rect 16153 2022 16162 2042
rect 16182 2022 16291 2042
rect 16153 2013 16291 2022
rect 15947 2012 15984 2013
rect 16003 1961 16039 2013
rect 16058 2012 16095 2013
rect 16154 2012 16191 2013
rect 15474 1959 15515 1960
rect 15366 1952 15515 1959
rect 15366 1932 15484 1952
rect 15504 1932 15515 1952
rect 15366 1924 15515 1932
rect 15582 1956 15941 1960
rect 15582 1951 15904 1956
rect 15582 1927 15695 1951
rect 15719 1932 15904 1951
rect 15928 1932 15941 1956
rect 15719 1927 15941 1932
rect 15582 1924 15941 1927
rect 16003 1924 16038 1961
rect 16106 1958 16206 1961
rect 16106 1954 16173 1958
rect 16106 1928 16118 1954
rect 16144 1932 16173 1954
rect 16199 1932 16206 1958
rect 16144 1928 16206 1932
rect 16106 1924 16206 1928
rect 15582 1903 15613 1924
rect 16003 1903 16039 1924
rect 15425 1902 15462 1903
rect 15424 1893 15462 1902
rect 15424 1873 15433 1893
rect 15453 1873 15462 1893
rect 15424 1865 15462 1873
rect 15528 1897 15613 1903
rect 15638 1902 15675 1903
rect 15528 1877 15536 1897
rect 15556 1877 15613 1897
rect 15528 1869 15613 1877
rect 15637 1893 15675 1902
rect 15637 1873 15646 1893
rect 15666 1873 15675 1893
rect 15528 1868 15564 1869
rect 15637 1865 15675 1873
rect 15741 1897 15826 1903
rect 15846 1902 15883 1903
rect 15741 1877 15749 1897
rect 15769 1896 15826 1897
rect 15769 1877 15798 1896
rect 15741 1876 15798 1877
rect 15819 1876 15826 1896
rect 15741 1869 15826 1876
rect 15845 1893 15883 1902
rect 15845 1873 15854 1893
rect 15874 1873 15883 1893
rect 15741 1868 15777 1869
rect 15845 1865 15883 1873
rect 15949 1897 16093 1903
rect 15949 1877 15957 1897
rect 15977 1894 16065 1897
rect 15977 1877 16008 1894
rect 15949 1874 16008 1877
rect 16031 1877 16065 1894
rect 16085 1877 16093 1897
rect 16031 1874 16093 1877
rect 15949 1869 16093 1874
rect 15949 1868 15985 1869
rect 16057 1868 16093 1869
rect 16159 1902 16196 1903
rect 16159 1901 16197 1902
rect 16159 1893 16223 1901
rect 16159 1873 16168 1893
rect 16188 1879 16223 1893
rect 16243 1879 16246 1899
rect 16188 1874 16246 1879
rect 16188 1873 16223 1874
rect 15425 1836 15462 1865
rect 15426 1834 15462 1836
rect 15638 1834 15675 1865
rect 15426 1812 15675 1834
rect 15846 1833 15883 1865
rect 16159 1861 16223 1873
rect 16263 1835 16290 2013
rect 18818 1991 18845 2169
rect 18885 2131 18949 2143
rect 19225 2139 19262 2171
rect 19433 2170 19682 2192
rect 19723 2171 19909 2203
rect 19737 2170 19909 2171
rect 19433 2139 19470 2170
rect 19646 2168 19682 2170
rect 19646 2139 19683 2168
rect 19875 2142 19909 2170
rect 18885 2130 18920 2131
rect 18862 2125 18920 2130
rect 18862 2105 18865 2125
rect 18885 2111 18920 2125
rect 18940 2111 18949 2131
rect 18885 2103 18949 2111
rect 18911 2102 18949 2103
rect 18912 2101 18949 2102
rect 19015 2135 19051 2136
rect 19123 2135 19159 2136
rect 19015 2128 19159 2135
rect 19015 2127 19075 2128
rect 19015 2107 19023 2127
rect 19043 2108 19075 2127
rect 19100 2127 19159 2128
rect 19100 2108 19131 2127
rect 19043 2107 19131 2108
rect 19151 2107 19159 2127
rect 19015 2101 19159 2107
rect 19225 2131 19263 2139
rect 19331 2135 19367 2136
rect 19225 2111 19234 2131
rect 19254 2111 19263 2131
rect 19225 2102 19263 2111
rect 19282 2128 19367 2135
rect 19282 2108 19289 2128
rect 19310 2127 19367 2128
rect 19310 2108 19339 2127
rect 19282 2107 19339 2108
rect 19359 2107 19367 2127
rect 19225 2101 19262 2102
rect 19282 2101 19367 2107
rect 19433 2131 19471 2139
rect 19544 2135 19580 2136
rect 19433 2111 19442 2131
rect 19462 2111 19471 2131
rect 19433 2102 19471 2111
rect 19495 2127 19580 2135
rect 19495 2107 19552 2127
rect 19572 2107 19580 2127
rect 19433 2101 19470 2102
rect 19495 2101 19580 2107
rect 19646 2131 19684 2139
rect 19646 2111 19655 2131
rect 19675 2111 19684 2131
rect 19646 2102 19684 2111
rect 19873 2132 19910 2142
rect 19873 2114 19883 2132
rect 19901 2114 19910 2132
rect 19873 2105 19910 2114
rect 19875 2104 19909 2105
rect 19646 2101 19683 2102
rect 19069 2080 19105 2101
rect 19495 2080 19526 2101
rect 18902 2076 19002 2080
rect 18902 2072 18964 2076
rect 18902 2046 18909 2072
rect 18935 2050 18964 2072
rect 18990 2050 19002 2076
rect 18935 2046 19002 2050
rect 18902 2043 19002 2046
rect 19070 2043 19105 2080
rect 19167 2077 19526 2080
rect 19167 2072 19389 2077
rect 19167 2048 19180 2072
rect 19204 2053 19389 2072
rect 19413 2053 19526 2077
rect 19204 2048 19526 2053
rect 19167 2044 19526 2048
rect 19593 2072 19742 2080
rect 19593 2052 19604 2072
rect 19624 2052 19742 2072
rect 19593 2045 19742 2052
rect 19593 2044 19634 2045
rect 18917 1991 18954 1992
rect 19013 1991 19050 1992
rect 19069 1991 19105 2043
rect 19124 1991 19161 1992
rect 18817 1982 18955 1991
rect 18412 1961 18523 1976
rect 18412 1959 18454 1961
rect 18082 1938 18187 1940
rect 17740 1930 17908 1931
rect 18082 1930 18131 1938
rect 17740 1911 18131 1930
rect 18162 1911 18187 1938
rect 18412 1939 18419 1959
rect 18438 1939 18454 1959
rect 18412 1931 18454 1939
rect 18482 1959 18523 1961
rect 18482 1939 18496 1959
rect 18515 1939 18523 1959
rect 18817 1962 18926 1982
rect 18946 1962 18955 1982
rect 18817 1955 18955 1962
rect 19013 1982 19161 1991
rect 19013 1962 19022 1982
rect 19042 1962 19132 1982
rect 19152 1962 19161 1982
rect 18817 1953 18913 1955
rect 19013 1952 19161 1962
rect 19220 1982 19257 1992
rect 19332 1991 19369 1992
rect 19313 1989 19369 1991
rect 19220 1962 19228 1982
rect 19248 1962 19257 1982
rect 19069 1951 19105 1952
rect 18482 1931 18523 1939
rect 18412 1925 18523 1931
rect 17740 1904 18187 1911
rect 17740 1902 17908 1904
rect 16588 1871 16698 1885
rect 16588 1868 16631 1871
rect 16588 1863 16592 1868
rect 16122 1833 16290 1835
rect 15846 1830 16290 1833
rect 15507 1806 15618 1812
rect 15507 1798 15548 1806
rect 15196 1743 15235 1787
rect 15507 1778 15515 1798
rect 15534 1778 15548 1798
rect 15507 1776 15548 1778
rect 15576 1798 15618 1806
rect 15576 1778 15592 1798
rect 15611 1778 15618 1798
rect 15576 1776 15618 1778
rect 15507 1761 15618 1776
rect 15844 1807 16290 1830
rect 15196 1719 15236 1743
rect 15536 1719 15583 1721
rect 15844 1719 15882 1807
rect 16122 1806 16290 1807
rect 16510 1841 16592 1863
rect 16621 1841 16631 1868
rect 16659 1844 16666 1871
rect 16695 1863 16698 1871
rect 16695 1844 16760 1863
rect 16659 1841 16760 1844
rect 16510 1839 16760 1841
rect 16510 1760 16547 1839
rect 16588 1826 16698 1839
rect 16662 1770 16693 1771
rect 16510 1740 16519 1760
rect 16539 1740 16547 1760
rect 16510 1730 16547 1740
rect 16606 1760 16693 1770
rect 16606 1740 16615 1760
rect 16635 1740 16693 1760
rect 16606 1731 16693 1740
rect 16606 1730 16643 1731
rect 15196 1686 15882 1719
rect 15196 1629 15235 1686
rect 15844 1684 15882 1686
rect 16662 1678 16693 1731
rect 16723 1760 16760 1839
rect 16931 1852 17324 1856
rect 16931 1835 16950 1852
rect 16970 1836 17324 1852
rect 17344 1836 17347 1856
rect 16970 1835 17347 1836
rect 16931 1831 17347 1835
rect 16931 1830 17272 1831
rect 16875 1770 16906 1771
rect 16723 1740 16732 1760
rect 16752 1740 16760 1760
rect 16723 1730 16760 1740
rect 16819 1763 16906 1770
rect 16819 1760 16880 1763
rect 16819 1740 16828 1760
rect 16848 1743 16880 1760
rect 16901 1743 16906 1763
rect 16848 1740 16906 1743
rect 16819 1733 16906 1740
rect 16931 1760 16968 1830
rect 17234 1829 17271 1830
rect 17083 1770 17119 1771
rect 16931 1740 16940 1760
rect 16960 1740 16968 1760
rect 16819 1731 16875 1733
rect 16819 1730 16856 1731
rect 16931 1730 16968 1740
rect 17027 1760 17175 1770
rect 17343 1769 17372 1770
rect 17275 1767 17372 1769
rect 17027 1740 17036 1760
rect 17056 1756 17146 1760
rect 17056 1740 17089 1756
rect 17027 1731 17089 1740
rect 17027 1730 17064 1731
rect 17083 1718 17089 1731
rect 17112 1740 17146 1756
rect 17166 1740 17175 1760
rect 17112 1731 17175 1740
rect 17233 1760 17372 1767
rect 17233 1740 17242 1760
rect 17262 1740 17372 1760
rect 17233 1731 17372 1740
rect 17112 1718 17119 1731
rect 17138 1730 17175 1731
rect 17234 1730 17271 1731
rect 17083 1679 17119 1718
rect 16554 1677 16595 1678
rect 16446 1670 16595 1677
rect 16446 1650 16564 1670
rect 16584 1650 16595 1670
rect 16446 1642 16595 1650
rect 16662 1674 17021 1678
rect 16662 1669 16984 1674
rect 16662 1645 16775 1669
rect 16799 1650 16984 1669
rect 17008 1650 17021 1674
rect 16799 1645 17021 1650
rect 16662 1642 17021 1645
rect 17083 1642 17118 1679
rect 17186 1676 17286 1679
rect 17186 1672 17253 1676
rect 17186 1646 17198 1672
rect 17224 1650 17253 1672
rect 17279 1650 17286 1676
rect 17224 1646 17286 1650
rect 17186 1642 17286 1646
rect 15196 1627 15244 1629
rect 15196 1609 15207 1627
rect 15225 1609 15244 1627
rect 16662 1621 16693 1642
rect 17083 1621 17119 1642
rect 16505 1620 16542 1621
rect 15196 1600 15244 1609
rect 15197 1599 15244 1600
rect 15510 1604 15620 1618
rect 15510 1601 15553 1604
rect 15510 1596 15514 1601
rect 15432 1574 15514 1596
rect 15543 1574 15553 1601
rect 15581 1577 15588 1604
rect 15617 1596 15620 1604
rect 16504 1611 16542 1620
rect 15617 1577 15682 1596
rect 16504 1591 16513 1611
rect 16533 1591 16542 1611
rect 15581 1574 15682 1577
rect 15432 1572 15682 1574
rect 15200 1536 15237 1537
rect 14818 1429 14828 1447
rect 14846 1429 14858 1447
rect 14818 1424 14858 1429
rect 15196 1533 15237 1536
rect 15196 1528 15238 1533
rect 15196 1510 15209 1528
rect 15227 1510 15238 1528
rect 15196 1496 15238 1510
rect 15276 1496 15323 1500
rect 15196 1490 15323 1496
rect 15196 1461 15284 1490
rect 15313 1461 15323 1490
rect 15432 1493 15469 1572
rect 15510 1559 15620 1572
rect 15584 1503 15615 1504
rect 15432 1473 15441 1493
rect 15461 1473 15469 1493
rect 15432 1463 15469 1473
rect 15528 1493 15615 1503
rect 15528 1473 15537 1493
rect 15557 1473 15615 1493
rect 15528 1464 15615 1473
rect 15528 1463 15565 1464
rect 15196 1457 15323 1461
rect 15196 1440 15235 1457
rect 15276 1456 15323 1457
rect 14818 1420 14855 1424
rect 15196 1422 15207 1440
rect 15225 1422 15235 1440
rect 15196 1413 15235 1422
rect 15197 1412 15234 1413
rect 15584 1411 15615 1464
rect 15645 1493 15682 1572
rect 15853 1569 16246 1589
rect 16266 1569 16269 1589
rect 16504 1583 16542 1591
rect 16608 1615 16693 1621
rect 16718 1620 16755 1621
rect 16608 1595 16616 1615
rect 16636 1595 16693 1615
rect 16608 1587 16693 1595
rect 16717 1611 16755 1620
rect 16717 1591 16726 1611
rect 16746 1591 16755 1611
rect 16608 1586 16644 1587
rect 16717 1583 16755 1591
rect 16821 1615 16906 1621
rect 16926 1620 16963 1621
rect 16821 1595 16829 1615
rect 16849 1614 16906 1615
rect 16849 1595 16878 1614
rect 16821 1594 16878 1595
rect 16899 1594 16906 1614
rect 16821 1587 16906 1594
rect 16925 1611 16963 1620
rect 16925 1591 16934 1611
rect 16954 1591 16963 1611
rect 16821 1586 16857 1587
rect 16925 1583 16963 1591
rect 17029 1615 17173 1621
rect 17029 1595 17037 1615
rect 17057 1595 17145 1615
rect 17165 1595 17173 1615
rect 17029 1587 17173 1595
rect 17029 1586 17065 1587
rect 17137 1586 17173 1587
rect 17239 1620 17276 1621
rect 17239 1619 17277 1620
rect 17239 1611 17303 1619
rect 17239 1591 17248 1611
rect 17268 1597 17303 1611
rect 17323 1597 17326 1617
rect 17268 1592 17326 1597
rect 17268 1591 17303 1592
rect 15853 1564 16269 1569
rect 15853 1563 16194 1564
rect 15797 1503 15828 1504
rect 15645 1473 15654 1493
rect 15674 1473 15682 1493
rect 15645 1463 15682 1473
rect 15741 1496 15828 1503
rect 15741 1493 15802 1496
rect 15741 1473 15750 1493
rect 15770 1476 15802 1493
rect 15823 1476 15828 1496
rect 15770 1473 15828 1476
rect 15741 1466 15828 1473
rect 15853 1493 15890 1563
rect 16156 1562 16193 1563
rect 16505 1554 16542 1583
rect 16506 1552 16542 1554
rect 16718 1552 16755 1583
rect 16506 1530 16755 1552
rect 16926 1551 16963 1583
rect 17239 1579 17303 1591
rect 17343 1553 17372 1731
rect 17740 1724 17767 1902
rect 17807 1864 17871 1876
rect 18147 1872 18184 1904
rect 18355 1903 18604 1925
rect 18355 1872 18392 1903
rect 18568 1901 18604 1903
rect 18568 1872 18605 1901
rect 18917 1892 18954 1893
rect 19220 1892 19257 1962
rect 19282 1982 19369 1989
rect 19282 1979 19340 1982
rect 19282 1959 19287 1979
rect 19308 1962 19340 1979
rect 19360 1962 19369 1982
rect 19308 1959 19369 1962
rect 19282 1952 19369 1959
rect 19428 1982 19465 1992
rect 19428 1962 19436 1982
rect 19456 1962 19465 1982
rect 19282 1951 19313 1952
rect 18916 1891 19257 1892
rect 18841 1886 19257 1891
rect 17807 1863 17842 1864
rect 17784 1858 17842 1863
rect 17784 1838 17787 1858
rect 17807 1844 17842 1858
rect 17862 1844 17871 1864
rect 17807 1836 17871 1844
rect 17833 1835 17871 1836
rect 17834 1834 17871 1835
rect 17937 1868 17973 1869
rect 18045 1868 18081 1869
rect 17937 1863 18081 1868
rect 17937 1860 17997 1863
rect 17937 1840 17945 1860
rect 17965 1842 17997 1860
rect 18024 1860 18081 1863
rect 18024 1842 18053 1860
rect 17965 1840 18053 1842
rect 18073 1840 18081 1860
rect 17937 1834 18081 1840
rect 18147 1864 18185 1872
rect 18253 1868 18289 1869
rect 18147 1844 18156 1864
rect 18176 1844 18185 1864
rect 18147 1835 18185 1844
rect 18204 1861 18289 1868
rect 18204 1841 18211 1861
rect 18232 1860 18289 1861
rect 18232 1841 18261 1860
rect 18204 1840 18261 1841
rect 18281 1840 18289 1860
rect 18147 1834 18184 1835
rect 18204 1834 18289 1840
rect 18355 1864 18393 1872
rect 18466 1868 18502 1869
rect 18355 1844 18364 1864
rect 18384 1844 18393 1864
rect 18355 1835 18393 1844
rect 18417 1860 18502 1868
rect 18417 1840 18474 1860
rect 18494 1840 18502 1860
rect 18355 1834 18392 1835
rect 18417 1834 18502 1840
rect 18568 1864 18606 1872
rect 18841 1866 18844 1886
rect 18864 1866 19257 1886
rect 19428 1883 19465 1962
rect 19495 1991 19526 2044
rect 19876 2042 19913 2043
rect 19875 2033 19914 2042
rect 19875 2015 19885 2033
rect 19903 2015 19914 2033
rect 19787 1998 19834 1999
rect 19875 1998 19914 2015
rect 19787 1994 19914 1998
rect 19545 1991 19582 1992
rect 19495 1982 19582 1991
rect 19495 1962 19553 1982
rect 19573 1962 19582 1982
rect 19495 1952 19582 1962
rect 19641 1982 19678 1992
rect 19641 1962 19649 1982
rect 19669 1962 19678 1982
rect 19495 1951 19526 1952
rect 19490 1883 19600 1896
rect 19641 1883 19678 1962
rect 19787 1965 19797 1994
rect 19826 1965 19914 1994
rect 19787 1959 19914 1965
rect 19787 1955 19834 1959
rect 19872 1945 19914 1959
rect 19872 1927 19883 1945
rect 19901 1927 19914 1945
rect 19872 1922 19914 1927
rect 19873 1919 19914 1922
rect 19873 1918 19910 1919
rect 19428 1881 19678 1883
rect 19428 1878 19529 1881
rect 18568 1844 18577 1864
rect 18597 1844 18606 1864
rect 19428 1859 19493 1878
rect 18568 1835 18606 1844
rect 19490 1851 19493 1859
rect 19522 1851 19529 1878
rect 19557 1854 19567 1881
rect 19596 1859 19678 1881
rect 19596 1854 19600 1859
rect 19557 1851 19600 1854
rect 19490 1837 19600 1851
rect 19866 1855 19913 1856
rect 19866 1846 19914 1855
rect 18568 1834 18605 1835
rect 17991 1813 18027 1834
rect 18417 1813 18448 1834
rect 19866 1828 19885 1846
rect 19903 1828 19914 1846
rect 19866 1826 19914 1828
rect 17824 1809 17924 1813
rect 17824 1805 17886 1809
rect 17824 1779 17831 1805
rect 17857 1783 17886 1805
rect 17912 1783 17924 1809
rect 17857 1779 17924 1783
rect 17824 1776 17924 1779
rect 17992 1776 18027 1813
rect 18089 1810 18448 1813
rect 18089 1805 18311 1810
rect 18089 1781 18102 1805
rect 18126 1786 18311 1805
rect 18335 1786 18448 1810
rect 18126 1781 18448 1786
rect 18089 1777 18448 1781
rect 18515 1805 18664 1813
rect 18515 1785 18526 1805
rect 18546 1785 18664 1805
rect 18515 1778 18664 1785
rect 18515 1777 18556 1778
rect 17839 1724 17876 1725
rect 17935 1724 17972 1725
rect 17991 1724 18027 1776
rect 18046 1724 18083 1725
rect 17739 1715 17877 1724
rect 17739 1695 17848 1715
rect 17868 1695 17877 1715
rect 17739 1688 17877 1695
rect 17935 1715 18083 1724
rect 17935 1695 17944 1715
rect 17964 1695 18054 1715
rect 18074 1695 18083 1715
rect 17739 1686 17835 1688
rect 17935 1685 18083 1695
rect 18142 1715 18179 1725
rect 18254 1724 18291 1725
rect 18235 1722 18291 1724
rect 18142 1695 18150 1715
rect 18170 1695 18179 1715
rect 17991 1684 18027 1685
rect 17839 1625 17876 1626
rect 18142 1625 18179 1695
rect 18204 1715 18291 1722
rect 18204 1712 18262 1715
rect 18204 1692 18209 1712
rect 18230 1695 18262 1712
rect 18282 1695 18291 1715
rect 18230 1692 18291 1695
rect 18204 1685 18291 1692
rect 18350 1715 18387 1725
rect 18350 1695 18358 1715
rect 18378 1695 18387 1715
rect 18204 1684 18235 1685
rect 17838 1624 18179 1625
rect 17763 1620 18179 1624
rect 17763 1619 18140 1620
rect 17763 1599 17766 1619
rect 17786 1603 18140 1619
rect 18160 1603 18179 1620
rect 17786 1599 18179 1603
rect 18350 1616 18387 1695
rect 18417 1724 18448 1777
rect 19228 1769 19266 1771
rect 19875 1769 19914 1826
rect 19228 1736 19914 1769
rect 18467 1724 18504 1725
rect 18417 1715 18504 1724
rect 18417 1695 18475 1715
rect 18495 1695 18504 1715
rect 18417 1685 18504 1695
rect 18563 1715 18600 1725
rect 18563 1695 18571 1715
rect 18591 1695 18600 1715
rect 18417 1684 18448 1685
rect 18412 1616 18522 1629
rect 18563 1616 18600 1695
rect 18350 1614 18600 1616
rect 18350 1611 18451 1614
rect 18350 1592 18415 1611
rect 18412 1584 18415 1592
rect 18444 1584 18451 1611
rect 18479 1587 18489 1614
rect 18518 1592 18600 1614
rect 18820 1648 18988 1649
rect 19228 1648 19266 1736
rect 19527 1734 19574 1736
rect 19874 1712 19914 1736
rect 18820 1625 19266 1648
rect 19492 1679 19603 1694
rect 19492 1677 19534 1679
rect 19492 1657 19499 1677
rect 19518 1657 19534 1677
rect 19492 1649 19534 1657
rect 19562 1677 19603 1679
rect 19562 1657 19576 1677
rect 19595 1657 19603 1677
rect 19875 1668 19914 1712
rect 19562 1649 19603 1657
rect 19492 1643 19603 1649
rect 18820 1622 19264 1625
rect 18820 1620 18988 1622
rect 18518 1587 18522 1592
rect 18479 1584 18522 1587
rect 18412 1570 18522 1584
rect 17202 1551 17372 1553
rect 16923 1544 17372 1551
rect 16587 1524 16698 1530
rect 16587 1516 16628 1524
rect 16005 1503 16041 1504
rect 15853 1473 15862 1493
rect 15882 1473 15890 1493
rect 15741 1464 15797 1466
rect 15741 1463 15778 1464
rect 15853 1463 15890 1473
rect 15949 1493 16097 1503
rect 16197 1500 16293 1502
rect 15949 1473 15958 1493
rect 15978 1473 16068 1493
rect 16088 1473 16097 1493
rect 15949 1464 16097 1473
rect 16155 1493 16293 1500
rect 16155 1473 16164 1493
rect 16184 1473 16293 1493
rect 16587 1496 16595 1516
rect 16614 1496 16628 1516
rect 16587 1494 16628 1496
rect 16656 1516 16698 1524
rect 16656 1496 16672 1516
rect 16691 1496 16698 1516
rect 16923 1517 16948 1544
rect 16979 1525 17372 1544
rect 16979 1517 17028 1525
rect 17202 1524 17372 1525
rect 16923 1515 17028 1517
rect 16656 1494 16698 1496
rect 16587 1479 16698 1494
rect 16155 1464 16293 1473
rect 15949 1463 15986 1464
rect 16005 1412 16041 1464
rect 16060 1463 16097 1464
rect 16156 1463 16193 1464
rect 15476 1410 15517 1411
rect 15368 1403 15517 1410
rect 14491 1401 14528 1402
rect 14441 1392 14528 1401
rect 14441 1372 14499 1392
rect 14519 1372 14528 1392
rect 14441 1362 14528 1372
rect 14587 1392 14624 1402
rect 14587 1372 14595 1392
rect 14615 1372 14624 1392
rect 15368 1383 15486 1403
rect 15506 1383 15517 1403
rect 15368 1375 15517 1383
rect 15584 1407 15943 1411
rect 15584 1402 15906 1407
rect 15584 1378 15697 1402
rect 15721 1383 15906 1402
rect 15930 1383 15943 1407
rect 15721 1378 15943 1383
rect 15584 1375 15943 1378
rect 16005 1375 16040 1412
rect 16108 1409 16208 1412
rect 16108 1405 16175 1409
rect 16108 1379 16120 1405
rect 16146 1383 16175 1405
rect 16201 1383 16208 1409
rect 16146 1379 16208 1383
rect 16108 1375 16208 1379
rect 14441 1361 14472 1362
rect 14436 1293 14546 1306
rect 14587 1293 14624 1372
rect 14821 1357 14858 1358
rect 14817 1348 14858 1357
rect 15584 1354 15615 1375
rect 16005 1354 16041 1375
rect 15427 1353 15464 1354
rect 15201 1350 15235 1351
rect 14817 1330 14830 1348
rect 14848 1330 14858 1348
rect 14817 1321 14858 1330
rect 15200 1341 15237 1350
rect 15200 1323 15209 1341
rect 15227 1323 15237 1341
rect 14817 1301 14857 1321
rect 15200 1313 15237 1323
rect 15426 1344 15464 1353
rect 15426 1324 15435 1344
rect 15455 1324 15464 1344
rect 15426 1316 15464 1324
rect 15530 1348 15615 1354
rect 15640 1353 15677 1354
rect 15530 1328 15538 1348
rect 15558 1328 15615 1348
rect 15530 1320 15615 1328
rect 15639 1344 15677 1353
rect 15639 1324 15648 1344
rect 15668 1324 15677 1344
rect 15530 1319 15566 1320
rect 15639 1316 15677 1324
rect 15743 1348 15828 1354
rect 15848 1353 15885 1354
rect 15743 1328 15751 1348
rect 15771 1347 15828 1348
rect 15771 1328 15800 1347
rect 15743 1327 15800 1328
rect 15821 1327 15828 1347
rect 15743 1320 15828 1327
rect 15847 1344 15885 1353
rect 15847 1324 15856 1344
rect 15876 1324 15885 1344
rect 15743 1319 15779 1320
rect 15847 1316 15885 1324
rect 15951 1348 16095 1354
rect 15951 1328 15959 1348
rect 15979 1347 16067 1348
rect 15979 1328 16010 1347
rect 15951 1327 16010 1328
rect 16035 1328 16067 1347
rect 16087 1328 16095 1348
rect 16035 1327 16095 1328
rect 15951 1320 16095 1327
rect 15951 1319 15987 1320
rect 16059 1319 16095 1320
rect 16161 1353 16198 1354
rect 16161 1352 16199 1353
rect 16161 1344 16225 1352
rect 16161 1324 16170 1344
rect 16190 1330 16225 1344
rect 16245 1330 16248 1350
rect 16190 1325 16248 1330
rect 16190 1324 16225 1325
rect 14374 1291 14624 1293
rect 14374 1288 14475 1291
rect 12892 1231 12956 1243
rect 13232 1239 13269 1266
rect 13440 1239 13477 1270
rect 13653 1268 13689 1270
rect 14374 1269 14439 1288
rect 13653 1239 13690 1268
rect 14436 1261 14439 1269
rect 14468 1261 14475 1288
rect 14503 1264 14513 1291
rect 14542 1269 14624 1291
rect 14732 1291 14857 1301
rect 14732 1272 14740 1291
rect 14765 1272 14857 1291
rect 14542 1264 14546 1269
rect 14732 1265 14857 1272
rect 14503 1261 14546 1264
rect 14436 1247 14546 1261
rect 12892 1230 12927 1231
rect 12869 1225 12927 1230
rect 12869 1205 12872 1225
rect 12892 1211 12927 1225
rect 12947 1211 12956 1231
rect 12892 1203 12956 1211
rect 12918 1202 12956 1203
rect 12919 1201 12956 1202
rect 13022 1235 13058 1236
rect 13130 1235 13166 1236
rect 13022 1227 13166 1235
rect 13022 1207 13030 1227
rect 13050 1224 13138 1227
rect 13050 1207 13082 1224
rect 13102 1207 13138 1224
rect 13158 1207 13166 1227
rect 13022 1201 13166 1207
rect 13232 1231 13270 1239
rect 13338 1235 13374 1236
rect 13232 1211 13241 1231
rect 13261 1211 13270 1231
rect 13232 1202 13270 1211
rect 13289 1228 13374 1235
rect 13289 1208 13296 1228
rect 13317 1227 13374 1228
rect 13317 1208 13346 1227
rect 13289 1207 13346 1208
rect 13366 1207 13374 1227
rect 13232 1201 13269 1202
rect 13289 1201 13374 1207
rect 13440 1231 13478 1239
rect 13551 1235 13587 1236
rect 13440 1211 13449 1231
rect 13469 1211 13478 1231
rect 13440 1202 13478 1211
rect 13502 1227 13587 1235
rect 13502 1207 13559 1227
rect 13579 1207 13587 1227
rect 13440 1201 13477 1202
rect 13502 1201 13587 1207
rect 13653 1231 13691 1239
rect 13653 1211 13662 1231
rect 13682 1211 13691 1231
rect 13653 1202 13691 1211
rect 14817 1217 14857 1265
rect 15201 1285 15235 1313
rect 15427 1287 15464 1316
rect 15428 1285 15464 1287
rect 15640 1285 15677 1316
rect 15201 1284 15373 1285
rect 15201 1252 15387 1284
rect 15428 1263 15677 1285
rect 15848 1284 15885 1316
rect 16161 1312 16225 1324
rect 16265 1286 16292 1464
rect 18820 1442 18847 1620
rect 18887 1582 18951 1594
rect 19227 1590 19264 1622
rect 19435 1621 19684 1643
rect 19435 1590 19472 1621
rect 19648 1619 19684 1621
rect 19648 1590 19685 1619
rect 18887 1581 18922 1582
rect 18864 1576 18922 1581
rect 18864 1556 18867 1576
rect 18887 1562 18922 1576
rect 18942 1562 18951 1582
rect 18887 1554 18951 1562
rect 18913 1553 18951 1554
rect 18914 1552 18951 1553
rect 19017 1586 19053 1587
rect 19125 1586 19161 1587
rect 19017 1581 19161 1586
rect 19017 1578 19079 1581
rect 19017 1558 19025 1578
rect 19045 1561 19079 1578
rect 19102 1578 19161 1581
rect 19102 1561 19133 1578
rect 19045 1558 19133 1561
rect 19153 1558 19161 1578
rect 19017 1552 19161 1558
rect 19227 1582 19265 1590
rect 19333 1586 19369 1587
rect 19227 1562 19236 1582
rect 19256 1562 19265 1582
rect 19227 1553 19265 1562
rect 19284 1579 19369 1586
rect 19284 1559 19291 1579
rect 19312 1578 19369 1579
rect 19312 1559 19341 1578
rect 19284 1558 19341 1559
rect 19361 1558 19369 1578
rect 19227 1552 19264 1553
rect 19284 1552 19369 1558
rect 19435 1582 19473 1590
rect 19546 1586 19582 1587
rect 19435 1562 19444 1582
rect 19464 1562 19473 1582
rect 19435 1553 19473 1562
rect 19497 1578 19582 1586
rect 19497 1558 19554 1578
rect 19574 1558 19582 1578
rect 19435 1552 19472 1553
rect 19497 1552 19582 1558
rect 19648 1582 19686 1590
rect 19648 1562 19657 1582
rect 19677 1562 19686 1582
rect 19648 1553 19686 1562
rect 19648 1552 19685 1553
rect 19071 1531 19107 1552
rect 19497 1531 19528 1552
rect 18904 1527 19004 1531
rect 18904 1523 18966 1527
rect 18904 1497 18911 1523
rect 18937 1501 18966 1523
rect 18992 1501 19004 1527
rect 18937 1497 19004 1501
rect 18904 1494 19004 1497
rect 19072 1494 19107 1531
rect 19169 1528 19528 1531
rect 19169 1523 19391 1528
rect 19169 1499 19182 1523
rect 19206 1504 19391 1523
rect 19415 1504 19528 1528
rect 19206 1499 19528 1504
rect 19169 1495 19528 1499
rect 19595 1523 19744 1531
rect 19595 1503 19606 1523
rect 19626 1503 19744 1523
rect 19595 1496 19744 1503
rect 19595 1495 19636 1496
rect 18919 1442 18956 1443
rect 19015 1442 19052 1443
rect 19071 1442 19107 1494
rect 19126 1442 19163 1443
rect 18819 1433 18957 1442
rect 18819 1413 18928 1433
rect 18948 1413 18957 1433
rect 18819 1406 18957 1413
rect 19015 1433 19163 1442
rect 19015 1413 19024 1433
rect 19044 1413 19134 1433
rect 19154 1413 19163 1433
rect 18819 1404 18915 1406
rect 19015 1403 19163 1413
rect 19222 1433 19259 1443
rect 19334 1442 19371 1443
rect 19315 1440 19371 1442
rect 19222 1413 19230 1433
rect 19250 1413 19259 1433
rect 19071 1402 19107 1403
rect 16448 1360 16558 1374
rect 16448 1357 16491 1360
rect 16448 1352 16452 1357
rect 16124 1284 16292 1286
rect 15848 1278 16292 1284
rect 15201 1220 15235 1252
rect 13653 1201 13690 1202
rect 13076 1180 13112 1201
rect 13502 1180 13533 1201
rect 14817 1199 14828 1217
rect 14846 1199 14857 1217
rect 14817 1191 14857 1199
rect 15197 1211 15235 1220
rect 15197 1193 15207 1211
rect 15225 1193 15235 1211
rect 14818 1190 14855 1191
rect 15197 1187 15235 1193
rect 15353 1189 15387 1252
rect 15509 1257 15620 1263
rect 15509 1249 15550 1257
rect 15509 1229 15517 1249
rect 15536 1229 15550 1249
rect 15509 1227 15550 1229
rect 15578 1249 15620 1257
rect 15578 1229 15594 1249
rect 15613 1229 15620 1249
rect 15578 1227 15620 1229
rect 15509 1212 15620 1227
rect 15847 1258 16292 1278
rect 15847 1189 15885 1258
rect 16124 1257 16292 1258
rect 16370 1330 16452 1352
rect 16481 1330 16491 1357
rect 16519 1333 16526 1360
rect 16555 1352 16558 1360
rect 18553 1369 18664 1384
rect 18553 1367 18595 1369
rect 16555 1333 16620 1352
rect 16519 1330 16620 1333
rect 16370 1328 16620 1330
rect 16370 1249 16407 1328
rect 16448 1315 16558 1328
rect 16522 1259 16553 1260
rect 16370 1229 16379 1249
rect 16399 1229 16407 1249
rect 16370 1219 16407 1229
rect 16466 1249 16553 1259
rect 16466 1229 16475 1249
rect 16495 1229 16553 1249
rect 16466 1220 16553 1229
rect 16466 1219 16503 1220
rect 15197 1183 15234 1187
rect 12909 1176 13009 1180
rect 12909 1172 12971 1176
rect 12909 1146 12916 1172
rect 12942 1150 12971 1172
rect 12997 1150 13009 1176
rect 12942 1146 13009 1150
rect 12909 1143 13009 1146
rect 13077 1143 13112 1180
rect 13174 1177 13533 1180
rect 13174 1172 13396 1177
rect 13174 1148 13187 1172
rect 13211 1153 13396 1172
rect 13420 1153 13533 1177
rect 13211 1148 13533 1153
rect 13174 1144 13533 1148
rect 13600 1172 13749 1180
rect 15353 1178 15885 1189
rect 13600 1152 13611 1172
rect 13631 1152 13749 1172
rect 15352 1162 15885 1178
rect 16522 1167 16553 1220
rect 16583 1249 16620 1328
rect 16791 1338 17184 1345
rect 16791 1321 16799 1338
rect 16831 1325 17184 1338
rect 17204 1325 17207 1345
rect 18286 1340 18327 1349
rect 16831 1321 17207 1325
rect 16791 1320 17207 1321
rect 17881 1338 18049 1339
rect 18286 1338 18295 1340
rect 16791 1319 17132 1320
rect 16735 1259 16766 1260
rect 16583 1229 16592 1249
rect 16612 1229 16620 1249
rect 16583 1219 16620 1229
rect 16679 1252 16766 1259
rect 16679 1249 16740 1252
rect 16679 1229 16688 1249
rect 16708 1232 16740 1249
rect 16761 1232 16766 1252
rect 16708 1229 16766 1232
rect 16679 1222 16766 1229
rect 16791 1249 16828 1319
rect 17094 1318 17131 1319
rect 17881 1318 18295 1338
rect 18321 1318 18327 1340
rect 18553 1347 18560 1367
rect 18579 1347 18595 1367
rect 18553 1339 18595 1347
rect 18623 1367 18664 1369
rect 18623 1347 18637 1367
rect 18656 1347 18664 1367
rect 18623 1339 18664 1347
rect 18919 1343 18956 1344
rect 19222 1343 19259 1413
rect 19284 1433 19371 1440
rect 19284 1430 19342 1433
rect 19284 1410 19289 1430
rect 19310 1413 19342 1430
rect 19362 1413 19371 1433
rect 19310 1410 19371 1413
rect 19284 1403 19371 1410
rect 19430 1433 19467 1443
rect 19430 1413 19438 1433
rect 19458 1413 19467 1433
rect 19284 1402 19315 1403
rect 18918 1342 19259 1343
rect 18553 1333 18664 1339
rect 18843 1337 19259 1342
rect 17881 1312 18327 1318
rect 17881 1310 18049 1312
rect 16943 1259 16979 1260
rect 16791 1229 16800 1249
rect 16820 1229 16828 1249
rect 16679 1220 16735 1222
rect 16679 1219 16716 1220
rect 16791 1219 16828 1229
rect 16887 1249 17035 1259
rect 17135 1256 17231 1258
rect 16887 1229 16896 1249
rect 16916 1244 17006 1249
rect 16916 1229 16951 1244
rect 16887 1220 16951 1229
rect 16887 1219 16924 1220
rect 16943 1203 16951 1220
rect 16972 1229 17006 1244
rect 17026 1229 17035 1249
rect 16972 1220 17035 1229
rect 17093 1249 17231 1256
rect 17093 1229 17102 1249
rect 17122 1229 17231 1249
rect 17093 1220 17231 1229
rect 16972 1203 16979 1220
rect 16998 1219 17035 1220
rect 17094 1219 17131 1220
rect 16943 1168 16979 1203
rect 16414 1166 16455 1167
rect 15352 1161 15866 1162
rect 13600 1145 13749 1152
rect 16306 1159 16455 1166
rect 14189 1149 14703 1150
rect 13600 1144 13641 1145
rect 12924 1091 12961 1092
rect 13020 1091 13057 1092
rect 13076 1091 13112 1143
rect 13131 1091 13168 1092
rect 12824 1082 12962 1091
rect 12824 1062 12933 1082
rect 12953 1062 12962 1082
rect 12824 1055 12962 1062
rect 13020 1082 13168 1091
rect 13020 1062 13029 1082
rect 13049 1062 13139 1082
rect 13159 1062 13168 1082
rect 12824 1053 12920 1055
rect 13020 1052 13168 1062
rect 13227 1082 13264 1092
rect 13339 1091 13376 1092
rect 13320 1089 13376 1091
rect 13227 1062 13235 1082
rect 13255 1062 13264 1082
rect 13076 1051 13112 1052
rect 12006 999 12174 1001
rect 11728 993 12174 999
rect 10796 969 11212 974
rect 11391 972 11502 978
rect 10796 968 11137 969
rect 10740 908 10771 909
rect 10588 878 10597 898
rect 10617 878 10625 898
rect 10588 868 10625 878
rect 10684 901 10771 908
rect 10684 898 10745 901
rect 10684 878 10693 898
rect 10713 881 10745 898
rect 10766 881 10771 901
rect 10713 878 10771 881
rect 10684 871 10771 878
rect 10796 898 10833 968
rect 11099 967 11136 968
rect 11391 964 11432 972
rect 11391 944 11399 964
rect 11418 944 11432 964
rect 11391 942 11432 944
rect 11460 964 11502 972
rect 11460 944 11476 964
rect 11495 944 11502 964
rect 11728 971 11734 993
rect 11760 973 12174 993
rect 12924 992 12961 993
rect 13227 992 13264 1062
rect 13289 1082 13376 1089
rect 13289 1079 13347 1082
rect 13289 1059 13294 1079
rect 13315 1062 13347 1079
rect 13367 1062 13376 1082
rect 13315 1059 13376 1062
rect 13289 1052 13376 1059
rect 13435 1082 13472 1092
rect 13435 1062 13443 1082
rect 13463 1062 13472 1082
rect 13289 1051 13320 1052
rect 12923 991 13264 992
rect 11760 971 11769 973
rect 12006 972 12174 973
rect 12848 986 13264 991
rect 11728 962 11769 971
rect 12848 966 12851 986
rect 12871 966 13264 986
rect 13435 983 13472 1062
rect 13502 1091 13533 1144
rect 14170 1133 14703 1149
rect 16306 1139 16424 1159
rect 16444 1139 16455 1159
rect 14170 1122 14702 1133
rect 16306 1131 16455 1139
rect 16522 1163 16881 1167
rect 16522 1158 16844 1163
rect 16522 1134 16635 1158
rect 16659 1139 16844 1158
rect 16868 1139 16881 1163
rect 16659 1134 16881 1139
rect 16522 1131 16881 1134
rect 16943 1131 16978 1168
rect 17046 1165 17146 1168
rect 17046 1161 17113 1165
rect 17046 1135 17058 1161
rect 17084 1139 17113 1161
rect 17139 1139 17146 1165
rect 17084 1135 17146 1139
rect 17046 1131 17146 1135
rect 14821 1124 14858 1128
rect 13552 1091 13589 1092
rect 13502 1082 13589 1091
rect 13502 1062 13560 1082
rect 13580 1062 13589 1082
rect 13502 1052 13589 1062
rect 13648 1082 13685 1092
rect 13648 1062 13656 1082
rect 13676 1062 13685 1082
rect 13502 1051 13533 1052
rect 13497 983 13607 996
rect 13648 983 13685 1062
rect 13435 981 13685 983
rect 13435 978 13536 981
rect 13435 959 13500 978
rect 11460 942 11502 944
rect 11391 927 11502 942
rect 13497 951 13500 959
rect 13529 951 13536 978
rect 13564 954 13574 981
rect 13603 959 13685 981
rect 13763 1053 13931 1054
rect 14170 1053 14208 1122
rect 13763 1033 14208 1053
rect 14435 1084 14546 1099
rect 14435 1082 14477 1084
rect 14435 1062 14442 1082
rect 14461 1062 14477 1082
rect 14435 1054 14477 1062
rect 14505 1082 14546 1084
rect 14505 1062 14519 1082
rect 14538 1062 14546 1082
rect 14505 1054 14546 1062
rect 14435 1048 14546 1054
rect 14668 1059 14702 1122
rect 14820 1118 14858 1124
rect 15200 1120 15237 1121
rect 14820 1100 14830 1118
rect 14848 1100 14858 1118
rect 14820 1091 14858 1100
rect 15198 1112 15238 1120
rect 15198 1094 15209 1112
rect 15227 1094 15238 1112
rect 16522 1110 16553 1131
rect 16943 1110 16979 1131
rect 16365 1109 16402 1110
rect 14820 1059 14854 1091
rect 13763 1027 14207 1033
rect 13763 1025 13931 1027
rect 13603 954 13607 959
rect 13564 951 13607 954
rect 13497 937 13607 951
rect 10948 908 10984 909
rect 10796 878 10805 898
rect 10825 878 10833 898
rect 10684 869 10740 871
rect 10684 868 10721 869
rect 10796 868 10833 878
rect 10892 898 11040 908
rect 11140 905 11236 907
rect 10892 878 10901 898
rect 10921 878 11011 898
rect 11031 878 11040 898
rect 10892 869 11040 878
rect 11098 898 11236 905
rect 11098 878 11107 898
rect 11127 878 11236 898
rect 11098 869 11236 878
rect 10892 868 10929 869
rect 10948 817 10984 869
rect 11003 868 11040 869
rect 11099 868 11136 869
rect 10419 815 10460 816
rect 10311 808 10460 815
rect 10311 788 10429 808
rect 10449 788 10460 808
rect 10311 780 10460 788
rect 10527 812 10886 816
rect 10527 807 10849 812
rect 10527 783 10640 807
rect 10664 788 10849 807
rect 10873 788 10886 812
rect 10664 783 10886 788
rect 10527 780 10886 783
rect 10948 780 10983 817
rect 11051 814 11151 817
rect 11051 810 11118 814
rect 11051 784 11063 810
rect 11089 788 11118 810
rect 11144 788 11151 814
rect 11089 784 11151 788
rect 11051 780 11151 784
rect 10527 759 10558 780
rect 10948 759 10984 780
rect 10370 758 10407 759
rect 10369 749 10407 758
rect 10369 729 10378 749
rect 10398 729 10407 749
rect 10369 721 10407 729
rect 10473 753 10558 759
rect 10583 758 10620 759
rect 10473 733 10481 753
rect 10501 733 10558 753
rect 10473 725 10558 733
rect 10582 749 10620 758
rect 10582 729 10591 749
rect 10611 729 10620 749
rect 10473 724 10509 725
rect 10582 721 10620 729
rect 10686 753 10771 759
rect 10791 758 10828 759
rect 10686 733 10694 753
rect 10714 752 10771 753
rect 10714 733 10743 752
rect 10686 732 10743 733
rect 10764 732 10771 752
rect 10686 725 10771 732
rect 10790 749 10828 758
rect 10790 729 10799 749
rect 10819 729 10828 749
rect 10686 724 10722 725
rect 10790 721 10828 729
rect 10894 753 11038 759
rect 10894 733 10902 753
rect 10922 750 11010 753
rect 10922 733 10953 750
rect 10894 730 10953 733
rect 10976 733 11010 750
rect 11030 733 11038 753
rect 10976 730 11038 733
rect 10894 725 11038 730
rect 10894 724 10930 725
rect 11002 724 11038 725
rect 11104 758 11141 759
rect 11104 757 11142 758
rect 11104 749 11168 757
rect 11104 729 11113 749
rect 11133 735 11168 749
rect 11188 735 11191 755
rect 11133 730 11191 735
rect 11133 729 11168 730
rect 10370 692 10407 721
rect 10371 690 10407 692
rect 10583 690 10620 721
rect 10371 668 10620 690
rect 10791 689 10828 721
rect 11104 717 11168 729
rect 11208 691 11235 869
rect 13763 847 13790 1025
rect 13830 987 13894 999
rect 14170 995 14207 1027
rect 14378 1026 14627 1048
rect 14668 1027 14854 1059
rect 14682 1026 14854 1027
rect 14378 995 14415 1026
rect 14591 1024 14627 1026
rect 14591 995 14628 1024
rect 14820 998 14854 1026
rect 15198 1046 15238 1094
rect 16364 1100 16402 1109
rect 16364 1080 16373 1100
rect 16393 1080 16402 1100
rect 16364 1072 16402 1080
rect 16468 1104 16553 1110
rect 16578 1109 16615 1110
rect 16468 1084 16476 1104
rect 16496 1084 16553 1104
rect 16468 1076 16553 1084
rect 16577 1100 16615 1109
rect 16577 1080 16586 1100
rect 16606 1080 16615 1100
rect 16468 1075 16504 1076
rect 16577 1072 16615 1080
rect 16681 1104 16766 1110
rect 16786 1109 16823 1110
rect 16681 1084 16689 1104
rect 16709 1103 16766 1104
rect 16709 1084 16738 1103
rect 16681 1083 16738 1084
rect 16759 1083 16766 1103
rect 16681 1076 16766 1083
rect 16785 1100 16823 1109
rect 16785 1080 16794 1100
rect 16814 1080 16823 1100
rect 16681 1075 16717 1076
rect 16785 1072 16823 1080
rect 16889 1104 17033 1110
rect 16889 1084 16897 1104
rect 16917 1084 17005 1104
rect 17025 1084 17033 1104
rect 16889 1076 17033 1084
rect 16889 1075 16925 1076
rect 16997 1075 17033 1076
rect 17099 1109 17136 1110
rect 17099 1108 17137 1109
rect 17099 1100 17163 1108
rect 17099 1080 17108 1100
rect 17128 1086 17163 1100
rect 17183 1086 17186 1106
rect 17128 1081 17186 1086
rect 17128 1080 17163 1081
rect 15509 1050 15619 1064
rect 15509 1047 15552 1050
rect 15198 1039 15323 1046
rect 15509 1042 15513 1047
rect 15198 1020 15290 1039
rect 15315 1020 15323 1039
rect 15198 1010 15323 1020
rect 15431 1020 15513 1042
rect 15542 1020 15552 1047
rect 15580 1023 15587 1050
rect 15616 1042 15619 1050
rect 16365 1043 16402 1072
rect 15616 1023 15681 1042
rect 16366 1041 16402 1043
rect 16578 1041 16615 1072
rect 16786 1045 16823 1072
rect 17099 1068 17163 1080
rect 15580 1020 15681 1023
rect 15431 1018 15681 1020
rect 13830 986 13865 987
rect 13807 981 13865 986
rect 13807 961 13810 981
rect 13830 967 13865 981
rect 13885 967 13894 987
rect 13830 959 13894 967
rect 13856 958 13894 959
rect 13857 957 13894 958
rect 13960 991 13996 992
rect 14068 991 14104 992
rect 13960 984 14104 991
rect 13960 983 14020 984
rect 13960 963 13968 983
rect 13988 964 14020 983
rect 14045 983 14104 984
rect 14045 964 14076 983
rect 13988 963 14076 964
rect 14096 963 14104 983
rect 13960 957 14104 963
rect 14170 987 14208 995
rect 14276 991 14312 992
rect 14170 967 14179 987
rect 14199 967 14208 987
rect 14170 958 14208 967
rect 14227 984 14312 991
rect 14227 964 14234 984
rect 14255 983 14312 984
rect 14255 964 14284 983
rect 14227 963 14284 964
rect 14304 963 14312 983
rect 14170 957 14207 958
rect 14227 957 14312 963
rect 14378 987 14416 995
rect 14489 991 14525 992
rect 14378 967 14387 987
rect 14407 967 14416 987
rect 14378 958 14416 967
rect 14440 983 14525 991
rect 14440 963 14497 983
rect 14517 963 14525 983
rect 14378 957 14415 958
rect 14440 957 14525 963
rect 14591 987 14629 995
rect 14591 967 14600 987
rect 14620 967 14629 987
rect 14591 958 14629 967
rect 14818 988 14855 998
rect 15198 990 15238 1010
rect 14818 970 14828 988
rect 14846 970 14855 988
rect 14818 961 14855 970
rect 15197 981 15238 990
rect 15197 963 15207 981
rect 15225 963 15238 981
rect 14820 960 14854 961
rect 14591 957 14628 958
rect 14014 936 14050 957
rect 14440 936 14471 957
rect 15197 954 15238 963
rect 15197 953 15234 954
rect 15431 939 15468 1018
rect 15509 1005 15619 1018
rect 15583 949 15614 950
rect 13847 932 13947 936
rect 13847 928 13909 932
rect 13847 902 13854 928
rect 13880 906 13909 928
rect 13935 906 13947 932
rect 13880 902 13947 906
rect 13847 899 13947 902
rect 14015 899 14050 936
rect 14112 933 14471 936
rect 14112 928 14334 933
rect 14112 904 14125 928
rect 14149 909 14334 928
rect 14358 909 14471 933
rect 14149 904 14471 909
rect 14112 900 14471 904
rect 14538 928 14687 936
rect 14538 908 14549 928
rect 14569 908 14687 928
rect 15431 919 15440 939
rect 15460 919 15468 939
rect 15431 909 15468 919
rect 15527 939 15614 949
rect 15527 919 15536 939
rect 15556 919 15614 939
rect 15527 910 15614 919
rect 15527 909 15564 910
rect 14538 901 14687 908
rect 14538 900 14579 901
rect 13862 847 13899 848
rect 13958 847 13995 848
rect 14014 847 14050 899
rect 14069 847 14106 848
rect 13762 838 13900 847
rect 13762 818 13871 838
rect 13891 818 13900 838
rect 13762 811 13900 818
rect 13958 838 14106 847
rect 13958 818 13967 838
rect 13987 818 14077 838
rect 14097 818 14106 838
rect 13762 809 13858 811
rect 13958 808 14106 818
rect 14165 838 14202 848
rect 14277 847 14314 848
rect 14258 845 14314 847
rect 14165 818 14173 838
rect 14193 818 14202 838
rect 14014 807 14050 808
rect 13862 748 13899 749
rect 14165 748 14202 818
rect 14227 838 14314 845
rect 14227 835 14285 838
rect 14227 815 14232 835
rect 14253 818 14285 835
rect 14305 818 14314 838
rect 14253 815 14314 818
rect 14227 808 14314 815
rect 14373 838 14410 848
rect 14373 818 14381 838
rect 14401 818 14410 838
rect 14227 807 14258 808
rect 13861 747 14202 748
rect 13786 742 14202 747
rect 13786 722 13789 742
rect 13809 722 14202 742
rect 14373 739 14410 818
rect 14440 847 14471 900
rect 14821 898 14858 899
rect 14820 889 14859 898
rect 14820 871 14830 889
rect 14848 871 14859 889
rect 15200 887 15237 891
rect 14732 854 14779 855
rect 14820 854 14859 871
rect 14732 850 14859 854
rect 14490 847 14527 848
rect 14440 838 14527 847
rect 14440 818 14498 838
rect 14518 818 14527 838
rect 14440 808 14527 818
rect 14586 838 14623 848
rect 14586 818 14594 838
rect 14614 818 14623 838
rect 14440 807 14471 808
rect 14435 739 14545 752
rect 14586 739 14623 818
rect 14732 821 14742 850
rect 14771 821 14859 850
rect 14732 815 14859 821
rect 14732 811 14779 815
rect 14817 801 14859 815
rect 14817 783 14828 801
rect 14846 783 14859 801
rect 14817 778 14859 783
rect 14818 775 14859 778
rect 15197 882 15237 887
rect 15197 864 15209 882
rect 15227 864 15237 882
rect 14818 774 14855 775
rect 14373 737 14623 739
rect 14373 734 14474 737
rect 14373 715 14438 734
rect 14435 707 14438 715
rect 14467 707 14474 734
rect 14502 710 14512 737
rect 14541 715 14623 737
rect 14541 710 14545 715
rect 14502 707 14545 710
rect 14435 693 14545 707
rect 14811 711 14858 712
rect 14811 702 14859 711
rect 11067 689 11235 691
rect 10791 686 11235 689
rect 10452 662 10563 668
rect 10452 654 10493 662
rect 10141 599 10180 643
rect 10452 634 10460 654
rect 10479 634 10493 654
rect 10452 632 10493 634
rect 10521 656 10563 662
rect 10789 663 11235 686
rect 14811 684 14830 702
rect 14848 684 14859 702
rect 14811 682 14859 684
rect 14820 663 14859 682
rect 15197 684 15237 864
rect 15583 857 15614 910
rect 15644 939 15681 1018
rect 15852 1015 16245 1035
rect 16265 1015 16268 1035
rect 16366 1019 16615 1041
rect 16784 1040 16825 1045
rect 17203 1042 17230 1220
rect 17881 1132 17908 1310
rect 18286 1307 18327 1312
rect 18496 1311 18745 1333
rect 18843 1317 18846 1337
rect 18866 1317 19259 1337
rect 19430 1334 19467 1413
rect 19497 1442 19528 1495
rect 19874 1488 19914 1668
rect 19874 1470 19884 1488
rect 19902 1470 19914 1488
rect 19874 1465 19914 1470
rect 19874 1461 19911 1465
rect 19547 1442 19584 1443
rect 19497 1433 19584 1442
rect 19497 1413 19555 1433
rect 19575 1413 19584 1433
rect 19497 1403 19584 1413
rect 19643 1433 19680 1443
rect 19643 1413 19651 1433
rect 19671 1413 19680 1433
rect 19497 1402 19528 1403
rect 19492 1334 19602 1347
rect 19643 1334 19680 1413
rect 19877 1398 19914 1399
rect 19873 1389 19914 1398
rect 19873 1371 19886 1389
rect 19904 1371 19914 1389
rect 19873 1362 19914 1371
rect 19873 1342 19913 1362
rect 19430 1332 19680 1334
rect 19430 1329 19531 1332
rect 17948 1272 18012 1284
rect 18288 1280 18325 1307
rect 18496 1280 18533 1311
rect 18709 1309 18745 1311
rect 19430 1310 19495 1329
rect 18709 1280 18746 1309
rect 19492 1302 19495 1310
rect 19524 1302 19531 1329
rect 19559 1305 19569 1332
rect 19598 1310 19680 1332
rect 19788 1332 19913 1342
rect 19788 1313 19796 1332
rect 19821 1313 19913 1332
rect 19598 1305 19602 1310
rect 19788 1306 19913 1313
rect 19559 1302 19602 1305
rect 19492 1288 19602 1302
rect 17948 1271 17983 1272
rect 17925 1266 17983 1271
rect 17925 1246 17928 1266
rect 17948 1252 17983 1266
rect 18003 1252 18012 1272
rect 17948 1244 18012 1252
rect 17974 1243 18012 1244
rect 17975 1242 18012 1243
rect 18078 1276 18114 1277
rect 18186 1276 18222 1277
rect 18078 1268 18222 1276
rect 18078 1248 18086 1268
rect 18106 1265 18194 1268
rect 18106 1248 18138 1265
rect 18158 1248 18194 1265
rect 18214 1248 18222 1268
rect 18078 1242 18222 1248
rect 18288 1272 18326 1280
rect 18394 1276 18430 1277
rect 18288 1252 18297 1272
rect 18317 1252 18326 1272
rect 18288 1243 18326 1252
rect 18345 1269 18430 1276
rect 18345 1249 18352 1269
rect 18373 1268 18430 1269
rect 18373 1249 18402 1268
rect 18345 1248 18402 1249
rect 18422 1248 18430 1268
rect 18288 1242 18325 1243
rect 18345 1242 18430 1248
rect 18496 1272 18534 1280
rect 18607 1276 18643 1277
rect 18496 1252 18505 1272
rect 18525 1252 18534 1272
rect 18496 1243 18534 1252
rect 18558 1268 18643 1276
rect 18558 1248 18615 1268
rect 18635 1248 18643 1268
rect 18496 1242 18533 1243
rect 18558 1242 18643 1248
rect 18709 1272 18747 1280
rect 18709 1252 18718 1272
rect 18738 1252 18747 1272
rect 18709 1243 18747 1252
rect 19873 1258 19913 1306
rect 18709 1242 18746 1243
rect 18132 1221 18168 1242
rect 18558 1221 18589 1242
rect 19873 1240 19884 1258
rect 19902 1240 19913 1258
rect 19873 1232 19913 1240
rect 19874 1231 19911 1232
rect 17965 1217 18065 1221
rect 17965 1213 18027 1217
rect 17965 1187 17972 1213
rect 17998 1191 18027 1213
rect 18053 1191 18065 1217
rect 17998 1187 18065 1191
rect 17965 1184 18065 1187
rect 18133 1184 18168 1221
rect 18230 1218 18589 1221
rect 18230 1213 18452 1218
rect 18230 1189 18243 1213
rect 18267 1194 18452 1213
rect 18476 1194 18589 1218
rect 18267 1189 18589 1194
rect 18230 1185 18589 1189
rect 18656 1213 18805 1221
rect 18656 1193 18667 1213
rect 18687 1193 18805 1213
rect 18656 1186 18805 1193
rect 19245 1190 19759 1191
rect 18656 1185 18697 1186
rect 17980 1132 18017 1133
rect 18076 1132 18113 1133
rect 18132 1132 18168 1184
rect 18187 1132 18224 1133
rect 17880 1123 18018 1132
rect 17880 1103 17989 1123
rect 18009 1103 18018 1123
rect 17880 1096 18018 1103
rect 18076 1123 18224 1132
rect 18076 1103 18085 1123
rect 18105 1103 18195 1123
rect 18215 1103 18224 1123
rect 17880 1094 17976 1096
rect 18076 1093 18224 1103
rect 18283 1123 18320 1133
rect 18395 1132 18432 1133
rect 18376 1130 18432 1132
rect 18283 1103 18291 1123
rect 18311 1103 18320 1123
rect 18132 1092 18168 1093
rect 17062 1040 17230 1042
rect 16784 1034 17230 1040
rect 15852 1010 16268 1015
rect 16447 1013 16558 1019
rect 15852 1009 16193 1010
rect 15796 949 15827 950
rect 15644 919 15653 939
rect 15673 919 15681 939
rect 15644 909 15681 919
rect 15740 942 15827 949
rect 15740 939 15801 942
rect 15740 919 15749 939
rect 15769 922 15801 939
rect 15822 922 15827 942
rect 15769 919 15827 922
rect 15740 912 15827 919
rect 15852 939 15889 1009
rect 16155 1008 16192 1009
rect 16447 1005 16488 1013
rect 16447 985 16455 1005
rect 16474 985 16488 1005
rect 16447 983 16488 985
rect 16516 1005 16558 1013
rect 16516 985 16532 1005
rect 16551 985 16558 1005
rect 16784 1012 16790 1034
rect 16816 1014 17230 1034
rect 17980 1033 18017 1034
rect 18283 1033 18320 1103
rect 18345 1123 18432 1130
rect 18345 1120 18403 1123
rect 18345 1100 18350 1120
rect 18371 1103 18403 1120
rect 18423 1103 18432 1123
rect 18371 1100 18432 1103
rect 18345 1093 18432 1100
rect 18491 1123 18528 1133
rect 18491 1103 18499 1123
rect 18519 1103 18528 1123
rect 18345 1092 18376 1093
rect 17979 1032 18320 1033
rect 16816 1012 16825 1014
rect 17062 1013 17230 1014
rect 17904 1027 18320 1032
rect 16784 1003 16825 1012
rect 17904 1007 17907 1027
rect 17927 1007 18320 1027
rect 18491 1024 18528 1103
rect 18558 1132 18589 1185
rect 19226 1174 19759 1190
rect 19226 1163 19758 1174
rect 19877 1165 19914 1169
rect 18608 1132 18645 1133
rect 18558 1123 18645 1132
rect 18558 1103 18616 1123
rect 18636 1103 18645 1123
rect 18558 1093 18645 1103
rect 18704 1123 18741 1133
rect 18704 1103 18712 1123
rect 18732 1103 18741 1123
rect 18558 1092 18589 1093
rect 18553 1024 18663 1037
rect 18704 1024 18741 1103
rect 18491 1022 18741 1024
rect 18491 1019 18592 1022
rect 18491 1000 18556 1019
rect 16516 983 16558 985
rect 16447 968 16558 983
rect 18553 992 18556 1000
rect 18585 992 18592 1019
rect 18620 995 18630 1022
rect 18659 1000 18741 1022
rect 18819 1094 18987 1095
rect 19226 1094 19264 1163
rect 18819 1074 19264 1094
rect 19491 1125 19602 1140
rect 19491 1123 19533 1125
rect 19491 1103 19498 1123
rect 19517 1103 19533 1123
rect 19491 1095 19533 1103
rect 19561 1123 19602 1125
rect 19561 1103 19575 1123
rect 19594 1103 19602 1123
rect 19561 1095 19602 1103
rect 19491 1089 19602 1095
rect 19724 1100 19758 1163
rect 19876 1159 19914 1165
rect 19876 1141 19886 1159
rect 19904 1141 19914 1159
rect 19876 1132 19914 1141
rect 19876 1100 19910 1132
rect 18819 1068 19263 1074
rect 18819 1066 18987 1068
rect 18659 995 18663 1000
rect 18620 992 18663 995
rect 18553 978 18663 992
rect 16004 949 16040 950
rect 15852 919 15861 939
rect 15881 919 15889 939
rect 15740 910 15796 912
rect 15740 909 15777 910
rect 15852 909 15889 919
rect 15948 939 16096 949
rect 16196 946 16292 948
rect 15948 919 15957 939
rect 15977 919 16067 939
rect 16087 919 16096 939
rect 15948 910 16096 919
rect 16154 939 16292 946
rect 16154 919 16163 939
rect 16183 919 16292 939
rect 16154 910 16292 919
rect 15948 909 15985 910
rect 16004 858 16040 910
rect 16059 909 16096 910
rect 16155 909 16192 910
rect 15475 856 15516 857
rect 15367 849 15516 856
rect 15367 829 15485 849
rect 15505 829 15516 849
rect 15367 821 15516 829
rect 15583 853 15942 857
rect 15583 848 15905 853
rect 15583 824 15696 848
rect 15720 829 15905 848
rect 15929 829 15942 853
rect 15720 824 15942 829
rect 15583 821 15942 824
rect 16004 821 16039 858
rect 16107 855 16207 858
rect 16107 851 16174 855
rect 16107 825 16119 851
rect 16145 829 16174 851
rect 16200 829 16207 855
rect 16145 825 16207 829
rect 16107 821 16207 825
rect 15583 800 15614 821
rect 16004 800 16040 821
rect 15426 799 15463 800
rect 15425 790 15463 799
rect 15425 770 15434 790
rect 15454 770 15463 790
rect 15425 762 15463 770
rect 15529 794 15614 800
rect 15639 799 15676 800
rect 15529 774 15537 794
rect 15557 774 15614 794
rect 15529 766 15614 774
rect 15638 790 15676 799
rect 15638 770 15647 790
rect 15667 770 15676 790
rect 15529 765 15565 766
rect 15638 762 15676 770
rect 15742 794 15827 800
rect 15847 799 15884 800
rect 15742 774 15750 794
rect 15770 793 15827 794
rect 15770 774 15799 793
rect 15742 773 15799 774
rect 15820 773 15827 793
rect 15742 766 15827 773
rect 15846 790 15884 799
rect 15846 770 15855 790
rect 15875 770 15884 790
rect 15742 765 15778 766
rect 15846 762 15884 770
rect 15950 794 16094 800
rect 15950 774 15958 794
rect 15978 791 16066 794
rect 15978 774 16009 791
rect 15950 771 16009 774
rect 16032 774 16066 791
rect 16086 774 16094 794
rect 16032 771 16094 774
rect 15950 766 16094 771
rect 15950 765 15986 766
rect 16058 765 16094 766
rect 16160 799 16197 800
rect 16160 798 16198 799
rect 16160 790 16224 798
rect 16160 770 16169 790
rect 16189 776 16224 790
rect 16244 776 16247 796
rect 16189 771 16247 776
rect 16189 770 16224 771
rect 15426 733 15463 762
rect 15427 731 15463 733
rect 15639 731 15676 762
rect 15427 709 15676 731
rect 15847 730 15884 762
rect 16160 758 16224 770
rect 16264 732 16291 910
rect 18819 888 18846 1066
rect 18886 1028 18950 1040
rect 19226 1036 19263 1068
rect 19434 1067 19683 1089
rect 19724 1068 19910 1100
rect 19738 1067 19910 1068
rect 19434 1036 19471 1067
rect 19647 1065 19683 1067
rect 19647 1036 19684 1065
rect 19876 1039 19910 1067
rect 18886 1027 18921 1028
rect 18863 1022 18921 1027
rect 18863 1002 18866 1022
rect 18886 1008 18921 1022
rect 18941 1008 18950 1028
rect 18886 1000 18950 1008
rect 18912 999 18950 1000
rect 18913 998 18950 999
rect 19016 1032 19052 1033
rect 19124 1032 19160 1033
rect 19016 1025 19160 1032
rect 19016 1024 19076 1025
rect 19016 1004 19024 1024
rect 19044 1005 19076 1024
rect 19101 1024 19160 1025
rect 19101 1005 19132 1024
rect 19044 1004 19132 1005
rect 19152 1004 19160 1024
rect 19016 998 19160 1004
rect 19226 1028 19264 1036
rect 19332 1032 19368 1033
rect 19226 1008 19235 1028
rect 19255 1008 19264 1028
rect 19226 999 19264 1008
rect 19283 1025 19368 1032
rect 19283 1005 19290 1025
rect 19311 1024 19368 1025
rect 19311 1005 19340 1024
rect 19283 1004 19340 1005
rect 19360 1004 19368 1024
rect 19226 998 19263 999
rect 19283 998 19368 1004
rect 19434 1028 19472 1036
rect 19545 1032 19581 1033
rect 19434 1008 19443 1028
rect 19463 1008 19472 1028
rect 19434 999 19472 1008
rect 19496 1024 19581 1032
rect 19496 1004 19553 1024
rect 19573 1004 19581 1024
rect 19434 998 19471 999
rect 19496 998 19581 1004
rect 19647 1028 19685 1036
rect 19647 1008 19656 1028
rect 19676 1008 19685 1028
rect 19647 999 19685 1008
rect 19874 1029 19911 1039
rect 19874 1011 19884 1029
rect 19902 1011 19911 1029
rect 19874 1002 19911 1011
rect 19876 1001 19910 1002
rect 19647 998 19684 999
rect 19070 977 19106 998
rect 19496 977 19527 998
rect 18903 973 19003 977
rect 18903 969 18965 973
rect 18903 943 18910 969
rect 18936 947 18965 969
rect 18991 947 19003 973
rect 18936 943 19003 947
rect 18903 940 19003 943
rect 19071 940 19106 977
rect 19168 974 19527 977
rect 19168 969 19390 974
rect 19168 945 19181 969
rect 19205 950 19390 969
rect 19414 950 19527 974
rect 19205 945 19527 950
rect 19168 941 19527 945
rect 19594 969 19743 977
rect 19594 949 19605 969
rect 19625 949 19743 969
rect 19594 942 19743 949
rect 19594 941 19635 942
rect 18918 888 18955 889
rect 19014 888 19051 889
rect 19070 888 19106 940
rect 19125 888 19162 889
rect 18818 879 18956 888
rect 18818 859 18927 879
rect 18947 859 18956 879
rect 18818 852 18956 859
rect 19014 879 19162 888
rect 19014 859 19023 879
rect 19043 859 19133 879
rect 19153 859 19162 879
rect 18818 850 18914 852
rect 19014 849 19162 859
rect 19221 879 19258 889
rect 19333 888 19370 889
rect 19314 886 19370 888
rect 19221 859 19229 879
rect 19249 859 19258 879
rect 19070 848 19106 849
rect 18918 789 18955 790
rect 19221 789 19258 859
rect 19283 879 19370 886
rect 19283 876 19341 879
rect 19283 856 19288 876
rect 19309 859 19341 876
rect 19361 859 19370 879
rect 19309 856 19370 859
rect 19283 849 19370 856
rect 19429 879 19466 889
rect 19429 859 19437 879
rect 19457 859 19466 879
rect 19283 848 19314 849
rect 18917 788 19258 789
rect 18842 783 19258 788
rect 18842 763 18845 783
rect 18865 763 19258 783
rect 19429 780 19466 859
rect 19496 888 19527 941
rect 19877 939 19914 940
rect 19876 930 19915 939
rect 19876 912 19886 930
rect 19904 912 19915 930
rect 19788 895 19835 896
rect 19876 895 19915 912
rect 19788 891 19915 895
rect 19546 888 19583 889
rect 19496 879 19583 888
rect 19496 859 19554 879
rect 19574 859 19583 879
rect 19496 849 19583 859
rect 19642 879 19679 889
rect 19642 859 19650 879
rect 19670 859 19679 879
rect 19496 848 19527 849
rect 19491 780 19601 793
rect 19642 780 19679 859
rect 19788 862 19798 891
rect 19827 862 19915 891
rect 19788 856 19915 862
rect 19788 852 19835 856
rect 19873 842 19915 856
rect 19873 824 19884 842
rect 19902 824 19915 842
rect 19873 819 19915 824
rect 19874 816 19915 819
rect 19874 815 19911 816
rect 19429 778 19679 780
rect 19429 775 19530 778
rect 19429 756 19494 775
rect 19491 748 19494 756
rect 19523 748 19530 775
rect 19558 751 19568 778
rect 19597 756 19679 778
rect 19597 751 19601 756
rect 19558 748 19601 751
rect 19491 734 19601 748
rect 19867 752 19914 753
rect 19867 743 19915 752
rect 16123 730 16291 732
rect 15847 727 16291 730
rect 15508 703 15619 709
rect 15508 695 15549 703
rect 10521 654 10562 656
rect 10521 634 10537 654
rect 10556 634 10562 654
rect 10521 632 10562 634
rect 10452 617 10562 632
rect 4787 550 4792 571
rect 4821 550 4831 571
rect 5774 568 5853 578
rect 10141 575 10181 599
rect 10789 589 10827 663
rect 11067 662 11235 663
rect 10749 575 10828 589
rect 10141 574 10431 575
rect 10597 574 10828 575
rect 10141 572 10828 574
rect 4787 537 4831 550
rect 10141 551 10788 572
rect 10817 551 10828 572
rect 10141 542 10828 551
rect 14818 576 14862 663
rect 15197 640 15236 684
rect 15508 675 15516 695
rect 15535 675 15549 695
rect 15508 673 15549 675
rect 15577 697 15619 703
rect 15845 704 16291 727
rect 19867 725 19886 743
rect 19904 725 19915 743
rect 19867 723 19915 725
rect 19876 704 19915 723
rect 15577 695 15618 697
rect 15577 675 15593 695
rect 15612 675 15618 695
rect 15577 673 15618 675
rect 15508 658 15618 673
rect 15197 616 15237 640
rect 15845 630 15883 704
rect 16123 703 16291 704
rect 15805 616 15884 630
rect 15197 615 15487 616
rect 15653 615 15884 616
rect 15197 613 15884 615
rect 15197 592 15844 613
rect 15873 592 15884 613
rect 15197 583 15884 592
rect 19874 617 19918 704
rect 19874 596 19879 617
rect 19908 596 19918 617
rect 19874 583 19918 596
rect 14818 555 14823 576
rect 14852 555 14862 576
rect 15805 573 15884 583
rect 14818 542 14862 555
rect 718 527 797 537
rect 10749 532 10828 542
rect 6725 486 6835 500
rect 6725 483 6768 486
rect 6725 478 6729 483
rect 1669 445 1779 459
rect 1669 442 1712 445
rect 1669 437 1673 442
rect 1591 415 1673 437
rect 1702 415 1712 442
rect 1740 418 1747 445
rect 1776 437 1779 445
rect 6647 456 6729 478
rect 6758 456 6768 483
rect 6796 459 6803 486
rect 6832 478 6835 486
rect 16756 491 16866 505
rect 16756 488 16799 491
rect 16756 483 16760 488
rect 6832 459 6897 478
rect 6796 456 6897 459
rect 6647 454 6897 456
rect 1776 418 1841 437
rect 1740 415 1841 418
rect 1591 413 1841 415
rect 1591 334 1628 413
rect 1669 400 1779 413
rect 1743 344 1774 345
rect 1591 314 1600 334
rect 1620 314 1628 334
rect 1591 304 1628 314
rect 1687 334 1774 344
rect 1687 314 1696 334
rect 1716 314 1774 334
rect 1687 305 1774 314
rect 1687 304 1724 305
rect 1743 252 1774 305
rect 1804 334 1841 413
rect 2012 410 2405 430
rect 2425 410 2428 430
rect 4619 425 4729 439
rect 4619 422 4662 425
rect 4619 417 4623 422
rect 2012 405 2428 410
rect 2012 404 2353 405
rect 1956 344 1987 345
rect 1804 314 1813 334
rect 1833 314 1841 334
rect 1804 304 1841 314
rect 1900 337 1987 344
rect 1900 334 1961 337
rect 1900 314 1909 334
rect 1929 317 1961 334
rect 1982 317 1987 337
rect 1929 314 1987 317
rect 1900 307 1987 314
rect 2012 334 2049 404
rect 2315 403 2352 404
rect 4541 395 4623 417
rect 4652 395 4662 422
rect 4690 398 4697 425
rect 4726 417 4729 425
rect 4726 398 4791 417
rect 4690 395 4791 398
rect 4541 393 4791 395
rect 2164 344 2200 345
rect 2012 314 2021 334
rect 2041 314 2049 334
rect 1900 305 1956 307
rect 1900 304 1937 305
rect 2012 304 2049 314
rect 2108 334 2256 344
rect 2356 341 2452 343
rect 2108 314 2117 334
rect 2137 314 2227 334
rect 2247 314 2256 334
rect 2108 305 2256 314
rect 2314 334 2452 341
rect 2314 314 2323 334
rect 2343 314 2452 334
rect 2314 305 2452 314
rect 4541 314 4578 393
rect 4619 380 4729 393
rect 4693 324 4724 325
rect 2108 304 2145 305
rect 2164 253 2200 305
rect 2219 304 2256 305
rect 2315 304 2352 305
rect 1635 251 1676 252
rect 1527 244 1676 251
rect 1527 224 1645 244
rect 1665 224 1676 244
rect 1527 216 1676 224
rect 1743 248 2102 252
rect 1743 243 2065 248
rect 1743 219 1856 243
rect 1880 224 2065 243
rect 2089 224 2102 248
rect 1880 219 2102 224
rect 1743 216 2102 219
rect 2164 216 2199 253
rect 2267 250 2367 253
rect 2267 246 2334 250
rect 2267 220 2279 246
rect 2305 224 2334 246
rect 2360 224 2367 250
rect 2305 220 2367 224
rect 2267 216 2367 220
rect 1743 195 1774 216
rect 2164 195 2200 216
rect 1586 194 1623 195
rect 1585 185 1623 194
rect 1585 165 1594 185
rect 1614 165 1623 185
rect 1585 157 1623 165
rect 1689 189 1774 195
rect 1799 194 1836 195
rect 1689 169 1697 189
rect 1717 169 1774 189
rect 1689 161 1774 169
rect 1798 185 1836 194
rect 1798 165 1807 185
rect 1827 165 1836 185
rect 1689 160 1725 161
rect 1798 157 1836 165
rect 1902 189 1987 195
rect 2007 194 2044 195
rect 1902 169 1910 189
rect 1930 188 1987 189
rect 1930 169 1959 188
rect 1902 168 1959 169
rect 1980 168 1987 188
rect 1902 161 1987 168
rect 2006 185 2044 194
rect 2006 165 2015 185
rect 2035 165 2044 185
rect 1902 160 1938 161
rect 2006 157 2044 165
rect 2110 189 2254 195
rect 2110 169 2118 189
rect 2138 187 2226 189
rect 2138 169 2165 187
rect 2110 167 2165 169
rect 2199 169 2226 187
rect 2246 169 2254 189
rect 2199 167 2254 169
rect 2110 161 2254 167
rect 2110 160 2146 161
rect 2218 160 2254 161
rect 2320 194 2357 195
rect 2320 193 2358 194
rect 2320 185 2384 193
rect 2320 165 2329 185
rect 2349 171 2384 185
rect 2404 171 2407 191
rect 2349 166 2407 171
rect 2349 165 2384 166
rect 1586 128 1623 157
rect 1587 126 1623 128
rect 1799 126 1836 157
rect 1587 104 1836 126
rect 2007 125 2044 157
rect 2320 153 2384 165
rect 2424 136 2451 305
rect 4541 294 4550 314
rect 4570 294 4578 314
rect 4541 284 4578 294
rect 4637 314 4724 324
rect 4637 294 4646 314
rect 4666 294 4724 314
rect 4637 285 4724 294
rect 4637 284 4674 285
rect 4693 232 4724 285
rect 4754 314 4791 393
rect 4962 390 5355 410
rect 5375 390 5378 410
rect 4962 385 5378 390
rect 4962 384 5303 385
rect 4906 324 4937 325
rect 4754 294 4763 314
rect 4783 294 4791 314
rect 4754 284 4791 294
rect 4850 317 4937 324
rect 4850 314 4911 317
rect 4850 294 4859 314
rect 4879 297 4911 314
rect 4932 297 4937 317
rect 4879 294 4937 297
rect 4850 287 4937 294
rect 4962 314 4999 384
rect 5265 383 5302 384
rect 6647 375 6684 454
rect 6725 441 6835 454
rect 6799 385 6830 386
rect 6647 355 6656 375
rect 6676 355 6684 375
rect 6647 345 6684 355
rect 6743 375 6830 385
rect 6743 355 6752 375
rect 6772 355 6830 375
rect 6743 346 6830 355
rect 6743 345 6780 346
rect 5114 324 5150 325
rect 4962 294 4971 314
rect 4991 294 4999 314
rect 4850 285 4906 287
rect 4850 284 4887 285
rect 4962 284 4999 294
rect 5058 314 5206 324
rect 5306 321 5402 323
rect 5058 294 5067 314
rect 5087 294 5177 314
rect 5197 294 5206 314
rect 5058 285 5206 294
rect 5264 314 5402 321
rect 5264 294 5273 314
rect 5293 294 5402 314
rect 5264 285 5402 294
rect 6799 293 6830 346
rect 6860 375 6897 454
rect 7068 451 7461 471
rect 7481 451 7484 471
rect 7068 446 7484 451
rect 11700 450 11810 464
rect 11700 447 11743 450
rect 7068 445 7409 446
rect 7012 385 7043 386
rect 6860 355 6869 375
rect 6889 355 6897 375
rect 6860 345 6897 355
rect 6956 378 7043 385
rect 6956 375 7017 378
rect 6956 355 6965 375
rect 6985 358 7017 375
rect 7038 358 7043 378
rect 6985 355 7043 358
rect 6956 348 7043 355
rect 7068 375 7105 445
rect 7371 444 7408 445
rect 11700 442 11704 447
rect 11622 420 11704 442
rect 11733 420 11743 447
rect 11771 423 11778 450
rect 11807 442 11810 450
rect 16678 461 16760 483
rect 16789 461 16799 488
rect 16827 464 16834 491
rect 16863 483 16866 491
rect 16863 464 16928 483
rect 16827 461 16928 464
rect 16678 459 16928 461
rect 11807 423 11872 442
rect 11771 420 11872 423
rect 11622 418 11872 420
rect 7220 385 7256 386
rect 7068 355 7077 375
rect 7097 355 7105 375
rect 6956 346 7012 348
rect 6956 345 6993 346
rect 7068 345 7105 355
rect 7164 375 7312 385
rect 7412 382 7508 384
rect 7164 355 7173 375
rect 7193 355 7283 375
rect 7303 355 7312 375
rect 7164 346 7312 355
rect 7370 375 7508 382
rect 7370 355 7379 375
rect 7399 355 7508 375
rect 7370 346 7508 355
rect 7164 345 7201 346
rect 7220 294 7256 346
rect 7275 345 7312 346
rect 7371 345 7408 346
rect 6691 292 6732 293
rect 6583 285 6732 292
rect 5058 284 5095 285
rect 5114 264 5150 285
rect 5169 284 5206 285
rect 5265 284 5302 285
rect 5112 234 5150 264
rect 5114 233 5150 234
rect 4585 231 4626 232
rect 4477 224 4626 231
rect 4477 204 4595 224
rect 4615 204 4626 224
rect 4477 196 4626 204
rect 4693 228 5052 232
rect 4693 223 5015 228
rect 4693 199 4806 223
rect 4830 204 5015 223
rect 5039 204 5052 228
rect 4830 199 5052 204
rect 4693 196 5052 199
rect 5114 196 5149 233
rect 5217 230 5317 233
rect 5217 226 5284 230
rect 5217 200 5229 226
rect 5255 204 5284 226
rect 5310 204 5317 230
rect 5255 200 5317 204
rect 5217 196 5317 200
rect 4693 175 4724 196
rect 5114 175 5150 196
rect 4536 174 4573 175
rect 4535 165 4573 174
rect 4535 145 4544 165
rect 4564 145 4573 165
rect 4535 137 4573 145
rect 4639 169 4724 175
rect 4749 174 4786 175
rect 4639 149 4647 169
rect 4667 149 4724 169
rect 4639 141 4724 149
rect 4748 165 4786 174
rect 4748 145 4757 165
rect 4777 145 4786 165
rect 4639 140 4675 141
rect 4748 137 4786 145
rect 4852 169 4937 175
rect 4957 174 4994 175
rect 4852 149 4860 169
rect 4880 168 4937 169
rect 4880 149 4909 168
rect 4852 148 4909 149
rect 4930 148 4937 168
rect 4852 141 4937 148
rect 4956 165 4994 174
rect 4956 145 4965 165
rect 4985 145 4994 165
rect 4852 140 4888 141
rect 4956 137 4994 145
rect 5060 169 5204 175
rect 5060 149 5068 169
rect 5088 167 5176 169
rect 5088 149 5109 167
rect 5060 147 5109 149
rect 5150 149 5176 167
rect 5196 149 5204 169
rect 5150 147 5204 149
rect 5060 141 5204 147
rect 5060 140 5096 141
rect 5168 140 5204 141
rect 5270 174 5307 175
rect 5270 173 5308 174
rect 5270 165 5334 173
rect 5270 145 5279 165
rect 5299 151 5334 165
rect 5354 151 5357 171
rect 5299 146 5357 151
rect 5299 145 5334 146
rect 2397 130 2525 136
rect 2397 127 2486 130
rect 2283 125 2486 127
rect 2007 109 2486 125
rect 2513 109 2525 130
rect 1668 98 1779 104
rect 2007 99 2525 109
rect 4536 108 4573 137
rect 2283 98 2525 99
rect 1668 90 1709 98
rect 1668 70 1676 90
rect 1695 70 1709 90
rect 1668 68 1709 70
rect 1737 90 1779 98
rect 2397 96 2525 98
rect 4537 106 4573 108
rect 4749 106 4786 137
rect 1737 70 1753 90
rect 1772 70 1779 90
rect 4537 84 4786 106
rect 4957 105 4994 137
rect 5270 133 5334 145
rect 5374 125 5401 285
rect 6583 265 6701 285
rect 6721 265 6732 285
rect 6583 257 6732 265
rect 6799 289 7158 293
rect 6799 284 7121 289
rect 6799 260 6912 284
rect 6936 265 7121 284
rect 7145 265 7158 289
rect 6936 260 7158 265
rect 6799 257 7158 260
rect 7220 257 7255 294
rect 7323 291 7423 294
rect 7323 287 7390 291
rect 7323 261 7335 287
rect 7361 265 7390 287
rect 7416 265 7423 291
rect 7361 261 7423 265
rect 7323 257 7423 261
rect 6799 236 6830 257
rect 7220 236 7256 257
rect 6642 235 6679 236
rect 6641 226 6679 235
rect 6641 206 6650 226
rect 6670 206 6679 226
rect 6641 198 6679 206
rect 6745 230 6830 236
rect 6855 235 6892 236
rect 6745 210 6753 230
rect 6773 210 6830 230
rect 6745 202 6830 210
rect 6854 226 6892 235
rect 6854 206 6863 226
rect 6883 206 6892 226
rect 6745 201 6781 202
rect 6854 198 6892 206
rect 6958 230 7043 236
rect 7063 235 7100 236
rect 6958 210 6966 230
rect 6986 229 7043 230
rect 6986 210 7015 229
rect 6958 209 7015 210
rect 7036 209 7043 229
rect 6958 202 7043 209
rect 7062 226 7100 235
rect 7062 206 7071 226
rect 7091 206 7100 226
rect 6958 201 6994 202
rect 7062 198 7100 206
rect 7166 230 7310 236
rect 7166 210 7174 230
rect 7194 228 7282 230
rect 7194 210 7221 228
rect 7166 208 7221 210
rect 7255 210 7282 228
rect 7302 210 7310 230
rect 7255 208 7310 210
rect 7166 202 7310 208
rect 7166 201 7202 202
rect 7274 201 7310 202
rect 7376 235 7413 236
rect 7376 234 7414 235
rect 7376 226 7440 234
rect 7376 206 7385 226
rect 7405 212 7440 226
rect 7460 212 7463 232
rect 7405 207 7463 212
rect 7405 206 7440 207
rect 6642 169 6679 198
rect 6643 167 6679 169
rect 6855 167 6892 198
rect 6643 145 6892 167
rect 7063 166 7100 198
rect 7376 194 7440 206
rect 7480 177 7507 346
rect 11622 339 11659 418
rect 11700 405 11810 418
rect 11774 349 11805 350
rect 9553 309 9663 323
rect 11622 319 11631 339
rect 11651 319 11659 339
rect 11622 309 11659 319
rect 11718 339 11805 349
rect 11718 319 11727 339
rect 11747 319 11805 339
rect 11718 310 11805 319
rect 11718 309 11755 310
rect 9553 306 9596 309
rect 9553 301 9557 306
rect 9475 279 9557 301
rect 9586 279 9596 306
rect 9624 282 9631 309
rect 9660 301 9663 309
rect 9660 282 9725 301
rect 9624 279 9725 282
rect 9475 277 9725 279
rect 9475 198 9512 277
rect 9553 264 9663 277
rect 9627 208 9658 209
rect 9475 178 9484 198
rect 9504 178 9512 198
rect 7453 171 7581 177
rect 7453 168 7542 171
rect 7339 166 7542 168
rect 7063 150 7542 166
rect 7569 150 7581 171
rect 9475 168 9512 178
rect 9571 198 9658 208
rect 9571 178 9580 198
rect 9600 178 9658 198
rect 9571 169 9658 178
rect 9571 168 9608 169
rect 6724 139 6835 145
rect 7063 140 7581 150
rect 7339 139 7581 140
rect 6724 131 6765 139
rect 5370 111 5493 125
rect 5370 107 5422 111
rect 5233 105 5422 107
rect 4957 85 5422 105
rect 5481 85 5493 111
rect 6724 111 6732 131
rect 6751 111 6765 131
rect 6724 109 6765 111
rect 6793 131 6835 139
rect 7453 137 7581 139
rect 6793 111 6809 131
rect 6828 111 6835 131
rect 9627 116 9658 169
rect 9688 198 9725 277
rect 9896 274 10289 294
rect 10309 274 10312 294
rect 9896 269 10312 274
rect 9896 268 10237 269
rect 9840 208 9871 209
rect 9688 178 9697 198
rect 9717 178 9725 198
rect 9688 168 9725 178
rect 9784 201 9871 208
rect 9784 198 9845 201
rect 9784 178 9793 198
rect 9813 181 9845 198
rect 9866 181 9871 201
rect 9813 178 9871 181
rect 9784 171 9871 178
rect 9896 198 9933 268
rect 10199 267 10236 268
rect 11774 257 11805 310
rect 11835 339 11872 418
rect 12043 415 12436 435
rect 12456 415 12459 435
rect 14650 430 14760 444
rect 14650 427 14693 430
rect 14650 422 14654 427
rect 12043 410 12459 415
rect 12043 409 12384 410
rect 11987 349 12018 350
rect 11835 319 11844 339
rect 11864 319 11872 339
rect 11835 309 11872 319
rect 11931 342 12018 349
rect 11931 339 11992 342
rect 11931 319 11940 339
rect 11960 322 11992 339
rect 12013 322 12018 342
rect 11960 319 12018 322
rect 11931 312 12018 319
rect 12043 339 12080 409
rect 12346 408 12383 409
rect 14572 400 14654 422
rect 14683 400 14693 427
rect 14721 403 14728 430
rect 14757 422 14760 430
rect 14757 403 14822 422
rect 14721 400 14822 403
rect 14572 398 14822 400
rect 12195 349 12231 350
rect 12043 319 12052 339
rect 12072 319 12080 339
rect 11931 310 11987 312
rect 11931 309 11968 310
rect 12043 309 12080 319
rect 12139 339 12287 349
rect 12387 346 12483 348
rect 12139 319 12148 339
rect 12168 319 12258 339
rect 12278 319 12287 339
rect 12139 310 12287 319
rect 12345 339 12483 346
rect 12345 319 12354 339
rect 12374 319 12483 339
rect 12345 310 12483 319
rect 14572 319 14609 398
rect 14650 385 14760 398
rect 14724 329 14755 330
rect 12139 309 12176 310
rect 12195 258 12231 310
rect 12250 309 12287 310
rect 12346 309 12383 310
rect 11666 256 11707 257
rect 11558 249 11707 256
rect 11558 229 11676 249
rect 11696 229 11707 249
rect 11558 221 11707 229
rect 11774 253 12133 257
rect 11774 248 12096 253
rect 11774 224 11887 248
rect 11911 229 12096 248
rect 12120 229 12133 253
rect 11911 224 12133 229
rect 11774 221 12133 224
rect 12195 221 12230 258
rect 12298 255 12398 258
rect 12298 251 12365 255
rect 12298 225 12310 251
rect 12336 229 12365 251
rect 12391 229 12398 255
rect 12336 225 12398 229
rect 12298 221 12398 225
rect 10048 208 10084 209
rect 9896 178 9905 198
rect 9925 178 9933 198
rect 9784 169 9840 171
rect 9784 168 9821 169
rect 9896 168 9933 178
rect 9992 198 10140 208
rect 10240 205 10336 207
rect 9992 178 10001 198
rect 10021 178 10111 198
rect 10131 178 10140 198
rect 9992 169 10140 178
rect 10198 198 10336 205
rect 11774 200 11805 221
rect 12195 200 12231 221
rect 11617 199 11654 200
rect 10198 178 10207 198
rect 10227 178 10336 198
rect 10198 169 10336 178
rect 11616 190 11654 199
rect 11616 170 11625 190
rect 11645 170 11654 190
rect 9992 168 10029 169
rect 10048 117 10084 169
rect 10103 168 10140 169
rect 10199 168 10236 169
rect 9519 115 9560 116
rect 6793 109 6835 111
rect 6724 94 6835 109
rect 9411 108 9560 115
rect 1737 68 1779 70
rect 1668 53 1779 68
rect 4618 78 4729 84
rect 4957 79 5493 85
rect 9411 88 9529 108
rect 9549 88 9560 108
rect 9411 80 9560 88
rect 9627 112 9986 116
rect 9627 107 9949 112
rect 9627 83 9740 107
rect 9764 88 9949 107
rect 9973 88 9986 112
rect 9764 83 9986 88
rect 9627 80 9986 83
rect 10048 80 10083 117
rect 10151 114 10251 117
rect 10151 110 10218 114
rect 10151 84 10163 110
rect 10189 88 10218 110
rect 10244 88 10251 114
rect 10189 84 10251 88
rect 10151 80 10251 84
rect 5233 78 5493 79
rect 4618 70 4659 78
rect 4618 50 4626 70
rect 4645 50 4659 70
rect 4618 48 4659 50
rect 4687 70 4729 78
rect 5361 76 5493 78
rect 5404 74 5493 76
rect 4687 50 4703 70
rect 4722 50 4729 70
rect 9627 59 9658 80
rect 10048 59 10084 80
rect 9470 58 9507 59
rect 4687 48 4729 50
rect 4618 33 4729 48
rect 9469 49 9507 58
rect 9469 29 9478 49
rect 9498 29 9507 49
rect 9469 21 9507 29
rect 9573 53 9658 59
rect 9683 58 9720 59
rect 9573 33 9581 53
rect 9601 33 9658 53
rect 9573 25 9658 33
rect 9682 49 9720 58
rect 9682 29 9691 49
rect 9711 29 9720 49
rect 9573 24 9609 25
rect 9682 21 9720 29
rect 9786 53 9871 59
rect 9891 58 9928 59
rect 9786 33 9794 53
rect 9814 52 9871 53
rect 9814 33 9843 52
rect 9786 32 9843 33
rect 9864 32 9871 52
rect 9786 25 9871 32
rect 9890 49 9928 58
rect 9890 29 9899 49
rect 9919 29 9928 49
rect 9786 24 9822 25
rect 9890 21 9928 29
rect 9994 53 10138 59
rect 9994 33 10002 53
rect 10022 52 10110 53
rect 10022 33 10050 52
rect 9994 28 10050 33
rect 10083 33 10110 52
rect 10130 33 10138 53
rect 10083 28 10138 33
rect 9994 25 10138 28
rect 9994 24 10030 25
rect 10102 24 10138 25
rect 10204 58 10241 59
rect 10204 57 10242 58
rect 10204 49 10268 57
rect 10204 29 10213 49
rect 10233 35 10268 49
rect 10288 35 10291 55
rect 10233 30 10291 35
rect 10233 29 10268 30
rect 9470 -8 9507 21
rect 9471 -10 9507 -8
rect 9683 -10 9720 21
rect 9471 -32 9720 -10
rect 9891 -11 9928 21
rect 10204 17 10268 29
rect 10308 -2 10335 169
rect 11616 162 11654 170
rect 11720 194 11805 200
rect 11830 199 11867 200
rect 11720 174 11728 194
rect 11748 174 11805 194
rect 11720 166 11805 174
rect 11829 190 11867 199
rect 11829 170 11838 190
rect 11858 170 11867 190
rect 11720 165 11756 166
rect 11829 162 11867 170
rect 11933 194 12018 200
rect 12038 199 12075 200
rect 11933 174 11941 194
rect 11961 193 12018 194
rect 11961 174 11990 193
rect 11933 173 11990 174
rect 12011 173 12018 193
rect 11933 166 12018 173
rect 12037 190 12075 199
rect 12037 170 12046 190
rect 12066 170 12075 190
rect 11933 165 11969 166
rect 12037 162 12075 170
rect 12141 194 12285 200
rect 12141 174 12149 194
rect 12169 192 12257 194
rect 12169 174 12196 192
rect 12141 172 12196 174
rect 12230 174 12257 192
rect 12277 174 12285 194
rect 12230 172 12285 174
rect 12141 166 12285 172
rect 12141 165 12177 166
rect 12249 165 12285 166
rect 12351 199 12388 200
rect 12351 198 12389 199
rect 12351 190 12415 198
rect 12351 170 12360 190
rect 12380 176 12415 190
rect 12435 176 12438 196
rect 12380 171 12438 176
rect 12380 170 12415 171
rect 11617 133 11654 162
rect 11618 131 11654 133
rect 11830 131 11867 162
rect 11618 109 11867 131
rect 12038 130 12075 162
rect 12351 158 12415 170
rect 12455 141 12482 310
rect 14572 299 14581 319
rect 14601 299 14609 319
rect 14572 289 14609 299
rect 14668 319 14755 329
rect 14668 299 14677 319
rect 14697 299 14755 319
rect 14668 290 14755 299
rect 14668 289 14705 290
rect 14724 237 14755 290
rect 14785 319 14822 398
rect 14993 395 15386 415
rect 15406 395 15409 415
rect 14993 390 15409 395
rect 14993 389 15334 390
rect 14937 329 14968 330
rect 14785 299 14794 319
rect 14814 299 14822 319
rect 14785 289 14822 299
rect 14881 322 14968 329
rect 14881 319 14942 322
rect 14881 299 14890 319
rect 14910 302 14942 319
rect 14963 302 14968 322
rect 14910 299 14968 302
rect 14881 292 14968 299
rect 14993 319 15030 389
rect 15296 388 15333 389
rect 16678 380 16715 459
rect 16756 446 16866 459
rect 16830 390 16861 391
rect 16678 360 16687 380
rect 16707 360 16715 380
rect 16678 350 16715 360
rect 16774 380 16861 390
rect 16774 360 16783 380
rect 16803 360 16861 380
rect 16774 351 16861 360
rect 16774 350 16811 351
rect 15145 329 15181 330
rect 14993 299 15002 319
rect 15022 299 15030 319
rect 14881 290 14937 292
rect 14881 289 14918 290
rect 14993 289 15030 299
rect 15089 319 15237 329
rect 15337 326 15433 328
rect 15089 299 15098 319
rect 15118 299 15208 319
rect 15228 299 15237 319
rect 15089 290 15237 299
rect 15295 319 15433 326
rect 15295 299 15304 319
rect 15324 299 15433 319
rect 15295 290 15433 299
rect 16830 298 16861 351
rect 16891 380 16928 459
rect 17099 456 17492 476
rect 17512 456 17515 476
rect 17099 451 17515 456
rect 17099 450 17440 451
rect 17043 390 17074 391
rect 16891 360 16900 380
rect 16920 360 16928 380
rect 16891 350 16928 360
rect 16987 383 17074 390
rect 16987 380 17048 383
rect 16987 360 16996 380
rect 17016 363 17048 380
rect 17069 363 17074 383
rect 17016 360 17074 363
rect 16987 353 17074 360
rect 17099 380 17136 450
rect 17402 449 17439 450
rect 17251 390 17287 391
rect 17099 360 17108 380
rect 17128 360 17136 380
rect 16987 351 17043 353
rect 16987 350 17024 351
rect 17099 350 17136 360
rect 17195 380 17343 390
rect 17443 387 17539 389
rect 17195 360 17204 380
rect 17224 360 17314 380
rect 17334 360 17343 380
rect 17195 351 17343 360
rect 17401 380 17539 387
rect 17401 360 17410 380
rect 17430 360 17539 380
rect 17401 351 17539 360
rect 17195 350 17232 351
rect 17251 332 17287 351
rect 17306 350 17343 351
rect 17402 350 17439 351
rect 17248 307 17287 332
rect 17251 299 17287 307
rect 16722 297 16763 298
rect 16614 290 16763 297
rect 15089 289 15126 290
rect 15145 270 15181 290
rect 15200 289 15237 290
rect 15296 289 15333 290
rect 15135 241 15181 270
rect 15145 238 15181 241
rect 14616 236 14657 237
rect 14508 229 14657 236
rect 14508 209 14626 229
rect 14646 209 14657 229
rect 14508 201 14657 209
rect 14724 233 15083 237
rect 14724 228 15046 233
rect 14724 204 14837 228
rect 14861 209 15046 228
rect 15070 209 15083 233
rect 14861 204 15083 209
rect 14724 201 15083 204
rect 15145 201 15180 238
rect 15248 235 15348 238
rect 15248 231 15315 235
rect 15248 205 15260 231
rect 15286 209 15315 231
rect 15341 209 15348 235
rect 15286 205 15348 209
rect 15248 201 15348 205
rect 14724 180 14755 201
rect 15145 180 15181 201
rect 14567 179 14604 180
rect 14566 170 14604 179
rect 14566 150 14575 170
rect 14595 150 14604 170
rect 14566 142 14604 150
rect 14670 174 14755 180
rect 14780 179 14817 180
rect 14670 154 14678 174
rect 14698 154 14755 174
rect 14670 146 14755 154
rect 14779 170 14817 179
rect 14779 150 14788 170
rect 14808 150 14817 170
rect 14670 145 14706 146
rect 14779 142 14817 150
rect 14883 174 14968 180
rect 14988 179 15025 180
rect 14883 154 14891 174
rect 14911 173 14968 174
rect 14911 154 14940 173
rect 14883 153 14940 154
rect 14961 153 14968 173
rect 14883 146 14968 153
rect 14987 170 15025 179
rect 14987 150 14996 170
rect 15016 150 15025 170
rect 14883 145 14919 146
rect 14987 142 15025 150
rect 15091 174 15235 180
rect 15091 154 15099 174
rect 15119 173 15207 174
rect 15119 154 15137 173
rect 15091 149 15137 154
rect 15178 154 15207 173
rect 15227 154 15235 174
rect 15178 149 15235 154
rect 15091 146 15235 149
rect 15091 145 15127 146
rect 15199 145 15235 146
rect 15301 179 15338 180
rect 15301 178 15339 179
rect 15301 170 15365 178
rect 15301 150 15310 170
rect 15330 156 15365 170
rect 15385 156 15388 176
rect 15330 151 15388 156
rect 15330 150 15365 151
rect 12428 135 12556 141
rect 12428 132 12517 135
rect 12314 130 12517 132
rect 12038 114 12517 130
rect 12544 114 12556 135
rect 11699 103 11810 109
rect 12038 104 12556 114
rect 14567 113 14604 142
rect 12314 103 12556 104
rect 11699 95 11740 103
rect 11699 75 11707 95
rect 11726 75 11740 95
rect 11699 73 11740 75
rect 11768 95 11810 103
rect 12428 101 12556 103
rect 14568 111 14604 113
rect 14780 111 14817 142
rect 11768 75 11784 95
rect 11803 75 11810 95
rect 14568 89 14817 111
rect 14988 110 15025 142
rect 15301 138 15365 150
rect 15405 130 15432 290
rect 16614 270 16732 290
rect 16752 270 16763 290
rect 16614 262 16763 270
rect 16830 294 17189 298
rect 16830 289 17152 294
rect 16830 265 16943 289
rect 16967 270 17152 289
rect 17176 270 17189 294
rect 16967 265 17189 270
rect 16830 262 17189 265
rect 17251 262 17286 299
rect 17354 296 17454 299
rect 17354 292 17421 296
rect 17354 266 17366 292
rect 17392 270 17421 292
rect 17447 270 17454 296
rect 17392 266 17454 270
rect 17354 262 17454 266
rect 16830 241 16861 262
rect 17251 241 17287 262
rect 16673 240 16710 241
rect 16672 231 16710 240
rect 16672 211 16681 231
rect 16701 211 16710 231
rect 16672 203 16710 211
rect 16776 235 16861 241
rect 16886 240 16923 241
rect 16776 215 16784 235
rect 16804 215 16861 235
rect 16776 207 16861 215
rect 16885 231 16923 240
rect 16885 211 16894 231
rect 16914 211 16923 231
rect 16776 206 16812 207
rect 16885 203 16923 211
rect 16989 235 17074 241
rect 17094 240 17131 241
rect 16989 215 16997 235
rect 17017 234 17074 235
rect 17017 215 17046 234
rect 16989 214 17046 215
rect 17067 214 17074 234
rect 16989 207 17074 214
rect 17093 231 17131 240
rect 17093 211 17102 231
rect 17122 211 17131 231
rect 16989 206 17025 207
rect 17093 203 17131 211
rect 17197 235 17341 241
rect 17197 215 17205 235
rect 17225 233 17313 235
rect 17225 215 17252 233
rect 17197 213 17252 215
rect 17286 215 17313 233
rect 17333 215 17341 235
rect 17286 213 17341 215
rect 17197 207 17341 213
rect 17197 206 17233 207
rect 17305 206 17341 207
rect 17407 240 17444 241
rect 17407 239 17445 240
rect 17407 231 17471 239
rect 17407 211 17416 231
rect 17436 217 17471 231
rect 17491 217 17494 237
rect 17436 212 17494 217
rect 17436 211 17471 212
rect 16673 174 16710 203
rect 16674 172 16710 174
rect 16886 172 16923 203
rect 16674 150 16923 172
rect 17094 171 17131 203
rect 17407 199 17471 211
rect 17511 182 17538 351
rect 17484 176 17612 182
rect 17484 173 17573 176
rect 17370 171 17573 173
rect 17094 155 17573 171
rect 17600 155 17612 176
rect 16755 144 16866 150
rect 17094 145 17612 155
rect 17370 144 17612 145
rect 16755 136 16796 144
rect 15401 116 15524 130
rect 15401 112 15453 116
rect 15264 110 15453 112
rect 14988 90 15453 110
rect 15512 90 15524 116
rect 16755 116 16763 136
rect 16782 116 16796 136
rect 16755 114 16796 116
rect 16824 136 16866 144
rect 17484 142 17612 144
rect 16824 116 16840 136
rect 16859 116 16866 136
rect 16824 114 16866 116
rect 16755 99 16866 114
rect 11768 73 11810 75
rect 11699 58 11810 73
rect 14649 83 14760 89
rect 14988 84 15524 90
rect 15264 83 15524 84
rect 14649 75 14690 83
rect 14649 55 14657 75
rect 14676 55 14690 75
rect 14649 53 14690 55
rect 14718 75 14760 83
rect 15392 81 15524 83
rect 15435 79 15524 81
rect 14718 55 14734 75
rect 14753 55 14760 75
rect 14718 53 14760 55
rect 14649 38 14760 53
rect 10273 -9 10335 -2
rect 10167 -11 10335 -9
rect 9891 -12 10335 -11
rect 9552 -38 9663 -32
rect 9891 -37 10282 -12
rect 10167 -38 10282 -37
rect 9552 -46 9593 -38
rect 9552 -66 9560 -46
rect 9579 -66 9593 -46
rect 9552 -68 9593 -66
rect 9621 -46 9663 -38
rect 9621 -66 9637 -46
rect 9656 -66 9663 -46
rect 10273 -42 10282 -38
rect 10323 -38 10335 -12
rect 10323 -42 10333 -38
rect 10273 -52 10333 -42
rect 9621 -68 9663 -66
rect 9552 -83 9663 -68
<< viali >>
rect 4408 9332 4427 9352
rect 4485 9332 4504 9352
rect 423 9249 452 9276
rect 497 9252 526 9279
rect 193 9136 222 9165
rect 1155 9244 1175 9264
rect 711 9151 732 9171
rect 1084 9058 1110 9084
rect 709 9002 730 9022
rect 919 9002 944 9022
rect 1134 9005 1154 9025
rect 3776 9231 3796 9251
rect 3988 9236 4011 9256
rect 4200 9234 4221 9254
rect 3820 9172 3846 9198
rect 426 8904 445 8924
rect 503 8904 522 8924
rect 1361 9005 1390 9032
rect 1435 9008 1464 9035
rect 2093 9000 2113 9020
rect 1649 8907 1670 8927
rect 3204 8993 3230 9015
rect 3469 9022 3488 9042
rect 3546 9022 3565 9042
rect 4198 9085 4219 9105
rect 2022 8814 2048 8840
rect 1647 8758 1668 8778
rect 1862 8762 1882 8779
rect 2072 8761 2092 8781
rect 199 8695 224 8714
rect 422 8695 451 8722
rect 496 8698 525 8725
rect 1154 8690 1174 8710
rect 3755 8992 3775 9012
rect 9464 9373 9483 9393
rect 9541 9373 9560 9393
rect 5479 9290 5508 9317
rect 5553 9293 5582 9320
rect 5249 9177 5278 9206
rect 6211 9285 6231 9305
rect 5767 9192 5788 9212
rect 6140 9099 6166 9125
rect 5765 9043 5786 9063
rect 5975 9043 6000 9063
rect 6190 9046 6210 9066
rect 4404 8977 4433 9004
rect 4478 8980 4507 9007
rect 4705 8988 4730 9007
rect 2837 8921 2857 8941
rect 3261 8924 3282 8944
rect 8832 9272 8852 9292
rect 9044 9277 9067 9297
rect 9256 9275 9277 9295
rect 8876 9213 8902 9239
rect 5482 8945 5501 8965
rect 5559 8945 5578 8965
rect 6417 9046 6446 9073
rect 6491 9049 6520 9076
rect 2881 8862 2907 8888
rect 7149 9041 7169 9061
rect 6705 8948 6726 8968
rect 8260 9034 8286 9056
rect 8525 9063 8544 9083
rect 8602 9063 8621 9083
rect 9254 9126 9275 9146
rect 3048 8783 3069 8824
rect 710 8597 731 8617
rect 1364 8660 1383 8680
rect 1441 8660 1460 8680
rect 1699 8687 1725 8709
rect 3259 8775 3280 8795
rect 2816 8682 2836 8702
rect 3189 8689 3221 8706
rect 7078 8855 7104 8881
rect 3465 8667 3494 8694
rect 3539 8670 3568 8697
rect 4407 8778 4426 8798
rect 4484 8778 4503 8798
rect 1083 8504 1109 8530
rect 708 8448 729 8468
rect 918 8446 941 8466
rect 1133 8451 1153 8471
rect 6703 8799 6724 8819
rect 6918 8803 6938 8820
rect 7128 8802 7148 8822
rect 5255 8736 5280 8755
rect 5478 8736 5507 8763
rect 5552 8739 5581 8766
rect 3775 8677 3795 8697
rect 3985 8680 4010 8700
rect 4199 8680 4220 8700
rect 3819 8618 3845 8644
rect 3041 8483 3072 8510
rect 3329 8511 3348 8531
rect 3406 8511 3425 8531
rect 425 8350 444 8370
rect 502 8350 521 8370
rect 1502 8413 1531 8440
rect 1576 8416 1605 8443
rect 1860 8407 1880 8424
rect 2234 8408 2254 8428
rect 1790 8315 1811 8335
rect 2163 8222 2189 8248
rect 424 8146 453 8173
rect 498 8149 527 8176
rect 194 8033 223 8062
rect 1156 8141 1176 8161
rect 1788 8166 1809 8186
rect 1996 8164 2023 8185
rect 2213 8169 2233 8189
rect 712 8048 733 8068
rect 4197 8531 4218 8551
rect 2697 8410 2717 8430
rect 3121 8413 3142 8433
rect 3754 8438 3774 8458
rect 4707 8537 4736 8566
rect 4403 8423 4432 8450
rect 4477 8426 4506 8453
rect 2741 8351 2767 8377
rect 2908 8271 2931 8309
rect 3119 8264 3140 8284
rect 2676 8171 2696 8191
rect 3050 8175 3070 8192
rect 3325 8156 3354 8183
rect 3399 8159 3428 8186
rect 4409 8229 4428 8249
rect 4486 8229 4505 8249
rect 1505 8068 1524 8088
rect 1582 8068 1601 8088
rect 1858 8089 1889 8116
rect 1085 7955 1111 7981
rect 710 7899 731 7919
rect 920 7899 945 7919
rect 1135 7902 1155 7922
rect 3777 8128 3797 8148
rect 3989 8133 4012 8153
rect 4201 8131 4222 8151
rect 3821 8069 3847 8095
rect 427 7801 446 7821
rect 504 7801 523 7821
rect 1362 7902 1391 7929
rect 1436 7905 1465 7932
rect 1709 7893 1741 7910
rect 2094 7897 2114 7917
rect 1650 7804 1671 7824
rect 3205 7890 3231 7912
rect 3470 7919 3489 7939
rect 3547 7919 3566 7939
rect 4199 7982 4220 8002
rect 1861 7775 1882 7816
rect 2023 7711 2049 7737
rect 1648 7655 1669 7675
rect 2073 7658 2093 7678
rect 200 7592 225 7611
rect 423 7592 452 7619
rect 497 7595 526 7622
rect 1155 7587 1175 7607
rect 3756 7889 3776 7909
rect 6210 8731 6230 8751
rect 8811 9033 8831 9053
rect 14439 9337 14458 9357
rect 14516 9337 14535 9357
rect 10454 9254 10483 9281
rect 10528 9257 10557 9284
rect 10224 9141 10253 9170
rect 11186 9249 11206 9269
rect 10742 9156 10763 9176
rect 9460 9018 9489 9045
rect 9534 9021 9563 9048
rect 11115 9063 11141 9089
rect 9761 9029 9786 9048
rect 7893 8962 7913 8982
rect 8317 8965 8338 8985
rect 10740 9007 10761 9027
rect 10950 9007 10975 9027
rect 11165 9010 11185 9030
rect 7937 8903 7963 8929
rect 13807 9236 13827 9256
rect 14019 9241 14042 9261
rect 14231 9239 14252 9259
rect 13851 9177 13877 9203
rect 8104 8824 8125 8865
rect 5766 8638 5787 8658
rect 6420 8701 6439 8721
rect 6497 8701 6516 8721
rect 6755 8728 6781 8750
rect 8315 8816 8336 8836
rect 7872 8723 7892 8743
rect 8245 8730 8277 8747
rect 8521 8708 8550 8735
rect 8595 8711 8624 8738
rect 9463 8819 9482 8839
rect 9540 8819 9559 8839
rect 10457 8909 10476 8929
rect 10534 8909 10553 8929
rect 11392 9010 11421 9037
rect 11466 9013 11495 9040
rect 12124 9005 12144 9025
rect 11680 8912 11701 8932
rect 13235 8998 13261 9020
rect 13500 9027 13519 9047
rect 13577 9027 13596 9047
rect 14229 9090 14250 9110
rect 6139 8545 6165 8571
rect 5764 8489 5785 8509
rect 5974 8487 5997 8507
rect 6189 8492 6209 8512
rect 12053 8819 12079 8845
rect 8831 8718 8851 8738
rect 9041 8721 9066 8741
rect 9255 8721 9276 8741
rect 11678 8763 11699 8783
rect 11893 8767 11913 8784
rect 12103 8766 12123 8786
rect 10230 8700 10255 8719
rect 8875 8659 8901 8685
rect 10453 8700 10482 8727
rect 10527 8703 10556 8730
rect 8097 8524 8128 8551
rect 8385 8552 8404 8572
rect 8462 8552 8481 8572
rect 5481 8391 5500 8411
rect 5558 8391 5577 8411
rect 6558 8454 6587 8481
rect 6632 8457 6661 8484
rect 6916 8448 6936 8465
rect 7290 8449 7310 8469
rect 6846 8356 6867 8376
rect 7219 8263 7245 8289
rect 5480 8187 5509 8214
rect 5554 8190 5583 8217
rect 5250 8074 5279 8103
rect 6212 8182 6232 8202
rect 6844 8207 6865 8227
rect 7052 8205 7079 8226
rect 7269 8210 7289 8230
rect 5768 8089 5789 8109
rect 9253 8572 9274 8592
rect 7753 8451 7773 8471
rect 8177 8454 8198 8474
rect 8810 8479 8830 8499
rect 9763 8578 9792 8607
rect 9459 8464 9488 8491
rect 9533 8467 9562 8494
rect 7797 8392 7823 8418
rect 7964 8312 7987 8350
rect 8175 8305 8196 8325
rect 7732 8212 7752 8232
rect 8106 8216 8126 8233
rect 8381 8197 8410 8224
rect 8455 8200 8484 8227
rect 9465 8270 9484 8290
rect 9542 8270 9561 8290
rect 6561 8109 6580 8129
rect 6638 8109 6657 8129
rect 6914 8130 6945 8157
rect 6141 7996 6167 8022
rect 5766 7940 5787 7960
rect 5976 7940 6001 7960
rect 6191 7943 6211 7963
rect 4405 7874 4434 7901
rect 4479 7877 4508 7904
rect 4706 7885 4731 7904
rect 2838 7818 2858 7838
rect 3048 7820 3068 7837
rect 3262 7821 3283 7841
rect 8833 8169 8853 8189
rect 9045 8174 9068 8194
rect 9257 8172 9278 8192
rect 8877 8110 8903 8136
rect 5483 7842 5502 7862
rect 5560 7842 5579 7862
rect 6418 7943 6447 7970
rect 6492 7946 6521 7973
rect 2882 7759 2908 7785
rect 6765 7934 6797 7951
rect 7150 7938 7170 7958
rect 6706 7845 6727 7865
rect 8261 7931 8287 7953
rect 8526 7960 8545 7980
rect 8603 7960 8622 7980
rect 9255 8023 9276 8043
rect 6917 7816 6938 7857
rect 711 7494 732 7514
rect 1365 7557 1384 7577
rect 1442 7557 1461 7577
rect 1700 7584 1726 7606
rect 3260 7672 3281 7692
rect 2817 7579 2837 7599
rect 7079 7752 7105 7778
rect 3466 7564 3495 7591
rect 3540 7567 3569 7594
rect 4408 7675 4427 7695
rect 4485 7675 4504 7695
rect 1084 7401 1110 7427
rect 709 7345 730 7365
rect 919 7343 942 7363
rect 1134 7348 1154 7368
rect 6704 7696 6725 7716
rect 7129 7699 7149 7719
rect 5256 7633 5281 7652
rect 5479 7633 5508 7660
rect 5553 7636 5582 7663
rect 3776 7574 3796 7594
rect 3986 7577 4011 7597
rect 4200 7577 4221 7597
rect 3820 7515 3846 7541
rect 2707 7367 2755 7396
rect 3360 7395 3379 7415
rect 3437 7395 3456 7415
rect 426 7247 445 7267
rect 503 7247 522 7267
rect 1472 7323 1501 7350
rect 1546 7326 1575 7353
rect 2204 7318 2224 7338
rect 1760 7225 1781 7245
rect 2133 7132 2159 7158
rect 424 7043 453 7070
rect 498 7046 527 7073
rect 1758 7076 1779 7096
rect 1966 7076 1995 7095
rect 2183 7079 2203 7099
rect 194 6930 223 6959
rect 1156 7038 1176 7058
rect 712 6945 733 6965
rect 4198 7428 4219 7448
rect 3755 7335 3775 7355
rect 4708 7434 4737 7463
rect 2728 7294 2748 7314
rect 3152 7297 3173 7317
rect 4404 7320 4433 7347
rect 4478 7323 4507 7350
rect 2772 7235 2798 7261
rect 6211 7628 6231 7648
rect 8812 7930 8832 7950
rect 11185 8695 11205 8715
rect 13786 8997 13806 9017
rect 19495 9378 19514 9398
rect 19572 9378 19591 9398
rect 15510 9295 15539 9322
rect 15584 9298 15613 9325
rect 15280 9182 15309 9211
rect 16242 9290 16262 9310
rect 15798 9197 15819 9217
rect 16171 9104 16197 9130
rect 15796 9048 15817 9068
rect 16006 9048 16031 9068
rect 16221 9051 16241 9071
rect 14435 8982 14464 9009
rect 14509 8985 14538 9012
rect 14736 8993 14761 9012
rect 12868 8926 12888 8946
rect 13292 8929 13313 8949
rect 18863 9277 18883 9297
rect 19075 9282 19098 9302
rect 19287 9280 19308 9300
rect 18907 9218 18933 9244
rect 15513 8950 15532 8970
rect 15590 8950 15609 8970
rect 16448 9051 16477 9078
rect 16522 9054 16551 9081
rect 12912 8867 12938 8893
rect 17180 9046 17200 9066
rect 16736 8953 16757 8973
rect 18291 9039 18317 9061
rect 18556 9068 18575 9088
rect 18633 9068 18652 9088
rect 19285 9131 19306 9151
rect 13079 8788 13100 8829
rect 10741 8602 10762 8622
rect 11395 8665 11414 8685
rect 11472 8665 11491 8685
rect 11730 8692 11756 8714
rect 13290 8780 13311 8800
rect 12847 8687 12867 8707
rect 13220 8694 13252 8711
rect 17109 8860 17135 8886
rect 13496 8672 13525 8699
rect 13570 8675 13599 8702
rect 14438 8783 14457 8803
rect 14515 8783 14534 8803
rect 11114 8509 11140 8535
rect 10739 8453 10760 8473
rect 10949 8451 10972 8471
rect 11164 8456 11184 8476
rect 16734 8804 16755 8824
rect 16949 8808 16969 8825
rect 17159 8807 17179 8827
rect 15286 8741 15311 8760
rect 15509 8741 15538 8768
rect 15583 8744 15612 8771
rect 13806 8682 13826 8702
rect 14016 8685 14041 8705
rect 14230 8685 14251 8705
rect 13850 8623 13876 8649
rect 13072 8488 13103 8515
rect 13360 8516 13379 8536
rect 13437 8516 13456 8536
rect 10456 8355 10475 8375
rect 10533 8355 10552 8375
rect 11533 8418 11562 8445
rect 11607 8421 11636 8448
rect 11891 8412 11911 8429
rect 12265 8413 12285 8433
rect 11821 8320 11842 8340
rect 12194 8227 12220 8253
rect 10455 8151 10484 8178
rect 10529 8154 10558 8181
rect 10225 8038 10254 8067
rect 11187 8146 11207 8166
rect 11819 8171 11840 8191
rect 12027 8169 12054 8190
rect 12244 8174 12264 8194
rect 10743 8053 10764 8073
rect 14228 8536 14249 8556
rect 12728 8415 12748 8435
rect 13152 8418 13173 8438
rect 13785 8443 13805 8463
rect 14738 8542 14767 8571
rect 14434 8428 14463 8455
rect 14508 8431 14537 8458
rect 12772 8356 12798 8382
rect 12939 8276 12962 8314
rect 13150 8269 13171 8289
rect 12707 8176 12727 8196
rect 13081 8180 13101 8197
rect 13356 8161 13385 8188
rect 13430 8164 13459 8191
rect 14440 8234 14459 8254
rect 14517 8234 14536 8254
rect 11536 8073 11555 8093
rect 11613 8073 11632 8093
rect 11889 8094 11920 8121
rect 9461 7915 9490 7942
rect 9535 7918 9564 7945
rect 11116 7960 11142 7986
rect 9762 7926 9787 7945
rect 7894 7859 7914 7879
rect 8104 7861 8124 7878
rect 8318 7862 8339 7882
rect 10741 7904 10762 7924
rect 10951 7904 10976 7924
rect 11166 7907 11186 7927
rect 7938 7800 7964 7826
rect 13808 8133 13828 8153
rect 14020 8138 14043 8158
rect 14232 8136 14253 8156
rect 13852 8074 13878 8100
rect 5767 7535 5788 7555
rect 6421 7598 6440 7618
rect 6498 7598 6517 7618
rect 6756 7625 6782 7647
rect 8316 7713 8337 7733
rect 7873 7620 7893 7640
rect 8522 7605 8551 7632
rect 8596 7608 8625 7635
rect 9464 7716 9483 7736
rect 9541 7716 9560 7736
rect 10458 7806 10477 7826
rect 10535 7806 10554 7826
rect 11393 7907 11422 7934
rect 11467 7910 11496 7937
rect 11740 7898 11772 7915
rect 12125 7902 12145 7922
rect 11681 7809 11702 7829
rect 13236 7895 13262 7917
rect 13501 7924 13520 7944
rect 13578 7924 13597 7944
rect 14230 7987 14251 8007
rect 11892 7780 11913 7821
rect 6140 7442 6166 7468
rect 5765 7386 5786 7406
rect 5975 7384 5998 7404
rect 6190 7389 6210 7409
rect 12054 7716 12080 7742
rect 8832 7615 8852 7635
rect 9042 7618 9067 7638
rect 9256 7618 9277 7638
rect 11679 7660 11700 7680
rect 12104 7663 12124 7683
rect 10231 7597 10256 7616
rect 8876 7556 8902 7582
rect 10454 7597 10483 7624
rect 10528 7600 10557 7627
rect 7763 7408 7811 7437
rect 8416 7436 8435 7456
rect 8493 7436 8512 7456
rect 5482 7288 5501 7308
rect 5559 7288 5578 7308
rect 2937 7160 2964 7192
rect 3150 7148 3171 7168
rect 2707 7057 2727 7075
rect 3097 7053 3118 7073
rect 3356 7040 3385 7067
rect 3430 7043 3459 7070
rect 6528 7364 6557 7391
rect 6602 7367 6631 7394
rect 7260 7359 7280 7379
rect 6816 7266 6837 7286
rect 4409 7126 4428 7146
rect 4486 7126 4505 7146
rect 1475 6978 1494 6998
rect 1552 6978 1571 6998
rect 1085 6852 1111 6878
rect 710 6796 731 6816
rect 920 6796 945 6816
rect 1135 6799 1155 6819
rect 3777 7025 3797 7045
rect 3989 7030 4012 7050
rect 4201 7028 4222 7048
rect 3821 6966 3847 6992
rect 2176 6857 2224 6886
rect 427 6698 446 6718
rect 504 6698 523 6718
rect 1362 6799 1391 6826
rect 1436 6802 1465 6829
rect 2094 6794 2114 6814
rect 1650 6701 1671 6721
rect 3205 6787 3231 6809
rect 3470 6816 3489 6836
rect 3547 6816 3566 6836
rect 4199 6879 4220 6899
rect 2023 6608 2049 6634
rect 1648 6552 1669 6572
rect 1863 6556 1883 6573
rect 2073 6555 2093 6575
rect 200 6489 225 6508
rect 423 6489 452 6516
rect 497 6492 526 6519
rect 1155 6484 1175 6504
rect 3756 6786 3776 6806
rect 7189 7173 7215 7199
rect 5480 7084 5509 7111
rect 5554 7087 5583 7114
rect 6814 7117 6835 7137
rect 7022 7117 7051 7136
rect 7239 7120 7259 7140
rect 5250 6971 5279 7000
rect 6212 7079 6232 7099
rect 5768 6986 5789 7006
rect 9254 7469 9275 7489
rect 8811 7376 8831 7396
rect 9764 7475 9793 7504
rect 7784 7335 7804 7355
rect 8208 7338 8229 7358
rect 9460 7361 9489 7388
rect 9534 7364 9563 7391
rect 7828 7276 7854 7302
rect 7993 7201 8020 7233
rect 8206 7189 8227 7209
rect 7763 7098 7783 7116
rect 8153 7094 8174 7114
rect 8412 7081 8441 7108
rect 8486 7084 8515 7111
rect 9465 7167 9484 7187
rect 9542 7167 9561 7187
rect 6531 7019 6550 7039
rect 6608 7019 6627 7039
rect 6141 6893 6167 6919
rect 5766 6837 5787 6857
rect 5976 6837 6001 6857
rect 6191 6840 6211 6860
rect 4405 6771 4434 6798
rect 4479 6774 4508 6801
rect 4706 6782 4731 6801
rect 2838 6715 2858 6735
rect 3262 6718 3283 6738
rect 8833 7066 8853 7086
rect 9045 7071 9068 7091
rect 9257 7069 9278 7089
rect 8877 7007 8903 7033
rect 7232 6898 7280 6927
rect 5483 6739 5502 6759
rect 5560 6739 5579 6759
rect 6418 6840 6447 6867
rect 6492 6843 6521 6870
rect 2882 6656 2908 6682
rect 7150 6835 7170 6855
rect 6706 6742 6727 6762
rect 8261 6828 8287 6850
rect 8526 6857 8545 6877
rect 8603 6857 8622 6877
rect 9255 6920 9276 6940
rect 3049 6577 3070 6618
rect 711 6391 732 6411
rect 1365 6454 1384 6474
rect 1442 6454 1461 6474
rect 1700 6481 1726 6503
rect 3260 6569 3281 6589
rect 2817 6476 2837 6496
rect 3190 6483 3222 6500
rect 7079 6649 7105 6675
rect 3466 6461 3495 6488
rect 3540 6464 3569 6491
rect 4408 6572 4427 6592
rect 4485 6572 4504 6592
rect 1084 6298 1110 6324
rect 709 6242 730 6262
rect 919 6240 942 6260
rect 1134 6245 1154 6265
rect 6704 6593 6725 6613
rect 6919 6597 6939 6614
rect 7129 6596 7149 6616
rect 5256 6530 5281 6549
rect 5479 6530 5508 6557
rect 5553 6533 5582 6560
rect 3776 6471 3796 6491
rect 3986 6474 4011 6494
rect 4200 6474 4221 6494
rect 3820 6412 3846 6438
rect 3042 6277 3073 6304
rect 3330 6305 3349 6325
rect 3407 6305 3426 6325
rect 426 6144 445 6164
rect 503 6144 522 6164
rect 1503 6207 1532 6234
rect 1577 6210 1606 6237
rect 1861 6201 1881 6218
rect 2235 6202 2255 6222
rect 1791 6109 1812 6129
rect 2000 6084 2023 6122
rect 2164 6016 2190 6042
rect 425 5940 454 5967
rect 499 5943 528 5970
rect 195 5827 224 5856
rect 1157 5935 1177 5955
rect 1789 5960 1810 5980
rect 2214 5963 2234 5983
rect 713 5842 734 5862
rect 4198 6325 4219 6345
rect 2698 6204 2718 6224
rect 2908 6208 2935 6229
rect 3122 6207 3143 6227
rect 3755 6232 3775 6252
rect 4708 6331 4737 6360
rect 4404 6217 4433 6244
rect 4478 6220 4507 6247
rect 2742 6145 2768 6171
rect 3120 6058 3141 6078
rect 2677 5965 2697 5985
rect 3051 5969 3071 5986
rect 3326 5950 3355 5977
rect 3400 5953 3429 5980
rect 4410 6023 4429 6043
rect 4487 6023 4506 6043
rect 1506 5862 1525 5882
rect 1583 5862 1602 5882
rect 1859 5883 1890 5910
rect 1086 5749 1112 5775
rect 711 5693 732 5713
rect 921 5693 946 5713
rect 1136 5696 1156 5716
rect 3778 5922 3798 5942
rect 3990 5927 4013 5947
rect 4202 5925 4223 5945
rect 3822 5863 3848 5889
rect 428 5595 447 5615
rect 505 5595 524 5615
rect 1363 5696 1392 5723
rect 1437 5699 1466 5726
rect 1710 5687 1742 5704
rect 2095 5691 2115 5711
rect 1651 5598 1672 5618
rect 3206 5684 3232 5706
rect 3471 5713 3490 5733
rect 3548 5713 3567 5733
rect 4200 5776 4221 5796
rect 1862 5569 1883 5610
rect 2024 5505 2050 5531
rect 1649 5449 1670 5469
rect 2074 5452 2094 5472
rect 201 5386 226 5405
rect 424 5386 453 5413
rect 498 5389 527 5416
rect 1156 5381 1176 5401
rect 3757 5683 3777 5703
rect 6211 6525 6231 6545
rect 8812 6827 8832 6847
rect 11186 7592 11206 7612
rect 13787 7894 13807 7914
rect 16241 8736 16261 8756
rect 18842 9038 18862 9058
rect 19491 9023 19520 9050
rect 19565 9026 19594 9053
rect 19792 9034 19817 9053
rect 17924 8967 17944 8987
rect 18348 8970 18369 8990
rect 17968 8908 17994 8934
rect 18135 8829 18156 8870
rect 15797 8643 15818 8663
rect 16451 8706 16470 8726
rect 16528 8706 16547 8726
rect 16786 8733 16812 8755
rect 18346 8821 18367 8841
rect 17903 8728 17923 8748
rect 18276 8735 18308 8752
rect 18552 8713 18581 8740
rect 18626 8716 18655 8743
rect 19494 8824 19513 8844
rect 19571 8824 19590 8844
rect 16170 8550 16196 8576
rect 15795 8494 15816 8514
rect 16005 8492 16028 8512
rect 16220 8497 16240 8517
rect 18862 8723 18882 8743
rect 19072 8726 19097 8746
rect 19286 8726 19307 8746
rect 18906 8664 18932 8690
rect 18128 8529 18159 8556
rect 18416 8557 18435 8577
rect 18493 8557 18512 8577
rect 15512 8396 15531 8416
rect 15589 8396 15608 8416
rect 16589 8459 16618 8486
rect 16663 8462 16692 8489
rect 16947 8453 16967 8470
rect 17321 8454 17341 8474
rect 16877 8361 16898 8381
rect 17250 8268 17276 8294
rect 15511 8192 15540 8219
rect 15585 8195 15614 8222
rect 15281 8079 15310 8108
rect 16243 8187 16263 8207
rect 16875 8212 16896 8232
rect 17083 8210 17110 8231
rect 17300 8215 17320 8235
rect 15799 8094 15820 8114
rect 19284 8577 19305 8597
rect 17784 8456 17804 8476
rect 18208 8459 18229 8479
rect 18841 8484 18861 8504
rect 19794 8583 19823 8612
rect 19490 8469 19519 8496
rect 19564 8472 19593 8499
rect 17828 8397 17854 8423
rect 17995 8317 18018 8355
rect 18206 8310 18227 8330
rect 17763 8217 17783 8237
rect 18137 8221 18157 8238
rect 18412 8202 18441 8229
rect 18486 8205 18515 8232
rect 19496 8275 19515 8295
rect 19573 8275 19592 8295
rect 16592 8114 16611 8134
rect 16669 8114 16688 8134
rect 16945 8135 16976 8162
rect 16172 8001 16198 8027
rect 15797 7945 15818 7965
rect 16007 7945 16032 7965
rect 16222 7948 16242 7968
rect 14436 7879 14465 7906
rect 14510 7882 14539 7909
rect 14737 7890 14762 7909
rect 12869 7823 12889 7843
rect 13079 7825 13099 7842
rect 13293 7826 13314 7846
rect 18864 8174 18884 8194
rect 19076 8179 19099 8199
rect 19288 8177 19309 8197
rect 18908 8115 18934 8141
rect 15514 7847 15533 7867
rect 15591 7847 15610 7867
rect 16449 7948 16478 7975
rect 16523 7951 16552 7978
rect 12913 7764 12939 7790
rect 16796 7939 16828 7956
rect 17181 7943 17201 7963
rect 16737 7850 16758 7870
rect 18292 7936 18318 7958
rect 18557 7965 18576 7985
rect 18634 7965 18653 7985
rect 19286 8028 19307 8048
rect 16948 7821 16969 7862
rect 10742 7499 10763 7519
rect 11396 7562 11415 7582
rect 11473 7562 11492 7582
rect 11731 7589 11757 7611
rect 13291 7677 13312 7697
rect 12848 7584 12868 7604
rect 17110 7757 17136 7783
rect 13497 7569 13526 7596
rect 13571 7572 13600 7599
rect 14439 7680 14458 7700
rect 14516 7680 14535 7700
rect 11115 7406 11141 7432
rect 10740 7350 10761 7370
rect 10950 7348 10973 7368
rect 11165 7353 11185 7373
rect 16735 7701 16756 7721
rect 17160 7704 17180 7724
rect 15287 7638 15312 7657
rect 15510 7638 15539 7665
rect 15584 7641 15613 7668
rect 13807 7579 13827 7599
rect 14017 7582 14042 7602
rect 14231 7582 14252 7602
rect 13851 7520 13877 7546
rect 12738 7372 12786 7401
rect 13391 7400 13410 7420
rect 13468 7400 13487 7420
rect 10457 7252 10476 7272
rect 10534 7252 10553 7272
rect 11503 7328 11532 7355
rect 11577 7331 11606 7358
rect 12235 7323 12255 7343
rect 11791 7230 11812 7250
rect 12164 7137 12190 7163
rect 10455 7048 10484 7075
rect 10529 7051 10558 7078
rect 11789 7081 11810 7101
rect 11997 7081 12026 7100
rect 12214 7084 12234 7104
rect 10225 6935 10254 6964
rect 11187 7043 11207 7063
rect 10743 6950 10764 6970
rect 14229 7433 14250 7453
rect 13786 7340 13806 7360
rect 14739 7439 14768 7468
rect 12759 7299 12779 7319
rect 13183 7302 13204 7322
rect 14435 7325 14464 7352
rect 14509 7328 14538 7355
rect 12803 7240 12829 7266
rect 16242 7633 16262 7653
rect 18843 7935 18863 7955
rect 19492 7920 19521 7947
rect 19566 7923 19595 7950
rect 19793 7931 19818 7950
rect 17925 7864 17945 7884
rect 18135 7866 18155 7883
rect 18349 7867 18370 7887
rect 17969 7805 17995 7831
rect 15798 7540 15819 7560
rect 16452 7603 16471 7623
rect 16529 7603 16548 7623
rect 16787 7630 16813 7652
rect 18347 7718 18368 7738
rect 17904 7625 17924 7645
rect 18553 7610 18582 7637
rect 18627 7613 18656 7640
rect 19495 7721 19514 7741
rect 19572 7721 19591 7741
rect 16171 7447 16197 7473
rect 15796 7391 15817 7411
rect 16006 7389 16029 7409
rect 16221 7394 16241 7414
rect 18863 7620 18883 7640
rect 19073 7623 19098 7643
rect 19287 7623 19308 7643
rect 18907 7561 18933 7587
rect 17794 7413 17842 7442
rect 18447 7441 18466 7461
rect 18524 7441 18543 7461
rect 15513 7293 15532 7313
rect 15590 7293 15609 7313
rect 12968 7165 12995 7197
rect 13181 7153 13202 7173
rect 12738 7062 12758 7080
rect 13128 7058 13149 7078
rect 13387 7045 13416 7072
rect 13461 7048 13490 7075
rect 16559 7369 16588 7396
rect 16633 7372 16662 7399
rect 17291 7364 17311 7384
rect 16847 7271 16868 7291
rect 14440 7131 14459 7151
rect 14517 7131 14536 7151
rect 11506 6983 11525 7003
rect 11583 6983 11602 7003
rect 9461 6812 9490 6839
rect 9535 6815 9564 6842
rect 11116 6857 11142 6883
rect 9762 6823 9787 6842
rect 7894 6756 7914 6776
rect 8318 6759 8339 6779
rect 10741 6801 10762 6821
rect 10951 6801 10976 6821
rect 11166 6804 11186 6824
rect 7938 6697 7964 6723
rect 13808 7030 13828 7050
rect 14020 7035 14043 7055
rect 14232 7033 14253 7053
rect 13852 6971 13878 6997
rect 12207 6862 12255 6891
rect 8105 6618 8126 6659
rect 5767 6432 5788 6452
rect 6421 6495 6440 6515
rect 6498 6495 6517 6515
rect 6756 6522 6782 6544
rect 8316 6610 8337 6630
rect 7873 6517 7893 6537
rect 8246 6524 8278 6541
rect 8522 6502 8551 6529
rect 8596 6505 8625 6532
rect 9464 6613 9483 6633
rect 9541 6613 9560 6633
rect 10458 6703 10477 6723
rect 10535 6703 10554 6723
rect 11393 6804 11422 6831
rect 11467 6807 11496 6834
rect 12125 6799 12145 6819
rect 11681 6706 11702 6726
rect 13236 6792 13262 6814
rect 13501 6821 13520 6841
rect 13578 6821 13597 6841
rect 14230 6884 14251 6904
rect 6140 6339 6166 6365
rect 5765 6283 5786 6303
rect 5975 6281 5998 6301
rect 6190 6286 6210 6306
rect 12054 6613 12080 6639
rect 8832 6512 8852 6532
rect 9042 6515 9067 6535
rect 9256 6515 9277 6535
rect 11679 6557 11700 6577
rect 11894 6561 11914 6578
rect 12104 6560 12124 6580
rect 10231 6494 10256 6513
rect 8876 6453 8902 6479
rect 10454 6494 10483 6521
rect 10528 6497 10557 6524
rect 8098 6318 8129 6345
rect 8386 6346 8405 6366
rect 8463 6346 8482 6366
rect 5482 6185 5501 6205
rect 5559 6185 5578 6205
rect 6559 6248 6588 6275
rect 6633 6251 6662 6278
rect 6917 6242 6937 6259
rect 7291 6243 7311 6263
rect 6847 6150 6868 6170
rect 7056 6125 7079 6163
rect 7220 6057 7246 6083
rect 5481 5981 5510 6008
rect 5555 5984 5584 6011
rect 5251 5868 5280 5897
rect 6213 5976 6233 5996
rect 6845 6001 6866 6021
rect 7270 6004 7290 6024
rect 5769 5883 5790 5903
rect 9254 6366 9275 6386
rect 7754 6245 7774 6265
rect 7964 6249 7991 6270
rect 8178 6248 8199 6268
rect 8811 6273 8831 6293
rect 9764 6372 9793 6401
rect 9460 6258 9489 6285
rect 9534 6261 9563 6288
rect 7798 6186 7824 6212
rect 8176 6099 8197 6119
rect 7733 6006 7753 6026
rect 8107 6010 8127 6027
rect 8382 5991 8411 6018
rect 8456 5994 8485 6021
rect 9466 6064 9485 6084
rect 9543 6064 9562 6084
rect 6562 5903 6581 5923
rect 6639 5903 6658 5923
rect 6915 5924 6946 5951
rect 6142 5790 6168 5816
rect 5767 5734 5788 5754
rect 5977 5734 6002 5754
rect 6192 5737 6212 5757
rect 4406 5668 4435 5695
rect 4480 5671 4509 5698
rect 4707 5679 4732 5698
rect 2839 5612 2859 5632
rect 3049 5614 3069 5631
rect 3263 5615 3284 5635
rect 8834 5963 8854 5983
rect 9046 5968 9069 5988
rect 9258 5966 9279 5986
rect 8878 5904 8904 5930
rect 5484 5636 5503 5656
rect 5561 5636 5580 5656
rect 6419 5737 6448 5764
rect 6493 5740 6522 5767
rect 2883 5553 2909 5579
rect 6766 5728 6798 5745
rect 7151 5732 7171 5752
rect 6707 5639 6728 5659
rect 8262 5725 8288 5747
rect 8527 5754 8546 5774
rect 8604 5754 8623 5774
rect 9256 5817 9277 5837
rect 6918 5610 6939 5651
rect 712 5288 733 5308
rect 1366 5351 1385 5371
rect 1443 5351 1462 5371
rect 1701 5378 1727 5400
rect 3261 5466 3282 5486
rect 2818 5373 2838 5393
rect 7080 5546 7106 5572
rect 3467 5358 3496 5385
rect 3541 5361 3570 5388
rect 4409 5469 4428 5489
rect 4486 5469 4505 5489
rect 2567 5300 2594 5340
rect 1085 5195 1111 5221
rect 710 5139 731 5159
rect 920 5137 943 5157
rect 1135 5142 1155 5162
rect 6705 5490 6726 5510
rect 7130 5493 7150 5513
rect 5257 5427 5282 5446
rect 5480 5427 5509 5454
rect 5554 5430 5583 5457
rect 3777 5368 3797 5388
rect 3987 5371 4012 5391
rect 4201 5371 4222 5391
rect 3821 5309 3847 5335
rect 3362 5183 3381 5203
rect 3439 5183 3458 5203
rect 427 5041 446 5061
rect 504 5041 523 5061
rect 1472 5123 1501 5150
rect 1546 5126 1575 5153
rect 2204 5118 2224 5138
rect 1760 5025 1781 5045
rect 2133 4932 2159 4958
rect 425 4837 454 4864
rect 499 4840 528 4867
rect 1758 4876 1779 4896
rect 1966 4875 1992 4899
rect 2183 4879 2203 4899
rect 195 4724 224 4753
rect 1157 4832 1177 4852
rect 713 4739 734 4759
rect 4199 5222 4220 5242
rect 3756 5129 3776 5149
rect 4709 5228 4738 5257
rect 2730 5082 2750 5102
rect 2937 5085 2962 5105
rect 3154 5085 3175 5105
rect 4405 5114 4434 5141
rect 4479 5117 4508 5144
rect 2774 5023 2800 5049
rect 6212 5422 6232 5442
rect 8813 5724 8833 5744
rect 11186 6489 11206 6509
rect 13787 6791 13807 6811
rect 17220 7178 17246 7204
rect 15511 7089 15540 7116
rect 15585 7092 15614 7119
rect 16845 7122 16866 7142
rect 17053 7122 17082 7141
rect 17270 7125 17290 7145
rect 15281 6976 15310 7005
rect 16243 7084 16263 7104
rect 15799 6991 15820 7011
rect 19285 7474 19306 7494
rect 18842 7381 18862 7401
rect 19795 7480 19824 7509
rect 17815 7340 17835 7360
rect 18239 7343 18260 7363
rect 19491 7366 19520 7393
rect 19565 7369 19594 7396
rect 17859 7281 17885 7307
rect 18024 7206 18051 7238
rect 18237 7194 18258 7214
rect 17794 7103 17814 7121
rect 18184 7099 18205 7119
rect 18443 7086 18472 7113
rect 18517 7089 18546 7116
rect 19496 7172 19515 7192
rect 19573 7172 19592 7192
rect 16562 7024 16581 7044
rect 16639 7024 16658 7044
rect 16172 6898 16198 6924
rect 15797 6842 15818 6862
rect 16007 6842 16032 6862
rect 16222 6845 16242 6865
rect 14436 6776 14465 6803
rect 14510 6779 14539 6806
rect 14737 6787 14762 6806
rect 12869 6720 12889 6740
rect 13293 6723 13314 6743
rect 18864 7071 18884 7091
rect 19076 7076 19099 7096
rect 19288 7074 19309 7094
rect 18908 7012 18934 7038
rect 17263 6903 17311 6932
rect 15514 6744 15533 6764
rect 15591 6744 15610 6764
rect 16449 6845 16478 6872
rect 16523 6848 16552 6875
rect 12913 6661 12939 6687
rect 17181 6840 17201 6860
rect 16737 6747 16758 6767
rect 18292 6833 18318 6855
rect 18557 6862 18576 6882
rect 18634 6862 18653 6882
rect 19286 6925 19307 6945
rect 13080 6582 13101 6623
rect 10742 6396 10763 6416
rect 11396 6459 11415 6479
rect 11473 6459 11492 6479
rect 11731 6486 11757 6508
rect 13291 6574 13312 6594
rect 12848 6481 12868 6501
rect 13221 6488 13253 6505
rect 17110 6654 17136 6680
rect 13497 6466 13526 6493
rect 13571 6469 13600 6496
rect 14439 6577 14458 6597
rect 14516 6577 14535 6597
rect 11115 6303 11141 6329
rect 10740 6247 10761 6267
rect 10950 6245 10973 6265
rect 11165 6250 11185 6270
rect 16735 6598 16756 6618
rect 16950 6602 16970 6619
rect 17160 6601 17180 6621
rect 15287 6535 15312 6554
rect 15510 6535 15539 6562
rect 15584 6538 15613 6565
rect 13807 6476 13827 6496
rect 14017 6479 14042 6499
rect 14231 6479 14252 6499
rect 13851 6417 13877 6443
rect 13073 6282 13104 6309
rect 13361 6310 13380 6330
rect 13438 6310 13457 6330
rect 10457 6149 10476 6169
rect 10534 6149 10553 6169
rect 11534 6212 11563 6239
rect 11608 6215 11637 6242
rect 11892 6206 11912 6223
rect 12266 6207 12286 6227
rect 11822 6114 11843 6134
rect 12031 6089 12054 6127
rect 12195 6021 12221 6047
rect 10456 5945 10485 5972
rect 10530 5948 10559 5975
rect 10226 5832 10255 5861
rect 11188 5940 11208 5960
rect 11820 5965 11841 5985
rect 12245 5968 12265 5988
rect 10744 5847 10765 5867
rect 14229 6330 14250 6350
rect 12729 6209 12749 6229
rect 12939 6213 12966 6234
rect 13153 6212 13174 6232
rect 13786 6237 13806 6257
rect 14739 6336 14768 6365
rect 14435 6222 14464 6249
rect 14509 6225 14538 6252
rect 12773 6150 12799 6176
rect 13151 6063 13172 6083
rect 12708 5970 12728 5990
rect 13082 5974 13102 5991
rect 13357 5955 13386 5982
rect 13431 5958 13460 5985
rect 14441 6028 14460 6048
rect 14518 6028 14537 6048
rect 11537 5867 11556 5887
rect 11614 5867 11633 5887
rect 11890 5888 11921 5915
rect 9462 5709 9491 5736
rect 9536 5712 9565 5739
rect 11117 5754 11143 5780
rect 9763 5720 9788 5739
rect 7895 5653 7915 5673
rect 8105 5655 8125 5672
rect 8319 5656 8340 5676
rect 10742 5698 10763 5718
rect 10952 5698 10977 5718
rect 11167 5701 11187 5721
rect 7939 5594 7965 5620
rect 13809 5927 13829 5947
rect 14021 5932 14044 5952
rect 14233 5930 14254 5950
rect 13853 5868 13879 5894
rect 5768 5329 5789 5349
rect 6422 5392 6441 5412
rect 6499 5392 6518 5412
rect 6757 5419 6783 5441
rect 8317 5507 8338 5527
rect 7874 5414 7894 5434
rect 8523 5399 8552 5426
rect 8597 5402 8626 5429
rect 9465 5510 9484 5530
rect 9542 5510 9561 5530
rect 10459 5600 10478 5620
rect 10536 5600 10555 5620
rect 11394 5701 11423 5728
rect 11468 5704 11497 5731
rect 11741 5692 11773 5709
rect 12126 5696 12146 5716
rect 11682 5603 11703 5623
rect 13237 5689 13263 5711
rect 13502 5718 13521 5738
rect 13579 5718 13598 5738
rect 14231 5781 14252 5801
rect 11893 5574 11914 5615
rect 7623 5341 7650 5381
rect 6141 5236 6167 5262
rect 5766 5180 5787 5200
rect 5976 5178 5999 5198
rect 6191 5183 6211 5203
rect 12055 5510 12081 5536
rect 8833 5409 8853 5429
rect 9043 5412 9068 5432
rect 9257 5412 9278 5432
rect 11680 5454 11701 5474
rect 12105 5457 12125 5477
rect 10232 5391 10257 5410
rect 8877 5350 8903 5376
rect 10455 5391 10484 5418
rect 10529 5394 10558 5421
rect 8418 5224 8437 5244
rect 8495 5224 8514 5244
rect 3152 4936 3173 4956
rect 2709 4843 2729 4863
rect 5483 5082 5502 5102
rect 5560 5082 5579 5102
rect 6528 5164 6557 5191
rect 6602 5167 6631 5194
rect 3358 4828 3387 4855
rect 3432 4831 3461 4858
rect 4410 4920 4429 4940
rect 4487 4920 4506 4940
rect 7260 5159 7280 5179
rect 6816 5066 6837 5086
rect 1475 4778 1494 4798
rect 1552 4778 1571 4798
rect 1086 4646 1112 4672
rect 711 4590 732 4610
rect 921 4590 946 4610
rect 1136 4593 1156 4613
rect 3778 4819 3798 4839
rect 3990 4824 4013 4844
rect 4202 4822 4223 4842
rect 3822 4760 3848 4786
rect 2339 4641 2366 4681
rect 428 4492 447 4512
rect 505 4492 524 4512
rect 1363 4593 1392 4620
rect 1437 4596 1466 4623
rect 2095 4588 2115 4608
rect 1651 4495 1672 4515
rect 3206 4581 3232 4603
rect 3471 4610 3490 4630
rect 3548 4610 3567 4630
rect 4200 4673 4221 4693
rect 2024 4402 2050 4428
rect 1649 4346 1670 4366
rect 1864 4350 1884 4367
rect 2074 4349 2094 4369
rect 201 4283 226 4302
rect 424 4283 453 4310
rect 498 4286 527 4313
rect 1156 4278 1176 4298
rect 3757 4580 3777 4600
rect 7189 4973 7215 4999
rect 5481 4878 5510 4905
rect 5555 4881 5584 4908
rect 6814 4917 6835 4937
rect 7022 4916 7048 4940
rect 7239 4920 7259 4940
rect 5251 4765 5280 4794
rect 6213 4873 6233 4893
rect 5769 4780 5790 4800
rect 9255 5263 9276 5283
rect 8812 5170 8832 5190
rect 9765 5269 9794 5298
rect 7786 5123 7806 5143
rect 7993 5126 8018 5146
rect 8210 5126 8231 5146
rect 9461 5155 9490 5182
rect 9535 5158 9564 5185
rect 7830 5064 7856 5090
rect 8208 4977 8229 4997
rect 7765 4884 7785 4904
rect 11187 5386 11207 5406
rect 13788 5688 13808 5708
rect 16242 6530 16262 6550
rect 18843 6832 18863 6852
rect 19492 6817 19521 6844
rect 19566 6820 19595 6847
rect 19793 6828 19818 6847
rect 17925 6761 17945 6781
rect 18349 6764 18370 6784
rect 17969 6702 17995 6728
rect 18136 6623 18157 6664
rect 15798 6437 15819 6457
rect 16452 6500 16471 6520
rect 16529 6500 16548 6520
rect 16787 6527 16813 6549
rect 18347 6615 18368 6635
rect 17904 6522 17924 6542
rect 18277 6529 18309 6546
rect 18553 6507 18582 6534
rect 18627 6510 18656 6537
rect 19495 6618 19514 6638
rect 19572 6618 19591 6638
rect 16171 6344 16197 6370
rect 15796 6288 15817 6308
rect 16006 6286 16029 6306
rect 16221 6291 16241 6311
rect 18863 6517 18883 6537
rect 19073 6520 19098 6540
rect 19287 6520 19308 6540
rect 18907 6458 18933 6484
rect 18129 6323 18160 6350
rect 18417 6351 18436 6371
rect 18494 6351 18513 6371
rect 15513 6190 15532 6210
rect 15590 6190 15609 6210
rect 16590 6253 16619 6280
rect 16664 6256 16693 6283
rect 16948 6247 16968 6264
rect 17322 6248 17342 6268
rect 16878 6155 16899 6175
rect 17087 6130 17110 6168
rect 17251 6062 17277 6088
rect 15512 5986 15541 6013
rect 15586 5989 15615 6016
rect 15282 5873 15311 5902
rect 16244 5981 16264 6001
rect 16876 6006 16897 6026
rect 17301 6009 17321 6029
rect 15800 5888 15821 5908
rect 19285 6371 19306 6391
rect 17785 6250 17805 6270
rect 17995 6254 18022 6275
rect 18209 6253 18230 6273
rect 18842 6278 18862 6298
rect 19795 6377 19824 6406
rect 19491 6263 19520 6290
rect 19565 6266 19594 6293
rect 17829 6191 17855 6217
rect 18207 6104 18228 6124
rect 17764 6011 17784 6031
rect 18138 6015 18158 6032
rect 18413 5996 18442 6023
rect 18487 5999 18516 6026
rect 19497 6069 19516 6089
rect 19574 6069 19593 6089
rect 16593 5908 16612 5928
rect 16670 5908 16689 5928
rect 16946 5929 16977 5956
rect 16173 5795 16199 5821
rect 15798 5739 15819 5759
rect 16008 5739 16033 5759
rect 16223 5742 16243 5762
rect 14437 5673 14466 5700
rect 14511 5676 14540 5703
rect 14738 5684 14763 5703
rect 12870 5617 12890 5637
rect 13080 5619 13100 5636
rect 13294 5620 13315 5640
rect 18865 5968 18885 5988
rect 19077 5973 19100 5993
rect 19289 5971 19310 5991
rect 18909 5909 18935 5935
rect 15515 5641 15534 5661
rect 15592 5641 15611 5661
rect 16450 5742 16479 5769
rect 16524 5745 16553 5772
rect 12914 5558 12940 5584
rect 16797 5733 16829 5750
rect 17182 5737 17202 5757
rect 16738 5644 16759 5664
rect 18293 5730 18319 5752
rect 18558 5759 18577 5779
rect 18635 5759 18654 5779
rect 19287 5822 19308 5842
rect 16949 5615 16970 5656
rect 10743 5293 10764 5313
rect 11397 5356 11416 5376
rect 11474 5356 11493 5376
rect 11732 5383 11758 5405
rect 13292 5471 13313 5491
rect 12849 5378 12869 5398
rect 17111 5551 17137 5577
rect 13498 5363 13527 5390
rect 13572 5366 13601 5393
rect 14440 5474 14459 5494
rect 14517 5474 14536 5494
rect 12598 5305 12625 5345
rect 11116 5200 11142 5226
rect 10741 5144 10762 5164
rect 10951 5142 10974 5162
rect 11166 5147 11186 5167
rect 16736 5495 16757 5515
rect 17161 5498 17181 5518
rect 15288 5432 15313 5451
rect 15511 5432 15540 5459
rect 15585 5435 15614 5462
rect 13808 5373 13828 5393
rect 14018 5376 14043 5396
rect 14232 5376 14253 5396
rect 13852 5314 13878 5340
rect 13393 5188 13412 5208
rect 13470 5188 13489 5208
rect 8414 4869 8443 4896
rect 8488 4872 8517 4899
rect 9466 4961 9485 4981
rect 9543 4961 9562 4981
rect 10458 5046 10477 5066
rect 10535 5046 10554 5066
rect 11503 5128 11532 5155
rect 11577 5131 11606 5158
rect 6531 4819 6550 4839
rect 6608 4819 6627 4839
rect 6142 4687 6168 4713
rect 5767 4631 5788 4651
rect 5977 4631 6002 4651
rect 6192 4634 6212 4654
rect 4406 4565 4435 4592
rect 4480 4568 4509 4595
rect 4707 4576 4732 4595
rect 2839 4509 2859 4529
rect 3263 4512 3284 4532
rect 8834 4860 8854 4880
rect 9046 4865 9069 4885
rect 9258 4863 9279 4883
rect 8878 4801 8904 4827
rect 7395 4682 7422 4722
rect 5484 4533 5503 4553
rect 5561 4533 5580 4553
rect 6419 4634 6448 4661
rect 6493 4637 6522 4664
rect 2883 4450 2909 4476
rect 7151 4629 7171 4649
rect 6707 4536 6728 4556
rect 8262 4622 8288 4644
rect 8527 4651 8546 4671
rect 8604 4651 8623 4671
rect 9256 4714 9277 4734
rect 3050 4371 3071 4412
rect 712 4185 733 4205
rect 1366 4248 1385 4268
rect 1443 4248 1462 4268
rect 1701 4275 1727 4297
rect 3261 4363 3282 4383
rect 2818 4270 2838 4290
rect 3191 4277 3223 4294
rect 7080 4443 7106 4469
rect 3467 4255 3496 4282
rect 3541 4258 3570 4285
rect 4409 4366 4428 4386
rect 4486 4366 4505 4386
rect 1085 4092 1111 4118
rect 710 4036 731 4056
rect 920 4034 943 4054
rect 1135 4039 1155 4059
rect 6705 4387 6726 4407
rect 6920 4391 6940 4408
rect 7130 4390 7150 4410
rect 5257 4324 5282 4343
rect 5480 4324 5509 4351
rect 5554 4327 5583 4354
rect 3777 4265 3797 4285
rect 3987 4268 4012 4288
rect 4201 4268 4222 4288
rect 3821 4206 3847 4232
rect 3043 4071 3074 4098
rect 3331 4099 3350 4119
rect 3408 4099 3427 4119
rect 427 3938 446 3958
rect 504 3938 523 3958
rect 1504 4001 1533 4028
rect 1578 4004 1607 4031
rect 1862 3995 1882 4012
rect 2236 3996 2256 4016
rect 1792 3903 1813 3923
rect 2165 3810 2191 3836
rect 426 3734 455 3761
rect 500 3737 529 3764
rect 196 3621 225 3650
rect 1158 3729 1178 3749
rect 1790 3754 1811 3774
rect 1998 3752 2025 3773
rect 2215 3757 2235 3777
rect 714 3636 735 3656
rect 4199 4119 4220 4139
rect 2699 3998 2719 4018
rect 3123 4001 3144 4021
rect 3756 4026 3776 4046
rect 4709 4125 4738 4154
rect 4405 4011 4434 4038
rect 4479 4014 4508 4041
rect 2743 3939 2769 3965
rect 2910 3859 2933 3897
rect 3121 3852 3142 3872
rect 2678 3759 2698 3779
rect 3052 3763 3072 3780
rect 3327 3744 3356 3771
rect 3401 3747 3430 3774
rect 4411 3817 4430 3837
rect 4488 3817 4507 3837
rect 1507 3656 1526 3676
rect 1584 3656 1603 3676
rect 1860 3677 1891 3704
rect 1087 3543 1113 3569
rect 712 3487 733 3507
rect 922 3487 947 3507
rect 1137 3490 1157 3510
rect 3779 3716 3799 3736
rect 3991 3721 4014 3741
rect 4203 3719 4224 3739
rect 3823 3657 3849 3683
rect 429 3389 448 3409
rect 506 3389 525 3409
rect 1364 3490 1393 3517
rect 1438 3493 1467 3520
rect 1711 3481 1743 3498
rect 2096 3485 2116 3505
rect 1652 3392 1673 3412
rect 3207 3478 3233 3500
rect 3472 3507 3491 3527
rect 3549 3507 3568 3527
rect 4201 3570 4222 3590
rect 1863 3363 1884 3404
rect 2025 3299 2051 3325
rect 1650 3243 1671 3263
rect 2075 3246 2095 3266
rect 202 3180 227 3199
rect 425 3180 454 3207
rect 499 3183 528 3210
rect 1157 3175 1177 3195
rect 3758 3477 3778 3497
rect 6212 4319 6232 4339
rect 8813 4621 8833 4641
rect 12235 5123 12255 5143
rect 11791 5030 11812 5050
rect 12164 4937 12190 4963
rect 10456 4842 10485 4869
rect 10530 4845 10559 4872
rect 11789 4881 11810 4901
rect 11997 4880 12023 4904
rect 12214 4884 12234 4904
rect 10226 4729 10255 4758
rect 11188 4837 11208 4857
rect 10744 4744 10765 4764
rect 14230 5227 14251 5247
rect 13787 5134 13807 5154
rect 14740 5233 14769 5262
rect 12761 5087 12781 5107
rect 12968 5090 12993 5110
rect 13185 5090 13206 5110
rect 14436 5119 14465 5146
rect 14510 5122 14539 5149
rect 12805 5028 12831 5054
rect 16243 5427 16263 5447
rect 18844 5729 18864 5749
rect 19493 5714 19522 5741
rect 19567 5717 19596 5744
rect 19794 5725 19819 5744
rect 17926 5658 17946 5678
rect 18136 5660 18156 5677
rect 18350 5661 18371 5681
rect 17970 5599 17996 5625
rect 15799 5334 15820 5354
rect 16453 5397 16472 5417
rect 16530 5397 16549 5417
rect 16788 5424 16814 5446
rect 18348 5512 18369 5532
rect 17905 5419 17925 5439
rect 18554 5404 18583 5431
rect 18628 5407 18657 5434
rect 19496 5515 19515 5535
rect 19573 5515 19592 5535
rect 17654 5346 17681 5386
rect 16172 5241 16198 5267
rect 15797 5185 15818 5205
rect 16007 5183 16030 5203
rect 16222 5188 16242 5208
rect 18864 5414 18884 5434
rect 19074 5417 19099 5437
rect 19288 5417 19309 5437
rect 18908 5355 18934 5381
rect 18449 5229 18468 5249
rect 18526 5229 18545 5249
rect 13183 4941 13204 4961
rect 12740 4848 12760 4868
rect 15514 5087 15533 5107
rect 15591 5087 15610 5107
rect 16559 5169 16588 5196
rect 16633 5172 16662 5199
rect 13389 4833 13418 4860
rect 13463 4836 13492 4863
rect 14441 4925 14460 4945
rect 14518 4925 14537 4945
rect 17291 5164 17311 5184
rect 16847 5071 16868 5091
rect 11506 4783 11525 4803
rect 11583 4783 11602 4803
rect 9462 4606 9491 4633
rect 9536 4609 9565 4636
rect 11117 4651 11143 4677
rect 9763 4617 9788 4636
rect 7895 4550 7915 4570
rect 8319 4553 8340 4573
rect 10742 4595 10763 4615
rect 10952 4595 10977 4615
rect 11167 4598 11187 4618
rect 7939 4491 7965 4517
rect 13809 4824 13829 4844
rect 14021 4829 14044 4849
rect 14233 4827 14254 4847
rect 13853 4765 13879 4791
rect 12370 4646 12397 4686
rect 8106 4412 8127 4453
rect 5768 4226 5789 4246
rect 6422 4289 6441 4309
rect 6499 4289 6518 4309
rect 6757 4316 6783 4338
rect 8317 4404 8338 4424
rect 7874 4311 7894 4331
rect 8247 4318 8279 4335
rect 8523 4296 8552 4323
rect 8597 4299 8626 4326
rect 9465 4407 9484 4427
rect 9542 4407 9561 4427
rect 10459 4497 10478 4517
rect 10536 4497 10555 4517
rect 11394 4598 11423 4625
rect 11468 4601 11497 4628
rect 12126 4593 12146 4613
rect 11682 4500 11703 4520
rect 13237 4586 13263 4608
rect 13502 4615 13521 4635
rect 13579 4615 13598 4635
rect 14231 4678 14252 4698
rect 6141 4133 6167 4159
rect 5766 4077 5787 4097
rect 5976 4075 5999 4095
rect 6191 4080 6211 4100
rect 12055 4407 12081 4433
rect 8833 4306 8853 4326
rect 9043 4309 9068 4329
rect 9257 4309 9278 4329
rect 11680 4351 11701 4371
rect 11895 4355 11915 4372
rect 12105 4354 12125 4374
rect 10232 4288 10257 4307
rect 8877 4247 8903 4273
rect 10455 4288 10484 4315
rect 10529 4291 10558 4318
rect 8099 4112 8130 4139
rect 8387 4140 8406 4160
rect 8464 4140 8483 4160
rect 5483 3979 5502 3999
rect 5560 3979 5579 3999
rect 6560 4042 6589 4069
rect 6634 4045 6663 4072
rect 6918 4036 6938 4053
rect 7292 4037 7312 4057
rect 6848 3944 6869 3964
rect 7221 3851 7247 3877
rect 5482 3775 5511 3802
rect 5556 3778 5585 3805
rect 5252 3662 5281 3691
rect 6214 3770 6234 3790
rect 6846 3795 6867 3815
rect 7054 3793 7081 3814
rect 7271 3798 7291 3818
rect 5770 3677 5791 3697
rect 9255 4160 9276 4180
rect 7755 4039 7775 4059
rect 8179 4042 8200 4062
rect 8812 4067 8832 4087
rect 9765 4166 9794 4195
rect 9461 4052 9490 4079
rect 9535 4055 9564 4082
rect 7799 3980 7825 4006
rect 7966 3900 7989 3938
rect 8177 3893 8198 3913
rect 7734 3800 7754 3820
rect 8108 3804 8128 3821
rect 8383 3785 8412 3812
rect 8457 3788 8486 3815
rect 9467 3858 9486 3878
rect 9544 3858 9563 3878
rect 6563 3697 6582 3717
rect 6640 3697 6659 3717
rect 6916 3718 6947 3745
rect 6143 3584 6169 3610
rect 5768 3528 5789 3548
rect 5978 3528 6003 3548
rect 6193 3531 6213 3551
rect 4407 3462 4436 3489
rect 4481 3465 4510 3492
rect 4708 3473 4733 3492
rect 2840 3406 2860 3426
rect 3050 3408 3070 3425
rect 3264 3409 3285 3429
rect 8835 3757 8855 3777
rect 9047 3762 9070 3782
rect 9259 3760 9280 3780
rect 8879 3698 8905 3724
rect 5485 3430 5504 3450
rect 5562 3430 5581 3450
rect 6420 3531 6449 3558
rect 6494 3534 6523 3561
rect 2884 3347 2910 3373
rect 6767 3522 6799 3539
rect 7152 3526 7172 3546
rect 6708 3433 6729 3453
rect 8263 3519 8289 3541
rect 8528 3548 8547 3568
rect 8605 3548 8624 3568
rect 9257 3611 9278 3631
rect 6919 3404 6940 3445
rect 713 3082 734 3102
rect 1367 3145 1386 3165
rect 1444 3145 1463 3165
rect 1702 3172 1728 3194
rect 3262 3260 3283 3280
rect 2819 3167 2839 3187
rect 7081 3340 7107 3366
rect 3468 3152 3497 3179
rect 3542 3155 3571 3182
rect 4410 3263 4429 3283
rect 4487 3263 4506 3283
rect 2709 3095 2757 3124
rect 1086 2989 1112 3015
rect 711 2933 732 2953
rect 921 2931 944 2951
rect 1136 2936 1156 2956
rect 6706 3284 6727 3304
rect 7131 3287 7151 3307
rect 5258 3221 5283 3240
rect 5481 3221 5510 3248
rect 5555 3224 5584 3251
rect 3778 3162 3798 3182
rect 3988 3165 4013 3185
rect 4202 3165 4223 3185
rect 3822 3103 3848 3129
rect 3362 2983 3381 3003
rect 3439 2983 3458 3003
rect 428 2835 447 2855
rect 505 2835 524 2855
rect 1474 2911 1503 2938
rect 1548 2914 1577 2941
rect 1815 2908 1836 2928
rect 2206 2906 2226 2924
rect 1762 2813 1783 2833
rect 1969 2789 1996 2821
rect 2135 2720 2161 2746
rect 426 2631 455 2658
rect 500 2634 529 2661
rect 1760 2664 1781 2684
rect 2185 2667 2205 2687
rect 196 2518 225 2547
rect 1158 2626 1178 2646
rect 714 2533 735 2553
rect 4200 3016 4221 3036
rect 3757 2923 3777 2943
rect 4710 3022 4739 3051
rect 2730 2882 2750 2902
rect 2938 2886 2967 2905
rect 3154 2885 3175 2905
rect 4406 2908 4435 2935
rect 4480 2911 4509 2938
rect 2774 2823 2800 2849
rect 6213 3216 6233 3236
rect 8814 3518 8834 3538
rect 11187 4283 11207 4303
rect 13788 4585 13808 4605
rect 17220 4978 17246 5004
rect 15512 4883 15541 4910
rect 15586 4886 15615 4913
rect 16845 4922 16866 4942
rect 17053 4921 17079 4945
rect 17270 4925 17290 4945
rect 15282 4770 15311 4799
rect 16244 4878 16264 4898
rect 15800 4785 15821 4805
rect 19286 5268 19307 5288
rect 18843 5175 18863 5195
rect 19796 5274 19825 5303
rect 17817 5128 17837 5148
rect 18024 5131 18049 5151
rect 18241 5131 18262 5151
rect 19492 5160 19521 5187
rect 19566 5163 19595 5190
rect 17861 5069 17887 5095
rect 18239 4982 18260 5002
rect 17796 4889 17816 4909
rect 18445 4874 18474 4901
rect 18519 4877 18548 4904
rect 19497 4966 19516 4986
rect 19574 4966 19593 4986
rect 16562 4824 16581 4844
rect 16639 4824 16658 4844
rect 16173 4692 16199 4718
rect 15798 4636 15819 4656
rect 16008 4636 16033 4656
rect 16223 4639 16243 4659
rect 14437 4570 14466 4597
rect 14511 4573 14540 4600
rect 14738 4581 14763 4600
rect 12870 4514 12890 4534
rect 13294 4517 13315 4537
rect 18865 4865 18885 4885
rect 19077 4870 19100 4890
rect 19289 4868 19310 4888
rect 18909 4806 18935 4832
rect 17426 4687 17453 4727
rect 15515 4538 15534 4558
rect 15592 4538 15611 4558
rect 16450 4639 16479 4666
rect 16524 4642 16553 4669
rect 12914 4455 12940 4481
rect 17182 4634 17202 4654
rect 16738 4541 16759 4561
rect 18293 4627 18319 4649
rect 18558 4656 18577 4676
rect 18635 4656 18654 4676
rect 19287 4719 19308 4739
rect 13081 4376 13102 4417
rect 10743 4190 10764 4210
rect 11397 4253 11416 4273
rect 11474 4253 11493 4273
rect 11732 4280 11758 4302
rect 13292 4368 13313 4388
rect 12849 4275 12869 4295
rect 13222 4282 13254 4299
rect 17111 4448 17137 4474
rect 13498 4260 13527 4287
rect 13572 4263 13601 4290
rect 14440 4371 14459 4391
rect 14517 4371 14536 4391
rect 11116 4097 11142 4123
rect 10741 4041 10762 4061
rect 10951 4039 10974 4059
rect 11166 4044 11186 4064
rect 16736 4392 16757 4412
rect 16951 4396 16971 4413
rect 17161 4395 17181 4415
rect 15288 4329 15313 4348
rect 15511 4329 15540 4356
rect 15585 4332 15614 4359
rect 13808 4270 13828 4290
rect 14018 4273 14043 4293
rect 14232 4273 14253 4293
rect 13852 4211 13878 4237
rect 13074 4076 13105 4103
rect 13362 4104 13381 4124
rect 13439 4104 13458 4124
rect 10458 3943 10477 3963
rect 10535 3943 10554 3963
rect 11535 4006 11564 4033
rect 11609 4009 11638 4036
rect 11893 4000 11913 4017
rect 12267 4001 12287 4021
rect 11823 3908 11844 3928
rect 12196 3815 12222 3841
rect 10457 3739 10486 3766
rect 10531 3742 10560 3769
rect 10227 3626 10256 3655
rect 11189 3734 11209 3754
rect 11821 3759 11842 3779
rect 12029 3757 12056 3778
rect 12246 3762 12266 3782
rect 10745 3641 10766 3661
rect 14230 4124 14251 4144
rect 12730 4003 12750 4023
rect 13154 4006 13175 4026
rect 13787 4031 13807 4051
rect 14740 4130 14769 4159
rect 14436 4016 14465 4043
rect 14510 4019 14539 4046
rect 12774 3944 12800 3970
rect 12941 3864 12964 3902
rect 13152 3857 13173 3877
rect 12709 3764 12729 3784
rect 13083 3768 13103 3785
rect 13358 3749 13387 3776
rect 13432 3752 13461 3779
rect 14442 3822 14461 3842
rect 14519 3822 14538 3842
rect 11538 3661 11557 3681
rect 11615 3661 11634 3681
rect 11891 3682 11922 3709
rect 9463 3503 9492 3530
rect 9537 3506 9566 3533
rect 11118 3548 11144 3574
rect 9764 3514 9789 3533
rect 7896 3447 7916 3467
rect 8106 3449 8126 3466
rect 8320 3450 8341 3470
rect 10743 3492 10764 3512
rect 10953 3492 10978 3512
rect 11168 3495 11188 3515
rect 7940 3388 7966 3414
rect 13810 3721 13830 3741
rect 14022 3726 14045 3746
rect 14234 3724 14255 3744
rect 13854 3662 13880 3688
rect 5769 3123 5790 3143
rect 6423 3186 6442 3206
rect 6500 3186 6519 3206
rect 6758 3213 6784 3235
rect 8318 3301 8339 3321
rect 7875 3208 7895 3228
rect 8524 3193 8553 3220
rect 8598 3196 8627 3223
rect 9466 3304 9485 3324
rect 9543 3304 9562 3324
rect 10460 3394 10479 3414
rect 10537 3394 10556 3414
rect 11395 3495 11424 3522
rect 11469 3498 11498 3525
rect 11742 3486 11774 3503
rect 12127 3490 12147 3510
rect 11683 3397 11704 3417
rect 13238 3483 13264 3505
rect 13503 3512 13522 3532
rect 13580 3512 13599 3532
rect 14232 3575 14253 3595
rect 11894 3368 11915 3409
rect 7765 3136 7813 3165
rect 6142 3030 6168 3056
rect 5767 2974 5788 2994
rect 5977 2972 6000 2992
rect 6192 2977 6212 2997
rect 12056 3304 12082 3330
rect 8834 3203 8854 3223
rect 9044 3206 9069 3226
rect 9258 3206 9279 3226
rect 11681 3248 11702 3268
rect 12106 3251 12126 3271
rect 10233 3185 10258 3204
rect 8878 3144 8904 3170
rect 10456 3185 10485 3212
rect 10530 3188 10559 3215
rect 8418 3024 8437 3044
rect 8495 3024 8514 3044
rect 5484 2876 5503 2896
rect 5561 2876 5580 2896
rect 3152 2736 3173 2756
rect 2709 2643 2729 2663
rect 3358 2628 3387 2655
rect 3432 2631 3461 2658
rect 6530 2952 6559 2979
rect 6604 2955 6633 2982
rect 6871 2949 6892 2969
rect 7262 2947 7282 2965
rect 6818 2854 6839 2874
rect 7025 2830 7052 2862
rect 4411 2714 4430 2734
rect 4488 2714 4507 2734
rect 1477 2566 1496 2586
rect 1554 2566 1573 2586
rect 2178 2585 2226 2614
rect 1087 2440 1113 2466
rect 712 2384 733 2404
rect 922 2384 947 2404
rect 1137 2387 1157 2407
rect 3779 2613 3799 2633
rect 3991 2618 4014 2638
rect 4203 2616 4224 2636
rect 3823 2554 3849 2580
rect 429 2286 448 2306
rect 506 2286 525 2306
rect 1364 2387 1393 2414
rect 1438 2390 1467 2417
rect 2096 2382 2116 2402
rect 1652 2289 1673 2309
rect 3207 2375 3233 2397
rect 3472 2404 3491 2424
rect 3549 2404 3568 2424
rect 4201 2467 4222 2487
rect 2025 2196 2051 2222
rect 1650 2140 1671 2160
rect 1865 2144 1885 2161
rect 2075 2143 2095 2163
rect 202 2077 227 2096
rect 425 2077 454 2104
rect 499 2080 528 2107
rect 1157 2072 1177 2092
rect 3758 2374 3778 2394
rect 7191 2761 7217 2787
rect 5482 2672 5511 2699
rect 5556 2675 5585 2702
rect 6816 2705 6837 2725
rect 7241 2708 7261 2728
rect 5252 2559 5281 2588
rect 6214 2667 6234 2687
rect 5770 2574 5791 2594
rect 9256 3057 9277 3077
rect 8813 2964 8833 2984
rect 9766 3063 9795 3092
rect 7786 2923 7806 2943
rect 7994 2927 8023 2946
rect 8210 2926 8231 2946
rect 9462 2949 9491 2976
rect 9536 2952 9565 2979
rect 7830 2864 7856 2890
rect 8208 2777 8229 2797
rect 7765 2684 7785 2704
rect 8414 2669 8443 2696
rect 8488 2672 8517 2699
rect 9467 2755 9486 2775
rect 9544 2755 9563 2775
rect 6533 2607 6552 2627
rect 6610 2607 6629 2627
rect 7234 2626 7282 2655
rect 6143 2481 6169 2507
rect 5768 2425 5789 2445
rect 5978 2425 6003 2445
rect 6193 2428 6213 2448
rect 4407 2359 4436 2386
rect 4481 2362 4510 2389
rect 4708 2370 4733 2389
rect 2840 2303 2860 2323
rect 3264 2306 3285 2326
rect 8835 2654 8855 2674
rect 9047 2659 9070 2679
rect 9259 2657 9280 2677
rect 8879 2595 8905 2621
rect 5485 2327 5504 2347
rect 5562 2327 5581 2347
rect 6420 2428 6449 2455
rect 6494 2431 6523 2458
rect 2884 2244 2910 2270
rect 7152 2423 7172 2443
rect 6708 2330 6729 2350
rect 8263 2416 8289 2438
rect 8528 2445 8547 2465
rect 8605 2445 8624 2465
rect 9257 2508 9278 2528
rect 3051 2165 3072 2206
rect 713 1979 734 1999
rect 1367 2042 1386 2062
rect 1444 2042 1463 2062
rect 1702 2069 1728 2091
rect 3262 2157 3283 2177
rect 2819 2064 2839 2084
rect 3192 2071 3224 2088
rect 7081 2237 7107 2263
rect 3468 2049 3497 2076
rect 3542 2052 3571 2079
rect 4410 2160 4429 2180
rect 4487 2160 4506 2180
rect 1086 1886 1112 1912
rect 711 1830 732 1850
rect 921 1828 944 1848
rect 1136 1833 1156 1853
rect 6706 2181 6727 2201
rect 6921 2185 6941 2202
rect 7131 2184 7151 2204
rect 5258 2118 5283 2137
rect 5481 2118 5510 2145
rect 5555 2121 5584 2148
rect 3778 2059 3798 2079
rect 3988 2062 4013 2082
rect 4202 2062 4223 2082
rect 3822 2000 3848 2026
rect 3044 1865 3075 1892
rect 3332 1893 3351 1913
rect 3409 1893 3428 1913
rect 428 1732 447 1752
rect 505 1732 524 1752
rect 1505 1795 1534 1822
rect 1579 1798 1608 1825
rect 1863 1789 1883 1806
rect 2237 1790 2257 1810
rect 1793 1697 1814 1717
rect 2002 1672 2025 1710
rect 2166 1604 2192 1630
rect 427 1528 456 1555
rect 501 1531 530 1558
rect 197 1415 226 1444
rect 1159 1523 1179 1543
rect 1791 1548 1812 1568
rect 2216 1551 2236 1571
rect 715 1430 736 1450
rect 4200 1913 4221 1933
rect 2700 1792 2720 1812
rect 2910 1796 2937 1817
rect 3124 1795 3145 1815
rect 3757 1820 3777 1840
rect 4710 1919 4739 1948
rect 4406 1805 4435 1832
rect 4480 1808 4509 1835
rect 2744 1733 2770 1759
rect 3122 1646 3143 1666
rect 2679 1553 2699 1573
rect 3053 1557 3073 1574
rect 3328 1538 3357 1565
rect 3402 1541 3431 1568
rect 4412 1611 4431 1631
rect 4489 1611 4508 1631
rect 1508 1450 1527 1470
rect 1585 1450 1604 1470
rect 1861 1471 1892 1498
rect 1088 1337 1114 1363
rect 713 1281 734 1301
rect 923 1281 948 1301
rect 1138 1284 1158 1304
rect 3780 1510 3800 1530
rect 3992 1515 4015 1535
rect 4204 1513 4225 1533
rect 3824 1451 3850 1477
rect 430 1183 449 1203
rect 507 1183 526 1203
rect 1365 1284 1394 1311
rect 1439 1287 1468 1314
rect 1712 1275 1744 1292
rect 2097 1279 2117 1299
rect 1653 1186 1674 1206
rect 3208 1272 3234 1294
rect 3473 1301 3492 1321
rect 3550 1301 3569 1321
rect 4202 1364 4223 1384
rect 1864 1157 1885 1198
rect 2026 1093 2052 1119
rect 1651 1037 1672 1057
rect 2076 1040 2096 1060
rect 203 974 228 993
rect 426 974 455 1001
rect 500 977 529 1004
rect 1158 969 1178 989
rect 3759 1271 3779 1291
rect 6213 2113 6233 2133
rect 8814 2415 8834 2435
rect 11188 3180 11208 3200
rect 13789 3482 13809 3502
rect 16243 4324 16263 4344
rect 18844 4626 18864 4646
rect 19493 4611 19522 4638
rect 19567 4614 19596 4641
rect 19794 4622 19819 4641
rect 17926 4555 17946 4575
rect 18350 4558 18371 4578
rect 17970 4496 17996 4522
rect 18137 4417 18158 4458
rect 15799 4231 15820 4251
rect 16453 4294 16472 4314
rect 16530 4294 16549 4314
rect 16788 4321 16814 4343
rect 18348 4409 18369 4429
rect 17905 4316 17925 4336
rect 18278 4323 18310 4340
rect 18554 4301 18583 4328
rect 18628 4304 18657 4331
rect 19496 4412 19515 4432
rect 19573 4412 19592 4432
rect 16172 4138 16198 4164
rect 15797 4082 15818 4102
rect 16007 4080 16030 4100
rect 16222 4085 16242 4105
rect 18864 4311 18884 4331
rect 19074 4314 19099 4334
rect 19288 4314 19309 4334
rect 18908 4252 18934 4278
rect 18130 4117 18161 4144
rect 18418 4145 18437 4165
rect 18495 4145 18514 4165
rect 15514 3984 15533 4004
rect 15591 3984 15610 4004
rect 16591 4047 16620 4074
rect 16665 4050 16694 4077
rect 16949 4041 16969 4058
rect 17323 4042 17343 4062
rect 16879 3949 16900 3969
rect 17252 3856 17278 3882
rect 15513 3780 15542 3807
rect 15587 3783 15616 3810
rect 15283 3667 15312 3696
rect 16245 3775 16265 3795
rect 16877 3800 16898 3820
rect 17085 3798 17112 3819
rect 17302 3803 17322 3823
rect 15801 3682 15822 3702
rect 19286 4165 19307 4185
rect 17786 4044 17806 4064
rect 18210 4047 18231 4067
rect 18843 4072 18863 4092
rect 19796 4171 19825 4200
rect 19492 4057 19521 4084
rect 19566 4060 19595 4087
rect 17830 3985 17856 4011
rect 17997 3905 18020 3943
rect 18208 3898 18229 3918
rect 17765 3805 17785 3825
rect 18139 3809 18159 3826
rect 18414 3790 18443 3817
rect 18488 3793 18517 3820
rect 19498 3863 19517 3883
rect 19575 3863 19594 3883
rect 16594 3702 16613 3722
rect 16671 3702 16690 3722
rect 16947 3723 16978 3750
rect 16174 3589 16200 3615
rect 15799 3533 15820 3553
rect 16009 3533 16034 3553
rect 16224 3536 16244 3556
rect 14438 3467 14467 3494
rect 14512 3470 14541 3497
rect 14739 3478 14764 3497
rect 12871 3411 12891 3431
rect 13081 3413 13101 3430
rect 13295 3414 13316 3434
rect 18866 3762 18886 3782
rect 19078 3767 19101 3787
rect 19290 3765 19311 3785
rect 18910 3703 18936 3729
rect 15516 3435 15535 3455
rect 15593 3435 15612 3455
rect 16451 3536 16480 3563
rect 16525 3539 16554 3566
rect 12915 3352 12941 3378
rect 16798 3527 16830 3544
rect 17183 3531 17203 3551
rect 16739 3438 16760 3458
rect 18294 3524 18320 3546
rect 18559 3553 18578 3573
rect 18636 3553 18655 3573
rect 19288 3616 19309 3636
rect 16950 3409 16971 3450
rect 10744 3087 10765 3107
rect 11398 3150 11417 3170
rect 11475 3150 11494 3170
rect 11733 3177 11759 3199
rect 13293 3265 13314 3285
rect 12850 3172 12870 3192
rect 17112 3345 17138 3371
rect 13499 3157 13528 3184
rect 13573 3160 13602 3187
rect 14441 3268 14460 3288
rect 14518 3268 14537 3288
rect 12740 3100 12788 3129
rect 11117 2994 11143 3020
rect 10742 2938 10763 2958
rect 10952 2936 10975 2956
rect 11167 2941 11187 2961
rect 16737 3289 16758 3309
rect 17162 3292 17182 3312
rect 15289 3226 15314 3245
rect 15512 3226 15541 3253
rect 15586 3229 15615 3256
rect 13809 3167 13829 3187
rect 14019 3170 14044 3190
rect 14233 3170 14254 3190
rect 13853 3108 13879 3134
rect 13393 2988 13412 3008
rect 13470 2988 13489 3008
rect 10459 2840 10478 2860
rect 10536 2840 10555 2860
rect 11505 2916 11534 2943
rect 11579 2919 11608 2946
rect 11846 2913 11867 2933
rect 12237 2911 12257 2929
rect 11793 2818 11814 2838
rect 12000 2794 12027 2826
rect 12166 2725 12192 2751
rect 10457 2636 10486 2663
rect 10531 2639 10560 2666
rect 11791 2669 11812 2689
rect 12216 2672 12236 2692
rect 10227 2523 10256 2552
rect 11189 2631 11209 2651
rect 10745 2538 10766 2558
rect 14231 3021 14252 3041
rect 13788 2928 13808 2948
rect 14741 3027 14770 3056
rect 12761 2887 12781 2907
rect 12969 2891 12998 2910
rect 13185 2890 13206 2910
rect 14437 2913 14466 2940
rect 14511 2916 14540 2943
rect 12805 2828 12831 2854
rect 16244 3221 16264 3241
rect 18845 3523 18865 3543
rect 19494 3508 19523 3535
rect 19568 3511 19597 3538
rect 19795 3519 19820 3538
rect 17927 3452 17947 3472
rect 18137 3454 18157 3471
rect 18351 3455 18372 3475
rect 17971 3393 17997 3419
rect 15800 3128 15821 3148
rect 16454 3191 16473 3211
rect 16531 3191 16550 3211
rect 16789 3218 16815 3240
rect 18349 3306 18370 3326
rect 17906 3213 17926 3233
rect 18555 3198 18584 3225
rect 18629 3201 18658 3228
rect 19497 3309 19516 3329
rect 19574 3309 19593 3329
rect 17796 3141 17844 3170
rect 16173 3035 16199 3061
rect 15798 2979 15819 2999
rect 16008 2977 16031 2997
rect 16223 2982 16243 3002
rect 18865 3208 18885 3228
rect 19075 3211 19100 3231
rect 19289 3211 19310 3231
rect 18909 3149 18935 3175
rect 18449 3029 18468 3049
rect 18526 3029 18545 3049
rect 15515 2881 15534 2901
rect 15592 2881 15611 2901
rect 13183 2741 13204 2761
rect 12740 2648 12760 2668
rect 13389 2633 13418 2660
rect 13463 2636 13492 2663
rect 16561 2957 16590 2984
rect 16635 2960 16664 2987
rect 16902 2954 16923 2974
rect 17293 2952 17313 2970
rect 16849 2859 16870 2879
rect 17056 2835 17083 2867
rect 14442 2719 14461 2739
rect 14519 2719 14538 2739
rect 11508 2571 11527 2591
rect 11585 2571 11604 2591
rect 12209 2590 12257 2619
rect 9463 2400 9492 2427
rect 9537 2403 9566 2430
rect 11118 2445 11144 2471
rect 9764 2411 9789 2430
rect 7896 2344 7916 2364
rect 8320 2347 8341 2367
rect 10743 2389 10764 2409
rect 10953 2389 10978 2409
rect 11168 2392 11188 2412
rect 7940 2285 7966 2311
rect 13810 2618 13830 2638
rect 14022 2623 14045 2643
rect 14234 2621 14255 2641
rect 13854 2559 13880 2585
rect 8107 2206 8128 2247
rect 5769 2020 5790 2040
rect 6423 2083 6442 2103
rect 6500 2083 6519 2103
rect 6758 2110 6784 2132
rect 8318 2198 8339 2218
rect 7875 2105 7895 2125
rect 8248 2112 8280 2129
rect 8524 2090 8553 2117
rect 8598 2093 8627 2120
rect 9466 2201 9485 2221
rect 9543 2201 9562 2221
rect 10460 2291 10479 2311
rect 10537 2291 10556 2311
rect 11395 2392 11424 2419
rect 11469 2395 11498 2422
rect 12127 2387 12147 2407
rect 11683 2294 11704 2314
rect 13238 2380 13264 2402
rect 13503 2409 13522 2429
rect 13580 2409 13599 2429
rect 14232 2472 14253 2492
rect 6142 1927 6168 1953
rect 5767 1871 5788 1891
rect 5977 1869 6000 1889
rect 6192 1874 6212 1894
rect 12056 2201 12082 2227
rect 8834 2100 8854 2120
rect 9044 2103 9069 2123
rect 9258 2103 9279 2123
rect 11681 2145 11702 2165
rect 11896 2149 11916 2166
rect 12106 2148 12126 2168
rect 10233 2082 10258 2101
rect 8878 2041 8904 2067
rect 10456 2082 10485 2109
rect 10530 2085 10559 2112
rect 8100 1906 8131 1933
rect 8388 1934 8407 1954
rect 8465 1934 8484 1954
rect 5484 1773 5503 1793
rect 5561 1773 5580 1793
rect 6561 1836 6590 1863
rect 6635 1839 6664 1866
rect 6919 1830 6939 1847
rect 7293 1831 7313 1851
rect 6849 1738 6870 1758
rect 7058 1713 7081 1751
rect 7222 1645 7248 1671
rect 5483 1569 5512 1596
rect 5557 1572 5586 1599
rect 5253 1456 5282 1485
rect 6215 1564 6235 1584
rect 6847 1589 6868 1609
rect 7272 1592 7292 1612
rect 5771 1471 5792 1491
rect 9256 1954 9277 1974
rect 7756 1833 7776 1853
rect 7966 1837 7993 1858
rect 8180 1836 8201 1856
rect 8813 1861 8833 1881
rect 9766 1960 9795 1989
rect 9462 1846 9491 1873
rect 9536 1849 9565 1876
rect 7800 1774 7826 1800
rect 8178 1687 8199 1707
rect 7735 1594 7755 1614
rect 8109 1598 8129 1615
rect 8384 1579 8413 1606
rect 8458 1582 8487 1609
rect 9468 1652 9487 1672
rect 9545 1652 9564 1672
rect 6564 1491 6583 1511
rect 6641 1491 6660 1511
rect 6917 1512 6948 1539
rect 6144 1378 6170 1404
rect 5769 1322 5790 1342
rect 5979 1322 6004 1342
rect 6194 1325 6214 1345
rect 4408 1256 4437 1283
rect 4482 1259 4511 1286
rect 4709 1267 4734 1286
rect 2841 1200 2861 1220
rect 3051 1202 3071 1219
rect 3265 1203 3286 1223
rect 8836 1551 8856 1571
rect 9048 1556 9071 1576
rect 9260 1554 9281 1574
rect 8880 1492 8906 1518
rect 5486 1224 5505 1244
rect 5563 1224 5582 1244
rect 6421 1325 6450 1352
rect 6495 1328 6524 1355
rect 2885 1141 2911 1167
rect 6768 1316 6800 1333
rect 7153 1320 7173 1340
rect 6709 1227 6730 1247
rect 8264 1313 8290 1335
rect 8529 1342 8548 1362
rect 8606 1342 8625 1362
rect 9258 1405 9279 1425
rect 6920 1198 6941 1239
rect 714 876 735 896
rect 1368 939 1387 959
rect 1445 939 1464 959
rect 1703 966 1729 988
rect 3263 1054 3284 1074
rect 2820 961 2840 981
rect 7082 1134 7108 1160
rect 3469 946 3498 973
rect 3543 949 3572 976
rect 4411 1057 4430 1077
rect 4488 1057 4507 1077
rect 1087 783 1113 809
rect 712 727 733 747
rect 922 725 945 745
rect 1137 730 1157 750
rect 6707 1078 6728 1098
rect 7132 1081 7152 1101
rect 5259 1015 5284 1034
rect 5482 1015 5511 1042
rect 5556 1018 5585 1045
rect 3779 956 3799 976
rect 3989 959 4014 979
rect 4203 959 4224 979
rect 3823 897 3849 923
rect 4201 810 4222 830
rect 3758 717 3778 737
rect 4711 816 4740 845
rect 4407 702 4436 729
rect 4481 705 4510 732
rect 429 629 448 649
rect 6214 1010 6234 1030
rect 8815 1312 8835 1332
rect 11188 2077 11208 2097
rect 13789 2379 13809 2399
rect 17222 2766 17248 2792
rect 15513 2677 15542 2704
rect 15587 2680 15616 2707
rect 16847 2710 16868 2730
rect 17272 2713 17292 2733
rect 15283 2564 15312 2593
rect 16245 2672 16265 2692
rect 15801 2579 15822 2599
rect 19287 3062 19308 3082
rect 18844 2969 18864 2989
rect 19797 3068 19826 3097
rect 17817 2928 17837 2948
rect 18025 2932 18054 2951
rect 18241 2931 18262 2951
rect 19493 2954 19522 2981
rect 19567 2957 19596 2984
rect 17861 2869 17887 2895
rect 18239 2782 18260 2802
rect 17796 2689 17816 2709
rect 18445 2674 18474 2701
rect 18519 2677 18548 2704
rect 19498 2760 19517 2780
rect 19575 2760 19594 2780
rect 16564 2612 16583 2632
rect 16641 2612 16660 2632
rect 17265 2631 17313 2660
rect 16174 2486 16200 2512
rect 15799 2430 15820 2450
rect 16009 2430 16034 2450
rect 16224 2433 16244 2453
rect 14438 2364 14467 2391
rect 14512 2367 14541 2394
rect 14739 2375 14764 2394
rect 12871 2308 12891 2328
rect 13295 2311 13316 2331
rect 18866 2659 18886 2679
rect 19078 2664 19101 2684
rect 19290 2662 19311 2682
rect 18910 2600 18936 2626
rect 15516 2332 15535 2352
rect 15593 2332 15612 2352
rect 16451 2433 16480 2460
rect 16525 2436 16554 2463
rect 12915 2249 12941 2275
rect 17183 2428 17203 2448
rect 16739 2335 16760 2355
rect 18294 2421 18320 2443
rect 18559 2450 18578 2470
rect 18636 2450 18655 2470
rect 19288 2513 19309 2533
rect 13082 2170 13103 2211
rect 10744 1984 10765 2004
rect 11398 2047 11417 2067
rect 11475 2047 11494 2067
rect 11733 2074 11759 2096
rect 13293 2162 13314 2182
rect 12850 2069 12870 2089
rect 13223 2076 13255 2093
rect 17112 2242 17138 2268
rect 13499 2054 13528 2081
rect 13573 2057 13602 2084
rect 14441 2165 14460 2185
rect 14518 2165 14537 2185
rect 11117 1891 11143 1917
rect 10742 1835 10763 1855
rect 10952 1833 10975 1853
rect 11167 1838 11187 1858
rect 16737 2186 16758 2206
rect 16952 2190 16972 2207
rect 17162 2189 17182 2209
rect 15289 2123 15314 2142
rect 15512 2123 15541 2150
rect 15586 2126 15615 2153
rect 13809 2064 13829 2084
rect 14019 2067 14044 2087
rect 14233 2067 14254 2087
rect 13853 2005 13879 2031
rect 13075 1870 13106 1897
rect 13363 1898 13382 1918
rect 13440 1898 13459 1918
rect 10459 1737 10478 1757
rect 10536 1737 10555 1757
rect 11536 1800 11565 1827
rect 11610 1803 11639 1830
rect 11894 1794 11914 1811
rect 12268 1795 12288 1815
rect 11824 1702 11845 1722
rect 12033 1677 12056 1715
rect 12197 1609 12223 1635
rect 10458 1533 10487 1560
rect 10532 1536 10561 1563
rect 10228 1420 10257 1449
rect 11190 1528 11210 1548
rect 11822 1553 11843 1573
rect 12247 1556 12267 1576
rect 10746 1435 10767 1455
rect 14231 1918 14252 1938
rect 12731 1797 12751 1817
rect 12941 1801 12968 1822
rect 13155 1800 13176 1820
rect 13788 1825 13808 1845
rect 14741 1924 14770 1953
rect 14437 1810 14466 1837
rect 14511 1813 14540 1840
rect 12775 1738 12801 1764
rect 13153 1651 13174 1671
rect 12710 1558 12730 1578
rect 13084 1562 13104 1579
rect 13359 1543 13388 1570
rect 13433 1546 13462 1573
rect 14443 1616 14462 1636
rect 14520 1616 14539 1636
rect 11539 1455 11558 1475
rect 11616 1455 11635 1475
rect 11892 1476 11923 1503
rect 9464 1297 9493 1324
rect 9538 1300 9567 1327
rect 11119 1342 11145 1368
rect 9765 1308 9790 1327
rect 7897 1241 7917 1261
rect 8107 1243 8127 1260
rect 8321 1244 8342 1264
rect 10744 1286 10765 1306
rect 10954 1286 10979 1306
rect 11169 1289 11189 1309
rect 7941 1182 7967 1208
rect 13811 1515 13831 1535
rect 14023 1520 14046 1540
rect 14235 1518 14256 1538
rect 13855 1456 13881 1482
rect 5770 917 5791 937
rect 6424 980 6443 1000
rect 6501 980 6520 1000
rect 6759 1007 6785 1029
rect 8319 1095 8340 1115
rect 7876 1002 7896 1022
rect 8525 987 8554 1014
rect 8599 990 8628 1017
rect 9467 1098 9486 1118
rect 9544 1098 9563 1118
rect 10461 1188 10480 1208
rect 10538 1188 10557 1208
rect 11396 1289 11425 1316
rect 11470 1292 11499 1319
rect 11743 1280 11775 1297
rect 12128 1284 12148 1304
rect 11684 1191 11705 1211
rect 13239 1277 13265 1299
rect 13504 1306 13523 1326
rect 13581 1306 13600 1326
rect 14233 1369 14254 1389
rect 11895 1162 11916 1203
rect 6143 824 6169 850
rect 5768 768 5789 788
rect 5978 766 6001 786
rect 6193 771 6213 791
rect 12057 1098 12083 1124
rect 8835 997 8855 1017
rect 9045 1000 9070 1020
rect 9259 1000 9280 1020
rect 11682 1042 11703 1062
rect 12107 1045 12127 1065
rect 10234 979 10259 998
rect 8879 938 8905 964
rect 10457 979 10486 1006
rect 10531 982 10560 1009
rect 9257 851 9278 871
rect 8814 758 8834 778
rect 9767 857 9796 886
rect 9463 743 9492 770
rect 9537 746 9566 773
rect 506 629 525 649
rect 757 546 786 567
rect 5485 670 5504 690
rect 5562 670 5581 690
rect 5813 587 5842 608
rect 9848 591 9877 612
rect 11189 974 11209 994
rect 13790 1276 13810 1296
rect 16244 2118 16264 2138
rect 18845 2420 18865 2440
rect 19494 2405 19523 2432
rect 19568 2408 19597 2435
rect 19795 2416 19820 2435
rect 17927 2349 17947 2369
rect 18351 2352 18372 2372
rect 17971 2290 17997 2316
rect 18138 2211 18159 2252
rect 15800 2025 15821 2045
rect 16454 2088 16473 2108
rect 16531 2088 16550 2108
rect 16789 2115 16815 2137
rect 18349 2203 18370 2223
rect 17906 2110 17926 2130
rect 18279 2117 18311 2134
rect 18555 2095 18584 2122
rect 18629 2098 18658 2125
rect 19497 2206 19516 2226
rect 19574 2206 19593 2226
rect 16173 1932 16199 1958
rect 15798 1876 15819 1896
rect 16008 1874 16031 1894
rect 16223 1879 16243 1899
rect 18865 2105 18885 2125
rect 19075 2108 19100 2128
rect 19289 2108 19310 2128
rect 18909 2046 18935 2072
rect 18131 1911 18162 1938
rect 18419 1939 18438 1959
rect 18496 1939 18515 1959
rect 15515 1778 15534 1798
rect 15592 1778 15611 1798
rect 16592 1841 16621 1868
rect 16666 1844 16695 1871
rect 16950 1835 16970 1852
rect 17324 1836 17344 1856
rect 16880 1743 16901 1763
rect 17089 1718 17112 1756
rect 17253 1650 17279 1676
rect 15514 1574 15543 1601
rect 15588 1577 15617 1604
rect 15284 1461 15313 1490
rect 16246 1569 16266 1589
rect 16878 1594 16899 1614
rect 17303 1597 17323 1617
rect 15802 1476 15823 1496
rect 19287 1959 19308 1979
rect 17787 1838 17807 1858
rect 17997 1842 18024 1863
rect 18211 1841 18232 1861
rect 18844 1866 18864 1886
rect 19797 1965 19826 1994
rect 19493 1851 19522 1878
rect 19567 1854 19596 1881
rect 17831 1779 17857 1805
rect 18209 1692 18230 1712
rect 17766 1599 17786 1619
rect 18140 1603 18160 1620
rect 18415 1584 18444 1611
rect 18489 1587 18518 1614
rect 19499 1657 19518 1677
rect 19576 1657 19595 1677
rect 16595 1496 16614 1516
rect 16672 1496 16691 1516
rect 16948 1517 16979 1544
rect 16175 1383 16201 1409
rect 15800 1327 15821 1347
rect 16010 1327 16035 1347
rect 16225 1330 16245 1350
rect 14439 1261 14468 1288
rect 14513 1264 14542 1291
rect 14740 1272 14765 1291
rect 12872 1205 12892 1225
rect 13082 1207 13102 1224
rect 13296 1208 13317 1228
rect 18867 1556 18887 1576
rect 19079 1561 19102 1581
rect 19291 1559 19312 1579
rect 18911 1497 18937 1523
rect 15517 1229 15536 1249
rect 15594 1229 15613 1249
rect 16452 1330 16481 1357
rect 16526 1333 16555 1360
rect 12916 1146 12942 1172
rect 16799 1321 16831 1338
rect 17184 1325 17204 1345
rect 16740 1232 16761 1252
rect 18295 1318 18321 1340
rect 18560 1347 18579 1367
rect 18637 1347 18656 1367
rect 19289 1410 19310 1430
rect 16951 1203 16972 1244
rect 10745 881 10766 901
rect 11399 944 11418 964
rect 11476 944 11495 964
rect 11734 971 11760 993
rect 13294 1059 13315 1079
rect 12851 966 12871 986
rect 17113 1139 17139 1165
rect 13500 951 13529 978
rect 13574 954 13603 981
rect 14442 1062 14461 1082
rect 14519 1062 14538 1082
rect 11118 788 11144 814
rect 10743 732 10764 752
rect 10953 730 10976 750
rect 11168 735 11188 755
rect 16738 1083 16759 1103
rect 17163 1086 17183 1106
rect 15290 1020 15315 1039
rect 15513 1020 15542 1047
rect 15587 1023 15616 1050
rect 13810 961 13830 981
rect 14020 964 14045 984
rect 14234 964 14255 984
rect 13854 902 13880 928
rect 14232 815 14253 835
rect 13789 722 13809 742
rect 14742 821 14771 850
rect 14438 707 14467 734
rect 14512 710 14541 737
rect 10460 634 10479 654
rect 16245 1015 16265 1035
rect 18846 1317 18866 1337
rect 19495 1302 19524 1329
rect 19569 1305 19598 1332
rect 19796 1313 19821 1332
rect 17928 1246 17948 1266
rect 18138 1248 18158 1265
rect 18352 1249 18373 1269
rect 17972 1187 17998 1213
rect 15801 922 15822 942
rect 16455 985 16474 1005
rect 16532 985 16551 1005
rect 16790 1012 16816 1034
rect 18350 1100 18371 1120
rect 17907 1007 17927 1027
rect 18556 992 18585 1019
rect 18630 995 18659 1022
rect 19498 1103 19517 1123
rect 19575 1103 19594 1123
rect 16174 829 16200 855
rect 15799 773 15820 793
rect 16009 771 16032 791
rect 16224 776 16244 796
rect 18866 1002 18886 1022
rect 19076 1005 19101 1025
rect 19290 1005 19311 1025
rect 18910 943 18936 969
rect 19288 856 19309 876
rect 18845 763 18865 783
rect 19798 862 19827 891
rect 19494 748 19523 775
rect 19568 751 19597 778
rect 10537 634 10556 654
rect 4792 550 4821 571
rect 10788 551 10817 572
rect 15516 675 15535 695
rect 15593 675 15612 695
rect 15844 592 15873 613
rect 19879 596 19908 617
rect 14823 555 14852 576
rect 1673 415 1702 442
rect 1747 418 1776 445
rect 6729 456 6758 483
rect 6803 459 6832 486
rect 2405 410 2425 430
rect 1961 317 1982 337
rect 4623 395 4652 422
rect 4697 398 4726 425
rect 2334 224 2360 250
rect 1959 168 1980 188
rect 2165 167 2199 187
rect 2384 171 2404 191
rect 5355 390 5375 410
rect 4911 297 4932 317
rect 7461 451 7481 471
rect 7017 358 7038 378
rect 11704 420 11733 447
rect 11778 423 11807 450
rect 16760 461 16789 488
rect 16834 464 16863 491
rect 5284 204 5310 230
rect 4909 148 4930 168
rect 5109 147 5150 167
rect 5334 151 5354 171
rect 2486 109 2513 130
rect 1676 70 1695 90
rect 1753 70 1772 90
rect 7390 265 7416 291
rect 7015 209 7036 229
rect 7221 208 7255 228
rect 7440 212 7460 232
rect 9557 279 9586 306
rect 9631 282 9660 309
rect 7542 150 7569 171
rect 5422 85 5481 111
rect 6732 111 6751 131
rect 6809 111 6828 131
rect 10289 274 10309 294
rect 9845 181 9866 201
rect 12436 415 12456 435
rect 11992 322 12013 342
rect 14654 400 14683 427
rect 14728 403 14757 430
rect 12365 229 12391 255
rect 10218 88 10244 114
rect 4626 50 4645 70
rect 4703 50 4722 70
rect 9843 32 9864 52
rect 10050 28 10083 52
rect 10268 35 10288 55
rect 11990 173 12011 193
rect 12196 172 12230 192
rect 12415 176 12435 196
rect 15386 395 15406 415
rect 14942 302 14963 322
rect 17492 456 17512 476
rect 17048 363 17069 383
rect 15315 209 15341 235
rect 14940 153 14961 173
rect 15137 149 15178 173
rect 15365 156 15385 176
rect 12517 114 12544 135
rect 11707 75 11726 95
rect 11784 75 11803 95
rect 17421 270 17447 296
rect 17046 214 17067 234
rect 17252 213 17286 233
rect 17471 217 17491 237
rect 17573 155 17600 176
rect 15453 90 15512 116
rect 16763 116 16782 136
rect 16840 116 16859 136
rect 14657 55 14676 75
rect 14734 55 14753 75
rect 9560 -66 9579 -46
rect 9637 -66 9656 -46
rect 10282 -42 10323 -12
<< metal1 >>
rect 18806 9416 19108 9418
rect 8775 9411 9077 9413
rect 6206 9388 6241 9390
rect 5242 9385 6241 9388
rect 3719 9370 4021 9372
rect 1150 9347 1185 9349
rect 186 9344 1185 9347
rect 185 9320 1185 9344
rect 185 9165 233 9320
rect 419 9279 529 9293
rect 419 9276 497 9279
rect 419 9249 423 9276
rect 452 9252 497 9276
rect 526 9252 529 9279
rect 1150 9269 1185 9320
rect 452 9249 529 9252
rect 419 9234 529 9249
rect 1148 9264 1185 9269
rect 1148 9244 1155 9264
rect 1175 9244 1185 9264
rect 1148 9237 1185 9244
rect 3658 9341 4021 9370
rect 3658 9339 3719 9341
rect 1148 9236 1183 9237
rect 185 9136 193 9165
rect 222 9136 233 9165
rect 185 9131 233 9136
rect 704 9171 736 9178
rect 704 9151 711 9171
rect 732 9151 736 9171
rect 704 9086 736 9151
rect 1074 9086 1114 9087
rect 704 9084 1116 9086
rect 704 9058 1084 9084
rect 1110 9058 1116 9084
rect 704 9050 1116 9058
rect 704 9022 736 9050
rect 1149 9030 1183 9236
rect 3200 9119 3237 9121
rect 3658 9119 3691 9339
rect 3979 9260 4021 9341
rect 4401 9352 4512 9369
rect 4401 9332 4408 9352
rect 4427 9332 4485 9352
rect 4504 9332 4512 9352
rect 4401 9310 4512 9332
rect 5241 9361 6241 9385
rect 3768 9258 3803 9259
rect 2087 9103 2121 9104
rect 1218 9068 2122 9103
rect 3200 9090 3691 9119
rect 704 9002 709 9022
rect 730 9002 736 9022
rect 704 8995 736 9002
rect 911 9022 950 9028
rect 911 9002 919 9022
rect 944 9002 950 9022
rect 911 8995 950 9002
rect 1127 9025 1183 9030
rect 1127 9005 1134 9025
rect 1154 9005 1183 9025
rect 1127 8998 1183 9005
rect 1127 8997 1162 8998
rect 919 8949 950 8995
rect 418 8924 529 8946
rect 418 8904 426 8924
rect 445 8904 503 8924
rect 522 8904 529 8924
rect 918 8932 950 8949
rect 1219 8932 1256 9068
rect 1357 9035 1467 9049
rect 1357 9032 1435 9035
rect 1357 9005 1361 9032
rect 1390 9008 1435 9032
rect 1464 9008 1467 9035
rect 2087 9025 2121 9068
rect 1390 9005 1467 9008
rect 1357 8990 1467 9005
rect 2086 9020 2121 9025
rect 3200 9024 3237 9090
rect 3658 9089 3691 9090
rect 3747 9251 3803 9258
rect 3747 9231 3776 9251
rect 3796 9231 3803 9251
rect 3747 9226 3803 9231
rect 3977 9256 4021 9260
rect 3977 9236 3988 9256
rect 4011 9236 4021 9256
rect 3977 9229 4021 9236
rect 4194 9254 4226 9261
rect 4194 9234 4200 9254
rect 4221 9234 4226 9254
rect 3977 9227 4020 9229
rect 2086 9000 2093 9020
rect 2113 9000 2121 9020
rect 2086 8992 2121 9000
rect 918 8919 1256 8932
rect 418 8887 529 8904
rect 919 8900 1256 8919
rect 1198 8899 1256 8900
rect 1642 8927 1674 8934
rect 1642 8907 1649 8927
rect 1670 8907 1674 8927
rect 1642 8842 1674 8907
rect 2012 8842 2052 8843
rect 1642 8840 2054 8842
rect 1642 8814 2022 8840
rect 2048 8814 2054 8840
rect 1642 8806 2054 8814
rect 188 8767 1184 8793
rect 1642 8778 1674 8806
rect 190 8714 232 8767
rect 190 8695 199 8714
rect 224 8695 232 8714
rect 190 8685 232 8695
rect 418 8725 528 8739
rect 418 8722 496 8725
rect 418 8695 422 8722
rect 451 8698 496 8722
rect 525 8698 528 8725
rect 1148 8715 1182 8767
rect 1642 8758 1647 8778
rect 1668 8758 1674 8778
rect 1642 8751 1674 8758
rect 1852 8779 1890 8789
rect 2087 8786 2121 8992
rect 3195 9015 3237 9024
rect 3195 8993 3204 9015
rect 3230 8993 3237 9015
rect 3462 9042 3573 9059
rect 3462 9022 3469 9042
rect 3488 9022 3546 9042
rect 3565 9022 3573 9042
rect 3462 9000 3573 9022
rect 3747 9020 3781 9226
rect 4194 9206 4226 9234
rect 3814 9198 4226 9206
rect 3814 9172 3820 9198
rect 3846 9172 4226 9198
rect 5241 9206 5289 9361
rect 5475 9320 5585 9334
rect 5475 9317 5553 9320
rect 5475 9290 5479 9317
rect 5508 9293 5553 9317
rect 5582 9293 5585 9320
rect 6206 9310 6241 9361
rect 5508 9290 5585 9293
rect 5475 9275 5585 9290
rect 6204 9305 6241 9310
rect 6204 9285 6211 9305
rect 6231 9285 6241 9305
rect 6204 9278 6241 9285
rect 8714 9382 9077 9411
rect 8714 9380 8775 9382
rect 6204 9277 6239 9278
rect 5241 9177 5249 9206
rect 5278 9177 5289 9206
rect 5241 9172 5289 9177
rect 5760 9212 5792 9219
rect 5760 9192 5767 9212
rect 5788 9192 5792 9212
rect 3814 9170 4226 9172
rect 3816 9169 3856 9170
rect 4194 9105 4226 9170
rect 4194 9085 4198 9105
rect 4219 9085 4226 9105
rect 4194 9078 4226 9085
rect 5760 9127 5792 9192
rect 6130 9127 6170 9128
rect 5760 9125 6172 9127
rect 5760 9099 6140 9125
rect 6166 9099 6172 9125
rect 5760 9091 6172 9099
rect 5760 9063 5792 9091
rect 6205 9071 6239 9277
rect 8256 9160 8293 9162
rect 8714 9160 8747 9380
rect 9035 9301 9077 9382
rect 9457 9393 9568 9408
rect 16237 9393 16272 9395
rect 9457 9373 9464 9393
rect 9483 9373 9541 9393
rect 9560 9373 9568 9393
rect 15273 9390 16272 9393
rect 13750 9375 14052 9377
rect 9457 9351 9568 9373
rect 11181 9352 11216 9354
rect 10217 9349 11216 9352
rect 10216 9325 11216 9349
rect 8824 9299 8859 9300
rect 7143 9144 7177 9145
rect 6274 9109 7178 9144
rect 8256 9131 8747 9160
rect 5760 9043 5765 9063
rect 5786 9043 5792 9063
rect 5760 9036 5792 9043
rect 5967 9063 6006 9069
rect 5967 9043 5975 9063
rect 6000 9043 6006 9063
rect 5967 9036 6006 9043
rect 6183 9066 6239 9071
rect 6183 9046 6190 9066
rect 6210 9046 6239 9066
rect 6183 9039 6239 9046
rect 6183 9038 6218 9039
rect 3747 9012 3782 9020
rect 3195 8983 3237 8993
rect 3747 8992 3755 9012
rect 3775 8992 3782 9012
rect 3747 8987 3782 8992
rect 4401 9007 4511 9022
rect 4401 9004 4478 9007
rect 3195 8982 3236 8983
rect 2829 8948 2864 8949
rect 1852 8762 1862 8779
rect 1882 8762 1890 8779
rect 1693 8719 1734 8720
rect 451 8695 528 8698
rect 418 8680 528 8695
rect 1147 8710 1182 8715
rect 1147 8690 1154 8710
rect 1174 8690 1182 8710
rect 1692 8709 1734 8719
rect 1147 8682 1182 8690
rect 703 8617 735 8624
rect 703 8597 710 8617
rect 731 8597 735 8617
rect 703 8532 735 8597
rect 1073 8532 1113 8533
rect 703 8530 1115 8532
rect 703 8504 1083 8530
rect 1109 8504 1115 8530
rect 703 8496 1115 8504
rect 703 8468 735 8496
rect 1148 8476 1182 8682
rect 1356 8680 1467 8702
rect 1356 8660 1364 8680
rect 1383 8660 1441 8680
rect 1460 8660 1467 8680
rect 1356 8643 1467 8660
rect 1692 8687 1699 8709
rect 1725 8687 1734 8709
rect 1692 8678 1734 8687
rect 909 8473 952 8475
rect 703 8448 708 8468
rect 729 8448 735 8468
rect 703 8441 735 8448
rect 908 8466 952 8473
rect 908 8446 918 8466
rect 941 8446 952 8466
rect 908 8442 952 8446
rect 1126 8471 1182 8476
rect 1126 8451 1133 8471
rect 1153 8451 1182 8471
rect 1126 8444 1182 8451
rect 1238 8612 1271 8613
rect 1692 8612 1729 8678
rect 1238 8583 1729 8612
rect 1126 8443 1161 8444
rect 417 8370 528 8392
rect 417 8350 425 8370
rect 444 8350 502 8370
rect 521 8350 528 8370
rect 417 8333 528 8350
rect 908 8361 950 8442
rect 1238 8363 1271 8583
rect 1692 8581 1729 8583
rect 1498 8443 1608 8457
rect 1498 8440 1576 8443
rect 1498 8413 1502 8440
rect 1531 8416 1576 8440
rect 1605 8416 1608 8443
rect 1531 8413 1608 8416
rect 1498 8398 1608 8413
rect 1852 8424 1890 8762
rect 2065 8781 2121 8786
rect 2065 8761 2072 8781
rect 2092 8761 2121 8781
rect 2065 8754 2121 8761
rect 2808 8941 2864 8948
rect 2808 8921 2837 8941
rect 2857 8921 2864 8941
rect 2808 8916 2864 8921
rect 3255 8944 3287 8951
rect 3255 8924 3261 8944
rect 3282 8924 3287 8944
rect 3747 8935 3781 8987
rect 4401 8977 4404 9004
rect 4433 8980 4478 9004
rect 4507 8980 4511 9007
rect 4433 8977 4511 8980
rect 4401 8963 4511 8977
rect 4697 9007 4739 9017
rect 4697 8988 4705 9007
rect 4730 8988 4739 9007
rect 5975 8990 6006 9036
rect 4697 8935 4739 8988
rect 5474 8965 5585 8987
rect 5474 8945 5482 8965
rect 5501 8945 5559 8965
rect 5578 8945 5585 8965
rect 5974 8973 6006 8990
rect 6275 8973 6312 9109
rect 6413 9076 6523 9090
rect 6413 9073 6491 9076
rect 6413 9046 6417 9073
rect 6446 9049 6491 9073
rect 6520 9049 6523 9076
rect 7143 9066 7177 9109
rect 6446 9046 6523 9049
rect 6413 9031 6523 9046
rect 7142 9061 7177 9066
rect 8256 9065 8293 9131
rect 8714 9130 8747 9131
rect 8803 9292 8859 9299
rect 8803 9272 8832 9292
rect 8852 9272 8859 9292
rect 8803 9267 8859 9272
rect 9033 9297 9077 9301
rect 9033 9277 9044 9297
rect 9067 9277 9077 9297
rect 9033 9270 9077 9277
rect 9250 9295 9282 9302
rect 9250 9275 9256 9295
rect 9277 9275 9282 9295
rect 9033 9268 9076 9270
rect 7142 9041 7149 9061
rect 7169 9041 7177 9061
rect 7142 9033 7177 9041
rect 5974 8960 6312 8973
rect 2065 8753 2100 8754
rect 2808 8710 2842 8916
rect 3255 8896 3287 8924
rect 3745 8909 4741 8935
rect 5474 8928 5585 8945
rect 5975 8941 6312 8960
rect 6254 8940 6312 8941
rect 6698 8968 6730 8975
rect 6698 8948 6705 8968
rect 6726 8948 6730 8968
rect 2875 8888 3287 8896
rect 2875 8862 2881 8888
rect 2907 8862 3287 8888
rect 2875 8860 3287 8862
rect 2877 8859 2917 8860
rect 3037 8824 3076 8839
rect 3037 8783 3048 8824
rect 3069 8783 3076 8824
rect 2807 8702 2843 8710
rect 2807 8682 2816 8702
rect 2836 8682 2843 8702
rect 2807 8681 2843 8682
rect 2807 8670 2841 8681
rect 3037 8510 3076 8783
rect 3255 8795 3287 8860
rect 6698 8883 6730 8948
rect 7068 8883 7108 8884
rect 6698 8881 7110 8883
rect 6698 8855 7078 8881
rect 7104 8855 7110 8881
rect 6698 8847 7110 8855
rect 3255 8775 3259 8795
rect 3280 8775 3287 8795
rect 3255 8768 3287 8775
rect 3673 8802 3731 8803
rect 3673 8783 4010 8802
rect 4400 8798 4511 8815
rect 5244 8808 6240 8834
rect 6698 8819 6730 8847
rect 3673 8770 4011 8783
rect 3177 8706 3230 8709
rect 3177 8689 3189 8706
rect 3221 8689 3230 8706
rect 3177 8681 3230 8689
rect 3176 8634 3230 8681
rect 3462 8697 3572 8712
rect 3462 8694 3539 8697
rect 3462 8667 3465 8694
rect 3494 8670 3539 8694
rect 3568 8670 3572 8697
rect 3494 8667 3572 8670
rect 3462 8653 3572 8667
rect 3673 8634 3710 8770
rect 3979 8753 4011 8770
rect 4400 8778 4407 8798
rect 4426 8778 4484 8798
rect 4503 8778 4511 8798
rect 4400 8756 4511 8778
rect 5246 8755 5288 8808
rect 3979 8707 4010 8753
rect 5246 8736 5255 8755
rect 5280 8736 5288 8755
rect 5246 8726 5288 8736
rect 5474 8766 5584 8780
rect 5474 8763 5552 8766
rect 5474 8736 5478 8763
rect 5507 8739 5552 8763
rect 5581 8739 5584 8766
rect 6204 8756 6238 8808
rect 6698 8799 6703 8819
rect 6724 8799 6730 8819
rect 6698 8792 6730 8799
rect 6908 8820 6946 8830
rect 7143 8827 7177 9033
rect 8251 9056 8293 9065
rect 8251 9034 8260 9056
rect 8286 9034 8293 9056
rect 8518 9083 8629 9100
rect 8518 9063 8525 9083
rect 8544 9063 8602 9083
rect 8621 9063 8629 9083
rect 8518 9041 8629 9063
rect 8803 9061 8837 9267
rect 9250 9247 9282 9275
rect 8870 9239 9282 9247
rect 8870 9213 8876 9239
rect 8902 9213 9282 9239
rect 8870 9211 9282 9213
rect 8872 9210 8912 9211
rect 9250 9146 9282 9211
rect 9250 9126 9254 9146
rect 9275 9126 9282 9146
rect 10216 9170 10264 9325
rect 10450 9284 10560 9298
rect 10450 9281 10528 9284
rect 10450 9254 10454 9281
rect 10483 9257 10528 9281
rect 10557 9257 10560 9284
rect 11181 9274 11216 9325
rect 10483 9254 10560 9257
rect 10450 9239 10560 9254
rect 11179 9269 11216 9274
rect 11179 9249 11186 9269
rect 11206 9249 11216 9269
rect 11179 9242 11216 9249
rect 13689 9346 14052 9375
rect 13689 9344 13750 9346
rect 11179 9241 11214 9242
rect 10216 9141 10224 9170
rect 10253 9141 10264 9170
rect 10216 9136 10264 9141
rect 10735 9176 10767 9183
rect 10735 9156 10742 9176
rect 10763 9156 10767 9176
rect 9250 9119 9282 9126
rect 10735 9091 10767 9156
rect 11105 9091 11145 9092
rect 10735 9089 11147 9091
rect 10735 9063 11115 9089
rect 11141 9063 11147 9089
rect 8803 9053 8838 9061
rect 8251 9024 8293 9034
rect 8803 9033 8811 9053
rect 8831 9033 8838 9053
rect 8803 9028 8838 9033
rect 9457 9048 9567 9063
rect 9457 9045 9534 9048
rect 8251 9023 8292 9024
rect 7885 8989 7920 8990
rect 6908 8803 6918 8820
rect 6938 8803 6946 8820
rect 6749 8760 6790 8761
rect 5507 8736 5584 8739
rect 5474 8721 5584 8736
rect 6203 8751 6238 8756
rect 6203 8731 6210 8751
rect 6230 8731 6238 8751
rect 6748 8750 6790 8760
rect 6203 8723 6238 8731
rect 3767 8704 3802 8705
rect 3746 8697 3802 8704
rect 3746 8677 3775 8697
rect 3795 8677 3802 8697
rect 3746 8672 3802 8677
rect 3979 8700 4018 8707
rect 3979 8680 3985 8700
rect 4010 8680 4018 8700
rect 3979 8674 4018 8680
rect 4193 8700 4225 8707
rect 4193 8680 4199 8700
rect 4220 8680 4225 8700
rect 3176 8599 3711 8634
rect 3176 8595 3229 8599
rect 3037 8483 3041 8510
rect 3072 8483 3076 8510
rect 3322 8531 3433 8548
rect 3322 8511 3329 8531
rect 3348 8511 3406 8531
rect 3425 8511 3433 8531
rect 3322 8489 3433 8511
rect 3037 8476 3076 8483
rect 3746 8466 3780 8672
rect 4193 8652 4225 8680
rect 3813 8644 4225 8652
rect 3813 8618 3819 8644
rect 3845 8618 4225 8644
rect 3813 8616 4225 8618
rect 3815 8615 3855 8616
rect 4193 8551 4225 8616
rect 5759 8658 5791 8665
rect 5759 8638 5766 8658
rect 5787 8638 5791 8658
rect 5759 8573 5791 8638
rect 6129 8573 6169 8574
rect 5759 8571 6171 8573
rect 4193 8531 4197 8551
rect 4218 8531 4225 8551
rect 4193 8524 4225 8531
rect 4696 8566 4744 8571
rect 4696 8537 4707 8566
rect 4736 8537 4744 8566
rect 3746 8465 3781 8466
rect 3744 8458 3781 8465
rect 2689 8437 2724 8438
rect 2230 8433 2262 8434
rect 1852 8407 1860 8424
rect 1880 8407 1890 8424
rect 1852 8401 1890 8407
rect 2227 8428 2262 8433
rect 2227 8408 2234 8428
rect 2254 8408 2262 8428
rect 2227 8400 2262 8408
rect 1210 8361 1271 8363
rect 908 8332 1271 8361
rect 1783 8335 1815 8342
rect 908 8330 1210 8332
rect 1783 8315 1790 8335
rect 1811 8315 1815 8335
rect 1783 8250 1815 8315
rect 2153 8250 2193 8251
rect 1783 8248 2195 8250
rect 1151 8244 1186 8246
rect 187 8241 1186 8244
rect 186 8217 1186 8241
rect 186 8062 234 8217
rect 420 8176 530 8190
rect 420 8173 498 8176
rect 420 8146 424 8173
rect 453 8149 498 8173
rect 527 8149 530 8176
rect 1151 8166 1186 8217
rect 453 8146 530 8149
rect 420 8131 530 8146
rect 1149 8161 1186 8166
rect 1149 8141 1156 8161
rect 1176 8141 1186 8161
rect 1783 8222 2163 8248
rect 2189 8222 2195 8248
rect 1783 8214 2195 8222
rect 1783 8186 1815 8214
rect 1783 8166 1788 8186
rect 1809 8166 1815 8186
rect 1783 8159 1815 8166
rect 1989 8185 2031 8196
rect 2228 8194 2262 8400
rect 2666 8430 2724 8437
rect 2666 8410 2697 8430
rect 2717 8410 2724 8430
rect 2666 8405 2724 8410
rect 3115 8433 3147 8440
rect 3115 8413 3121 8433
rect 3142 8413 3147 8433
rect 2666 8257 2702 8405
rect 3115 8385 3147 8413
rect 2735 8377 3147 8385
rect 2735 8351 2741 8377
rect 2767 8351 3147 8377
rect 3744 8438 3754 8458
rect 3774 8438 3781 8458
rect 3744 8433 3781 8438
rect 4400 8453 4510 8468
rect 4400 8450 4477 8453
rect 3744 8382 3779 8433
rect 4400 8423 4403 8450
rect 4432 8426 4477 8450
rect 4506 8426 4510 8453
rect 4432 8423 4510 8426
rect 4400 8409 4510 8423
rect 4696 8382 4744 8537
rect 5759 8545 6139 8571
rect 6165 8545 6171 8571
rect 5759 8537 6171 8545
rect 5759 8509 5791 8537
rect 6204 8517 6238 8723
rect 6412 8721 6523 8743
rect 6412 8701 6420 8721
rect 6439 8701 6497 8721
rect 6516 8701 6523 8721
rect 6412 8684 6523 8701
rect 6748 8728 6755 8750
rect 6781 8728 6790 8750
rect 6748 8719 6790 8728
rect 5965 8514 6008 8516
rect 5759 8489 5764 8509
rect 5785 8489 5791 8509
rect 5759 8482 5791 8489
rect 5964 8507 6008 8514
rect 5964 8487 5974 8507
rect 5997 8487 6008 8507
rect 5964 8483 6008 8487
rect 6182 8512 6238 8517
rect 6182 8492 6189 8512
rect 6209 8492 6238 8512
rect 6182 8485 6238 8492
rect 6294 8653 6327 8654
rect 6748 8653 6785 8719
rect 6294 8624 6785 8653
rect 6182 8484 6217 8485
rect 3744 8358 4744 8382
rect 5473 8411 5584 8433
rect 5473 8391 5481 8411
rect 5500 8391 5558 8411
rect 5577 8391 5584 8411
rect 5473 8374 5584 8391
rect 5964 8402 6006 8483
rect 6294 8404 6327 8624
rect 6748 8622 6785 8624
rect 6554 8484 6664 8498
rect 6554 8481 6632 8484
rect 6554 8454 6558 8481
rect 6587 8457 6632 8481
rect 6661 8457 6664 8484
rect 6587 8454 6664 8457
rect 6554 8439 6664 8454
rect 6908 8465 6946 8803
rect 7121 8822 7177 8827
rect 7121 8802 7128 8822
rect 7148 8802 7177 8822
rect 7121 8795 7177 8802
rect 7864 8982 7920 8989
rect 7864 8962 7893 8982
rect 7913 8962 7920 8982
rect 7864 8957 7920 8962
rect 8311 8985 8343 8992
rect 8311 8965 8317 8985
rect 8338 8965 8343 8985
rect 8803 8976 8837 9028
rect 9457 9018 9460 9045
rect 9489 9021 9534 9045
rect 9563 9021 9567 9048
rect 9489 9018 9567 9021
rect 9457 9004 9567 9018
rect 9753 9048 9795 9058
rect 9753 9029 9761 9048
rect 9786 9029 9795 9048
rect 9753 8976 9795 9029
rect 10735 9055 11147 9063
rect 10735 9027 10767 9055
rect 11180 9035 11214 9241
rect 13231 9124 13268 9126
rect 13689 9124 13722 9344
rect 14010 9265 14052 9346
rect 14432 9357 14543 9374
rect 14432 9337 14439 9357
rect 14458 9337 14516 9357
rect 14535 9337 14543 9357
rect 14432 9315 14543 9337
rect 15272 9366 16272 9390
rect 13799 9263 13834 9264
rect 12118 9108 12152 9109
rect 11249 9073 12153 9108
rect 13231 9095 13722 9124
rect 10735 9007 10740 9027
rect 10761 9007 10767 9027
rect 10735 9000 10767 9007
rect 10942 9027 10981 9033
rect 10942 9007 10950 9027
rect 10975 9007 10981 9027
rect 10942 9000 10981 9007
rect 11158 9030 11214 9035
rect 11158 9010 11165 9030
rect 11185 9010 11214 9030
rect 11158 9003 11214 9010
rect 11158 9002 11193 9003
rect 7121 8794 7156 8795
rect 7864 8751 7898 8957
rect 8311 8937 8343 8965
rect 8801 8950 9797 8976
rect 10950 8954 10981 9000
rect 7931 8929 8343 8937
rect 7931 8903 7937 8929
rect 7963 8903 8343 8929
rect 7931 8901 8343 8903
rect 7933 8900 7973 8901
rect 8093 8865 8132 8880
rect 8093 8824 8104 8865
rect 8125 8824 8132 8865
rect 7863 8743 7899 8751
rect 7863 8723 7872 8743
rect 7892 8723 7899 8743
rect 7863 8722 7899 8723
rect 7863 8711 7897 8722
rect 8093 8551 8132 8824
rect 8311 8836 8343 8901
rect 10449 8929 10560 8951
rect 10449 8909 10457 8929
rect 10476 8909 10534 8929
rect 10553 8909 10560 8929
rect 10949 8937 10981 8954
rect 11250 8937 11287 9073
rect 11388 9040 11498 9054
rect 11388 9037 11466 9040
rect 11388 9010 11392 9037
rect 11421 9013 11466 9037
rect 11495 9013 11498 9040
rect 12118 9030 12152 9073
rect 11421 9010 11498 9013
rect 11388 8995 11498 9010
rect 12117 9025 12152 9030
rect 13231 9029 13268 9095
rect 13689 9094 13722 9095
rect 13778 9256 13834 9263
rect 13778 9236 13807 9256
rect 13827 9236 13834 9256
rect 13778 9231 13834 9236
rect 14008 9261 14052 9265
rect 14008 9241 14019 9261
rect 14042 9241 14052 9261
rect 14008 9234 14052 9241
rect 14225 9259 14257 9266
rect 14225 9239 14231 9259
rect 14252 9239 14257 9259
rect 14008 9232 14051 9234
rect 12117 9005 12124 9025
rect 12144 9005 12152 9025
rect 12117 8997 12152 9005
rect 10949 8924 11287 8937
rect 10449 8892 10560 8909
rect 10950 8905 11287 8924
rect 11229 8904 11287 8905
rect 11673 8932 11705 8939
rect 11673 8912 11680 8932
rect 11701 8912 11705 8932
rect 8311 8816 8315 8836
rect 8336 8816 8343 8836
rect 8311 8809 8343 8816
rect 8729 8843 8787 8844
rect 8729 8824 9066 8843
rect 9456 8839 9567 8856
rect 8729 8811 9067 8824
rect 8233 8747 8286 8750
rect 8233 8730 8245 8747
rect 8277 8730 8286 8747
rect 8233 8722 8286 8730
rect 8232 8675 8286 8722
rect 8518 8738 8628 8753
rect 8518 8735 8595 8738
rect 8518 8708 8521 8735
rect 8550 8711 8595 8735
rect 8624 8711 8628 8738
rect 8550 8708 8628 8711
rect 8518 8694 8628 8708
rect 8729 8675 8766 8811
rect 9035 8794 9067 8811
rect 9456 8819 9463 8839
rect 9482 8819 9540 8839
rect 9559 8819 9567 8839
rect 9456 8797 9567 8819
rect 11673 8847 11705 8912
rect 12043 8847 12083 8848
rect 11673 8845 12085 8847
rect 11673 8819 12053 8845
rect 12079 8819 12085 8845
rect 11673 8811 12085 8819
rect 9035 8748 9066 8794
rect 10219 8772 11215 8798
rect 11673 8783 11705 8811
rect 8823 8745 8858 8746
rect 8802 8738 8858 8745
rect 8802 8718 8831 8738
rect 8851 8718 8858 8738
rect 8802 8713 8858 8718
rect 9035 8741 9074 8748
rect 9035 8721 9041 8741
rect 9066 8721 9074 8741
rect 9035 8715 9074 8721
rect 9249 8741 9281 8748
rect 9249 8721 9255 8741
rect 9276 8721 9281 8741
rect 8232 8640 8767 8675
rect 8232 8636 8285 8640
rect 8093 8524 8097 8551
rect 8128 8524 8132 8551
rect 8378 8572 8489 8589
rect 8378 8552 8385 8572
rect 8404 8552 8462 8572
rect 8481 8552 8489 8572
rect 8378 8530 8489 8552
rect 8093 8517 8132 8524
rect 8802 8507 8836 8713
rect 9249 8693 9281 8721
rect 8869 8685 9281 8693
rect 10221 8719 10263 8772
rect 10221 8700 10230 8719
rect 10255 8700 10263 8719
rect 10221 8690 10263 8700
rect 10449 8730 10559 8744
rect 10449 8727 10527 8730
rect 10449 8700 10453 8727
rect 10482 8703 10527 8727
rect 10556 8703 10559 8730
rect 11179 8720 11213 8772
rect 11673 8763 11678 8783
rect 11699 8763 11705 8783
rect 11673 8756 11705 8763
rect 11883 8784 11921 8794
rect 12118 8791 12152 8997
rect 13226 9020 13268 9029
rect 13226 8998 13235 9020
rect 13261 8998 13268 9020
rect 13493 9047 13604 9064
rect 13493 9027 13500 9047
rect 13519 9027 13577 9047
rect 13596 9027 13604 9047
rect 13493 9005 13604 9027
rect 13778 9025 13812 9231
rect 14225 9211 14257 9239
rect 13845 9203 14257 9211
rect 13845 9177 13851 9203
rect 13877 9177 14257 9203
rect 15272 9211 15320 9366
rect 15506 9325 15616 9339
rect 15506 9322 15584 9325
rect 15506 9295 15510 9322
rect 15539 9298 15584 9322
rect 15613 9298 15616 9325
rect 16237 9315 16272 9366
rect 15539 9295 15616 9298
rect 15506 9280 15616 9295
rect 16235 9310 16272 9315
rect 16235 9290 16242 9310
rect 16262 9290 16272 9310
rect 16235 9283 16272 9290
rect 18745 9387 19108 9416
rect 18745 9385 18806 9387
rect 16235 9282 16270 9283
rect 15272 9182 15280 9211
rect 15309 9182 15320 9211
rect 15272 9177 15320 9182
rect 15791 9217 15823 9224
rect 15791 9197 15798 9217
rect 15819 9197 15823 9217
rect 13845 9175 14257 9177
rect 13847 9174 13887 9175
rect 14225 9110 14257 9175
rect 14225 9090 14229 9110
rect 14250 9090 14257 9110
rect 14225 9083 14257 9090
rect 15791 9132 15823 9197
rect 16161 9132 16201 9133
rect 15791 9130 16203 9132
rect 15791 9104 16171 9130
rect 16197 9104 16203 9130
rect 15791 9096 16203 9104
rect 15791 9068 15823 9096
rect 16236 9076 16270 9282
rect 18287 9165 18324 9167
rect 18745 9165 18778 9385
rect 19066 9306 19108 9387
rect 19488 9398 19599 9415
rect 19488 9378 19495 9398
rect 19514 9378 19572 9398
rect 19591 9378 19599 9398
rect 19488 9356 19599 9378
rect 18855 9304 18890 9305
rect 17174 9149 17208 9150
rect 16305 9114 17209 9149
rect 18287 9136 18778 9165
rect 15791 9048 15796 9068
rect 15817 9048 15823 9068
rect 15791 9041 15823 9048
rect 15998 9068 16037 9074
rect 15998 9048 16006 9068
rect 16031 9048 16037 9068
rect 15998 9041 16037 9048
rect 16214 9071 16270 9076
rect 16214 9051 16221 9071
rect 16241 9051 16270 9071
rect 16214 9044 16270 9051
rect 16214 9043 16249 9044
rect 13778 9017 13813 9025
rect 13226 8988 13268 8998
rect 13778 8997 13786 9017
rect 13806 8997 13813 9017
rect 13778 8992 13813 8997
rect 14432 9012 14542 9027
rect 14432 9009 14509 9012
rect 13226 8987 13267 8988
rect 12860 8953 12895 8954
rect 11883 8767 11893 8784
rect 11913 8767 11921 8784
rect 11724 8724 11765 8725
rect 10482 8700 10559 8703
rect 10449 8685 10559 8700
rect 11178 8715 11213 8720
rect 11178 8695 11185 8715
rect 11205 8695 11213 8715
rect 11723 8714 11765 8724
rect 11178 8687 11213 8695
rect 8869 8659 8875 8685
rect 8901 8659 9281 8685
rect 8869 8657 9281 8659
rect 8871 8656 8911 8657
rect 9249 8592 9281 8657
rect 10734 8622 10766 8629
rect 9249 8572 9253 8592
rect 9274 8572 9281 8592
rect 9249 8565 9281 8572
rect 9752 8607 9800 8612
rect 9752 8578 9763 8607
rect 9792 8578 9800 8607
rect 8802 8506 8837 8507
rect 8800 8499 8837 8506
rect 7745 8478 7780 8479
rect 7286 8474 7318 8475
rect 6908 8448 6916 8465
rect 6936 8448 6946 8465
rect 6908 8442 6946 8448
rect 7283 8469 7318 8474
rect 7283 8449 7290 8469
rect 7310 8449 7318 8469
rect 7283 8441 7318 8449
rect 6266 8402 6327 8404
rect 5964 8373 6327 8402
rect 6839 8376 6871 8383
rect 5964 8371 6266 8373
rect 3744 8355 4743 8358
rect 6839 8356 6846 8376
rect 6867 8356 6871 8376
rect 3744 8353 3779 8355
rect 2735 8349 3147 8351
rect 2737 8348 2777 8349
rect 1989 8164 1996 8185
rect 2023 8164 2031 8185
rect 1149 8134 1186 8141
rect 1149 8133 1184 8134
rect 186 8033 194 8062
rect 223 8033 234 8062
rect 186 8028 234 8033
rect 705 8068 737 8075
rect 705 8048 712 8068
rect 733 8048 737 8068
rect 705 7983 737 8048
rect 1075 7983 1115 7984
rect 705 7981 1117 7983
rect 705 7955 1085 7981
rect 1111 7955 1117 7981
rect 705 7947 1117 7955
rect 705 7919 737 7947
rect 1150 7927 1184 8133
rect 1854 8116 1893 8123
rect 1497 8088 1608 8110
rect 1497 8068 1505 8088
rect 1524 8068 1582 8088
rect 1601 8068 1608 8088
rect 1497 8051 1608 8068
rect 1854 8089 1858 8116
rect 1889 8089 1893 8116
rect 1701 8000 1754 8004
rect 1219 7965 1754 8000
rect 705 7899 710 7919
rect 731 7899 737 7919
rect 705 7892 737 7899
rect 912 7919 951 7925
rect 912 7899 920 7919
rect 945 7899 951 7919
rect 912 7892 951 7899
rect 1128 7922 1184 7927
rect 1128 7902 1135 7922
rect 1155 7902 1184 7922
rect 1128 7895 1184 7902
rect 1128 7894 1163 7895
rect 920 7846 951 7892
rect 419 7821 530 7843
rect 419 7801 427 7821
rect 446 7801 504 7821
rect 523 7801 530 7821
rect 919 7829 951 7846
rect 1220 7829 1257 7965
rect 1358 7932 1468 7946
rect 1358 7929 1436 7932
rect 1358 7902 1362 7929
rect 1391 7905 1436 7929
rect 1465 7905 1468 7932
rect 1391 7902 1468 7905
rect 1358 7887 1468 7902
rect 1700 7918 1754 7965
rect 1700 7910 1753 7918
rect 1700 7893 1709 7910
rect 1741 7893 1753 7910
rect 1700 7890 1753 7893
rect 919 7816 1257 7829
rect 419 7784 530 7801
rect 920 7797 1257 7816
rect 1199 7796 1257 7797
rect 1643 7824 1675 7831
rect 1643 7804 1650 7824
rect 1671 7804 1675 7824
rect 1643 7739 1675 7804
rect 1854 7816 1893 8089
rect 1989 7993 2031 8164
rect 2206 8189 2262 8194
rect 2206 8169 2213 8189
rect 2233 8169 2262 8189
rect 2206 8162 2262 8169
rect 2669 8199 2702 8257
rect 2899 8309 2937 8319
rect 2899 8271 2908 8309
rect 2931 8271 2937 8309
rect 2669 8191 2703 8199
rect 2669 8171 2676 8191
rect 2696 8171 2703 8191
rect 2669 8166 2703 8171
rect 2669 8165 2700 8166
rect 2206 8161 2241 8162
rect 2899 8135 2937 8271
rect 3115 8284 3147 8349
rect 6839 8291 6871 8356
rect 7209 8291 7249 8292
rect 6839 8289 7251 8291
rect 6207 8285 6242 8287
rect 3115 8264 3119 8284
rect 3140 8264 3147 8284
rect 5243 8282 6242 8285
rect 3720 8267 4022 8269
rect 3115 8257 3147 8264
rect 3659 8238 4022 8267
rect 3659 8236 3720 8238
rect 3040 8192 3078 8198
rect 3040 8175 3050 8192
rect 3070 8175 3078 8192
rect 1989 7959 2233 7993
rect 2899 7981 2943 8135
rect 2736 7979 2943 7981
rect 2196 7951 2233 7959
rect 2089 7918 2123 7929
rect 2087 7917 2123 7918
rect 2087 7897 2094 7917
rect 2114 7897 2123 7917
rect 2087 7889 2123 7897
rect 1854 7775 1861 7816
rect 1882 7775 1893 7816
rect 1854 7760 1893 7775
rect 2013 7739 2053 7740
rect 1643 7737 2055 7739
rect 1643 7711 2023 7737
rect 2049 7711 2055 7737
rect 1643 7703 2055 7711
rect 189 7664 1185 7690
rect 1643 7675 1675 7703
rect 2088 7683 2122 7889
rect 191 7611 233 7664
rect 191 7592 200 7611
rect 225 7592 233 7611
rect 191 7582 233 7592
rect 419 7622 529 7636
rect 419 7619 497 7622
rect 419 7592 423 7619
rect 452 7595 497 7619
rect 526 7595 529 7622
rect 1149 7612 1183 7664
rect 1643 7655 1648 7675
rect 1669 7655 1675 7675
rect 1643 7648 1675 7655
rect 2066 7678 2122 7683
rect 2066 7658 2073 7678
rect 2093 7658 2122 7678
rect 2066 7651 2122 7658
rect 2066 7650 2101 7651
rect 1694 7616 1735 7617
rect 452 7592 529 7595
rect 419 7577 529 7592
rect 1148 7607 1183 7612
rect 1148 7587 1155 7607
rect 1175 7587 1183 7607
rect 1693 7606 1735 7616
rect 1148 7579 1183 7587
rect 704 7514 736 7521
rect 704 7494 711 7514
rect 732 7494 736 7514
rect 704 7429 736 7494
rect 1074 7429 1114 7430
rect 704 7427 1116 7429
rect 704 7401 1084 7427
rect 1110 7401 1116 7427
rect 704 7393 1116 7401
rect 704 7365 736 7393
rect 1149 7373 1183 7579
rect 1357 7577 1468 7599
rect 1357 7557 1365 7577
rect 1384 7557 1442 7577
rect 1461 7557 1468 7577
rect 1357 7540 1468 7557
rect 1693 7584 1700 7606
rect 1726 7584 1735 7606
rect 1693 7575 1735 7584
rect 910 7370 953 7372
rect 704 7345 709 7365
rect 730 7345 736 7365
rect 704 7338 736 7345
rect 909 7363 953 7370
rect 909 7343 919 7363
rect 942 7343 953 7363
rect 909 7339 953 7343
rect 1127 7368 1183 7373
rect 1127 7348 1134 7368
rect 1154 7348 1183 7368
rect 1127 7341 1183 7348
rect 1239 7509 1272 7510
rect 1693 7509 1730 7575
rect 1239 7480 1730 7509
rect 1127 7340 1162 7341
rect 418 7267 529 7289
rect 418 7247 426 7267
rect 445 7247 503 7267
rect 522 7247 529 7267
rect 418 7231 529 7247
rect 909 7258 951 7339
rect 1239 7260 1272 7480
rect 1693 7478 1730 7480
rect 1468 7353 1578 7367
rect 1468 7350 1546 7353
rect 1468 7323 1472 7350
rect 1501 7326 1546 7350
rect 1575 7326 1578 7353
rect 1501 7323 1578 7326
rect 1468 7308 1578 7323
rect 2196 7338 2234 7951
rect 2712 7946 2943 7979
rect 2712 7405 2762 7946
rect 2899 7942 2943 7946
rect 2830 7845 2865 7846
rect 2809 7838 2865 7845
rect 2809 7818 2838 7838
rect 2858 7818 2865 7838
rect 2809 7813 2865 7818
rect 3040 7837 3078 8175
rect 3322 8186 3432 8201
rect 3322 8183 3399 8186
rect 3322 8156 3325 8183
rect 3354 8159 3399 8183
rect 3428 8159 3432 8186
rect 3354 8156 3432 8159
rect 3322 8142 3432 8156
rect 3201 8016 3238 8018
rect 3659 8016 3692 8236
rect 3980 8157 4022 8238
rect 4402 8249 4513 8266
rect 4402 8229 4409 8249
rect 4428 8229 4486 8249
rect 4505 8229 4513 8249
rect 4402 8207 4513 8229
rect 5242 8258 6242 8282
rect 3769 8155 3804 8156
rect 3201 7987 3692 8016
rect 3201 7921 3238 7987
rect 3659 7986 3692 7987
rect 3748 8148 3804 8155
rect 3748 8128 3777 8148
rect 3797 8128 3804 8148
rect 3748 8123 3804 8128
rect 3978 8153 4022 8157
rect 3978 8133 3989 8153
rect 4012 8133 4022 8153
rect 3978 8126 4022 8133
rect 4195 8151 4227 8158
rect 4195 8131 4201 8151
rect 4222 8131 4227 8151
rect 3978 8124 4021 8126
rect 3196 7912 3238 7921
rect 3196 7890 3205 7912
rect 3231 7890 3238 7912
rect 3463 7939 3574 7956
rect 3463 7919 3470 7939
rect 3489 7919 3547 7939
rect 3566 7919 3574 7939
rect 3463 7897 3574 7919
rect 3748 7917 3782 8123
rect 4195 8103 4227 8131
rect 3815 8095 4227 8103
rect 3815 8069 3821 8095
rect 3847 8069 4227 8095
rect 5242 8103 5290 8258
rect 5476 8217 5586 8231
rect 5476 8214 5554 8217
rect 5476 8187 5480 8214
rect 5509 8190 5554 8214
rect 5583 8190 5586 8217
rect 6207 8207 6242 8258
rect 5509 8187 5586 8190
rect 5476 8172 5586 8187
rect 6205 8202 6242 8207
rect 6205 8182 6212 8202
rect 6232 8182 6242 8202
rect 6839 8263 7219 8289
rect 7245 8263 7251 8289
rect 6839 8255 7251 8263
rect 6839 8227 6871 8255
rect 6839 8207 6844 8227
rect 6865 8207 6871 8227
rect 6839 8200 6871 8207
rect 7045 8226 7087 8237
rect 7284 8235 7318 8441
rect 7722 8471 7780 8478
rect 7722 8451 7753 8471
rect 7773 8451 7780 8471
rect 7722 8446 7780 8451
rect 8171 8474 8203 8481
rect 8171 8454 8177 8474
rect 8198 8454 8203 8474
rect 7722 8298 7758 8446
rect 8171 8426 8203 8454
rect 7791 8418 8203 8426
rect 7791 8392 7797 8418
rect 7823 8392 8203 8418
rect 8800 8479 8810 8499
rect 8830 8479 8837 8499
rect 8800 8474 8837 8479
rect 9456 8494 9566 8509
rect 9456 8491 9533 8494
rect 8800 8423 8835 8474
rect 9456 8464 9459 8491
rect 9488 8467 9533 8491
rect 9562 8467 9566 8494
rect 9488 8464 9566 8467
rect 9456 8450 9566 8464
rect 9752 8423 9800 8578
rect 10734 8602 10741 8622
rect 10762 8602 10766 8622
rect 10734 8537 10766 8602
rect 11104 8537 11144 8538
rect 10734 8535 11146 8537
rect 10734 8509 11114 8535
rect 11140 8509 11146 8535
rect 10734 8501 11146 8509
rect 10734 8473 10766 8501
rect 11179 8481 11213 8687
rect 11387 8685 11498 8707
rect 11387 8665 11395 8685
rect 11414 8665 11472 8685
rect 11491 8665 11498 8685
rect 11387 8648 11498 8665
rect 11723 8692 11730 8714
rect 11756 8692 11765 8714
rect 11723 8683 11765 8692
rect 10940 8478 10983 8480
rect 10734 8453 10739 8473
rect 10760 8453 10766 8473
rect 10734 8446 10766 8453
rect 10939 8471 10983 8478
rect 10939 8451 10949 8471
rect 10972 8451 10983 8471
rect 10939 8447 10983 8451
rect 11157 8476 11213 8481
rect 11157 8456 11164 8476
rect 11184 8456 11213 8476
rect 11157 8449 11213 8456
rect 11269 8617 11302 8618
rect 11723 8617 11760 8683
rect 11269 8588 11760 8617
rect 11157 8448 11192 8449
rect 8800 8399 9800 8423
rect 8800 8396 9799 8399
rect 8800 8394 8835 8396
rect 7791 8390 8203 8392
rect 7793 8389 7833 8390
rect 7045 8205 7052 8226
rect 7079 8205 7087 8226
rect 6205 8175 6242 8182
rect 6205 8174 6240 8175
rect 5242 8074 5250 8103
rect 5279 8074 5290 8103
rect 5242 8069 5290 8074
rect 5761 8109 5793 8116
rect 5761 8089 5768 8109
rect 5789 8089 5793 8109
rect 3815 8067 4227 8069
rect 3817 8066 3857 8067
rect 4195 8002 4227 8067
rect 4195 7982 4199 8002
rect 4220 7982 4227 8002
rect 4195 7975 4227 7982
rect 5761 8024 5793 8089
rect 6131 8024 6171 8025
rect 5761 8022 6173 8024
rect 5761 7996 6141 8022
rect 6167 7996 6173 8022
rect 5761 7988 6173 7996
rect 5761 7960 5793 7988
rect 6206 7968 6240 8174
rect 6910 8157 6949 8164
rect 6553 8129 6664 8151
rect 6553 8109 6561 8129
rect 6580 8109 6638 8129
rect 6657 8109 6664 8129
rect 6553 8092 6664 8109
rect 6910 8130 6914 8157
rect 6945 8130 6949 8157
rect 6757 8041 6810 8045
rect 6275 8006 6810 8041
rect 5761 7940 5766 7960
rect 5787 7940 5793 7960
rect 5761 7933 5793 7940
rect 5968 7960 6007 7966
rect 5968 7940 5976 7960
rect 6001 7940 6007 7960
rect 5968 7933 6007 7940
rect 6184 7963 6240 7968
rect 6184 7943 6191 7963
rect 6211 7943 6240 7963
rect 6184 7936 6240 7943
rect 6184 7935 6219 7936
rect 3748 7909 3783 7917
rect 3196 7880 3238 7890
rect 3748 7889 3756 7909
rect 3776 7889 3783 7909
rect 3748 7884 3783 7889
rect 4402 7904 4512 7919
rect 4402 7901 4479 7904
rect 3196 7879 3237 7880
rect 3040 7820 3048 7837
rect 3068 7820 3078 7837
rect 2809 7607 2843 7813
rect 3040 7810 3078 7820
rect 3256 7841 3288 7848
rect 3256 7821 3262 7841
rect 3283 7821 3288 7841
rect 3748 7832 3782 7884
rect 4402 7874 4405 7901
rect 4434 7877 4479 7901
rect 4508 7877 4512 7904
rect 4434 7874 4512 7877
rect 4402 7860 4512 7874
rect 4698 7904 4740 7914
rect 4698 7885 4706 7904
rect 4731 7885 4740 7904
rect 5976 7887 6007 7933
rect 4698 7832 4740 7885
rect 5475 7862 5586 7884
rect 5475 7842 5483 7862
rect 5502 7842 5560 7862
rect 5579 7842 5586 7862
rect 5975 7870 6007 7887
rect 6276 7870 6313 8006
rect 6414 7973 6524 7987
rect 6414 7970 6492 7973
rect 6414 7943 6418 7970
rect 6447 7946 6492 7970
rect 6521 7946 6524 7973
rect 6447 7943 6524 7946
rect 6414 7928 6524 7943
rect 6756 7959 6810 8006
rect 6756 7951 6809 7959
rect 6756 7934 6765 7951
rect 6797 7934 6809 7951
rect 6756 7931 6809 7934
rect 5975 7857 6313 7870
rect 3256 7793 3288 7821
rect 3746 7806 4742 7832
rect 5475 7825 5586 7842
rect 5976 7838 6313 7857
rect 6255 7837 6313 7838
rect 6699 7865 6731 7872
rect 6699 7845 6706 7865
rect 6727 7845 6731 7865
rect 2876 7785 3288 7793
rect 2876 7759 2882 7785
rect 2908 7759 3288 7785
rect 2876 7757 3288 7759
rect 2878 7756 2918 7757
rect 3256 7692 3288 7757
rect 6699 7780 6731 7845
rect 6910 7857 6949 8130
rect 7045 8034 7087 8205
rect 7262 8230 7318 8235
rect 7262 8210 7269 8230
rect 7289 8210 7318 8230
rect 7262 8203 7318 8210
rect 7725 8240 7758 8298
rect 7955 8350 7993 8360
rect 7955 8312 7964 8350
rect 7987 8312 7993 8350
rect 7725 8232 7759 8240
rect 7725 8212 7732 8232
rect 7752 8212 7759 8232
rect 7725 8207 7759 8212
rect 7725 8206 7756 8207
rect 7262 8202 7297 8203
rect 7955 8176 7993 8312
rect 8171 8325 8203 8390
rect 10448 8375 10559 8397
rect 10448 8355 10456 8375
rect 10475 8355 10533 8375
rect 10552 8355 10559 8375
rect 10448 8338 10559 8355
rect 10939 8366 10981 8447
rect 11269 8368 11302 8588
rect 11723 8586 11760 8588
rect 11529 8448 11639 8462
rect 11529 8445 11607 8448
rect 11529 8418 11533 8445
rect 11562 8421 11607 8445
rect 11636 8421 11639 8448
rect 11562 8418 11639 8421
rect 11529 8403 11639 8418
rect 11883 8429 11921 8767
rect 12096 8786 12152 8791
rect 12096 8766 12103 8786
rect 12123 8766 12152 8786
rect 12096 8759 12152 8766
rect 12839 8946 12895 8953
rect 12839 8926 12868 8946
rect 12888 8926 12895 8946
rect 12839 8921 12895 8926
rect 13286 8949 13318 8956
rect 13286 8929 13292 8949
rect 13313 8929 13318 8949
rect 13778 8940 13812 8992
rect 14432 8982 14435 9009
rect 14464 8985 14509 9009
rect 14538 8985 14542 9012
rect 14464 8982 14542 8985
rect 14432 8968 14542 8982
rect 14728 9012 14770 9022
rect 14728 8993 14736 9012
rect 14761 8993 14770 9012
rect 16006 8995 16037 9041
rect 14728 8940 14770 8993
rect 15505 8970 15616 8992
rect 15505 8950 15513 8970
rect 15532 8950 15590 8970
rect 15609 8950 15616 8970
rect 16005 8978 16037 8995
rect 16306 8978 16343 9114
rect 16444 9081 16554 9095
rect 16444 9078 16522 9081
rect 16444 9051 16448 9078
rect 16477 9054 16522 9078
rect 16551 9054 16554 9081
rect 17174 9071 17208 9114
rect 16477 9051 16554 9054
rect 16444 9036 16554 9051
rect 17173 9066 17208 9071
rect 18287 9070 18324 9136
rect 18745 9135 18778 9136
rect 18834 9297 18890 9304
rect 18834 9277 18863 9297
rect 18883 9277 18890 9297
rect 18834 9272 18890 9277
rect 19064 9302 19108 9306
rect 19064 9282 19075 9302
rect 19098 9282 19108 9302
rect 19064 9275 19108 9282
rect 19281 9300 19313 9307
rect 19281 9280 19287 9300
rect 19308 9280 19313 9300
rect 19064 9273 19107 9275
rect 17173 9046 17180 9066
rect 17200 9046 17208 9066
rect 17173 9038 17208 9046
rect 16005 8965 16343 8978
rect 12096 8758 12131 8759
rect 12839 8715 12873 8921
rect 13286 8901 13318 8929
rect 13776 8914 14772 8940
rect 15505 8933 15616 8950
rect 16006 8946 16343 8965
rect 16285 8945 16343 8946
rect 16729 8973 16761 8980
rect 16729 8953 16736 8973
rect 16757 8953 16761 8973
rect 12906 8893 13318 8901
rect 12906 8867 12912 8893
rect 12938 8867 13318 8893
rect 12906 8865 13318 8867
rect 12908 8864 12948 8865
rect 13068 8829 13107 8844
rect 13068 8788 13079 8829
rect 13100 8788 13107 8829
rect 12838 8707 12874 8715
rect 12838 8687 12847 8707
rect 12867 8687 12874 8707
rect 12838 8686 12874 8687
rect 12838 8675 12872 8686
rect 13068 8515 13107 8788
rect 13286 8800 13318 8865
rect 16729 8888 16761 8953
rect 17099 8888 17139 8889
rect 16729 8886 17141 8888
rect 16729 8860 17109 8886
rect 17135 8860 17141 8886
rect 16729 8852 17141 8860
rect 13286 8780 13290 8800
rect 13311 8780 13318 8800
rect 13286 8773 13318 8780
rect 13704 8807 13762 8808
rect 13704 8788 14041 8807
rect 14431 8803 14542 8820
rect 15275 8813 16271 8839
rect 16729 8824 16761 8852
rect 13704 8775 14042 8788
rect 13208 8711 13261 8714
rect 13208 8694 13220 8711
rect 13252 8694 13261 8711
rect 13208 8686 13261 8694
rect 13207 8639 13261 8686
rect 13493 8702 13603 8717
rect 13493 8699 13570 8702
rect 13493 8672 13496 8699
rect 13525 8675 13570 8699
rect 13599 8675 13603 8702
rect 13525 8672 13603 8675
rect 13493 8658 13603 8672
rect 13704 8639 13741 8775
rect 14010 8758 14042 8775
rect 14431 8783 14438 8803
rect 14457 8783 14515 8803
rect 14534 8783 14542 8803
rect 14431 8761 14542 8783
rect 15277 8760 15319 8813
rect 14010 8712 14041 8758
rect 15277 8741 15286 8760
rect 15311 8741 15319 8760
rect 15277 8731 15319 8741
rect 15505 8771 15615 8785
rect 15505 8768 15583 8771
rect 15505 8741 15509 8768
rect 15538 8744 15583 8768
rect 15612 8744 15615 8771
rect 16235 8761 16269 8813
rect 16729 8804 16734 8824
rect 16755 8804 16761 8824
rect 16729 8797 16761 8804
rect 16939 8825 16977 8835
rect 17174 8832 17208 9038
rect 18282 9061 18324 9070
rect 18282 9039 18291 9061
rect 18317 9039 18324 9061
rect 18549 9088 18660 9105
rect 18549 9068 18556 9088
rect 18575 9068 18633 9088
rect 18652 9068 18660 9088
rect 18549 9046 18660 9068
rect 18834 9066 18868 9272
rect 19281 9252 19313 9280
rect 18901 9244 19313 9252
rect 18901 9218 18907 9244
rect 18933 9218 19313 9244
rect 18901 9216 19313 9218
rect 18903 9215 18943 9216
rect 19281 9151 19313 9216
rect 19281 9131 19285 9151
rect 19306 9131 19313 9151
rect 19281 9124 19313 9131
rect 18834 9058 18869 9066
rect 18282 9029 18324 9039
rect 18834 9038 18842 9058
rect 18862 9038 18869 9058
rect 18834 9033 18869 9038
rect 19488 9053 19598 9068
rect 19488 9050 19565 9053
rect 18282 9028 18323 9029
rect 17916 8994 17951 8995
rect 16939 8808 16949 8825
rect 16969 8808 16977 8825
rect 16780 8765 16821 8766
rect 15538 8741 15615 8744
rect 15505 8726 15615 8741
rect 16234 8756 16269 8761
rect 16234 8736 16241 8756
rect 16261 8736 16269 8756
rect 16779 8755 16821 8765
rect 16234 8728 16269 8736
rect 13798 8709 13833 8710
rect 13777 8702 13833 8709
rect 13777 8682 13806 8702
rect 13826 8682 13833 8702
rect 13777 8677 13833 8682
rect 14010 8705 14049 8712
rect 14010 8685 14016 8705
rect 14041 8685 14049 8705
rect 14010 8679 14049 8685
rect 14224 8705 14256 8712
rect 14224 8685 14230 8705
rect 14251 8685 14256 8705
rect 13207 8604 13742 8639
rect 13207 8600 13260 8604
rect 13068 8488 13072 8515
rect 13103 8488 13107 8515
rect 13353 8536 13464 8553
rect 13353 8516 13360 8536
rect 13379 8516 13437 8536
rect 13456 8516 13464 8536
rect 13353 8494 13464 8516
rect 13068 8481 13107 8488
rect 13777 8471 13811 8677
rect 14224 8657 14256 8685
rect 13844 8649 14256 8657
rect 13844 8623 13850 8649
rect 13876 8623 14256 8649
rect 13844 8621 14256 8623
rect 13846 8620 13886 8621
rect 14224 8556 14256 8621
rect 15790 8663 15822 8670
rect 15790 8643 15797 8663
rect 15818 8643 15822 8663
rect 15790 8578 15822 8643
rect 16160 8578 16200 8579
rect 15790 8576 16202 8578
rect 14224 8536 14228 8556
rect 14249 8536 14256 8556
rect 14224 8529 14256 8536
rect 14727 8571 14775 8576
rect 14727 8542 14738 8571
rect 14767 8542 14775 8571
rect 13777 8470 13812 8471
rect 13775 8463 13812 8470
rect 12720 8442 12755 8443
rect 12261 8438 12293 8439
rect 11883 8412 11891 8429
rect 11911 8412 11921 8429
rect 11883 8406 11921 8412
rect 12258 8433 12293 8438
rect 12258 8413 12265 8433
rect 12285 8413 12293 8433
rect 12258 8405 12293 8413
rect 11241 8366 11302 8368
rect 10939 8337 11302 8366
rect 11814 8340 11846 8347
rect 10939 8335 11241 8337
rect 8171 8305 8175 8325
rect 8196 8305 8203 8325
rect 11814 8320 11821 8340
rect 11842 8320 11846 8340
rect 8776 8308 9078 8310
rect 8171 8298 8203 8305
rect 8715 8279 9078 8308
rect 8715 8277 8776 8279
rect 8096 8233 8134 8239
rect 8096 8216 8106 8233
rect 8126 8216 8134 8233
rect 7045 8000 7289 8034
rect 7955 8022 7999 8176
rect 7792 8020 7999 8022
rect 7252 7992 7289 8000
rect 7145 7959 7179 7970
rect 7143 7958 7179 7959
rect 7143 7938 7150 7958
rect 7170 7938 7179 7958
rect 7143 7930 7179 7938
rect 6910 7816 6917 7857
rect 6938 7816 6949 7857
rect 6910 7801 6949 7816
rect 7069 7780 7109 7781
rect 6699 7778 7111 7780
rect 6699 7752 7079 7778
rect 7105 7752 7111 7778
rect 6699 7744 7111 7752
rect 3256 7672 3260 7692
rect 3281 7672 3288 7692
rect 3256 7665 3288 7672
rect 3674 7699 3732 7700
rect 3674 7680 4011 7699
rect 4401 7695 4512 7712
rect 5245 7705 6241 7731
rect 6699 7716 6731 7744
rect 7144 7724 7178 7930
rect 3674 7667 4012 7680
rect 2809 7599 2844 7607
rect 2809 7579 2817 7599
rect 2837 7579 2844 7599
rect 2809 7574 2844 7579
rect 3463 7594 3573 7609
rect 3463 7591 3540 7594
rect 2809 7531 2843 7574
rect 3463 7564 3466 7591
rect 3495 7567 3540 7591
rect 3569 7567 3573 7594
rect 3495 7564 3573 7567
rect 3463 7550 3573 7564
rect 3674 7531 3711 7667
rect 3980 7650 4012 7667
rect 4401 7675 4408 7695
rect 4427 7675 4485 7695
rect 4504 7675 4512 7695
rect 4401 7653 4512 7675
rect 5247 7652 5289 7705
rect 3980 7604 4011 7650
rect 5247 7633 5256 7652
rect 5281 7633 5289 7652
rect 5247 7623 5289 7633
rect 5475 7663 5585 7677
rect 5475 7660 5553 7663
rect 5475 7633 5479 7660
rect 5508 7636 5553 7660
rect 5582 7636 5585 7663
rect 6205 7653 6239 7705
rect 6699 7696 6704 7716
rect 6725 7696 6731 7716
rect 6699 7689 6731 7696
rect 7122 7719 7178 7724
rect 7122 7699 7129 7719
rect 7149 7699 7178 7719
rect 7122 7692 7178 7699
rect 7122 7691 7157 7692
rect 6750 7657 6791 7658
rect 5508 7633 5585 7636
rect 5475 7618 5585 7633
rect 6204 7648 6239 7653
rect 6204 7628 6211 7648
rect 6231 7628 6239 7648
rect 6749 7647 6791 7657
rect 6204 7620 6239 7628
rect 3768 7601 3803 7602
rect 3747 7594 3803 7601
rect 3747 7574 3776 7594
rect 3796 7574 3803 7594
rect 3747 7569 3803 7574
rect 3980 7597 4019 7604
rect 3980 7577 3986 7597
rect 4011 7577 4019 7597
rect 3980 7571 4019 7577
rect 4194 7597 4226 7604
rect 4194 7577 4200 7597
rect 4221 7577 4226 7597
rect 2808 7496 3712 7531
rect 2809 7495 2843 7496
rect 2690 7396 2762 7405
rect 2690 7367 2707 7396
rect 2755 7367 2762 7396
rect 3353 7415 3464 7432
rect 3353 7395 3360 7415
rect 3379 7395 3437 7415
rect 3456 7395 3464 7415
rect 3353 7373 3464 7395
rect 2690 7360 2762 7367
rect 3747 7363 3781 7569
rect 4194 7549 4226 7577
rect 3814 7541 4226 7549
rect 3814 7515 3820 7541
rect 3846 7515 4226 7541
rect 3814 7513 4226 7515
rect 3816 7512 3856 7513
rect 4194 7448 4226 7513
rect 5760 7555 5792 7562
rect 5760 7535 5767 7555
rect 5788 7535 5792 7555
rect 5760 7470 5792 7535
rect 6130 7470 6170 7471
rect 5760 7468 6172 7470
rect 4194 7428 4198 7448
rect 4219 7428 4226 7448
rect 4194 7421 4226 7428
rect 4697 7463 4745 7468
rect 4697 7434 4708 7463
rect 4737 7434 4745 7463
rect 3747 7362 3782 7363
rect 2690 7350 2760 7360
rect 3745 7355 3782 7362
rect 2196 7318 2204 7338
rect 2224 7318 2234 7338
rect 3745 7335 3755 7355
rect 3775 7335 3782 7355
rect 3745 7330 3782 7335
rect 4401 7350 4511 7365
rect 4401 7347 4478 7350
rect 2720 7321 2755 7322
rect 2196 7311 2234 7318
rect 2699 7314 2755 7321
rect 2197 7310 2232 7311
rect 1211 7258 1272 7260
rect 909 7229 1272 7258
rect 1753 7245 1785 7252
rect 909 7227 1211 7229
rect 1753 7225 1760 7245
rect 1781 7225 1785 7245
rect 1753 7160 1785 7225
rect 2123 7160 2163 7161
rect 1753 7158 2165 7160
rect 1151 7141 1186 7143
rect 187 7138 1186 7141
rect 186 7114 1186 7138
rect 186 6959 234 7114
rect 420 7073 530 7087
rect 420 7070 498 7073
rect 420 7043 424 7070
rect 453 7046 498 7070
rect 527 7046 530 7073
rect 1151 7063 1186 7114
rect 1753 7132 2133 7158
rect 2159 7132 2165 7158
rect 1753 7124 2165 7132
rect 1753 7096 1785 7124
rect 1753 7076 1758 7096
rect 1779 7076 1785 7096
rect 1753 7069 1785 7076
rect 1959 7095 2004 7107
rect 2198 7104 2232 7310
rect 1959 7076 1966 7095
rect 1995 7076 2004 7095
rect 453 7043 530 7046
rect 420 7028 530 7043
rect 1149 7058 1186 7063
rect 1149 7038 1156 7058
rect 1176 7038 1186 7058
rect 1149 7031 1186 7038
rect 1149 7030 1184 7031
rect 186 6930 194 6959
rect 223 6930 234 6959
rect 186 6925 234 6930
rect 705 6965 737 6972
rect 705 6945 712 6965
rect 733 6945 737 6965
rect 705 6880 737 6945
rect 1075 6880 1115 6881
rect 705 6878 1117 6880
rect 705 6852 1085 6878
rect 1111 6852 1117 6878
rect 705 6844 1117 6852
rect 705 6816 737 6844
rect 1150 6824 1184 7030
rect 1467 6998 1578 7020
rect 1467 6978 1475 6998
rect 1494 6978 1552 6998
rect 1571 6978 1578 6998
rect 1467 6961 1578 6978
rect 1959 6993 2004 7076
rect 2176 7099 2232 7104
rect 2176 7079 2183 7099
rect 2203 7079 2232 7099
rect 2699 7294 2728 7314
rect 2748 7294 2755 7314
rect 2699 7289 2755 7294
rect 3146 7317 3178 7324
rect 3146 7297 3152 7317
rect 3173 7297 3178 7317
rect 2699 7083 2733 7289
rect 3146 7269 3178 7297
rect 2766 7261 3178 7269
rect 2766 7235 2772 7261
rect 2798 7235 3178 7261
rect 3745 7279 3780 7330
rect 4401 7320 4404 7347
rect 4433 7323 4478 7347
rect 4507 7323 4511 7350
rect 4433 7320 4511 7323
rect 4401 7306 4511 7320
rect 4697 7279 4745 7434
rect 5760 7442 6140 7468
rect 6166 7442 6172 7468
rect 5760 7434 6172 7442
rect 5760 7406 5792 7434
rect 6205 7414 6239 7620
rect 6413 7618 6524 7640
rect 6413 7598 6421 7618
rect 6440 7598 6498 7618
rect 6517 7598 6524 7618
rect 6413 7581 6524 7598
rect 6749 7625 6756 7647
rect 6782 7625 6791 7647
rect 6749 7616 6791 7625
rect 5966 7411 6009 7413
rect 5760 7386 5765 7406
rect 5786 7386 5792 7406
rect 5760 7379 5792 7386
rect 5965 7404 6009 7411
rect 5965 7384 5975 7404
rect 5998 7384 6009 7404
rect 5965 7380 6009 7384
rect 6183 7409 6239 7414
rect 6183 7389 6190 7409
rect 6210 7389 6239 7409
rect 6183 7382 6239 7389
rect 6295 7550 6328 7551
rect 6749 7550 6786 7616
rect 6295 7521 6786 7550
rect 6183 7381 6218 7382
rect 3745 7255 4745 7279
rect 5474 7308 5585 7330
rect 5474 7288 5482 7308
rect 5501 7288 5559 7308
rect 5578 7288 5585 7308
rect 5474 7272 5585 7288
rect 5965 7299 6007 7380
rect 6295 7301 6328 7521
rect 6749 7519 6786 7521
rect 6524 7394 6634 7408
rect 6524 7391 6602 7394
rect 6524 7364 6528 7391
rect 6557 7367 6602 7391
rect 6631 7367 6634 7394
rect 6557 7364 6634 7367
rect 6524 7349 6634 7364
rect 7252 7379 7290 7992
rect 7768 7987 7999 8020
rect 7768 7446 7818 7987
rect 7955 7983 7999 7987
rect 7886 7886 7921 7887
rect 7865 7879 7921 7886
rect 7865 7859 7894 7879
rect 7914 7859 7921 7879
rect 7865 7854 7921 7859
rect 8096 7878 8134 8216
rect 8378 8227 8488 8242
rect 8378 8224 8455 8227
rect 8378 8197 8381 8224
rect 8410 8200 8455 8224
rect 8484 8200 8488 8227
rect 8410 8197 8488 8200
rect 8378 8183 8488 8197
rect 8257 8057 8294 8059
rect 8715 8057 8748 8277
rect 9036 8198 9078 8279
rect 9458 8290 9569 8307
rect 9458 8270 9465 8290
rect 9484 8270 9542 8290
rect 9561 8270 9569 8290
rect 9458 8248 9569 8270
rect 11814 8255 11846 8320
rect 12184 8255 12224 8256
rect 11814 8253 12226 8255
rect 11182 8249 11217 8251
rect 10218 8246 11217 8249
rect 10217 8222 11217 8246
rect 8825 8196 8860 8197
rect 8257 8028 8748 8057
rect 8257 7962 8294 8028
rect 8715 8027 8748 8028
rect 8804 8189 8860 8196
rect 8804 8169 8833 8189
rect 8853 8169 8860 8189
rect 8804 8164 8860 8169
rect 9034 8194 9078 8198
rect 9034 8174 9045 8194
rect 9068 8174 9078 8194
rect 9034 8167 9078 8174
rect 9251 8192 9283 8199
rect 9251 8172 9257 8192
rect 9278 8172 9283 8192
rect 9034 8165 9077 8167
rect 8252 7953 8294 7962
rect 8252 7931 8261 7953
rect 8287 7931 8294 7953
rect 8519 7980 8630 7997
rect 8519 7960 8526 7980
rect 8545 7960 8603 7980
rect 8622 7960 8630 7980
rect 8519 7938 8630 7960
rect 8804 7958 8838 8164
rect 9251 8144 9283 8172
rect 8871 8136 9283 8144
rect 8871 8110 8877 8136
rect 8903 8110 9283 8136
rect 8871 8108 9283 8110
rect 8873 8107 8913 8108
rect 9251 8043 9283 8108
rect 9251 8023 9255 8043
rect 9276 8023 9283 8043
rect 10217 8067 10265 8222
rect 10451 8181 10561 8195
rect 10451 8178 10529 8181
rect 10451 8151 10455 8178
rect 10484 8154 10529 8178
rect 10558 8154 10561 8181
rect 11182 8171 11217 8222
rect 10484 8151 10561 8154
rect 10451 8136 10561 8151
rect 11180 8166 11217 8171
rect 11180 8146 11187 8166
rect 11207 8146 11217 8166
rect 11814 8227 12194 8253
rect 12220 8227 12226 8253
rect 11814 8219 12226 8227
rect 11814 8191 11846 8219
rect 11814 8171 11819 8191
rect 11840 8171 11846 8191
rect 11814 8164 11846 8171
rect 12020 8190 12062 8201
rect 12259 8199 12293 8405
rect 12697 8435 12755 8442
rect 12697 8415 12728 8435
rect 12748 8415 12755 8435
rect 12697 8410 12755 8415
rect 13146 8438 13178 8445
rect 13146 8418 13152 8438
rect 13173 8418 13178 8438
rect 12697 8262 12733 8410
rect 13146 8390 13178 8418
rect 12766 8382 13178 8390
rect 12766 8356 12772 8382
rect 12798 8356 13178 8382
rect 13775 8443 13785 8463
rect 13805 8443 13812 8463
rect 13775 8438 13812 8443
rect 14431 8458 14541 8473
rect 14431 8455 14508 8458
rect 13775 8387 13810 8438
rect 14431 8428 14434 8455
rect 14463 8431 14508 8455
rect 14537 8431 14541 8458
rect 14463 8428 14541 8431
rect 14431 8414 14541 8428
rect 14727 8387 14775 8542
rect 15790 8550 16170 8576
rect 16196 8550 16202 8576
rect 15790 8542 16202 8550
rect 15790 8514 15822 8542
rect 16235 8522 16269 8728
rect 16443 8726 16554 8748
rect 16443 8706 16451 8726
rect 16470 8706 16528 8726
rect 16547 8706 16554 8726
rect 16443 8689 16554 8706
rect 16779 8733 16786 8755
rect 16812 8733 16821 8755
rect 16779 8724 16821 8733
rect 15996 8519 16039 8521
rect 15790 8494 15795 8514
rect 15816 8494 15822 8514
rect 15790 8487 15822 8494
rect 15995 8512 16039 8519
rect 15995 8492 16005 8512
rect 16028 8492 16039 8512
rect 15995 8488 16039 8492
rect 16213 8517 16269 8522
rect 16213 8497 16220 8517
rect 16240 8497 16269 8517
rect 16213 8490 16269 8497
rect 16325 8658 16358 8659
rect 16779 8658 16816 8724
rect 16325 8629 16816 8658
rect 16213 8489 16248 8490
rect 13775 8363 14775 8387
rect 15504 8416 15615 8438
rect 15504 8396 15512 8416
rect 15531 8396 15589 8416
rect 15608 8396 15615 8416
rect 15504 8379 15615 8396
rect 15995 8407 16037 8488
rect 16325 8409 16358 8629
rect 16779 8627 16816 8629
rect 16585 8489 16695 8503
rect 16585 8486 16663 8489
rect 16585 8459 16589 8486
rect 16618 8462 16663 8486
rect 16692 8462 16695 8489
rect 16618 8459 16695 8462
rect 16585 8444 16695 8459
rect 16939 8470 16977 8808
rect 17152 8827 17208 8832
rect 17152 8807 17159 8827
rect 17179 8807 17208 8827
rect 17152 8800 17208 8807
rect 17895 8987 17951 8994
rect 17895 8967 17924 8987
rect 17944 8967 17951 8987
rect 17895 8962 17951 8967
rect 18342 8990 18374 8997
rect 18342 8970 18348 8990
rect 18369 8970 18374 8990
rect 18834 8981 18868 9033
rect 19488 9023 19491 9050
rect 19520 9026 19565 9050
rect 19594 9026 19598 9053
rect 19520 9023 19598 9026
rect 19488 9009 19598 9023
rect 19784 9053 19826 9063
rect 19784 9034 19792 9053
rect 19817 9034 19826 9053
rect 19784 8981 19826 9034
rect 17152 8799 17187 8800
rect 17895 8756 17929 8962
rect 18342 8942 18374 8970
rect 18832 8955 19828 8981
rect 17962 8934 18374 8942
rect 17962 8908 17968 8934
rect 17994 8908 18374 8934
rect 17962 8906 18374 8908
rect 17964 8905 18004 8906
rect 18124 8870 18163 8885
rect 18124 8829 18135 8870
rect 18156 8829 18163 8870
rect 17894 8748 17930 8756
rect 17894 8728 17903 8748
rect 17923 8728 17930 8748
rect 17894 8727 17930 8728
rect 17894 8716 17928 8727
rect 18124 8556 18163 8829
rect 18342 8841 18374 8906
rect 18342 8821 18346 8841
rect 18367 8821 18374 8841
rect 18342 8814 18374 8821
rect 18760 8848 18818 8849
rect 18760 8829 19097 8848
rect 19487 8844 19598 8861
rect 18760 8816 19098 8829
rect 18264 8752 18317 8755
rect 18264 8735 18276 8752
rect 18308 8735 18317 8752
rect 18264 8727 18317 8735
rect 18263 8680 18317 8727
rect 18549 8743 18659 8758
rect 18549 8740 18626 8743
rect 18549 8713 18552 8740
rect 18581 8716 18626 8740
rect 18655 8716 18659 8743
rect 18581 8713 18659 8716
rect 18549 8699 18659 8713
rect 18760 8680 18797 8816
rect 19066 8799 19098 8816
rect 19487 8824 19494 8844
rect 19513 8824 19571 8844
rect 19590 8824 19598 8844
rect 19487 8802 19598 8824
rect 19066 8753 19097 8799
rect 18854 8750 18889 8751
rect 18833 8743 18889 8750
rect 18833 8723 18862 8743
rect 18882 8723 18889 8743
rect 18833 8718 18889 8723
rect 19066 8746 19105 8753
rect 19066 8726 19072 8746
rect 19097 8726 19105 8746
rect 19066 8720 19105 8726
rect 19280 8746 19312 8753
rect 19280 8726 19286 8746
rect 19307 8726 19312 8746
rect 18263 8645 18798 8680
rect 18263 8641 18316 8645
rect 18124 8529 18128 8556
rect 18159 8529 18163 8556
rect 18409 8577 18520 8594
rect 18409 8557 18416 8577
rect 18435 8557 18493 8577
rect 18512 8557 18520 8577
rect 18409 8535 18520 8557
rect 18124 8522 18163 8529
rect 18833 8512 18867 8718
rect 19280 8698 19312 8726
rect 18900 8690 19312 8698
rect 18900 8664 18906 8690
rect 18932 8664 19312 8690
rect 18900 8662 19312 8664
rect 18902 8661 18942 8662
rect 19280 8597 19312 8662
rect 19280 8577 19284 8597
rect 19305 8577 19312 8597
rect 19280 8570 19312 8577
rect 19783 8612 19831 8617
rect 19783 8583 19794 8612
rect 19823 8583 19831 8612
rect 18833 8511 18868 8512
rect 18831 8504 18868 8511
rect 17776 8483 17811 8484
rect 17317 8479 17349 8480
rect 16939 8453 16947 8470
rect 16967 8453 16977 8470
rect 16939 8447 16977 8453
rect 17314 8474 17349 8479
rect 17314 8454 17321 8474
rect 17341 8454 17349 8474
rect 17314 8446 17349 8454
rect 16297 8407 16358 8409
rect 15995 8378 16358 8407
rect 16870 8381 16902 8388
rect 15995 8376 16297 8378
rect 13775 8360 14774 8363
rect 16870 8361 16877 8381
rect 16898 8361 16902 8381
rect 13775 8358 13810 8360
rect 12766 8354 13178 8356
rect 12768 8353 12808 8354
rect 12020 8169 12027 8190
rect 12054 8169 12062 8190
rect 11180 8139 11217 8146
rect 11180 8138 11215 8139
rect 10217 8038 10225 8067
rect 10254 8038 10265 8067
rect 10217 8033 10265 8038
rect 10736 8073 10768 8080
rect 10736 8053 10743 8073
rect 10764 8053 10768 8073
rect 9251 8016 9283 8023
rect 10736 7988 10768 8053
rect 11106 7988 11146 7989
rect 10736 7986 11148 7988
rect 10736 7960 11116 7986
rect 11142 7960 11148 7986
rect 8804 7950 8839 7958
rect 8252 7921 8294 7931
rect 8804 7930 8812 7950
rect 8832 7930 8839 7950
rect 8804 7925 8839 7930
rect 9458 7945 9568 7960
rect 9458 7942 9535 7945
rect 8252 7920 8293 7921
rect 8096 7861 8104 7878
rect 8124 7861 8134 7878
rect 7865 7648 7899 7854
rect 8096 7851 8134 7861
rect 8312 7882 8344 7889
rect 8312 7862 8318 7882
rect 8339 7862 8344 7882
rect 8804 7873 8838 7925
rect 9458 7915 9461 7942
rect 9490 7918 9535 7942
rect 9564 7918 9568 7945
rect 9490 7915 9568 7918
rect 9458 7901 9568 7915
rect 9754 7945 9796 7955
rect 9754 7926 9762 7945
rect 9787 7926 9796 7945
rect 9754 7873 9796 7926
rect 10736 7952 11148 7960
rect 10736 7924 10768 7952
rect 11181 7932 11215 8138
rect 11885 8121 11924 8128
rect 11528 8093 11639 8115
rect 11528 8073 11536 8093
rect 11555 8073 11613 8093
rect 11632 8073 11639 8093
rect 11528 8056 11639 8073
rect 11885 8094 11889 8121
rect 11920 8094 11924 8121
rect 11732 8005 11785 8009
rect 11250 7970 11785 8005
rect 10736 7904 10741 7924
rect 10762 7904 10768 7924
rect 10736 7897 10768 7904
rect 10943 7924 10982 7930
rect 10943 7904 10951 7924
rect 10976 7904 10982 7924
rect 10943 7897 10982 7904
rect 11159 7927 11215 7932
rect 11159 7907 11166 7927
rect 11186 7907 11215 7927
rect 11159 7900 11215 7907
rect 11159 7899 11194 7900
rect 8312 7834 8344 7862
rect 8802 7847 9798 7873
rect 10951 7851 10982 7897
rect 7932 7826 8344 7834
rect 7932 7800 7938 7826
rect 7964 7800 8344 7826
rect 7932 7798 8344 7800
rect 7934 7797 7974 7798
rect 8312 7733 8344 7798
rect 10450 7826 10561 7848
rect 10450 7806 10458 7826
rect 10477 7806 10535 7826
rect 10554 7806 10561 7826
rect 10950 7834 10982 7851
rect 11251 7834 11288 7970
rect 11389 7937 11499 7951
rect 11389 7934 11467 7937
rect 11389 7907 11393 7934
rect 11422 7910 11467 7934
rect 11496 7910 11499 7937
rect 11422 7907 11499 7910
rect 11389 7892 11499 7907
rect 11731 7923 11785 7970
rect 11731 7915 11784 7923
rect 11731 7898 11740 7915
rect 11772 7898 11784 7915
rect 11731 7895 11784 7898
rect 10950 7821 11288 7834
rect 10450 7789 10561 7806
rect 10951 7802 11288 7821
rect 11230 7801 11288 7802
rect 11674 7829 11706 7836
rect 11674 7809 11681 7829
rect 11702 7809 11706 7829
rect 8312 7713 8316 7733
rect 8337 7713 8344 7733
rect 8312 7706 8344 7713
rect 8730 7740 8788 7741
rect 8730 7721 9067 7740
rect 9457 7736 9568 7753
rect 8730 7708 9068 7721
rect 7865 7640 7900 7648
rect 7865 7620 7873 7640
rect 7893 7620 7900 7640
rect 7865 7615 7900 7620
rect 8519 7635 8629 7650
rect 8519 7632 8596 7635
rect 7865 7572 7899 7615
rect 8519 7605 8522 7632
rect 8551 7608 8596 7632
rect 8625 7608 8629 7635
rect 8551 7605 8629 7608
rect 8519 7591 8629 7605
rect 8730 7572 8767 7708
rect 9036 7691 9068 7708
rect 9457 7716 9464 7736
rect 9483 7716 9541 7736
rect 9560 7716 9568 7736
rect 9457 7694 9568 7716
rect 11674 7744 11706 7809
rect 11885 7821 11924 8094
rect 12020 7998 12062 8169
rect 12237 8194 12293 8199
rect 12237 8174 12244 8194
rect 12264 8174 12293 8194
rect 12237 8167 12293 8174
rect 12700 8204 12733 8262
rect 12930 8314 12968 8324
rect 12930 8276 12939 8314
rect 12962 8276 12968 8314
rect 12700 8196 12734 8204
rect 12700 8176 12707 8196
rect 12727 8176 12734 8196
rect 12700 8171 12734 8176
rect 12700 8170 12731 8171
rect 12237 8166 12272 8167
rect 12930 8140 12968 8276
rect 13146 8289 13178 8354
rect 16870 8296 16902 8361
rect 17240 8296 17280 8297
rect 16870 8294 17282 8296
rect 16238 8290 16273 8292
rect 13146 8269 13150 8289
rect 13171 8269 13178 8289
rect 15274 8287 16273 8290
rect 13751 8272 14053 8274
rect 13146 8262 13178 8269
rect 13690 8243 14053 8272
rect 13690 8241 13751 8243
rect 13071 8197 13109 8203
rect 13071 8180 13081 8197
rect 13101 8180 13109 8197
rect 12020 7964 12264 7998
rect 12930 7986 12974 8140
rect 12767 7984 12974 7986
rect 12227 7956 12264 7964
rect 12120 7923 12154 7934
rect 12118 7922 12154 7923
rect 12118 7902 12125 7922
rect 12145 7902 12154 7922
rect 12118 7894 12154 7902
rect 11885 7780 11892 7821
rect 11913 7780 11924 7821
rect 11885 7765 11924 7780
rect 12044 7744 12084 7745
rect 11674 7742 12086 7744
rect 11674 7716 12054 7742
rect 12080 7716 12086 7742
rect 11674 7708 12086 7716
rect 9036 7645 9067 7691
rect 10220 7669 11216 7695
rect 11674 7680 11706 7708
rect 12119 7688 12153 7894
rect 8824 7642 8859 7643
rect 8803 7635 8859 7642
rect 8803 7615 8832 7635
rect 8852 7615 8859 7635
rect 8803 7610 8859 7615
rect 9036 7638 9075 7645
rect 9036 7618 9042 7638
rect 9067 7618 9075 7638
rect 9036 7612 9075 7618
rect 9250 7638 9282 7645
rect 9250 7618 9256 7638
rect 9277 7618 9282 7638
rect 7864 7537 8768 7572
rect 7865 7536 7899 7537
rect 7746 7437 7818 7446
rect 7746 7408 7763 7437
rect 7811 7408 7818 7437
rect 8409 7456 8520 7473
rect 8409 7436 8416 7456
rect 8435 7436 8493 7456
rect 8512 7436 8520 7456
rect 8409 7414 8520 7436
rect 7746 7401 7818 7408
rect 8803 7404 8837 7610
rect 9250 7590 9282 7618
rect 8870 7582 9282 7590
rect 10222 7616 10264 7669
rect 10222 7597 10231 7616
rect 10256 7597 10264 7616
rect 10222 7587 10264 7597
rect 10450 7627 10560 7641
rect 10450 7624 10528 7627
rect 10450 7597 10454 7624
rect 10483 7600 10528 7624
rect 10557 7600 10560 7627
rect 11180 7617 11214 7669
rect 11674 7660 11679 7680
rect 11700 7660 11706 7680
rect 11674 7653 11706 7660
rect 12097 7683 12153 7688
rect 12097 7663 12104 7683
rect 12124 7663 12153 7683
rect 12097 7656 12153 7663
rect 12097 7655 12132 7656
rect 11725 7621 11766 7622
rect 10483 7597 10560 7600
rect 10450 7582 10560 7597
rect 11179 7612 11214 7617
rect 11179 7592 11186 7612
rect 11206 7592 11214 7612
rect 11724 7611 11766 7621
rect 11179 7584 11214 7592
rect 8870 7556 8876 7582
rect 8902 7556 9282 7582
rect 8870 7554 9282 7556
rect 8872 7553 8912 7554
rect 9250 7489 9282 7554
rect 10735 7519 10767 7526
rect 9250 7469 9254 7489
rect 9275 7469 9282 7489
rect 9250 7462 9282 7469
rect 9753 7504 9801 7509
rect 9753 7475 9764 7504
rect 9793 7475 9801 7504
rect 8803 7403 8838 7404
rect 7746 7391 7816 7401
rect 8801 7396 8838 7403
rect 7252 7359 7260 7379
rect 7280 7359 7290 7379
rect 8801 7376 8811 7396
rect 8831 7376 8838 7396
rect 8801 7371 8838 7376
rect 9457 7391 9567 7406
rect 9457 7388 9534 7391
rect 7776 7362 7811 7363
rect 7252 7352 7290 7359
rect 7755 7355 7811 7362
rect 7253 7351 7288 7352
rect 6267 7299 6328 7301
rect 5965 7270 6328 7299
rect 6809 7286 6841 7293
rect 5965 7268 6267 7270
rect 6809 7266 6816 7286
rect 6837 7266 6841 7286
rect 3745 7252 4744 7255
rect 3745 7250 3780 7252
rect 2766 7233 3178 7235
rect 2768 7232 2808 7233
rect 2934 7192 2969 7210
rect 2934 7160 2937 7192
rect 2964 7160 2969 7192
rect 2699 7082 2734 7083
rect 2176 7072 2232 7079
rect 2697 7075 2735 7082
rect 2176 7071 2211 7072
rect 2697 7071 2707 7075
rect 2691 7057 2707 7071
rect 2727 7071 2735 7075
rect 2727 7057 2741 7071
rect 2691 7050 2741 7057
rect 2324 6993 2374 6995
rect 1959 6959 2374 6993
rect 2088 6897 2122 6898
rect 1219 6862 2123 6897
rect 2171 6886 2239 6897
rect 2171 6865 2176 6886
rect 705 6796 710 6816
rect 731 6796 737 6816
rect 705 6789 737 6796
rect 912 6816 951 6822
rect 912 6796 920 6816
rect 945 6796 951 6816
rect 912 6789 951 6796
rect 1128 6819 1184 6824
rect 1128 6799 1135 6819
rect 1155 6799 1184 6819
rect 1128 6792 1184 6799
rect 1128 6791 1163 6792
rect 920 6743 951 6789
rect 419 6718 530 6740
rect 419 6698 427 6718
rect 446 6698 504 6718
rect 523 6698 530 6718
rect 919 6726 951 6743
rect 1220 6726 1257 6862
rect 1358 6829 1468 6843
rect 1358 6826 1436 6829
rect 1358 6799 1362 6826
rect 1391 6802 1436 6826
rect 1465 6802 1468 6829
rect 2088 6819 2122 6862
rect 1391 6799 1468 6802
rect 1358 6784 1468 6799
rect 2087 6814 2122 6819
rect 2087 6794 2094 6814
rect 2114 6794 2122 6814
rect 2087 6786 2122 6794
rect 919 6713 1257 6726
rect 419 6681 530 6698
rect 920 6694 1257 6713
rect 1199 6693 1257 6694
rect 1643 6721 1675 6728
rect 1643 6701 1650 6721
rect 1671 6701 1675 6721
rect 1643 6636 1675 6701
rect 2013 6636 2053 6637
rect 1643 6634 2055 6636
rect 1643 6608 2023 6634
rect 2049 6608 2055 6634
rect 1643 6600 2055 6608
rect 189 6561 1185 6587
rect 1643 6572 1675 6600
rect 191 6508 233 6561
rect 191 6489 200 6508
rect 225 6489 233 6508
rect 191 6479 233 6489
rect 419 6519 529 6533
rect 419 6516 497 6519
rect 419 6489 423 6516
rect 452 6492 497 6516
rect 526 6492 529 6519
rect 1149 6509 1183 6561
rect 1643 6552 1648 6572
rect 1669 6552 1675 6572
rect 1643 6545 1675 6552
rect 1853 6573 1891 6583
rect 2088 6580 2122 6786
rect 1853 6556 1863 6573
rect 1883 6556 1891 6573
rect 1694 6513 1735 6514
rect 452 6489 529 6492
rect 419 6474 529 6489
rect 1148 6504 1183 6509
rect 1148 6484 1155 6504
rect 1175 6484 1183 6504
rect 1693 6503 1735 6513
rect 1148 6476 1183 6484
rect 704 6411 736 6418
rect 704 6391 711 6411
rect 732 6391 736 6411
rect 704 6326 736 6391
rect 1074 6326 1114 6327
rect 704 6324 1116 6326
rect 704 6298 1084 6324
rect 1110 6298 1116 6324
rect 704 6290 1116 6298
rect 704 6262 736 6290
rect 1149 6270 1183 6476
rect 1357 6474 1468 6496
rect 1357 6454 1365 6474
rect 1384 6454 1442 6474
rect 1461 6454 1468 6474
rect 1357 6437 1468 6454
rect 1693 6481 1700 6503
rect 1726 6481 1735 6503
rect 1693 6472 1735 6481
rect 910 6267 953 6269
rect 704 6242 709 6262
rect 730 6242 736 6262
rect 704 6235 736 6242
rect 909 6260 953 6267
rect 909 6240 919 6260
rect 942 6240 953 6260
rect 909 6236 953 6240
rect 1127 6265 1183 6270
rect 1127 6245 1134 6265
rect 1154 6245 1183 6265
rect 1127 6238 1183 6245
rect 1239 6406 1272 6407
rect 1693 6406 1730 6472
rect 1239 6377 1730 6406
rect 1127 6237 1162 6238
rect 418 6164 529 6186
rect 418 6144 426 6164
rect 445 6144 503 6164
rect 522 6144 529 6164
rect 418 6127 529 6144
rect 909 6155 951 6236
rect 1239 6157 1272 6377
rect 1693 6375 1730 6377
rect 1499 6237 1609 6251
rect 1499 6234 1577 6237
rect 1499 6207 1503 6234
rect 1532 6210 1577 6234
rect 1606 6210 1609 6237
rect 1532 6207 1609 6210
rect 1499 6192 1609 6207
rect 1853 6218 1891 6556
rect 2066 6575 2122 6580
rect 2066 6555 2073 6575
rect 2093 6555 2122 6575
rect 2066 6548 2122 6555
rect 2169 6857 2176 6865
rect 2224 6857 2239 6886
rect 2169 6848 2239 6857
rect 2066 6547 2101 6548
rect 1988 6447 2032 6451
rect 2169 6447 2219 6848
rect 2324 6831 2374 6959
rect 2557 6972 2667 6974
rect 2934 6972 2969 7160
rect 3146 7168 3178 7233
rect 6809 7201 6841 7266
rect 7179 7201 7219 7202
rect 6809 7199 7221 7201
rect 6207 7182 6242 7184
rect 5243 7179 6242 7182
rect 3146 7148 3150 7168
rect 3171 7148 3178 7168
rect 3720 7164 4022 7166
rect 3146 7141 3178 7148
rect 3659 7135 4022 7164
rect 3659 7133 3720 7135
rect 2557 6942 2969 6972
rect 2557 6917 2601 6942
rect 2640 6939 2969 6942
rect 3088 7073 3122 7079
rect 3088 7053 3097 7073
rect 3118 7053 3122 7073
rect 1988 6414 2219 6447
rect 1988 6412 2195 6414
rect 1988 6258 2032 6412
rect 1853 6201 1861 6218
rect 1881 6201 1891 6218
rect 1853 6195 1891 6201
rect 1211 6155 1272 6157
rect 909 6126 1272 6155
rect 1784 6129 1816 6136
rect 909 6124 1211 6126
rect 1784 6109 1791 6129
rect 1812 6109 1816 6129
rect 1784 6044 1816 6109
rect 1994 6122 2032 6258
rect 2231 6227 2262 6228
rect 2228 6222 2262 6227
rect 2228 6202 2235 6222
rect 2255 6202 2262 6222
rect 2228 6194 2262 6202
rect 1994 6084 2000 6122
rect 2023 6084 2032 6122
rect 1994 6074 2032 6084
rect 2229 6136 2262 6194
rect 2154 6044 2194 6045
rect 1784 6042 2196 6044
rect 1152 6038 1187 6040
rect 188 6035 1187 6038
rect 187 6011 1187 6035
rect 187 5856 235 6011
rect 421 5970 531 5984
rect 421 5967 499 5970
rect 421 5940 425 5967
rect 454 5943 499 5967
rect 528 5943 531 5970
rect 1152 5960 1187 6011
rect 454 5940 531 5943
rect 421 5925 531 5940
rect 1150 5955 1187 5960
rect 1150 5935 1157 5955
rect 1177 5935 1187 5955
rect 1784 6016 2164 6042
rect 2190 6016 2196 6042
rect 1784 6008 2196 6016
rect 1784 5980 1816 6008
rect 2229 5988 2265 6136
rect 1784 5960 1789 5980
rect 1810 5960 1816 5980
rect 1784 5953 1816 5960
rect 2207 5983 2265 5988
rect 2207 5963 2214 5983
rect 2234 5963 2265 5983
rect 2207 5956 2265 5963
rect 2207 5955 2242 5956
rect 1150 5928 1187 5935
rect 1150 5927 1185 5928
rect 187 5827 195 5856
rect 224 5827 235 5856
rect 187 5822 235 5827
rect 706 5862 738 5869
rect 706 5842 713 5862
rect 734 5842 738 5862
rect 706 5777 738 5842
rect 1076 5777 1116 5778
rect 706 5775 1118 5777
rect 706 5749 1086 5775
rect 1112 5749 1118 5775
rect 706 5741 1118 5749
rect 706 5713 738 5741
rect 1151 5721 1185 5927
rect 1855 5910 1894 5917
rect 1498 5882 1609 5904
rect 1498 5862 1506 5882
rect 1525 5862 1583 5882
rect 1602 5862 1609 5882
rect 1498 5845 1609 5862
rect 1855 5883 1859 5910
rect 1890 5883 1894 5910
rect 1702 5794 1755 5798
rect 1220 5759 1755 5794
rect 706 5693 711 5713
rect 732 5693 738 5713
rect 706 5686 738 5693
rect 913 5713 952 5719
rect 913 5693 921 5713
rect 946 5693 952 5713
rect 913 5686 952 5693
rect 1129 5716 1185 5721
rect 1129 5696 1136 5716
rect 1156 5696 1185 5716
rect 1129 5689 1185 5696
rect 1129 5688 1164 5689
rect 921 5640 952 5686
rect 420 5615 531 5637
rect 420 5595 428 5615
rect 447 5595 505 5615
rect 524 5595 531 5615
rect 920 5623 952 5640
rect 1221 5623 1258 5759
rect 1359 5726 1469 5740
rect 1359 5723 1437 5726
rect 1359 5696 1363 5723
rect 1392 5699 1437 5723
rect 1466 5699 1469 5726
rect 1392 5696 1469 5699
rect 1359 5681 1469 5696
rect 1701 5712 1755 5759
rect 1701 5704 1754 5712
rect 1701 5687 1710 5704
rect 1742 5687 1754 5704
rect 1701 5684 1754 5687
rect 920 5610 1258 5623
rect 420 5578 531 5595
rect 921 5591 1258 5610
rect 1200 5590 1258 5591
rect 1644 5618 1676 5625
rect 1644 5598 1651 5618
rect 1672 5598 1676 5618
rect 1644 5533 1676 5598
rect 1855 5610 1894 5883
rect 2090 5712 2124 5723
rect 2088 5711 2124 5712
rect 2088 5691 2095 5711
rect 2115 5691 2124 5711
rect 2088 5683 2124 5691
rect 1855 5569 1862 5610
rect 1883 5569 1894 5610
rect 1855 5554 1894 5569
rect 2014 5533 2054 5534
rect 1644 5531 2056 5533
rect 1644 5505 2024 5531
rect 2050 5505 2056 5531
rect 1644 5497 2056 5505
rect 190 5458 1186 5484
rect 1644 5469 1676 5497
rect 2089 5477 2123 5683
rect 192 5405 234 5458
rect 192 5386 201 5405
rect 226 5386 234 5405
rect 192 5376 234 5386
rect 420 5416 530 5430
rect 420 5413 498 5416
rect 420 5386 424 5413
rect 453 5389 498 5413
rect 527 5389 530 5416
rect 1150 5406 1184 5458
rect 1644 5449 1649 5469
rect 1670 5449 1676 5469
rect 1644 5442 1676 5449
rect 2067 5472 2123 5477
rect 2067 5452 2074 5472
rect 2094 5452 2123 5472
rect 2067 5445 2123 5452
rect 2067 5444 2102 5445
rect 1695 5410 1736 5411
rect 453 5386 530 5389
rect 420 5371 530 5386
rect 1149 5401 1184 5406
rect 1149 5381 1156 5401
rect 1176 5381 1184 5401
rect 1694 5400 1736 5410
rect 1149 5373 1184 5381
rect 705 5308 737 5315
rect 705 5288 712 5308
rect 733 5288 737 5308
rect 705 5223 737 5288
rect 1075 5223 1115 5224
rect 705 5221 1117 5223
rect 705 5195 1085 5221
rect 1111 5195 1117 5221
rect 705 5187 1117 5195
rect 705 5159 737 5187
rect 1150 5167 1184 5373
rect 1358 5371 1469 5393
rect 1358 5351 1366 5371
rect 1385 5351 1443 5371
rect 1462 5351 1469 5371
rect 1358 5334 1469 5351
rect 1694 5378 1701 5400
rect 1727 5378 1736 5400
rect 1694 5369 1736 5378
rect 911 5164 954 5166
rect 705 5139 710 5159
rect 731 5139 737 5159
rect 705 5132 737 5139
rect 910 5157 954 5164
rect 910 5137 920 5157
rect 943 5137 954 5157
rect 910 5133 954 5137
rect 1128 5162 1184 5167
rect 1128 5142 1135 5162
rect 1155 5142 1184 5162
rect 1128 5135 1184 5142
rect 1240 5303 1273 5304
rect 1694 5303 1731 5369
rect 2326 5346 2372 6831
rect 1240 5274 1731 5303
rect 1128 5134 1163 5135
rect 419 5061 530 5083
rect 419 5041 427 5061
rect 446 5041 504 5061
rect 523 5041 530 5061
rect 419 5024 530 5041
rect 910 5052 952 5133
rect 1240 5054 1273 5274
rect 1694 5272 1731 5274
rect 2324 5322 2372 5346
rect 2554 5340 2601 6917
rect 3088 6874 3122 7053
rect 3353 7070 3463 7085
rect 3353 7067 3430 7070
rect 3353 7040 3356 7067
rect 3385 7043 3430 7067
rect 3459 7043 3463 7070
rect 3385 7040 3463 7043
rect 3353 7026 3463 7040
rect 2697 6849 3122 6874
rect 3201 6913 3238 6915
rect 3659 6913 3692 7133
rect 3980 7054 4022 7135
rect 4402 7146 4513 7162
rect 4402 7126 4409 7146
rect 4428 7126 4486 7146
rect 4505 7126 4513 7146
rect 4402 7104 4513 7126
rect 5242 7155 6242 7179
rect 3769 7052 3804 7053
rect 3201 6884 3692 6913
rect 2697 6833 3121 6849
rect 2697 6442 2735 6833
rect 3201 6818 3238 6884
rect 3659 6883 3692 6884
rect 3748 7045 3804 7052
rect 3748 7025 3777 7045
rect 3797 7025 3804 7045
rect 3748 7020 3804 7025
rect 3978 7050 4022 7054
rect 3978 7030 3989 7050
rect 4012 7030 4022 7050
rect 3978 7023 4022 7030
rect 4195 7048 4227 7055
rect 4195 7028 4201 7048
rect 4222 7028 4227 7048
rect 3978 7021 4021 7023
rect 3196 6809 3238 6818
rect 3196 6787 3205 6809
rect 3231 6787 3238 6809
rect 3463 6836 3574 6853
rect 3463 6816 3470 6836
rect 3489 6816 3547 6836
rect 3566 6816 3574 6836
rect 3463 6794 3574 6816
rect 3748 6814 3782 7020
rect 4195 7000 4227 7028
rect 3815 6992 4227 7000
rect 3815 6966 3821 6992
rect 3847 6966 4227 6992
rect 5242 7000 5290 7155
rect 5476 7114 5586 7128
rect 5476 7111 5554 7114
rect 5476 7084 5480 7111
rect 5509 7087 5554 7111
rect 5583 7087 5586 7114
rect 6207 7104 6242 7155
rect 6809 7173 7189 7199
rect 7215 7173 7221 7199
rect 6809 7165 7221 7173
rect 6809 7137 6841 7165
rect 6809 7117 6814 7137
rect 6835 7117 6841 7137
rect 6809 7110 6841 7117
rect 7015 7136 7060 7148
rect 7254 7145 7288 7351
rect 7015 7117 7022 7136
rect 7051 7117 7060 7136
rect 5509 7084 5586 7087
rect 5476 7069 5586 7084
rect 6205 7099 6242 7104
rect 6205 7079 6212 7099
rect 6232 7079 6242 7099
rect 6205 7072 6242 7079
rect 6205 7071 6240 7072
rect 5242 6971 5250 7000
rect 5279 6971 5290 7000
rect 5242 6966 5290 6971
rect 5761 7006 5793 7013
rect 5761 6986 5768 7006
rect 5789 6986 5793 7006
rect 3815 6964 4227 6966
rect 3817 6963 3857 6964
rect 4195 6899 4227 6964
rect 4195 6879 4199 6899
rect 4220 6879 4227 6899
rect 4195 6872 4227 6879
rect 5761 6921 5793 6986
rect 6131 6921 6171 6922
rect 5761 6919 6173 6921
rect 5761 6893 6141 6919
rect 6167 6893 6173 6919
rect 5761 6885 6173 6893
rect 5761 6857 5793 6885
rect 6206 6865 6240 7071
rect 6523 7039 6634 7061
rect 6523 7019 6531 7039
rect 6550 7019 6608 7039
rect 6627 7019 6634 7039
rect 6523 7002 6634 7019
rect 7015 7034 7060 7117
rect 7232 7140 7288 7145
rect 7232 7120 7239 7140
rect 7259 7120 7288 7140
rect 7755 7335 7784 7355
rect 7804 7335 7811 7355
rect 7755 7330 7811 7335
rect 8202 7358 8234 7365
rect 8202 7338 8208 7358
rect 8229 7338 8234 7358
rect 7755 7124 7789 7330
rect 8202 7310 8234 7338
rect 7822 7302 8234 7310
rect 7822 7276 7828 7302
rect 7854 7276 8234 7302
rect 8801 7320 8836 7371
rect 9457 7361 9460 7388
rect 9489 7364 9534 7388
rect 9563 7364 9567 7391
rect 9489 7361 9567 7364
rect 9457 7347 9567 7361
rect 9753 7320 9801 7475
rect 10735 7499 10742 7519
rect 10763 7499 10767 7519
rect 10735 7434 10767 7499
rect 11105 7434 11145 7435
rect 10735 7432 11147 7434
rect 10735 7406 11115 7432
rect 11141 7406 11147 7432
rect 10735 7398 11147 7406
rect 10735 7370 10767 7398
rect 11180 7378 11214 7584
rect 11388 7582 11499 7604
rect 11388 7562 11396 7582
rect 11415 7562 11473 7582
rect 11492 7562 11499 7582
rect 11388 7545 11499 7562
rect 11724 7589 11731 7611
rect 11757 7589 11766 7611
rect 11724 7580 11766 7589
rect 10941 7375 10984 7377
rect 10735 7350 10740 7370
rect 10761 7350 10767 7370
rect 10735 7343 10767 7350
rect 10940 7368 10984 7375
rect 10940 7348 10950 7368
rect 10973 7348 10984 7368
rect 10940 7344 10984 7348
rect 11158 7373 11214 7378
rect 11158 7353 11165 7373
rect 11185 7353 11214 7373
rect 11158 7346 11214 7353
rect 11270 7514 11303 7515
rect 11724 7514 11761 7580
rect 11270 7485 11761 7514
rect 11158 7345 11193 7346
rect 8801 7296 9801 7320
rect 8801 7293 9800 7296
rect 8801 7291 8836 7293
rect 7822 7274 8234 7276
rect 7824 7273 7864 7274
rect 7990 7233 8025 7251
rect 7990 7201 7993 7233
rect 8020 7201 8025 7233
rect 7755 7123 7790 7124
rect 7232 7113 7288 7120
rect 7753 7116 7791 7123
rect 7232 7112 7267 7113
rect 7753 7112 7763 7116
rect 7747 7098 7763 7112
rect 7783 7112 7791 7116
rect 7783 7098 7797 7112
rect 7747 7091 7797 7098
rect 7380 7034 7430 7036
rect 7015 7000 7430 7034
rect 7144 6938 7178 6939
rect 6275 6903 7179 6938
rect 7227 6927 7295 6938
rect 7227 6906 7232 6927
rect 5761 6837 5766 6857
rect 5787 6837 5793 6857
rect 5761 6830 5793 6837
rect 5968 6857 6007 6863
rect 5968 6837 5976 6857
rect 6001 6837 6007 6857
rect 5968 6830 6007 6837
rect 6184 6860 6240 6865
rect 6184 6840 6191 6860
rect 6211 6840 6240 6860
rect 6184 6833 6240 6840
rect 6184 6832 6219 6833
rect 3748 6806 3783 6814
rect 3196 6777 3238 6787
rect 3748 6786 3756 6806
rect 3776 6786 3783 6806
rect 3748 6781 3783 6786
rect 4402 6801 4512 6816
rect 4402 6798 4479 6801
rect 3196 6776 3237 6777
rect 2830 6742 2865 6743
rect 2809 6735 2865 6742
rect 2809 6715 2838 6735
rect 2858 6715 2865 6735
rect 2809 6710 2865 6715
rect 3256 6738 3288 6745
rect 3256 6718 3262 6738
rect 3283 6718 3288 6738
rect 3748 6729 3782 6781
rect 4402 6771 4405 6798
rect 4434 6774 4479 6798
rect 4508 6774 4512 6801
rect 4434 6771 4512 6774
rect 4402 6757 4512 6771
rect 4698 6801 4740 6811
rect 4698 6782 4706 6801
rect 4731 6782 4740 6801
rect 5976 6784 6007 6830
rect 4698 6729 4740 6782
rect 5475 6759 5586 6781
rect 5475 6739 5483 6759
rect 5502 6739 5560 6759
rect 5579 6739 5586 6759
rect 5975 6767 6007 6784
rect 6276 6767 6313 6903
rect 6414 6870 6524 6884
rect 6414 6867 6492 6870
rect 6414 6840 6418 6867
rect 6447 6843 6492 6867
rect 6521 6843 6524 6870
rect 7144 6860 7178 6903
rect 6447 6840 6524 6843
rect 6414 6825 6524 6840
rect 7143 6855 7178 6860
rect 7143 6835 7150 6855
rect 7170 6835 7178 6855
rect 7143 6827 7178 6835
rect 5975 6754 6313 6767
rect 2809 6504 2843 6710
rect 3256 6690 3288 6718
rect 3746 6703 4742 6729
rect 5475 6722 5586 6739
rect 5976 6735 6313 6754
rect 6255 6734 6313 6735
rect 6699 6762 6731 6769
rect 6699 6742 6706 6762
rect 6727 6742 6731 6762
rect 2876 6682 3288 6690
rect 2876 6656 2882 6682
rect 2908 6656 3288 6682
rect 2876 6654 3288 6656
rect 2878 6653 2918 6654
rect 3038 6618 3077 6633
rect 3038 6577 3049 6618
rect 3070 6577 3077 6618
rect 2808 6496 2844 6504
rect 2808 6476 2817 6496
rect 2837 6476 2844 6496
rect 2808 6475 2844 6476
rect 2808 6464 2842 6475
rect 2698 6434 2735 6442
rect 2698 6400 2942 6434
rect 2690 6231 2725 6232
rect 2669 6224 2725 6231
rect 2669 6204 2698 6224
rect 2718 6204 2725 6224
rect 2669 6199 2725 6204
rect 2900 6229 2942 6400
rect 3038 6304 3077 6577
rect 3256 6589 3288 6654
rect 6699 6677 6731 6742
rect 7069 6677 7109 6678
rect 6699 6675 7111 6677
rect 6699 6649 7079 6675
rect 7105 6649 7111 6675
rect 6699 6641 7111 6649
rect 3256 6569 3260 6589
rect 3281 6569 3288 6589
rect 3256 6562 3288 6569
rect 3674 6596 3732 6597
rect 3674 6577 4011 6596
rect 4401 6592 4512 6609
rect 5245 6602 6241 6628
rect 6699 6613 6731 6641
rect 3674 6564 4012 6577
rect 3178 6500 3231 6503
rect 3178 6483 3190 6500
rect 3222 6483 3231 6500
rect 3178 6475 3231 6483
rect 3177 6428 3231 6475
rect 3463 6491 3573 6506
rect 3463 6488 3540 6491
rect 3463 6461 3466 6488
rect 3495 6464 3540 6488
rect 3569 6464 3573 6491
rect 3495 6461 3573 6464
rect 3463 6447 3573 6461
rect 3674 6428 3711 6564
rect 3980 6547 4012 6564
rect 4401 6572 4408 6592
rect 4427 6572 4485 6592
rect 4504 6572 4512 6592
rect 4401 6550 4512 6572
rect 5247 6549 5289 6602
rect 3980 6501 4011 6547
rect 5247 6530 5256 6549
rect 5281 6530 5289 6549
rect 5247 6520 5289 6530
rect 5475 6560 5585 6574
rect 5475 6557 5553 6560
rect 5475 6530 5479 6557
rect 5508 6533 5553 6557
rect 5582 6533 5585 6560
rect 6205 6550 6239 6602
rect 6699 6593 6704 6613
rect 6725 6593 6731 6613
rect 6699 6586 6731 6593
rect 6909 6614 6947 6624
rect 7144 6621 7178 6827
rect 6909 6597 6919 6614
rect 6939 6597 6947 6614
rect 6750 6554 6791 6555
rect 5508 6530 5585 6533
rect 5475 6515 5585 6530
rect 6204 6545 6239 6550
rect 6204 6525 6211 6545
rect 6231 6525 6239 6545
rect 6749 6544 6791 6554
rect 6204 6517 6239 6525
rect 3768 6498 3803 6499
rect 3747 6491 3803 6498
rect 3747 6471 3776 6491
rect 3796 6471 3803 6491
rect 3747 6466 3803 6471
rect 3980 6494 4019 6501
rect 3980 6474 3986 6494
rect 4011 6474 4019 6494
rect 3980 6468 4019 6474
rect 4194 6494 4226 6501
rect 4194 6474 4200 6494
rect 4221 6474 4226 6494
rect 3177 6393 3712 6428
rect 3177 6389 3230 6393
rect 3038 6277 3042 6304
rect 3073 6277 3077 6304
rect 3323 6325 3434 6342
rect 3323 6305 3330 6325
rect 3349 6305 3407 6325
rect 3426 6305 3434 6325
rect 3323 6283 3434 6305
rect 3038 6270 3077 6277
rect 3747 6260 3781 6466
rect 4194 6446 4226 6474
rect 3814 6438 4226 6446
rect 3814 6412 3820 6438
rect 3846 6412 4226 6438
rect 3814 6410 4226 6412
rect 3816 6409 3856 6410
rect 4194 6345 4226 6410
rect 5760 6452 5792 6459
rect 5760 6432 5767 6452
rect 5788 6432 5792 6452
rect 5760 6367 5792 6432
rect 6130 6367 6170 6368
rect 5760 6365 6172 6367
rect 4194 6325 4198 6345
rect 4219 6325 4226 6345
rect 4194 6318 4226 6325
rect 4697 6360 4745 6365
rect 4697 6331 4708 6360
rect 4737 6331 4745 6360
rect 3747 6259 3782 6260
rect 3745 6252 3782 6259
rect 2900 6208 2908 6229
rect 2935 6208 2942 6229
rect 2669 5993 2703 6199
rect 2900 6197 2942 6208
rect 3116 6227 3148 6234
rect 3116 6207 3122 6227
rect 3143 6207 3148 6227
rect 3116 6179 3148 6207
rect 2736 6171 3148 6179
rect 2736 6145 2742 6171
rect 2768 6145 3148 6171
rect 3745 6232 3755 6252
rect 3775 6232 3782 6252
rect 3745 6227 3782 6232
rect 4401 6247 4511 6262
rect 4401 6244 4478 6247
rect 3745 6176 3780 6227
rect 4401 6217 4404 6244
rect 4433 6220 4478 6244
rect 4507 6220 4511 6247
rect 4433 6217 4511 6220
rect 4401 6203 4511 6217
rect 4697 6176 4745 6331
rect 5760 6339 6140 6365
rect 6166 6339 6172 6365
rect 5760 6331 6172 6339
rect 5760 6303 5792 6331
rect 6205 6311 6239 6517
rect 6413 6515 6524 6537
rect 6413 6495 6421 6515
rect 6440 6495 6498 6515
rect 6517 6495 6524 6515
rect 6413 6478 6524 6495
rect 6749 6522 6756 6544
rect 6782 6522 6791 6544
rect 6749 6513 6791 6522
rect 5966 6308 6009 6310
rect 5760 6283 5765 6303
rect 5786 6283 5792 6303
rect 5760 6276 5792 6283
rect 5965 6301 6009 6308
rect 5965 6281 5975 6301
rect 5998 6281 6009 6301
rect 5965 6277 6009 6281
rect 6183 6306 6239 6311
rect 6183 6286 6190 6306
rect 6210 6286 6239 6306
rect 6183 6279 6239 6286
rect 6295 6447 6328 6448
rect 6749 6447 6786 6513
rect 6295 6418 6786 6447
rect 6183 6278 6218 6279
rect 3745 6152 4745 6176
rect 5474 6205 5585 6227
rect 5474 6185 5482 6205
rect 5501 6185 5559 6205
rect 5578 6185 5585 6205
rect 5474 6168 5585 6185
rect 5965 6196 6007 6277
rect 6295 6198 6328 6418
rect 6749 6416 6786 6418
rect 6555 6278 6665 6292
rect 6555 6275 6633 6278
rect 6555 6248 6559 6275
rect 6588 6251 6633 6275
rect 6662 6251 6665 6278
rect 6588 6248 6665 6251
rect 6555 6233 6665 6248
rect 6909 6259 6947 6597
rect 7122 6616 7178 6621
rect 7122 6596 7129 6616
rect 7149 6596 7178 6616
rect 7122 6589 7178 6596
rect 7225 6898 7232 6906
rect 7280 6898 7295 6927
rect 7225 6889 7295 6898
rect 7122 6588 7157 6589
rect 7044 6488 7088 6492
rect 7225 6488 7275 6889
rect 7380 6872 7430 7000
rect 7613 7013 7723 7015
rect 7990 7013 8025 7201
rect 8202 7209 8234 7274
rect 10449 7272 10560 7294
rect 10449 7252 10457 7272
rect 10476 7252 10534 7272
rect 10553 7252 10560 7272
rect 10449 7236 10560 7252
rect 10940 7263 10982 7344
rect 11270 7265 11303 7485
rect 11724 7483 11761 7485
rect 11499 7358 11609 7372
rect 11499 7355 11577 7358
rect 11499 7328 11503 7355
rect 11532 7331 11577 7355
rect 11606 7331 11609 7358
rect 11532 7328 11609 7331
rect 11499 7313 11609 7328
rect 12227 7343 12265 7956
rect 12743 7951 12974 7984
rect 12743 7410 12793 7951
rect 12930 7947 12974 7951
rect 12861 7850 12896 7851
rect 12840 7843 12896 7850
rect 12840 7823 12869 7843
rect 12889 7823 12896 7843
rect 12840 7818 12896 7823
rect 13071 7842 13109 8180
rect 13353 8191 13463 8206
rect 13353 8188 13430 8191
rect 13353 8161 13356 8188
rect 13385 8164 13430 8188
rect 13459 8164 13463 8191
rect 13385 8161 13463 8164
rect 13353 8147 13463 8161
rect 13232 8021 13269 8023
rect 13690 8021 13723 8241
rect 14011 8162 14053 8243
rect 14433 8254 14544 8271
rect 14433 8234 14440 8254
rect 14459 8234 14517 8254
rect 14536 8234 14544 8254
rect 14433 8212 14544 8234
rect 15273 8263 16273 8287
rect 13800 8160 13835 8161
rect 13232 7992 13723 8021
rect 13232 7926 13269 7992
rect 13690 7991 13723 7992
rect 13779 8153 13835 8160
rect 13779 8133 13808 8153
rect 13828 8133 13835 8153
rect 13779 8128 13835 8133
rect 14009 8158 14053 8162
rect 14009 8138 14020 8158
rect 14043 8138 14053 8158
rect 14009 8131 14053 8138
rect 14226 8156 14258 8163
rect 14226 8136 14232 8156
rect 14253 8136 14258 8156
rect 14009 8129 14052 8131
rect 13227 7917 13269 7926
rect 13227 7895 13236 7917
rect 13262 7895 13269 7917
rect 13494 7944 13605 7961
rect 13494 7924 13501 7944
rect 13520 7924 13578 7944
rect 13597 7924 13605 7944
rect 13494 7902 13605 7924
rect 13779 7922 13813 8128
rect 14226 8108 14258 8136
rect 13846 8100 14258 8108
rect 13846 8074 13852 8100
rect 13878 8074 14258 8100
rect 15273 8108 15321 8263
rect 15507 8222 15617 8236
rect 15507 8219 15585 8222
rect 15507 8192 15511 8219
rect 15540 8195 15585 8219
rect 15614 8195 15617 8222
rect 16238 8212 16273 8263
rect 15540 8192 15617 8195
rect 15507 8177 15617 8192
rect 16236 8207 16273 8212
rect 16236 8187 16243 8207
rect 16263 8187 16273 8207
rect 16870 8268 17250 8294
rect 17276 8268 17282 8294
rect 16870 8260 17282 8268
rect 16870 8232 16902 8260
rect 16870 8212 16875 8232
rect 16896 8212 16902 8232
rect 16870 8205 16902 8212
rect 17076 8231 17118 8242
rect 17315 8240 17349 8446
rect 17753 8476 17811 8483
rect 17753 8456 17784 8476
rect 17804 8456 17811 8476
rect 17753 8451 17811 8456
rect 18202 8479 18234 8486
rect 18202 8459 18208 8479
rect 18229 8459 18234 8479
rect 17753 8303 17789 8451
rect 18202 8431 18234 8459
rect 17822 8423 18234 8431
rect 17822 8397 17828 8423
rect 17854 8397 18234 8423
rect 18831 8484 18841 8504
rect 18861 8484 18868 8504
rect 18831 8479 18868 8484
rect 19487 8499 19597 8514
rect 19487 8496 19564 8499
rect 18831 8428 18866 8479
rect 19487 8469 19490 8496
rect 19519 8472 19564 8496
rect 19593 8472 19597 8499
rect 19519 8469 19597 8472
rect 19487 8455 19597 8469
rect 19783 8428 19831 8583
rect 18831 8404 19831 8428
rect 18831 8401 19830 8404
rect 18831 8399 18866 8401
rect 17822 8395 18234 8397
rect 17824 8394 17864 8395
rect 17076 8210 17083 8231
rect 17110 8210 17118 8231
rect 16236 8180 16273 8187
rect 16236 8179 16271 8180
rect 15273 8079 15281 8108
rect 15310 8079 15321 8108
rect 15273 8074 15321 8079
rect 15792 8114 15824 8121
rect 15792 8094 15799 8114
rect 15820 8094 15824 8114
rect 13846 8072 14258 8074
rect 13848 8071 13888 8072
rect 14226 8007 14258 8072
rect 14226 7987 14230 8007
rect 14251 7987 14258 8007
rect 14226 7980 14258 7987
rect 15792 8029 15824 8094
rect 16162 8029 16202 8030
rect 15792 8027 16204 8029
rect 15792 8001 16172 8027
rect 16198 8001 16204 8027
rect 15792 7993 16204 8001
rect 15792 7965 15824 7993
rect 16237 7973 16271 8179
rect 16941 8162 16980 8169
rect 16584 8134 16695 8156
rect 16584 8114 16592 8134
rect 16611 8114 16669 8134
rect 16688 8114 16695 8134
rect 16584 8097 16695 8114
rect 16941 8135 16945 8162
rect 16976 8135 16980 8162
rect 16788 8046 16841 8050
rect 16306 8011 16841 8046
rect 15792 7945 15797 7965
rect 15818 7945 15824 7965
rect 15792 7938 15824 7945
rect 15999 7965 16038 7971
rect 15999 7945 16007 7965
rect 16032 7945 16038 7965
rect 15999 7938 16038 7945
rect 16215 7968 16271 7973
rect 16215 7948 16222 7968
rect 16242 7948 16271 7968
rect 16215 7941 16271 7948
rect 16215 7940 16250 7941
rect 13779 7914 13814 7922
rect 13227 7885 13269 7895
rect 13779 7894 13787 7914
rect 13807 7894 13814 7914
rect 13779 7889 13814 7894
rect 14433 7909 14543 7924
rect 14433 7906 14510 7909
rect 13227 7884 13268 7885
rect 13071 7825 13079 7842
rect 13099 7825 13109 7842
rect 12840 7612 12874 7818
rect 13071 7815 13109 7825
rect 13287 7846 13319 7853
rect 13287 7826 13293 7846
rect 13314 7826 13319 7846
rect 13779 7837 13813 7889
rect 14433 7879 14436 7906
rect 14465 7882 14510 7906
rect 14539 7882 14543 7909
rect 14465 7879 14543 7882
rect 14433 7865 14543 7879
rect 14729 7909 14771 7919
rect 14729 7890 14737 7909
rect 14762 7890 14771 7909
rect 16007 7892 16038 7938
rect 14729 7837 14771 7890
rect 15506 7867 15617 7889
rect 15506 7847 15514 7867
rect 15533 7847 15591 7867
rect 15610 7847 15617 7867
rect 16006 7875 16038 7892
rect 16307 7875 16344 8011
rect 16445 7978 16555 7992
rect 16445 7975 16523 7978
rect 16445 7948 16449 7975
rect 16478 7951 16523 7975
rect 16552 7951 16555 7978
rect 16478 7948 16555 7951
rect 16445 7933 16555 7948
rect 16787 7964 16841 8011
rect 16787 7956 16840 7964
rect 16787 7939 16796 7956
rect 16828 7939 16840 7956
rect 16787 7936 16840 7939
rect 16006 7862 16344 7875
rect 13287 7798 13319 7826
rect 13777 7811 14773 7837
rect 15506 7830 15617 7847
rect 16007 7843 16344 7862
rect 16286 7842 16344 7843
rect 16730 7870 16762 7877
rect 16730 7850 16737 7870
rect 16758 7850 16762 7870
rect 12907 7790 13319 7798
rect 12907 7764 12913 7790
rect 12939 7764 13319 7790
rect 12907 7762 13319 7764
rect 12909 7761 12949 7762
rect 13287 7697 13319 7762
rect 16730 7785 16762 7850
rect 16941 7862 16980 8135
rect 17076 8039 17118 8210
rect 17293 8235 17349 8240
rect 17293 8215 17300 8235
rect 17320 8215 17349 8235
rect 17293 8208 17349 8215
rect 17756 8245 17789 8303
rect 17986 8355 18024 8365
rect 17986 8317 17995 8355
rect 18018 8317 18024 8355
rect 17756 8237 17790 8245
rect 17756 8217 17763 8237
rect 17783 8217 17790 8237
rect 17756 8212 17790 8217
rect 17756 8211 17787 8212
rect 17293 8207 17328 8208
rect 17986 8181 18024 8317
rect 18202 8330 18234 8395
rect 18202 8310 18206 8330
rect 18227 8310 18234 8330
rect 18807 8313 19109 8315
rect 18202 8303 18234 8310
rect 18746 8284 19109 8313
rect 18746 8282 18807 8284
rect 18127 8238 18165 8244
rect 18127 8221 18137 8238
rect 18157 8221 18165 8238
rect 17076 8005 17320 8039
rect 17986 8027 18030 8181
rect 17823 8025 18030 8027
rect 17283 7997 17320 8005
rect 17176 7964 17210 7975
rect 17174 7963 17210 7964
rect 17174 7943 17181 7963
rect 17201 7943 17210 7963
rect 17174 7935 17210 7943
rect 16941 7821 16948 7862
rect 16969 7821 16980 7862
rect 16941 7806 16980 7821
rect 17100 7785 17140 7786
rect 16730 7783 17142 7785
rect 16730 7757 17110 7783
rect 17136 7757 17142 7783
rect 16730 7749 17142 7757
rect 13287 7677 13291 7697
rect 13312 7677 13319 7697
rect 13287 7670 13319 7677
rect 13705 7704 13763 7705
rect 13705 7685 14042 7704
rect 14432 7700 14543 7717
rect 15276 7710 16272 7736
rect 16730 7721 16762 7749
rect 17175 7729 17209 7935
rect 13705 7672 14043 7685
rect 12840 7604 12875 7612
rect 12840 7584 12848 7604
rect 12868 7584 12875 7604
rect 12840 7579 12875 7584
rect 13494 7599 13604 7614
rect 13494 7596 13571 7599
rect 12840 7536 12874 7579
rect 13494 7569 13497 7596
rect 13526 7572 13571 7596
rect 13600 7572 13604 7599
rect 13526 7569 13604 7572
rect 13494 7555 13604 7569
rect 13705 7536 13742 7672
rect 14011 7655 14043 7672
rect 14432 7680 14439 7700
rect 14458 7680 14516 7700
rect 14535 7680 14543 7700
rect 14432 7658 14543 7680
rect 15278 7657 15320 7710
rect 14011 7609 14042 7655
rect 15278 7638 15287 7657
rect 15312 7638 15320 7657
rect 15278 7628 15320 7638
rect 15506 7668 15616 7682
rect 15506 7665 15584 7668
rect 15506 7638 15510 7665
rect 15539 7641 15584 7665
rect 15613 7641 15616 7668
rect 16236 7658 16270 7710
rect 16730 7701 16735 7721
rect 16756 7701 16762 7721
rect 16730 7694 16762 7701
rect 17153 7724 17209 7729
rect 17153 7704 17160 7724
rect 17180 7704 17209 7724
rect 17153 7697 17209 7704
rect 17153 7696 17188 7697
rect 16781 7662 16822 7663
rect 15539 7638 15616 7641
rect 15506 7623 15616 7638
rect 16235 7653 16270 7658
rect 16235 7633 16242 7653
rect 16262 7633 16270 7653
rect 16780 7652 16822 7662
rect 16235 7625 16270 7633
rect 13799 7606 13834 7607
rect 13778 7599 13834 7606
rect 13778 7579 13807 7599
rect 13827 7579 13834 7599
rect 13778 7574 13834 7579
rect 14011 7602 14050 7609
rect 14011 7582 14017 7602
rect 14042 7582 14050 7602
rect 14011 7576 14050 7582
rect 14225 7602 14257 7609
rect 14225 7582 14231 7602
rect 14252 7582 14257 7602
rect 12839 7501 13743 7536
rect 12840 7500 12874 7501
rect 12721 7401 12793 7410
rect 12721 7372 12738 7401
rect 12786 7372 12793 7401
rect 13384 7420 13495 7437
rect 13384 7400 13391 7420
rect 13410 7400 13468 7420
rect 13487 7400 13495 7420
rect 13384 7378 13495 7400
rect 12721 7365 12793 7372
rect 13778 7368 13812 7574
rect 14225 7554 14257 7582
rect 13845 7546 14257 7554
rect 13845 7520 13851 7546
rect 13877 7520 14257 7546
rect 13845 7518 14257 7520
rect 13847 7517 13887 7518
rect 14225 7453 14257 7518
rect 15791 7560 15823 7567
rect 15791 7540 15798 7560
rect 15819 7540 15823 7560
rect 15791 7475 15823 7540
rect 16161 7475 16201 7476
rect 15791 7473 16203 7475
rect 14225 7433 14229 7453
rect 14250 7433 14257 7453
rect 14225 7426 14257 7433
rect 14728 7468 14776 7473
rect 14728 7439 14739 7468
rect 14768 7439 14776 7468
rect 13778 7367 13813 7368
rect 12721 7355 12791 7365
rect 13776 7360 13813 7367
rect 12227 7323 12235 7343
rect 12255 7323 12265 7343
rect 13776 7340 13786 7360
rect 13806 7340 13813 7360
rect 13776 7335 13813 7340
rect 14432 7355 14542 7370
rect 14432 7352 14509 7355
rect 12751 7326 12786 7327
rect 12227 7316 12265 7323
rect 12730 7319 12786 7326
rect 12228 7315 12263 7316
rect 11242 7263 11303 7265
rect 10940 7234 11303 7263
rect 11784 7250 11816 7257
rect 10940 7232 11242 7234
rect 8202 7189 8206 7209
rect 8227 7189 8234 7209
rect 11784 7230 11791 7250
rect 11812 7230 11816 7250
rect 8776 7205 9078 7207
rect 8202 7182 8234 7189
rect 8715 7176 9078 7205
rect 8715 7174 8776 7176
rect 7613 6983 8025 7013
rect 7613 6958 7657 6983
rect 7696 6980 8025 6983
rect 8144 7114 8178 7120
rect 8144 7094 8153 7114
rect 8174 7094 8178 7114
rect 7044 6455 7275 6488
rect 7044 6453 7251 6455
rect 7044 6299 7088 6453
rect 6909 6242 6917 6259
rect 6937 6242 6947 6259
rect 6909 6236 6947 6242
rect 6267 6196 6328 6198
rect 5965 6167 6328 6196
rect 6840 6170 6872 6177
rect 5965 6165 6267 6167
rect 3745 6149 4744 6152
rect 6840 6150 6847 6170
rect 6868 6150 6872 6170
rect 3745 6147 3780 6149
rect 2736 6143 3148 6145
rect 2738 6142 2778 6143
rect 3116 6078 3148 6143
rect 6840 6085 6872 6150
rect 7050 6163 7088 6299
rect 7287 6268 7318 6269
rect 7284 6263 7318 6268
rect 7284 6243 7291 6263
rect 7311 6243 7318 6263
rect 7284 6235 7318 6243
rect 7050 6125 7056 6163
rect 7079 6125 7088 6163
rect 7050 6115 7088 6125
rect 7285 6177 7318 6235
rect 7210 6085 7250 6086
rect 6840 6083 7252 6085
rect 6208 6079 6243 6081
rect 3116 6058 3120 6078
rect 3141 6058 3148 6078
rect 5244 6076 6243 6079
rect 3721 6061 4023 6063
rect 3116 6051 3148 6058
rect 3660 6032 4023 6061
rect 3660 6030 3721 6032
rect 2669 5985 2704 5993
rect 2669 5965 2677 5985
rect 2697 5965 2704 5985
rect 2669 5960 2704 5965
rect 3041 5986 3079 5992
rect 3041 5969 3051 5986
rect 3071 5969 3079 5986
rect 2669 5959 2701 5960
rect 2831 5639 2866 5640
rect 1468 5153 1578 5167
rect 1468 5150 1546 5153
rect 1468 5123 1472 5150
rect 1501 5126 1546 5150
rect 1575 5126 1578 5153
rect 2324 5144 2371 5322
rect 2554 5300 2567 5340
rect 2594 5300 2601 5340
rect 2810 5632 2866 5639
rect 2810 5612 2839 5632
rect 2859 5612 2866 5632
rect 2810 5607 2866 5612
rect 3041 5631 3079 5969
rect 3323 5980 3433 5995
rect 3323 5977 3400 5980
rect 3323 5950 3326 5977
rect 3355 5953 3400 5977
rect 3429 5953 3433 5980
rect 3355 5950 3433 5953
rect 3323 5936 3433 5950
rect 3202 5810 3239 5812
rect 3660 5810 3693 6030
rect 3981 5951 4023 6032
rect 4403 6043 4514 6060
rect 4403 6023 4410 6043
rect 4429 6023 4487 6043
rect 4506 6023 4514 6043
rect 4403 6001 4514 6023
rect 5243 6052 6243 6076
rect 3770 5949 3805 5950
rect 3202 5781 3693 5810
rect 3202 5715 3239 5781
rect 3660 5780 3693 5781
rect 3749 5942 3805 5949
rect 3749 5922 3778 5942
rect 3798 5922 3805 5942
rect 3749 5917 3805 5922
rect 3979 5947 4023 5951
rect 3979 5927 3990 5947
rect 4013 5927 4023 5947
rect 3979 5920 4023 5927
rect 4196 5945 4228 5952
rect 4196 5925 4202 5945
rect 4223 5925 4228 5945
rect 3979 5918 4022 5920
rect 3197 5706 3239 5715
rect 3197 5684 3206 5706
rect 3232 5684 3239 5706
rect 3464 5733 3575 5750
rect 3464 5713 3471 5733
rect 3490 5713 3548 5733
rect 3567 5713 3575 5733
rect 3464 5691 3575 5713
rect 3749 5711 3783 5917
rect 4196 5897 4228 5925
rect 3816 5889 4228 5897
rect 3816 5863 3822 5889
rect 3848 5863 4228 5889
rect 5243 5897 5291 6052
rect 5477 6011 5587 6025
rect 5477 6008 5555 6011
rect 5477 5981 5481 6008
rect 5510 5984 5555 6008
rect 5584 5984 5587 6011
rect 6208 6001 6243 6052
rect 5510 5981 5587 5984
rect 5477 5966 5587 5981
rect 6206 5996 6243 6001
rect 6206 5976 6213 5996
rect 6233 5976 6243 5996
rect 6840 6057 7220 6083
rect 7246 6057 7252 6083
rect 6840 6049 7252 6057
rect 6840 6021 6872 6049
rect 7285 6029 7321 6177
rect 6840 6001 6845 6021
rect 6866 6001 6872 6021
rect 6840 5994 6872 6001
rect 7263 6024 7321 6029
rect 7263 6004 7270 6024
rect 7290 6004 7321 6024
rect 7263 5997 7321 6004
rect 7263 5996 7298 5997
rect 6206 5969 6243 5976
rect 6206 5968 6241 5969
rect 5243 5868 5251 5897
rect 5280 5868 5291 5897
rect 5243 5863 5291 5868
rect 5762 5903 5794 5910
rect 5762 5883 5769 5903
rect 5790 5883 5794 5903
rect 3816 5861 4228 5863
rect 3818 5860 3858 5861
rect 4196 5796 4228 5861
rect 4196 5776 4200 5796
rect 4221 5776 4228 5796
rect 4196 5769 4228 5776
rect 5762 5818 5794 5883
rect 6132 5818 6172 5819
rect 5762 5816 6174 5818
rect 5762 5790 6142 5816
rect 6168 5790 6174 5816
rect 5762 5782 6174 5790
rect 5762 5754 5794 5782
rect 6207 5762 6241 5968
rect 6911 5951 6950 5958
rect 6554 5923 6665 5945
rect 6554 5903 6562 5923
rect 6581 5903 6639 5923
rect 6658 5903 6665 5923
rect 6554 5886 6665 5903
rect 6911 5924 6915 5951
rect 6946 5924 6950 5951
rect 6758 5835 6811 5839
rect 6276 5800 6811 5835
rect 5762 5734 5767 5754
rect 5788 5734 5794 5754
rect 5762 5727 5794 5734
rect 5969 5754 6008 5760
rect 5969 5734 5977 5754
rect 6002 5734 6008 5754
rect 5969 5727 6008 5734
rect 6185 5757 6241 5762
rect 6185 5737 6192 5757
rect 6212 5737 6241 5757
rect 6185 5730 6241 5737
rect 6185 5729 6220 5730
rect 3749 5703 3784 5711
rect 3197 5674 3239 5684
rect 3749 5683 3757 5703
rect 3777 5683 3784 5703
rect 3749 5678 3784 5683
rect 4403 5698 4513 5713
rect 4403 5695 4480 5698
rect 3197 5673 3238 5674
rect 3041 5614 3049 5631
rect 3069 5614 3079 5631
rect 2810 5401 2844 5607
rect 3041 5604 3079 5614
rect 3257 5635 3289 5642
rect 3257 5615 3263 5635
rect 3284 5615 3289 5635
rect 3749 5626 3783 5678
rect 4403 5668 4406 5695
rect 4435 5671 4480 5695
rect 4509 5671 4513 5698
rect 4435 5668 4513 5671
rect 4403 5654 4513 5668
rect 4699 5698 4741 5708
rect 4699 5679 4707 5698
rect 4732 5679 4741 5698
rect 5977 5681 6008 5727
rect 4699 5626 4741 5679
rect 5476 5656 5587 5678
rect 5476 5636 5484 5656
rect 5503 5636 5561 5656
rect 5580 5636 5587 5656
rect 5976 5664 6008 5681
rect 6277 5664 6314 5800
rect 6415 5767 6525 5781
rect 6415 5764 6493 5767
rect 6415 5737 6419 5764
rect 6448 5740 6493 5764
rect 6522 5740 6525 5767
rect 6448 5737 6525 5740
rect 6415 5722 6525 5737
rect 6757 5753 6811 5800
rect 6757 5745 6810 5753
rect 6757 5728 6766 5745
rect 6798 5728 6810 5745
rect 6757 5725 6810 5728
rect 5976 5651 6314 5664
rect 3257 5587 3289 5615
rect 3747 5600 4743 5626
rect 5476 5619 5587 5636
rect 5977 5632 6314 5651
rect 6256 5631 6314 5632
rect 6700 5659 6732 5666
rect 6700 5639 6707 5659
rect 6728 5639 6732 5659
rect 2877 5579 3289 5587
rect 2877 5553 2883 5579
rect 2909 5553 3289 5579
rect 2877 5551 3289 5553
rect 2879 5550 2919 5551
rect 3257 5486 3289 5551
rect 6700 5574 6732 5639
rect 6911 5651 6950 5924
rect 7146 5753 7180 5764
rect 7144 5752 7180 5753
rect 7144 5732 7151 5752
rect 7171 5732 7180 5752
rect 7144 5724 7180 5732
rect 6911 5610 6918 5651
rect 6939 5610 6950 5651
rect 6911 5595 6950 5610
rect 7070 5574 7110 5575
rect 6700 5572 7112 5574
rect 6700 5546 7080 5572
rect 7106 5546 7112 5572
rect 6700 5538 7112 5546
rect 3257 5466 3261 5486
rect 3282 5466 3289 5486
rect 3257 5459 3289 5466
rect 3675 5493 3733 5494
rect 3675 5474 4012 5493
rect 4402 5489 4513 5506
rect 5246 5499 6242 5525
rect 6700 5510 6732 5538
rect 7145 5518 7179 5724
rect 3675 5461 4013 5474
rect 2810 5393 2845 5401
rect 2810 5373 2818 5393
rect 2838 5373 2845 5393
rect 2810 5368 2845 5373
rect 3464 5388 3574 5403
rect 3464 5385 3541 5388
rect 2810 5325 2844 5368
rect 3464 5358 3467 5385
rect 3496 5361 3541 5385
rect 3570 5361 3574 5388
rect 3496 5358 3574 5361
rect 3464 5344 3574 5358
rect 3675 5325 3712 5461
rect 3981 5444 4013 5461
rect 4402 5469 4409 5489
rect 4428 5469 4486 5489
rect 4505 5469 4513 5489
rect 4402 5447 4513 5469
rect 5248 5446 5290 5499
rect 3981 5398 4012 5444
rect 5248 5427 5257 5446
rect 5282 5427 5290 5446
rect 5248 5417 5290 5427
rect 5476 5457 5586 5471
rect 5476 5454 5554 5457
rect 5476 5427 5480 5454
rect 5509 5430 5554 5454
rect 5583 5430 5586 5457
rect 6206 5447 6240 5499
rect 6700 5490 6705 5510
rect 6726 5490 6732 5510
rect 6700 5483 6732 5490
rect 7123 5513 7179 5518
rect 7123 5493 7130 5513
rect 7150 5493 7179 5513
rect 7123 5486 7179 5493
rect 7123 5485 7158 5486
rect 6751 5451 6792 5452
rect 5509 5427 5586 5430
rect 5476 5412 5586 5427
rect 6205 5442 6240 5447
rect 6205 5422 6212 5442
rect 6232 5422 6240 5442
rect 6750 5441 6792 5451
rect 6205 5414 6240 5422
rect 3769 5395 3804 5396
rect 3748 5388 3804 5395
rect 3748 5368 3777 5388
rect 3797 5368 3804 5388
rect 3748 5363 3804 5368
rect 3981 5391 4020 5398
rect 3981 5371 3987 5391
rect 4012 5371 4020 5391
rect 3981 5365 4020 5371
rect 4195 5391 4227 5398
rect 4195 5371 4201 5391
rect 4222 5371 4227 5391
rect 2554 5282 2601 5300
rect 2809 5290 3713 5325
rect 2810 5289 2844 5290
rect 2471 5223 2523 5228
rect 2926 5223 2971 5225
rect 2471 5208 2971 5223
rect 2471 5155 2485 5208
rect 2516 5184 2971 5208
rect 2516 5183 2541 5184
rect 2516 5155 2523 5183
rect 1501 5123 1578 5126
rect 1468 5108 1578 5123
rect 2193 5138 2374 5144
rect 2193 5118 2204 5138
rect 2224 5118 2374 5138
rect 2471 5131 2523 5155
rect 2193 5112 2374 5118
rect 2197 5110 2232 5112
rect 1212 5052 1273 5054
rect 910 5023 1273 5052
rect 1753 5045 1785 5052
rect 1753 5025 1760 5045
rect 1781 5025 1785 5045
rect 910 5021 1212 5023
rect 1753 4960 1785 5025
rect 2123 4960 2163 4961
rect 1753 4958 2165 4960
rect 1152 4935 1187 4937
rect 188 4932 1187 4935
rect 187 4908 1187 4932
rect 187 4753 235 4908
rect 421 4867 531 4881
rect 421 4864 499 4867
rect 421 4837 425 4864
rect 454 4840 499 4864
rect 528 4840 531 4867
rect 1152 4857 1187 4908
rect 1753 4932 2133 4958
rect 2159 4932 2165 4958
rect 1753 4924 2165 4932
rect 1753 4896 1785 4924
rect 2198 4904 2232 5110
rect 2722 5109 2757 5110
rect 1753 4876 1758 4896
rect 1779 4876 1785 4896
rect 1753 4869 1785 4876
rect 1955 4899 2000 4904
rect 1955 4875 1966 4899
rect 1992 4875 2000 4899
rect 1955 4864 2000 4875
rect 2176 4899 2232 4904
rect 2176 4879 2183 4899
rect 2203 4879 2232 4899
rect 2176 4872 2232 4879
rect 2701 5102 2757 5109
rect 2701 5082 2730 5102
rect 2750 5082 2757 5102
rect 2701 5077 2757 5082
rect 2926 5105 2971 5184
rect 3355 5203 3466 5220
rect 3355 5183 3362 5203
rect 3381 5183 3439 5203
rect 3458 5183 3466 5203
rect 3355 5161 3466 5183
rect 3748 5157 3782 5363
rect 4195 5343 4227 5371
rect 3815 5335 4227 5343
rect 3815 5309 3821 5335
rect 3847 5309 4227 5335
rect 3815 5307 4227 5309
rect 3817 5306 3857 5307
rect 4195 5242 4227 5307
rect 5761 5349 5793 5356
rect 5761 5329 5768 5349
rect 5789 5329 5793 5349
rect 5761 5264 5793 5329
rect 6131 5264 6171 5265
rect 5761 5262 6173 5264
rect 4195 5222 4199 5242
rect 4220 5222 4227 5242
rect 4195 5215 4227 5222
rect 4698 5257 4746 5262
rect 4698 5228 4709 5257
rect 4738 5228 4746 5257
rect 3748 5156 3783 5157
rect 3746 5149 3783 5156
rect 3746 5129 3756 5149
rect 3776 5129 3783 5149
rect 3746 5124 3783 5129
rect 4402 5144 4512 5159
rect 4402 5141 4479 5144
rect 2926 5085 2937 5105
rect 2962 5085 2971 5105
rect 2926 5081 2971 5085
rect 3148 5105 3180 5112
rect 3148 5085 3154 5105
rect 3175 5085 3180 5105
rect 2176 4871 2211 4872
rect 2701 4871 2735 5077
rect 3148 5057 3180 5085
rect 2768 5049 3180 5057
rect 2768 5023 2774 5049
rect 2800 5023 3180 5049
rect 3746 5073 3781 5124
rect 4402 5114 4405 5141
rect 4434 5117 4479 5141
rect 4508 5117 4512 5144
rect 4434 5114 4512 5117
rect 4402 5100 4512 5114
rect 4698 5073 4746 5228
rect 5761 5236 6141 5262
rect 6167 5236 6173 5262
rect 5761 5228 6173 5236
rect 5761 5200 5793 5228
rect 6206 5208 6240 5414
rect 6414 5412 6525 5434
rect 6414 5392 6422 5412
rect 6441 5392 6499 5412
rect 6518 5392 6525 5412
rect 6414 5375 6525 5392
rect 6750 5419 6757 5441
rect 6783 5419 6792 5441
rect 6750 5410 6792 5419
rect 5967 5205 6010 5207
rect 5761 5180 5766 5200
rect 5787 5180 5793 5200
rect 5761 5173 5793 5180
rect 5966 5198 6010 5205
rect 5966 5178 5976 5198
rect 5999 5178 6010 5198
rect 5966 5174 6010 5178
rect 6184 5203 6240 5208
rect 6184 5183 6191 5203
rect 6211 5183 6240 5203
rect 6184 5176 6240 5183
rect 6296 5344 6329 5345
rect 6750 5344 6787 5410
rect 7382 5387 7428 6872
rect 6296 5315 6787 5344
rect 6184 5175 6219 5176
rect 3746 5049 4746 5073
rect 5475 5102 5586 5124
rect 5475 5082 5483 5102
rect 5502 5082 5560 5102
rect 5579 5082 5586 5102
rect 5475 5065 5586 5082
rect 5966 5093 6008 5174
rect 6296 5095 6329 5315
rect 6750 5313 6787 5315
rect 7380 5363 7428 5387
rect 7610 5381 7657 6958
rect 8144 6915 8178 7094
rect 8409 7111 8519 7126
rect 8409 7108 8486 7111
rect 8409 7081 8412 7108
rect 8441 7084 8486 7108
rect 8515 7084 8519 7111
rect 8441 7081 8519 7084
rect 8409 7067 8519 7081
rect 7753 6890 8178 6915
rect 8257 6954 8294 6956
rect 8715 6954 8748 7174
rect 9036 7095 9078 7176
rect 9458 7187 9569 7203
rect 9458 7167 9465 7187
rect 9484 7167 9542 7187
rect 9561 7167 9569 7187
rect 9458 7145 9569 7167
rect 11784 7165 11816 7230
rect 12154 7165 12194 7166
rect 11784 7163 12196 7165
rect 11182 7146 11217 7148
rect 10218 7143 11217 7146
rect 10217 7119 11217 7143
rect 8825 7093 8860 7094
rect 8257 6925 8748 6954
rect 7753 6874 8177 6890
rect 7753 6483 7791 6874
rect 8257 6859 8294 6925
rect 8715 6924 8748 6925
rect 8804 7086 8860 7093
rect 8804 7066 8833 7086
rect 8853 7066 8860 7086
rect 8804 7061 8860 7066
rect 9034 7091 9078 7095
rect 9034 7071 9045 7091
rect 9068 7071 9078 7091
rect 9034 7064 9078 7071
rect 9251 7089 9283 7096
rect 9251 7069 9257 7089
rect 9278 7069 9283 7089
rect 9034 7062 9077 7064
rect 8252 6850 8294 6859
rect 8252 6828 8261 6850
rect 8287 6828 8294 6850
rect 8519 6877 8630 6894
rect 8519 6857 8526 6877
rect 8545 6857 8603 6877
rect 8622 6857 8630 6877
rect 8519 6835 8630 6857
rect 8804 6855 8838 7061
rect 9251 7041 9283 7069
rect 8871 7033 9283 7041
rect 8871 7007 8877 7033
rect 8903 7007 9283 7033
rect 8871 7005 9283 7007
rect 8873 7004 8913 7005
rect 9251 6940 9283 7005
rect 9251 6920 9255 6940
rect 9276 6920 9283 6940
rect 10217 6964 10265 7119
rect 10451 7078 10561 7092
rect 10451 7075 10529 7078
rect 10451 7048 10455 7075
rect 10484 7051 10529 7075
rect 10558 7051 10561 7078
rect 11182 7068 11217 7119
rect 11784 7137 12164 7163
rect 12190 7137 12196 7163
rect 11784 7129 12196 7137
rect 11784 7101 11816 7129
rect 11784 7081 11789 7101
rect 11810 7081 11816 7101
rect 11784 7074 11816 7081
rect 11990 7100 12035 7112
rect 12229 7109 12263 7315
rect 11990 7081 11997 7100
rect 12026 7081 12035 7100
rect 10484 7048 10561 7051
rect 10451 7033 10561 7048
rect 11180 7063 11217 7068
rect 11180 7043 11187 7063
rect 11207 7043 11217 7063
rect 11180 7036 11217 7043
rect 11180 7035 11215 7036
rect 10217 6935 10225 6964
rect 10254 6935 10265 6964
rect 10217 6930 10265 6935
rect 10736 6970 10768 6977
rect 10736 6950 10743 6970
rect 10764 6950 10768 6970
rect 9251 6913 9283 6920
rect 10736 6885 10768 6950
rect 11106 6885 11146 6886
rect 10736 6883 11148 6885
rect 10736 6857 11116 6883
rect 11142 6857 11148 6883
rect 8804 6847 8839 6855
rect 8252 6818 8294 6828
rect 8804 6827 8812 6847
rect 8832 6827 8839 6847
rect 8804 6822 8839 6827
rect 9458 6842 9568 6857
rect 9458 6839 9535 6842
rect 8252 6817 8293 6818
rect 7886 6783 7921 6784
rect 7865 6776 7921 6783
rect 7865 6756 7894 6776
rect 7914 6756 7921 6776
rect 7865 6751 7921 6756
rect 8312 6779 8344 6786
rect 8312 6759 8318 6779
rect 8339 6759 8344 6779
rect 8804 6770 8838 6822
rect 9458 6812 9461 6839
rect 9490 6815 9535 6839
rect 9564 6815 9568 6842
rect 9490 6812 9568 6815
rect 9458 6798 9568 6812
rect 9754 6842 9796 6852
rect 9754 6823 9762 6842
rect 9787 6823 9796 6842
rect 9754 6770 9796 6823
rect 10736 6849 11148 6857
rect 10736 6821 10768 6849
rect 11181 6829 11215 7035
rect 11498 7003 11609 7025
rect 11498 6983 11506 7003
rect 11525 6983 11583 7003
rect 11602 6983 11609 7003
rect 11498 6966 11609 6983
rect 11990 6998 12035 7081
rect 12207 7104 12263 7109
rect 12207 7084 12214 7104
rect 12234 7084 12263 7104
rect 12730 7299 12759 7319
rect 12779 7299 12786 7319
rect 12730 7294 12786 7299
rect 13177 7322 13209 7329
rect 13177 7302 13183 7322
rect 13204 7302 13209 7322
rect 12730 7088 12764 7294
rect 13177 7274 13209 7302
rect 12797 7266 13209 7274
rect 12797 7240 12803 7266
rect 12829 7240 13209 7266
rect 13776 7284 13811 7335
rect 14432 7325 14435 7352
rect 14464 7328 14509 7352
rect 14538 7328 14542 7355
rect 14464 7325 14542 7328
rect 14432 7311 14542 7325
rect 14728 7284 14776 7439
rect 15791 7447 16171 7473
rect 16197 7447 16203 7473
rect 15791 7439 16203 7447
rect 15791 7411 15823 7439
rect 16236 7419 16270 7625
rect 16444 7623 16555 7645
rect 16444 7603 16452 7623
rect 16471 7603 16529 7623
rect 16548 7603 16555 7623
rect 16444 7586 16555 7603
rect 16780 7630 16787 7652
rect 16813 7630 16822 7652
rect 16780 7621 16822 7630
rect 15997 7416 16040 7418
rect 15791 7391 15796 7411
rect 15817 7391 15823 7411
rect 15791 7384 15823 7391
rect 15996 7409 16040 7416
rect 15996 7389 16006 7409
rect 16029 7389 16040 7409
rect 15996 7385 16040 7389
rect 16214 7414 16270 7419
rect 16214 7394 16221 7414
rect 16241 7394 16270 7414
rect 16214 7387 16270 7394
rect 16326 7555 16359 7556
rect 16780 7555 16817 7621
rect 16326 7526 16817 7555
rect 16214 7386 16249 7387
rect 13776 7260 14776 7284
rect 15505 7313 15616 7335
rect 15505 7293 15513 7313
rect 15532 7293 15590 7313
rect 15609 7293 15616 7313
rect 15505 7277 15616 7293
rect 15996 7304 16038 7385
rect 16326 7306 16359 7526
rect 16780 7524 16817 7526
rect 16555 7399 16665 7413
rect 16555 7396 16633 7399
rect 16555 7369 16559 7396
rect 16588 7372 16633 7396
rect 16662 7372 16665 7399
rect 16588 7369 16665 7372
rect 16555 7354 16665 7369
rect 17283 7384 17321 7997
rect 17799 7992 18030 8025
rect 17799 7451 17849 7992
rect 17986 7988 18030 7992
rect 17917 7891 17952 7892
rect 17896 7884 17952 7891
rect 17896 7864 17925 7884
rect 17945 7864 17952 7884
rect 17896 7859 17952 7864
rect 18127 7883 18165 8221
rect 18409 8232 18519 8247
rect 18409 8229 18486 8232
rect 18409 8202 18412 8229
rect 18441 8205 18486 8229
rect 18515 8205 18519 8232
rect 18441 8202 18519 8205
rect 18409 8188 18519 8202
rect 18288 8062 18325 8064
rect 18746 8062 18779 8282
rect 19067 8203 19109 8284
rect 19489 8295 19600 8312
rect 19489 8275 19496 8295
rect 19515 8275 19573 8295
rect 19592 8275 19600 8295
rect 19489 8253 19600 8275
rect 18856 8201 18891 8202
rect 18288 8033 18779 8062
rect 18288 7967 18325 8033
rect 18746 8032 18779 8033
rect 18835 8194 18891 8201
rect 18835 8174 18864 8194
rect 18884 8174 18891 8194
rect 18835 8169 18891 8174
rect 19065 8199 19109 8203
rect 19065 8179 19076 8199
rect 19099 8179 19109 8199
rect 19065 8172 19109 8179
rect 19282 8197 19314 8204
rect 19282 8177 19288 8197
rect 19309 8177 19314 8197
rect 19065 8170 19108 8172
rect 18283 7958 18325 7967
rect 18283 7936 18292 7958
rect 18318 7936 18325 7958
rect 18550 7985 18661 8002
rect 18550 7965 18557 7985
rect 18576 7965 18634 7985
rect 18653 7965 18661 7985
rect 18550 7943 18661 7965
rect 18835 7963 18869 8169
rect 19282 8149 19314 8177
rect 18902 8141 19314 8149
rect 18902 8115 18908 8141
rect 18934 8115 19314 8141
rect 18902 8113 19314 8115
rect 18904 8112 18944 8113
rect 19282 8048 19314 8113
rect 19282 8028 19286 8048
rect 19307 8028 19314 8048
rect 19282 8021 19314 8028
rect 18835 7955 18870 7963
rect 18283 7926 18325 7936
rect 18835 7935 18843 7955
rect 18863 7935 18870 7955
rect 18835 7930 18870 7935
rect 19489 7950 19599 7965
rect 19489 7947 19566 7950
rect 18283 7925 18324 7926
rect 18127 7866 18135 7883
rect 18155 7866 18165 7883
rect 17896 7653 17930 7859
rect 18127 7856 18165 7866
rect 18343 7887 18375 7894
rect 18343 7867 18349 7887
rect 18370 7867 18375 7887
rect 18835 7878 18869 7930
rect 19489 7920 19492 7947
rect 19521 7923 19566 7947
rect 19595 7923 19599 7950
rect 19521 7920 19599 7923
rect 19489 7906 19599 7920
rect 19785 7950 19827 7960
rect 19785 7931 19793 7950
rect 19818 7931 19827 7950
rect 19785 7878 19827 7931
rect 18343 7839 18375 7867
rect 18833 7852 19829 7878
rect 17963 7831 18375 7839
rect 17963 7805 17969 7831
rect 17995 7805 18375 7831
rect 17963 7803 18375 7805
rect 17965 7802 18005 7803
rect 18343 7738 18375 7803
rect 18343 7718 18347 7738
rect 18368 7718 18375 7738
rect 18343 7711 18375 7718
rect 18761 7745 18819 7746
rect 18761 7726 19098 7745
rect 19488 7741 19599 7758
rect 18761 7713 19099 7726
rect 17896 7645 17931 7653
rect 17896 7625 17904 7645
rect 17924 7625 17931 7645
rect 17896 7620 17931 7625
rect 18550 7640 18660 7655
rect 18550 7637 18627 7640
rect 17896 7577 17930 7620
rect 18550 7610 18553 7637
rect 18582 7613 18627 7637
rect 18656 7613 18660 7640
rect 18582 7610 18660 7613
rect 18550 7596 18660 7610
rect 18761 7577 18798 7713
rect 19067 7696 19099 7713
rect 19488 7721 19495 7741
rect 19514 7721 19572 7741
rect 19591 7721 19599 7741
rect 19488 7699 19599 7721
rect 19067 7650 19098 7696
rect 18855 7647 18890 7648
rect 18834 7640 18890 7647
rect 18834 7620 18863 7640
rect 18883 7620 18890 7640
rect 18834 7615 18890 7620
rect 19067 7643 19106 7650
rect 19067 7623 19073 7643
rect 19098 7623 19106 7643
rect 19067 7617 19106 7623
rect 19281 7643 19313 7650
rect 19281 7623 19287 7643
rect 19308 7623 19313 7643
rect 17895 7542 18799 7577
rect 17896 7541 17930 7542
rect 17777 7442 17849 7451
rect 17777 7413 17794 7442
rect 17842 7413 17849 7442
rect 18440 7461 18551 7478
rect 18440 7441 18447 7461
rect 18466 7441 18524 7461
rect 18543 7441 18551 7461
rect 18440 7419 18551 7441
rect 17777 7406 17849 7413
rect 18834 7409 18868 7615
rect 19281 7595 19313 7623
rect 18901 7587 19313 7595
rect 18901 7561 18907 7587
rect 18933 7561 19313 7587
rect 18901 7559 19313 7561
rect 18903 7558 18943 7559
rect 19281 7494 19313 7559
rect 19281 7474 19285 7494
rect 19306 7474 19313 7494
rect 19281 7467 19313 7474
rect 19784 7509 19832 7514
rect 19784 7480 19795 7509
rect 19824 7480 19832 7509
rect 18834 7408 18869 7409
rect 17777 7396 17847 7406
rect 18832 7401 18869 7408
rect 17283 7364 17291 7384
rect 17311 7364 17321 7384
rect 18832 7381 18842 7401
rect 18862 7381 18869 7401
rect 18832 7376 18869 7381
rect 19488 7396 19598 7411
rect 19488 7393 19565 7396
rect 17807 7367 17842 7368
rect 17283 7357 17321 7364
rect 17786 7360 17842 7367
rect 17284 7356 17319 7357
rect 16298 7304 16359 7306
rect 15996 7275 16359 7304
rect 16840 7291 16872 7298
rect 15996 7273 16298 7275
rect 16840 7271 16847 7291
rect 16868 7271 16872 7291
rect 13776 7257 14775 7260
rect 13776 7255 13811 7257
rect 12797 7238 13209 7240
rect 12799 7237 12839 7238
rect 12965 7197 13000 7215
rect 12965 7165 12968 7197
rect 12995 7165 13000 7197
rect 12730 7087 12765 7088
rect 12207 7077 12263 7084
rect 12728 7080 12766 7087
rect 12207 7076 12242 7077
rect 12728 7076 12738 7080
rect 12722 7062 12738 7076
rect 12758 7076 12766 7080
rect 12758 7062 12772 7076
rect 12722 7055 12772 7062
rect 12355 6998 12405 7000
rect 11990 6964 12405 6998
rect 12119 6902 12153 6903
rect 11250 6867 12154 6902
rect 12202 6891 12270 6902
rect 12202 6870 12207 6891
rect 10736 6801 10741 6821
rect 10762 6801 10768 6821
rect 10736 6794 10768 6801
rect 10943 6821 10982 6827
rect 10943 6801 10951 6821
rect 10976 6801 10982 6821
rect 10943 6794 10982 6801
rect 11159 6824 11215 6829
rect 11159 6804 11166 6824
rect 11186 6804 11215 6824
rect 11159 6797 11215 6804
rect 11159 6796 11194 6797
rect 7865 6545 7899 6751
rect 8312 6731 8344 6759
rect 8802 6744 9798 6770
rect 10951 6748 10982 6794
rect 7932 6723 8344 6731
rect 7932 6697 7938 6723
rect 7964 6697 8344 6723
rect 7932 6695 8344 6697
rect 7934 6694 7974 6695
rect 8094 6659 8133 6674
rect 8094 6618 8105 6659
rect 8126 6618 8133 6659
rect 7864 6537 7900 6545
rect 7864 6517 7873 6537
rect 7893 6517 7900 6537
rect 7864 6516 7900 6517
rect 7864 6505 7898 6516
rect 7754 6475 7791 6483
rect 7754 6441 7998 6475
rect 7746 6272 7781 6273
rect 7725 6265 7781 6272
rect 7725 6245 7754 6265
rect 7774 6245 7781 6265
rect 7725 6240 7781 6245
rect 7956 6270 7998 6441
rect 8094 6345 8133 6618
rect 8312 6630 8344 6695
rect 10450 6723 10561 6745
rect 10450 6703 10458 6723
rect 10477 6703 10535 6723
rect 10554 6703 10561 6723
rect 10950 6731 10982 6748
rect 11251 6731 11288 6867
rect 11389 6834 11499 6848
rect 11389 6831 11467 6834
rect 11389 6804 11393 6831
rect 11422 6807 11467 6831
rect 11496 6807 11499 6834
rect 12119 6824 12153 6867
rect 11422 6804 11499 6807
rect 11389 6789 11499 6804
rect 12118 6819 12153 6824
rect 12118 6799 12125 6819
rect 12145 6799 12153 6819
rect 12118 6791 12153 6799
rect 10950 6718 11288 6731
rect 10450 6686 10561 6703
rect 10951 6699 11288 6718
rect 11230 6698 11288 6699
rect 11674 6726 11706 6733
rect 11674 6706 11681 6726
rect 11702 6706 11706 6726
rect 8312 6610 8316 6630
rect 8337 6610 8344 6630
rect 8312 6603 8344 6610
rect 8730 6637 8788 6638
rect 8730 6618 9067 6637
rect 9457 6633 9568 6650
rect 8730 6605 9068 6618
rect 8234 6541 8287 6544
rect 8234 6524 8246 6541
rect 8278 6524 8287 6541
rect 8234 6516 8287 6524
rect 8233 6469 8287 6516
rect 8519 6532 8629 6547
rect 8519 6529 8596 6532
rect 8519 6502 8522 6529
rect 8551 6505 8596 6529
rect 8625 6505 8629 6532
rect 8551 6502 8629 6505
rect 8519 6488 8629 6502
rect 8730 6469 8767 6605
rect 9036 6588 9068 6605
rect 9457 6613 9464 6633
rect 9483 6613 9541 6633
rect 9560 6613 9568 6633
rect 9457 6591 9568 6613
rect 11674 6641 11706 6706
rect 12044 6641 12084 6642
rect 11674 6639 12086 6641
rect 11674 6613 12054 6639
rect 12080 6613 12086 6639
rect 11674 6605 12086 6613
rect 9036 6542 9067 6588
rect 10220 6566 11216 6592
rect 11674 6577 11706 6605
rect 8824 6539 8859 6540
rect 8803 6532 8859 6539
rect 8803 6512 8832 6532
rect 8852 6512 8859 6532
rect 8803 6507 8859 6512
rect 9036 6535 9075 6542
rect 9036 6515 9042 6535
rect 9067 6515 9075 6535
rect 9036 6509 9075 6515
rect 9250 6535 9282 6542
rect 9250 6515 9256 6535
rect 9277 6515 9282 6535
rect 8233 6434 8768 6469
rect 8233 6430 8286 6434
rect 8094 6318 8098 6345
rect 8129 6318 8133 6345
rect 8379 6366 8490 6383
rect 8379 6346 8386 6366
rect 8405 6346 8463 6366
rect 8482 6346 8490 6366
rect 8379 6324 8490 6346
rect 8094 6311 8133 6318
rect 8803 6301 8837 6507
rect 9250 6487 9282 6515
rect 8870 6479 9282 6487
rect 10222 6513 10264 6566
rect 10222 6494 10231 6513
rect 10256 6494 10264 6513
rect 10222 6484 10264 6494
rect 10450 6524 10560 6538
rect 10450 6521 10528 6524
rect 10450 6494 10454 6521
rect 10483 6497 10528 6521
rect 10557 6497 10560 6524
rect 11180 6514 11214 6566
rect 11674 6557 11679 6577
rect 11700 6557 11706 6577
rect 11674 6550 11706 6557
rect 11884 6578 11922 6588
rect 12119 6585 12153 6791
rect 11884 6561 11894 6578
rect 11914 6561 11922 6578
rect 11725 6518 11766 6519
rect 10483 6494 10560 6497
rect 10450 6479 10560 6494
rect 11179 6509 11214 6514
rect 11179 6489 11186 6509
rect 11206 6489 11214 6509
rect 11724 6508 11766 6518
rect 11179 6481 11214 6489
rect 8870 6453 8876 6479
rect 8902 6453 9282 6479
rect 8870 6451 9282 6453
rect 8872 6450 8912 6451
rect 9250 6386 9282 6451
rect 10735 6416 10767 6423
rect 9250 6366 9254 6386
rect 9275 6366 9282 6386
rect 9250 6359 9282 6366
rect 9753 6401 9801 6406
rect 9753 6372 9764 6401
rect 9793 6372 9801 6401
rect 8803 6300 8838 6301
rect 8801 6293 8838 6300
rect 7956 6249 7964 6270
rect 7991 6249 7998 6270
rect 7725 6034 7759 6240
rect 7956 6238 7998 6249
rect 8172 6268 8204 6275
rect 8172 6248 8178 6268
rect 8199 6248 8204 6268
rect 8172 6220 8204 6248
rect 7792 6212 8204 6220
rect 7792 6186 7798 6212
rect 7824 6186 8204 6212
rect 8801 6273 8811 6293
rect 8831 6273 8838 6293
rect 8801 6268 8838 6273
rect 9457 6288 9567 6303
rect 9457 6285 9534 6288
rect 8801 6217 8836 6268
rect 9457 6258 9460 6285
rect 9489 6261 9534 6285
rect 9563 6261 9567 6288
rect 9489 6258 9567 6261
rect 9457 6244 9567 6258
rect 9753 6217 9801 6372
rect 10735 6396 10742 6416
rect 10763 6396 10767 6416
rect 10735 6331 10767 6396
rect 11105 6331 11145 6332
rect 10735 6329 11147 6331
rect 10735 6303 11115 6329
rect 11141 6303 11147 6329
rect 10735 6295 11147 6303
rect 10735 6267 10767 6295
rect 11180 6275 11214 6481
rect 11388 6479 11499 6501
rect 11388 6459 11396 6479
rect 11415 6459 11473 6479
rect 11492 6459 11499 6479
rect 11388 6442 11499 6459
rect 11724 6486 11731 6508
rect 11757 6486 11766 6508
rect 11724 6477 11766 6486
rect 10941 6272 10984 6274
rect 10735 6247 10740 6267
rect 10761 6247 10767 6267
rect 10735 6240 10767 6247
rect 10940 6265 10984 6272
rect 10940 6245 10950 6265
rect 10973 6245 10984 6265
rect 10940 6241 10984 6245
rect 11158 6270 11214 6275
rect 11158 6250 11165 6270
rect 11185 6250 11214 6270
rect 11158 6243 11214 6250
rect 11270 6411 11303 6412
rect 11724 6411 11761 6477
rect 11270 6382 11761 6411
rect 11158 6242 11193 6243
rect 8801 6193 9801 6217
rect 8801 6190 9800 6193
rect 8801 6188 8836 6190
rect 7792 6184 8204 6186
rect 7794 6183 7834 6184
rect 8172 6119 8204 6184
rect 10449 6169 10560 6191
rect 10449 6149 10457 6169
rect 10476 6149 10534 6169
rect 10553 6149 10560 6169
rect 10449 6132 10560 6149
rect 10940 6160 10982 6241
rect 11270 6162 11303 6382
rect 11724 6380 11761 6382
rect 11530 6242 11640 6256
rect 11530 6239 11608 6242
rect 11530 6212 11534 6239
rect 11563 6215 11608 6239
rect 11637 6215 11640 6242
rect 11563 6212 11640 6215
rect 11530 6197 11640 6212
rect 11884 6223 11922 6561
rect 12097 6580 12153 6585
rect 12097 6560 12104 6580
rect 12124 6560 12153 6580
rect 12097 6553 12153 6560
rect 12200 6862 12207 6870
rect 12255 6862 12270 6891
rect 12200 6853 12270 6862
rect 12097 6552 12132 6553
rect 12019 6452 12063 6456
rect 12200 6452 12250 6853
rect 12355 6836 12405 6964
rect 12588 6977 12698 6979
rect 12965 6977 13000 7165
rect 13177 7173 13209 7238
rect 16840 7206 16872 7271
rect 17210 7206 17250 7207
rect 16840 7204 17252 7206
rect 16238 7187 16273 7189
rect 15274 7184 16273 7187
rect 13177 7153 13181 7173
rect 13202 7153 13209 7173
rect 13751 7169 14053 7171
rect 13177 7146 13209 7153
rect 13690 7140 14053 7169
rect 13690 7138 13751 7140
rect 12588 6947 13000 6977
rect 12588 6922 12632 6947
rect 12671 6944 13000 6947
rect 13119 7078 13153 7084
rect 13119 7058 13128 7078
rect 13149 7058 13153 7078
rect 12019 6419 12250 6452
rect 12019 6417 12226 6419
rect 12019 6263 12063 6417
rect 11884 6206 11892 6223
rect 11912 6206 11922 6223
rect 11884 6200 11922 6206
rect 11242 6160 11303 6162
rect 10940 6131 11303 6160
rect 11815 6134 11847 6141
rect 10940 6129 11242 6131
rect 8172 6099 8176 6119
rect 8197 6099 8204 6119
rect 11815 6114 11822 6134
rect 11843 6114 11847 6134
rect 8777 6102 9079 6104
rect 8172 6092 8204 6099
rect 8716 6073 9079 6102
rect 8716 6071 8777 6073
rect 7725 6026 7760 6034
rect 7725 6006 7733 6026
rect 7753 6006 7760 6026
rect 7725 6001 7760 6006
rect 8097 6027 8135 6033
rect 8097 6010 8107 6027
rect 8127 6010 8135 6027
rect 7725 6000 7757 6001
rect 7887 5680 7922 5681
rect 6524 5194 6634 5208
rect 6524 5191 6602 5194
rect 6524 5164 6528 5191
rect 6557 5167 6602 5191
rect 6631 5167 6634 5194
rect 7380 5185 7427 5363
rect 7610 5341 7623 5381
rect 7650 5341 7657 5381
rect 7866 5673 7922 5680
rect 7866 5653 7895 5673
rect 7915 5653 7922 5673
rect 7866 5648 7922 5653
rect 8097 5672 8135 6010
rect 8379 6021 8489 6036
rect 8379 6018 8456 6021
rect 8379 5991 8382 6018
rect 8411 5994 8456 6018
rect 8485 5994 8489 6021
rect 8411 5991 8489 5994
rect 8379 5977 8489 5991
rect 8258 5851 8295 5853
rect 8716 5851 8749 6071
rect 9037 5992 9079 6073
rect 9459 6084 9570 6101
rect 9459 6064 9466 6084
rect 9485 6064 9543 6084
rect 9562 6064 9570 6084
rect 9459 6042 9570 6064
rect 11815 6049 11847 6114
rect 12025 6127 12063 6263
rect 12262 6232 12293 6233
rect 12259 6227 12293 6232
rect 12259 6207 12266 6227
rect 12286 6207 12293 6227
rect 12259 6199 12293 6207
rect 12025 6089 12031 6127
rect 12054 6089 12063 6127
rect 12025 6079 12063 6089
rect 12260 6141 12293 6199
rect 12185 6049 12225 6050
rect 11815 6047 12227 6049
rect 11183 6043 11218 6045
rect 10219 6040 11218 6043
rect 10218 6016 11218 6040
rect 8826 5990 8861 5991
rect 8258 5822 8749 5851
rect 8258 5756 8295 5822
rect 8716 5821 8749 5822
rect 8805 5983 8861 5990
rect 8805 5963 8834 5983
rect 8854 5963 8861 5983
rect 8805 5958 8861 5963
rect 9035 5988 9079 5992
rect 9035 5968 9046 5988
rect 9069 5968 9079 5988
rect 9035 5961 9079 5968
rect 9252 5986 9284 5993
rect 9252 5966 9258 5986
rect 9279 5966 9284 5986
rect 9035 5959 9078 5961
rect 8253 5747 8295 5756
rect 8253 5725 8262 5747
rect 8288 5725 8295 5747
rect 8520 5774 8631 5791
rect 8520 5754 8527 5774
rect 8546 5754 8604 5774
rect 8623 5754 8631 5774
rect 8520 5732 8631 5754
rect 8805 5752 8839 5958
rect 9252 5938 9284 5966
rect 8872 5930 9284 5938
rect 8872 5904 8878 5930
rect 8904 5904 9284 5930
rect 8872 5902 9284 5904
rect 8874 5901 8914 5902
rect 9252 5837 9284 5902
rect 9252 5817 9256 5837
rect 9277 5817 9284 5837
rect 10218 5861 10266 6016
rect 10452 5975 10562 5989
rect 10452 5972 10530 5975
rect 10452 5945 10456 5972
rect 10485 5948 10530 5972
rect 10559 5948 10562 5975
rect 11183 5965 11218 6016
rect 10485 5945 10562 5948
rect 10452 5930 10562 5945
rect 11181 5960 11218 5965
rect 11181 5940 11188 5960
rect 11208 5940 11218 5960
rect 11815 6021 12195 6047
rect 12221 6021 12227 6047
rect 11815 6013 12227 6021
rect 11815 5985 11847 6013
rect 12260 5993 12296 6141
rect 11815 5965 11820 5985
rect 11841 5965 11847 5985
rect 11815 5958 11847 5965
rect 12238 5988 12296 5993
rect 12238 5968 12245 5988
rect 12265 5968 12296 5988
rect 12238 5961 12296 5968
rect 12238 5960 12273 5961
rect 11181 5933 11218 5940
rect 11181 5932 11216 5933
rect 10218 5832 10226 5861
rect 10255 5832 10266 5861
rect 10218 5827 10266 5832
rect 10737 5867 10769 5874
rect 10737 5847 10744 5867
rect 10765 5847 10769 5867
rect 9252 5810 9284 5817
rect 10737 5782 10769 5847
rect 11107 5782 11147 5783
rect 10737 5780 11149 5782
rect 10737 5754 11117 5780
rect 11143 5754 11149 5780
rect 8805 5744 8840 5752
rect 8253 5715 8295 5725
rect 8805 5724 8813 5744
rect 8833 5724 8840 5744
rect 8805 5719 8840 5724
rect 9459 5739 9569 5754
rect 9459 5736 9536 5739
rect 8253 5714 8294 5715
rect 8097 5655 8105 5672
rect 8125 5655 8135 5672
rect 7866 5442 7900 5648
rect 8097 5645 8135 5655
rect 8313 5676 8345 5683
rect 8313 5656 8319 5676
rect 8340 5656 8345 5676
rect 8805 5667 8839 5719
rect 9459 5709 9462 5736
rect 9491 5712 9536 5736
rect 9565 5712 9569 5739
rect 9491 5709 9569 5712
rect 9459 5695 9569 5709
rect 9755 5739 9797 5749
rect 9755 5720 9763 5739
rect 9788 5720 9797 5739
rect 9755 5667 9797 5720
rect 10737 5746 11149 5754
rect 10737 5718 10769 5746
rect 11182 5726 11216 5932
rect 11886 5915 11925 5922
rect 11529 5887 11640 5909
rect 11529 5867 11537 5887
rect 11556 5867 11614 5887
rect 11633 5867 11640 5887
rect 11529 5850 11640 5867
rect 11886 5888 11890 5915
rect 11921 5888 11925 5915
rect 11733 5799 11786 5803
rect 11251 5764 11786 5799
rect 10737 5698 10742 5718
rect 10763 5698 10769 5718
rect 10737 5691 10769 5698
rect 10944 5718 10983 5724
rect 10944 5698 10952 5718
rect 10977 5698 10983 5718
rect 10944 5691 10983 5698
rect 11160 5721 11216 5726
rect 11160 5701 11167 5721
rect 11187 5701 11216 5721
rect 11160 5694 11216 5701
rect 11160 5693 11195 5694
rect 8313 5628 8345 5656
rect 8803 5641 9799 5667
rect 10952 5645 10983 5691
rect 7933 5620 8345 5628
rect 7933 5594 7939 5620
rect 7965 5594 8345 5620
rect 7933 5592 8345 5594
rect 7935 5591 7975 5592
rect 8313 5527 8345 5592
rect 10451 5620 10562 5642
rect 10451 5600 10459 5620
rect 10478 5600 10536 5620
rect 10555 5600 10562 5620
rect 10951 5628 10983 5645
rect 11252 5628 11289 5764
rect 11390 5731 11500 5745
rect 11390 5728 11468 5731
rect 11390 5701 11394 5728
rect 11423 5704 11468 5728
rect 11497 5704 11500 5731
rect 11423 5701 11500 5704
rect 11390 5686 11500 5701
rect 11732 5717 11786 5764
rect 11732 5709 11785 5717
rect 11732 5692 11741 5709
rect 11773 5692 11785 5709
rect 11732 5689 11785 5692
rect 10951 5615 11289 5628
rect 10451 5583 10562 5600
rect 10952 5596 11289 5615
rect 11231 5595 11289 5596
rect 11675 5623 11707 5630
rect 11675 5603 11682 5623
rect 11703 5603 11707 5623
rect 8313 5507 8317 5527
rect 8338 5507 8345 5527
rect 8313 5500 8345 5507
rect 8731 5534 8789 5535
rect 8731 5515 9068 5534
rect 9458 5530 9569 5547
rect 8731 5502 9069 5515
rect 7866 5434 7901 5442
rect 7866 5414 7874 5434
rect 7894 5414 7901 5434
rect 7866 5409 7901 5414
rect 8520 5429 8630 5444
rect 8520 5426 8597 5429
rect 7866 5366 7900 5409
rect 8520 5399 8523 5426
rect 8552 5402 8597 5426
rect 8626 5402 8630 5429
rect 8552 5399 8630 5402
rect 8520 5385 8630 5399
rect 8731 5366 8768 5502
rect 9037 5485 9069 5502
rect 9458 5510 9465 5530
rect 9484 5510 9542 5530
rect 9561 5510 9569 5530
rect 9458 5488 9569 5510
rect 11675 5538 11707 5603
rect 11886 5615 11925 5888
rect 12121 5717 12155 5728
rect 12119 5716 12155 5717
rect 12119 5696 12126 5716
rect 12146 5696 12155 5716
rect 12119 5688 12155 5696
rect 11886 5574 11893 5615
rect 11914 5574 11925 5615
rect 11886 5559 11925 5574
rect 12045 5538 12085 5539
rect 11675 5536 12087 5538
rect 11675 5510 12055 5536
rect 12081 5510 12087 5536
rect 11675 5502 12087 5510
rect 9037 5439 9068 5485
rect 10221 5463 11217 5489
rect 11675 5474 11707 5502
rect 12120 5482 12154 5688
rect 8825 5436 8860 5437
rect 8804 5429 8860 5436
rect 8804 5409 8833 5429
rect 8853 5409 8860 5429
rect 8804 5404 8860 5409
rect 9037 5432 9076 5439
rect 9037 5412 9043 5432
rect 9068 5412 9076 5432
rect 9037 5406 9076 5412
rect 9251 5432 9283 5439
rect 9251 5412 9257 5432
rect 9278 5412 9283 5432
rect 7610 5323 7657 5341
rect 7865 5331 8769 5366
rect 7866 5330 7900 5331
rect 7527 5264 7579 5269
rect 7982 5264 8027 5266
rect 7527 5249 8027 5264
rect 7527 5196 7541 5249
rect 7572 5225 8027 5249
rect 7572 5224 7597 5225
rect 7572 5196 7579 5224
rect 6557 5164 6634 5167
rect 6524 5149 6634 5164
rect 7249 5179 7430 5185
rect 7249 5159 7260 5179
rect 7280 5159 7430 5179
rect 7527 5172 7579 5196
rect 7249 5153 7430 5159
rect 7253 5151 7288 5153
rect 6268 5093 6329 5095
rect 5966 5064 6329 5093
rect 6809 5086 6841 5093
rect 6809 5066 6816 5086
rect 6837 5066 6841 5086
rect 5966 5062 6268 5064
rect 3746 5046 4745 5049
rect 3746 5044 3781 5046
rect 2768 5021 3180 5023
rect 2770 5020 2810 5021
rect 3148 4956 3180 5021
rect 6809 5001 6841 5066
rect 7179 5001 7219 5002
rect 6809 4999 7221 5001
rect 6208 4976 6243 4978
rect 5244 4973 6243 4976
rect 3721 4958 4023 4960
rect 3148 4936 3152 4956
rect 3173 4936 3180 4956
rect 3148 4929 3180 4936
rect 3660 4929 4023 4958
rect 3660 4927 3721 4929
rect 2701 4869 2736 4871
rect 454 4837 531 4840
rect 421 4822 531 4837
rect 1150 4852 1187 4857
rect 1150 4832 1157 4852
rect 1177 4832 1187 4852
rect 1150 4825 1187 4832
rect 1956 4830 1994 4864
rect 2559 4863 2740 4869
rect 2559 4843 2709 4863
rect 2729 4843 2740 4863
rect 2559 4837 2740 4843
rect 3355 4858 3465 4873
rect 3355 4855 3432 4858
rect 2392 4830 2442 4834
rect 1150 4824 1185 4825
rect 187 4724 195 4753
rect 224 4724 235 4753
rect 187 4719 235 4724
rect 706 4759 738 4766
rect 706 4739 713 4759
rect 734 4739 738 4759
rect 706 4674 738 4739
rect 1076 4674 1116 4675
rect 706 4672 1118 4674
rect 706 4646 1086 4672
rect 1112 4646 1118 4672
rect 706 4638 1118 4646
rect 706 4610 738 4638
rect 1151 4618 1185 4824
rect 1956 4820 2442 4830
rect 1467 4798 1578 4820
rect 1467 4778 1475 4798
rect 1494 4778 1552 4798
rect 1571 4778 1578 4798
rect 1956 4788 2405 4820
rect 1467 4761 1578 4778
rect 2392 4767 2405 4788
rect 2436 4767 2442 4820
rect 2392 4750 2442 4767
rect 2089 4691 2123 4692
rect 1220 4656 2124 4691
rect 2332 4681 2379 4699
rect 706 4590 711 4610
rect 732 4590 738 4610
rect 706 4583 738 4590
rect 913 4610 952 4616
rect 913 4590 921 4610
rect 946 4590 952 4610
rect 913 4583 952 4590
rect 1129 4613 1185 4618
rect 1129 4593 1136 4613
rect 1156 4593 1185 4613
rect 1129 4586 1185 4593
rect 1129 4585 1164 4586
rect 921 4537 952 4583
rect 420 4512 531 4534
rect 420 4492 428 4512
rect 447 4492 505 4512
rect 524 4492 531 4512
rect 920 4520 952 4537
rect 1221 4520 1258 4656
rect 1359 4623 1469 4637
rect 1359 4620 1437 4623
rect 1359 4593 1363 4620
rect 1392 4596 1437 4620
rect 1466 4596 1469 4623
rect 2089 4613 2123 4656
rect 1392 4593 1469 4596
rect 1359 4578 1469 4593
rect 2088 4608 2123 4613
rect 2088 4588 2095 4608
rect 2115 4588 2123 4608
rect 2088 4580 2123 4588
rect 920 4507 1258 4520
rect 420 4475 531 4492
rect 921 4488 1258 4507
rect 1200 4487 1258 4488
rect 1644 4515 1676 4522
rect 1644 4495 1651 4515
rect 1672 4495 1676 4515
rect 1644 4430 1676 4495
rect 2014 4430 2054 4431
rect 1644 4428 2056 4430
rect 1644 4402 2024 4428
rect 2050 4402 2056 4428
rect 1644 4394 2056 4402
rect 190 4355 1186 4381
rect 1644 4366 1676 4394
rect 192 4302 234 4355
rect 192 4283 201 4302
rect 226 4283 234 4302
rect 192 4273 234 4283
rect 420 4313 530 4327
rect 420 4310 498 4313
rect 420 4283 424 4310
rect 453 4286 498 4310
rect 527 4286 530 4313
rect 1150 4303 1184 4355
rect 1644 4346 1649 4366
rect 1670 4346 1676 4366
rect 1644 4339 1676 4346
rect 1854 4367 1892 4377
rect 2089 4374 2123 4580
rect 1854 4350 1864 4367
rect 1884 4350 1892 4367
rect 1695 4307 1736 4308
rect 453 4283 530 4286
rect 420 4268 530 4283
rect 1149 4298 1184 4303
rect 1149 4278 1156 4298
rect 1176 4278 1184 4298
rect 1694 4297 1736 4307
rect 1149 4270 1184 4278
rect 705 4205 737 4212
rect 705 4185 712 4205
rect 733 4185 737 4205
rect 705 4120 737 4185
rect 1075 4120 1115 4121
rect 705 4118 1117 4120
rect 705 4092 1085 4118
rect 1111 4092 1117 4118
rect 705 4084 1117 4092
rect 705 4056 737 4084
rect 1150 4064 1184 4270
rect 1358 4268 1469 4290
rect 1358 4248 1366 4268
rect 1385 4248 1443 4268
rect 1462 4248 1469 4268
rect 1358 4231 1469 4248
rect 1694 4275 1701 4297
rect 1727 4275 1736 4297
rect 1694 4266 1736 4275
rect 911 4061 954 4063
rect 705 4036 710 4056
rect 731 4036 737 4056
rect 705 4029 737 4036
rect 910 4054 954 4061
rect 910 4034 920 4054
rect 943 4034 954 4054
rect 910 4030 954 4034
rect 1128 4059 1184 4064
rect 1128 4039 1135 4059
rect 1155 4039 1184 4059
rect 1128 4032 1184 4039
rect 1240 4200 1273 4201
rect 1694 4200 1731 4266
rect 1240 4171 1731 4200
rect 1128 4031 1163 4032
rect 419 3958 530 3980
rect 419 3938 427 3958
rect 446 3938 504 3958
rect 523 3938 530 3958
rect 419 3921 530 3938
rect 910 3949 952 4030
rect 1240 3951 1273 4171
rect 1694 4169 1731 4171
rect 1500 4031 1610 4045
rect 1500 4028 1578 4031
rect 1500 4001 1504 4028
rect 1533 4004 1578 4028
rect 1607 4004 1610 4031
rect 1533 4001 1610 4004
rect 1500 3986 1610 4001
rect 1854 4012 1892 4350
rect 2067 4369 2123 4374
rect 2067 4349 2074 4369
rect 2094 4349 2123 4369
rect 2067 4342 2123 4349
rect 2332 4641 2339 4681
rect 2366 4641 2379 4681
rect 2562 4659 2609 4837
rect 3355 4828 3358 4855
rect 3387 4831 3432 4855
rect 3461 4831 3465 4858
rect 3387 4828 3465 4831
rect 3355 4814 3465 4828
rect 2067 4341 2102 4342
rect 2232 4021 2264 4022
rect 1854 3995 1862 4012
rect 1882 3995 1892 4012
rect 1854 3989 1892 3995
rect 2229 4016 2264 4021
rect 2229 3996 2236 4016
rect 2256 3996 2264 4016
rect 2229 3988 2264 3996
rect 1212 3949 1273 3951
rect 910 3920 1273 3949
rect 1785 3923 1817 3930
rect 910 3918 1212 3920
rect 1785 3903 1792 3923
rect 1813 3903 1817 3923
rect 1785 3838 1817 3903
rect 2155 3838 2195 3839
rect 1785 3836 2197 3838
rect 1153 3832 1188 3834
rect 189 3829 1188 3832
rect 188 3805 1188 3829
rect 188 3650 236 3805
rect 422 3764 532 3778
rect 422 3761 500 3764
rect 422 3734 426 3761
rect 455 3737 500 3761
rect 529 3737 532 3764
rect 1153 3754 1188 3805
rect 455 3734 532 3737
rect 422 3719 532 3734
rect 1151 3749 1188 3754
rect 1151 3729 1158 3749
rect 1178 3729 1188 3749
rect 1785 3810 2165 3836
rect 2191 3810 2197 3836
rect 1785 3802 2197 3810
rect 1785 3774 1817 3802
rect 1785 3754 1790 3774
rect 1811 3754 1817 3774
rect 1785 3747 1817 3754
rect 1991 3773 2033 3784
rect 2230 3782 2264 3988
rect 1991 3752 1998 3773
rect 2025 3752 2033 3773
rect 1151 3722 1188 3729
rect 1151 3721 1186 3722
rect 188 3621 196 3650
rect 225 3621 236 3650
rect 188 3616 236 3621
rect 707 3656 739 3663
rect 707 3636 714 3656
rect 735 3636 739 3656
rect 707 3571 739 3636
rect 1077 3571 1117 3572
rect 707 3569 1119 3571
rect 707 3543 1087 3569
rect 1113 3543 1119 3569
rect 707 3535 1119 3543
rect 707 3507 739 3535
rect 1152 3515 1186 3721
rect 1856 3704 1895 3711
rect 1499 3676 1610 3698
rect 1499 3656 1507 3676
rect 1526 3656 1584 3676
rect 1603 3656 1610 3676
rect 1499 3639 1610 3656
rect 1856 3677 1860 3704
rect 1891 3677 1895 3704
rect 1703 3588 1756 3592
rect 1221 3553 1756 3588
rect 707 3487 712 3507
rect 733 3487 739 3507
rect 707 3480 739 3487
rect 914 3507 953 3513
rect 914 3487 922 3507
rect 947 3487 953 3507
rect 914 3480 953 3487
rect 1130 3510 1186 3515
rect 1130 3490 1137 3510
rect 1157 3490 1186 3510
rect 1130 3483 1186 3490
rect 1130 3482 1165 3483
rect 922 3434 953 3480
rect 421 3409 532 3431
rect 421 3389 429 3409
rect 448 3389 506 3409
rect 525 3389 532 3409
rect 921 3417 953 3434
rect 1222 3417 1259 3553
rect 1360 3520 1470 3534
rect 1360 3517 1438 3520
rect 1360 3490 1364 3517
rect 1393 3493 1438 3517
rect 1467 3493 1470 3520
rect 1393 3490 1470 3493
rect 1360 3475 1470 3490
rect 1702 3506 1756 3553
rect 1702 3498 1755 3506
rect 1702 3481 1711 3498
rect 1743 3481 1755 3498
rect 1702 3478 1755 3481
rect 921 3404 1259 3417
rect 421 3372 532 3389
rect 922 3385 1259 3404
rect 1201 3384 1259 3385
rect 1645 3412 1677 3419
rect 1645 3392 1652 3412
rect 1673 3392 1677 3412
rect 1645 3327 1677 3392
rect 1856 3404 1895 3677
rect 1991 3581 2033 3752
rect 2208 3777 2264 3782
rect 2208 3757 2215 3777
rect 2235 3757 2264 3777
rect 2208 3750 2264 3757
rect 2208 3749 2243 3750
rect 1991 3547 2235 3581
rect 2198 3539 2235 3547
rect 2091 3506 2125 3517
rect 2089 3505 2125 3506
rect 2089 3485 2096 3505
rect 2116 3485 2125 3505
rect 2089 3477 2125 3485
rect 1856 3363 1863 3404
rect 1884 3363 1895 3404
rect 1856 3348 1895 3363
rect 2015 3327 2055 3328
rect 1645 3325 2057 3327
rect 1645 3299 2025 3325
rect 2051 3299 2057 3325
rect 1645 3291 2057 3299
rect 191 3252 1187 3278
rect 1645 3263 1677 3291
rect 2090 3271 2124 3477
rect 193 3199 235 3252
rect 193 3180 202 3199
rect 227 3180 235 3199
rect 193 3170 235 3180
rect 421 3210 531 3224
rect 421 3207 499 3210
rect 421 3180 425 3207
rect 454 3183 499 3207
rect 528 3183 531 3210
rect 1151 3200 1185 3252
rect 1645 3243 1650 3263
rect 1671 3243 1677 3263
rect 1645 3236 1677 3243
rect 2068 3266 2124 3271
rect 2068 3246 2075 3266
rect 2095 3246 2124 3266
rect 2068 3239 2124 3246
rect 2068 3238 2103 3239
rect 1696 3204 1737 3205
rect 454 3180 531 3183
rect 421 3165 531 3180
rect 1150 3195 1185 3200
rect 1150 3175 1157 3195
rect 1177 3175 1185 3195
rect 1695 3194 1737 3204
rect 1150 3167 1185 3175
rect 706 3102 738 3109
rect 706 3082 713 3102
rect 734 3082 738 3102
rect 706 3017 738 3082
rect 1076 3017 1116 3018
rect 706 3015 1118 3017
rect 706 2989 1086 3015
rect 1112 2989 1118 3015
rect 706 2981 1118 2989
rect 706 2953 738 2981
rect 1151 2961 1185 3167
rect 1359 3165 1470 3187
rect 1359 3145 1367 3165
rect 1386 3145 1444 3165
rect 1463 3145 1470 3165
rect 1359 3128 1470 3145
rect 1695 3172 1702 3194
rect 1728 3172 1737 3194
rect 1695 3163 1737 3172
rect 912 2958 955 2960
rect 706 2933 711 2953
rect 732 2933 738 2953
rect 706 2926 738 2933
rect 911 2951 955 2958
rect 911 2931 921 2951
rect 944 2931 955 2951
rect 911 2927 955 2931
rect 1129 2956 1185 2961
rect 1129 2936 1136 2956
rect 1156 2936 1185 2956
rect 1129 2929 1185 2936
rect 1241 3097 1274 3098
rect 1695 3097 1732 3163
rect 2198 3148 2236 3539
rect 1812 3132 2236 3148
rect 1241 3068 1732 3097
rect 1129 2928 1164 2929
rect 420 2855 531 2877
rect 420 2835 428 2855
rect 447 2835 505 2855
rect 524 2835 531 2855
rect 420 2819 531 2835
rect 911 2846 953 2927
rect 1241 2848 1274 3068
rect 1695 3066 1732 3068
rect 1811 3107 2236 3132
rect 1470 2941 1580 2955
rect 1470 2938 1548 2941
rect 1470 2911 1474 2938
rect 1503 2914 1548 2938
rect 1577 2914 1580 2941
rect 1503 2911 1580 2914
rect 1470 2896 1580 2911
rect 1811 2928 1845 3107
rect 2332 3064 2379 4641
rect 2561 4635 2609 4659
rect 3202 4707 3239 4709
rect 3660 4707 3693 4927
rect 3981 4848 4023 4929
rect 4403 4940 4514 4957
rect 4403 4920 4410 4940
rect 4429 4920 4487 4940
rect 4506 4920 4514 4940
rect 4403 4898 4514 4920
rect 5243 4949 6243 4973
rect 3770 4846 3805 4847
rect 3202 4678 3693 4707
rect 2561 3150 2607 4635
rect 3202 4612 3239 4678
rect 3660 4677 3693 4678
rect 3749 4839 3805 4846
rect 3749 4819 3778 4839
rect 3798 4819 3805 4839
rect 3749 4814 3805 4819
rect 3979 4844 4023 4848
rect 3979 4824 3990 4844
rect 4013 4824 4023 4844
rect 3979 4817 4023 4824
rect 4196 4842 4228 4849
rect 4196 4822 4202 4842
rect 4223 4822 4228 4842
rect 3979 4815 4022 4817
rect 3197 4603 3239 4612
rect 3197 4581 3206 4603
rect 3232 4581 3239 4603
rect 3464 4630 3575 4647
rect 3464 4610 3471 4630
rect 3490 4610 3548 4630
rect 3567 4610 3575 4630
rect 3464 4588 3575 4610
rect 3749 4608 3783 4814
rect 4196 4794 4228 4822
rect 3816 4786 4228 4794
rect 3816 4760 3822 4786
rect 3848 4760 4228 4786
rect 5243 4794 5291 4949
rect 5477 4908 5587 4922
rect 5477 4905 5555 4908
rect 5477 4878 5481 4905
rect 5510 4881 5555 4905
rect 5584 4881 5587 4908
rect 6208 4898 6243 4949
rect 6809 4973 7189 4999
rect 7215 4973 7221 4999
rect 6809 4965 7221 4973
rect 6809 4937 6841 4965
rect 7254 4945 7288 5151
rect 7778 5150 7813 5151
rect 6809 4917 6814 4937
rect 6835 4917 6841 4937
rect 6809 4910 6841 4917
rect 7011 4940 7056 4945
rect 7011 4916 7022 4940
rect 7048 4916 7056 4940
rect 7011 4905 7056 4916
rect 7232 4940 7288 4945
rect 7232 4920 7239 4940
rect 7259 4920 7288 4940
rect 7232 4913 7288 4920
rect 7757 5143 7813 5150
rect 7757 5123 7786 5143
rect 7806 5123 7813 5143
rect 7757 5118 7813 5123
rect 7982 5146 8027 5225
rect 8411 5244 8522 5261
rect 8411 5224 8418 5244
rect 8437 5224 8495 5244
rect 8514 5224 8522 5244
rect 8411 5202 8522 5224
rect 8804 5198 8838 5404
rect 9251 5384 9283 5412
rect 8871 5376 9283 5384
rect 10223 5410 10265 5463
rect 10223 5391 10232 5410
rect 10257 5391 10265 5410
rect 10223 5381 10265 5391
rect 10451 5421 10561 5435
rect 10451 5418 10529 5421
rect 10451 5391 10455 5418
rect 10484 5394 10529 5418
rect 10558 5394 10561 5421
rect 11181 5411 11215 5463
rect 11675 5454 11680 5474
rect 11701 5454 11707 5474
rect 11675 5447 11707 5454
rect 12098 5477 12154 5482
rect 12098 5457 12105 5477
rect 12125 5457 12154 5477
rect 12098 5450 12154 5457
rect 12098 5449 12133 5450
rect 11726 5415 11767 5416
rect 10484 5391 10561 5394
rect 10451 5376 10561 5391
rect 11180 5406 11215 5411
rect 11180 5386 11187 5406
rect 11207 5386 11215 5406
rect 11725 5405 11767 5415
rect 11180 5378 11215 5386
rect 8871 5350 8877 5376
rect 8903 5350 9283 5376
rect 8871 5348 9283 5350
rect 8873 5347 8913 5348
rect 9251 5283 9283 5348
rect 10736 5313 10768 5320
rect 9251 5263 9255 5283
rect 9276 5263 9283 5283
rect 9251 5256 9283 5263
rect 9754 5298 9802 5303
rect 9754 5269 9765 5298
rect 9794 5269 9802 5298
rect 8804 5197 8839 5198
rect 8802 5190 8839 5197
rect 8802 5170 8812 5190
rect 8832 5170 8839 5190
rect 8802 5165 8839 5170
rect 9458 5185 9568 5200
rect 9458 5182 9535 5185
rect 7982 5126 7993 5146
rect 8018 5126 8027 5146
rect 7982 5122 8027 5126
rect 8204 5146 8236 5153
rect 8204 5126 8210 5146
rect 8231 5126 8236 5146
rect 7232 4912 7267 4913
rect 7757 4912 7791 5118
rect 8204 5098 8236 5126
rect 7824 5090 8236 5098
rect 7824 5064 7830 5090
rect 7856 5064 8236 5090
rect 8802 5114 8837 5165
rect 9458 5155 9461 5182
rect 9490 5158 9535 5182
rect 9564 5158 9568 5185
rect 9490 5155 9568 5158
rect 9458 5141 9568 5155
rect 9754 5114 9802 5269
rect 10736 5293 10743 5313
rect 10764 5293 10768 5313
rect 10736 5228 10768 5293
rect 11106 5228 11146 5229
rect 10736 5226 11148 5228
rect 10736 5200 11116 5226
rect 11142 5200 11148 5226
rect 10736 5192 11148 5200
rect 10736 5164 10768 5192
rect 11181 5172 11215 5378
rect 11389 5376 11500 5398
rect 11389 5356 11397 5376
rect 11416 5356 11474 5376
rect 11493 5356 11500 5376
rect 11389 5339 11500 5356
rect 11725 5383 11732 5405
rect 11758 5383 11767 5405
rect 11725 5374 11767 5383
rect 10942 5169 10985 5171
rect 10736 5144 10741 5164
rect 10762 5144 10768 5164
rect 10736 5137 10768 5144
rect 10941 5162 10985 5169
rect 10941 5142 10951 5162
rect 10974 5142 10985 5162
rect 10941 5138 10985 5142
rect 11159 5167 11215 5172
rect 11159 5147 11166 5167
rect 11186 5147 11215 5167
rect 11159 5140 11215 5147
rect 11271 5308 11304 5309
rect 11725 5308 11762 5374
rect 12357 5351 12403 6836
rect 11271 5279 11762 5308
rect 11159 5139 11194 5140
rect 8802 5090 9802 5114
rect 8802 5087 9801 5090
rect 8802 5085 8837 5087
rect 7824 5062 8236 5064
rect 7826 5061 7866 5062
rect 8204 4997 8236 5062
rect 10450 5066 10561 5088
rect 10450 5046 10458 5066
rect 10477 5046 10535 5066
rect 10554 5046 10561 5066
rect 10450 5029 10561 5046
rect 10941 5057 10983 5138
rect 11271 5059 11304 5279
rect 11725 5277 11762 5279
rect 12355 5327 12403 5351
rect 12585 5345 12632 6922
rect 13119 6879 13153 7058
rect 13384 7075 13494 7090
rect 13384 7072 13461 7075
rect 13384 7045 13387 7072
rect 13416 7048 13461 7072
rect 13490 7048 13494 7075
rect 13416 7045 13494 7048
rect 13384 7031 13494 7045
rect 12728 6854 13153 6879
rect 13232 6918 13269 6920
rect 13690 6918 13723 7138
rect 14011 7059 14053 7140
rect 14433 7151 14544 7167
rect 14433 7131 14440 7151
rect 14459 7131 14517 7151
rect 14536 7131 14544 7151
rect 14433 7109 14544 7131
rect 15273 7160 16273 7184
rect 13800 7057 13835 7058
rect 13232 6889 13723 6918
rect 12728 6838 13152 6854
rect 12728 6447 12766 6838
rect 13232 6823 13269 6889
rect 13690 6888 13723 6889
rect 13779 7050 13835 7057
rect 13779 7030 13808 7050
rect 13828 7030 13835 7050
rect 13779 7025 13835 7030
rect 14009 7055 14053 7059
rect 14009 7035 14020 7055
rect 14043 7035 14053 7055
rect 14009 7028 14053 7035
rect 14226 7053 14258 7060
rect 14226 7033 14232 7053
rect 14253 7033 14258 7053
rect 14009 7026 14052 7028
rect 13227 6814 13269 6823
rect 13227 6792 13236 6814
rect 13262 6792 13269 6814
rect 13494 6841 13605 6858
rect 13494 6821 13501 6841
rect 13520 6821 13578 6841
rect 13597 6821 13605 6841
rect 13494 6799 13605 6821
rect 13779 6819 13813 7025
rect 14226 7005 14258 7033
rect 13846 6997 14258 7005
rect 13846 6971 13852 6997
rect 13878 6971 14258 6997
rect 15273 7005 15321 7160
rect 15507 7119 15617 7133
rect 15507 7116 15585 7119
rect 15507 7089 15511 7116
rect 15540 7092 15585 7116
rect 15614 7092 15617 7119
rect 16238 7109 16273 7160
rect 16840 7178 17220 7204
rect 17246 7178 17252 7204
rect 16840 7170 17252 7178
rect 16840 7142 16872 7170
rect 16840 7122 16845 7142
rect 16866 7122 16872 7142
rect 16840 7115 16872 7122
rect 17046 7141 17091 7153
rect 17285 7150 17319 7356
rect 17046 7122 17053 7141
rect 17082 7122 17091 7141
rect 15540 7089 15617 7092
rect 15507 7074 15617 7089
rect 16236 7104 16273 7109
rect 16236 7084 16243 7104
rect 16263 7084 16273 7104
rect 16236 7077 16273 7084
rect 16236 7076 16271 7077
rect 15273 6976 15281 7005
rect 15310 6976 15321 7005
rect 15273 6971 15321 6976
rect 15792 7011 15824 7018
rect 15792 6991 15799 7011
rect 15820 6991 15824 7011
rect 13846 6969 14258 6971
rect 13848 6968 13888 6969
rect 14226 6904 14258 6969
rect 14226 6884 14230 6904
rect 14251 6884 14258 6904
rect 14226 6877 14258 6884
rect 15792 6926 15824 6991
rect 16162 6926 16202 6927
rect 15792 6924 16204 6926
rect 15792 6898 16172 6924
rect 16198 6898 16204 6924
rect 15792 6890 16204 6898
rect 15792 6862 15824 6890
rect 16237 6870 16271 7076
rect 16554 7044 16665 7066
rect 16554 7024 16562 7044
rect 16581 7024 16639 7044
rect 16658 7024 16665 7044
rect 16554 7007 16665 7024
rect 17046 7039 17091 7122
rect 17263 7145 17319 7150
rect 17263 7125 17270 7145
rect 17290 7125 17319 7145
rect 17786 7340 17815 7360
rect 17835 7340 17842 7360
rect 17786 7335 17842 7340
rect 18233 7363 18265 7370
rect 18233 7343 18239 7363
rect 18260 7343 18265 7363
rect 17786 7129 17820 7335
rect 18233 7315 18265 7343
rect 17853 7307 18265 7315
rect 17853 7281 17859 7307
rect 17885 7281 18265 7307
rect 18832 7325 18867 7376
rect 19488 7366 19491 7393
rect 19520 7369 19565 7393
rect 19594 7369 19598 7396
rect 19520 7366 19598 7369
rect 19488 7352 19598 7366
rect 19784 7325 19832 7480
rect 18832 7301 19832 7325
rect 18832 7298 19831 7301
rect 18832 7296 18867 7298
rect 17853 7279 18265 7281
rect 17855 7278 17895 7279
rect 18021 7238 18056 7256
rect 18021 7206 18024 7238
rect 18051 7206 18056 7238
rect 17786 7128 17821 7129
rect 17263 7118 17319 7125
rect 17784 7121 17822 7128
rect 17263 7117 17298 7118
rect 17784 7117 17794 7121
rect 17778 7103 17794 7117
rect 17814 7117 17822 7121
rect 17814 7103 17828 7117
rect 17778 7096 17828 7103
rect 17411 7039 17461 7041
rect 17046 7005 17461 7039
rect 17175 6943 17209 6944
rect 16306 6908 17210 6943
rect 17258 6932 17326 6943
rect 17258 6911 17263 6932
rect 15792 6842 15797 6862
rect 15818 6842 15824 6862
rect 15792 6835 15824 6842
rect 15999 6862 16038 6868
rect 15999 6842 16007 6862
rect 16032 6842 16038 6862
rect 15999 6835 16038 6842
rect 16215 6865 16271 6870
rect 16215 6845 16222 6865
rect 16242 6845 16271 6865
rect 16215 6838 16271 6845
rect 16215 6837 16250 6838
rect 13779 6811 13814 6819
rect 13227 6782 13269 6792
rect 13779 6791 13787 6811
rect 13807 6791 13814 6811
rect 13779 6786 13814 6791
rect 14433 6806 14543 6821
rect 14433 6803 14510 6806
rect 13227 6781 13268 6782
rect 12861 6747 12896 6748
rect 12840 6740 12896 6747
rect 12840 6720 12869 6740
rect 12889 6720 12896 6740
rect 12840 6715 12896 6720
rect 13287 6743 13319 6750
rect 13287 6723 13293 6743
rect 13314 6723 13319 6743
rect 13779 6734 13813 6786
rect 14433 6776 14436 6803
rect 14465 6779 14510 6803
rect 14539 6779 14543 6806
rect 14465 6776 14543 6779
rect 14433 6762 14543 6776
rect 14729 6806 14771 6816
rect 14729 6787 14737 6806
rect 14762 6787 14771 6806
rect 16007 6789 16038 6835
rect 14729 6734 14771 6787
rect 15506 6764 15617 6786
rect 15506 6744 15514 6764
rect 15533 6744 15591 6764
rect 15610 6744 15617 6764
rect 16006 6772 16038 6789
rect 16307 6772 16344 6908
rect 16445 6875 16555 6889
rect 16445 6872 16523 6875
rect 16445 6845 16449 6872
rect 16478 6848 16523 6872
rect 16552 6848 16555 6875
rect 17175 6865 17209 6908
rect 16478 6845 16555 6848
rect 16445 6830 16555 6845
rect 17174 6860 17209 6865
rect 17174 6840 17181 6860
rect 17201 6840 17209 6860
rect 17174 6832 17209 6840
rect 16006 6759 16344 6772
rect 12840 6509 12874 6715
rect 13287 6695 13319 6723
rect 13777 6708 14773 6734
rect 15506 6727 15617 6744
rect 16007 6740 16344 6759
rect 16286 6739 16344 6740
rect 16730 6767 16762 6774
rect 16730 6747 16737 6767
rect 16758 6747 16762 6767
rect 12907 6687 13319 6695
rect 12907 6661 12913 6687
rect 12939 6661 13319 6687
rect 12907 6659 13319 6661
rect 12909 6658 12949 6659
rect 13069 6623 13108 6638
rect 13069 6582 13080 6623
rect 13101 6582 13108 6623
rect 12839 6501 12875 6509
rect 12839 6481 12848 6501
rect 12868 6481 12875 6501
rect 12839 6480 12875 6481
rect 12839 6469 12873 6480
rect 12729 6439 12766 6447
rect 12729 6405 12973 6439
rect 12721 6236 12756 6237
rect 12700 6229 12756 6236
rect 12700 6209 12729 6229
rect 12749 6209 12756 6229
rect 12700 6204 12756 6209
rect 12931 6234 12973 6405
rect 13069 6309 13108 6582
rect 13287 6594 13319 6659
rect 16730 6682 16762 6747
rect 17100 6682 17140 6683
rect 16730 6680 17142 6682
rect 16730 6654 17110 6680
rect 17136 6654 17142 6680
rect 16730 6646 17142 6654
rect 13287 6574 13291 6594
rect 13312 6574 13319 6594
rect 13287 6567 13319 6574
rect 13705 6601 13763 6602
rect 13705 6582 14042 6601
rect 14432 6597 14543 6614
rect 15276 6607 16272 6633
rect 16730 6618 16762 6646
rect 13705 6569 14043 6582
rect 13209 6505 13262 6508
rect 13209 6488 13221 6505
rect 13253 6488 13262 6505
rect 13209 6480 13262 6488
rect 13208 6433 13262 6480
rect 13494 6496 13604 6511
rect 13494 6493 13571 6496
rect 13494 6466 13497 6493
rect 13526 6469 13571 6493
rect 13600 6469 13604 6496
rect 13526 6466 13604 6469
rect 13494 6452 13604 6466
rect 13705 6433 13742 6569
rect 14011 6552 14043 6569
rect 14432 6577 14439 6597
rect 14458 6577 14516 6597
rect 14535 6577 14543 6597
rect 14432 6555 14543 6577
rect 15278 6554 15320 6607
rect 14011 6506 14042 6552
rect 15278 6535 15287 6554
rect 15312 6535 15320 6554
rect 15278 6525 15320 6535
rect 15506 6565 15616 6579
rect 15506 6562 15584 6565
rect 15506 6535 15510 6562
rect 15539 6538 15584 6562
rect 15613 6538 15616 6565
rect 16236 6555 16270 6607
rect 16730 6598 16735 6618
rect 16756 6598 16762 6618
rect 16730 6591 16762 6598
rect 16940 6619 16978 6629
rect 17175 6626 17209 6832
rect 16940 6602 16950 6619
rect 16970 6602 16978 6619
rect 16781 6559 16822 6560
rect 15539 6535 15616 6538
rect 15506 6520 15616 6535
rect 16235 6550 16270 6555
rect 16235 6530 16242 6550
rect 16262 6530 16270 6550
rect 16780 6549 16822 6559
rect 16235 6522 16270 6530
rect 13799 6503 13834 6504
rect 13778 6496 13834 6503
rect 13778 6476 13807 6496
rect 13827 6476 13834 6496
rect 13778 6471 13834 6476
rect 14011 6499 14050 6506
rect 14011 6479 14017 6499
rect 14042 6479 14050 6499
rect 14011 6473 14050 6479
rect 14225 6499 14257 6506
rect 14225 6479 14231 6499
rect 14252 6479 14257 6499
rect 13208 6398 13743 6433
rect 13208 6394 13261 6398
rect 13069 6282 13073 6309
rect 13104 6282 13108 6309
rect 13354 6330 13465 6347
rect 13354 6310 13361 6330
rect 13380 6310 13438 6330
rect 13457 6310 13465 6330
rect 13354 6288 13465 6310
rect 13069 6275 13108 6282
rect 13778 6265 13812 6471
rect 14225 6451 14257 6479
rect 13845 6443 14257 6451
rect 13845 6417 13851 6443
rect 13877 6417 14257 6443
rect 13845 6415 14257 6417
rect 13847 6414 13887 6415
rect 14225 6350 14257 6415
rect 15791 6457 15823 6464
rect 15791 6437 15798 6457
rect 15819 6437 15823 6457
rect 15791 6372 15823 6437
rect 16161 6372 16201 6373
rect 15791 6370 16203 6372
rect 14225 6330 14229 6350
rect 14250 6330 14257 6350
rect 14225 6323 14257 6330
rect 14728 6365 14776 6370
rect 14728 6336 14739 6365
rect 14768 6336 14776 6365
rect 13778 6264 13813 6265
rect 13776 6257 13813 6264
rect 12931 6213 12939 6234
rect 12966 6213 12973 6234
rect 12700 5998 12734 6204
rect 12931 6202 12973 6213
rect 13147 6232 13179 6239
rect 13147 6212 13153 6232
rect 13174 6212 13179 6232
rect 13147 6184 13179 6212
rect 12767 6176 13179 6184
rect 12767 6150 12773 6176
rect 12799 6150 13179 6176
rect 13776 6237 13786 6257
rect 13806 6237 13813 6257
rect 13776 6232 13813 6237
rect 14432 6252 14542 6267
rect 14432 6249 14509 6252
rect 13776 6181 13811 6232
rect 14432 6222 14435 6249
rect 14464 6225 14509 6249
rect 14538 6225 14542 6252
rect 14464 6222 14542 6225
rect 14432 6208 14542 6222
rect 14728 6181 14776 6336
rect 15791 6344 16171 6370
rect 16197 6344 16203 6370
rect 15791 6336 16203 6344
rect 15791 6308 15823 6336
rect 16236 6316 16270 6522
rect 16444 6520 16555 6542
rect 16444 6500 16452 6520
rect 16471 6500 16529 6520
rect 16548 6500 16555 6520
rect 16444 6483 16555 6500
rect 16780 6527 16787 6549
rect 16813 6527 16822 6549
rect 16780 6518 16822 6527
rect 15997 6313 16040 6315
rect 15791 6288 15796 6308
rect 15817 6288 15823 6308
rect 15791 6281 15823 6288
rect 15996 6306 16040 6313
rect 15996 6286 16006 6306
rect 16029 6286 16040 6306
rect 15996 6282 16040 6286
rect 16214 6311 16270 6316
rect 16214 6291 16221 6311
rect 16241 6291 16270 6311
rect 16214 6284 16270 6291
rect 16326 6452 16359 6453
rect 16780 6452 16817 6518
rect 16326 6423 16817 6452
rect 16214 6283 16249 6284
rect 13776 6157 14776 6181
rect 15505 6210 15616 6232
rect 15505 6190 15513 6210
rect 15532 6190 15590 6210
rect 15609 6190 15616 6210
rect 15505 6173 15616 6190
rect 15996 6201 16038 6282
rect 16326 6203 16359 6423
rect 16780 6421 16817 6423
rect 16586 6283 16696 6297
rect 16586 6280 16664 6283
rect 16586 6253 16590 6280
rect 16619 6256 16664 6280
rect 16693 6256 16696 6283
rect 16619 6253 16696 6256
rect 16586 6238 16696 6253
rect 16940 6264 16978 6602
rect 17153 6621 17209 6626
rect 17153 6601 17160 6621
rect 17180 6601 17209 6621
rect 17153 6594 17209 6601
rect 17256 6903 17263 6911
rect 17311 6903 17326 6932
rect 17256 6894 17326 6903
rect 17153 6593 17188 6594
rect 17075 6493 17119 6497
rect 17256 6493 17306 6894
rect 17411 6877 17461 7005
rect 17644 7018 17754 7020
rect 18021 7018 18056 7206
rect 18233 7214 18265 7279
rect 18233 7194 18237 7214
rect 18258 7194 18265 7214
rect 18807 7210 19109 7212
rect 18233 7187 18265 7194
rect 18746 7181 19109 7210
rect 18746 7179 18807 7181
rect 17644 6988 18056 7018
rect 17644 6963 17688 6988
rect 17727 6985 18056 6988
rect 18175 7119 18209 7125
rect 18175 7099 18184 7119
rect 18205 7099 18209 7119
rect 17075 6460 17306 6493
rect 17075 6458 17282 6460
rect 17075 6304 17119 6458
rect 16940 6247 16948 6264
rect 16968 6247 16978 6264
rect 16940 6241 16978 6247
rect 16298 6201 16359 6203
rect 15996 6172 16359 6201
rect 16871 6175 16903 6182
rect 15996 6170 16298 6172
rect 13776 6154 14775 6157
rect 16871 6155 16878 6175
rect 16899 6155 16903 6175
rect 13776 6152 13811 6154
rect 12767 6148 13179 6150
rect 12769 6147 12809 6148
rect 13147 6083 13179 6148
rect 16871 6090 16903 6155
rect 17081 6168 17119 6304
rect 17318 6273 17349 6274
rect 17315 6268 17349 6273
rect 17315 6248 17322 6268
rect 17342 6248 17349 6268
rect 17315 6240 17349 6248
rect 17081 6130 17087 6168
rect 17110 6130 17119 6168
rect 17081 6120 17119 6130
rect 17316 6182 17349 6240
rect 17241 6090 17281 6091
rect 16871 6088 17283 6090
rect 16239 6084 16274 6086
rect 13147 6063 13151 6083
rect 13172 6063 13179 6083
rect 15275 6081 16274 6084
rect 13752 6066 14054 6068
rect 13147 6056 13179 6063
rect 13691 6037 14054 6066
rect 13691 6035 13752 6037
rect 12700 5990 12735 5998
rect 12700 5970 12708 5990
rect 12728 5970 12735 5990
rect 12700 5965 12735 5970
rect 13072 5991 13110 5997
rect 13072 5974 13082 5991
rect 13102 5974 13110 5991
rect 12700 5964 12732 5965
rect 12862 5644 12897 5645
rect 11499 5158 11609 5172
rect 11499 5155 11577 5158
rect 11499 5128 11503 5155
rect 11532 5131 11577 5155
rect 11606 5131 11609 5158
rect 12355 5149 12402 5327
rect 12585 5305 12598 5345
rect 12625 5305 12632 5345
rect 12841 5637 12897 5644
rect 12841 5617 12870 5637
rect 12890 5617 12897 5637
rect 12841 5612 12897 5617
rect 13072 5636 13110 5974
rect 13354 5985 13464 6000
rect 13354 5982 13431 5985
rect 13354 5955 13357 5982
rect 13386 5958 13431 5982
rect 13460 5958 13464 5985
rect 13386 5955 13464 5958
rect 13354 5941 13464 5955
rect 13233 5815 13270 5817
rect 13691 5815 13724 6035
rect 14012 5956 14054 6037
rect 14434 6048 14545 6065
rect 14434 6028 14441 6048
rect 14460 6028 14518 6048
rect 14537 6028 14545 6048
rect 14434 6006 14545 6028
rect 15274 6057 16274 6081
rect 13801 5954 13836 5955
rect 13233 5786 13724 5815
rect 13233 5720 13270 5786
rect 13691 5785 13724 5786
rect 13780 5947 13836 5954
rect 13780 5927 13809 5947
rect 13829 5927 13836 5947
rect 13780 5922 13836 5927
rect 14010 5952 14054 5956
rect 14010 5932 14021 5952
rect 14044 5932 14054 5952
rect 14010 5925 14054 5932
rect 14227 5950 14259 5957
rect 14227 5930 14233 5950
rect 14254 5930 14259 5950
rect 14010 5923 14053 5925
rect 13228 5711 13270 5720
rect 13228 5689 13237 5711
rect 13263 5689 13270 5711
rect 13495 5738 13606 5755
rect 13495 5718 13502 5738
rect 13521 5718 13579 5738
rect 13598 5718 13606 5738
rect 13495 5696 13606 5718
rect 13780 5716 13814 5922
rect 14227 5902 14259 5930
rect 13847 5894 14259 5902
rect 13847 5868 13853 5894
rect 13879 5868 14259 5894
rect 15274 5902 15322 6057
rect 15508 6016 15618 6030
rect 15508 6013 15586 6016
rect 15508 5986 15512 6013
rect 15541 5989 15586 6013
rect 15615 5989 15618 6016
rect 16239 6006 16274 6057
rect 15541 5986 15618 5989
rect 15508 5971 15618 5986
rect 16237 6001 16274 6006
rect 16237 5981 16244 6001
rect 16264 5981 16274 6001
rect 16871 6062 17251 6088
rect 17277 6062 17283 6088
rect 16871 6054 17283 6062
rect 16871 6026 16903 6054
rect 17316 6034 17352 6182
rect 16871 6006 16876 6026
rect 16897 6006 16903 6026
rect 16871 5999 16903 6006
rect 17294 6029 17352 6034
rect 17294 6009 17301 6029
rect 17321 6009 17352 6029
rect 17294 6002 17352 6009
rect 17294 6001 17329 6002
rect 16237 5974 16274 5981
rect 16237 5973 16272 5974
rect 15274 5873 15282 5902
rect 15311 5873 15322 5902
rect 15274 5868 15322 5873
rect 15793 5908 15825 5915
rect 15793 5888 15800 5908
rect 15821 5888 15825 5908
rect 13847 5866 14259 5868
rect 13849 5865 13889 5866
rect 14227 5801 14259 5866
rect 14227 5781 14231 5801
rect 14252 5781 14259 5801
rect 14227 5774 14259 5781
rect 15793 5823 15825 5888
rect 16163 5823 16203 5824
rect 15793 5821 16205 5823
rect 15793 5795 16173 5821
rect 16199 5795 16205 5821
rect 15793 5787 16205 5795
rect 15793 5759 15825 5787
rect 16238 5767 16272 5973
rect 16942 5956 16981 5963
rect 16585 5928 16696 5950
rect 16585 5908 16593 5928
rect 16612 5908 16670 5928
rect 16689 5908 16696 5928
rect 16585 5891 16696 5908
rect 16942 5929 16946 5956
rect 16977 5929 16981 5956
rect 16789 5840 16842 5844
rect 16307 5805 16842 5840
rect 15793 5739 15798 5759
rect 15819 5739 15825 5759
rect 15793 5732 15825 5739
rect 16000 5759 16039 5765
rect 16000 5739 16008 5759
rect 16033 5739 16039 5759
rect 16000 5732 16039 5739
rect 16216 5762 16272 5767
rect 16216 5742 16223 5762
rect 16243 5742 16272 5762
rect 16216 5735 16272 5742
rect 16216 5734 16251 5735
rect 13780 5708 13815 5716
rect 13228 5679 13270 5689
rect 13780 5688 13788 5708
rect 13808 5688 13815 5708
rect 13780 5683 13815 5688
rect 14434 5703 14544 5718
rect 14434 5700 14511 5703
rect 13228 5678 13269 5679
rect 13072 5619 13080 5636
rect 13100 5619 13110 5636
rect 12841 5406 12875 5612
rect 13072 5609 13110 5619
rect 13288 5640 13320 5647
rect 13288 5620 13294 5640
rect 13315 5620 13320 5640
rect 13780 5631 13814 5683
rect 14434 5673 14437 5700
rect 14466 5676 14511 5700
rect 14540 5676 14544 5703
rect 14466 5673 14544 5676
rect 14434 5659 14544 5673
rect 14730 5703 14772 5713
rect 14730 5684 14738 5703
rect 14763 5684 14772 5703
rect 16008 5686 16039 5732
rect 14730 5631 14772 5684
rect 15507 5661 15618 5683
rect 15507 5641 15515 5661
rect 15534 5641 15592 5661
rect 15611 5641 15618 5661
rect 16007 5669 16039 5686
rect 16308 5669 16345 5805
rect 16446 5772 16556 5786
rect 16446 5769 16524 5772
rect 16446 5742 16450 5769
rect 16479 5745 16524 5769
rect 16553 5745 16556 5772
rect 16479 5742 16556 5745
rect 16446 5727 16556 5742
rect 16788 5758 16842 5805
rect 16788 5750 16841 5758
rect 16788 5733 16797 5750
rect 16829 5733 16841 5750
rect 16788 5730 16841 5733
rect 16007 5656 16345 5669
rect 13288 5592 13320 5620
rect 13778 5605 14774 5631
rect 15507 5624 15618 5641
rect 16008 5637 16345 5656
rect 16287 5636 16345 5637
rect 16731 5664 16763 5671
rect 16731 5644 16738 5664
rect 16759 5644 16763 5664
rect 12908 5584 13320 5592
rect 12908 5558 12914 5584
rect 12940 5558 13320 5584
rect 12908 5556 13320 5558
rect 12910 5555 12950 5556
rect 13288 5491 13320 5556
rect 16731 5579 16763 5644
rect 16942 5656 16981 5929
rect 17177 5758 17211 5769
rect 17175 5757 17211 5758
rect 17175 5737 17182 5757
rect 17202 5737 17211 5757
rect 17175 5729 17211 5737
rect 16942 5615 16949 5656
rect 16970 5615 16981 5656
rect 16942 5600 16981 5615
rect 17101 5579 17141 5580
rect 16731 5577 17143 5579
rect 16731 5551 17111 5577
rect 17137 5551 17143 5577
rect 16731 5543 17143 5551
rect 13288 5471 13292 5491
rect 13313 5471 13320 5491
rect 13288 5464 13320 5471
rect 13706 5498 13764 5499
rect 13706 5479 14043 5498
rect 14433 5494 14544 5511
rect 15277 5504 16273 5530
rect 16731 5515 16763 5543
rect 17176 5523 17210 5729
rect 13706 5466 14044 5479
rect 12841 5398 12876 5406
rect 12841 5378 12849 5398
rect 12869 5378 12876 5398
rect 12841 5373 12876 5378
rect 13495 5393 13605 5408
rect 13495 5390 13572 5393
rect 12841 5330 12875 5373
rect 13495 5363 13498 5390
rect 13527 5366 13572 5390
rect 13601 5366 13605 5393
rect 13527 5363 13605 5366
rect 13495 5349 13605 5363
rect 13706 5330 13743 5466
rect 14012 5449 14044 5466
rect 14433 5474 14440 5494
rect 14459 5474 14517 5494
rect 14536 5474 14544 5494
rect 14433 5452 14544 5474
rect 15279 5451 15321 5504
rect 14012 5403 14043 5449
rect 15279 5432 15288 5451
rect 15313 5432 15321 5451
rect 15279 5422 15321 5432
rect 15507 5462 15617 5476
rect 15507 5459 15585 5462
rect 15507 5432 15511 5459
rect 15540 5435 15585 5459
rect 15614 5435 15617 5462
rect 16237 5452 16271 5504
rect 16731 5495 16736 5515
rect 16757 5495 16763 5515
rect 16731 5488 16763 5495
rect 17154 5518 17210 5523
rect 17154 5498 17161 5518
rect 17181 5498 17210 5518
rect 17154 5491 17210 5498
rect 17154 5490 17189 5491
rect 16782 5456 16823 5457
rect 15540 5432 15617 5435
rect 15507 5417 15617 5432
rect 16236 5447 16271 5452
rect 16236 5427 16243 5447
rect 16263 5427 16271 5447
rect 16781 5446 16823 5456
rect 16236 5419 16271 5427
rect 13800 5400 13835 5401
rect 13779 5393 13835 5400
rect 13779 5373 13808 5393
rect 13828 5373 13835 5393
rect 13779 5368 13835 5373
rect 14012 5396 14051 5403
rect 14012 5376 14018 5396
rect 14043 5376 14051 5396
rect 14012 5370 14051 5376
rect 14226 5396 14258 5403
rect 14226 5376 14232 5396
rect 14253 5376 14258 5396
rect 12585 5287 12632 5305
rect 12840 5295 13744 5330
rect 12841 5294 12875 5295
rect 12502 5228 12554 5233
rect 12957 5228 13002 5230
rect 12502 5213 13002 5228
rect 12502 5160 12516 5213
rect 12547 5189 13002 5213
rect 12547 5188 12572 5189
rect 12547 5160 12554 5188
rect 11532 5128 11609 5131
rect 11499 5113 11609 5128
rect 12224 5143 12405 5149
rect 12224 5123 12235 5143
rect 12255 5123 12405 5143
rect 12502 5136 12554 5160
rect 12224 5117 12405 5123
rect 12228 5115 12263 5117
rect 11243 5057 11304 5059
rect 10941 5028 11304 5057
rect 11784 5050 11816 5057
rect 11784 5030 11791 5050
rect 11812 5030 11816 5050
rect 10941 5026 11243 5028
rect 8777 4999 9079 5001
rect 8204 4977 8208 4997
rect 8229 4977 8236 4997
rect 8204 4970 8236 4977
rect 8716 4970 9079 4999
rect 8716 4968 8777 4970
rect 7757 4910 7792 4912
rect 5510 4878 5587 4881
rect 5477 4863 5587 4878
rect 6206 4893 6243 4898
rect 6206 4873 6213 4893
rect 6233 4873 6243 4893
rect 6206 4866 6243 4873
rect 7012 4871 7050 4905
rect 7615 4904 7796 4910
rect 7615 4884 7765 4904
rect 7785 4884 7796 4904
rect 7615 4878 7796 4884
rect 8411 4899 8521 4914
rect 8411 4896 8488 4899
rect 7448 4871 7498 4875
rect 6206 4865 6241 4866
rect 5243 4765 5251 4794
rect 5280 4765 5291 4794
rect 5243 4760 5291 4765
rect 5762 4800 5794 4807
rect 5762 4780 5769 4800
rect 5790 4780 5794 4800
rect 3816 4758 4228 4760
rect 3818 4757 3858 4758
rect 4196 4693 4228 4758
rect 4196 4673 4200 4693
rect 4221 4673 4228 4693
rect 4196 4666 4228 4673
rect 5762 4715 5794 4780
rect 6132 4715 6172 4716
rect 5762 4713 6174 4715
rect 5762 4687 6142 4713
rect 6168 4687 6174 4713
rect 5762 4679 6174 4687
rect 5762 4651 5794 4679
rect 6207 4659 6241 4865
rect 7012 4861 7498 4871
rect 6523 4839 6634 4861
rect 6523 4819 6531 4839
rect 6550 4819 6608 4839
rect 6627 4819 6634 4839
rect 7012 4829 7461 4861
rect 6523 4802 6634 4819
rect 7448 4808 7461 4829
rect 7492 4808 7498 4861
rect 7448 4791 7498 4808
rect 7145 4732 7179 4733
rect 6276 4697 7180 4732
rect 7388 4722 7435 4740
rect 5762 4631 5767 4651
rect 5788 4631 5794 4651
rect 5762 4624 5794 4631
rect 5969 4651 6008 4657
rect 5969 4631 5977 4651
rect 6002 4631 6008 4651
rect 5969 4624 6008 4631
rect 6185 4654 6241 4659
rect 6185 4634 6192 4654
rect 6212 4634 6241 4654
rect 6185 4627 6241 4634
rect 6185 4626 6220 4627
rect 3749 4600 3784 4608
rect 3197 4571 3239 4581
rect 3749 4580 3757 4600
rect 3777 4580 3784 4600
rect 3749 4575 3784 4580
rect 4403 4595 4513 4610
rect 4403 4592 4480 4595
rect 3197 4570 3238 4571
rect 2831 4536 2866 4537
rect 2810 4529 2866 4536
rect 2810 4509 2839 4529
rect 2859 4509 2866 4529
rect 2810 4504 2866 4509
rect 3257 4532 3289 4539
rect 3257 4512 3263 4532
rect 3284 4512 3289 4532
rect 3749 4523 3783 4575
rect 4403 4565 4406 4592
rect 4435 4568 4480 4592
rect 4509 4568 4513 4595
rect 4435 4565 4513 4568
rect 4403 4551 4513 4565
rect 4699 4595 4741 4605
rect 4699 4576 4707 4595
rect 4732 4576 4741 4595
rect 5977 4578 6008 4624
rect 4699 4523 4741 4576
rect 5476 4553 5587 4575
rect 5476 4533 5484 4553
rect 5503 4533 5561 4553
rect 5580 4533 5587 4553
rect 5976 4561 6008 4578
rect 6277 4561 6314 4697
rect 6415 4664 6525 4678
rect 6415 4661 6493 4664
rect 6415 4634 6419 4661
rect 6448 4637 6493 4661
rect 6522 4637 6525 4664
rect 7145 4654 7179 4697
rect 6448 4634 6525 4637
rect 6415 4619 6525 4634
rect 7144 4649 7179 4654
rect 7144 4629 7151 4649
rect 7171 4629 7179 4649
rect 7144 4621 7179 4629
rect 5976 4548 6314 4561
rect 2810 4298 2844 4504
rect 3257 4484 3289 4512
rect 3747 4497 4743 4523
rect 5476 4516 5587 4533
rect 5977 4529 6314 4548
rect 6256 4528 6314 4529
rect 6700 4556 6732 4563
rect 6700 4536 6707 4556
rect 6728 4536 6732 4556
rect 2877 4476 3289 4484
rect 2877 4450 2883 4476
rect 2909 4450 3289 4476
rect 2877 4448 3289 4450
rect 2879 4447 2919 4448
rect 3039 4412 3078 4427
rect 3039 4371 3050 4412
rect 3071 4371 3078 4412
rect 2809 4290 2845 4298
rect 2809 4270 2818 4290
rect 2838 4270 2845 4290
rect 2809 4269 2845 4270
rect 2809 4258 2843 4269
rect 3039 4098 3078 4371
rect 3257 4383 3289 4448
rect 6700 4471 6732 4536
rect 7070 4471 7110 4472
rect 6700 4469 7112 4471
rect 6700 4443 7080 4469
rect 7106 4443 7112 4469
rect 6700 4435 7112 4443
rect 3257 4363 3261 4383
rect 3282 4363 3289 4383
rect 3257 4356 3289 4363
rect 3675 4390 3733 4391
rect 3675 4371 4012 4390
rect 4402 4386 4513 4403
rect 5246 4396 6242 4422
rect 6700 4407 6732 4435
rect 3675 4358 4013 4371
rect 3179 4294 3232 4297
rect 3179 4277 3191 4294
rect 3223 4277 3232 4294
rect 3179 4269 3232 4277
rect 3178 4222 3232 4269
rect 3464 4285 3574 4300
rect 3464 4282 3541 4285
rect 3464 4255 3467 4282
rect 3496 4258 3541 4282
rect 3570 4258 3574 4285
rect 3496 4255 3574 4258
rect 3464 4241 3574 4255
rect 3675 4222 3712 4358
rect 3981 4341 4013 4358
rect 4402 4366 4409 4386
rect 4428 4366 4486 4386
rect 4505 4366 4513 4386
rect 4402 4344 4513 4366
rect 5248 4343 5290 4396
rect 3981 4295 4012 4341
rect 5248 4324 5257 4343
rect 5282 4324 5290 4343
rect 5248 4314 5290 4324
rect 5476 4354 5586 4368
rect 5476 4351 5554 4354
rect 5476 4324 5480 4351
rect 5509 4327 5554 4351
rect 5583 4327 5586 4354
rect 6206 4344 6240 4396
rect 6700 4387 6705 4407
rect 6726 4387 6732 4407
rect 6700 4380 6732 4387
rect 6910 4408 6948 4418
rect 7145 4415 7179 4621
rect 6910 4391 6920 4408
rect 6940 4391 6948 4408
rect 6751 4348 6792 4349
rect 5509 4324 5586 4327
rect 5476 4309 5586 4324
rect 6205 4339 6240 4344
rect 6205 4319 6212 4339
rect 6232 4319 6240 4339
rect 6750 4338 6792 4348
rect 6205 4311 6240 4319
rect 3769 4292 3804 4293
rect 3748 4285 3804 4292
rect 3748 4265 3777 4285
rect 3797 4265 3804 4285
rect 3748 4260 3804 4265
rect 3981 4288 4020 4295
rect 3981 4268 3987 4288
rect 4012 4268 4020 4288
rect 3981 4262 4020 4268
rect 4195 4288 4227 4295
rect 4195 4268 4201 4288
rect 4222 4268 4227 4288
rect 3178 4187 3713 4222
rect 3178 4183 3231 4187
rect 3039 4071 3043 4098
rect 3074 4071 3078 4098
rect 3324 4119 3435 4136
rect 3324 4099 3331 4119
rect 3350 4099 3408 4119
rect 3427 4099 3435 4119
rect 3324 4077 3435 4099
rect 3039 4064 3078 4071
rect 3748 4054 3782 4260
rect 4195 4240 4227 4268
rect 3815 4232 4227 4240
rect 3815 4206 3821 4232
rect 3847 4206 4227 4232
rect 3815 4204 4227 4206
rect 3817 4203 3857 4204
rect 4195 4139 4227 4204
rect 5761 4246 5793 4253
rect 5761 4226 5768 4246
rect 5789 4226 5793 4246
rect 5761 4161 5793 4226
rect 6131 4161 6171 4162
rect 5761 4159 6173 4161
rect 4195 4119 4199 4139
rect 4220 4119 4227 4139
rect 4195 4112 4227 4119
rect 4698 4154 4746 4159
rect 4698 4125 4709 4154
rect 4738 4125 4746 4154
rect 3748 4053 3783 4054
rect 3746 4046 3783 4053
rect 2691 4025 2726 4026
rect 2668 4018 2726 4025
rect 2668 3998 2699 4018
rect 2719 3998 2726 4018
rect 2668 3993 2726 3998
rect 3117 4021 3149 4028
rect 3117 4001 3123 4021
rect 3144 4001 3149 4021
rect 2668 3845 2704 3993
rect 3117 3973 3149 4001
rect 2737 3965 3149 3973
rect 2737 3939 2743 3965
rect 2769 3939 3149 3965
rect 3746 4026 3756 4046
rect 3776 4026 3783 4046
rect 3746 4021 3783 4026
rect 4402 4041 4512 4056
rect 4402 4038 4479 4041
rect 3746 3970 3781 4021
rect 4402 4011 4405 4038
rect 4434 4014 4479 4038
rect 4508 4014 4512 4041
rect 4434 4011 4512 4014
rect 4402 3997 4512 4011
rect 4698 3970 4746 4125
rect 5761 4133 6141 4159
rect 6167 4133 6173 4159
rect 5761 4125 6173 4133
rect 5761 4097 5793 4125
rect 6206 4105 6240 4311
rect 6414 4309 6525 4331
rect 6414 4289 6422 4309
rect 6441 4289 6499 4309
rect 6518 4289 6525 4309
rect 6414 4272 6525 4289
rect 6750 4316 6757 4338
rect 6783 4316 6792 4338
rect 6750 4307 6792 4316
rect 5967 4102 6010 4104
rect 5761 4077 5766 4097
rect 5787 4077 5793 4097
rect 5761 4070 5793 4077
rect 5966 4095 6010 4102
rect 5966 4075 5976 4095
rect 5999 4075 6010 4095
rect 5966 4071 6010 4075
rect 6184 4100 6240 4105
rect 6184 4080 6191 4100
rect 6211 4080 6240 4100
rect 6184 4073 6240 4080
rect 6296 4241 6329 4242
rect 6750 4241 6787 4307
rect 6296 4212 6787 4241
rect 6184 4072 6219 4073
rect 3746 3946 4746 3970
rect 5475 3999 5586 4021
rect 5475 3979 5483 3999
rect 5502 3979 5560 3999
rect 5579 3979 5586 3999
rect 5475 3962 5586 3979
rect 5966 3990 6008 4071
rect 6296 3992 6329 4212
rect 6750 4210 6787 4212
rect 6556 4072 6666 4086
rect 6556 4069 6634 4072
rect 6556 4042 6560 4069
rect 6589 4045 6634 4069
rect 6663 4045 6666 4072
rect 6589 4042 6666 4045
rect 6556 4027 6666 4042
rect 6910 4053 6948 4391
rect 7123 4410 7179 4415
rect 7123 4390 7130 4410
rect 7150 4390 7179 4410
rect 7123 4383 7179 4390
rect 7388 4682 7395 4722
rect 7422 4682 7435 4722
rect 7618 4700 7665 4878
rect 8411 4869 8414 4896
rect 8443 4872 8488 4896
rect 8517 4872 8521 4899
rect 8443 4869 8521 4872
rect 8411 4855 8521 4869
rect 7123 4382 7158 4383
rect 7288 4062 7320 4063
rect 6910 4036 6918 4053
rect 6938 4036 6948 4053
rect 6910 4030 6948 4036
rect 7285 4057 7320 4062
rect 7285 4037 7292 4057
rect 7312 4037 7320 4057
rect 7285 4029 7320 4037
rect 6268 3990 6329 3992
rect 5966 3961 6329 3990
rect 6841 3964 6873 3971
rect 5966 3959 6268 3961
rect 3746 3943 4745 3946
rect 6841 3944 6848 3964
rect 6869 3944 6873 3964
rect 3746 3941 3781 3943
rect 2737 3937 3149 3939
rect 2739 3936 2779 3937
rect 2671 3787 2704 3845
rect 2901 3897 2939 3907
rect 2901 3859 2910 3897
rect 2933 3859 2939 3897
rect 2671 3779 2705 3787
rect 2671 3759 2678 3779
rect 2698 3759 2705 3779
rect 2671 3754 2705 3759
rect 2671 3753 2702 3754
rect 2901 3723 2939 3859
rect 3117 3872 3149 3937
rect 6841 3879 6873 3944
rect 7211 3879 7251 3880
rect 6841 3877 7253 3879
rect 6209 3873 6244 3875
rect 3117 3852 3121 3872
rect 3142 3852 3149 3872
rect 5245 3870 6244 3873
rect 3722 3855 4024 3857
rect 3117 3845 3149 3852
rect 3661 3826 4024 3855
rect 3661 3824 3722 3826
rect 3042 3780 3080 3786
rect 3042 3763 3052 3780
rect 3072 3763 3080 3780
rect 2901 3569 2945 3723
rect 2738 3567 2945 3569
rect 2714 3534 2945 3567
rect 1811 2908 1815 2928
rect 1836 2908 1845 2928
rect 1811 2902 1845 2908
rect 1964 3039 2293 3042
rect 2332 3039 2376 3064
rect 1964 3009 2376 3039
rect 1213 2846 1274 2848
rect 911 2817 1274 2846
rect 1755 2833 1787 2840
rect 911 2815 1213 2817
rect 1755 2813 1762 2833
rect 1783 2813 1787 2833
rect 1755 2748 1787 2813
rect 1964 2821 1999 3009
rect 2266 3007 2376 3009
rect 2559 3022 2609 3150
rect 2714 3133 2764 3534
rect 2901 3530 2945 3534
rect 2832 3433 2867 3434
rect 2694 3124 2764 3133
rect 2694 3095 2709 3124
rect 2757 3116 2764 3124
rect 2811 3426 2867 3433
rect 2811 3406 2840 3426
rect 2860 3406 2867 3426
rect 2811 3401 2867 3406
rect 3042 3425 3080 3763
rect 3324 3774 3434 3789
rect 3324 3771 3401 3774
rect 3324 3744 3327 3771
rect 3356 3747 3401 3771
rect 3430 3747 3434 3774
rect 3356 3744 3434 3747
rect 3324 3730 3434 3744
rect 3203 3604 3240 3606
rect 3661 3604 3694 3824
rect 3982 3745 4024 3826
rect 4404 3837 4515 3854
rect 4404 3817 4411 3837
rect 4430 3817 4488 3837
rect 4507 3817 4515 3837
rect 4404 3795 4515 3817
rect 5244 3846 6244 3870
rect 3771 3743 3806 3744
rect 3203 3575 3694 3604
rect 3203 3509 3240 3575
rect 3661 3574 3694 3575
rect 3750 3736 3806 3743
rect 3750 3716 3779 3736
rect 3799 3716 3806 3736
rect 3750 3711 3806 3716
rect 3980 3741 4024 3745
rect 3980 3721 3991 3741
rect 4014 3721 4024 3741
rect 3980 3714 4024 3721
rect 4197 3739 4229 3746
rect 4197 3719 4203 3739
rect 4224 3719 4229 3739
rect 3980 3712 4023 3714
rect 3198 3500 3240 3509
rect 3198 3478 3207 3500
rect 3233 3478 3240 3500
rect 3465 3527 3576 3544
rect 3465 3507 3472 3527
rect 3491 3507 3549 3527
rect 3568 3507 3576 3527
rect 3465 3485 3576 3507
rect 3750 3505 3784 3711
rect 4197 3691 4229 3719
rect 3817 3683 4229 3691
rect 3817 3657 3823 3683
rect 3849 3657 4229 3683
rect 5244 3691 5292 3846
rect 5478 3805 5588 3819
rect 5478 3802 5556 3805
rect 5478 3775 5482 3802
rect 5511 3778 5556 3802
rect 5585 3778 5588 3805
rect 6209 3795 6244 3846
rect 5511 3775 5588 3778
rect 5478 3760 5588 3775
rect 6207 3790 6244 3795
rect 6207 3770 6214 3790
rect 6234 3770 6244 3790
rect 6841 3851 7221 3877
rect 7247 3851 7253 3877
rect 6841 3843 7253 3851
rect 6841 3815 6873 3843
rect 6841 3795 6846 3815
rect 6867 3795 6873 3815
rect 6841 3788 6873 3795
rect 7047 3814 7089 3825
rect 7286 3823 7320 4029
rect 7047 3793 7054 3814
rect 7081 3793 7089 3814
rect 6207 3763 6244 3770
rect 6207 3762 6242 3763
rect 5244 3662 5252 3691
rect 5281 3662 5292 3691
rect 5244 3657 5292 3662
rect 5763 3697 5795 3704
rect 5763 3677 5770 3697
rect 5791 3677 5795 3697
rect 3817 3655 4229 3657
rect 3819 3654 3859 3655
rect 4197 3590 4229 3655
rect 4197 3570 4201 3590
rect 4222 3570 4229 3590
rect 4197 3563 4229 3570
rect 5763 3612 5795 3677
rect 6133 3612 6173 3613
rect 5763 3610 6175 3612
rect 5763 3584 6143 3610
rect 6169 3584 6175 3610
rect 5763 3576 6175 3584
rect 5763 3548 5795 3576
rect 6208 3556 6242 3762
rect 6912 3745 6951 3752
rect 6555 3717 6666 3739
rect 6555 3697 6563 3717
rect 6582 3697 6640 3717
rect 6659 3697 6666 3717
rect 6555 3680 6666 3697
rect 6912 3718 6916 3745
rect 6947 3718 6951 3745
rect 6759 3629 6812 3633
rect 6277 3594 6812 3629
rect 5763 3528 5768 3548
rect 5789 3528 5795 3548
rect 5763 3521 5795 3528
rect 5970 3548 6009 3554
rect 5970 3528 5978 3548
rect 6003 3528 6009 3548
rect 5970 3521 6009 3528
rect 6186 3551 6242 3556
rect 6186 3531 6193 3551
rect 6213 3531 6242 3551
rect 6186 3524 6242 3531
rect 6186 3523 6221 3524
rect 3750 3497 3785 3505
rect 3198 3468 3240 3478
rect 3750 3477 3758 3497
rect 3778 3477 3785 3497
rect 3750 3472 3785 3477
rect 4404 3492 4514 3507
rect 4404 3489 4481 3492
rect 3198 3467 3239 3468
rect 3042 3408 3050 3425
rect 3070 3408 3080 3425
rect 2811 3195 2845 3401
rect 3042 3398 3080 3408
rect 3258 3429 3290 3436
rect 3258 3409 3264 3429
rect 3285 3409 3290 3429
rect 3750 3420 3784 3472
rect 4404 3462 4407 3489
rect 4436 3465 4481 3489
rect 4510 3465 4514 3492
rect 4436 3462 4514 3465
rect 4404 3448 4514 3462
rect 4700 3492 4742 3502
rect 4700 3473 4708 3492
rect 4733 3473 4742 3492
rect 5978 3475 6009 3521
rect 4700 3420 4742 3473
rect 5477 3450 5588 3472
rect 5477 3430 5485 3450
rect 5504 3430 5562 3450
rect 5581 3430 5588 3450
rect 5977 3458 6009 3475
rect 6278 3458 6315 3594
rect 6416 3561 6526 3575
rect 6416 3558 6494 3561
rect 6416 3531 6420 3558
rect 6449 3534 6494 3558
rect 6523 3534 6526 3561
rect 6449 3531 6526 3534
rect 6416 3516 6526 3531
rect 6758 3547 6812 3594
rect 6758 3539 6811 3547
rect 6758 3522 6767 3539
rect 6799 3522 6811 3539
rect 6758 3519 6811 3522
rect 5977 3445 6315 3458
rect 3258 3381 3290 3409
rect 3748 3394 4744 3420
rect 5477 3413 5588 3430
rect 5978 3426 6315 3445
rect 6257 3425 6315 3426
rect 6701 3453 6733 3460
rect 6701 3433 6708 3453
rect 6729 3433 6733 3453
rect 2878 3373 3290 3381
rect 2878 3347 2884 3373
rect 2910 3347 3290 3373
rect 2878 3345 3290 3347
rect 2880 3344 2920 3345
rect 3258 3280 3290 3345
rect 6701 3368 6733 3433
rect 6912 3445 6951 3718
rect 7047 3622 7089 3793
rect 7264 3818 7320 3823
rect 7264 3798 7271 3818
rect 7291 3798 7320 3818
rect 7264 3791 7320 3798
rect 7264 3790 7299 3791
rect 7047 3588 7291 3622
rect 7254 3580 7291 3588
rect 7147 3547 7181 3558
rect 7145 3546 7181 3547
rect 7145 3526 7152 3546
rect 7172 3526 7181 3546
rect 7145 3518 7181 3526
rect 6912 3404 6919 3445
rect 6940 3404 6951 3445
rect 6912 3389 6951 3404
rect 7071 3368 7111 3369
rect 6701 3366 7113 3368
rect 6701 3340 7081 3366
rect 7107 3340 7113 3366
rect 6701 3332 7113 3340
rect 3258 3260 3262 3280
rect 3283 3260 3290 3280
rect 3258 3253 3290 3260
rect 3676 3287 3734 3288
rect 3676 3268 4013 3287
rect 4403 3283 4514 3300
rect 5247 3293 6243 3319
rect 6701 3304 6733 3332
rect 7146 3312 7180 3518
rect 3676 3255 4014 3268
rect 2811 3187 2846 3195
rect 2811 3167 2819 3187
rect 2839 3167 2846 3187
rect 2811 3162 2846 3167
rect 3465 3182 3575 3197
rect 3465 3179 3542 3182
rect 2811 3119 2845 3162
rect 3465 3152 3468 3179
rect 3497 3155 3542 3179
rect 3571 3155 3575 3182
rect 3497 3152 3575 3155
rect 3465 3138 3575 3152
rect 3676 3119 3713 3255
rect 3982 3238 4014 3255
rect 4403 3263 4410 3283
rect 4429 3263 4487 3283
rect 4506 3263 4514 3283
rect 4403 3241 4514 3263
rect 5249 3240 5291 3293
rect 3982 3192 4013 3238
rect 5249 3221 5258 3240
rect 5283 3221 5291 3240
rect 5249 3211 5291 3221
rect 5477 3251 5587 3265
rect 5477 3248 5555 3251
rect 5477 3221 5481 3248
rect 5510 3224 5555 3248
rect 5584 3224 5587 3251
rect 6207 3241 6241 3293
rect 6701 3284 6706 3304
rect 6727 3284 6733 3304
rect 6701 3277 6733 3284
rect 7124 3307 7180 3312
rect 7124 3287 7131 3307
rect 7151 3287 7180 3307
rect 7124 3280 7180 3287
rect 7124 3279 7159 3280
rect 6752 3245 6793 3246
rect 5510 3221 5587 3224
rect 5477 3206 5587 3221
rect 6206 3236 6241 3241
rect 6206 3216 6213 3236
rect 6233 3216 6241 3236
rect 6751 3235 6793 3245
rect 6206 3208 6241 3216
rect 3770 3189 3805 3190
rect 3749 3182 3805 3189
rect 3749 3162 3778 3182
rect 3798 3162 3805 3182
rect 3749 3157 3805 3162
rect 3982 3185 4021 3192
rect 3982 3165 3988 3185
rect 4013 3165 4021 3185
rect 3982 3159 4021 3165
rect 4196 3185 4228 3192
rect 4196 3165 4202 3185
rect 4223 3165 4228 3185
rect 2757 3095 2762 3116
rect 2694 3084 2762 3095
rect 2810 3084 3714 3119
rect 2811 3083 2845 3084
rect 2559 2988 2974 3022
rect 2559 2986 2609 2988
rect 2192 2924 2242 2931
rect 2192 2910 2206 2924
rect 2198 2906 2206 2910
rect 2226 2910 2242 2924
rect 2226 2906 2236 2910
rect 2722 2909 2757 2910
rect 2198 2899 2236 2906
rect 2701 2902 2757 2909
rect 2199 2898 2234 2899
rect 1964 2789 1969 2821
rect 1996 2789 1999 2821
rect 1964 2771 1999 2789
rect 2125 2748 2165 2749
rect 1755 2746 2167 2748
rect 1153 2729 1188 2731
rect 189 2726 1188 2729
rect 188 2702 1188 2726
rect 188 2547 236 2702
rect 422 2661 532 2675
rect 422 2658 500 2661
rect 422 2631 426 2658
rect 455 2634 500 2658
rect 529 2634 532 2661
rect 1153 2651 1188 2702
rect 1755 2720 2135 2746
rect 2161 2720 2167 2746
rect 1755 2712 2167 2720
rect 1755 2684 1787 2712
rect 2200 2692 2234 2898
rect 1755 2664 1760 2684
rect 1781 2664 1787 2684
rect 1755 2657 1787 2664
rect 2178 2687 2234 2692
rect 2178 2667 2185 2687
rect 2205 2667 2234 2687
rect 2701 2882 2730 2902
rect 2750 2882 2757 2902
rect 2701 2877 2757 2882
rect 2929 2905 2974 2988
rect 3355 3003 3466 3020
rect 3355 2983 3362 3003
rect 3381 2983 3439 3003
rect 3458 2983 3466 3003
rect 3355 2961 3466 2983
rect 3749 2951 3783 3157
rect 4196 3137 4228 3165
rect 3816 3129 4228 3137
rect 3816 3103 3822 3129
rect 3848 3103 4228 3129
rect 3816 3101 4228 3103
rect 3818 3100 3858 3101
rect 4196 3036 4228 3101
rect 5762 3143 5794 3150
rect 5762 3123 5769 3143
rect 5790 3123 5794 3143
rect 5762 3058 5794 3123
rect 6132 3058 6172 3059
rect 5762 3056 6174 3058
rect 4196 3016 4200 3036
rect 4221 3016 4228 3036
rect 4196 3009 4228 3016
rect 4699 3051 4747 3056
rect 4699 3022 4710 3051
rect 4739 3022 4747 3051
rect 3749 2950 3784 2951
rect 3747 2943 3784 2950
rect 3747 2923 3757 2943
rect 3777 2923 3784 2943
rect 3747 2918 3784 2923
rect 4403 2938 4513 2953
rect 4403 2935 4480 2938
rect 2929 2886 2938 2905
rect 2967 2886 2974 2905
rect 2701 2671 2735 2877
rect 2929 2874 2974 2886
rect 3148 2905 3180 2912
rect 3148 2885 3154 2905
rect 3175 2885 3180 2905
rect 3148 2857 3180 2885
rect 2768 2849 3180 2857
rect 2768 2823 2774 2849
rect 2800 2823 3180 2849
rect 3747 2867 3782 2918
rect 4403 2908 4406 2935
rect 4435 2911 4480 2935
rect 4509 2911 4513 2938
rect 4435 2908 4513 2911
rect 4403 2894 4513 2908
rect 4699 2867 4747 3022
rect 5762 3030 6142 3056
rect 6168 3030 6174 3056
rect 5762 3022 6174 3030
rect 5762 2994 5794 3022
rect 6207 3002 6241 3208
rect 6415 3206 6526 3228
rect 6415 3186 6423 3206
rect 6442 3186 6500 3206
rect 6519 3186 6526 3206
rect 6415 3169 6526 3186
rect 6751 3213 6758 3235
rect 6784 3213 6793 3235
rect 6751 3204 6793 3213
rect 5968 2999 6011 3001
rect 5762 2974 5767 2994
rect 5788 2974 5794 2994
rect 5762 2967 5794 2974
rect 5967 2992 6011 2999
rect 5967 2972 5977 2992
rect 6000 2972 6011 2992
rect 5967 2968 6011 2972
rect 6185 2997 6241 3002
rect 6185 2977 6192 2997
rect 6212 2977 6241 2997
rect 6185 2970 6241 2977
rect 6297 3138 6330 3139
rect 6751 3138 6788 3204
rect 7254 3189 7292 3580
rect 6868 3173 7292 3189
rect 6297 3109 6788 3138
rect 6185 2969 6220 2970
rect 3747 2843 4747 2867
rect 5476 2896 5587 2918
rect 5476 2876 5484 2896
rect 5503 2876 5561 2896
rect 5580 2876 5587 2896
rect 5476 2860 5587 2876
rect 5967 2887 6009 2968
rect 6297 2889 6330 3109
rect 6751 3107 6788 3109
rect 6867 3148 7292 3173
rect 6526 2982 6636 2996
rect 6526 2979 6604 2982
rect 6526 2952 6530 2979
rect 6559 2955 6604 2979
rect 6633 2955 6636 2982
rect 6559 2952 6636 2955
rect 6526 2937 6636 2952
rect 6867 2969 6901 3148
rect 7388 3105 7435 4682
rect 7617 4676 7665 4700
rect 8258 4748 8295 4750
rect 8716 4748 8749 4968
rect 9037 4889 9079 4970
rect 9459 4981 9570 4998
rect 9459 4961 9466 4981
rect 9485 4961 9543 4981
rect 9562 4961 9570 4981
rect 9459 4939 9570 4961
rect 11784 4965 11816 5030
rect 12154 4965 12194 4966
rect 11784 4963 12196 4965
rect 11183 4940 11218 4942
rect 10219 4937 11218 4940
rect 10218 4913 11218 4937
rect 8826 4887 8861 4888
rect 8258 4719 8749 4748
rect 7617 3191 7663 4676
rect 8258 4653 8295 4719
rect 8716 4718 8749 4719
rect 8805 4880 8861 4887
rect 8805 4860 8834 4880
rect 8854 4860 8861 4880
rect 8805 4855 8861 4860
rect 9035 4885 9079 4889
rect 9035 4865 9046 4885
rect 9069 4865 9079 4885
rect 9035 4858 9079 4865
rect 9252 4883 9284 4890
rect 9252 4863 9258 4883
rect 9279 4863 9284 4883
rect 9035 4856 9078 4858
rect 8253 4644 8295 4653
rect 8253 4622 8262 4644
rect 8288 4622 8295 4644
rect 8520 4671 8631 4688
rect 8520 4651 8527 4671
rect 8546 4651 8604 4671
rect 8623 4651 8631 4671
rect 8520 4629 8631 4651
rect 8805 4649 8839 4855
rect 9252 4835 9284 4863
rect 8872 4827 9284 4835
rect 8872 4801 8878 4827
rect 8904 4801 9284 4827
rect 8872 4799 9284 4801
rect 8874 4798 8914 4799
rect 9252 4734 9284 4799
rect 9252 4714 9256 4734
rect 9277 4714 9284 4734
rect 10218 4758 10266 4913
rect 10452 4872 10562 4886
rect 10452 4869 10530 4872
rect 10452 4842 10456 4869
rect 10485 4845 10530 4869
rect 10559 4845 10562 4872
rect 11183 4862 11218 4913
rect 11784 4937 12164 4963
rect 12190 4937 12196 4963
rect 11784 4929 12196 4937
rect 11784 4901 11816 4929
rect 12229 4909 12263 5115
rect 12753 5114 12788 5115
rect 11784 4881 11789 4901
rect 11810 4881 11816 4901
rect 11784 4874 11816 4881
rect 11986 4904 12031 4909
rect 11986 4880 11997 4904
rect 12023 4880 12031 4904
rect 11986 4869 12031 4880
rect 12207 4904 12263 4909
rect 12207 4884 12214 4904
rect 12234 4884 12263 4904
rect 12207 4877 12263 4884
rect 12732 5107 12788 5114
rect 12732 5087 12761 5107
rect 12781 5087 12788 5107
rect 12732 5082 12788 5087
rect 12957 5110 13002 5189
rect 13386 5208 13497 5225
rect 13386 5188 13393 5208
rect 13412 5188 13470 5208
rect 13489 5188 13497 5208
rect 13386 5166 13497 5188
rect 13779 5162 13813 5368
rect 14226 5348 14258 5376
rect 13846 5340 14258 5348
rect 13846 5314 13852 5340
rect 13878 5314 14258 5340
rect 13846 5312 14258 5314
rect 13848 5311 13888 5312
rect 14226 5247 14258 5312
rect 15792 5354 15824 5361
rect 15792 5334 15799 5354
rect 15820 5334 15824 5354
rect 15792 5269 15824 5334
rect 16162 5269 16202 5270
rect 15792 5267 16204 5269
rect 14226 5227 14230 5247
rect 14251 5227 14258 5247
rect 14226 5220 14258 5227
rect 14729 5262 14777 5267
rect 14729 5233 14740 5262
rect 14769 5233 14777 5262
rect 13779 5161 13814 5162
rect 13777 5154 13814 5161
rect 13777 5134 13787 5154
rect 13807 5134 13814 5154
rect 13777 5129 13814 5134
rect 14433 5149 14543 5164
rect 14433 5146 14510 5149
rect 12957 5090 12968 5110
rect 12993 5090 13002 5110
rect 12957 5086 13002 5090
rect 13179 5110 13211 5117
rect 13179 5090 13185 5110
rect 13206 5090 13211 5110
rect 12207 4876 12242 4877
rect 12732 4876 12766 5082
rect 13179 5062 13211 5090
rect 12799 5054 13211 5062
rect 12799 5028 12805 5054
rect 12831 5028 13211 5054
rect 13777 5078 13812 5129
rect 14433 5119 14436 5146
rect 14465 5122 14510 5146
rect 14539 5122 14543 5149
rect 14465 5119 14543 5122
rect 14433 5105 14543 5119
rect 14729 5078 14777 5233
rect 15792 5241 16172 5267
rect 16198 5241 16204 5267
rect 15792 5233 16204 5241
rect 15792 5205 15824 5233
rect 16237 5213 16271 5419
rect 16445 5417 16556 5439
rect 16445 5397 16453 5417
rect 16472 5397 16530 5417
rect 16549 5397 16556 5417
rect 16445 5380 16556 5397
rect 16781 5424 16788 5446
rect 16814 5424 16823 5446
rect 16781 5415 16823 5424
rect 15998 5210 16041 5212
rect 15792 5185 15797 5205
rect 15818 5185 15824 5205
rect 15792 5178 15824 5185
rect 15997 5203 16041 5210
rect 15997 5183 16007 5203
rect 16030 5183 16041 5203
rect 15997 5179 16041 5183
rect 16215 5208 16271 5213
rect 16215 5188 16222 5208
rect 16242 5188 16271 5208
rect 16215 5181 16271 5188
rect 16327 5349 16360 5350
rect 16781 5349 16818 5415
rect 17413 5392 17459 6877
rect 16327 5320 16818 5349
rect 16215 5180 16250 5181
rect 13777 5054 14777 5078
rect 15506 5107 15617 5129
rect 15506 5087 15514 5107
rect 15533 5087 15591 5107
rect 15610 5087 15617 5107
rect 15506 5070 15617 5087
rect 15997 5098 16039 5179
rect 16327 5100 16360 5320
rect 16781 5318 16818 5320
rect 17411 5368 17459 5392
rect 17641 5386 17688 6963
rect 18175 6920 18209 7099
rect 18440 7116 18550 7131
rect 18440 7113 18517 7116
rect 18440 7086 18443 7113
rect 18472 7089 18517 7113
rect 18546 7089 18550 7116
rect 18472 7086 18550 7089
rect 18440 7072 18550 7086
rect 17784 6895 18209 6920
rect 18288 6959 18325 6961
rect 18746 6959 18779 7179
rect 19067 7100 19109 7181
rect 19489 7192 19600 7208
rect 19489 7172 19496 7192
rect 19515 7172 19573 7192
rect 19592 7172 19600 7192
rect 19489 7150 19600 7172
rect 18856 7098 18891 7099
rect 18288 6930 18779 6959
rect 17784 6879 18208 6895
rect 17784 6488 17822 6879
rect 18288 6864 18325 6930
rect 18746 6929 18779 6930
rect 18835 7091 18891 7098
rect 18835 7071 18864 7091
rect 18884 7071 18891 7091
rect 18835 7066 18891 7071
rect 19065 7096 19109 7100
rect 19065 7076 19076 7096
rect 19099 7076 19109 7096
rect 19065 7069 19109 7076
rect 19282 7094 19314 7101
rect 19282 7074 19288 7094
rect 19309 7074 19314 7094
rect 19065 7067 19108 7069
rect 18283 6855 18325 6864
rect 18283 6833 18292 6855
rect 18318 6833 18325 6855
rect 18550 6882 18661 6899
rect 18550 6862 18557 6882
rect 18576 6862 18634 6882
rect 18653 6862 18661 6882
rect 18550 6840 18661 6862
rect 18835 6860 18869 7066
rect 19282 7046 19314 7074
rect 18902 7038 19314 7046
rect 18902 7012 18908 7038
rect 18934 7012 19314 7038
rect 18902 7010 19314 7012
rect 18904 7009 18944 7010
rect 19282 6945 19314 7010
rect 19282 6925 19286 6945
rect 19307 6925 19314 6945
rect 19282 6918 19314 6925
rect 18835 6852 18870 6860
rect 18283 6823 18325 6833
rect 18835 6832 18843 6852
rect 18863 6832 18870 6852
rect 18835 6827 18870 6832
rect 19489 6847 19599 6862
rect 19489 6844 19566 6847
rect 18283 6822 18324 6823
rect 17917 6788 17952 6789
rect 17896 6781 17952 6788
rect 17896 6761 17925 6781
rect 17945 6761 17952 6781
rect 17896 6756 17952 6761
rect 18343 6784 18375 6791
rect 18343 6764 18349 6784
rect 18370 6764 18375 6784
rect 18835 6775 18869 6827
rect 19489 6817 19492 6844
rect 19521 6820 19566 6844
rect 19595 6820 19599 6847
rect 19521 6817 19599 6820
rect 19489 6803 19599 6817
rect 19785 6847 19827 6857
rect 19785 6828 19793 6847
rect 19818 6828 19827 6847
rect 19785 6775 19827 6828
rect 17896 6550 17930 6756
rect 18343 6736 18375 6764
rect 18833 6749 19829 6775
rect 17963 6728 18375 6736
rect 17963 6702 17969 6728
rect 17995 6702 18375 6728
rect 17963 6700 18375 6702
rect 17965 6699 18005 6700
rect 18125 6664 18164 6679
rect 18125 6623 18136 6664
rect 18157 6623 18164 6664
rect 17895 6542 17931 6550
rect 17895 6522 17904 6542
rect 17924 6522 17931 6542
rect 17895 6521 17931 6522
rect 17895 6510 17929 6521
rect 17785 6480 17822 6488
rect 17785 6446 18029 6480
rect 17777 6277 17812 6278
rect 17756 6270 17812 6277
rect 17756 6250 17785 6270
rect 17805 6250 17812 6270
rect 17756 6245 17812 6250
rect 17987 6275 18029 6446
rect 18125 6350 18164 6623
rect 18343 6635 18375 6700
rect 18343 6615 18347 6635
rect 18368 6615 18375 6635
rect 18343 6608 18375 6615
rect 18761 6642 18819 6643
rect 18761 6623 19098 6642
rect 19488 6638 19599 6655
rect 18761 6610 19099 6623
rect 18265 6546 18318 6549
rect 18265 6529 18277 6546
rect 18309 6529 18318 6546
rect 18265 6521 18318 6529
rect 18264 6474 18318 6521
rect 18550 6537 18660 6552
rect 18550 6534 18627 6537
rect 18550 6507 18553 6534
rect 18582 6510 18627 6534
rect 18656 6510 18660 6537
rect 18582 6507 18660 6510
rect 18550 6493 18660 6507
rect 18761 6474 18798 6610
rect 19067 6593 19099 6610
rect 19488 6618 19495 6638
rect 19514 6618 19572 6638
rect 19591 6618 19599 6638
rect 19488 6596 19599 6618
rect 19067 6547 19098 6593
rect 18855 6544 18890 6545
rect 18834 6537 18890 6544
rect 18834 6517 18863 6537
rect 18883 6517 18890 6537
rect 18834 6512 18890 6517
rect 19067 6540 19106 6547
rect 19067 6520 19073 6540
rect 19098 6520 19106 6540
rect 19067 6514 19106 6520
rect 19281 6540 19313 6547
rect 19281 6520 19287 6540
rect 19308 6520 19313 6540
rect 18264 6439 18799 6474
rect 18264 6435 18317 6439
rect 18125 6323 18129 6350
rect 18160 6323 18164 6350
rect 18410 6371 18521 6388
rect 18410 6351 18417 6371
rect 18436 6351 18494 6371
rect 18513 6351 18521 6371
rect 18410 6329 18521 6351
rect 18125 6316 18164 6323
rect 18834 6306 18868 6512
rect 19281 6492 19313 6520
rect 18901 6484 19313 6492
rect 18901 6458 18907 6484
rect 18933 6458 19313 6484
rect 18901 6456 19313 6458
rect 18903 6455 18943 6456
rect 19281 6391 19313 6456
rect 19281 6371 19285 6391
rect 19306 6371 19313 6391
rect 19281 6364 19313 6371
rect 19784 6406 19832 6411
rect 19784 6377 19795 6406
rect 19824 6377 19832 6406
rect 18834 6305 18869 6306
rect 18832 6298 18869 6305
rect 17987 6254 17995 6275
rect 18022 6254 18029 6275
rect 17756 6039 17790 6245
rect 17987 6243 18029 6254
rect 18203 6273 18235 6280
rect 18203 6253 18209 6273
rect 18230 6253 18235 6273
rect 18203 6225 18235 6253
rect 17823 6217 18235 6225
rect 17823 6191 17829 6217
rect 17855 6191 18235 6217
rect 18832 6278 18842 6298
rect 18862 6278 18869 6298
rect 18832 6273 18869 6278
rect 19488 6293 19598 6308
rect 19488 6290 19565 6293
rect 18832 6222 18867 6273
rect 19488 6263 19491 6290
rect 19520 6266 19565 6290
rect 19594 6266 19598 6293
rect 19520 6263 19598 6266
rect 19488 6249 19598 6263
rect 19784 6222 19832 6377
rect 18832 6198 19832 6222
rect 18832 6195 19831 6198
rect 18832 6193 18867 6195
rect 17823 6189 18235 6191
rect 17825 6188 17865 6189
rect 18203 6124 18235 6189
rect 18203 6104 18207 6124
rect 18228 6104 18235 6124
rect 18808 6107 19110 6109
rect 18203 6097 18235 6104
rect 18747 6078 19110 6107
rect 18747 6076 18808 6078
rect 17756 6031 17791 6039
rect 17756 6011 17764 6031
rect 17784 6011 17791 6031
rect 17756 6006 17791 6011
rect 18128 6032 18166 6038
rect 18128 6015 18138 6032
rect 18158 6015 18166 6032
rect 17756 6005 17788 6006
rect 17918 5685 17953 5686
rect 16555 5199 16665 5213
rect 16555 5196 16633 5199
rect 16555 5169 16559 5196
rect 16588 5172 16633 5196
rect 16662 5172 16665 5199
rect 17411 5190 17458 5368
rect 17641 5346 17654 5386
rect 17681 5346 17688 5386
rect 17897 5678 17953 5685
rect 17897 5658 17926 5678
rect 17946 5658 17953 5678
rect 17897 5653 17953 5658
rect 18128 5677 18166 6015
rect 18410 6026 18520 6041
rect 18410 6023 18487 6026
rect 18410 5996 18413 6023
rect 18442 5999 18487 6023
rect 18516 5999 18520 6026
rect 18442 5996 18520 5999
rect 18410 5982 18520 5996
rect 18289 5856 18326 5858
rect 18747 5856 18780 6076
rect 19068 5997 19110 6078
rect 19490 6089 19601 6106
rect 19490 6069 19497 6089
rect 19516 6069 19574 6089
rect 19593 6069 19601 6089
rect 19490 6047 19601 6069
rect 18857 5995 18892 5996
rect 18289 5827 18780 5856
rect 18289 5761 18326 5827
rect 18747 5826 18780 5827
rect 18836 5988 18892 5995
rect 18836 5968 18865 5988
rect 18885 5968 18892 5988
rect 18836 5963 18892 5968
rect 19066 5993 19110 5997
rect 19066 5973 19077 5993
rect 19100 5973 19110 5993
rect 19066 5966 19110 5973
rect 19283 5991 19315 5998
rect 19283 5971 19289 5991
rect 19310 5971 19315 5991
rect 19066 5964 19109 5966
rect 18284 5752 18326 5761
rect 18284 5730 18293 5752
rect 18319 5730 18326 5752
rect 18551 5779 18662 5796
rect 18551 5759 18558 5779
rect 18577 5759 18635 5779
rect 18654 5759 18662 5779
rect 18551 5737 18662 5759
rect 18836 5757 18870 5963
rect 19283 5943 19315 5971
rect 18903 5935 19315 5943
rect 18903 5909 18909 5935
rect 18935 5909 19315 5935
rect 18903 5907 19315 5909
rect 18905 5906 18945 5907
rect 19283 5842 19315 5907
rect 19283 5822 19287 5842
rect 19308 5822 19315 5842
rect 19283 5815 19315 5822
rect 18836 5749 18871 5757
rect 18284 5720 18326 5730
rect 18836 5729 18844 5749
rect 18864 5729 18871 5749
rect 18836 5724 18871 5729
rect 19490 5744 19600 5759
rect 19490 5741 19567 5744
rect 18284 5719 18325 5720
rect 18128 5660 18136 5677
rect 18156 5660 18166 5677
rect 17897 5447 17931 5653
rect 18128 5650 18166 5660
rect 18344 5681 18376 5688
rect 18344 5661 18350 5681
rect 18371 5661 18376 5681
rect 18836 5672 18870 5724
rect 19490 5714 19493 5741
rect 19522 5717 19567 5741
rect 19596 5717 19600 5744
rect 19522 5714 19600 5717
rect 19490 5700 19600 5714
rect 19786 5744 19828 5754
rect 19786 5725 19794 5744
rect 19819 5725 19828 5744
rect 19786 5672 19828 5725
rect 18344 5633 18376 5661
rect 18834 5646 19830 5672
rect 17964 5625 18376 5633
rect 17964 5599 17970 5625
rect 17996 5599 18376 5625
rect 17964 5597 18376 5599
rect 17966 5596 18006 5597
rect 18344 5532 18376 5597
rect 18344 5512 18348 5532
rect 18369 5512 18376 5532
rect 18344 5505 18376 5512
rect 18762 5539 18820 5540
rect 18762 5520 19099 5539
rect 19489 5535 19600 5552
rect 18762 5507 19100 5520
rect 17897 5439 17932 5447
rect 17897 5419 17905 5439
rect 17925 5419 17932 5439
rect 17897 5414 17932 5419
rect 18551 5434 18661 5449
rect 18551 5431 18628 5434
rect 17897 5371 17931 5414
rect 18551 5404 18554 5431
rect 18583 5407 18628 5431
rect 18657 5407 18661 5434
rect 18583 5404 18661 5407
rect 18551 5390 18661 5404
rect 18762 5371 18799 5507
rect 19068 5490 19100 5507
rect 19489 5515 19496 5535
rect 19515 5515 19573 5535
rect 19592 5515 19600 5535
rect 19489 5493 19600 5515
rect 19068 5444 19099 5490
rect 18856 5441 18891 5442
rect 18835 5434 18891 5441
rect 18835 5414 18864 5434
rect 18884 5414 18891 5434
rect 18835 5409 18891 5414
rect 19068 5437 19107 5444
rect 19068 5417 19074 5437
rect 19099 5417 19107 5437
rect 19068 5411 19107 5417
rect 19282 5437 19314 5444
rect 19282 5417 19288 5437
rect 19309 5417 19314 5437
rect 17641 5328 17688 5346
rect 17896 5336 18800 5371
rect 17897 5335 17931 5336
rect 17558 5269 17610 5274
rect 18013 5269 18058 5271
rect 17558 5254 18058 5269
rect 17558 5201 17572 5254
rect 17603 5230 18058 5254
rect 17603 5229 17628 5230
rect 17603 5201 17610 5229
rect 16588 5169 16665 5172
rect 16555 5154 16665 5169
rect 17280 5184 17461 5190
rect 17280 5164 17291 5184
rect 17311 5164 17461 5184
rect 17558 5177 17610 5201
rect 17280 5158 17461 5164
rect 17284 5156 17319 5158
rect 16299 5098 16360 5100
rect 15997 5069 16360 5098
rect 16840 5091 16872 5098
rect 16840 5071 16847 5091
rect 16868 5071 16872 5091
rect 15997 5067 16299 5069
rect 13777 5051 14776 5054
rect 13777 5049 13812 5051
rect 12799 5026 13211 5028
rect 12801 5025 12841 5026
rect 13179 4961 13211 5026
rect 16840 5006 16872 5071
rect 17210 5006 17250 5007
rect 16840 5004 17252 5006
rect 16239 4981 16274 4983
rect 15275 4978 16274 4981
rect 13752 4963 14054 4965
rect 13179 4941 13183 4961
rect 13204 4941 13211 4961
rect 13179 4934 13211 4941
rect 13691 4934 14054 4963
rect 13691 4932 13752 4934
rect 12732 4874 12767 4876
rect 10485 4842 10562 4845
rect 10452 4827 10562 4842
rect 11181 4857 11218 4862
rect 11181 4837 11188 4857
rect 11208 4837 11218 4857
rect 11181 4830 11218 4837
rect 11987 4835 12025 4869
rect 12590 4868 12771 4874
rect 12590 4848 12740 4868
rect 12760 4848 12771 4868
rect 12590 4842 12771 4848
rect 13386 4863 13496 4878
rect 13386 4860 13463 4863
rect 12423 4835 12473 4839
rect 11181 4829 11216 4830
rect 10218 4729 10226 4758
rect 10255 4729 10266 4758
rect 10218 4724 10266 4729
rect 10737 4764 10769 4771
rect 10737 4744 10744 4764
rect 10765 4744 10769 4764
rect 9252 4707 9284 4714
rect 10737 4679 10769 4744
rect 11107 4679 11147 4680
rect 10737 4677 11149 4679
rect 10737 4651 11117 4677
rect 11143 4651 11149 4677
rect 8805 4641 8840 4649
rect 8253 4612 8295 4622
rect 8805 4621 8813 4641
rect 8833 4621 8840 4641
rect 8805 4616 8840 4621
rect 9459 4636 9569 4651
rect 9459 4633 9536 4636
rect 8253 4611 8294 4612
rect 7887 4577 7922 4578
rect 7866 4570 7922 4577
rect 7866 4550 7895 4570
rect 7915 4550 7922 4570
rect 7866 4545 7922 4550
rect 8313 4573 8345 4580
rect 8313 4553 8319 4573
rect 8340 4553 8345 4573
rect 8805 4564 8839 4616
rect 9459 4606 9462 4633
rect 9491 4609 9536 4633
rect 9565 4609 9569 4636
rect 9491 4606 9569 4609
rect 9459 4592 9569 4606
rect 9755 4636 9797 4646
rect 9755 4617 9763 4636
rect 9788 4617 9797 4636
rect 9755 4564 9797 4617
rect 10737 4643 11149 4651
rect 10737 4615 10769 4643
rect 11182 4623 11216 4829
rect 11987 4825 12473 4835
rect 11498 4803 11609 4825
rect 11498 4783 11506 4803
rect 11525 4783 11583 4803
rect 11602 4783 11609 4803
rect 11987 4793 12436 4825
rect 11498 4766 11609 4783
rect 12423 4772 12436 4793
rect 12467 4772 12473 4825
rect 12423 4755 12473 4772
rect 12120 4696 12154 4697
rect 11251 4661 12155 4696
rect 12363 4686 12410 4704
rect 10737 4595 10742 4615
rect 10763 4595 10769 4615
rect 10737 4588 10769 4595
rect 10944 4615 10983 4621
rect 10944 4595 10952 4615
rect 10977 4595 10983 4615
rect 10944 4588 10983 4595
rect 11160 4618 11216 4623
rect 11160 4598 11167 4618
rect 11187 4598 11216 4618
rect 11160 4591 11216 4598
rect 11160 4590 11195 4591
rect 7866 4339 7900 4545
rect 8313 4525 8345 4553
rect 8803 4538 9799 4564
rect 10952 4542 10983 4588
rect 7933 4517 8345 4525
rect 7933 4491 7939 4517
rect 7965 4491 8345 4517
rect 7933 4489 8345 4491
rect 7935 4488 7975 4489
rect 8095 4453 8134 4468
rect 8095 4412 8106 4453
rect 8127 4412 8134 4453
rect 7865 4331 7901 4339
rect 7865 4311 7874 4331
rect 7894 4311 7901 4331
rect 7865 4310 7901 4311
rect 7865 4299 7899 4310
rect 8095 4139 8134 4412
rect 8313 4424 8345 4489
rect 10451 4517 10562 4539
rect 10451 4497 10459 4517
rect 10478 4497 10536 4517
rect 10555 4497 10562 4517
rect 10951 4525 10983 4542
rect 11252 4525 11289 4661
rect 11390 4628 11500 4642
rect 11390 4625 11468 4628
rect 11390 4598 11394 4625
rect 11423 4601 11468 4625
rect 11497 4601 11500 4628
rect 12120 4618 12154 4661
rect 11423 4598 11500 4601
rect 11390 4583 11500 4598
rect 12119 4613 12154 4618
rect 12119 4593 12126 4613
rect 12146 4593 12154 4613
rect 12119 4585 12154 4593
rect 10951 4512 11289 4525
rect 10451 4480 10562 4497
rect 10952 4493 11289 4512
rect 11231 4492 11289 4493
rect 11675 4520 11707 4527
rect 11675 4500 11682 4520
rect 11703 4500 11707 4520
rect 8313 4404 8317 4424
rect 8338 4404 8345 4424
rect 8313 4397 8345 4404
rect 8731 4431 8789 4432
rect 8731 4412 9068 4431
rect 9458 4427 9569 4444
rect 8731 4399 9069 4412
rect 8235 4335 8288 4338
rect 8235 4318 8247 4335
rect 8279 4318 8288 4335
rect 8235 4310 8288 4318
rect 8234 4263 8288 4310
rect 8520 4326 8630 4341
rect 8520 4323 8597 4326
rect 8520 4296 8523 4323
rect 8552 4299 8597 4323
rect 8626 4299 8630 4326
rect 8552 4296 8630 4299
rect 8520 4282 8630 4296
rect 8731 4263 8768 4399
rect 9037 4382 9069 4399
rect 9458 4407 9465 4427
rect 9484 4407 9542 4427
rect 9561 4407 9569 4427
rect 9458 4385 9569 4407
rect 11675 4435 11707 4500
rect 12045 4435 12085 4436
rect 11675 4433 12087 4435
rect 11675 4407 12055 4433
rect 12081 4407 12087 4433
rect 11675 4399 12087 4407
rect 9037 4336 9068 4382
rect 10221 4360 11217 4386
rect 11675 4371 11707 4399
rect 8825 4333 8860 4334
rect 8804 4326 8860 4333
rect 8804 4306 8833 4326
rect 8853 4306 8860 4326
rect 8804 4301 8860 4306
rect 9037 4329 9076 4336
rect 9037 4309 9043 4329
rect 9068 4309 9076 4329
rect 9037 4303 9076 4309
rect 9251 4329 9283 4336
rect 9251 4309 9257 4329
rect 9278 4309 9283 4329
rect 8234 4228 8769 4263
rect 8234 4224 8287 4228
rect 8095 4112 8099 4139
rect 8130 4112 8134 4139
rect 8380 4160 8491 4177
rect 8380 4140 8387 4160
rect 8406 4140 8464 4160
rect 8483 4140 8491 4160
rect 8380 4118 8491 4140
rect 8095 4105 8134 4112
rect 8804 4095 8838 4301
rect 9251 4281 9283 4309
rect 8871 4273 9283 4281
rect 10223 4307 10265 4360
rect 10223 4288 10232 4307
rect 10257 4288 10265 4307
rect 10223 4278 10265 4288
rect 10451 4318 10561 4332
rect 10451 4315 10529 4318
rect 10451 4288 10455 4315
rect 10484 4291 10529 4315
rect 10558 4291 10561 4318
rect 11181 4308 11215 4360
rect 11675 4351 11680 4371
rect 11701 4351 11707 4371
rect 11675 4344 11707 4351
rect 11885 4372 11923 4382
rect 12120 4379 12154 4585
rect 11885 4355 11895 4372
rect 11915 4355 11923 4372
rect 11726 4312 11767 4313
rect 10484 4288 10561 4291
rect 10451 4273 10561 4288
rect 11180 4303 11215 4308
rect 11180 4283 11187 4303
rect 11207 4283 11215 4303
rect 11725 4302 11767 4312
rect 11180 4275 11215 4283
rect 8871 4247 8877 4273
rect 8903 4247 9283 4273
rect 8871 4245 9283 4247
rect 8873 4244 8913 4245
rect 9251 4180 9283 4245
rect 10736 4210 10768 4217
rect 9251 4160 9255 4180
rect 9276 4160 9283 4180
rect 9251 4153 9283 4160
rect 9754 4195 9802 4200
rect 9754 4166 9765 4195
rect 9794 4166 9802 4195
rect 8804 4094 8839 4095
rect 8802 4087 8839 4094
rect 7747 4066 7782 4067
rect 7724 4059 7782 4066
rect 7724 4039 7755 4059
rect 7775 4039 7782 4059
rect 7724 4034 7782 4039
rect 8173 4062 8205 4069
rect 8173 4042 8179 4062
rect 8200 4042 8205 4062
rect 7724 3886 7760 4034
rect 8173 4014 8205 4042
rect 7793 4006 8205 4014
rect 7793 3980 7799 4006
rect 7825 3980 8205 4006
rect 8802 4067 8812 4087
rect 8832 4067 8839 4087
rect 8802 4062 8839 4067
rect 9458 4082 9568 4097
rect 9458 4079 9535 4082
rect 8802 4011 8837 4062
rect 9458 4052 9461 4079
rect 9490 4055 9535 4079
rect 9564 4055 9568 4082
rect 9490 4052 9568 4055
rect 9458 4038 9568 4052
rect 9754 4011 9802 4166
rect 10736 4190 10743 4210
rect 10764 4190 10768 4210
rect 10736 4125 10768 4190
rect 11106 4125 11146 4126
rect 10736 4123 11148 4125
rect 10736 4097 11116 4123
rect 11142 4097 11148 4123
rect 10736 4089 11148 4097
rect 10736 4061 10768 4089
rect 11181 4069 11215 4275
rect 11389 4273 11500 4295
rect 11389 4253 11397 4273
rect 11416 4253 11474 4273
rect 11493 4253 11500 4273
rect 11389 4236 11500 4253
rect 11725 4280 11732 4302
rect 11758 4280 11767 4302
rect 11725 4271 11767 4280
rect 10942 4066 10985 4068
rect 10736 4041 10741 4061
rect 10762 4041 10768 4061
rect 10736 4034 10768 4041
rect 10941 4059 10985 4066
rect 10941 4039 10951 4059
rect 10974 4039 10985 4059
rect 10941 4035 10985 4039
rect 11159 4064 11215 4069
rect 11159 4044 11166 4064
rect 11186 4044 11215 4064
rect 11159 4037 11215 4044
rect 11271 4205 11304 4206
rect 11725 4205 11762 4271
rect 11271 4176 11762 4205
rect 11159 4036 11194 4037
rect 8802 3987 9802 4011
rect 8802 3984 9801 3987
rect 8802 3982 8837 3984
rect 7793 3978 8205 3980
rect 7795 3977 7835 3978
rect 7727 3828 7760 3886
rect 7957 3938 7995 3948
rect 7957 3900 7966 3938
rect 7989 3900 7995 3938
rect 7727 3820 7761 3828
rect 7727 3800 7734 3820
rect 7754 3800 7761 3820
rect 7727 3795 7761 3800
rect 7727 3794 7758 3795
rect 7957 3764 7995 3900
rect 8173 3913 8205 3978
rect 10450 3963 10561 3985
rect 10450 3943 10458 3963
rect 10477 3943 10535 3963
rect 10554 3943 10561 3963
rect 10450 3926 10561 3943
rect 10941 3954 10983 4035
rect 11271 3956 11304 4176
rect 11725 4174 11762 4176
rect 11531 4036 11641 4050
rect 11531 4033 11609 4036
rect 11531 4006 11535 4033
rect 11564 4009 11609 4033
rect 11638 4009 11641 4036
rect 11564 4006 11641 4009
rect 11531 3991 11641 4006
rect 11885 4017 11923 4355
rect 12098 4374 12154 4379
rect 12098 4354 12105 4374
rect 12125 4354 12154 4374
rect 12098 4347 12154 4354
rect 12363 4646 12370 4686
rect 12397 4646 12410 4686
rect 12593 4664 12640 4842
rect 13386 4833 13389 4860
rect 13418 4836 13463 4860
rect 13492 4836 13496 4863
rect 13418 4833 13496 4836
rect 13386 4819 13496 4833
rect 12098 4346 12133 4347
rect 12263 4026 12295 4027
rect 11885 4000 11893 4017
rect 11913 4000 11923 4017
rect 11885 3994 11923 4000
rect 12260 4021 12295 4026
rect 12260 4001 12267 4021
rect 12287 4001 12295 4021
rect 12260 3993 12295 4001
rect 11243 3954 11304 3956
rect 10941 3925 11304 3954
rect 11816 3928 11848 3935
rect 10941 3923 11243 3925
rect 8173 3893 8177 3913
rect 8198 3893 8205 3913
rect 11816 3908 11823 3928
rect 11844 3908 11848 3928
rect 8778 3896 9080 3898
rect 8173 3886 8205 3893
rect 8717 3867 9080 3896
rect 8717 3865 8778 3867
rect 8098 3821 8136 3827
rect 8098 3804 8108 3821
rect 8128 3804 8136 3821
rect 7957 3610 8001 3764
rect 7794 3608 8001 3610
rect 7770 3575 8001 3608
rect 6867 2949 6871 2969
rect 6892 2949 6901 2969
rect 6867 2943 6901 2949
rect 7020 3080 7349 3083
rect 7388 3080 7432 3105
rect 7020 3050 7432 3080
rect 6269 2887 6330 2889
rect 5967 2858 6330 2887
rect 6811 2874 6843 2881
rect 5967 2856 6269 2858
rect 6811 2854 6818 2874
rect 6839 2854 6843 2874
rect 3747 2840 4746 2843
rect 3747 2838 3782 2840
rect 2768 2821 3180 2823
rect 2770 2820 2810 2821
rect 3148 2756 3180 2821
rect 6811 2789 6843 2854
rect 7020 2862 7055 3050
rect 7322 3048 7432 3050
rect 7615 3063 7665 3191
rect 7770 3174 7820 3575
rect 7957 3571 8001 3575
rect 7888 3474 7923 3475
rect 7750 3165 7820 3174
rect 7750 3136 7765 3165
rect 7813 3157 7820 3165
rect 7867 3467 7923 3474
rect 7867 3447 7896 3467
rect 7916 3447 7923 3467
rect 7867 3442 7923 3447
rect 8098 3466 8136 3804
rect 8380 3815 8490 3830
rect 8380 3812 8457 3815
rect 8380 3785 8383 3812
rect 8412 3788 8457 3812
rect 8486 3788 8490 3815
rect 8412 3785 8490 3788
rect 8380 3771 8490 3785
rect 8259 3645 8296 3647
rect 8717 3645 8750 3865
rect 9038 3786 9080 3867
rect 9460 3878 9571 3895
rect 9460 3858 9467 3878
rect 9486 3858 9544 3878
rect 9563 3858 9571 3878
rect 9460 3836 9571 3858
rect 11816 3843 11848 3908
rect 12186 3843 12226 3844
rect 11816 3841 12228 3843
rect 11184 3837 11219 3839
rect 10220 3834 11219 3837
rect 10219 3810 11219 3834
rect 8827 3784 8862 3785
rect 8259 3616 8750 3645
rect 8259 3550 8296 3616
rect 8717 3615 8750 3616
rect 8806 3777 8862 3784
rect 8806 3757 8835 3777
rect 8855 3757 8862 3777
rect 8806 3752 8862 3757
rect 9036 3782 9080 3786
rect 9036 3762 9047 3782
rect 9070 3762 9080 3782
rect 9036 3755 9080 3762
rect 9253 3780 9285 3787
rect 9253 3760 9259 3780
rect 9280 3760 9285 3780
rect 9036 3753 9079 3755
rect 8254 3541 8296 3550
rect 8254 3519 8263 3541
rect 8289 3519 8296 3541
rect 8521 3568 8632 3585
rect 8521 3548 8528 3568
rect 8547 3548 8605 3568
rect 8624 3548 8632 3568
rect 8521 3526 8632 3548
rect 8806 3546 8840 3752
rect 9253 3732 9285 3760
rect 8873 3724 9285 3732
rect 8873 3698 8879 3724
rect 8905 3698 9285 3724
rect 8873 3696 9285 3698
rect 8875 3695 8915 3696
rect 9253 3631 9285 3696
rect 9253 3611 9257 3631
rect 9278 3611 9285 3631
rect 10219 3655 10267 3810
rect 10453 3769 10563 3783
rect 10453 3766 10531 3769
rect 10453 3739 10457 3766
rect 10486 3742 10531 3766
rect 10560 3742 10563 3769
rect 11184 3759 11219 3810
rect 10486 3739 10563 3742
rect 10453 3724 10563 3739
rect 11182 3754 11219 3759
rect 11182 3734 11189 3754
rect 11209 3734 11219 3754
rect 11816 3815 12196 3841
rect 12222 3815 12228 3841
rect 11816 3807 12228 3815
rect 11816 3779 11848 3807
rect 11816 3759 11821 3779
rect 11842 3759 11848 3779
rect 11816 3752 11848 3759
rect 12022 3778 12064 3789
rect 12261 3787 12295 3993
rect 12022 3757 12029 3778
rect 12056 3757 12064 3778
rect 11182 3727 11219 3734
rect 11182 3726 11217 3727
rect 10219 3626 10227 3655
rect 10256 3626 10267 3655
rect 10219 3621 10267 3626
rect 10738 3661 10770 3668
rect 10738 3641 10745 3661
rect 10766 3641 10770 3661
rect 9253 3604 9285 3611
rect 10738 3576 10770 3641
rect 11108 3576 11148 3577
rect 10738 3574 11150 3576
rect 10738 3548 11118 3574
rect 11144 3548 11150 3574
rect 8806 3538 8841 3546
rect 8254 3509 8296 3519
rect 8806 3518 8814 3538
rect 8834 3518 8841 3538
rect 8806 3513 8841 3518
rect 9460 3533 9570 3548
rect 9460 3530 9537 3533
rect 8254 3508 8295 3509
rect 8098 3449 8106 3466
rect 8126 3449 8136 3466
rect 7867 3236 7901 3442
rect 8098 3439 8136 3449
rect 8314 3470 8346 3477
rect 8314 3450 8320 3470
rect 8341 3450 8346 3470
rect 8806 3461 8840 3513
rect 9460 3503 9463 3530
rect 9492 3506 9537 3530
rect 9566 3506 9570 3533
rect 9492 3503 9570 3506
rect 9460 3489 9570 3503
rect 9756 3533 9798 3543
rect 9756 3514 9764 3533
rect 9789 3514 9798 3533
rect 9756 3461 9798 3514
rect 10738 3540 11150 3548
rect 10738 3512 10770 3540
rect 11183 3520 11217 3726
rect 11887 3709 11926 3716
rect 11530 3681 11641 3703
rect 11530 3661 11538 3681
rect 11557 3661 11615 3681
rect 11634 3661 11641 3681
rect 11530 3644 11641 3661
rect 11887 3682 11891 3709
rect 11922 3682 11926 3709
rect 11734 3593 11787 3597
rect 11252 3558 11787 3593
rect 10738 3492 10743 3512
rect 10764 3492 10770 3512
rect 10738 3485 10770 3492
rect 10945 3512 10984 3518
rect 10945 3492 10953 3512
rect 10978 3492 10984 3512
rect 10945 3485 10984 3492
rect 11161 3515 11217 3520
rect 11161 3495 11168 3515
rect 11188 3495 11217 3515
rect 11161 3488 11217 3495
rect 11161 3487 11196 3488
rect 8314 3422 8346 3450
rect 8804 3435 9800 3461
rect 10953 3439 10984 3485
rect 7934 3414 8346 3422
rect 7934 3388 7940 3414
rect 7966 3388 8346 3414
rect 7934 3386 8346 3388
rect 7936 3385 7976 3386
rect 8314 3321 8346 3386
rect 10452 3414 10563 3436
rect 10452 3394 10460 3414
rect 10479 3394 10537 3414
rect 10556 3394 10563 3414
rect 10952 3422 10984 3439
rect 11253 3422 11290 3558
rect 11391 3525 11501 3539
rect 11391 3522 11469 3525
rect 11391 3495 11395 3522
rect 11424 3498 11469 3522
rect 11498 3498 11501 3525
rect 11424 3495 11501 3498
rect 11391 3480 11501 3495
rect 11733 3511 11787 3558
rect 11733 3503 11786 3511
rect 11733 3486 11742 3503
rect 11774 3486 11786 3503
rect 11733 3483 11786 3486
rect 10952 3409 11290 3422
rect 10452 3377 10563 3394
rect 10953 3390 11290 3409
rect 11232 3389 11290 3390
rect 11676 3417 11708 3424
rect 11676 3397 11683 3417
rect 11704 3397 11708 3417
rect 8314 3301 8318 3321
rect 8339 3301 8346 3321
rect 8314 3294 8346 3301
rect 8732 3328 8790 3329
rect 8732 3309 9069 3328
rect 9459 3324 9570 3341
rect 8732 3296 9070 3309
rect 7867 3228 7902 3236
rect 7867 3208 7875 3228
rect 7895 3208 7902 3228
rect 7867 3203 7902 3208
rect 8521 3223 8631 3238
rect 8521 3220 8598 3223
rect 7867 3160 7901 3203
rect 8521 3193 8524 3220
rect 8553 3196 8598 3220
rect 8627 3196 8631 3223
rect 8553 3193 8631 3196
rect 8521 3179 8631 3193
rect 8732 3160 8769 3296
rect 9038 3279 9070 3296
rect 9459 3304 9466 3324
rect 9485 3304 9543 3324
rect 9562 3304 9570 3324
rect 9459 3282 9570 3304
rect 11676 3332 11708 3397
rect 11887 3409 11926 3682
rect 12022 3586 12064 3757
rect 12239 3782 12295 3787
rect 12239 3762 12246 3782
rect 12266 3762 12295 3782
rect 12239 3755 12295 3762
rect 12239 3754 12274 3755
rect 12022 3552 12266 3586
rect 12229 3544 12266 3552
rect 12122 3511 12156 3522
rect 12120 3510 12156 3511
rect 12120 3490 12127 3510
rect 12147 3490 12156 3510
rect 12120 3482 12156 3490
rect 11887 3368 11894 3409
rect 11915 3368 11926 3409
rect 11887 3353 11926 3368
rect 12046 3332 12086 3333
rect 11676 3330 12088 3332
rect 11676 3304 12056 3330
rect 12082 3304 12088 3330
rect 11676 3296 12088 3304
rect 9038 3233 9069 3279
rect 10222 3257 11218 3283
rect 11676 3268 11708 3296
rect 12121 3276 12155 3482
rect 8826 3230 8861 3231
rect 8805 3223 8861 3230
rect 8805 3203 8834 3223
rect 8854 3203 8861 3223
rect 8805 3198 8861 3203
rect 9038 3226 9077 3233
rect 9038 3206 9044 3226
rect 9069 3206 9077 3226
rect 9038 3200 9077 3206
rect 9252 3226 9284 3233
rect 9252 3206 9258 3226
rect 9279 3206 9284 3226
rect 7813 3136 7818 3157
rect 7750 3125 7818 3136
rect 7866 3125 8770 3160
rect 7867 3124 7901 3125
rect 7615 3029 8030 3063
rect 7615 3027 7665 3029
rect 7248 2965 7298 2972
rect 7248 2951 7262 2965
rect 7254 2947 7262 2951
rect 7282 2951 7298 2965
rect 7282 2947 7292 2951
rect 7778 2950 7813 2951
rect 7254 2940 7292 2947
rect 7757 2943 7813 2950
rect 7255 2939 7290 2940
rect 7020 2830 7025 2862
rect 7052 2830 7055 2862
rect 7020 2812 7055 2830
rect 7181 2789 7221 2790
rect 6811 2787 7223 2789
rect 6209 2770 6244 2772
rect 5245 2767 6244 2770
rect 3148 2736 3152 2756
rect 3173 2736 3180 2756
rect 3722 2752 4024 2754
rect 3148 2729 3180 2736
rect 3661 2723 4024 2752
rect 3661 2721 3722 2723
rect 2701 2670 2736 2671
rect 2178 2660 2234 2667
rect 2699 2663 2737 2670
rect 2178 2659 2213 2660
rect 455 2631 532 2634
rect 422 2616 532 2631
rect 1151 2646 1188 2651
rect 1151 2626 1158 2646
rect 1178 2626 1188 2646
rect 2699 2643 2709 2663
rect 2729 2643 2737 2663
rect 1151 2619 1188 2626
rect 2173 2621 2243 2631
rect 1151 2618 1186 2619
rect 188 2518 196 2547
rect 225 2518 236 2547
rect 188 2513 236 2518
rect 707 2553 739 2560
rect 707 2533 714 2553
rect 735 2533 739 2553
rect 707 2468 739 2533
rect 1077 2468 1117 2469
rect 707 2466 1119 2468
rect 707 2440 1087 2466
rect 1113 2440 1119 2466
rect 707 2432 1119 2440
rect 707 2404 739 2432
rect 1152 2412 1186 2618
rect 2171 2614 2243 2621
rect 1469 2586 1580 2608
rect 1469 2566 1477 2586
rect 1496 2566 1554 2586
rect 1573 2566 1580 2586
rect 1469 2549 1580 2566
rect 2171 2585 2178 2614
rect 2226 2585 2243 2614
rect 2171 2576 2243 2585
rect 2090 2485 2124 2486
rect 1221 2450 2125 2485
rect 707 2384 712 2404
rect 733 2384 739 2404
rect 707 2377 739 2384
rect 914 2404 953 2410
rect 914 2384 922 2404
rect 947 2384 953 2404
rect 914 2377 953 2384
rect 1130 2407 1186 2412
rect 1130 2387 1137 2407
rect 1157 2387 1186 2407
rect 1130 2380 1186 2387
rect 1130 2379 1165 2380
rect 922 2331 953 2377
rect 421 2306 532 2328
rect 421 2286 429 2306
rect 448 2286 506 2306
rect 525 2286 532 2306
rect 921 2314 953 2331
rect 1222 2314 1259 2450
rect 1360 2417 1470 2431
rect 1360 2414 1438 2417
rect 1360 2387 1364 2414
rect 1393 2390 1438 2414
rect 1467 2390 1470 2417
rect 2090 2407 2124 2450
rect 1393 2387 1470 2390
rect 1360 2372 1470 2387
rect 2089 2402 2124 2407
rect 2089 2382 2096 2402
rect 2116 2382 2124 2402
rect 2089 2374 2124 2382
rect 921 2301 1259 2314
rect 421 2269 532 2286
rect 922 2282 1259 2301
rect 1201 2281 1259 2282
rect 1645 2309 1677 2316
rect 1645 2289 1652 2309
rect 1673 2289 1677 2309
rect 1645 2224 1677 2289
rect 2015 2224 2055 2225
rect 1645 2222 2057 2224
rect 1645 2196 2025 2222
rect 2051 2196 2057 2222
rect 1645 2188 2057 2196
rect 191 2149 1187 2175
rect 1645 2160 1677 2188
rect 193 2096 235 2149
rect 193 2077 202 2096
rect 227 2077 235 2096
rect 193 2067 235 2077
rect 421 2107 531 2121
rect 421 2104 499 2107
rect 421 2077 425 2104
rect 454 2080 499 2104
rect 528 2080 531 2107
rect 1151 2097 1185 2149
rect 1645 2140 1650 2160
rect 1671 2140 1677 2160
rect 1645 2133 1677 2140
rect 1855 2161 1893 2171
rect 2090 2168 2124 2374
rect 1855 2144 1865 2161
rect 1885 2144 1893 2161
rect 1696 2101 1737 2102
rect 454 2077 531 2080
rect 421 2062 531 2077
rect 1150 2092 1185 2097
rect 1150 2072 1157 2092
rect 1177 2072 1185 2092
rect 1695 2091 1737 2101
rect 1150 2064 1185 2072
rect 706 1999 738 2006
rect 706 1979 713 1999
rect 734 1979 738 1999
rect 706 1914 738 1979
rect 1076 1914 1116 1915
rect 706 1912 1118 1914
rect 706 1886 1086 1912
rect 1112 1886 1118 1912
rect 706 1878 1118 1886
rect 706 1850 738 1878
rect 1151 1858 1185 2064
rect 1359 2062 1470 2084
rect 1359 2042 1367 2062
rect 1386 2042 1444 2062
rect 1463 2042 1470 2062
rect 1359 2025 1470 2042
rect 1695 2069 1702 2091
rect 1728 2069 1737 2091
rect 1695 2060 1737 2069
rect 912 1855 955 1857
rect 706 1830 711 1850
rect 732 1830 738 1850
rect 706 1823 738 1830
rect 911 1848 955 1855
rect 911 1828 921 1848
rect 944 1828 955 1848
rect 911 1824 955 1828
rect 1129 1853 1185 1858
rect 1129 1833 1136 1853
rect 1156 1833 1185 1853
rect 1129 1826 1185 1833
rect 1241 1994 1274 1995
rect 1695 1994 1732 2060
rect 1241 1965 1732 1994
rect 1129 1825 1164 1826
rect 420 1752 531 1774
rect 420 1732 428 1752
rect 447 1732 505 1752
rect 524 1732 531 1752
rect 420 1715 531 1732
rect 911 1743 953 1824
rect 1241 1745 1274 1965
rect 1695 1963 1732 1965
rect 1501 1825 1611 1839
rect 1501 1822 1579 1825
rect 1501 1795 1505 1822
rect 1534 1798 1579 1822
rect 1608 1798 1611 1825
rect 1534 1795 1611 1798
rect 1501 1780 1611 1795
rect 1855 1806 1893 2144
rect 2068 2163 2124 2168
rect 2068 2143 2075 2163
rect 2095 2143 2124 2163
rect 2068 2136 2124 2143
rect 2068 2135 2103 2136
rect 1990 2035 2034 2039
rect 2171 2035 2221 2576
rect 1990 2002 2221 2035
rect 2699 2030 2737 2643
rect 3355 2658 3465 2673
rect 3355 2655 3432 2658
rect 3355 2628 3358 2655
rect 3387 2631 3432 2655
rect 3461 2631 3465 2658
rect 3387 2628 3465 2631
rect 3355 2614 3465 2628
rect 3203 2501 3240 2503
rect 3661 2501 3694 2721
rect 3982 2642 4024 2723
rect 4404 2734 4515 2750
rect 4404 2714 4411 2734
rect 4430 2714 4488 2734
rect 4507 2714 4515 2734
rect 4404 2692 4515 2714
rect 5244 2743 6244 2767
rect 3771 2640 3806 2641
rect 3203 2472 3694 2501
rect 3203 2406 3240 2472
rect 3661 2471 3694 2472
rect 3750 2633 3806 2640
rect 3750 2613 3779 2633
rect 3799 2613 3806 2633
rect 3750 2608 3806 2613
rect 3980 2638 4024 2642
rect 3980 2618 3991 2638
rect 4014 2618 4024 2638
rect 3980 2611 4024 2618
rect 4197 2636 4229 2643
rect 4197 2616 4203 2636
rect 4224 2616 4229 2636
rect 3980 2609 4023 2611
rect 3198 2397 3240 2406
rect 3198 2375 3207 2397
rect 3233 2375 3240 2397
rect 3465 2424 3576 2441
rect 3465 2404 3472 2424
rect 3491 2404 3549 2424
rect 3568 2404 3576 2424
rect 3465 2382 3576 2404
rect 3750 2402 3784 2608
rect 4197 2588 4229 2616
rect 3817 2580 4229 2588
rect 3817 2554 3823 2580
rect 3849 2554 4229 2580
rect 5244 2588 5292 2743
rect 5478 2702 5588 2716
rect 5478 2699 5556 2702
rect 5478 2672 5482 2699
rect 5511 2675 5556 2699
rect 5585 2675 5588 2702
rect 6209 2692 6244 2743
rect 6811 2761 7191 2787
rect 7217 2761 7223 2787
rect 6811 2753 7223 2761
rect 6811 2725 6843 2753
rect 7256 2733 7290 2939
rect 6811 2705 6816 2725
rect 6837 2705 6843 2725
rect 6811 2698 6843 2705
rect 7234 2728 7290 2733
rect 7234 2708 7241 2728
rect 7261 2708 7290 2728
rect 7757 2923 7786 2943
rect 7806 2923 7813 2943
rect 7757 2918 7813 2923
rect 7985 2946 8030 3029
rect 8411 3044 8522 3061
rect 8411 3024 8418 3044
rect 8437 3024 8495 3044
rect 8514 3024 8522 3044
rect 8411 3002 8522 3024
rect 8805 2992 8839 3198
rect 9252 3178 9284 3206
rect 8872 3170 9284 3178
rect 10224 3204 10266 3257
rect 10224 3185 10233 3204
rect 10258 3185 10266 3204
rect 10224 3175 10266 3185
rect 10452 3215 10562 3229
rect 10452 3212 10530 3215
rect 10452 3185 10456 3212
rect 10485 3188 10530 3212
rect 10559 3188 10562 3215
rect 11182 3205 11216 3257
rect 11676 3248 11681 3268
rect 11702 3248 11708 3268
rect 11676 3241 11708 3248
rect 12099 3271 12155 3276
rect 12099 3251 12106 3271
rect 12126 3251 12155 3271
rect 12099 3244 12155 3251
rect 12099 3243 12134 3244
rect 11727 3209 11768 3210
rect 10485 3185 10562 3188
rect 10452 3170 10562 3185
rect 11181 3200 11216 3205
rect 11181 3180 11188 3200
rect 11208 3180 11216 3200
rect 11726 3199 11768 3209
rect 11181 3172 11216 3180
rect 8872 3144 8878 3170
rect 8904 3144 9284 3170
rect 8872 3142 9284 3144
rect 8874 3141 8914 3142
rect 9252 3077 9284 3142
rect 10737 3107 10769 3114
rect 9252 3057 9256 3077
rect 9277 3057 9284 3077
rect 9252 3050 9284 3057
rect 9755 3092 9803 3097
rect 9755 3063 9766 3092
rect 9795 3063 9803 3092
rect 8805 2991 8840 2992
rect 8803 2984 8840 2991
rect 8803 2964 8813 2984
rect 8833 2964 8840 2984
rect 8803 2959 8840 2964
rect 9459 2979 9569 2994
rect 9459 2976 9536 2979
rect 7985 2927 7994 2946
rect 8023 2927 8030 2946
rect 7757 2712 7791 2918
rect 7985 2915 8030 2927
rect 8204 2946 8236 2953
rect 8204 2926 8210 2946
rect 8231 2926 8236 2946
rect 8204 2898 8236 2926
rect 7824 2890 8236 2898
rect 7824 2864 7830 2890
rect 7856 2864 8236 2890
rect 8803 2908 8838 2959
rect 9459 2949 9462 2976
rect 9491 2952 9536 2976
rect 9565 2952 9569 2979
rect 9491 2949 9569 2952
rect 9459 2935 9569 2949
rect 9755 2908 9803 3063
rect 10737 3087 10744 3107
rect 10765 3087 10769 3107
rect 10737 3022 10769 3087
rect 11107 3022 11147 3023
rect 10737 3020 11149 3022
rect 10737 2994 11117 3020
rect 11143 2994 11149 3020
rect 10737 2986 11149 2994
rect 10737 2958 10769 2986
rect 11182 2966 11216 3172
rect 11390 3170 11501 3192
rect 11390 3150 11398 3170
rect 11417 3150 11475 3170
rect 11494 3150 11501 3170
rect 11390 3133 11501 3150
rect 11726 3177 11733 3199
rect 11759 3177 11768 3199
rect 11726 3168 11768 3177
rect 10943 2963 10986 2965
rect 10737 2938 10742 2958
rect 10763 2938 10769 2958
rect 10737 2931 10769 2938
rect 10942 2956 10986 2963
rect 10942 2936 10952 2956
rect 10975 2936 10986 2956
rect 10942 2932 10986 2936
rect 11160 2961 11216 2966
rect 11160 2941 11167 2961
rect 11187 2941 11216 2961
rect 11160 2934 11216 2941
rect 11272 3102 11305 3103
rect 11726 3102 11763 3168
rect 12229 3153 12267 3544
rect 11843 3137 12267 3153
rect 11272 3073 11763 3102
rect 11160 2933 11195 2934
rect 8803 2884 9803 2908
rect 8803 2881 9802 2884
rect 8803 2879 8838 2881
rect 7824 2862 8236 2864
rect 7826 2861 7866 2862
rect 8204 2797 8236 2862
rect 10451 2860 10562 2882
rect 10451 2840 10459 2860
rect 10478 2840 10536 2860
rect 10555 2840 10562 2860
rect 10451 2824 10562 2840
rect 10942 2851 10984 2932
rect 11272 2853 11305 3073
rect 11726 3071 11763 3073
rect 11842 3112 12267 3137
rect 11501 2946 11611 2960
rect 11501 2943 11579 2946
rect 11501 2916 11505 2943
rect 11534 2919 11579 2943
rect 11608 2919 11611 2946
rect 11534 2916 11611 2919
rect 11501 2901 11611 2916
rect 11842 2933 11876 3112
rect 12363 3069 12410 4646
rect 12592 4640 12640 4664
rect 13233 4712 13270 4714
rect 13691 4712 13724 4932
rect 14012 4853 14054 4934
rect 14434 4945 14545 4962
rect 14434 4925 14441 4945
rect 14460 4925 14518 4945
rect 14537 4925 14545 4945
rect 14434 4903 14545 4925
rect 15274 4954 16274 4978
rect 13801 4851 13836 4852
rect 13233 4683 13724 4712
rect 12592 3155 12638 4640
rect 13233 4617 13270 4683
rect 13691 4682 13724 4683
rect 13780 4844 13836 4851
rect 13780 4824 13809 4844
rect 13829 4824 13836 4844
rect 13780 4819 13836 4824
rect 14010 4849 14054 4853
rect 14010 4829 14021 4849
rect 14044 4829 14054 4849
rect 14010 4822 14054 4829
rect 14227 4847 14259 4854
rect 14227 4827 14233 4847
rect 14254 4827 14259 4847
rect 14010 4820 14053 4822
rect 13228 4608 13270 4617
rect 13228 4586 13237 4608
rect 13263 4586 13270 4608
rect 13495 4635 13606 4652
rect 13495 4615 13502 4635
rect 13521 4615 13579 4635
rect 13598 4615 13606 4635
rect 13495 4593 13606 4615
rect 13780 4613 13814 4819
rect 14227 4799 14259 4827
rect 13847 4791 14259 4799
rect 13847 4765 13853 4791
rect 13879 4765 14259 4791
rect 15274 4799 15322 4954
rect 15508 4913 15618 4927
rect 15508 4910 15586 4913
rect 15508 4883 15512 4910
rect 15541 4886 15586 4910
rect 15615 4886 15618 4913
rect 16239 4903 16274 4954
rect 16840 4978 17220 5004
rect 17246 4978 17252 5004
rect 16840 4970 17252 4978
rect 16840 4942 16872 4970
rect 17285 4950 17319 5156
rect 17809 5155 17844 5156
rect 16840 4922 16845 4942
rect 16866 4922 16872 4942
rect 16840 4915 16872 4922
rect 17042 4945 17087 4950
rect 17042 4921 17053 4945
rect 17079 4921 17087 4945
rect 17042 4910 17087 4921
rect 17263 4945 17319 4950
rect 17263 4925 17270 4945
rect 17290 4925 17319 4945
rect 17263 4918 17319 4925
rect 17788 5148 17844 5155
rect 17788 5128 17817 5148
rect 17837 5128 17844 5148
rect 17788 5123 17844 5128
rect 18013 5151 18058 5230
rect 18442 5249 18553 5266
rect 18442 5229 18449 5249
rect 18468 5229 18526 5249
rect 18545 5229 18553 5249
rect 18442 5207 18553 5229
rect 18835 5203 18869 5409
rect 19282 5389 19314 5417
rect 18902 5381 19314 5389
rect 18902 5355 18908 5381
rect 18934 5355 19314 5381
rect 18902 5353 19314 5355
rect 18904 5352 18944 5353
rect 19282 5288 19314 5353
rect 19282 5268 19286 5288
rect 19307 5268 19314 5288
rect 19282 5261 19314 5268
rect 19785 5303 19833 5308
rect 19785 5274 19796 5303
rect 19825 5274 19833 5303
rect 18835 5202 18870 5203
rect 18833 5195 18870 5202
rect 18833 5175 18843 5195
rect 18863 5175 18870 5195
rect 18833 5170 18870 5175
rect 19489 5190 19599 5205
rect 19489 5187 19566 5190
rect 18013 5131 18024 5151
rect 18049 5131 18058 5151
rect 18013 5127 18058 5131
rect 18235 5151 18267 5158
rect 18235 5131 18241 5151
rect 18262 5131 18267 5151
rect 17263 4917 17298 4918
rect 17788 4917 17822 5123
rect 18235 5103 18267 5131
rect 17855 5095 18267 5103
rect 17855 5069 17861 5095
rect 17887 5069 18267 5095
rect 18833 5119 18868 5170
rect 19489 5160 19492 5187
rect 19521 5163 19566 5187
rect 19595 5163 19599 5190
rect 19521 5160 19599 5163
rect 19489 5146 19599 5160
rect 19785 5119 19833 5274
rect 18833 5095 19833 5119
rect 18833 5092 19832 5095
rect 18833 5090 18868 5092
rect 17855 5067 18267 5069
rect 17857 5066 17897 5067
rect 18235 5002 18267 5067
rect 18808 5004 19110 5006
rect 18235 4982 18239 5002
rect 18260 4982 18267 5002
rect 18235 4975 18267 4982
rect 18747 4975 19110 5004
rect 18747 4973 18808 4975
rect 17788 4915 17823 4917
rect 15541 4883 15618 4886
rect 15508 4868 15618 4883
rect 16237 4898 16274 4903
rect 16237 4878 16244 4898
rect 16264 4878 16274 4898
rect 16237 4871 16274 4878
rect 17043 4876 17081 4910
rect 17646 4909 17827 4915
rect 17646 4889 17796 4909
rect 17816 4889 17827 4909
rect 17646 4883 17827 4889
rect 18442 4904 18552 4919
rect 18442 4901 18519 4904
rect 17479 4876 17529 4880
rect 16237 4870 16272 4871
rect 15274 4770 15282 4799
rect 15311 4770 15322 4799
rect 15274 4765 15322 4770
rect 15793 4805 15825 4812
rect 15793 4785 15800 4805
rect 15821 4785 15825 4805
rect 13847 4763 14259 4765
rect 13849 4762 13889 4763
rect 14227 4698 14259 4763
rect 14227 4678 14231 4698
rect 14252 4678 14259 4698
rect 14227 4671 14259 4678
rect 15793 4720 15825 4785
rect 16163 4720 16203 4721
rect 15793 4718 16205 4720
rect 15793 4692 16173 4718
rect 16199 4692 16205 4718
rect 15793 4684 16205 4692
rect 15793 4656 15825 4684
rect 16238 4664 16272 4870
rect 17043 4866 17529 4876
rect 16554 4844 16665 4866
rect 16554 4824 16562 4844
rect 16581 4824 16639 4844
rect 16658 4824 16665 4844
rect 17043 4834 17492 4866
rect 16554 4807 16665 4824
rect 17479 4813 17492 4834
rect 17523 4813 17529 4866
rect 17479 4796 17529 4813
rect 17176 4737 17210 4738
rect 16307 4702 17211 4737
rect 17419 4727 17466 4745
rect 15793 4636 15798 4656
rect 15819 4636 15825 4656
rect 15793 4629 15825 4636
rect 16000 4656 16039 4662
rect 16000 4636 16008 4656
rect 16033 4636 16039 4656
rect 16000 4629 16039 4636
rect 16216 4659 16272 4664
rect 16216 4639 16223 4659
rect 16243 4639 16272 4659
rect 16216 4632 16272 4639
rect 16216 4631 16251 4632
rect 13780 4605 13815 4613
rect 13228 4576 13270 4586
rect 13780 4585 13788 4605
rect 13808 4585 13815 4605
rect 13780 4580 13815 4585
rect 14434 4600 14544 4615
rect 14434 4597 14511 4600
rect 13228 4575 13269 4576
rect 12862 4541 12897 4542
rect 12841 4534 12897 4541
rect 12841 4514 12870 4534
rect 12890 4514 12897 4534
rect 12841 4509 12897 4514
rect 13288 4537 13320 4544
rect 13288 4517 13294 4537
rect 13315 4517 13320 4537
rect 13780 4528 13814 4580
rect 14434 4570 14437 4597
rect 14466 4573 14511 4597
rect 14540 4573 14544 4600
rect 14466 4570 14544 4573
rect 14434 4556 14544 4570
rect 14730 4600 14772 4610
rect 14730 4581 14738 4600
rect 14763 4581 14772 4600
rect 16008 4583 16039 4629
rect 14730 4528 14772 4581
rect 15507 4558 15618 4580
rect 15507 4538 15515 4558
rect 15534 4538 15592 4558
rect 15611 4538 15618 4558
rect 16007 4566 16039 4583
rect 16308 4566 16345 4702
rect 16446 4669 16556 4683
rect 16446 4666 16524 4669
rect 16446 4639 16450 4666
rect 16479 4642 16524 4666
rect 16553 4642 16556 4669
rect 17176 4659 17210 4702
rect 16479 4639 16556 4642
rect 16446 4624 16556 4639
rect 17175 4654 17210 4659
rect 17175 4634 17182 4654
rect 17202 4634 17210 4654
rect 17175 4626 17210 4634
rect 16007 4553 16345 4566
rect 12841 4303 12875 4509
rect 13288 4489 13320 4517
rect 13778 4502 14774 4528
rect 15507 4521 15618 4538
rect 16008 4534 16345 4553
rect 16287 4533 16345 4534
rect 16731 4561 16763 4568
rect 16731 4541 16738 4561
rect 16759 4541 16763 4561
rect 12908 4481 13320 4489
rect 12908 4455 12914 4481
rect 12940 4455 13320 4481
rect 12908 4453 13320 4455
rect 12910 4452 12950 4453
rect 13070 4417 13109 4432
rect 13070 4376 13081 4417
rect 13102 4376 13109 4417
rect 12840 4295 12876 4303
rect 12840 4275 12849 4295
rect 12869 4275 12876 4295
rect 12840 4274 12876 4275
rect 12840 4263 12874 4274
rect 13070 4103 13109 4376
rect 13288 4388 13320 4453
rect 16731 4476 16763 4541
rect 17101 4476 17141 4477
rect 16731 4474 17143 4476
rect 16731 4448 17111 4474
rect 17137 4448 17143 4474
rect 16731 4440 17143 4448
rect 13288 4368 13292 4388
rect 13313 4368 13320 4388
rect 13288 4361 13320 4368
rect 13706 4395 13764 4396
rect 13706 4376 14043 4395
rect 14433 4391 14544 4408
rect 15277 4401 16273 4427
rect 16731 4412 16763 4440
rect 13706 4363 14044 4376
rect 13210 4299 13263 4302
rect 13210 4282 13222 4299
rect 13254 4282 13263 4299
rect 13210 4274 13263 4282
rect 13209 4227 13263 4274
rect 13495 4290 13605 4305
rect 13495 4287 13572 4290
rect 13495 4260 13498 4287
rect 13527 4263 13572 4287
rect 13601 4263 13605 4290
rect 13527 4260 13605 4263
rect 13495 4246 13605 4260
rect 13706 4227 13743 4363
rect 14012 4346 14044 4363
rect 14433 4371 14440 4391
rect 14459 4371 14517 4391
rect 14536 4371 14544 4391
rect 14433 4349 14544 4371
rect 15279 4348 15321 4401
rect 14012 4300 14043 4346
rect 15279 4329 15288 4348
rect 15313 4329 15321 4348
rect 15279 4319 15321 4329
rect 15507 4359 15617 4373
rect 15507 4356 15585 4359
rect 15507 4329 15511 4356
rect 15540 4332 15585 4356
rect 15614 4332 15617 4359
rect 16237 4349 16271 4401
rect 16731 4392 16736 4412
rect 16757 4392 16763 4412
rect 16731 4385 16763 4392
rect 16941 4413 16979 4423
rect 17176 4420 17210 4626
rect 16941 4396 16951 4413
rect 16971 4396 16979 4413
rect 16782 4353 16823 4354
rect 15540 4329 15617 4332
rect 15507 4314 15617 4329
rect 16236 4344 16271 4349
rect 16236 4324 16243 4344
rect 16263 4324 16271 4344
rect 16781 4343 16823 4353
rect 16236 4316 16271 4324
rect 13800 4297 13835 4298
rect 13779 4290 13835 4297
rect 13779 4270 13808 4290
rect 13828 4270 13835 4290
rect 13779 4265 13835 4270
rect 14012 4293 14051 4300
rect 14012 4273 14018 4293
rect 14043 4273 14051 4293
rect 14012 4267 14051 4273
rect 14226 4293 14258 4300
rect 14226 4273 14232 4293
rect 14253 4273 14258 4293
rect 13209 4192 13744 4227
rect 13209 4188 13262 4192
rect 13070 4076 13074 4103
rect 13105 4076 13109 4103
rect 13355 4124 13466 4141
rect 13355 4104 13362 4124
rect 13381 4104 13439 4124
rect 13458 4104 13466 4124
rect 13355 4082 13466 4104
rect 13070 4069 13109 4076
rect 13779 4059 13813 4265
rect 14226 4245 14258 4273
rect 13846 4237 14258 4245
rect 13846 4211 13852 4237
rect 13878 4211 14258 4237
rect 13846 4209 14258 4211
rect 13848 4208 13888 4209
rect 14226 4144 14258 4209
rect 15792 4251 15824 4258
rect 15792 4231 15799 4251
rect 15820 4231 15824 4251
rect 15792 4166 15824 4231
rect 16162 4166 16202 4167
rect 15792 4164 16204 4166
rect 14226 4124 14230 4144
rect 14251 4124 14258 4144
rect 14226 4117 14258 4124
rect 14729 4159 14777 4164
rect 14729 4130 14740 4159
rect 14769 4130 14777 4159
rect 13779 4058 13814 4059
rect 13777 4051 13814 4058
rect 12722 4030 12757 4031
rect 12699 4023 12757 4030
rect 12699 4003 12730 4023
rect 12750 4003 12757 4023
rect 12699 3998 12757 4003
rect 13148 4026 13180 4033
rect 13148 4006 13154 4026
rect 13175 4006 13180 4026
rect 12699 3850 12735 3998
rect 13148 3978 13180 4006
rect 12768 3970 13180 3978
rect 12768 3944 12774 3970
rect 12800 3944 13180 3970
rect 13777 4031 13787 4051
rect 13807 4031 13814 4051
rect 13777 4026 13814 4031
rect 14433 4046 14543 4061
rect 14433 4043 14510 4046
rect 13777 3975 13812 4026
rect 14433 4016 14436 4043
rect 14465 4019 14510 4043
rect 14539 4019 14543 4046
rect 14465 4016 14543 4019
rect 14433 4002 14543 4016
rect 14729 3975 14777 4130
rect 15792 4138 16172 4164
rect 16198 4138 16204 4164
rect 15792 4130 16204 4138
rect 15792 4102 15824 4130
rect 16237 4110 16271 4316
rect 16445 4314 16556 4336
rect 16445 4294 16453 4314
rect 16472 4294 16530 4314
rect 16549 4294 16556 4314
rect 16445 4277 16556 4294
rect 16781 4321 16788 4343
rect 16814 4321 16823 4343
rect 16781 4312 16823 4321
rect 15998 4107 16041 4109
rect 15792 4082 15797 4102
rect 15818 4082 15824 4102
rect 15792 4075 15824 4082
rect 15997 4100 16041 4107
rect 15997 4080 16007 4100
rect 16030 4080 16041 4100
rect 15997 4076 16041 4080
rect 16215 4105 16271 4110
rect 16215 4085 16222 4105
rect 16242 4085 16271 4105
rect 16215 4078 16271 4085
rect 16327 4246 16360 4247
rect 16781 4246 16818 4312
rect 16327 4217 16818 4246
rect 16215 4077 16250 4078
rect 13777 3951 14777 3975
rect 15506 4004 15617 4026
rect 15506 3984 15514 4004
rect 15533 3984 15591 4004
rect 15610 3984 15617 4004
rect 15506 3967 15617 3984
rect 15997 3995 16039 4076
rect 16327 3997 16360 4217
rect 16781 4215 16818 4217
rect 16587 4077 16697 4091
rect 16587 4074 16665 4077
rect 16587 4047 16591 4074
rect 16620 4050 16665 4074
rect 16694 4050 16697 4077
rect 16620 4047 16697 4050
rect 16587 4032 16697 4047
rect 16941 4058 16979 4396
rect 17154 4415 17210 4420
rect 17154 4395 17161 4415
rect 17181 4395 17210 4415
rect 17154 4388 17210 4395
rect 17419 4687 17426 4727
rect 17453 4687 17466 4727
rect 17649 4705 17696 4883
rect 18442 4874 18445 4901
rect 18474 4877 18519 4901
rect 18548 4877 18552 4904
rect 18474 4874 18552 4877
rect 18442 4860 18552 4874
rect 17154 4387 17189 4388
rect 17319 4067 17351 4068
rect 16941 4041 16949 4058
rect 16969 4041 16979 4058
rect 16941 4035 16979 4041
rect 17316 4062 17351 4067
rect 17316 4042 17323 4062
rect 17343 4042 17351 4062
rect 17316 4034 17351 4042
rect 16299 3995 16360 3997
rect 15997 3966 16360 3995
rect 16872 3969 16904 3976
rect 15997 3964 16299 3966
rect 13777 3948 14776 3951
rect 16872 3949 16879 3969
rect 16900 3949 16904 3969
rect 13777 3946 13812 3948
rect 12768 3942 13180 3944
rect 12770 3941 12810 3942
rect 12702 3792 12735 3850
rect 12932 3902 12970 3912
rect 12932 3864 12941 3902
rect 12964 3864 12970 3902
rect 12702 3784 12736 3792
rect 12702 3764 12709 3784
rect 12729 3764 12736 3784
rect 12702 3759 12736 3764
rect 12702 3758 12733 3759
rect 12932 3728 12970 3864
rect 13148 3877 13180 3942
rect 16872 3884 16904 3949
rect 17242 3884 17282 3885
rect 16872 3882 17284 3884
rect 16240 3878 16275 3880
rect 13148 3857 13152 3877
rect 13173 3857 13180 3877
rect 15276 3875 16275 3878
rect 13753 3860 14055 3862
rect 13148 3850 13180 3857
rect 13692 3831 14055 3860
rect 13692 3829 13753 3831
rect 13073 3785 13111 3791
rect 13073 3768 13083 3785
rect 13103 3768 13111 3785
rect 12932 3574 12976 3728
rect 12769 3572 12976 3574
rect 12745 3539 12976 3572
rect 11842 2913 11846 2933
rect 11867 2913 11876 2933
rect 11842 2907 11876 2913
rect 11995 3044 12324 3047
rect 12363 3044 12407 3069
rect 11995 3014 12407 3044
rect 11244 2851 11305 2853
rect 10942 2822 11305 2851
rect 11786 2838 11818 2845
rect 10942 2820 11244 2822
rect 8204 2777 8208 2797
rect 8229 2777 8236 2797
rect 11786 2818 11793 2838
rect 11814 2818 11818 2838
rect 8778 2793 9080 2795
rect 8204 2770 8236 2777
rect 8717 2764 9080 2793
rect 8717 2762 8778 2764
rect 7757 2711 7792 2712
rect 7234 2701 7290 2708
rect 7755 2704 7793 2711
rect 7234 2700 7269 2701
rect 5511 2672 5588 2675
rect 5478 2657 5588 2672
rect 6207 2687 6244 2692
rect 6207 2667 6214 2687
rect 6234 2667 6244 2687
rect 7755 2684 7765 2704
rect 7785 2684 7793 2704
rect 6207 2660 6244 2667
rect 7229 2662 7299 2672
rect 6207 2659 6242 2660
rect 5244 2559 5252 2588
rect 5281 2559 5292 2588
rect 5244 2554 5292 2559
rect 5763 2594 5795 2601
rect 5763 2574 5770 2594
rect 5791 2574 5795 2594
rect 3817 2552 4229 2554
rect 3819 2551 3859 2552
rect 4197 2487 4229 2552
rect 4197 2467 4201 2487
rect 4222 2467 4229 2487
rect 4197 2460 4229 2467
rect 5763 2509 5795 2574
rect 6133 2509 6173 2510
rect 5763 2507 6175 2509
rect 5763 2481 6143 2507
rect 6169 2481 6175 2507
rect 5763 2473 6175 2481
rect 5763 2445 5795 2473
rect 6208 2453 6242 2659
rect 7227 2655 7299 2662
rect 6525 2627 6636 2649
rect 6525 2607 6533 2627
rect 6552 2607 6610 2627
rect 6629 2607 6636 2627
rect 6525 2590 6636 2607
rect 7227 2626 7234 2655
rect 7282 2626 7299 2655
rect 7227 2617 7299 2626
rect 7146 2526 7180 2527
rect 6277 2491 7181 2526
rect 5763 2425 5768 2445
rect 5789 2425 5795 2445
rect 5763 2418 5795 2425
rect 5970 2445 6009 2451
rect 5970 2425 5978 2445
rect 6003 2425 6009 2445
rect 5970 2418 6009 2425
rect 6186 2448 6242 2453
rect 6186 2428 6193 2448
rect 6213 2428 6242 2448
rect 6186 2421 6242 2428
rect 6186 2420 6221 2421
rect 3750 2394 3785 2402
rect 3198 2365 3240 2375
rect 3750 2374 3758 2394
rect 3778 2374 3785 2394
rect 3750 2369 3785 2374
rect 4404 2389 4514 2404
rect 4404 2386 4481 2389
rect 3198 2364 3239 2365
rect 2832 2330 2867 2331
rect 2811 2323 2867 2330
rect 2811 2303 2840 2323
rect 2860 2303 2867 2323
rect 2811 2298 2867 2303
rect 3258 2326 3290 2333
rect 3258 2306 3264 2326
rect 3285 2306 3290 2326
rect 3750 2317 3784 2369
rect 4404 2359 4407 2386
rect 4436 2362 4481 2386
rect 4510 2362 4514 2389
rect 4436 2359 4514 2362
rect 4404 2345 4514 2359
rect 4700 2389 4742 2399
rect 4700 2370 4708 2389
rect 4733 2370 4742 2389
rect 5978 2372 6009 2418
rect 4700 2317 4742 2370
rect 5477 2347 5588 2369
rect 5477 2327 5485 2347
rect 5504 2327 5562 2347
rect 5581 2327 5588 2347
rect 5977 2355 6009 2372
rect 6278 2355 6315 2491
rect 6416 2458 6526 2472
rect 6416 2455 6494 2458
rect 6416 2428 6420 2455
rect 6449 2431 6494 2455
rect 6523 2431 6526 2458
rect 7146 2448 7180 2491
rect 6449 2428 6526 2431
rect 6416 2413 6526 2428
rect 7145 2443 7180 2448
rect 7145 2423 7152 2443
rect 7172 2423 7180 2443
rect 7145 2415 7180 2423
rect 5977 2342 6315 2355
rect 2811 2092 2845 2298
rect 3258 2278 3290 2306
rect 3748 2291 4744 2317
rect 5477 2310 5588 2327
rect 5978 2323 6315 2342
rect 6257 2322 6315 2323
rect 6701 2350 6733 2357
rect 6701 2330 6708 2350
rect 6729 2330 6733 2350
rect 2878 2270 3290 2278
rect 2878 2244 2884 2270
rect 2910 2244 3290 2270
rect 2878 2242 3290 2244
rect 2880 2241 2920 2242
rect 3040 2206 3079 2221
rect 3040 2165 3051 2206
rect 3072 2165 3079 2206
rect 2810 2084 2846 2092
rect 2810 2064 2819 2084
rect 2839 2064 2846 2084
rect 2810 2063 2846 2064
rect 2810 2052 2844 2063
rect 2700 2022 2737 2030
rect 1990 2000 2197 2002
rect 1990 1846 2034 2000
rect 2700 1988 2944 2022
rect 1855 1789 1863 1806
rect 1883 1789 1893 1806
rect 1855 1783 1893 1789
rect 1213 1743 1274 1745
rect 911 1714 1274 1743
rect 1786 1717 1818 1724
rect 911 1712 1213 1714
rect 1786 1697 1793 1717
rect 1814 1697 1818 1717
rect 1786 1632 1818 1697
rect 1996 1710 2034 1846
rect 2692 1819 2727 1820
rect 2233 1815 2264 1816
rect 2230 1810 2264 1815
rect 2230 1790 2237 1810
rect 2257 1790 2264 1810
rect 2230 1782 2264 1790
rect 1996 1672 2002 1710
rect 2025 1672 2034 1710
rect 1996 1662 2034 1672
rect 2231 1724 2264 1782
rect 2671 1812 2727 1819
rect 2671 1792 2700 1812
rect 2720 1792 2727 1812
rect 2671 1787 2727 1792
rect 2902 1817 2944 1988
rect 3040 1892 3079 2165
rect 3258 2177 3290 2242
rect 6701 2265 6733 2330
rect 7071 2265 7111 2266
rect 6701 2263 7113 2265
rect 6701 2237 7081 2263
rect 7107 2237 7113 2263
rect 6701 2229 7113 2237
rect 3258 2157 3262 2177
rect 3283 2157 3290 2177
rect 3258 2150 3290 2157
rect 3676 2184 3734 2185
rect 3676 2165 4013 2184
rect 4403 2180 4514 2197
rect 5247 2190 6243 2216
rect 6701 2201 6733 2229
rect 3676 2152 4014 2165
rect 3180 2088 3233 2091
rect 3180 2071 3192 2088
rect 3224 2071 3233 2088
rect 3180 2063 3233 2071
rect 3179 2016 3233 2063
rect 3465 2079 3575 2094
rect 3465 2076 3542 2079
rect 3465 2049 3468 2076
rect 3497 2052 3542 2076
rect 3571 2052 3575 2079
rect 3497 2049 3575 2052
rect 3465 2035 3575 2049
rect 3676 2016 3713 2152
rect 3982 2135 4014 2152
rect 4403 2160 4410 2180
rect 4429 2160 4487 2180
rect 4506 2160 4514 2180
rect 4403 2138 4514 2160
rect 5249 2137 5291 2190
rect 3982 2089 4013 2135
rect 5249 2118 5258 2137
rect 5283 2118 5291 2137
rect 5249 2108 5291 2118
rect 5477 2148 5587 2162
rect 5477 2145 5555 2148
rect 5477 2118 5481 2145
rect 5510 2121 5555 2145
rect 5584 2121 5587 2148
rect 6207 2138 6241 2190
rect 6701 2181 6706 2201
rect 6727 2181 6733 2201
rect 6701 2174 6733 2181
rect 6911 2202 6949 2212
rect 7146 2209 7180 2415
rect 6911 2185 6921 2202
rect 6941 2185 6949 2202
rect 6752 2142 6793 2143
rect 5510 2118 5587 2121
rect 5477 2103 5587 2118
rect 6206 2133 6241 2138
rect 6206 2113 6213 2133
rect 6233 2113 6241 2133
rect 6751 2132 6793 2142
rect 6206 2105 6241 2113
rect 3770 2086 3805 2087
rect 3749 2079 3805 2086
rect 3749 2059 3778 2079
rect 3798 2059 3805 2079
rect 3749 2054 3805 2059
rect 3982 2082 4021 2089
rect 3982 2062 3988 2082
rect 4013 2062 4021 2082
rect 3982 2056 4021 2062
rect 4196 2082 4228 2089
rect 4196 2062 4202 2082
rect 4223 2062 4228 2082
rect 3179 1981 3714 2016
rect 3179 1977 3232 1981
rect 3040 1865 3044 1892
rect 3075 1865 3079 1892
rect 3325 1913 3436 1930
rect 3325 1893 3332 1913
rect 3351 1893 3409 1913
rect 3428 1893 3436 1913
rect 3325 1871 3436 1893
rect 3040 1858 3079 1865
rect 3749 1848 3783 2054
rect 4196 2034 4228 2062
rect 3816 2026 4228 2034
rect 3816 2000 3822 2026
rect 3848 2000 4228 2026
rect 3816 1998 4228 2000
rect 3818 1997 3858 1998
rect 4196 1933 4228 1998
rect 5762 2040 5794 2047
rect 5762 2020 5769 2040
rect 5790 2020 5794 2040
rect 5762 1955 5794 2020
rect 6132 1955 6172 1956
rect 5762 1953 6174 1955
rect 4196 1913 4200 1933
rect 4221 1913 4228 1933
rect 4196 1906 4228 1913
rect 4699 1948 4747 1953
rect 4699 1919 4710 1948
rect 4739 1919 4747 1948
rect 3749 1847 3784 1848
rect 3747 1840 3784 1847
rect 2902 1796 2910 1817
rect 2937 1796 2944 1817
rect 2156 1632 2196 1633
rect 1786 1630 2198 1632
rect 1154 1626 1189 1628
rect 190 1623 1189 1626
rect 189 1599 1189 1623
rect 189 1444 237 1599
rect 423 1558 533 1572
rect 423 1555 501 1558
rect 423 1528 427 1555
rect 456 1531 501 1555
rect 530 1531 533 1558
rect 1154 1548 1189 1599
rect 456 1528 533 1531
rect 423 1513 533 1528
rect 1152 1543 1189 1548
rect 1152 1523 1159 1543
rect 1179 1523 1189 1543
rect 1786 1604 2166 1630
rect 2192 1604 2198 1630
rect 1786 1596 2198 1604
rect 1786 1568 1818 1596
rect 2231 1576 2267 1724
rect 1786 1548 1791 1568
rect 1812 1548 1818 1568
rect 1786 1541 1818 1548
rect 2209 1571 2267 1576
rect 2209 1551 2216 1571
rect 2236 1551 2267 1571
rect 2209 1544 2267 1551
rect 2671 1581 2705 1787
rect 2902 1785 2944 1796
rect 3118 1815 3150 1822
rect 3118 1795 3124 1815
rect 3145 1795 3150 1815
rect 3118 1767 3150 1795
rect 2738 1759 3150 1767
rect 2738 1733 2744 1759
rect 2770 1733 3150 1759
rect 3747 1820 3757 1840
rect 3777 1820 3784 1840
rect 3747 1815 3784 1820
rect 4403 1835 4513 1850
rect 4403 1832 4480 1835
rect 3747 1764 3782 1815
rect 4403 1805 4406 1832
rect 4435 1808 4480 1832
rect 4509 1808 4513 1835
rect 4435 1805 4513 1808
rect 4403 1791 4513 1805
rect 4699 1764 4747 1919
rect 5762 1927 6142 1953
rect 6168 1927 6174 1953
rect 5762 1919 6174 1927
rect 5762 1891 5794 1919
rect 6207 1899 6241 2105
rect 6415 2103 6526 2125
rect 6415 2083 6423 2103
rect 6442 2083 6500 2103
rect 6519 2083 6526 2103
rect 6415 2066 6526 2083
rect 6751 2110 6758 2132
rect 6784 2110 6793 2132
rect 6751 2101 6793 2110
rect 5968 1896 6011 1898
rect 5762 1871 5767 1891
rect 5788 1871 5794 1891
rect 5762 1864 5794 1871
rect 5967 1889 6011 1896
rect 5967 1869 5977 1889
rect 6000 1869 6011 1889
rect 5967 1865 6011 1869
rect 6185 1894 6241 1899
rect 6185 1874 6192 1894
rect 6212 1874 6241 1894
rect 6185 1867 6241 1874
rect 6297 2035 6330 2036
rect 6751 2035 6788 2101
rect 6297 2006 6788 2035
rect 6185 1866 6220 1867
rect 3747 1740 4747 1764
rect 5476 1793 5587 1815
rect 5476 1773 5484 1793
rect 5503 1773 5561 1793
rect 5580 1773 5587 1793
rect 5476 1756 5587 1773
rect 5967 1784 6009 1865
rect 6297 1786 6330 2006
rect 6751 2004 6788 2006
rect 6557 1866 6667 1880
rect 6557 1863 6635 1866
rect 6557 1836 6561 1863
rect 6590 1839 6635 1863
rect 6664 1839 6667 1866
rect 6590 1836 6667 1839
rect 6557 1821 6667 1836
rect 6911 1847 6949 2185
rect 7124 2204 7180 2209
rect 7124 2184 7131 2204
rect 7151 2184 7180 2204
rect 7124 2177 7180 2184
rect 7124 2176 7159 2177
rect 7046 2076 7090 2080
rect 7227 2076 7277 2617
rect 7046 2043 7277 2076
rect 7755 2071 7793 2684
rect 8411 2699 8521 2714
rect 8411 2696 8488 2699
rect 8411 2669 8414 2696
rect 8443 2672 8488 2696
rect 8517 2672 8521 2699
rect 8443 2669 8521 2672
rect 8411 2655 8521 2669
rect 8259 2542 8296 2544
rect 8717 2542 8750 2762
rect 9038 2683 9080 2764
rect 9460 2775 9571 2791
rect 9460 2755 9467 2775
rect 9486 2755 9544 2775
rect 9563 2755 9571 2775
rect 9460 2733 9571 2755
rect 11786 2753 11818 2818
rect 11995 2826 12030 3014
rect 12297 3012 12407 3014
rect 12590 3027 12640 3155
rect 12745 3138 12795 3539
rect 12932 3535 12976 3539
rect 12863 3438 12898 3439
rect 12725 3129 12795 3138
rect 12725 3100 12740 3129
rect 12788 3121 12795 3129
rect 12842 3431 12898 3438
rect 12842 3411 12871 3431
rect 12891 3411 12898 3431
rect 12842 3406 12898 3411
rect 13073 3430 13111 3768
rect 13355 3779 13465 3794
rect 13355 3776 13432 3779
rect 13355 3749 13358 3776
rect 13387 3752 13432 3776
rect 13461 3752 13465 3779
rect 13387 3749 13465 3752
rect 13355 3735 13465 3749
rect 13234 3609 13271 3611
rect 13692 3609 13725 3829
rect 14013 3750 14055 3831
rect 14435 3842 14546 3859
rect 14435 3822 14442 3842
rect 14461 3822 14519 3842
rect 14538 3822 14546 3842
rect 14435 3800 14546 3822
rect 15275 3851 16275 3875
rect 13802 3748 13837 3749
rect 13234 3580 13725 3609
rect 13234 3514 13271 3580
rect 13692 3579 13725 3580
rect 13781 3741 13837 3748
rect 13781 3721 13810 3741
rect 13830 3721 13837 3741
rect 13781 3716 13837 3721
rect 14011 3746 14055 3750
rect 14011 3726 14022 3746
rect 14045 3726 14055 3746
rect 14011 3719 14055 3726
rect 14228 3744 14260 3751
rect 14228 3724 14234 3744
rect 14255 3724 14260 3744
rect 14011 3717 14054 3719
rect 13229 3505 13271 3514
rect 13229 3483 13238 3505
rect 13264 3483 13271 3505
rect 13496 3532 13607 3549
rect 13496 3512 13503 3532
rect 13522 3512 13580 3532
rect 13599 3512 13607 3532
rect 13496 3490 13607 3512
rect 13781 3510 13815 3716
rect 14228 3696 14260 3724
rect 13848 3688 14260 3696
rect 13848 3662 13854 3688
rect 13880 3662 14260 3688
rect 15275 3696 15323 3851
rect 15509 3810 15619 3824
rect 15509 3807 15587 3810
rect 15509 3780 15513 3807
rect 15542 3783 15587 3807
rect 15616 3783 15619 3810
rect 16240 3800 16275 3851
rect 15542 3780 15619 3783
rect 15509 3765 15619 3780
rect 16238 3795 16275 3800
rect 16238 3775 16245 3795
rect 16265 3775 16275 3795
rect 16872 3856 17252 3882
rect 17278 3856 17284 3882
rect 16872 3848 17284 3856
rect 16872 3820 16904 3848
rect 16872 3800 16877 3820
rect 16898 3800 16904 3820
rect 16872 3793 16904 3800
rect 17078 3819 17120 3830
rect 17317 3828 17351 4034
rect 17078 3798 17085 3819
rect 17112 3798 17120 3819
rect 16238 3768 16275 3775
rect 16238 3767 16273 3768
rect 15275 3667 15283 3696
rect 15312 3667 15323 3696
rect 15275 3662 15323 3667
rect 15794 3702 15826 3709
rect 15794 3682 15801 3702
rect 15822 3682 15826 3702
rect 13848 3660 14260 3662
rect 13850 3659 13890 3660
rect 14228 3595 14260 3660
rect 14228 3575 14232 3595
rect 14253 3575 14260 3595
rect 14228 3568 14260 3575
rect 15794 3617 15826 3682
rect 16164 3617 16204 3618
rect 15794 3615 16206 3617
rect 15794 3589 16174 3615
rect 16200 3589 16206 3615
rect 15794 3581 16206 3589
rect 15794 3553 15826 3581
rect 16239 3561 16273 3767
rect 16943 3750 16982 3757
rect 16586 3722 16697 3744
rect 16586 3702 16594 3722
rect 16613 3702 16671 3722
rect 16690 3702 16697 3722
rect 16586 3685 16697 3702
rect 16943 3723 16947 3750
rect 16978 3723 16982 3750
rect 16790 3634 16843 3638
rect 16308 3599 16843 3634
rect 15794 3533 15799 3553
rect 15820 3533 15826 3553
rect 15794 3526 15826 3533
rect 16001 3553 16040 3559
rect 16001 3533 16009 3553
rect 16034 3533 16040 3553
rect 16001 3526 16040 3533
rect 16217 3556 16273 3561
rect 16217 3536 16224 3556
rect 16244 3536 16273 3556
rect 16217 3529 16273 3536
rect 16217 3528 16252 3529
rect 13781 3502 13816 3510
rect 13229 3473 13271 3483
rect 13781 3482 13789 3502
rect 13809 3482 13816 3502
rect 13781 3477 13816 3482
rect 14435 3497 14545 3512
rect 14435 3494 14512 3497
rect 13229 3472 13270 3473
rect 13073 3413 13081 3430
rect 13101 3413 13111 3430
rect 12842 3200 12876 3406
rect 13073 3403 13111 3413
rect 13289 3434 13321 3441
rect 13289 3414 13295 3434
rect 13316 3414 13321 3434
rect 13781 3425 13815 3477
rect 14435 3467 14438 3494
rect 14467 3470 14512 3494
rect 14541 3470 14545 3497
rect 14467 3467 14545 3470
rect 14435 3453 14545 3467
rect 14731 3497 14773 3507
rect 14731 3478 14739 3497
rect 14764 3478 14773 3497
rect 16009 3480 16040 3526
rect 14731 3425 14773 3478
rect 15508 3455 15619 3477
rect 15508 3435 15516 3455
rect 15535 3435 15593 3455
rect 15612 3435 15619 3455
rect 16008 3463 16040 3480
rect 16309 3463 16346 3599
rect 16447 3566 16557 3580
rect 16447 3563 16525 3566
rect 16447 3536 16451 3563
rect 16480 3539 16525 3563
rect 16554 3539 16557 3566
rect 16480 3536 16557 3539
rect 16447 3521 16557 3536
rect 16789 3552 16843 3599
rect 16789 3544 16842 3552
rect 16789 3527 16798 3544
rect 16830 3527 16842 3544
rect 16789 3524 16842 3527
rect 16008 3450 16346 3463
rect 13289 3386 13321 3414
rect 13779 3399 14775 3425
rect 15508 3418 15619 3435
rect 16009 3431 16346 3450
rect 16288 3430 16346 3431
rect 16732 3458 16764 3465
rect 16732 3438 16739 3458
rect 16760 3438 16764 3458
rect 12909 3378 13321 3386
rect 12909 3352 12915 3378
rect 12941 3352 13321 3378
rect 12909 3350 13321 3352
rect 12911 3349 12951 3350
rect 13289 3285 13321 3350
rect 16732 3373 16764 3438
rect 16943 3450 16982 3723
rect 17078 3627 17120 3798
rect 17295 3823 17351 3828
rect 17295 3803 17302 3823
rect 17322 3803 17351 3823
rect 17295 3796 17351 3803
rect 17295 3795 17330 3796
rect 17078 3593 17322 3627
rect 17285 3585 17322 3593
rect 17178 3552 17212 3563
rect 17176 3551 17212 3552
rect 17176 3531 17183 3551
rect 17203 3531 17212 3551
rect 17176 3523 17212 3531
rect 16943 3409 16950 3450
rect 16971 3409 16982 3450
rect 16943 3394 16982 3409
rect 17102 3373 17142 3374
rect 16732 3371 17144 3373
rect 16732 3345 17112 3371
rect 17138 3345 17144 3371
rect 16732 3337 17144 3345
rect 13289 3265 13293 3285
rect 13314 3265 13321 3285
rect 13289 3258 13321 3265
rect 13707 3292 13765 3293
rect 13707 3273 14044 3292
rect 14434 3288 14545 3305
rect 15278 3298 16274 3324
rect 16732 3309 16764 3337
rect 17177 3317 17211 3523
rect 13707 3260 14045 3273
rect 12842 3192 12877 3200
rect 12842 3172 12850 3192
rect 12870 3172 12877 3192
rect 12842 3167 12877 3172
rect 13496 3187 13606 3202
rect 13496 3184 13573 3187
rect 12842 3124 12876 3167
rect 13496 3157 13499 3184
rect 13528 3160 13573 3184
rect 13602 3160 13606 3187
rect 13528 3157 13606 3160
rect 13496 3143 13606 3157
rect 13707 3124 13744 3260
rect 14013 3243 14045 3260
rect 14434 3268 14441 3288
rect 14460 3268 14518 3288
rect 14537 3268 14545 3288
rect 14434 3246 14545 3268
rect 15280 3245 15322 3298
rect 14013 3197 14044 3243
rect 15280 3226 15289 3245
rect 15314 3226 15322 3245
rect 15280 3216 15322 3226
rect 15508 3256 15618 3270
rect 15508 3253 15586 3256
rect 15508 3226 15512 3253
rect 15541 3229 15586 3253
rect 15615 3229 15618 3256
rect 16238 3246 16272 3298
rect 16732 3289 16737 3309
rect 16758 3289 16764 3309
rect 16732 3282 16764 3289
rect 17155 3312 17211 3317
rect 17155 3292 17162 3312
rect 17182 3292 17211 3312
rect 17155 3285 17211 3292
rect 17155 3284 17190 3285
rect 16783 3250 16824 3251
rect 15541 3226 15618 3229
rect 15508 3211 15618 3226
rect 16237 3241 16272 3246
rect 16237 3221 16244 3241
rect 16264 3221 16272 3241
rect 16782 3240 16824 3250
rect 16237 3213 16272 3221
rect 13801 3194 13836 3195
rect 13780 3187 13836 3194
rect 13780 3167 13809 3187
rect 13829 3167 13836 3187
rect 13780 3162 13836 3167
rect 14013 3190 14052 3197
rect 14013 3170 14019 3190
rect 14044 3170 14052 3190
rect 14013 3164 14052 3170
rect 14227 3190 14259 3197
rect 14227 3170 14233 3190
rect 14254 3170 14259 3190
rect 12788 3100 12793 3121
rect 12725 3089 12793 3100
rect 12841 3089 13745 3124
rect 12842 3088 12876 3089
rect 12590 2993 13005 3027
rect 12590 2991 12640 2993
rect 12223 2929 12273 2936
rect 12223 2915 12237 2929
rect 12229 2911 12237 2915
rect 12257 2915 12273 2929
rect 12257 2911 12267 2915
rect 12753 2914 12788 2915
rect 12229 2904 12267 2911
rect 12732 2907 12788 2914
rect 12230 2903 12265 2904
rect 11995 2794 12000 2826
rect 12027 2794 12030 2826
rect 11995 2776 12030 2794
rect 12156 2753 12196 2754
rect 11786 2751 12198 2753
rect 11184 2734 11219 2736
rect 10220 2731 11219 2734
rect 10219 2707 11219 2731
rect 8827 2681 8862 2682
rect 8259 2513 8750 2542
rect 8259 2447 8296 2513
rect 8717 2512 8750 2513
rect 8806 2674 8862 2681
rect 8806 2654 8835 2674
rect 8855 2654 8862 2674
rect 8806 2649 8862 2654
rect 9036 2679 9080 2683
rect 9036 2659 9047 2679
rect 9070 2659 9080 2679
rect 9036 2652 9080 2659
rect 9253 2677 9285 2684
rect 9253 2657 9259 2677
rect 9280 2657 9285 2677
rect 9036 2650 9079 2652
rect 8254 2438 8296 2447
rect 8254 2416 8263 2438
rect 8289 2416 8296 2438
rect 8521 2465 8632 2482
rect 8521 2445 8528 2465
rect 8547 2445 8605 2465
rect 8624 2445 8632 2465
rect 8521 2423 8632 2445
rect 8806 2443 8840 2649
rect 9253 2629 9285 2657
rect 8873 2621 9285 2629
rect 8873 2595 8879 2621
rect 8905 2595 9285 2621
rect 8873 2593 9285 2595
rect 8875 2592 8915 2593
rect 9253 2528 9285 2593
rect 9253 2508 9257 2528
rect 9278 2508 9285 2528
rect 10219 2552 10267 2707
rect 10453 2666 10563 2680
rect 10453 2663 10531 2666
rect 10453 2636 10457 2663
rect 10486 2639 10531 2663
rect 10560 2639 10563 2666
rect 11184 2656 11219 2707
rect 11786 2725 12166 2751
rect 12192 2725 12198 2751
rect 11786 2717 12198 2725
rect 11786 2689 11818 2717
rect 12231 2697 12265 2903
rect 11786 2669 11791 2689
rect 11812 2669 11818 2689
rect 11786 2662 11818 2669
rect 12209 2692 12265 2697
rect 12209 2672 12216 2692
rect 12236 2672 12265 2692
rect 12732 2887 12761 2907
rect 12781 2887 12788 2907
rect 12732 2882 12788 2887
rect 12960 2910 13005 2993
rect 13386 3008 13497 3025
rect 13386 2988 13393 3008
rect 13412 2988 13470 3008
rect 13489 2988 13497 3008
rect 13386 2966 13497 2988
rect 13780 2956 13814 3162
rect 14227 3142 14259 3170
rect 13847 3134 14259 3142
rect 13847 3108 13853 3134
rect 13879 3108 14259 3134
rect 13847 3106 14259 3108
rect 13849 3105 13889 3106
rect 14227 3041 14259 3106
rect 15793 3148 15825 3155
rect 15793 3128 15800 3148
rect 15821 3128 15825 3148
rect 15793 3063 15825 3128
rect 16163 3063 16203 3064
rect 15793 3061 16205 3063
rect 14227 3021 14231 3041
rect 14252 3021 14259 3041
rect 14227 3014 14259 3021
rect 14730 3056 14778 3061
rect 14730 3027 14741 3056
rect 14770 3027 14778 3056
rect 13780 2955 13815 2956
rect 13778 2948 13815 2955
rect 13778 2928 13788 2948
rect 13808 2928 13815 2948
rect 13778 2923 13815 2928
rect 14434 2943 14544 2958
rect 14434 2940 14511 2943
rect 12960 2891 12969 2910
rect 12998 2891 13005 2910
rect 12732 2676 12766 2882
rect 12960 2879 13005 2891
rect 13179 2910 13211 2917
rect 13179 2890 13185 2910
rect 13206 2890 13211 2910
rect 13179 2862 13211 2890
rect 12799 2854 13211 2862
rect 12799 2828 12805 2854
rect 12831 2828 13211 2854
rect 13778 2872 13813 2923
rect 14434 2913 14437 2940
rect 14466 2916 14511 2940
rect 14540 2916 14544 2943
rect 14466 2913 14544 2916
rect 14434 2899 14544 2913
rect 14730 2872 14778 3027
rect 15793 3035 16173 3061
rect 16199 3035 16205 3061
rect 15793 3027 16205 3035
rect 15793 2999 15825 3027
rect 16238 3007 16272 3213
rect 16446 3211 16557 3233
rect 16446 3191 16454 3211
rect 16473 3191 16531 3211
rect 16550 3191 16557 3211
rect 16446 3174 16557 3191
rect 16782 3218 16789 3240
rect 16815 3218 16824 3240
rect 16782 3209 16824 3218
rect 15999 3004 16042 3006
rect 15793 2979 15798 2999
rect 15819 2979 15825 2999
rect 15793 2972 15825 2979
rect 15998 2997 16042 3004
rect 15998 2977 16008 2997
rect 16031 2977 16042 2997
rect 15998 2973 16042 2977
rect 16216 3002 16272 3007
rect 16216 2982 16223 3002
rect 16243 2982 16272 3002
rect 16216 2975 16272 2982
rect 16328 3143 16361 3144
rect 16782 3143 16819 3209
rect 17285 3194 17323 3585
rect 16899 3178 17323 3194
rect 16328 3114 16819 3143
rect 16216 2974 16251 2975
rect 13778 2848 14778 2872
rect 15507 2901 15618 2923
rect 15507 2881 15515 2901
rect 15534 2881 15592 2901
rect 15611 2881 15618 2901
rect 15507 2865 15618 2881
rect 15998 2892 16040 2973
rect 16328 2894 16361 3114
rect 16782 3112 16819 3114
rect 16898 3153 17323 3178
rect 16557 2987 16667 3001
rect 16557 2984 16635 2987
rect 16557 2957 16561 2984
rect 16590 2960 16635 2984
rect 16664 2960 16667 2987
rect 16590 2957 16667 2960
rect 16557 2942 16667 2957
rect 16898 2974 16932 3153
rect 17419 3110 17466 4687
rect 17648 4681 17696 4705
rect 18289 4753 18326 4755
rect 18747 4753 18780 4973
rect 19068 4894 19110 4975
rect 19490 4986 19601 5003
rect 19490 4966 19497 4986
rect 19516 4966 19574 4986
rect 19593 4966 19601 4986
rect 19490 4944 19601 4966
rect 18857 4892 18892 4893
rect 18289 4724 18780 4753
rect 17648 3196 17694 4681
rect 18289 4658 18326 4724
rect 18747 4723 18780 4724
rect 18836 4885 18892 4892
rect 18836 4865 18865 4885
rect 18885 4865 18892 4885
rect 18836 4860 18892 4865
rect 19066 4890 19110 4894
rect 19066 4870 19077 4890
rect 19100 4870 19110 4890
rect 19066 4863 19110 4870
rect 19283 4888 19315 4895
rect 19283 4868 19289 4888
rect 19310 4868 19315 4888
rect 19066 4861 19109 4863
rect 18284 4649 18326 4658
rect 18284 4627 18293 4649
rect 18319 4627 18326 4649
rect 18551 4676 18662 4693
rect 18551 4656 18558 4676
rect 18577 4656 18635 4676
rect 18654 4656 18662 4676
rect 18551 4634 18662 4656
rect 18836 4654 18870 4860
rect 19283 4840 19315 4868
rect 18903 4832 19315 4840
rect 18903 4806 18909 4832
rect 18935 4806 19315 4832
rect 18903 4804 19315 4806
rect 18905 4803 18945 4804
rect 19283 4739 19315 4804
rect 19283 4719 19287 4739
rect 19308 4719 19315 4739
rect 19283 4712 19315 4719
rect 18836 4646 18871 4654
rect 18284 4617 18326 4627
rect 18836 4626 18844 4646
rect 18864 4626 18871 4646
rect 18836 4621 18871 4626
rect 19490 4641 19600 4656
rect 19490 4638 19567 4641
rect 18284 4616 18325 4617
rect 17918 4582 17953 4583
rect 17897 4575 17953 4582
rect 17897 4555 17926 4575
rect 17946 4555 17953 4575
rect 17897 4550 17953 4555
rect 18344 4578 18376 4585
rect 18344 4558 18350 4578
rect 18371 4558 18376 4578
rect 18836 4569 18870 4621
rect 19490 4611 19493 4638
rect 19522 4614 19567 4638
rect 19596 4614 19600 4641
rect 19522 4611 19600 4614
rect 19490 4597 19600 4611
rect 19786 4641 19828 4651
rect 19786 4622 19794 4641
rect 19819 4622 19828 4641
rect 19786 4569 19828 4622
rect 17897 4344 17931 4550
rect 18344 4530 18376 4558
rect 18834 4543 19830 4569
rect 17964 4522 18376 4530
rect 17964 4496 17970 4522
rect 17996 4496 18376 4522
rect 17964 4494 18376 4496
rect 17966 4493 18006 4494
rect 18126 4458 18165 4473
rect 18126 4417 18137 4458
rect 18158 4417 18165 4458
rect 17896 4336 17932 4344
rect 17896 4316 17905 4336
rect 17925 4316 17932 4336
rect 17896 4315 17932 4316
rect 17896 4304 17930 4315
rect 18126 4144 18165 4417
rect 18344 4429 18376 4494
rect 18344 4409 18348 4429
rect 18369 4409 18376 4429
rect 18344 4402 18376 4409
rect 18762 4436 18820 4437
rect 18762 4417 19099 4436
rect 19489 4432 19600 4449
rect 18762 4404 19100 4417
rect 18266 4340 18319 4343
rect 18266 4323 18278 4340
rect 18310 4323 18319 4340
rect 18266 4315 18319 4323
rect 18265 4268 18319 4315
rect 18551 4331 18661 4346
rect 18551 4328 18628 4331
rect 18551 4301 18554 4328
rect 18583 4304 18628 4328
rect 18657 4304 18661 4331
rect 18583 4301 18661 4304
rect 18551 4287 18661 4301
rect 18762 4268 18799 4404
rect 19068 4387 19100 4404
rect 19489 4412 19496 4432
rect 19515 4412 19573 4432
rect 19592 4412 19600 4432
rect 19489 4390 19600 4412
rect 19068 4341 19099 4387
rect 18856 4338 18891 4339
rect 18835 4331 18891 4338
rect 18835 4311 18864 4331
rect 18884 4311 18891 4331
rect 18835 4306 18891 4311
rect 19068 4334 19107 4341
rect 19068 4314 19074 4334
rect 19099 4314 19107 4334
rect 19068 4308 19107 4314
rect 19282 4334 19314 4341
rect 19282 4314 19288 4334
rect 19309 4314 19314 4334
rect 18265 4233 18800 4268
rect 18265 4229 18318 4233
rect 18126 4117 18130 4144
rect 18161 4117 18165 4144
rect 18411 4165 18522 4182
rect 18411 4145 18418 4165
rect 18437 4145 18495 4165
rect 18514 4145 18522 4165
rect 18411 4123 18522 4145
rect 18126 4110 18165 4117
rect 18835 4100 18869 4306
rect 19282 4286 19314 4314
rect 18902 4278 19314 4286
rect 18902 4252 18908 4278
rect 18934 4252 19314 4278
rect 18902 4250 19314 4252
rect 18904 4249 18944 4250
rect 19282 4185 19314 4250
rect 19282 4165 19286 4185
rect 19307 4165 19314 4185
rect 19282 4158 19314 4165
rect 19785 4200 19833 4205
rect 19785 4171 19796 4200
rect 19825 4171 19833 4200
rect 18835 4099 18870 4100
rect 18833 4092 18870 4099
rect 17778 4071 17813 4072
rect 17755 4064 17813 4071
rect 17755 4044 17786 4064
rect 17806 4044 17813 4064
rect 17755 4039 17813 4044
rect 18204 4067 18236 4074
rect 18204 4047 18210 4067
rect 18231 4047 18236 4067
rect 17755 3891 17791 4039
rect 18204 4019 18236 4047
rect 17824 4011 18236 4019
rect 17824 3985 17830 4011
rect 17856 3985 18236 4011
rect 18833 4072 18843 4092
rect 18863 4072 18870 4092
rect 18833 4067 18870 4072
rect 19489 4087 19599 4102
rect 19489 4084 19566 4087
rect 18833 4016 18868 4067
rect 19489 4057 19492 4084
rect 19521 4060 19566 4084
rect 19595 4060 19599 4087
rect 19521 4057 19599 4060
rect 19489 4043 19599 4057
rect 19785 4016 19833 4171
rect 18833 3992 19833 4016
rect 18833 3989 19832 3992
rect 18833 3987 18868 3989
rect 17824 3983 18236 3985
rect 17826 3982 17866 3983
rect 17758 3833 17791 3891
rect 17988 3943 18026 3953
rect 17988 3905 17997 3943
rect 18020 3905 18026 3943
rect 17758 3825 17792 3833
rect 17758 3805 17765 3825
rect 17785 3805 17792 3825
rect 17758 3800 17792 3805
rect 17758 3799 17789 3800
rect 17988 3769 18026 3905
rect 18204 3918 18236 3983
rect 18204 3898 18208 3918
rect 18229 3898 18236 3918
rect 18809 3901 19111 3903
rect 18204 3891 18236 3898
rect 18748 3872 19111 3901
rect 18748 3870 18809 3872
rect 18129 3826 18167 3832
rect 18129 3809 18139 3826
rect 18159 3809 18167 3826
rect 17988 3615 18032 3769
rect 17825 3613 18032 3615
rect 17801 3580 18032 3613
rect 16898 2954 16902 2974
rect 16923 2954 16932 2974
rect 16898 2948 16932 2954
rect 17051 3085 17380 3088
rect 17419 3085 17463 3110
rect 17051 3055 17463 3085
rect 16300 2892 16361 2894
rect 15998 2863 16361 2892
rect 16842 2879 16874 2886
rect 15998 2861 16300 2863
rect 16842 2859 16849 2879
rect 16870 2859 16874 2879
rect 13778 2845 14777 2848
rect 13778 2843 13813 2845
rect 12799 2826 13211 2828
rect 12801 2825 12841 2826
rect 13179 2761 13211 2826
rect 16842 2794 16874 2859
rect 17051 2867 17086 3055
rect 17353 3053 17463 3055
rect 17646 3068 17696 3196
rect 17801 3179 17851 3580
rect 17988 3576 18032 3580
rect 17919 3479 17954 3480
rect 17781 3170 17851 3179
rect 17781 3141 17796 3170
rect 17844 3162 17851 3170
rect 17898 3472 17954 3479
rect 17898 3452 17927 3472
rect 17947 3452 17954 3472
rect 17898 3447 17954 3452
rect 18129 3471 18167 3809
rect 18411 3820 18521 3835
rect 18411 3817 18488 3820
rect 18411 3790 18414 3817
rect 18443 3793 18488 3817
rect 18517 3793 18521 3820
rect 18443 3790 18521 3793
rect 18411 3776 18521 3790
rect 18290 3650 18327 3652
rect 18748 3650 18781 3870
rect 19069 3791 19111 3872
rect 19491 3883 19602 3900
rect 19491 3863 19498 3883
rect 19517 3863 19575 3883
rect 19594 3863 19602 3883
rect 19491 3841 19602 3863
rect 18858 3789 18893 3790
rect 18290 3621 18781 3650
rect 18290 3555 18327 3621
rect 18748 3620 18781 3621
rect 18837 3782 18893 3789
rect 18837 3762 18866 3782
rect 18886 3762 18893 3782
rect 18837 3757 18893 3762
rect 19067 3787 19111 3791
rect 19067 3767 19078 3787
rect 19101 3767 19111 3787
rect 19067 3760 19111 3767
rect 19284 3785 19316 3792
rect 19284 3765 19290 3785
rect 19311 3765 19316 3785
rect 19067 3758 19110 3760
rect 18285 3546 18327 3555
rect 18285 3524 18294 3546
rect 18320 3524 18327 3546
rect 18552 3573 18663 3590
rect 18552 3553 18559 3573
rect 18578 3553 18636 3573
rect 18655 3553 18663 3573
rect 18552 3531 18663 3553
rect 18837 3551 18871 3757
rect 19284 3737 19316 3765
rect 18904 3729 19316 3737
rect 18904 3703 18910 3729
rect 18936 3703 19316 3729
rect 18904 3701 19316 3703
rect 18906 3700 18946 3701
rect 19284 3636 19316 3701
rect 19284 3616 19288 3636
rect 19309 3616 19316 3636
rect 19284 3609 19316 3616
rect 18837 3543 18872 3551
rect 18285 3514 18327 3524
rect 18837 3523 18845 3543
rect 18865 3523 18872 3543
rect 18837 3518 18872 3523
rect 19491 3538 19601 3553
rect 19491 3535 19568 3538
rect 18285 3513 18326 3514
rect 18129 3454 18137 3471
rect 18157 3454 18167 3471
rect 17898 3241 17932 3447
rect 18129 3444 18167 3454
rect 18345 3475 18377 3482
rect 18345 3455 18351 3475
rect 18372 3455 18377 3475
rect 18837 3466 18871 3518
rect 19491 3508 19494 3535
rect 19523 3511 19568 3535
rect 19597 3511 19601 3538
rect 19523 3508 19601 3511
rect 19491 3494 19601 3508
rect 19787 3538 19829 3548
rect 19787 3519 19795 3538
rect 19820 3519 19829 3538
rect 19787 3466 19829 3519
rect 18345 3427 18377 3455
rect 18835 3440 19831 3466
rect 17965 3419 18377 3427
rect 17965 3393 17971 3419
rect 17997 3393 18377 3419
rect 17965 3391 18377 3393
rect 17967 3390 18007 3391
rect 18345 3326 18377 3391
rect 18345 3306 18349 3326
rect 18370 3306 18377 3326
rect 18345 3299 18377 3306
rect 18763 3333 18821 3334
rect 18763 3314 19100 3333
rect 19490 3329 19601 3346
rect 18763 3301 19101 3314
rect 17898 3233 17933 3241
rect 17898 3213 17906 3233
rect 17926 3213 17933 3233
rect 17898 3208 17933 3213
rect 18552 3228 18662 3243
rect 18552 3225 18629 3228
rect 17898 3165 17932 3208
rect 18552 3198 18555 3225
rect 18584 3201 18629 3225
rect 18658 3201 18662 3228
rect 18584 3198 18662 3201
rect 18552 3184 18662 3198
rect 18763 3165 18800 3301
rect 19069 3284 19101 3301
rect 19490 3309 19497 3329
rect 19516 3309 19574 3329
rect 19593 3309 19601 3329
rect 19490 3287 19601 3309
rect 19069 3238 19100 3284
rect 18857 3235 18892 3236
rect 18836 3228 18892 3235
rect 18836 3208 18865 3228
rect 18885 3208 18892 3228
rect 18836 3203 18892 3208
rect 19069 3231 19108 3238
rect 19069 3211 19075 3231
rect 19100 3211 19108 3231
rect 19069 3205 19108 3211
rect 19283 3231 19315 3238
rect 19283 3211 19289 3231
rect 19310 3211 19315 3231
rect 17844 3141 17849 3162
rect 17781 3130 17849 3141
rect 17897 3130 18801 3165
rect 17898 3129 17932 3130
rect 17646 3034 18061 3068
rect 17646 3032 17696 3034
rect 17279 2970 17329 2977
rect 17279 2956 17293 2970
rect 17285 2952 17293 2956
rect 17313 2956 17329 2970
rect 17313 2952 17323 2956
rect 17809 2955 17844 2956
rect 17285 2945 17323 2952
rect 17788 2948 17844 2955
rect 17286 2944 17321 2945
rect 17051 2835 17056 2867
rect 17083 2835 17086 2867
rect 17051 2817 17086 2835
rect 17212 2794 17252 2795
rect 16842 2792 17254 2794
rect 16240 2775 16275 2777
rect 15276 2772 16275 2775
rect 13179 2741 13183 2761
rect 13204 2741 13211 2761
rect 13753 2757 14055 2759
rect 13179 2734 13211 2741
rect 13692 2728 14055 2757
rect 13692 2726 13753 2728
rect 12732 2675 12767 2676
rect 12209 2665 12265 2672
rect 12730 2668 12768 2675
rect 12209 2664 12244 2665
rect 10486 2636 10563 2639
rect 10453 2621 10563 2636
rect 11182 2651 11219 2656
rect 11182 2631 11189 2651
rect 11209 2631 11219 2651
rect 12730 2648 12740 2668
rect 12760 2648 12768 2668
rect 11182 2624 11219 2631
rect 12204 2626 12274 2636
rect 11182 2623 11217 2624
rect 10219 2523 10227 2552
rect 10256 2523 10267 2552
rect 10219 2518 10267 2523
rect 10738 2558 10770 2565
rect 10738 2538 10745 2558
rect 10766 2538 10770 2558
rect 9253 2501 9285 2508
rect 10738 2473 10770 2538
rect 11108 2473 11148 2474
rect 10738 2471 11150 2473
rect 10738 2445 11118 2471
rect 11144 2445 11150 2471
rect 8806 2435 8841 2443
rect 8254 2406 8296 2416
rect 8806 2415 8814 2435
rect 8834 2415 8841 2435
rect 8806 2410 8841 2415
rect 9460 2430 9570 2445
rect 9460 2427 9537 2430
rect 8254 2405 8295 2406
rect 7888 2371 7923 2372
rect 7867 2364 7923 2371
rect 7867 2344 7896 2364
rect 7916 2344 7923 2364
rect 7867 2339 7923 2344
rect 8314 2367 8346 2374
rect 8314 2347 8320 2367
rect 8341 2347 8346 2367
rect 8806 2358 8840 2410
rect 9460 2400 9463 2427
rect 9492 2403 9537 2427
rect 9566 2403 9570 2430
rect 9492 2400 9570 2403
rect 9460 2386 9570 2400
rect 9756 2430 9798 2440
rect 9756 2411 9764 2430
rect 9789 2411 9798 2430
rect 9756 2358 9798 2411
rect 10738 2437 11150 2445
rect 10738 2409 10770 2437
rect 11183 2417 11217 2623
rect 12202 2619 12274 2626
rect 11500 2591 11611 2613
rect 11500 2571 11508 2591
rect 11527 2571 11585 2591
rect 11604 2571 11611 2591
rect 11500 2554 11611 2571
rect 12202 2590 12209 2619
rect 12257 2590 12274 2619
rect 12202 2581 12274 2590
rect 12121 2490 12155 2491
rect 11252 2455 12156 2490
rect 10738 2389 10743 2409
rect 10764 2389 10770 2409
rect 10738 2382 10770 2389
rect 10945 2409 10984 2415
rect 10945 2389 10953 2409
rect 10978 2389 10984 2409
rect 10945 2382 10984 2389
rect 11161 2412 11217 2417
rect 11161 2392 11168 2412
rect 11188 2392 11217 2412
rect 11161 2385 11217 2392
rect 11161 2384 11196 2385
rect 7867 2133 7901 2339
rect 8314 2319 8346 2347
rect 8804 2332 9800 2358
rect 10953 2336 10984 2382
rect 7934 2311 8346 2319
rect 7934 2285 7940 2311
rect 7966 2285 8346 2311
rect 7934 2283 8346 2285
rect 7936 2282 7976 2283
rect 8096 2247 8135 2262
rect 8096 2206 8107 2247
rect 8128 2206 8135 2247
rect 7866 2125 7902 2133
rect 7866 2105 7875 2125
rect 7895 2105 7902 2125
rect 7866 2104 7902 2105
rect 7866 2093 7900 2104
rect 7756 2063 7793 2071
rect 7046 2041 7253 2043
rect 7046 1887 7090 2041
rect 7756 2029 8000 2063
rect 6911 1830 6919 1847
rect 6939 1830 6949 1847
rect 6911 1824 6949 1830
rect 6269 1784 6330 1786
rect 5967 1755 6330 1784
rect 6842 1758 6874 1765
rect 5967 1753 6269 1755
rect 3747 1737 4746 1740
rect 6842 1738 6849 1758
rect 6870 1738 6874 1758
rect 3747 1735 3782 1737
rect 2738 1731 3150 1733
rect 2740 1730 2780 1731
rect 3118 1666 3150 1731
rect 6842 1673 6874 1738
rect 7052 1751 7090 1887
rect 7748 1860 7783 1861
rect 7289 1856 7320 1857
rect 7286 1851 7320 1856
rect 7286 1831 7293 1851
rect 7313 1831 7320 1851
rect 7286 1823 7320 1831
rect 7052 1713 7058 1751
rect 7081 1713 7090 1751
rect 7052 1703 7090 1713
rect 7287 1765 7320 1823
rect 7727 1853 7783 1860
rect 7727 1833 7756 1853
rect 7776 1833 7783 1853
rect 7727 1828 7783 1833
rect 7958 1858 8000 2029
rect 8096 1933 8135 2206
rect 8314 2218 8346 2283
rect 10452 2311 10563 2333
rect 10452 2291 10460 2311
rect 10479 2291 10537 2311
rect 10556 2291 10563 2311
rect 10952 2319 10984 2336
rect 11253 2319 11290 2455
rect 11391 2422 11501 2436
rect 11391 2419 11469 2422
rect 11391 2392 11395 2419
rect 11424 2395 11469 2419
rect 11498 2395 11501 2422
rect 12121 2412 12155 2455
rect 11424 2392 11501 2395
rect 11391 2377 11501 2392
rect 12120 2407 12155 2412
rect 12120 2387 12127 2407
rect 12147 2387 12155 2407
rect 12120 2379 12155 2387
rect 10952 2306 11290 2319
rect 10452 2274 10563 2291
rect 10953 2287 11290 2306
rect 11232 2286 11290 2287
rect 11676 2314 11708 2321
rect 11676 2294 11683 2314
rect 11704 2294 11708 2314
rect 8314 2198 8318 2218
rect 8339 2198 8346 2218
rect 8314 2191 8346 2198
rect 8732 2225 8790 2226
rect 8732 2206 9069 2225
rect 9459 2221 9570 2238
rect 8732 2193 9070 2206
rect 8236 2129 8289 2132
rect 8236 2112 8248 2129
rect 8280 2112 8289 2129
rect 8236 2104 8289 2112
rect 8235 2057 8289 2104
rect 8521 2120 8631 2135
rect 8521 2117 8598 2120
rect 8521 2090 8524 2117
rect 8553 2093 8598 2117
rect 8627 2093 8631 2120
rect 8553 2090 8631 2093
rect 8521 2076 8631 2090
rect 8732 2057 8769 2193
rect 9038 2176 9070 2193
rect 9459 2201 9466 2221
rect 9485 2201 9543 2221
rect 9562 2201 9570 2221
rect 9459 2179 9570 2201
rect 11676 2229 11708 2294
rect 12046 2229 12086 2230
rect 11676 2227 12088 2229
rect 11676 2201 12056 2227
rect 12082 2201 12088 2227
rect 11676 2193 12088 2201
rect 9038 2130 9069 2176
rect 10222 2154 11218 2180
rect 11676 2165 11708 2193
rect 8826 2127 8861 2128
rect 8805 2120 8861 2127
rect 8805 2100 8834 2120
rect 8854 2100 8861 2120
rect 8805 2095 8861 2100
rect 9038 2123 9077 2130
rect 9038 2103 9044 2123
rect 9069 2103 9077 2123
rect 9038 2097 9077 2103
rect 9252 2123 9284 2130
rect 9252 2103 9258 2123
rect 9279 2103 9284 2123
rect 8235 2022 8770 2057
rect 8235 2018 8288 2022
rect 8096 1906 8100 1933
rect 8131 1906 8135 1933
rect 8381 1954 8492 1971
rect 8381 1934 8388 1954
rect 8407 1934 8465 1954
rect 8484 1934 8492 1954
rect 8381 1912 8492 1934
rect 8096 1899 8135 1906
rect 8805 1889 8839 2095
rect 9252 2075 9284 2103
rect 8872 2067 9284 2075
rect 10224 2101 10266 2154
rect 10224 2082 10233 2101
rect 10258 2082 10266 2101
rect 10224 2072 10266 2082
rect 10452 2112 10562 2126
rect 10452 2109 10530 2112
rect 10452 2082 10456 2109
rect 10485 2085 10530 2109
rect 10559 2085 10562 2112
rect 11182 2102 11216 2154
rect 11676 2145 11681 2165
rect 11702 2145 11708 2165
rect 11676 2138 11708 2145
rect 11886 2166 11924 2176
rect 12121 2173 12155 2379
rect 11886 2149 11896 2166
rect 11916 2149 11924 2166
rect 11727 2106 11768 2107
rect 10485 2082 10562 2085
rect 10452 2067 10562 2082
rect 11181 2097 11216 2102
rect 11181 2077 11188 2097
rect 11208 2077 11216 2097
rect 11726 2096 11768 2106
rect 11181 2069 11216 2077
rect 8872 2041 8878 2067
rect 8904 2041 9284 2067
rect 8872 2039 9284 2041
rect 8874 2038 8914 2039
rect 9252 1974 9284 2039
rect 10737 2004 10769 2011
rect 9252 1954 9256 1974
rect 9277 1954 9284 1974
rect 9252 1947 9284 1954
rect 9755 1989 9803 1994
rect 9755 1960 9766 1989
rect 9795 1960 9803 1989
rect 8805 1888 8840 1889
rect 8803 1881 8840 1888
rect 7958 1837 7966 1858
rect 7993 1837 8000 1858
rect 7212 1673 7252 1674
rect 6842 1671 7254 1673
rect 6210 1667 6245 1669
rect 3118 1646 3122 1666
rect 3143 1646 3150 1666
rect 5246 1664 6245 1667
rect 3723 1649 4025 1651
rect 3118 1639 3150 1646
rect 3662 1620 4025 1649
rect 3662 1618 3723 1620
rect 2671 1573 2706 1581
rect 2671 1553 2679 1573
rect 2699 1553 2706 1573
rect 2671 1548 2706 1553
rect 3043 1574 3081 1580
rect 3043 1557 3053 1574
rect 3073 1557 3081 1574
rect 2671 1547 2703 1548
rect 2209 1543 2244 1544
rect 1152 1516 1189 1523
rect 1152 1515 1187 1516
rect 189 1415 197 1444
rect 226 1415 237 1444
rect 189 1410 237 1415
rect 708 1450 740 1457
rect 708 1430 715 1450
rect 736 1430 740 1450
rect 708 1365 740 1430
rect 1078 1365 1118 1366
rect 708 1363 1120 1365
rect 708 1337 1088 1363
rect 1114 1337 1120 1363
rect 708 1329 1120 1337
rect 708 1301 740 1329
rect 1153 1309 1187 1515
rect 1857 1498 1896 1505
rect 1500 1470 1611 1492
rect 1500 1450 1508 1470
rect 1527 1450 1585 1470
rect 1604 1450 1611 1470
rect 1500 1433 1611 1450
rect 1857 1471 1861 1498
rect 1892 1471 1896 1498
rect 1704 1382 1757 1386
rect 1222 1347 1757 1382
rect 708 1281 713 1301
rect 734 1281 740 1301
rect 708 1274 740 1281
rect 915 1301 954 1307
rect 915 1281 923 1301
rect 948 1281 954 1301
rect 915 1274 954 1281
rect 1131 1304 1187 1309
rect 1131 1284 1138 1304
rect 1158 1284 1187 1304
rect 1131 1277 1187 1284
rect 1131 1276 1166 1277
rect 923 1228 954 1274
rect 422 1203 533 1225
rect 422 1183 430 1203
rect 449 1183 507 1203
rect 526 1183 533 1203
rect 922 1211 954 1228
rect 1223 1211 1260 1347
rect 1361 1314 1471 1328
rect 1361 1311 1439 1314
rect 1361 1284 1365 1311
rect 1394 1287 1439 1311
rect 1468 1287 1471 1314
rect 1394 1284 1471 1287
rect 1361 1269 1471 1284
rect 1703 1300 1757 1347
rect 1703 1292 1756 1300
rect 1703 1275 1712 1292
rect 1744 1275 1756 1292
rect 1703 1272 1756 1275
rect 922 1198 1260 1211
rect 422 1166 533 1183
rect 923 1179 1260 1198
rect 1202 1178 1260 1179
rect 1646 1206 1678 1213
rect 1646 1186 1653 1206
rect 1674 1186 1678 1206
rect 1646 1121 1678 1186
rect 1857 1198 1896 1471
rect 2092 1300 2126 1311
rect 2090 1299 2126 1300
rect 2090 1279 2097 1299
rect 2117 1279 2126 1299
rect 2090 1271 2126 1279
rect 1857 1157 1864 1198
rect 1885 1157 1896 1198
rect 1857 1142 1896 1157
rect 2016 1121 2056 1122
rect 1646 1119 2058 1121
rect 1646 1093 2026 1119
rect 2052 1093 2058 1119
rect 1646 1085 2058 1093
rect 192 1046 1188 1072
rect 1646 1057 1678 1085
rect 2091 1065 2125 1271
rect 2833 1227 2868 1228
rect 194 993 236 1046
rect 194 974 203 993
rect 228 974 236 993
rect 194 964 236 974
rect 422 1004 532 1018
rect 422 1001 500 1004
rect 422 974 426 1001
rect 455 977 500 1001
rect 529 977 532 1004
rect 1152 994 1186 1046
rect 1646 1037 1651 1057
rect 1672 1037 1678 1057
rect 1646 1030 1678 1037
rect 2069 1060 2125 1065
rect 2069 1040 2076 1060
rect 2096 1040 2125 1060
rect 2069 1033 2125 1040
rect 2812 1220 2868 1227
rect 2812 1200 2841 1220
rect 2861 1200 2868 1220
rect 2812 1195 2868 1200
rect 3043 1219 3081 1557
rect 3325 1568 3435 1583
rect 3325 1565 3402 1568
rect 3325 1538 3328 1565
rect 3357 1541 3402 1565
rect 3431 1541 3435 1568
rect 3357 1538 3435 1541
rect 3325 1524 3435 1538
rect 3204 1398 3241 1400
rect 3662 1398 3695 1618
rect 3983 1539 4025 1620
rect 4405 1631 4516 1648
rect 4405 1611 4412 1631
rect 4431 1611 4489 1631
rect 4508 1611 4516 1631
rect 4405 1589 4516 1611
rect 5245 1640 6245 1664
rect 3772 1537 3807 1538
rect 3204 1369 3695 1398
rect 3204 1303 3241 1369
rect 3662 1368 3695 1369
rect 3751 1530 3807 1537
rect 3751 1510 3780 1530
rect 3800 1510 3807 1530
rect 3751 1505 3807 1510
rect 3981 1535 4025 1539
rect 3981 1515 3992 1535
rect 4015 1515 4025 1535
rect 3981 1508 4025 1515
rect 4198 1533 4230 1540
rect 4198 1513 4204 1533
rect 4225 1513 4230 1533
rect 3981 1506 4024 1508
rect 3199 1294 3241 1303
rect 3199 1272 3208 1294
rect 3234 1272 3241 1294
rect 3466 1321 3577 1338
rect 3466 1301 3473 1321
rect 3492 1301 3550 1321
rect 3569 1301 3577 1321
rect 3466 1279 3577 1301
rect 3751 1299 3785 1505
rect 4198 1485 4230 1513
rect 3818 1477 4230 1485
rect 3818 1451 3824 1477
rect 3850 1451 4230 1477
rect 5245 1485 5293 1640
rect 5479 1599 5589 1613
rect 5479 1596 5557 1599
rect 5479 1569 5483 1596
rect 5512 1572 5557 1596
rect 5586 1572 5589 1599
rect 6210 1589 6245 1640
rect 5512 1569 5589 1572
rect 5479 1554 5589 1569
rect 6208 1584 6245 1589
rect 6208 1564 6215 1584
rect 6235 1564 6245 1584
rect 6842 1645 7222 1671
rect 7248 1645 7254 1671
rect 6842 1637 7254 1645
rect 6842 1609 6874 1637
rect 7287 1617 7323 1765
rect 6842 1589 6847 1609
rect 6868 1589 6874 1609
rect 6842 1582 6874 1589
rect 7265 1612 7323 1617
rect 7265 1592 7272 1612
rect 7292 1592 7323 1612
rect 7265 1585 7323 1592
rect 7727 1622 7761 1828
rect 7958 1826 8000 1837
rect 8174 1856 8206 1863
rect 8174 1836 8180 1856
rect 8201 1836 8206 1856
rect 8174 1808 8206 1836
rect 7794 1800 8206 1808
rect 7794 1774 7800 1800
rect 7826 1774 8206 1800
rect 8803 1861 8813 1881
rect 8833 1861 8840 1881
rect 8803 1856 8840 1861
rect 9459 1876 9569 1891
rect 9459 1873 9536 1876
rect 8803 1805 8838 1856
rect 9459 1846 9462 1873
rect 9491 1849 9536 1873
rect 9565 1849 9569 1876
rect 9491 1846 9569 1849
rect 9459 1832 9569 1846
rect 9755 1805 9803 1960
rect 10737 1984 10744 2004
rect 10765 1984 10769 2004
rect 10737 1919 10769 1984
rect 11107 1919 11147 1920
rect 10737 1917 11149 1919
rect 10737 1891 11117 1917
rect 11143 1891 11149 1917
rect 10737 1883 11149 1891
rect 10737 1855 10769 1883
rect 11182 1863 11216 2069
rect 11390 2067 11501 2089
rect 11390 2047 11398 2067
rect 11417 2047 11475 2067
rect 11494 2047 11501 2067
rect 11390 2030 11501 2047
rect 11726 2074 11733 2096
rect 11759 2074 11768 2096
rect 11726 2065 11768 2074
rect 10943 1860 10986 1862
rect 10737 1835 10742 1855
rect 10763 1835 10769 1855
rect 10737 1828 10769 1835
rect 10942 1853 10986 1860
rect 10942 1833 10952 1853
rect 10975 1833 10986 1853
rect 10942 1829 10986 1833
rect 11160 1858 11216 1863
rect 11160 1838 11167 1858
rect 11187 1838 11216 1858
rect 11160 1831 11216 1838
rect 11272 1999 11305 2000
rect 11726 1999 11763 2065
rect 11272 1970 11763 1999
rect 11160 1830 11195 1831
rect 8803 1781 9803 1805
rect 8803 1778 9802 1781
rect 8803 1776 8838 1778
rect 7794 1772 8206 1774
rect 7796 1771 7836 1772
rect 8174 1707 8206 1772
rect 10451 1757 10562 1779
rect 10451 1737 10459 1757
rect 10478 1737 10536 1757
rect 10555 1737 10562 1757
rect 10451 1720 10562 1737
rect 10942 1748 10984 1829
rect 11272 1750 11305 1970
rect 11726 1968 11763 1970
rect 11532 1830 11642 1844
rect 11532 1827 11610 1830
rect 11532 1800 11536 1827
rect 11565 1803 11610 1827
rect 11639 1803 11642 1830
rect 11565 1800 11642 1803
rect 11532 1785 11642 1800
rect 11886 1811 11924 2149
rect 12099 2168 12155 2173
rect 12099 2148 12106 2168
rect 12126 2148 12155 2168
rect 12099 2141 12155 2148
rect 12099 2140 12134 2141
rect 12021 2040 12065 2044
rect 12202 2040 12252 2581
rect 12021 2007 12252 2040
rect 12730 2035 12768 2648
rect 13386 2663 13496 2678
rect 13386 2660 13463 2663
rect 13386 2633 13389 2660
rect 13418 2636 13463 2660
rect 13492 2636 13496 2663
rect 13418 2633 13496 2636
rect 13386 2619 13496 2633
rect 13234 2506 13271 2508
rect 13692 2506 13725 2726
rect 14013 2647 14055 2728
rect 14435 2739 14546 2755
rect 14435 2719 14442 2739
rect 14461 2719 14519 2739
rect 14538 2719 14546 2739
rect 14435 2697 14546 2719
rect 15275 2748 16275 2772
rect 13802 2645 13837 2646
rect 13234 2477 13725 2506
rect 13234 2411 13271 2477
rect 13692 2476 13725 2477
rect 13781 2638 13837 2645
rect 13781 2618 13810 2638
rect 13830 2618 13837 2638
rect 13781 2613 13837 2618
rect 14011 2643 14055 2647
rect 14011 2623 14022 2643
rect 14045 2623 14055 2643
rect 14011 2616 14055 2623
rect 14228 2641 14260 2648
rect 14228 2621 14234 2641
rect 14255 2621 14260 2641
rect 14011 2614 14054 2616
rect 13229 2402 13271 2411
rect 13229 2380 13238 2402
rect 13264 2380 13271 2402
rect 13496 2429 13607 2446
rect 13496 2409 13503 2429
rect 13522 2409 13580 2429
rect 13599 2409 13607 2429
rect 13496 2387 13607 2409
rect 13781 2407 13815 2613
rect 14228 2593 14260 2621
rect 13848 2585 14260 2593
rect 13848 2559 13854 2585
rect 13880 2559 14260 2585
rect 15275 2593 15323 2748
rect 15509 2707 15619 2721
rect 15509 2704 15587 2707
rect 15509 2677 15513 2704
rect 15542 2680 15587 2704
rect 15616 2680 15619 2707
rect 16240 2697 16275 2748
rect 16842 2766 17222 2792
rect 17248 2766 17254 2792
rect 16842 2758 17254 2766
rect 16842 2730 16874 2758
rect 17287 2738 17321 2944
rect 16842 2710 16847 2730
rect 16868 2710 16874 2730
rect 16842 2703 16874 2710
rect 17265 2733 17321 2738
rect 17265 2713 17272 2733
rect 17292 2713 17321 2733
rect 17788 2928 17817 2948
rect 17837 2928 17844 2948
rect 17788 2923 17844 2928
rect 18016 2951 18061 3034
rect 18442 3049 18553 3066
rect 18442 3029 18449 3049
rect 18468 3029 18526 3049
rect 18545 3029 18553 3049
rect 18442 3007 18553 3029
rect 18836 2997 18870 3203
rect 19283 3183 19315 3211
rect 18903 3175 19315 3183
rect 18903 3149 18909 3175
rect 18935 3149 19315 3175
rect 18903 3147 19315 3149
rect 18905 3146 18945 3147
rect 19283 3082 19315 3147
rect 19283 3062 19287 3082
rect 19308 3062 19315 3082
rect 19283 3055 19315 3062
rect 19786 3097 19834 3102
rect 19786 3068 19797 3097
rect 19826 3068 19834 3097
rect 18836 2996 18871 2997
rect 18834 2989 18871 2996
rect 18834 2969 18844 2989
rect 18864 2969 18871 2989
rect 18834 2964 18871 2969
rect 19490 2984 19600 2999
rect 19490 2981 19567 2984
rect 18016 2932 18025 2951
rect 18054 2932 18061 2951
rect 17788 2717 17822 2923
rect 18016 2920 18061 2932
rect 18235 2951 18267 2958
rect 18235 2931 18241 2951
rect 18262 2931 18267 2951
rect 18235 2903 18267 2931
rect 17855 2895 18267 2903
rect 17855 2869 17861 2895
rect 17887 2869 18267 2895
rect 18834 2913 18869 2964
rect 19490 2954 19493 2981
rect 19522 2957 19567 2981
rect 19596 2957 19600 2984
rect 19522 2954 19600 2957
rect 19490 2940 19600 2954
rect 19786 2913 19834 3068
rect 18834 2889 19834 2913
rect 18834 2886 19833 2889
rect 18834 2884 18869 2886
rect 17855 2867 18267 2869
rect 17857 2866 17897 2867
rect 18235 2802 18267 2867
rect 18235 2782 18239 2802
rect 18260 2782 18267 2802
rect 18809 2798 19111 2800
rect 18235 2775 18267 2782
rect 18748 2769 19111 2798
rect 18748 2767 18809 2769
rect 17788 2716 17823 2717
rect 17265 2706 17321 2713
rect 17786 2709 17824 2716
rect 17265 2705 17300 2706
rect 15542 2677 15619 2680
rect 15509 2662 15619 2677
rect 16238 2692 16275 2697
rect 16238 2672 16245 2692
rect 16265 2672 16275 2692
rect 17786 2689 17796 2709
rect 17816 2689 17824 2709
rect 16238 2665 16275 2672
rect 17260 2667 17330 2677
rect 16238 2664 16273 2665
rect 15275 2564 15283 2593
rect 15312 2564 15323 2593
rect 15275 2559 15323 2564
rect 15794 2599 15826 2606
rect 15794 2579 15801 2599
rect 15822 2579 15826 2599
rect 13848 2557 14260 2559
rect 13850 2556 13890 2557
rect 14228 2492 14260 2557
rect 14228 2472 14232 2492
rect 14253 2472 14260 2492
rect 14228 2465 14260 2472
rect 15794 2514 15826 2579
rect 16164 2514 16204 2515
rect 15794 2512 16206 2514
rect 15794 2486 16174 2512
rect 16200 2486 16206 2512
rect 15794 2478 16206 2486
rect 15794 2450 15826 2478
rect 16239 2458 16273 2664
rect 17258 2660 17330 2667
rect 16556 2632 16667 2654
rect 16556 2612 16564 2632
rect 16583 2612 16641 2632
rect 16660 2612 16667 2632
rect 16556 2595 16667 2612
rect 17258 2631 17265 2660
rect 17313 2631 17330 2660
rect 17258 2622 17330 2631
rect 17177 2531 17211 2532
rect 16308 2496 17212 2531
rect 15794 2430 15799 2450
rect 15820 2430 15826 2450
rect 15794 2423 15826 2430
rect 16001 2450 16040 2456
rect 16001 2430 16009 2450
rect 16034 2430 16040 2450
rect 16001 2423 16040 2430
rect 16217 2453 16273 2458
rect 16217 2433 16224 2453
rect 16244 2433 16273 2453
rect 16217 2426 16273 2433
rect 16217 2425 16252 2426
rect 13781 2399 13816 2407
rect 13229 2370 13271 2380
rect 13781 2379 13789 2399
rect 13809 2379 13816 2399
rect 13781 2374 13816 2379
rect 14435 2394 14545 2409
rect 14435 2391 14512 2394
rect 13229 2369 13270 2370
rect 12863 2335 12898 2336
rect 12842 2328 12898 2335
rect 12842 2308 12871 2328
rect 12891 2308 12898 2328
rect 12842 2303 12898 2308
rect 13289 2331 13321 2338
rect 13289 2311 13295 2331
rect 13316 2311 13321 2331
rect 13781 2322 13815 2374
rect 14435 2364 14438 2391
rect 14467 2367 14512 2391
rect 14541 2367 14545 2394
rect 14467 2364 14545 2367
rect 14435 2350 14545 2364
rect 14731 2394 14773 2404
rect 14731 2375 14739 2394
rect 14764 2375 14773 2394
rect 16009 2377 16040 2423
rect 14731 2322 14773 2375
rect 15508 2352 15619 2374
rect 15508 2332 15516 2352
rect 15535 2332 15593 2352
rect 15612 2332 15619 2352
rect 16008 2360 16040 2377
rect 16309 2360 16346 2496
rect 16447 2463 16557 2477
rect 16447 2460 16525 2463
rect 16447 2433 16451 2460
rect 16480 2436 16525 2460
rect 16554 2436 16557 2463
rect 17177 2453 17211 2496
rect 16480 2433 16557 2436
rect 16447 2418 16557 2433
rect 17176 2448 17211 2453
rect 17176 2428 17183 2448
rect 17203 2428 17211 2448
rect 17176 2420 17211 2428
rect 16008 2347 16346 2360
rect 12842 2097 12876 2303
rect 13289 2283 13321 2311
rect 13779 2296 14775 2322
rect 15508 2315 15619 2332
rect 16009 2328 16346 2347
rect 16288 2327 16346 2328
rect 16732 2355 16764 2362
rect 16732 2335 16739 2355
rect 16760 2335 16764 2355
rect 12909 2275 13321 2283
rect 12909 2249 12915 2275
rect 12941 2249 13321 2275
rect 12909 2247 13321 2249
rect 12911 2246 12951 2247
rect 13071 2211 13110 2226
rect 13071 2170 13082 2211
rect 13103 2170 13110 2211
rect 12841 2089 12877 2097
rect 12841 2069 12850 2089
rect 12870 2069 12877 2089
rect 12841 2068 12877 2069
rect 12841 2057 12875 2068
rect 12731 2027 12768 2035
rect 12021 2005 12228 2007
rect 12021 1851 12065 2005
rect 12731 1993 12975 2027
rect 11886 1794 11894 1811
rect 11914 1794 11924 1811
rect 11886 1788 11924 1794
rect 11244 1748 11305 1750
rect 10942 1719 11305 1748
rect 11817 1722 11849 1729
rect 10942 1717 11244 1719
rect 8174 1687 8178 1707
rect 8199 1687 8206 1707
rect 11817 1702 11824 1722
rect 11845 1702 11849 1722
rect 8779 1690 9081 1692
rect 8174 1680 8206 1687
rect 8718 1661 9081 1690
rect 8718 1659 8779 1661
rect 7727 1614 7762 1622
rect 7727 1594 7735 1614
rect 7755 1594 7762 1614
rect 7727 1589 7762 1594
rect 8099 1615 8137 1621
rect 8099 1598 8109 1615
rect 8129 1598 8137 1615
rect 7727 1588 7759 1589
rect 7265 1584 7300 1585
rect 6208 1557 6245 1564
rect 6208 1556 6243 1557
rect 5245 1456 5253 1485
rect 5282 1456 5293 1485
rect 5245 1451 5293 1456
rect 5764 1491 5796 1498
rect 5764 1471 5771 1491
rect 5792 1471 5796 1491
rect 3818 1449 4230 1451
rect 3820 1448 3860 1449
rect 4198 1384 4230 1449
rect 4198 1364 4202 1384
rect 4223 1364 4230 1384
rect 4198 1357 4230 1364
rect 5764 1406 5796 1471
rect 6134 1406 6174 1407
rect 5764 1404 6176 1406
rect 5764 1378 6144 1404
rect 6170 1378 6176 1404
rect 5764 1370 6176 1378
rect 5764 1342 5796 1370
rect 6209 1350 6243 1556
rect 6913 1539 6952 1546
rect 6556 1511 6667 1533
rect 6556 1491 6564 1511
rect 6583 1491 6641 1511
rect 6660 1491 6667 1511
rect 6556 1474 6667 1491
rect 6913 1512 6917 1539
rect 6948 1512 6952 1539
rect 6760 1423 6813 1427
rect 6278 1388 6813 1423
rect 5764 1322 5769 1342
rect 5790 1322 5796 1342
rect 5764 1315 5796 1322
rect 5971 1342 6010 1348
rect 5971 1322 5979 1342
rect 6004 1322 6010 1342
rect 5971 1315 6010 1322
rect 6187 1345 6243 1350
rect 6187 1325 6194 1345
rect 6214 1325 6243 1345
rect 6187 1318 6243 1325
rect 6187 1317 6222 1318
rect 3751 1291 3786 1299
rect 3199 1262 3241 1272
rect 3751 1271 3759 1291
rect 3779 1271 3786 1291
rect 3751 1266 3786 1271
rect 4405 1286 4515 1301
rect 4405 1283 4482 1286
rect 3199 1261 3240 1262
rect 3043 1202 3051 1219
rect 3071 1202 3081 1219
rect 2069 1032 2104 1033
rect 1697 998 1738 999
rect 455 974 532 977
rect 422 959 532 974
rect 1151 989 1186 994
rect 1151 969 1158 989
rect 1178 969 1186 989
rect 1696 988 1738 998
rect 1151 961 1186 969
rect 707 896 739 903
rect 707 876 714 896
rect 735 876 739 896
rect 707 811 739 876
rect 1077 811 1117 812
rect 707 809 1119 811
rect 707 783 1087 809
rect 1113 783 1119 809
rect 707 775 1119 783
rect 707 747 739 775
rect 1152 755 1186 961
rect 1360 959 1471 981
rect 1360 939 1368 959
rect 1387 939 1445 959
rect 1464 939 1471 959
rect 1360 922 1471 939
rect 1696 966 1703 988
rect 1729 966 1738 988
rect 1696 957 1738 966
rect 2812 989 2846 1195
rect 3043 1192 3081 1202
rect 3259 1223 3291 1230
rect 3259 1203 3265 1223
rect 3286 1203 3291 1223
rect 3751 1214 3785 1266
rect 4405 1256 4408 1283
rect 4437 1259 4482 1283
rect 4511 1259 4515 1286
rect 4437 1256 4515 1259
rect 4405 1242 4515 1256
rect 4701 1286 4743 1296
rect 4701 1267 4709 1286
rect 4734 1267 4743 1286
rect 5979 1269 6010 1315
rect 4701 1214 4743 1267
rect 5478 1244 5589 1266
rect 5478 1224 5486 1244
rect 5505 1224 5563 1244
rect 5582 1224 5589 1244
rect 5978 1252 6010 1269
rect 6279 1252 6316 1388
rect 6417 1355 6527 1369
rect 6417 1352 6495 1355
rect 6417 1325 6421 1352
rect 6450 1328 6495 1352
rect 6524 1328 6527 1355
rect 6450 1325 6527 1328
rect 6417 1310 6527 1325
rect 6759 1341 6813 1388
rect 6759 1333 6812 1341
rect 6759 1316 6768 1333
rect 6800 1316 6812 1333
rect 6759 1313 6812 1316
rect 5978 1239 6316 1252
rect 3259 1175 3291 1203
rect 3749 1188 4745 1214
rect 5478 1207 5589 1224
rect 5979 1220 6316 1239
rect 6258 1219 6316 1220
rect 6702 1247 6734 1254
rect 6702 1227 6709 1247
rect 6730 1227 6734 1247
rect 2879 1167 3291 1175
rect 2879 1141 2885 1167
rect 2911 1141 3291 1167
rect 2879 1139 3291 1141
rect 2881 1138 2921 1139
rect 3259 1074 3291 1139
rect 6702 1162 6734 1227
rect 6913 1239 6952 1512
rect 7148 1341 7182 1352
rect 7146 1340 7182 1341
rect 7146 1320 7153 1340
rect 7173 1320 7182 1340
rect 7146 1312 7182 1320
rect 6913 1198 6920 1239
rect 6941 1198 6952 1239
rect 6913 1183 6952 1198
rect 7072 1162 7112 1163
rect 6702 1160 7114 1162
rect 6702 1134 7082 1160
rect 7108 1134 7114 1160
rect 6702 1126 7114 1134
rect 3259 1054 3263 1074
rect 3284 1054 3291 1074
rect 3259 1047 3291 1054
rect 3677 1081 3735 1082
rect 3677 1062 4014 1081
rect 4404 1077 4515 1094
rect 5248 1087 6244 1113
rect 6702 1098 6734 1126
rect 7147 1106 7181 1312
rect 7889 1268 7924 1269
rect 3677 1049 4015 1062
rect 2812 981 2847 989
rect 2812 961 2820 981
rect 2840 961 2847 981
rect 913 752 956 754
rect 707 727 712 747
rect 733 727 739 747
rect 707 720 739 727
rect 912 745 956 752
rect 912 725 922 745
rect 945 725 956 745
rect 912 721 956 725
rect 1130 750 1186 755
rect 1130 730 1137 750
rect 1157 730 1186 750
rect 1130 723 1186 730
rect 1242 891 1275 892
rect 1696 891 1733 957
rect 2812 956 2847 961
rect 3466 976 3576 991
rect 3466 973 3543 976
rect 2812 913 2846 956
rect 3466 946 3469 973
rect 3498 949 3543 973
rect 3572 949 3576 976
rect 3498 946 3576 949
rect 3466 932 3576 946
rect 3677 913 3714 1049
rect 3983 1032 4015 1049
rect 4404 1057 4411 1077
rect 4430 1057 4488 1077
rect 4507 1057 4515 1077
rect 4404 1035 4515 1057
rect 5250 1034 5292 1087
rect 3983 986 4014 1032
rect 5250 1015 5259 1034
rect 5284 1015 5292 1034
rect 5250 1005 5292 1015
rect 5478 1045 5588 1059
rect 5478 1042 5556 1045
rect 5478 1015 5482 1042
rect 5511 1018 5556 1042
rect 5585 1018 5588 1045
rect 6208 1035 6242 1087
rect 6702 1078 6707 1098
rect 6728 1078 6734 1098
rect 6702 1071 6734 1078
rect 7125 1101 7181 1106
rect 7125 1081 7132 1101
rect 7152 1081 7181 1101
rect 7125 1074 7181 1081
rect 7868 1261 7924 1268
rect 7868 1241 7897 1261
rect 7917 1241 7924 1261
rect 7868 1236 7924 1241
rect 8099 1260 8137 1598
rect 8381 1609 8491 1624
rect 8381 1606 8458 1609
rect 8381 1579 8384 1606
rect 8413 1582 8458 1606
rect 8487 1582 8491 1609
rect 8413 1579 8491 1582
rect 8381 1565 8491 1579
rect 8260 1439 8297 1441
rect 8718 1439 8751 1659
rect 9039 1580 9081 1661
rect 9461 1672 9572 1689
rect 9461 1652 9468 1672
rect 9487 1652 9545 1672
rect 9564 1652 9572 1672
rect 9461 1630 9572 1652
rect 11817 1637 11849 1702
rect 12027 1715 12065 1851
rect 12723 1824 12758 1825
rect 12264 1820 12295 1821
rect 12261 1815 12295 1820
rect 12261 1795 12268 1815
rect 12288 1795 12295 1815
rect 12261 1787 12295 1795
rect 12027 1677 12033 1715
rect 12056 1677 12065 1715
rect 12027 1667 12065 1677
rect 12262 1729 12295 1787
rect 12702 1817 12758 1824
rect 12702 1797 12731 1817
rect 12751 1797 12758 1817
rect 12702 1792 12758 1797
rect 12933 1822 12975 1993
rect 13071 1897 13110 2170
rect 13289 2182 13321 2247
rect 16732 2270 16764 2335
rect 17102 2270 17142 2271
rect 16732 2268 17144 2270
rect 16732 2242 17112 2268
rect 17138 2242 17144 2268
rect 16732 2234 17144 2242
rect 13289 2162 13293 2182
rect 13314 2162 13321 2182
rect 13289 2155 13321 2162
rect 13707 2189 13765 2190
rect 13707 2170 14044 2189
rect 14434 2185 14545 2202
rect 15278 2195 16274 2221
rect 16732 2206 16764 2234
rect 13707 2157 14045 2170
rect 13211 2093 13264 2096
rect 13211 2076 13223 2093
rect 13255 2076 13264 2093
rect 13211 2068 13264 2076
rect 13210 2021 13264 2068
rect 13496 2084 13606 2099
rect 13496 2081 13573 2084
rect 13496 2054 13499 2081
rect 13528 2057 13573 2081
rect 13602 2057 13606 2084
rect 13528 2054 13606 2057
rect 13496 2040 13606 2054
rect 13707 2021 13744 2157
rect 14013 2140 14045 2157
rect 14434 2165 14441 2185
rect 14460 2165 14518 2185
rect 14537 2165 14545 2185
rect 14434 2143 14545 2165
rect 15280 2142 15322 2195
rect 14013 2094 14044 2140
rect 15280 2123 15289 2142
rect 15314 2123 15322 2142
rect 15280 2113 15322 2123
rect 15508 2153 15618 2167
rect 15508 2150 15586 2153
rect 15508 2123 15512 2150
rect 15541 2126 15586 2150
rect 15615 2126 15618 2153
rect 16238 2143 16272 2195
rect 16732 2186 16737 2206
rect 16758 2186 16764 2206
rect 16732 2179 16764 2186
rect 16942 2207 16980 2217
rect 17177 2214 17211 2420
rect 16942 2190 16952 2207
rect 16972 2190 16980 2207
rect 16783 2147 16824 2148
rect 15541 2123 15618 2126
rect 15508 2108 15618 2123
rect 16237 2138 16272 2143
rect 16237 2118 16244 2138
rect 16264 2118 16272 2138
rect 16782 2137 16824 2147
rect 16237 2110 16272 2118
rect 13801 2091 13836 2092
rect 13780 2084 13836 2091
rect 13780 2064 13809 2084
rect 13829 2064 13836 2084
rect 13780 2059 13836 2064
rect 14013 2087 14052 2094
rect 14013 2067 14019 2087
rect 14044 2067 14052 2087
rect 14013 2061 14052 2067
rect 14227 2087 14259 2094
rect 14227 2067 14233 2087
rect 14254 2067 14259 2087
rect 13210 1986 13745 2021
rect 13210 1982 13263 1986
rect 13071 1870 13075 1897
rect 13106 1870 13110 1897
rect 13356 1918 13467 1935
rect 13356 1898 13363 1918
rect 13382 1898 13440 1918
rect 13459 1898 13467 1918
rect 13356 1876 13467 1898
rect 13071 1863 13110 1870
rect 13780 1853 13814 2059
rect 14227 2039 14259 2067
rect 13847 2031 14259 2039
rect 13847 2005 13853 2031
rect 13879 2005 14259 2031
rect 13847 2003 14259 2005
rect 13849 2002 13889 2003
rect 14227 1938 14259 2003
rect 15793 2045 15825 2052
rect 15793 2025 15800 2045
rect 15821 2025 15825 2045
rect 15793 1960 15825 2025
rect 16163 1960 16203 1961
rect 15793 1958 16205 1960
rect 14227 1918 14231 1938
rect 14252 1918 14259 1938
rect 14227 1911 14259 1918
rect 14730 1953 14778 1958
rect 14730 1924 14741 1953
rect 14770 1924 14778 1953
rect 13780 1852 13815 1853
rect 13778 1845 13815 1852
rect 12933 1801 12941 1822
rect 12968 1801 12975 1822
rect 12187 1637 12227 1638
rect 11817 1635 12229 1637
rect 11185 1631 11220 1633
rect 10221 1628 11220 1631
rect 10220 1604 11220 1628
rect 8828 1578 8863 1579
rect 8260 1410 8751 1439
rect 8260 1344 8297 1410
rect 8718 1409 8751 1410
rect 8807 1571 8863 1578
rect 8807 1551 8836 1571
rect 8856 1551 8863 1571
rect 8807 1546 8863 1551
rect 9037 1576 9081 1580
rect 9037 1556 9048 1576
rect 9071 1556 9081 1576
rect 9037 1549 9081 1556
rect 9254 1574 9286 1581
rect 9254 1554 9260 1574
rect 9281 1554 9286 1574
rect 9037 1547 9080 1549
rect 8255 1335 8297 1344
rect 8255 1313 8264 1335
rect 8290 1313 8297 1335
rect 8522 1362 8633 1379
rect 8522 1342 8529 1362
rect 8548 1342 8606 1362
rect 8625 1342 8633 1362
rect 8522 1320 8633 1342
rect 8807 1340 8841 1546
rect 9254 1526 9286 1554
rect 8874 1518 9286 1526
rect 8874 1492 8880 1518
rect 8906 1492 9286 1518
rect 8874 1490 9286 1492
rect 8876 1489 8916 1490
rect 9254 1425 9286 1490
rect 9254 1405 9258 1425
rect 9279 1405 9286 1425
rect 10220 1449 10268 1604
rect 10454 1563 10564 1577
rect 10454 1560 10532 1563
rect 10454 1533 10458 1560
rect 10487 1536 10532 1560
rect 10561 1536 10564 1563
rect 11185 1553 11220 1604
rect 10487 1533 10564 1536
rect 10454 1518 10564 1533
rect 11183 1548 11220 1553
rect 11183 1528 11190 1548
rect 11210 1528 11220 1548
rect 11817 1609 12197 1635
rect 12223 1609 12229 1635
rect 11817 1601 12229 1609
rect 11817 1573 11849 1601
rect 12262 1581 12298 1729
rect 11817 1553 11822 1573
rect 11843 1553 11849 1573
rect 11817 1546 11849 1553
rect 12240 1576 12298 1581
rect 12240 1556 12247 1576
rect 12267 1556 12298 1576
rect 12240 1549 12298 1556
rect 12702 1586 12736 1792
rect 12933 1790 12975 1801
rect 13149 1820 13181 1827
rect 13149 1800 13155 1820
rect 13176 1800 13181 1820
rect 13149 1772 13181 1800
rect 12769 1764 13181 1772
rect 12769 1738 12775 1764
rect 12801 1738 13181 1764
rect 13778 1825 13788 1845
rect 13808 1825 13815 1845
rect 13778 1820 13815 1825
rect 14434 1840 14544 1855
rect 14434 1837 14511 1840
rect 13778 1769 13813 1820
rect 14434 1810 14437 1837
rect 14466 1813 14511 1837
rect 14540 1813 14544 1840
rect 14466 1810 14544 1813
rect 14434 1796 14544 1810
rect 14730 1769 14778 1924
rect 15793 1932 16173 1958
rect 16199 1932 16205 1958
rect 15793 1924 16205 1932
rect 15793 1896 15825 1924
rect 16238 1904 16272 2110
rect 16446 2108 16557 2130
rect 16446 2088 16454 2108
rect 16473 2088 16531 2108
rect 16550 2088 16557 2108
rect 16446 2071 16557 2088
rect 16782 2115 16789 2137
rect 16815 2115 16824 2137
rect 16782 2106 16824 2115
rect 15999 1901 16042 1903
rect 15793 1876 15798 1896
rect 15819 1876 15825 1896
rect 15793 1869 15825 1876
rect 15998 1894 16042 1901
rect 15998 1874 16008 1894
rect 16031 1874 16042 1894
rect 15998 1870 16042 1874
rect 16216 1899 16272 1904
rect 16216 1879 16223 1899
rect 16243 1879 16272 1899
rect 16216 1872 16272 1879
rect 16328 2040 16361 2041
rect 16782 2040 16819 2106
rect 16328 2011 16819 2040
rect 16216 1871 16251 1872
rect 13778 1745 14778 1769
rect 15507 1798 15618 1820
rect 15507 1778 15515 1798
rect 15534 1778 15592 1798
rect 15611 1778 15618 1798
rect 15507 1761 15618 1778
rect 15998 1789 16040 1870
rect 16328 1791 16361 2011
rect 16782 2009 16819 2011
rect 16588 1871 16698 1885
rect 16588 1868 16666 1871
rect 16588 1841 16592 1868
rect 16621 1844 16666 1868
rect 16695 1844 16698 1871
rect 16621 1841 16698 1844
rect 16588 1826 16698 1841
rect 16942 1852 16980 2190
rect 17155 2209 17211 2214
rect 17155 2189 17162 2209
rect 17182 2189 17211 2209
rect 17155 2182 17211 2189
rect 17155 2181 17190 2182
rect 17077 2081 17121 2085
rect 17258 2081 17308 2622
rect 17077 2048 17308 2081
rect 17786 2076 17824 2689
rect 18442 2704 18552 2719
rect 18442 2701 18519 2704
rect 18442 2674 18445 2701
rect 18474 2677 18519 2701
rect 18548 2677 18552 2704
rect 18474 2674 18552 2677
rect 18442 2660 18552 2674
rect 18290 2547 18327 2549
rect 18748 2547 18781 2767
rect 19069 2688 19111 2769
rect 19491 2780 19602 2796
rect 19491 2760 19498 2780
rect 19517 2760 19575 2780
rect 19594 2760 19602 2780
rect 19491 2738 19602 2760
rect 18858 2686 18893 2687
rect 18290 2518 18781 2547
rect 18290 2452 18327 2518
rect 18748 2517 18781 2518
rect 18837 2679 18893 2686
rect 18837 2659 18866 2679
rect 18886 2659 18893 2679
rect 18837 2654 18893 2659
rect 19067 2684 19111 2688
rect 19067 2664 19078 2684
rect 19101 2664 19111 2684
rect 19067 2657 19111 2664
rect 19284 2682 19316 2689
rect 19284 2662 19290 2682
rect 19311 2662 19316 2682
rect 19067 2655 19110 2657
rect 18285 2443 18327 2452
rect 18285 2421 18294 2443
rect 18320 2421 18327 2443
rect 18552 2470 18663 2487
rect 18552 2450 18559 2470
rect 18578 2450 18636 2470
rect 18655 2450 18663 2470
rect 18552 2428 18663 2450
rect 18837 2448 18871 2654
rect 19284 2634 19316 2662
rect 18904 2626 19316 2634
rect 18904 2600 18910 2626
rect 18936 2600 19316 2626
rect 18904 2598 19316 2600
rect 18906 2597 18946 2598
rect 19284 2533 19316 2598
rect 19284 2513 19288 2533
rect 19309 2513 19316 2533
rect 19284 2506 19316 2513
rect 18837 2440 18872 2448
rect 18285 2411 18327 2421
rect 18837 2420 18845 2440
rect 18865 2420 18872 2440
rect 18837 2415 18872 2420
rect 19491 2435 19601 2450
rect 19491 2432 19568 2435
rect 18285 2410 18326 2411
rect 17919 2376 17954 2377
rect 17898 2369 17954 2376
rect 17898 2349 17927 2369
rect 17947 2349 17954 2369
rect 17898 2344 17954 2349
rect 18345 2372 18377 2379
rect 18345 2352 18351 2372
rect 18372 2352 18377 2372
rect 18837 2363 18871 2415
rect 19491 2405 19494 2432
rect 19523 2408 19568 2432
rect 19597 2408 19601 2435
rect 19523 2405 19601 2408
rect 19491 2391 19601 2405
rect 19787 2435 19829 2445
rect 19787 2416 19795 2435
rect 19820 2416 19829 2435
rect 19787 2363 19829 2416
rect 17898 2138 17932 2344
rect 18345 2324 18377 2352
rect 18835 2337 19831 2363
rect 17965 2316 18377 2324
rect 17965 2290 17971 2316
rect 17997 2290 18377 2316
rect 17965 2288 18377 2290
rect 17967 2287 18007 2288
rect 18127 2252 18166 2267
rect 18127 2211 18138 2252
rect 18159 2211 18166 2252
rect 17897 2130 17933 2138
rect 17897 2110 17906 2130
rect 17926 2110 17933 2130
rect 17897 2109 17933 2110
rect 17897 2098 17931 2109
rect 17787 2068 17824 2076
rect 17077 2046 17284 2048
rect 17077 1892 17121 2046
rect 17787 2034 18031 2068
rect 16942 1835 16950 1852
rect 16970 1835 16980 1852
rect 16942 1829 16980 1835
rect 16300 1789 16361 1791
rect 15998 1760 16361 1789
rect 16873 1763 16905 1770
rect 15998 1758 16300 1760
rect 13778 1742 14777 1745
rect 16873 1743 16880 1763
rect 16901 1743 16905 1763
rect 13778 1740 13813 1742
rect 12769 1736 13181 1738
rect 12771 1735 12811 1736
rect 13149 1671 13181 1736
rect 16873 1678 16905 1743
rect 17083 1756 17121 1892
rect 17779 1865 17814 1866
rect 17320 1861 17351 1862
rect 17317 1856 17351 1861
rect 17317 1836 17324 1856
rect 17344 1836 17351 1856
rect 17317 1828 17351 1836
rect 17083 1718 17089 1756
rect 17112 1718 17121 1756
rect 17083 1708 17121 1718
rect 17318 1770 17351 1828
rect 17758 1858 17814 1865
rect 17758 1838 17787 1858
rect 17807 1838 17814 1858
rect 17758 1833 17814 1838
rect 17989 1863 18031 2034
rect 18127 1938 18166 2211
rect 18345 2223 18377 2288
rect 18345 2203 18349 2223
rect 18370 2203 18377 2223
rect 18345 2196 18377 2203
rect 18763 2230 18821 2231
rect 18763 2211 19100 2230
rect 19490 2226 19601 2243
rect 18763 2198 19101 2211
rect 18267 2134 18320 2137
rect 18267 2117 18279 2134
rect 18311 2117 18320 2134
rect 18267 2109 18320 2117
rect 18266 2062 18320 2109
rect 18552 2125 18662 2140
rect 18552 2122 18629 2125
rect 18552 2095 18555 2122
rect 18584 2098 18629 2122
rect 18658 2098 18662 2125
rect 18584 2095 18662 2098
rect 18552 2081 18662 2095
rect 18763 2062 18800 2198
rect 19069 2181 19101 2198
rect 19490 2206 19497 2226
rect 19516 2206 19574 2226
rect 19593 2206 19601 2226
rect 19490 2184 19601 2206
rect 19069 2135 19100 2181
rect 18857 2132 18892 2133
rect 18836 2125 18892 2132
rect 18836 2105 18865 2125
rect 18885 2105 18892 2125
rect 18836 2100 18892 2105
rect 19069 2128 19108 2135
rect 19069 2108 19075 2128
rect 19100 2108 19108 2128
rect 19069 2102 19108 2108
rect 19283 2128 19315 2135
rect 19283 2108 19289 2128
rect 19310 2108 19315 2128
rect 18266 2027 18801 2062
rect 18266 2023 18319 2027
rect 18127 1911 18131 1938
rect 18162 1911 18166 1938
rect 18412 1959 18523 1976
rect 18412 1939 18419 1959
rect 18438 1939 18496 1959
rect 18515 1939 18523 1959
rect 18412 1917 18523 1939
rect 18127 1904 18166 1911
rect 18836 1894 18870 2100
rect 19283 2080 19315 2108
rect 18903 2072 19315 2080
rect 18903 2046 18909 2072
rect 18935 2046 19315 2072
rect 18903 2044 19315 2046
rect 18905 2043 18945 2044
rect 19283 1979 19315 2044
rect 19283 1959 19287 1979
rect 19308 1959 19315 1979
rect 19283 1952 19315 1959
rect 19786 1994 19834 1999
rect 19786 1965 19797 1994
rect 19826 1965 19834 1994
rect 18836 1893 18871 1894
rect 18834 1886 18871 1893
rect 17989 1842 17997 1863
rect 18024 1842 18031 1863
rect 17243 1678 17283 1679
rect 16873 1676 17285 1678
rect 16241 1672 16276 1674
rect 13149 1651 13153 1671
rect 13174 1651 13181 1671
rect 15277 1669 16276 1672
rect 13754 1654 14056 1656
rect 13149 1644 13181 1651
rect 13693 1625 14056 1654
rect 13693 1623 13754 1625
rect 12702 1578 12737 1586
rect 12702 1558 12710 1578
rect 12730 1558 12737 1578
rect 12702 1553 12737 1558
rect 13074 1579 13112 1585
rect 13074 1562 13084 1579
rect 13104 1562 13112 1579
rect 12702 1552 12734 1553
rect 12240 1548 12275 1549
rect 11183 1521 11220 1528
rect 11183 1520 11218 1521
rect 10220 1420 10228 1449
rect 10257 1420 10268 1449
rect 10220 1415 10268 1420
rect 10739 1455 10771 1462
rect 10739 1435 10746 1455
rect 10767 1435 10771 1455
rect 9254 1398 9286 1405
rect 10739 1370 10771 1435
rect 11109 1370 11149 1371
rect 10739 1368 11151 1370
rect 10739 1342 11119 1368
rect 11145 1342 11151 1368
rect 8807 1332 8842 1340
rect 8255 1303 8297 1313
rect 8807 1312 8815 1332
rect 8835 1312 8842 1332
rect 8807 1307 8842 1312
rect 9461 1327 9571 1342
rect 9461 1324 9538 1327
rect 8255 1302 8296 1303
rect 8099 1243 8107 1260
rect 8127 1243 8137 1260
rect 7125 1073 7160 1074
rect 6753 1039 6794 1040
rect 5511 1015 5588 1018
rect 5478 1000 5588 1015
rect 6207 1030 6242 1035
rect 6207 1010 6214 1030
rect 6234 1010 6242 1030
rect 6752 1029 6794 1039
rect 6207 1002 6242 1010
rect 3771 983 3806 984
rect 3750 976 3806 983
rect 3750 956 3779 976
rect 3799 956 3806 976
rect 3750 951 3806 956
rect 3983 979 4022 986
rect 3983 959 3989 979
rect 4014 959 4022 979
rect 3983 953 4022 959
rect 4197 979 4229 986
rect 4197 959 4203 979
rect 4224 959 4229 979
rect 1242 862 1733 891
rect 2811 878 3715 913
rect 2812 877 2846 878
rect 1130 722 1165 723
rect 421 651 532 671
rect 421 649 531 651
rect 421 629 429 649
rect 448 629 506 649
rect 525 629 531 649
rect 421 612 531 629
rect 912 640 954 721
rect 1242 642 1275 862
rect 1696 860 1733 862
rect 3750 745 3784 951
rect 4197 931 4229 959
rect 3817 923 4229 931
rect 3817 897 3823 923
rect 3849 897 4229 923
rect 3817 895 4229 897
rect 3819 894 3859 895
rect 4197 830 4229 895
rect 5763 937 5795 944
rect 5763 917 5770 937
rect 5791 917 5795 937
rect 5763 852 5795 917
rect 6133 852 6173 853
rect 5763 850 6175 852
rect 4197 810 4201 830
rect 4222 810 4229 830
rect 4197 803 4229 810
rect 4700 845 4748 850
rect 4700 816 4711 845
rect 4740 816 4748 845
rect 3750 744 3785 745
rect 1214 640 1275 642
rect 912 611 1275 640
rect 3748 737 3785 744
rect 3748 717 3758 737
rect 3778 717 3785 737
rect 3748 712 3785 717
rect 4404 732 4514 747
rect 4404 729 4481 732
rect 3748 661 3783 712
rect 4404 702 4407 729
rect 4436 705 4481 729
rect 4510 705 4514 732
rect 4436 702 4514 705
rect 4404 688 4514 702
rect 4700 661 4748 816
rect 5763 824 6143 850
rect 6169 824 6175 850
rect 5763 816 6175 824
rect 5763 788 5795 816
rect 6208 796 6242 1002
rect 6416 1000 6527 1022
rect 6416 980 6424 1000
rect 6443 980 6501 1000
rect 6520 980 6527 1000
rect 6416 963 6527 980
rect 6752 1007 6759 1029
rect 6785 1007 6794 1029
rect 6752 998 6794 1007
rect 7868 1030 7902 1236
rect 8099 1233 8137 1243
rect 8315 1264 8347 1271
rect 8315 1244 8321 1264
rect 8342 1244 8347 1264
rect 8807 1255 8841 1307
rect 9461 1297 9464 1324
rect 9493 1300 9538 1324
rect 9567 1300 9571 1327
rect 9493 1297 9571 1300
rect 9461 1283 9571 1297
rect 9757 1327 9799 1337
rect 9757 1308 9765 1327
rect 9790 1308 9799 1327
rect 9757 1255 9799 1308
rect 10739 1334 11151 1342
rect 10739 1306 10771 1334
rect 11184 1314 11218 1520
rect 11888 1503 11927 1510
rect 11531 1475 11642 1497
rect 11531 1455 11539 1475
rect 11558 1455 11616 1475
rect 11635 1455 11642 1475
rect 11531 1438 11642 1455
rect 11888 1476 11892 1503
rect 11923 1476 11927 1503
rect 11735 1387 11788 1391
rect 11253 1352 11788 1387
rect 10739 1286 10744 1306
rect 10765 1286 10771 1306
rect 10739 1279 10771 1286
rect 10946 1306 10985 1312
rect 10946 1286 10954 1306
rect 10979 1286 10985 1306
rect 10946 1279 10985 1286
rect 11162 1309 11218 1314
rect 11162 1289 11169 1309
rect 11189 1289 11218 1309
rect 11162 1282 11218 1289
rect 11162 1281 11197 1282
rect 8315 1216 8347 1244
rect 8805 1229 9801 1255
rect 10954 1233 10985 1279
rect 7935 1208 8347 1216
rect 7935 1182 7941 1208
rect 7967 1182 8347 1208
rect 7935 1180 8347 1182
rect 7937 1179 7977 1180
rect 8315 1115 8347 1180
rect 10453 1208 10564 1230
rect 10453 1188 10461 1208
rect 10480 1188 10538 1208
rect 10557 1188 10564 1208
rect 10953 1216 10985 1233
rect 11254 1216 11291 1352
rect 11392 1319 11502 1333
rect 11392 1316 11470 1319
rect 11392 1289 11396 1316
rect 11425 1292 11470 1316
rect 11499 1292 11502 1319
rect 11425 1289 11502 1292
rect 11392 1274 11502 1289
rect 11734 1305 11788 1352
rect 11734 1297 11787 1305
rect 11734 1280 11743 1297
rect 11775 1280 11787 1297
rect 11734 1277 11787 1280
rect 10953 1203 11291 1216
rect 10453 1171 10564 1188
rect 10954 1184 11291 1203
rect 11233 1183 11291 1184
rect 11677 1211 11709 1218
rect 11677 1191 11684 1211
rect 11705 1191 11709 1211
rect 8315 1095 8319 1115
rect 8340 1095 8347 1115
rect 8315 1088 8347 1095
rect 8733 1122 8791 1123
rect 8733 1103 9070 1122
rect 9460 1118 9571 1135
rect 8733 1090 9071 1103
rect 7868 1022 7903 1030
rect 7868 1002 7876 1022
rect 7896 1002 7903 1022
rect 5969 793 6012 795
rect 5763 768 5768 788
rect 5789 768 5795 788
rect 5763 761 5795 768
rect 5968 786 6012 793
rect 5968 766 5978 786
rect 6001 766 6012 786
rect 5968 762 6012 766
rect 6186 791 6242 796
rect 6186 771 6193 791
rect 6213 771 6242 791
rect 6186 764 6242 771
rect 6298 932 6331 933
rect 6752 932 6789 998
rect 7868 997 7903 1002
rect 8522 1017 8632 1032
rect 8522 1014 8599 1017
rect 7868 954 7902 997
rect 8522 987 8525 1014
rect 8554 990 8599 1014
rect 8628 990 8632 1017
rect 8554 987 8632 990
rect 8522 973 8632 987
rect 8733 954 8770 1090
rect 9039 1073 9071 1090
rect 9460 1098 9467 1118
rect 9486 1098 9544 1118
rect 9563 1098 9571 1118
rect 9460 1076 9571 1098
rect 11677 1126 11709 1191
rect 11888 1203 11927 1476
rect 12123 1305 12157 1316
rect 12121 1304 12157 1305
rect 12121 1284 12128 1304
rect 12148 1284 12157 1304
rect 12121 1276 12157 1284
rect 11888 1162 11895 1203
rect 11916 1162 11927 1203
rect 11888 1147 11927 1162
rect 12047 1126 12087 1127
rect 11677 1124 12089 1126
rect 11677 1098 12057 1124
rect 12083 1098 12089 1124
rect 11677 1090 12089 1098
rect 9039 1027 9070 1073
rect 10223 1051 11219 1077
rect 11677 1062 11709 1090
rect 12122 1070 12156 1276
rect 12864 1232 12899 1233
rect 8827 1024 8862 1025
rect 8806 1017 8862 1024
rect 8806 997 8835 1017
rect 8855 997 8862 1017
rect 8806 992 8862 997
rect 9039 1020 9078 1027
rect 9039 1000 9045 1020
rect 9070 1000 9078 1020
rect 9039 994 9078 1000
rect 9253 1020 9285 1027
rect 9253 1000 9259 1020
rect 9280 1000 9285 1020
rect 6298 903 6789 932
rect 7867 919 8771 954
rect 7868 918 7902 919
rect 6186 763 6221 764
rect 3748 637 4748 661
rect 5477 692 5588 712
rect 5477 690 5587 692
rect 5477 670 5485 690
rect 5504 670 5562 690
rect 5581 670 5587 690
rect 5477 653 5587 670
rect 5968 681 6010 762
rect 6298 683 6331 903
rect 6752 901 6789 903
rect 8806 786 8840 992
rect 9253 972 9285 1000
rect 8873 964 9285 972
rect 10225 998 10267 1051
rect 10225 979 10234 998
rect 10259 979 10267 998
rect 10225 969 10267 979
rect 10453 1009 10563 1023
rect 10453 1006 10531 1009
rect 10453 979 10457 1006
rect 10486 982 10531 1006
rect 10560 982 10563 1009
rect 11183 999 11217 1051
rect 11677 1042 11682 1062
rect 11703 1042 11709 1062
rect 11677 1035 11709 1042
rect 12100 1065 12156 1070
rect 12100 1045 12107 1065
rect 12127 1045 12156 1065
rect 12100 1038 12156 1045
rect 12843 1225 12899 1232
rect 12843 1205 12872 1225
rect 12892 1205 12899 1225
rect 12843 1200 12899 1205
rect 13074 1224 13112 1562
rect 13356 1573 13466 1588
rect 13356 1570 13433 1573
rect 13356 1543 13359 1570
rect 13388 1546 13433 1570
rect 13462 1546 13466 1573
rect 13388 1543 13466 1546
rect 13356 1529 13466 1543
rect 13235 1403 13272 1405
rect 13693 1403 13726 1623
rect 14014 1544 14056 1625
rect 14436 1636 14547 1653
rect 14436 1616 14443 1636
rect 14462 1616 14520 1636
rect 14539 1616 14547 1636
rect 14436 1594 14547 1616
rect 15276 1645 16276 1669
rect 13803 1542 13838 1543
rect 13235 1374 13726 1403
rect 13235 1308 13272 1374
rect 13693 1373 13726 1374
rect 13782 1535 13838 1542
rect 13782 1515 13811 1535
rect 13831 1515 13838 1535
rect 13782 1510 13838 1515
rect 14012 1540 14056 1544
rect 14012 1520 14023 1540
rect 14046 1520 14056 1540
rect 14012 1513 14056 1520
rect 14229 1538 14261 1545
rect 14229 1518 14235 1538
rect 14256 1518 14261 1538
rect 14012 1511 14055 1513
rect 13230 1299 13272 1308
rect 13230 1277 13239 1299
rect 13265 1277 13272 1299
rect 13497 1326 13608 1343
rect 13497 1306 13504 1326
rect 13523 1306 13581 1326
rect 13600 1306 13608 1326
rect 13497 1284 13608 1306
rect 13782 1304 13816 1510
rect 14229 1490 14261 1518
rect 13849 1482 14261 1490
rect 13849 1456 13855 1482
rect 13881 1456 14261 1482
rect 15276 1490 15324 1645
rect 15510 1604 15620 1618
rect 15510 1601 15588 1604
rect 15510 1574 15514 1601
rect 15543 1577 15588 1601
rect 15617 1577 15620 1604
rect 16241 1594 16276 1645
rect 15543 1574 15620 1577
rect 15510 1559 15620 1574
rect 16239 1589 16276 1594
rect 16239 1569 16246 1589
rect 16266 1569 16276 1589
rect 16873 1650 17253 1676
rect 17279 1650 17285 1676
rect 16873 1642 17285 1650
rect 16873 1614 16905 1642
rect 17318 1622 17354 1770
rect 16873 1594 16878 1614
rect 16899 1594 16905 1614
rect 16873 1587 16905 1594
rect 17296 1617 17354 1622
rect 17296 1597 17303 1617
rect 17323 1597 17354 1617
rect 17296 1590 17354 1597
rect 17758 1627 17792 1833
rect 17989 1831 18031 1842
rect 18205 1861 18237 1868
rect 18205 1841 18211 1861
rect 18232 1841 18237 1861
rect 18205 1813 18237 1841
rect 17825 1805 18237 1813
rect 17825 1779 17831 1805
rect 17857 1779 18237 1805
rect 18834 1866 18844 1886
rect 18864 1866 18871 1886
rect 18834 1861 18871 1866
rect 19490 1881 19600 1896
rect 19490 1878 19567 1881
rect 18834 1810 18869 1861
rect 19490 1851 19493 1878
rect 19522 1854 19567 1878
rect 19596 1854 19600 1881
rect 19522 1851 19600 1854
rect 19490 1837 19600 1851
rect 19786 1810 19834 1965
rect 18834 1786 19834 1810
rect 18834 1783 19833 1786
rect 18834 1781 18869 1783
rect 17825 1777 18237 1779
rect 17827 1776 17867 1777
rect 18205 1712 18237 1777
rect 18205 1692 18209 1712
rect 18230 1692 18237 1712
rect 18810 1695 19112 1697
rect 18205 1685 18237 1692
rect 18749 1666 19112 1695
rect 18749 1664 18810 1666
rect 17758 1619 17793 1627
rect 17758 1599 17766 1619
rect 17786 1599 17793 1619
rect 17758 1594 17793 1599
rect 18130 1620 18168 1626
rect 18130 1603 18140 1620
rect 18160 1603 18168 1620
rect 17758 1593 17790 1594
rect 17296 1589 17331 1590
rect 16239 1562 16276 1569
rect 16239 1561 16274 1562
rect 15276 1461 15284 1490
rect 15313 1461 15324 1490
rect 15276 1456 15324 1461
rect 15795 1496 15827 1503
rect 15795 1476 15802 1496
rect 15823 1476 15827 1496
rect 13849 1454 14261 1456
rect 13851 1453 13891 1454
rect 14229 1389 14261 1454
rect 14229 1369 14233 1389
rect 14254 1369 14261 1389
rect 14229 1362 14261 1369
rect 15795 1411 15827 1476
rect 16165 1411 16205 1412
rect 15795 1409 16207 1411
rect 15795 1383 16175 1409
rect 16201 1383 16207 1409
rect 15795 1375 16207 1383
rect 15795 1347 15827 1375
rect 16240 1355 16274 1561
rect 16944 1544 16983 1551
rect 16587 1516 16698 1538
rect 16587 1496 16595 1516
rect 16614 1496 16672 1516
rect 16691 1496 16698 1516
rect 16587 1479 16698 1496
rect 16944 1517 16948 1544
rect 16979 1517 16983 1544
rect 16791 1428 16844 1432
rect 16309 1393 16844 1428
rect 15795 1327 15800 1347
rect 15821 1327 15827 1347
rect 15795 1320 15827 1327
rect 16002 1347 16041 1353
rect 16002 1327 16010 1347
rect 16035 1327 16041 1347
rect 16002 1320 16041 1327
rect 16218 1350 16274 1355
rect 16218 1330 16225 1350
rect 16245 1330 16274 1350
rect 16218 1323 16274 1330
rect 16218 1322 16253 1323
rect 13782 1296 13817 1304
rect 13230 1267 13272 1277
rect 13782 1276 13790 1296
rect 13810 1276 13817 1296
rect 13782 1271 13817 1276
rect 14436 1291 14546 1306
rect 14436 1288 14513 1291
rect 13230 1266 13271 1267
rect 13074 1207 13082 1224
rect 13102 1207 13112 1224
rect 12100 1037 12135 1038
rect 11728 1003 11769 1004
rect 10486 979 10563 982
rect 10453 964 10563 979
rect 11182 994 11217 999
rect 11182 974 11189 994
rect 11209 974 11217 994
rect 11727 993 11769 1003
rect 11182 966 11217 974
rect 8873 938 8879 964
rect 8905 938 9285 964
rect 8873 936 9285 938
rect 8875 935 8915 936
rect 9253 871 9285 936
rect 10738 901 10770 908
rect 9253 851 9257 871
rect 9278 851 9285 871
rect 9253 844 9285 851
rect 9756 886 9804 891
rect 9756 857 9767 886
rect 9796 857 9804 886
rect 8806 785 8841 786
rect 6270 681 6331 683
rect 5968 652 6331 681
rect 8804 778 8841 785
rect 8804 758 8814 778
rect 8834 758 8841 778
rect 8804 753 8841 758
rect 9460 773 9570 788
rect 9460 770 9537 773
rect 8804 702 8839 753
rect 9460 743 9463 770
rect 9492 746 9537 770
rect 9566 746 9570 773
rect 9492 743 9570 746
rect 9460 729 9570 743
rect 9756 702 9804 857
rect 10738 881 10745 901
rect 10766 881 10770 901
rect 10738 816 10770 881
rect 11108 816 11148 817
rect 10738 814 11150 816
rect 10738 788 11118 814
rect 11144 788 11150 814
rect 10738 780 11150 788
rect 10738 752 10770 780
rect 11183 760 11217 966
rect 11391 964 11502 986
rect 11391 944 11399 964
rect 11418 944 11476 964
rect 11495 944 11502 964
rect 11391 927 11502 944
rect 11727 971 11734 993
rect 11760 971 11769 993
rect 11727 962 11769 971
rect 12843 994 12877 1200
rect 13074 1197 13112 1207
rect 13290 1228 13322 1235
rect 13290 1208 13296 1228
rect 13317 1208 13322 1228
rect 13782 1219 13816 1271
rect 14436 1261 14439 1288
rect 14468 1264 14513 1288
rect 14542 1264 14546 1291
rect 14468 1261 14546 1264
rect 14436 1247 14546 1261
rect 14732 1291 14774 1301
rect 14732 1272 14740 1291
rect 14765 1272 14774 1291
rect 16010 1274 16041 1320
rect 14732 1219 14774 1272
rect 15509 1249 15620 1271
rect 15509 1229 15517 1249
rect 15536 1229 15594 1249
rect 15613 1229 15620 1249
rect 16009 1257 16041 1274
rect 16310 1257 16347 1393
rect 16448 1360 16558 1374
rect 16448 1357 16526 1360
rect 16448 1330 16452 1357
rect 16481 1333 16526 1357
rect 16555 1333 16558 1360
rect 16481 1330 16558 1333
rect 16448 1315 16558 1330
rect 16790 1346 16844 1393
rect 16790 1338 16843 1346
rect 16790 1321 16799 1338
rect 16831 1321 16843 1338
rect 16790 1318 16843 1321
rect 16009 1244 16347 1257
rect 13290 1180 13322 1208
rect 13780 1193 14776 1219
rect 15509 1212 15620 1229
rect 16010 1225 16347 1244
rect 16289 1224 16347 1225
rect 16733 1252 16765 1259
rect 16733 1232 16740 1252
rect 16761 1232 16765 1252
rect 12910 1172 13322 1180
rect 12910 1146 12916 1172
rect 12942 1146 13322 1172
rect 12910 1144 13322 1146
rect 12912 1143 12952 1144
rect 13290 1079 13322 1144
rect 16733 1167 16765 1232
rect 16944 1244 16983 1517
rect 17179 1346 17213 1357
rect 17177 1345 17213 1346
rect 17177 1325 17184 1345
rect 17204 1325 17213 1345
rect 17177 1317 17213 1325
rect 16944 1203 16951 1244
rect 16972 1203 16983 1244
rect 16944 1188 16983 1203
rect 17103 1167 17143 1168
rect 16733 1165 17145 1167
rect 16733 1139 17113 1165
rect 17139 1139 17145 1165
rect 16733 1131 17145 1139
rect 13290 1059 13294 1079
rect 13315 1059 13322 1079
rect 13290 1052 13322 1059
rect 13708 1086 13766 1087
rect 13708 1067 14045 1086
rect 14435 1082 14546 1099
rect 15279 1092 16275 1118
rect 16733 1103 16765 1131
rect 17178 1111 17212 1317
rect 17920 1273 17955 1274
rect 13708 1054 14046 1067
rect 12843 986 12878 994
rect 12843 966 12851 986
rect 12871 966 12878 986
rect 10944 757 10987 759
rect 10738 732 10743 752
rect 10764 732 10770 752
rect 10738 725 10770 732
rect 10943 750 10987 757
rect 10943 730 10953 750
rect 10976 730 10987 750
rect 10943 726 10987 730
rect 11161 755 11217 760
rect 11161 735 11168 755
rect 11188 735 11217 755
rect 11161 728 11217 735
rect 11273 896 11306 897
rect 11727 896 11764 962
rect 12843 961 12878 966
rect 13497 981 13607 996
rect 13497 978 13574 981
rect 12843 918 12877 961
rect 13497 951 13500 978
rect 13529 954 13574 978
rect 13603 954 13607 981
rect 13529 951 13607 954
rect 13497 937 13607 951
rect 13708 918 13745 1054
rect 14014 1037 14046 1054
rect 14435 1062 14442 1082
rect 14461 1062 14519 1082
rect 14538 1062 14546 1082
rect 14435 1040 14546 1062
rect 15281 1039 15323 1092
rect 14014 991 14045 1037
rect 15281 1020 15290 1039
rect 15315 1020 15323 1039
rect 15281 1010 15323 1020
rect 15509 1050 15619 1064
rect 15509 1047 15587 1050
rect 15509 1020 15513 1047
rect 15542 1023 15587 1047
rect 15616 1023 15619 1050
rect 16239 1040 16273 1092
rect 16733 1083 16738 1103
rect 16759 1083 16765 1103
rect 16733 1076 16765 1083
rect 17156 1106 17212 1111
rect 17156 1086 17163 1106
rect 17183 1086 17212 1106
rect 17156 1079 17212 1086
rect 17899 1266 17955 1273
rect 17899 1246 17928 1266
rect 17948 1246 17955 1266
rect 17899 1241 17955 1246
rect 18130 1265 18168 1603
rect 18412 1614 18522 1629
rect 18412 1611 18489 1614
rect 18412 1584 18415 1611
rect 18444 1587 18489 1611
rect 18518 1587 18522 1614
rect 18444 1584 18522 1587
rect 18412 1570 18522 1584
rect 18291 1444 18328 1446
rect 18749 1444 18782 1664
rect 19070 1585 19112 1666
rect 19492 1677 19603 1694
rect 19492 1657 19499 1677
rect 19518 1657 19576 1677
rect 19595 1657 19603 1677
rect 19492 1635 19603 1657
rect 18859 1583 18894 1584
rect 18291 1415 18782 1444
rect 18291 1349 18328 1415
rect 18749 1414 18782 1415
rect 18838 1576 18894 1583
rect 18838 1556 18867 1576
rect 18887 1556 18894 1576
rect 18838 1551 18894 1556
rect 19068 1581 19112 1585
rect 19068 1561 19079 1581
rect 19102 1561 19112 1581
rect 19068 1554 19112 1561
rect 19285 1579 19317 1586
rect 19285 1559 19291 1579
rect 19312 1559 19317 1579
rect 19068 1552 19111 1554
rect 18286 1340 18328 1349
rect 18286 1318 18295 1340
rect 18321 1318 18328 1340
rect 18553 1367 18664 1384
rect 18553 1347 18560 1367
rect 18579 1347 18637 1367
rect 18656 1347 18664 1367
rect 18553 1325 18664 1347
rect 18838 1345 18872 1551
rect 19285 1531 19317 1559
rect 18905 1523 19317 1531
rect 18905 1497 18911 1523
rect 18937 1497 19317 1523
rect 18905 1495 19317 1497
rect 18907 1494 18947 1495
rect 19285 1430 19317 1495
rect 19285 1410 19289 1430
rect 19310 1410 19317 1430
rect 19285 1403 19317 1410
rect 18838 1337 18873 1345
rect 18286 1308 18328 1318
rect 18838 1317 18846 1337
rect 18866 1317 18873 1337
rect 18838 1312 18873 1317
rect 19492 1332 19602 1347
rect 19492 1329 19569 1332
rect 18286 1307 18327 1308
rect 18130 1248 18138 1265
rect 18158 1248 18168 1265
rect 17156 1078 17191 1079
rect 16784 1044 16825 1045
rect 15542 1020 15619 1023
rect 15509 1005 15619 1020
rect 16238 1035 16273 1040
rect 16238 1015 16245 1035
rect 16265 1015 16273 1035
rect 16783 1034 16825 1044
rect 16238 1007 16273 1015
rect 13802 988 13837 989
rect 13781 981 13837 988
rect 13781 961 13810 981
rect 13830 961 13837 981
rect 13781 956 13837 961
rect 14014 984 14053 991
rect 14014 964 14020 984
rect 14045 964 14053 984
rect 14014 958 14053 964
rect 14228 984 14260 991
rect 14228 964 14234 984
rect 14255 964 14260 984
rect 11273 867 11764 896
rect 12842 883 13746 918
rect 12843 882 12877 883
rect 11161 727 11196 728
rect 8804 678 9804 702
rect 8804 675 9803 678
rect 8804 673 8839 675
rect 10452 656 10563 676
rect 10452 654 10562 656
rect 5968 650 6270 652
rect 3748 634 4747 637
rect 10452 634 10460 654
rect 10479 634 10537 654
rect 10556 634 10562 654
rect 3748 632 3783 634
rect 5774 621 5853 625
rect 5774 612 9885 621
rect 10452 617 10562 634
rect 10943 645 10985 726
rect 11273 647 11306 867
rect 11727 865 11764 867
rect 13781 750 13815 956
rect 14228 936 14260 964
rect 13848 928 14260 936
rect 13848 902 13854 928
rect 13880 902 14260 928
rect 13848 900 14260 902
rect 13850 899 13890 900
rect 14228 835 14260 900
rect 15794 942 15826 949
rect 15794 922 15801 942
rect 15822 922 15826 942
rect 15794 857 15826 922
rect 16164 857 16204 858
rect 15794 855 16206 857
rect 14228 815 14232 835
rect 14253 815 14260 835
rect 14228 808 14260 815
rect 14731 850 14779 855
rect 14731 821 14742 850
rect 14771 821 14779 850
rect 13781 749 13816 750
rect 11245 645 11306 647
rect 10943 616 11306 645
rect 13779 742 13816 749
rect 13779 722 13789 742
rect 13809 722 13816 742
rect 13779 717 13816 722
rect 14435 737 14545 752
rect 14435 734 14512 737
rect 13779 666 13814 717
rect 14435 707 14438 734
rect 14467 710 14512 734
rect 14541 710 14545 737
rect 14467 707 14545 710
rect 14435 693 14545 707
rect 14731 666 14779 821
rect 15794 829 16174 855
rect 16200 829 16206 855
rect 15794 821 16206 829
rect 15794 793 15826 821
rect 16239 801 16273 1007
rect 16447 1005 16558 1027
rect 16447 985 16455 1005
rect 16474 985 16532 1005
rect 16551 985 16558 1005
rect 16447 968 16558 985
rect 16783 1012 16790 1034
rect 16816 1012 16825 1034
rect 16783 1003 16825 1012
rect 17899 1035 17933 1241
rect 18130 1238 18168 1248
rect 18346 1269 18378 1276
rect 18346 1249 18352 1269
rect 18373 1249 18378 1269
rect 18838 1260 18872 1312
rect 19492 1302 19495 1329
rect 19524 1305 19569 1329
rect 19598 1305 19602 1332
rect 19524 1302 19602 1305
rect 19492 1288 19602 1302
rect 19788 1332 19830 1342
rect 19788 1313 19796 1332
rect 19821 1313 19830 1332
rect 19788 1260 19830 1313
rect 18346 1221 18378 1249
rect 18836 1234 19832 1260
rect 17966 1213 18378 1221
rect 17966 1187 17972 1213
rect 17998 1187 18378 1213
rect 17966 1185 18378 1187
rect 17968 1184 18008 1185
rect 18346 1120 18378 1185
rect 18346 1100 18350 1120
rect 18371 1100 18378 1120
rect 18346 1093 18378 1100
rect 18764 1127 18822 1128
rect 18764 1108 19101 1127
rect 19491 1123 19602 1140
rect 18764 1095 19102 1108
rect 17899 1027 17934 1035
rect 17899 1007 17907 1027
rect 17927 1007 17934 1027
rect 16000 798 16043 800
rect 15794 773 15799 793
rect 15820 773 15826 793
rect 15794 766 15826 773
rect 15999 791 16043 798
rect 15999 771 16009 791
rect 16032 771 16043 791
rect 15999 767 16043 771
rect 16217 796 16273 801
rect 16217 776 16224 796
rect 16244 776 16273 796
rect 16217 769 16273 776
rect 16329 937 16362 938
rect 16783 937 16820 1003
rect 17899 1002 17934 1007
rect 18553 1022 18663 1037
rect 18553 1019 18630 1022
rect 17899 959 17933 1002
rect 18553 992 18556 1019
rect 18585 995 18630 1019
rect 18659 995 18663 1022
rect 18585 992 18663 995
rect 18553 978 18663 992
rect 18764 959 18801 1095
rect 19070 1078 19102 1095
rect 19491 1103 19498 1123
rect 19517 1103 19575 1123
rect 19594 1103 19602 1123
rect 19491 1081 19602 1103
rect 19070 1032 19101 1078
rect 18858 1029 18893 1030
rect 18837 1022 18893 1029
rect 18837 1002 18866 1022
rect 18886 1002 18893 1022
rect 18837 997 18893 1002
rect 19070 1025 19109 1032
rect 19070 1005 19076 1025
rect 19101 1005 19109 1025
rect 19070 999 19109 1005
rect 19284 1025 19316 1032
rect 19284 1005 19290 1025
rect 19311 1005 19316 1025
rect 16329 908 16820 937
rect 17898 924 18802 959
rect 17899 923 17933 924
rect 16217 768 16252 769
rect 13779 642 14779 666
rect 15508 697 15619 717
rect 15508 695 15618 697
rect 15508 675 15516 695
rect 15535 675 15593 695
rect 15612 675 15618 695
rect 15508 658 15618 675
rect 15999 686 16041 767
rect 16329 688 16362 908
rect 16783 906 16820 908
rect 18837 791 18871 997
rect 19284 977 19316 1005
rect 18904 969 19316 977
rect 18904 943 18910 969
rect 18936 943 19316 969
rect 18904 941 19316 943
rect 18906 940 18946 941
rect 19284 876 19316 941
rect 19284 856 19288 876
rect 19309 856 19316 876
rect 19284 849 19316 856
rect 19787 891 19835 896
rect 19787 862 19798 891
rect 19827 862 19835 891
rect 18837 790 18872 791
rect 16301 686 16362 688
rect 15999 657 16362 686
rect 18835 783 18872 790
rect 18835 763 18845 783
rect 18865 763 18872 783
rect 18835 758 18872 763
rect 19491 778 19601 793
rect 19491 775 19568 778
rect 18835 707 18870 758
rect 19491 748 19494 775
rect 19523 751 19568 775
rect 19597 751 19601 778
rect 19523 748 19601 751
rect 19491 734 19601 748
rect 19787 707 19835 862
rect 18835 683 19835 707
rect 18835 680 19834 683
rect 18835 678 18870 680
rect 15999 655 16301 657
rect 13779 639 14778 642
rect 13779 637 13814 639
rect 15805 626 15884 630
rect 15805 617 19916 626
rect 10943 614 11245 616
rect 912 609 1214 611
rect 5774 608 9848 612
rect 5774 587 5813 608
rect 5842 591 9848 608
rect 9877 591 9885 612
rect 5842 587 9885 591
rect 15805 613 19879 617
rect 15805 592 15844 613
rect 15873 596 19879 613
rect 19908 596 19916 617
rect 15873 592 19916 596
rect 718 580 797 584
rect 718 571 4829 580
rect 718 567 4792 571
rect 718 546 757 567
rect 786 550 4792 567
rect 4821 550 4829 571
rect 5774 579 9885 587
rect 10749 585 10828 589
rect 5774 568 5853 579
rect 10749 576 14860 585
rect 10749 572 14823 576
rect 786 546 4829 550
rect 10749 551 10788 572
rect 10817 555 14823 572
rect 14852 555 14860 576
rect 15805 584 19916 592
rect 15805 573 15884 584
rect 10817 551 14860 555
rect 718 538 4829 546
rect 718 527 797 538
rect 7440 529 7499 545
rect 2384 488 2443 504
rect 1669 445 1779 459
rect 1669 442 1747 445
rect 1669 415 1673 442
rect 1702 418 1747 442
rect 1776 418 1779 445
rect 1702 415 1779 418
rect 1669 400 1779 415
rect 2384 446 2403 488
rect 2435 446 2443 488
rect 2384 430 2443 446
rect 2384 410 2405 430
rect 2425 410 2443 430
rect 2384 405 2443 410
rect 2472 485 2532 505
rect 5351 494 5389 496
rect 2472 422 2484 485
rect 2515 422 2532 485
rect 4311 460 5391 494
rect 6725 486 6835 500
rect 6725 483 6803 486
rect 2472 407 2532 422
rect 2398 402 2433 405
rect 1954 337 1986 344
rect 1954 317 1961 337
rect 1982 317 1986 337
rect 1954 252 1986 317
rect 2324 252 2364 253
rect 1954 250 2366 252
rect 1954 224 2334 250
rect 2360 224 2366 250
rect 1954 216 2366 224
rect 1954 188 1986 216
rect 2399 196 2433 402
rect 1954 168 1959 188
rect 1980 168 1986 188
rect 1954 161 1986 168
rect 2154 187 2212 194
rect 2154 167 2165 187
rect 2199 167 2212 187
rect 1668 90 1779 112
rect 1668 70 1676 90
rect 1695 70 1753 90
rect 1772 70 1779 90
rect 1668 53 1779 70
rect 2154 94 2212 167
rect 2377 191 2433 196
rect 2377 171 2384 191
rect 2404 171 2433 191
rect 2377 164 2433 171
rect 2377 163 2412 164
rect 2472 130 2527 407
rect 2472 109 2486 130
rect 2513 109 2527 130
rect 2472 99 2527 109
rect 2154 83 2215 94
rect 4315 83 4367 460
rect 4619 425 4729 439
rect 4619 422 4697 425
rect 4619 395 4623 422
rect 4652 398 4697 422
rect 4726 398 4729 425
rect 5351 415 5389 460
rect 6725 456 6729 483
rect 6758 459 6803 483
rect 6832 459 6835 486
rect 6758 456 6835 459
rect 6725 441 6835 456
rect 7440 487 7459 529
rect 7491 487 7499 529
rect 7440 471 7499 487
rect 7440 451 7461 471
rect 7481 451 7499 471
rect 7440 446 7499 451
rect 7528 526 7588 546
rect 10749 543 14860 551
rect 10749 532 10828 543
rect 17471 534 17530 550
rect 7528 463 7540 526
rect 7571 463 7588 526
rect 7898 491 10266 494
rect 12415 493 12474 509
rect 7898 485 10321 491
rect 7528 448 7588 463
rect 7454 443 7489 446
rect 4652 395 4729 398
rect 4619 380 4729 395
rect 5348 410 5389 415
rect 5348 390 5355 410
rect 5375 390 5389 410
rect 5348 388 5389 390
rect 5348 382 5383 388
rect 4904 317 4936 324
rect 4904 297 4911 317
rect 4932 297 4936 317
rect 4904 232 4936 297
rect 5274 232 5314 233
rect 4904 230 5316 232
rect 4904 204 5284 230
rect 5310 204 5316 230
rect 4904 196 5316 204
rect 4904 168 4936 196
rect 4904 148 4909 168
rect 4930 148 4936 168
rect 4904 141 4936 148
rect 5099 167 5162 177
rect 5349 176 5383 382
rect 7010 378 7042 385
rect 7010 358 7017 378
rect 7038 358 7042 378
rect 7010 293 7042 358
rect 7380 293 7420 294
rect 7010 291 7422 293
rect 7010 265 7390 291
rect 7416 265 7422 291
rect 7010 257 7422 265
rect 7010 229 7042 257
rect 7455 237 7489 443
rect 7010 209 7015 229
rect 7036 209 7042 229
rect 7010 202 7042 209
rect 7210 228 7268 235
rect 7210 208 7221 228
rect 7255 208 7268 228
rect 5099 147 5109 167
rect 5150 147 5162 167
rect 2154 66 4367 83
rect 2155 42 4367 66
rect 4315 38 4367 42
rect 4618 70 4729 92
rect 4618 50 4626 70
rect 4645 50 4703 70
rect 4722 50 4729 70
rect 4618 33 4729 50
rect 5099 4 5162 147
rect 5327 171 5383 176
rect 5327 151 5334 171
rect 5354 151 5383 171
rect 5327 144 5383 151
rect 5327 143 5362 144
rect 6724 131 6835 153
rect 5413 111 5486 123
rect 5413 85 5422 111
rect 5481 85 5486 111
rect 6724 111 6732 131
rect 6751 111 6809 131
rect 6828 111 6835 131
rect 6724 94 6835 111
rect 5413 52 5486 85
rect 7210 76 7268 208
rect 7433 232 7489 237
rect 7433 212 7440 232
rect 7460 212 7489 232
rect 7433 205 7489 212
rect 7433 204 7468 205
rect 7528 171 7583 448
rect 7528 150 7542 171
rect 7569 150 7583 171
rect 7528 140 7583 150
rect 7893 419 10321 485
rect 7205 52 7270 76
rect 5100 -34 5161 4
rect 5406 0 7275 52
rect 7893 -26 7996 419
rect 9553 309 9663 323
rect 9553 306 9631 309
rect 9553 279 9557 306
rect 9586 282 9631 306
rect 9660 282 9663 309
rect 10283 299 10321 419
rect 11700 450 11810 464
rect 11700 447 11778 450
rect 11700 420 11704 447
rect 11733 423 11778 447
rect 11807 423 11810 450
rect 11733 420 11810 423
rect 11700 405 11810 420
rect 12415 451 12434 493
rect 12466 451 12474 493
rect 12415 435 12474 451
rect 12415 415 12436 435
rect 12456 415 12474 435
rect 12415 410 12474 415
rect 12503 490 12563 510
rect 15382 499 15420 501
rect 12503 427 12515 490
rect 12546 427 12563 490
rect 14342 465 15422 499
rect 16756 491 16866 505
rect 16756 488 16834 491
rect 12503 412 12563 427
rect 12429 407 12464 410
rect 9586 279 9663 282
rect 9553 264 9663 279
rect 10282 294 10321 299
rect 10282 274 10289 294
rect 10309 274 10321 294
rect 10282 270 10321 274
rect 11985 342 12017 349
rect 11985 322 11992 342
rect 12013 322 12017 342
rect 10282 266 10317 270
rect 9838 201 9870 208
rect 9838 181 9845 201
rect 9866 181 9870 201
rect 9838 116 9870 181
rect 10208 116 10248 117
rect 9838 114 10250 116
rect 9838 88 10218 114
rect 10244 88 10250 114
rect 9838 80 10250 88
rect 9838 52 9870 80
rect 10283 60 10317 266
rect 11985 257 12017 322
rect 12355 257 12395 258
rect 11985 255 12397 257
rect 11985 229 12365 255
rect 12391 229 12397 255
rect 11985 221 12397 229
rect 11985 193 12017 221
rect 12430 201 12464 407
rect 11985 173 11990 193
rect 12011 173 12017 193
rect 11985 166 12017 173
rect 12185 192 12243 199
rect 12185 172 12196 192
rect 12230 172 12243 192
rect 9838 32 9843 52
rect 9864 32 9870 52
rect 9838 25 9870 32
rect 10035 52 10100 58
rect 10035 28 10050 52
rect 10083 28 10100 52
rect 5564 -34 7996 -26
rect 5100 -78 7996 -34
rect 5564 -80 7996 -78
rect 7893 -87 7996 -80
rect 9552 -46 9663 -24
rect 9552 -66 9560 -46
rect 9579 -66 9637 -46
rect 9656 -66 9663 -46
rect 9552 -83 9663 -66
rect 10035 -190 10100 28
rect 10261 55 10317 60
rect 11699 95 11810 117
rect 11699 75 11707 95
rect 11726 75 11784 95
rect 11803 75 11810 95
rect 11699 58 11810 75
rect 12185 99 12243 172
rect 12408 196 12464 201
rect 12408 176 12415 196
rect 12435 176 12464 196
rect 12408 169 12464 176
rect 12408 168 12443 169
rect 12503 135 12558 412
rect 12503 114 12517 135
rect 12544 114 12558 135
rect 12503 104 12558 114
rect 12185 88 12246 99
rect 14346 88 14398 465
rect 14650 430 14760 444
rect 14650 427 14728 430
rect 14650 400 14654 427
rect 14683 403 14728 427
rect 14757 403 14760 430
rect 15382 420 15420 465
rect 16756 461 16760 488
rect 16789 464 16834 488
rect 16863 464 16866 491
rect 16789 461 16866 464
rect 16756 446 16866 461
rect 17471 492 17490 534
rect 17522 492 17530 534
rect 17471 476 17530 492
rect 17471 456 17492 476
rect 17512 456 17530 476
rect 17471 451 17530 456
rect 17559 531 17619 551
rect 17559 468 17571 531
rect 17602 468 17619 531
rect 17559 453 17619 468
rect 17485 448 17520 451
rect 14683 400 14760 403
rect 14650 385 14760 400
rect 15379 415 15420 420
rect 15379 395 15386 415
rect 15406 395 15420 415
rect 15379 393 15420 395
rect 15379 387 15414 393
rect 14935 322 14967 329
rect 14935 302 14942 322
rect 14963 302 14967 322
rect 14935 237 14967 302
rect 15305 237 15345 238
rect 14935 235 15347 237
rect 14935 209 15315 235
rect 15341 209 15347 235
rect 14935 201 15347 209
rect 14935 173 14967 201
rect 15380 181 15414 387
rect 17041 383 17073 390
rect 17041 363 17048 383
rect 17069 363 17073 383
rect 17041 298 17073 363
rect 17411 298 17451 299
rect 17041 296 17453 298
rect 17041 270 17421 296
rect 17447 270 17453 296
rect 17041 262 17453 270
rect 17041 234 17073 262
rect 17486 242 17520 448
rect 17041 214 17046 234
rect 17067 214 17073 234
rect 17041 207 17073 214
rect 17241 233 17299 240
rect 17241 213 17252 233
rect 17286 213 17299 233
rect 14935 153 14940 173
rect 14961 153 14967 173
rect 14935 146 14967 153
rect 15121 173 15192 180
rect 15121 149 15137 173
rect 15178 149 15192 173
rect 12185 71 14398 88
rect 10261 35 10268 55
rect 10288 35 10317 55
rect 12186 47 14398 71
rect 14346 43 14398 47
rect 14649 75 14760 97
rect 14649 55 14657 75
rect 14676 55 14734 75
rect 14753 55 14760 75
rect 14649 38 14760 55
rect 10261 28 10317 35
rect 10261 27 10296 28
rect 10273 -12 10333 -2
rect 10273 -42 10282 -12
rect 10323 -42 10333 -12
rect 10273 -52 10333 -42
rect 10280 -126 10333 -52
rect 10280 -127 10664 -126
rect 15121 -127 15192 149
rect 15358 176 15414 181
rect 15358 156 15365 176
rect 15385 156 15414 176
rect 15358 149 15414 156
rect 15358 148 15393 149
rect 16755 136 16866 158
rect 15444 116 15517 128
rect 15444 90 15453 116
rect 15512 90 15517 116
rect 16755 116 16763 136
rect 16782 116 16840 136
rect 16859 116 16866 136
rect 16755 99 16866 116
rect 15444 57 15517 90
rect 17241 81 17299 213
rect 17464 237 17520 242
rect 17464 217 17471 237
rect 17491 217 17520 237
rect 17464 210 17520 217
rect 17464 209 17499 210
rect 17559 176 17614 453
rect 17559 155 17573 176
rect 17600 155 17614 176
rect 17559 145 17614 155
rect 17236 57 17301 81
rect 15437 5 17306 57
rect 10280 -189 15192 -127
rect 10280 -193 10664 -189
<< via1 >>
rect 2485 5155 2516 5208
rect 7541 5196 7572 5249
rect 2405 4767 2436 4820
rect 12516 5160 12547 5213
rect 7461 4808 7492 4861
rect 17572 5201 17603 5254
rect 12436 4772 12467 4825
rect 17492 4813 17523 4866
rect 2403 446 2435 488
rect 2484 422 2515 485
rect 7459 487 7491 529
rect 7540 463 7571 526
rect 12434 451 12466 493
rect 12515 427 12546 490
rect 17490 492 17522 534
rect 17571 468 17602 531
<< metal2 >>
rect 7529 5249 7577 5268
rect 2473 5208 2521 5227
rect 2473 5155 2485 5208
rect 2516 5155 2521 5208
rect 2394 4820 2442 4835
rect 2394 4767 2405 4820
rect 2436 4767 2442 4820
rect 2394 504 2442 4767
rect 2473 505 2521 5155
rect 7529 5196 7541 5249
rect 7572 5196 7577 5249
rect 17560 5254 17608 5273
rect 7450 4861 7498 4876
rect 7450 4808 7461 4861
rect 7492 4808 7498 4861
rect 7450 545 7498 4808
rect 7529 546 7577 5196
rect 12504 5213 12552 5232
rect 12504 5160 12516 5213
rect 12547 5160 12552 5213
rect 12425 4825 12473 4840
rect 12425 4772 12436 4825
rect 12467 4772 12473 4825
rect 7440 529 7499 545
rect 2384 488 2443 504
rect 2384 446 2403 488
rect 2435 446 2443 488
rect 2384 405 2443 446
rect 2472 485 2532 505
rect 2472 422 2484 485
rect 2515 422 2532 485
rect 7440 487 7459 529
rect 7491 487 7499 529
rect 7440 446 7499 487
rect 7528 526 7588 546
rect 7528 463 7540 526
rect 7571 463 7588 526
rect 12425 509 12473 4772
rect 12504 510 12552 5160
rect 17560 5201 17572 5254
rect 17603 5201 17608 5254
rect 17481 4866 17529 4881
rect 17481 4813 17492 4866
rect 17523 4813 17529 4866
rect 17481 550 17529 4813
rect 17560 551 17608 5201
rect 17471 534 17530 550
rect 7528 448 7588 463
rect 12415 493 12474 509
rect 12415 451 12434 493
rect 12466 451 12474 493
rect 2472 407 2532 422
rect 12415 410 12474 451
rect 12503 490 12563 510
rect 12503 427 12515 490
rect 12546 427 12563 490
rect 17471 492 17490 534
rect 17522 492 17530 534
rect 17471 451 17530 492
rect 17559 531 17619 551
rect 17559 468 17571 531
rect 17602 468 17619 531
rect 17559 453 17619 468
rect 12503 412 12563 427
<< labels >>
rlabel locali 290 9060 312 9075 1 d0
rlabel metal1 459 9283 487 9288 1 vdd
rlabel metal1 456 8890 490 8896 1 gnd
rlabel locali 1227 8812 1255 8833 1 d1
rlabel metal1 1394 8646 1428 8652 1 gnd
rlabel metal1 1397 9039 1425 9044 1 vdd
rlabel locali 289 8506 311 8521 1 d0
rlabel metal1 458 8729 486 8734 1 vdd
rlabel metal1 455 8336 489 8342 1 gnd
rlabel locali 110 9345 138 9353 1 vref
rlabel locali 291 7957 313 7972 1 d0
rlabel metal1 460 8180 488 8185 1 vdd
rlabel metal1 457 7787 491 7793 1 gnd
rlabel locali 1228 7709 1256 7730 1 d1
rlabel metal1 1395 7543 1429 7549 1 gnd
rlabel metal1 1398 7936 1426 7941 1 vdd
rlabel locali 290 7403 312 7418 1 d0
rlabel metal1 459 7626 487 7631 1 vdd
rlabel metal1 456 7233 490 7239 1 gnd
rlabel metal1 1538 8447 1566 8452 1 vdd
rlabel metal1 1535 8054 1569 8060 1 gnd
rlabel locali 1366 8219 1387 8238 1 d2
rlabel locali 291 6854 313 6869 1 d0
rlabel metal1 460 7077 488 7082 1 vdd
rlabel metal1 457 6684 491 6690 1 gnd
rlabel locali 1228 6606 1256 6627 1 d1
rlabel metal1 1395 6440 1429 6446 1 gnd
rlabel metal1 1398 6833 1426 6838 1 vdd
rlabel locali 290 6300 312 6315 1 d0
rlabel metal1 459 6523 487 6528 1 vdd
rlabel metal1 456 6130 490 6136 1 gnd
rlabel locali 292 5751 314 5766 1 d0
rlabel metal1 461 5974 489 5979 1 vdd
rlabel metal1 458 5581 492 5587 1 gnd
rlabel locali 1229 5503 1257 5524 1 d1
rlabel metal1 1396 5337 1430 5343 1 gnd
rlabel metal1 1399 5730 1427 5735 1 vdd
rlabel locali 291 5197 313 5212 1 d0
rlabel metal1 460 5420 488 5425 1 vdd
rlabel metal1 457 5027 491 5033 1 gnd
rlabel metal1 1539 6241 1567 6246 1 vdd
rlabel metal1 1536 5848 1570 5854 1 gnd
rlabel locali 1367 6013 1388 6032 1 d2
rlabel metal1 1508 7357 1536 7362 1 vdd
rlabel metal1 1505 6964 1539 6970 1 gnd
rlabel locali 1338 7133 1364 7150 1 d3
rlabel locali 1340 2721 1366 2738 1 d3
rlabel metal1 1507 2552 1541 2558 1 gnd
rlabel metal1 1510 2945 1538 2950 1 vdd
rlabel locali 1369 1601 1390 1620 1 d2
rlabel metal1 1538 1436 1572 1442 1 gnd
rlabel metal1 1541 1829 1569 1834 1 vdd
rlabel metal1 459 615 493 621 1 gnd
rlabel metal1 462 1008 490 1013 1 vdd
rlabel locali 293 785 315 800 1 d0
rlabel metal1 1401 1318 1429 1323 1 vdd
rlabel metal1 1398 925 1432 931 1 gnd
rlabel locali 1231 1091 1259 1112 1 d1
rlabel metal1 460 1169 494 1175 1 gnd
rlabel metal1 463 1562 491 1567 1 vdd
rlabel locali 294 1339 316 1354 1 d0
rlabel metal1 458 1718 492 1724 1 gnd
rlabel metal1 461 2111 489 2116 1 vdd
rlabel locali 292 1888 314 1903 1 d0
rlabel metal1 1400 2421 1428 2426 1 vdd
rlabel metal1 1397 2028 1431 2034 1 gnd
rlabel locali 1230 2194 1258 2215 1 d1
rlabel metal1 459 2272 493 2278 1 gnd
rlabel metal1 462 2665 490 2670 1 vdd
rlabel locali 293 2442 315 2457 1 d0
rlabel locali 1368 3807 1389 3826 1 d2
rlabel metal1 1537 3642 1571 3648 1 gnd
rlabel metal1 1540 4035 1568 4040 1 vdd
rlabel metal1 458 2821 492 2827 1 gnd
rlabel metal1 461 3214 489 3219 1 vdd
rlabel locali 292 2991 314 3006 1 d0
rlabel metal1 1400 3524 1428 3529 1 vdd
rlabel metal1 1397 3131 1431 3137 1 gnd
rlabel locali 1230 3297 1258 3318 1 d1
rlabel metal1 459 3375 493 3381 1 gnd
rlabel metal1 462 3768 490 3773 1 vdd
rlabel locali 293 3545 315 3560 1 d0
rlabel metal1 457 3924 491 3930 1 gnd
rlabel metal1 460 4317 488 4322 1 vdd
rlabel locali 291 4094 313 4109 1 d0
rlabel metal1 1399 4627 1427 4632 1 vdd
rlabel metal1 1396 4234 1430 4240 1 gnd
rlabel locali 1229 4400 1257 4421 1 d1
rlabel metal1 458 4478 492 4484 1 gnd
rlabel metal1 461 4871 489 4876 1 vdd
rlabel locali 292 4648 314 4663 1 d0
rlabel metal1 1508 5157 1536 5162 1 vdd
rlabel metal1 1505 4764 1539 4770 1 gnd
rlabel locali 1332 4926 1367 4952 1 d4
rlabel locali 4621 906 4643 921 5 d0
rlabel metal1 4446 693 4474 698 5 vdd
rlabel metal1 4443 1085 4477 1091 5 gnd
rlabel locali 3678 1148 3706 1169 5 d1
rlabel metal1 3505 1329 3539 1335 5 gnd
rlabel metal1 3508 937 3536 942 5 vdd
rlabel locali 4622 1460 4644 1475 5 d0
rlabel metal1 4447 1247 4475 1252 5 vdd
rlabel metal1 4444 1639 4478 1645 5 gnd
rlabel locali 4620 2009 4642 2024 5 d0
rlabel metal1 4445 1796 4473 1801 5 vdd
rlabel metal1 4442 2188 4476 2194 5 gnd
rlabel locali 3677 2251 3705 2272 5 d1
rlabel metal1 3504 2432 3538 2438 5 gnd
rlabel metal1 3507 2040 3535 2045 5 vdd
rlabel locali 4621 2563 4643 2578 5 d0
rlabel metal1 4446 2350 4474 2355 5 vdd
rlabel metal1 4443 2742 4477 2748 5 gnd
rlabel metal1 3367 1529 3395 1534 5 vdd
rlabel metal1 3364 1921 3398 1927 5 gnd
rlabel locali 3546 1743 3567 1762 5 d2
rlabel locali 4620 3112 4642 3127 5 d0
rlabel metal1 4445 2899 4473 2904 5 vdd
rlabel metal1 4442 3291 4476 3297 5 gnd
rlabel locali 3677 3354 3705 3375 5 d1
rlabel metal1 3504 3535 3538 3541 5 gnd
rlabel metal1 3507 3143 3535 3148 5 vdd
rlabel locali 4621 3666 4643 3681 5 d0
rlabel metal1 4446 3453 4474 3458 5 vdd
rlabel metal1 4443 3845 4477 3851 5 gnd
rlabel locali 4619 4215 4641 4230 5 d0
rlabel metal1 4444 4002 4472 4007 5 vdd
rlabel metal1 4441 4394 4475 4400 5 gnd
rlabel locali 3676 4457 3704 4478 5 d1
rlabel metal1 3503 4638 3537 4644 5 gnd
rlabel metal1 3506 4246 3534 4251 5 vdd
rlabel locali 4620 4769 4642 4784 5 d0
rlabel metal1 4445 4556 4473 4561 5 vdd
rlabel metal1 4442 4948 4476 4954 5 gnd
rlabel metal1 3366 3735 3394 3740 5 vdd
rlabel metal1 3363 4127 3397 4133 5 gnd
rlabel locali 3545 3949 3566 3968 5 d2
rlabel metal1 3397 2619 3425 2624 5 vdd
rlabel metal1 3394 3011 3428 3017 5 gnd
rlabel locali 3569 2831 3595 2848 5 d3
rlabel locali 3567 7243 3593 7260 5 d3
rlabel metal1 3392 7423 3426 7429 5 gnd
rlabel metal1 3395 7031 3423 7036 5 vdd
rlabel locali 3543 8361 3564 8380 5 d2
rlabel metal1 3361 8539 3395 8545 5 gnd
rlabel metal1 3364 8147 3392 8152 5 vdd
rlabel metal1 4440 9360 4474 9366 5 gnd
rlabel metal1 4443 8968 4471 8973 5 vdd
rlabel locali 4618 9181 4640 9196 5 d0
rlabel metal1 3504 8658 3532 8663 5 vdd
rlabel metal1 3501 9050 3535 9056 5 gnd
rlabel locali 3674 8869 3702 8890 5 d1
rlabel metal1 4439 8806 4473 8812 5 gnd
rlabel metal1 4442 8414 4470 8419 5 vdd
rlabel locali 4617 8627 4639 8642 5 d0
rlabel metal1 4441 8257 4475 8263 5 gnd
rlabel metal1 4444 7865 4472 7870 5 vdd
rlabel locali 4619 8078 4641 8093 5 d0
rlabel metal1 3505 7555 3533 7560 5 vdd
rlabel metal1 3502 7947 3536 7953 5 gnd
rlabel locali 3675 7766 3703 7787 5 d1
rlabel metal1 4440 7703 4474 7709 5 gnd
rlabel metal1 4443 7311 4471 7316 5 vdd
rlabel locali 4618 7524 4640 7539 5 d0
rlabel locali 3544 6155 3565 6174 5 d2
rlabel metal1 3362 6333 3396 6339 5 gnd
rlabel metal1 3365 5941 3393 5946 5 vdd
rlabel metal1 4441 7154 4475 7160 5 gnd
rlabel metal1 4444 6762 4472 6767 5 vdd
rlabel locali 4619 6975 4641 6990 5 d0
rlabel metal1 3505 6452 3533 6457 5 vdd
rlabel metal1 3502 6844 3536 6850 5 gnd
rlabel locali 3675 6663 3703 6684 5 d1
rlabel metal1 4440 6600 4474 6606 5 gnd
rlabel metal1 4443 6208 4471 6213 5 vdd
rlabel locali 4618 6421 4640 6436 5 d0
rlabel metal1 4442 6051 4476 6057 5 gnd
rlabel metal1 4445 5659 4473 5664 5 vdd
rlabel locali 4620 5872 4642 5887 5 d0
rlabel metal1 3506 5349 3534 5354 5 vdd
rlabel metal1 3503 5741 3537 5747 5 gnd
rlabel locali 3676 5560 3704 5581 5 d1
rlabel metal1 4441 5497 4475 5503 5 gnd
rlabel metal1 4444 5105 4472 5110 5 vdd
rlabel locali 4619 5318 4641 5333 5 d0
rlabel metal1 3397 4819 3425 4824 5 vdd
rlabel metal1 3394 5211 3428 5217 5 gnd
rlabel locali 3566 5029 3601 5055 5 d4
rlabel metal1 1709 449 1737 454 1 vdd
rlabel metal1 1706 56 1740 62 1 gnd
rlabel locali 1535 220 1563 242 1 d5
rlabel locali 5346 9101 5368 9116 1 d0
rlabel metal1 5515 9324 5543 9329 1 vdd
rlabel metal1 5512 8931 5546 8937 1 gnd
rlabel locali 6283 8853 6311 8874 1 d1
rlabel metal1 6450 8687 6484 8693 1 gnd
rlabel metal1 6453 9080 6481 9085 1 vdd
rlabel locali 5345 8547 5367 8562 1 d0
rlabel metal1 5514 8770 5542 8775 1 vdd
rlabel metal1 5511 8377 5545 8383 1 gnd
rlabel locali 5347 7998 5369 8013 1 d0
rlabel metal1 5516 8221 5544 8226 1 vdd
rlabel metal1 5513 7828 5547 7834 1 gnd
rlabel locali 6284 7750 6312 7771 1 d1
rlabel metal1 6451 7584 6485 7590 1 gnd
rlabel metal1 6454 7977 6482 7982 1 vdd
rlabel locali 5346 7444 5368 7459 1 d0
rlabel metal1 5515 7667 5543 7672 1 vdd
rlabel metal1 5512 7274 5546 7280 1 gnd
rlabel metal1 6594 8488 6622 8493 1 vdd
rlabel metal1 6591 8095 6625 8101 1 gnd
rlabel locali 6422 8260 6443 8279 1 d2
rlabel locali 5347 6895 5369 6910 1 d0
rlabel metal1 5516 7118 5544 7123 1 vdd
rlabel metal1 5513 6725 5547 6731 1 gnd
rlabel locali 6284 6647 6312 6668 1 d1
rlabel metal1 6451 6481 6485 6487 1 gnd
rlabel metal1 6454 6874 6482 6879 1 vdd
rlabel locali 5346 6341 5368 6356 1 d0
rlabel metal1 5515 6564 5543 6569 1 vdd
rlabel metal1 5512 6171 5546 6177 1 gnd
rlabel locali 5348 5792 5370 5807 1 d0
rlabel metal1 5517 6015 5545 6020 1 vdd
rlabel metal1 5514 5622 5548 5628 1 gnd
rlabel locali 6285 5544 6313 5565 1 d1
rlabel metal1 6452 5378 6486 5384 1 gnd
rlabel metal1 6455 5771 6483 5776 1 vdd
rlabel locali 5347 5238 5369 5253 1 d0
rlabel metal1 5516 5461 5544 5466 1 vdd
rlabel metal1 5513 5068 5547 5074 1 gnd
rlabel metal1 6595 6282 6623 6287 1 vdd
rlabel metal1 6592 5889 6626 5895 1 gnd
rlabel locali 6423 6054 6444 6073 1 d2
rlabel metal1 6564 7398 6592 7403 1 vdd
rlabel metal1 6561 7005 6595 7011 1 gnd
rlabel locali 6394 7174 6420 7191 1 d3
rlabel locali 6396 2762 6422 2779 1 d3
rlabel metal1 6563 2593 6597 2599 1 gnd
rlabel metal1 6566 2986 6594 2991 1 vdd
rlabel locali 6425 1642 6446 1661 1 d2
rlabel metal1 6594 1477 6628 1483 1 gnd
rlabel metal1 6597 1870 6625 1875 1 vdd
rlabel metal1 5515 656 5549 662 1 gnd
rlabel metal1 5518 1049 5546 1054 1 vdd
rlabel locali 5349 826 5371 841 1 d0
rlabel metal1 6457 1359 6485 1364 1 vdd
rlabel metal1 6454 966 6488 972 1 gnd
rlabel locali 6287 1132 6315 1153 1 d1
rlabel metal1 5516 1210 5550 1216 1 gnd
rlabel metal1 5519 1603 5547 1608 1 vdd
rlabel locali 5350 1380 5372 1395 1 d0
rlabel metal1 5514 1759 5548 1765 1 gnd
rlabel metal1 5517 2152 5545 2157 1 vdd
rlabel locali 5348 1929 5370 1944 1 d0
rlabel metal1 6456 2462 6484 2467 1 vdd
rlabel metal1 6453 2069 6487 2075 1 gnd
rlabel locali 6286 2235 6314 2256 1 d1
rlabel metal1 5515 2313 5549 2319 1 gnd
rlabel metal1 5518 2706 5546 2711 1 vdd
rlabel locali 5349 2483 5371 2498 1 d0
rlabel locali 6424 3848 6445 3867 1 d2
rlabel metal1 6593 3683 6627 3689 1 gnd
rlabel metal1 6596 4076 6624 4081 1 vdd
rlabel metal1 5514 2862 5548 2868 1 gnd
rlabel metal1 5517 3255 5545 3260 1 vdd
rlabel locali 5348 3032 5370 3047 1 d0
rlabel metal1 6456 3565 6484 3570 1 vdd
rlabel metal1 6453 3172 6487 3178 1 gnd
rlabel locali 6286 3338 6314 3359 1 d1
rlabel metal1 5515 3416 5549 3422 1 gnd
rlabel metal1 5518 3809 5546 3814 1 vdd
rlabel locali 5349 3586 5371 3601 1 d0
rlabel metal1 5513 3965 5547 3971 1 gnd
rlabel metal1 5516 4358 5544 4363 1 vdd
rlabel locali 5347 4135 5369 4150 1 d0
rlabel metal1 6455 4668 6483 4673 1 vdd
rlabel metal1 6452 4275 6486 4281 1 gnd
rlabel locali 6285 4441 6313 4462 1 d1
rlabel metal1 5514 4519 5548 4525 1 gnd
rlabel metal1 5517 4912 5545 4917 1 vdd
rlabel locali 5348 4689 5370 4704 1 d0
rlabel metal1 6564 5198 6592 5203 1 vdd
rlabel metal1 6561 4805 6595 4811 1 gnd
rlabel locali 6388 4967 6423 4993 1 d4
rlabel locali 9677 947 9699 962 5 d0
rlabel metal1 9502 734 9530 739 5 vdd
rlabel metal1 9499 1126 9533 1132 5 gnd
rlabel locali 8734 1189 8762 1210 5 d1
rlabel metal1 8561 1370 8595 1376 5 gnd
rlabel metal1 8564 978 8592 983 5 vdd
rlabel locali 9678 1501 9700 1516 5 d0
rlabel metal1 9503 1288 9531 1293 5 vdd
rlabel metal1 9500 1680 9534 1686 5 gnd
rlabel locali 9676 2050 9698 2065 5 d0
rlabel metal1 9501 1837 9529 1842 5 vdd
rlabel metal1 9498 2229 9532 2235 5 gnd
rlabel locali 8733 2292 8761 2313 5 d1
rlabel metal1 8560 2473 8594 2479 5 gnd
rlabel metal1 8563 2081 8591 2086 5 vdd
rlabel locali 9677 2604 9699 2619 5 d0
rlabel metal1 9502 2391 9530 2396 5 vdd
rlabel metal1 9499 2783 9533 2789 5 gnd
rlabel metal1 8423 1570 8451 1575 5 vdd
rlabel metal1 8420 1962 8454 1968 5 gnd
rlabel locali 8602 1784 8623 1803 5 d2
rlabel locali 9676 3153 9698 3168 5 d0
rlabel metal1 9501 2940 9529 2945 5 vdd
rlabel metal1 9498 3332 9532 3338 5 gnd
rlabel locali 8733 3395 8761 3416 5 d1
rlabel metal1 8560 3576 8594 3582 5 gnd
rlabel metal1 8563 3184 8591 3189 5 vdd
rlabel locali 9677 3707 9699 3722 5 d0
rlabel metal1 9502 3494 9530 3499 5 vdd
rlabel metal1 9499 3886 9533 3892 5 gnd
rlabel locali 9675 4256 9697 4271 5 d0
rlabel metal1 9500 4043 9528 4048 5 vdd
rlabel metal1 9497 4435 9531 4441 5 gnd
rlabel locali 8732 4498 8760 4519 5 d1
rlabel metal1 8559 4679 8593 4685 5 gnd
rlabel metal1 8562 4287 8590 4292 5 vdd
rlabel locali 9676 4810 9698 4825 5 d0
rlabel metal1 9501 4597 9529 4602 5 vdd
rlabel metal1 9498 4989 9532 4995 5 gnd
rlabel metal1 8422 3776 8450 3781 5 vdd
rlabel metal1 8419 4168 8453 4174 5 gnd
rlabel locali 8601 3990 8622 4009 5 d2
rlabel metal1 8453 2660 8481 2665 5 vdd
rlabel metal1 8450 3052 8484 3058 5 gnd
rlabel locali 8625 2872 8651 2889 5 d3
rlabel locali 8623 7284 8649 7301 5 d3
rlabel metal1 8448 7464 8482 7470 5 gnd
rlabel metal1 8451 7072 8479 7077 5 vdd
rlabel locali 8599 8402 8620 8421 5 d2
rlabel metal1 8417 8580 8451 8586 5 gnd
rlabel metal1 8420 8188 8448 8193 5 vdd
rlabel metal1 9496 9401 9530 9407 5 gnd
rlabel metal1 9499 9009 9527 9014 5 vdd
rlabel locali 9674 9222 9696 9237 5 d0
rlabel metal1 8560 8699 8588 8704 5 vdd
rlabel metal1 8557 9091 8591 9097 5 gnd
rlabel locali 8730 8910 8758 8931 5 d1
rlabel metal1 9495 8847 9529 8853 5 gnd
rlabel metal1 9498 8455 9526 8460 5 vdd
rlabel locali 9673 8668 9695 8683 5 d0
rlabel metal1 9497 8298 9531 8304 5 gnd
rlabel metal1 9500 7906 9528 7911 5 vdd
rlabel locali 9675 8119 9697 8134 5 d0
rlabel metal1 8561 7596 8589 7601 5 vdd
rlabel metal1 8558 7988 8592 7994 5 gnd
rlabel locali 8731 7807 8759 7828 5 d1
rlabel metal1 9496 7744 9530 7750 5 gnd
rlabel metal1 9499 7352 9527 7357 5 vdd
rlabel locali 9674 7565 9696 7580 5 d0
rlabel locali 8600 6196 8621 6215 5 d2
rlabel metal1 8418 6374 8452 6380 5 gnd
rlabel metal1 8421 5982 8449 5987 5 vdd
rlabel metal1 9497 7195 9531 7201 5 gnd
rlabel metal1 9500 6803 9528 6808 5 vdd
rlabel locali 9675 7016 9697 7031 5 d0
rlabel metal1 8561 6493 8589 6498 5 vdd
rlabel metal1 8558 6885 8592 6891 5 gnd
rlabel locali 8731 6704 8759 6725 5 d1
rlabel metal1 9496 6641 9530 6647 5 gnd
rlabel metal1 9499 6249 9527 6254 5 vdd
rlabel locali 9674 6462 9696 6477 5 d0
rlabel metal1 9498 6092 9532 6098 5 gnd
rlabel metal1 9501 5700 9529 5705 5 vdd
rlabel locali 9676 5913 9698 5928 5 d0
rlabel metal1 8562 5390 8590 5395 5 vdd
rlabel metal1 8559 5782 8593 5788 5 gnd
rlabel locali 8732 5601 8760 5622 5 d1
rlabel metal1 9497 5538 9531 5544 5 gnd
rlabel metal1 9500 5146 9528 5151 5 vdd
rlabel locali 9675 5359 9697 5374 5 d0
rlabel metal1 8453 4860 8481 4865 5 vdd
rlabel metal1 8450 5252 8484 5258 5 gnd
rlabel locali 8622 5070 8657 5096 5 d4
rlabel metal1 6765 490 6793 495 1 vdd
rlabel metal1 6762 97 6796 103 1 gnd
rlabel locali 6591 261 6619 283 1 d5
rlabel metal1 4659 429 4687 434 1 vdd
rlabel metal1 4656 36 4690 42 1 gnd
rlabel locali 4488 199 4515 225 1 d6
rlabel locali 10321 9065 10343 9080 1 d0
rlabel metal1 10490 9288 10518 9293 1 vdd
rlabel metal1 10487 8895 10521 8901 1 gnd
rlabel locali 11258 8817 11286 8838 1 d1
rlabel metal1 11425 8651 11459 8657 1 gnd
rlabel metal1 11428 9044 11456 9049 1 vdd
rlabel locali 10320 8511 10342 8526 1 d0
rlabel metal1 10489 8734 10517 8739 1 vdd
rlabel metal1 10486 8341 10520 8347 1 gnd
rlabel locali 10322 7962 10344 7977 1 d0
rlabel metal1 10491 8185 10519 8190 1 vdd
rlabel metal1 10488 7792 10522 7798 1 gnd
rlabel locali 11259 7714 11287 7735 1 d1
rlabel metal1 11426 7548 11460 7554 1 gnd
rlabel metal1 11429 7941 11457 7946 1 vdd
rlabel locali 10321 7408 10343 7423 1 d0
rlabel metal1 10490 7631 10518 7636 1 vdd
rlabel metal1 10487 7238 10521 7244 1 gnd
rlabel metal1 11569 8452 11597 8457 1 vdd
rlabel metal1 11566 8059 11600 8065 1 gnd
rlabel locali 11397 8224 11418 8243 1 d2
rlabel locali 10322 6859 10344 6874 1 d0
rlabel metal1 10491 7082 10519 7087 1 vdd
rlabel metal1 10488 6689 10522 6695 1 gnd
rlabel locali 11259 6611 11287 6632 1 d1
rlabel metal1 11426 6445 11460 6451 1 gnd
rlabel metal1 11429 6838 11457 6843 1 vdd
rlabel locali 10321 6305 10343 6320 1 d0
rlabel metal1 10490 6528 10518 6533 1 vdd
rlabel metal1 10487 6135 10521 6141 1 gnd
rlabel locali 10323 5756 10345 5771 1 d0
rlabel metal1 10492 5979 10520 5984 1 vdd
rlabel metal1 10489 5586 10523 5592 1 gnd
rlabel locali 11260 5508 11288 5529 1 d1
rlabel metal1 11427 5342 11461 5348 1 gnd
rlabel metal1 11430 5735 11458 5740 1 vdd
rlabel locali 10322 5202 10344 5217 1 d0
rlabel metal1 10491 5425 10519 5430 1 vdd
rlabel metal1 10488 5032 10522 5038 1 gnd
rlabel metal1 11570 6246 11598 6251 1 vdd
rlabel metal1 11567 5853 11601 5859 1 gnd
rlabel locali 11398 6018 11419 6037 1 d2
rlabel metal1 11539 7362 11567 7367 1 vdd
rlabel metal1 11536 6969 11570 6975 1 gnd
rlabel locali 11369 7138 11395 7155 1 d3
rlabel locali 11371 2726 11397 2743 1 d3
rlabel metal1 11538 2557 11572 2563 1 gnd
rlabel metal1 11541 2950 11569 2955 1 vdd
rlabel locali 11400 1606 11421 1625 1 d2
rlabel metal1 11569 1441 11603 1447 1 gnd
rlabel metal1 11572 1834 11600 1839 1 vdd
rlabel metal1 10490 620 10524 626 1 gnd
rlabel metal1 10493 1013 10521 1018 1 vdd
rlabel locali 10324 790 10346 805 1 d0
rlabel metal1 11432 1323 11460 1328 1 vdd
rlabel metal1 11429 930 11463 936 1 gnd
rlabel locali 11262 1096 11290 1117 1 d1
rlabel metal1 10491 1174 10525 1180 1 gnd
rlabel metal1 10494 1567 10522 1572 1 vdd
rlabel locali 10325 1344 10347 1359 1 d0
rlabel metal1 10489 1723 10523 1729 1 gnd
rlabel metal1 10492 2116 10520 2121 1 vdd
rlabel locali 10323 1893 10345 1908 1 d0
rlabel metal1 11431 2426 11459 2431 1 vdd
rlabel metal1 11428 2033 11462 2039 1 gnd
rlabel locali 11261 2199 11289 2220 1 d1
rlabel metal1 10490 2277 10524 2283 1 gnd
rlabel metal1 10493 2670 10521 2675 1 vdd
rlabel locali 10324 2447 10346 2462 1 d0
rlabel locali 11399 3812 11420 3831 1 d2
rlabel metal1 11568 3647 11602 3653 1 gnd
rlabel metal1 11571 4040 11599 4045 1 vdd
rlabel metal1 10489 2826 10523 2832 1 gnd
rlabel metal1 10492 3219 10520 3224 1 vdd
rlabel locali 10323 2996 10345 3011 1 d0
rlabel metal1 11431 3529 11459 3534 1 vdd
rlabel metal1 11428 3136 11462 3142 1 gnd
rlabel locali 11261 3302 11289 3323 1 d1
rlabel metal1 10490 3380 10524 3386 1 gnd
rlabel metal1 10493 3773 10521 3778 1 vdd
rlabel locali 10324 3550 10346 3565 1 d0
rlabel metal1 10488 3929 10522 3935 1 gnd
rlabel metal1 10491 4322 10519 4327 1 vdd
rlabel locali 10322 4099 10344 4114 1 d0
rlabel metal1 11430 4632 11458 4637 1 vdd
rlabel metal1 11427 4239 11461 4245 1 gnd
rlabel locali 11260 4405 11288 4426 1 d1
rlabel metal1 10489 4483 10523 4489 1 gnd
rlabel metal1 10492 4876 10520 4881 1 vdd
rlabel locali 10323 4653 10345 4668 1 d0
rlabel metal1 11539 5162 11567 5167 1 vdd
rlabel metal1 11536 4769 11570 4775 1 gnd
rlabel locali 11363 4931 11398 4957 1 d4
rlabel locali 14652 911 14674 926 5 d0
rlabel metal1 14477 698 14505 703 5 vdd
rlabel metal1 14474 1090 14508 1096 5 gnd
rlabel locali 13709 1153 13737 1174 5 d1
rlabel metal1 13536 1334 13570 1340 5 gnd
rlabel metal1 13539 942 13567 947 5 vdd
rlabel locali 14653 1465 14675 1480 5 d0
rlabel metal1 14478 1252 14506 1257 5 vdd
rlabel metal1 14475 1644 14509 1650 5 gnd
rlabel locali 14651 2014 14673 2029 5 d0
rlabel metal1 14476 1801 14504 1806 5 vdd
rlabel metal1 14473 2193 14507 2199 5 gnd
rlabel locali 13708 2256 13736 2277 5 d1
rlabel metal1 13535 2437 13569 2443 5 gnd
rlabel metal1 13538 2045 13566 2050 5 vdd
rlabel locali 14652 2568 14674 2583 5 d0
rlabel metal1 14477 2355 14505 2360 5 vdd
rlabel metal1 14474 2747 14508 2753 5 gnd
rlabel metal1 13398 1534 13426 1539 5 vdd
rlabel metal1 13395 1926 13429 1932 5 gnd
rlabel locali 13577 1748 13598 1767 5 d2
rlabel locali 14651 3117 14673 3132 5 d0
rlabel metal1 14476 2904 14504 2909 5 vdd
rlabel metal1 14473 3296 14507 3302 5 gnd
rlabel locali 13708 3359 13736 3380 5 d1
rlabel metal1 13535 3540 13569 3546 5 gnd
rlabel metal1 13538 3148 13566 3153 5 vdd
rlabel locali 14652 3671 14674 3686 5 d0
rlabel metal1 14477 3458 14505 3463 5 vdd
rlabel metal1 14474 3850 14508 3856 5 gnd
rlabel locali 14650 4220 14672 4235 5 d0
rlabel metal1 14475 4007 14503 4012 5 vdd
rlabel metal1 14472 4399 14506 4405 5 gnd
rlabel locali 13707 4462 13735 4483 5 d1
rlabel metal1 13534 4643 13568 4649 5 gnd
rlabel metal1 13537 4251 13565 4256 5 vdd
rlabel locali 14651 4774 14673 4789 5 d0
rlabel metal1 14476 4561 14504 4566 5 vdd
rlabel metal1 14473 4953 14507 4959 5 gnd
rlabel metal1 13397 3740 13425 3745 5 vdd
rlabel metal1 13394 4132 13428 4138 5 gnd
rlabel locali 13576 3954 13597 3973 5 d2
rlabel metal1 13428 2624 13456 2629 5 vdd
rlabel metal1 13425 3016 13459 3022 5 gnd
rlabel locali 13600 2836 13626 2853 5 d3
rlabel locali 13598 7248 13624 7265 5 d3
rlabel metal1 13423 7428 13457 7434 5 gnd
rlabel metal1 13426 7036 13454 7041 5 vdd
rlabel locali 13574 8366 13595 8385 5 d2
rlabel metal1 13392 8544 13426 8550 5 gnd
rlabel metal1 13395 8152 13423 8157 5 vdd
rlabel metal1 14471 9365 14505 9371 5 gnd
rlabel metal1 14474 8973 14502 8978 5 vdd
rlabel locali 14649 9186 14671 9201 5 d0
rlabel metal1 13535 8663 13563 8668 5 vdd
rlabel metal1 13532 9055 13566 9061 5 gnd
rlabel locali 13705 8874 13733 8895 5 d1
rlabel metal1 14470 8811 14504 8817 5 gnd
rlabel metal1 14473 8419 14501 8424 5 vdd
rlabel locali 14648 8632 14670 8647 5 d0
rlabel metal1 14472 8262 14506 8268 5 gnd
rlabel metal1 14475 7870 14503 7875 5 vdd
rlabel locali 14650 8083 14672 8098 5 d0
rlabel metal1 13536 7560 13564 7565 5 vdd
rlabel metal1 13533 7952 13567 7958 5 gnd
rlabel locali 13706 7771 13734 7792 5 d1
rlabel metal1 14471 7708 14505 7714 5 gnd
rlabel metal1 14474 7316 14502 7321 5 vdd
rlabel locali 14649 7529 14671 7544 5 d0
rlabel locali 13575 6160 13596 6179 5 d2
rlabel metal1 13393 6338 13427 6344 5 gnd
rlabel metal1 13396 5946 13424 5951 5 vdd
rlabel metal1 14472 7159 14506 7165 5 gnd
rlabel metal1 14475 6767 14503 6772 5 vdd
rlabel locali 14650 6980 14672 6995 5 d0
rlabel metal1 13536 6457 13564 6462 5 vdd
rlabel metal1 13533 6849 13567 6855 5 gnd
rlabel locali 13706 6668 13734 6689 5 d1
rlabel metal1 14471 6605 14505 6611 5 gnd
rlabel metal1 14474 6213 14502 6218 5 vdd
rlabel locali 14649 6426 14671 6441 5 d0
rlabel metal1 14473 6056 14507 6062 5 gnd
rlabel metal1 14476 5664 14504 5669 5 vdd
rlabel locali 14651 5877 14673 5892 5 d0
rlabel metal1 13537 5354 13565 5359 5 vdd
rlabel metal1 13534 5746 13568 5752 5 gnd
rlabel locali 13707 5565 13735 5586 5 d1
rlabel metal1 14472 5502 14506 5508 5 gnd
rlabel metal1 14475 5110 14503 5115 5 vdd
rlabel locali 14650 5323 14672 5338 5 d0
rlabel metal1 13428 4824 13456 4829 5 vdd
rlabel metal1 13425 5216 13459 5222 5 gnd
rlabel locali 13597 5034 13632 5060 5 d4
rlabel metal1 11740 454 11768 459 1 vdd
rlabel metal1 11737 61 11771 67 1 gnd
rlabel locali 11566 225 11594 247 1 d5
rlabel locali 15377 9106 15399 9121 1 d0
rlabel metal1 15546 9329 15574 9334 1 vdd
rlabel metal1 15543 8936 15577 8942 1 gnd
rlabel locali 16314 8858 16342 8879 1 d1
rlabel metal1 16481 8692 16515 8698 1 gnd
rlabel metal1 16484 9085 16512 9090 1 vdd
rlabel locali 15376 8552 15398 8567 1 d0
rlabel metal1 15545 8775 15573 8780 1 vdd
rlabel metal1 15542 8382 15576 8388 1 gnd
rlabel locali 15378 8003 15400 8018 1 d0
rlabel metal1 15547 8226 15575 8231 1 vdd
rlabel metal1 15544 7833 15578 7839 1 gnd
rlabel locali 16315 7755 16343 7776 1 d1
rlabel metal1 16482 7589 16516 7595 1 gnd
rlabel metal1 16485 7982 16513 7987 1 vdd
rlabel locali 15377 7449 15399 7464 1 d0
rlabel metal1 15546 7672 15574 7677 1 vdd
rlabel metal1 15543 7279 15577 7285 1 gnd
rlabel metal1 16625 8493 16653 8498 1 vdd
rlabel metal1 16622 8100 16656 8106 1 gnd
rlabel locali 16453 8265 16474 8284 1 d2
rlabel locali 15378 6900 15400 6915 1 d0
rlabel metal1 15547 7123 15575 7128 1 vdd
rlabel metal1 15544 6730 15578 6736 1 gnd
rlabel locali 16315 6652 16343 6673 1 d1
rlabel metal1 16482 6486 16516 6492 1 gnd
rlabel metal1 16485 6879 16513 6884 1 vdd
rlabel locali 15377 6346 15399 6361 1 d0
rlabel metal1 15546 6569 15574 6574 1 vdd
rlabel metal1 15543 6176 15577 6182 1 gnd
rlabel locali 15379 5797 15401 5812 1 d0
rlabel metal1 15548 6020 15576 6025 1 vdd
rlabel metal1 15545 5627 15579 5633 1 gnd
rlabel locali 16316 5549 16344 5570 1 d1
rlabel metal1 16483 5383 16517 5389 1 gnd
rlabel metal1 16486 5776 16514 5781 1 vdd
rlabel locali 15378 5243 15400 5258 1 d0
rlabel metal1 15547 5466 15575 5471 1 vdd
rlabel metal1 15544 5073 15578 5079 1 gnd
rlabel metal1 16626 6287 16654 6292 1 vdd
rlabel metal1 16623 5894 16657 5900 1 gnd
rlabel locali 16454 6059 16475 6078 1 d2
rlabel metal1 16595 7403 16623 7408 1 vdd
rlabel metal1 16592 7010 16626 7016 1 gnd
rlabel locali 16425 7179 16451 7196 1 d3
rlabel locali 16427 2767 16453 2784 1 d3
rlabel metal1 16594 2598 16628 2604 1 gnd
rlabel metal1 16597 2991 16625 2996 1 vdd
rlabel locali 16456 1647 16477 1666 1 d2
rlabel metal1 16625 1482 16659 1488 1 gnd
rlabel metal1 16628 1875 16656 1880 1 vdd
rlabel metal1 15546 661 15580 667 1 gnd
rlabel metal1 15549 1054 15577 1059 1 vdd
rlabel locali 15380 831 15402 846 1 d0
rlabel metal1 16488 1364 16516 1369 1 vdd
rlabel metal1 16485 971 16519 977 1 gnd
rlabel locali 16318 1137 16346 1158 1 d1
rlabel metal1 15547 1215 15581 1221 1 gnd
rlabel metal1 15550 1608 15578 1613 1 vdd
rlabel locali 15381 1385 15403 1400 1 d0
rlabel metal1 15545 1764 15579 1770 1 gnd
rlabel metal1 15548 2157 15576 2162 1 vdd
rlabel locali 15379 1934 15401 1949 1 d0
rlabel metal1 16487 2467 16515 2472 1 vdd
rlabel metal1 16484 2074 16518 2080 1 gnd
rlabel locali 16317 2240 16345 2261 1 d1
rlabel metal1 15546 2318 15580 2324 1 gnd
rlabel metal1 15549 2711 15577 2716 1 vdd
rlabel locali 15380 2488 15402 2503 1 d0
rlabel locali 16455 3853 16476 3872 1 d2
rlabel metal1 16624 3688 16658 3694 1 gnd
rlabel metal1 16627 4081 16655 4086 1 vdd
rlabel metal1 15545 2867 15579 2873 1 gnd
rlabel metal1 15548 3260 15576 3265 1 vdd
rlabel locali 15379 3037 15401 3052 1 d0
rlabel metal1 16487 3570 16515 3575 1 vdd
rlabel metal1 16484 3177 16518 3183 1 gnd
rlabel locali 16317 3343 16345 3364 1 d1
rlabel metal1 15546 3421 15580 3427 1 gnd
rlabel metal1 15549 3814 15577 3819 1 vdd
rlabel locali 15380 3591 15402 3606 1 d0
rlabel metal1 15544 3970 15578 3976 1 gnd
rlabel metal1 15547 4363 15575 4368 1 vdd
rlabel locali 15378 4140 15400 4155 1 d0
rlabel metal1 16486 4673 16514 4678 1 vdd
rlabel metal1 16483 4280 16517 4286 1 gnd
rlabel locali 16316 4446 16344 4467 1 d1
rlabel metal1 15545 4524 15579 4530 1 gnd
rlabel metal1 15548 4917 15576 4922 1 vdd
rlabel locali 15379 4694 15401 4709 1 d0
rlabel metal1 16595 5203 16623 5208 1 vdd
rlabel metal1 16592 4810 16626 4816 1 gnd
rlabel locali 16419 4972 16454 4998 1 d4
rlabel locali 19708 952 19730 967 5 d0
rlabel metal1 19533 739 19561 744 5 vdd
rlabel metal1 19530 1131 19564 1137 5 gnd
rlabel locali 18765 1194 18793 1215 5 d1
rlabel metal1 18592 1375 18626 1381 5 gnd
rlabel metal1 18595 983 18623 988 5 vdd
rlabel locali 19709 1506 19731 1521 5 d0
rlabel metal1 19534 1293 19562 1298 5 vdd
rlabel metal1 19531 1685 19565 1691 5 gnd
rlabel locali 19707 2055 19729 2070 5 d0
rlabel metal1 19532 1842 19560 1847 5 vdd
rlabel metal1 19529 2234 19563 2240 5 gnd
rlabel locali 18764 2297 18792 2318 5 d1
rlabel metal1 18591 2478 18625 2484 5 gnd
rlabel metal1 18594 2086 18622 2091 5 vdd
rlabel locali 19708 2609 19730 2624 5 d0
rlabel metal1 19533 2396 19561 2401 5 vdd
rlabel metal1 19530 2788 19564 2794 5 gnd
rlabel metal1 18454 1575 18482 1580 5 vdd
rlabel metal1 18451 1967 18485 1973 5 gnd
rlabel locali 18633 1789 18654 1808 5 d2
rlabel locali 19707 3158 19729 3173 5 d0
rlabel metal1 19532 2945 19560 2950 5 vdd
rlabel metal1 19529 3337 19563 3343 5 gnd
rlabel locali 18764 3400 18792 3421 5 d1
rlabel metal1 18591 3581 18625 3587 5 gnd
rlabel metal1 18594 3189 18622 3194 5 vdd
rlabel locali 19708 3712 19730 3727 5 d0
rlabel metal1 19533 3499 19561 3504 5 vdd
rlabel metal1 19530 3891 19564 3897 5 gnd
rlabel locali 19706 4261 19728 4276 5 d0
rlabel metal1 19531 4048 19559 4053 5 vdd
rlabel metal1 19528 4440 19562 4446 5 gnd
rlabel locali 18763 4503 18791 4524 5 d1
rlabel metal1 18590 4684 18624 4690 5 gnd
rlabel metal1 18593 4292 18621 4297 5 vdd
rlabel locali 19707 4815 19729 4830 5 d0
rlabel metal1 19532 4602 19560 4607 5 vdd
rlabel metal1 19529 4994 19563 5000 5 gnd
rlabel metal1 18453 3781 18481 3786 5 vdd
rlabel metal1 18450 4173 18484 4179 5 gnd
rlabel locali 18632 3995 18653 4014 5 d2
rlabel metal1 18484 2665 18512 2670 5 vdd
rlabel metal1 18481 3057 18515 3063 5 gnd
rlabel locali 18656 2877 18682 2894 5 d3
rlabel locali 18654 7289 18680 7306 5 d3
rlabel metal1 18479 7469 18513 7475 5 gnd
rlabel metal1 18482 7077 18510 7082 5 vdd
rlabel locali 18630 8407 18651 8426 5 d2
rlabel metal1 18448 8585 18482 8591 5 gnd
rlabel metal1 18451 8193 18479 8198 5 vdd
rlabel metal1 19527 9406 19561 9412 5 gnd
rlabel metal1 19530 9014 19558 9019 5 vdd
rlabel locali 19705 9227 19727 9242 5 d0
rlabel metal1 18591 8704 18619 8709 5 vdd
rlabel metal1 18588 9096 18622 9102 5 gnd
rlabel locali 18761 8915 18789 8936 5 d1
rlabel metal1 19526 8852 19560 8858 5 gnd
rlabel metal1 19529 8460 19557 8465 5 vdd
rlabel locali 19704 8673 19726 8688 5 d0
rlabel metal1 19528 8303 19562 8309 5 gnd
rlabel metal1 19531 7911 19559 7916 5 vdd
rlabel locali 19706 8124 19728 8139 5 d0
rlabel metal1 18592 7601 18620 7606 5 vdd
rlabel metal1 18589 7993 18623 7999 5 gnd
rlabel locali 18762 7812 18790 7833 5 d1
rlabel metal1 19527 7749 19561 7755 5 gnd
rlabel metal1 19530 7357 19558 7362 5 vdd
rlabel locali 19705 7570 19727 7585 5 d0
rlabel locali 18631 6201 18652 6220 5 d2
rlabel metal1 18449 6379 18483 6385 5 gnd
rlabel metal1 18452 5987 18480 5992 5 vdd
rlabel metal1 19528 7200 19562 7206 5 gnd
rlabel metal1 19531 6808 19559 6813 5 vdd
rlabel locali 19706 7021 19728 7036 5 d0
rlabel metal1 18592 6498 18620 6503 5 vdd
rlabel metal1 18589 6890 18623 6896 5 gnd
rlabel locali 18762 6709 18790 6730 5 d1
rlabel metal1 19527 6646 19561 6652 5 gnd
rlabel metal1 19530 6254 19558 6259 5 vdd
rlabel locali 19705 6467 19727 6482 5 d0
rlabel metal1 19529 6097 19563 6103 5 gnd
rlabel metal1 19532 5705 19560 5710 5 vdd
rlabel locali 19707 5918 19729 5933 5 d0
rlabel metal1 18593 5395 18621 5400 5 vdd
rlabel metal1 18590 5787 18624 5793 5 gnd
rlabel locali 18763 5606 18791 5627 5 d1
rlabel metal1 19528 5543 19562 5549 5 gnd
rlabel metal1 19531 5151 19559 5156 5 vdd
rlabel locali 19706 5364 19728 5379 5 d0
rlabel metal1 18484 4865 18512 4870 5 vdd
rlabel metal1 18481 5257 18515 5263 5 gnd
rlabel locali 18653 5075 18688 5101 5 d4
rlabel metal1 16796 495 16824 500 1 vdd
rlabel metal1 16793 102 16827 108 1 gnd
rlabel locali 16622 266 16650 288 1 d5
rlabel metal1 14690 434 14718 439 1 vdd
rlabel metal1 14687 41 14721 47 1 gnd
rlabel locali 14519 204 14546 230 1 d6
rlabel metal1 9593 313 9621 318 1 vdd
rlabel metal1 9590 -80 9624 -74 1 gnd
rlabel locali 9415 89 9446 108 1 d7
rlabel locali 10052 130 10076 159 1 vout
<< end >>
