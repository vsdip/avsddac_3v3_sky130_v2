magic
tech sky130A
timestamp 1633172786
<< nwell >>
rect 869 13580 1680 13804
rect 1917 13576 2728 13800
rect 11577 13574 12388 13798
rect 12625 13570 13436 13794
rect 22542 13578 23353 13802
rect 23590 13574 24401 13798
rect 33250 13572 34061 13796
rect 34298 13568 35109 13792
rect 9155 13325 9966 13549
rect 19863 13319 20674 13543
rect 30828 13323 31639 13547
rect 41536 13317 42347 13541
rect 869 12901 1680 13125
rect 3364 12896 4175 13120
rect 11577 12895 12388 13119
rect 14072 12890 14883 13114
rect 22542 12899 23353 13123
rect 25037 12894 25848 13118
rect 33250 12893 34061 13117
rect 35745 12888 36556 13112
rect 8107 12650 8918 12874
rect 9155 12646 9966 12870
rect 18815 12644 19626 12868
rect 19863 12640 20674 12864
rect 29780 12648 30591 12872
rect 30828 12644 31639 12868
rect 40488 12642 41299 12866
rect 41536 12638 42347 12862
rect 869 12133 1680 12357
rect 1917 12129 2728 12353
rect 11577 12127 12388 12351
rect 12625 12123 13436 12347
rect 22542 12131 23353 12355
rect 23590 12127 24401 12351
rect 33250 12125 34061 12349
rect 34298 12121 35109 12345
rect 6660 11883 7471 12107
rect 9155 11878 9966 12102
rect 17368 11877 18179 12101
rect 19863 11872 20674 12096
rect 28333 11881 29144 12105
rect 30828 11876 31639 12100
rect 39041 11875 39852 12099
rect 41536 11870 42347 12094
rect 869 11454 1680 11678
rect 3407 11451 4218 11675
rect 11577 11448 12388 11672
rect 14115 11445 14926 11669
rect 22542 11452 23353 11676
rect 25080 11449 25891 11673
rect 33250 11446 34061 11670
rect 35788 11443 36599 11667
rect 8107 11203 8918 11427
rect 9155 11199 9966 11423
rect 18815 11197 19626 11421
rect 19863 11193 20674 11417
rect 29780 11201 30591 11425
rect 30828 11197 31639 11421
rect 40488 11195 41299 11419
rect 41536 11191 42347 11415
rect 870 10613 1681 10837
rect 1918 10609 2729 10833
rect 11578 10607 12389 10831
rect 12626 10603 13437 10827
rect 22543 10611 23354 10835
rect 23591 10607 24402 10831
rect 33251 10605 34062 10829
rect 34299 10601 35110 10825
rect 6618 10361 7429 10585
rect 9156 10358 9967 10582
rect 17326 10355 18137 10579
rect 19864 10352 20675 10576
rect 28291 10359 29102 10583
rect 30829 10356 31640 10580
rect 38999 10353 39810 10577
rect 41537 10350 42348 10574
rect 870 9934 1681 10158
rect 3365 9929 4176 10153
rect 11578 9928 12389 10152
rect 14073 9923 14884 10147
rect 22543 9932 23354 10156
rect 25038 9927 25849 10151
rect 33251 9926 34062 10150
rect 35746 9921 36557 10145
rect 8108 9683 8919 9907
rect 9156 9679 9967 9903
rect 18816 9677 19627 9901
rect 19864 9673 20675 9897
rect 29781 9681 30592 9905
rect 30829 9677 31640 9901
rect 40489 9675 41300 9899
rect 41537 9671 42348 9895
rect 870 9166 1681 9390
rect 1918 9162 2729 9386
rect 11578 9160 12389 9384
rect 12626 9156 13437 9380
rect 22543 9164 23354 9388
rect 23591 9160 24402 9384
rect 33251 9158 34062 9382
rect 34299 9154 35110 9378
rect 6661 8916 7472 9140
rect 9156 8911 9967 9135
rect 17369 8910 18180 9134
rect 19864 8905 20675 9129
rect 28334 8914 29145 9138
rect 30829 8909 31640 9133
rect 39042 8908 39853 9132
rect 41537 8903 42348 9127
rect 870 8487 1681 8711
rect 4473 8478 5284 8702
rect 11578 8481 12389 8705
rect 15181 8472 15992 8696
rect 22543 8485 23354 8709
rect 26146 8476 26957 8700
rect 33251 8479 34062 8703
rect 36854 8470 37665 8694
rect 8108 8236 8919 8460
rect 9156 8232 9967 8456
rect 18816 8230 19627 8454
rect 19864 8226 20675 8450
rect 29781 8234 30592 8458
rect 30829 8230 31640 8454
rect 40489 8228 41300 8452
rect 41537 8224 42348 8448
rect 867 7572 1678 7796
rect 1915 7568 2726 7792
rect 11575 7566 12386 7790
rect 12623 7562 13434 7786
rect 22540 7570 23351 7794
rect 23588 7566 24399 7790
rect 33248 7564 34059 7788
rect 34296 7560 35107 7784
rect 5550 7326 6361 7550
rect 9153 7317 9964 7541
rect 16258 7320 17069 7544
rect 19861 7311 20672 7535
rect 27223 7324 28034 7548
rect 30826 7315 31637 7539
rect 37931 7318 38742 7542
rect 41534 7309 42345 7533
rect 867 6893 1678 7117
rect 3362 6888 4173 7112
rect 11575 6887 12386 7111
rect 14070 6882 14881 7106
rect 22540 6891 23351 7115
rect 25035 6886 25846 7110
rect 33248 6885 34059 7109
rect 35743 6880 36554 7104
rect 8105 6642 8916 6866
rect 9153 6638 9964 6862
rect 18813 6636 19624 6860
rect 19861 6632 20672 6856
rect 29778 6640 30589 6864
rect 30826 6636 31637 6860
rect 40486 6634 41297 6858
rect 41534 6630 42345 6854
rect 867 6125 1678 6349
rect 1915 6121 2726 6345
rect 11575 6119 12386 6343
rect 12623 6115 13434 6339
rect 22540 6123 23351 6347
rect 23588 6119 24399 6343
rect 33248 6117 34059 6341
rect 34296 6113 35107 6337
rect 6658 5875 7469 6099
rect 9153 5870 9964 6094
rect 17366 5869 18177 6093
rect 19861 5864 20672 6088
rect 28331 5873 29142 6097
rect 30826 5868 31637 6092
rect 39039 5867 39850 6091
rect 41534 5862 42345 6086
rect 867 5446 1678 5670
rect 3405 5443 4216 5667
rect 11575 5440 12386 5664
rect 14113 5437 14924 5661
rect 22540 5444 23351 5668
rect 25078 5441 25889 5665
rect 33248 5438 34059 5662
rect 35786 5435 36597 5659
rect 8105 5195 8916 5419
rect 9153 5191 9964 5415
rect 18813 5189 19624 5413
rect 19861 5185 20672 5409
rect 29778 5193 30589 5417
rect 30826 5189 31637 5413
rect 40486 5187 41297 5411
rect 41534 5183 42345 5407
rect 868 4605 1679 4829
rect 1916 4601 2727 4825
rect 4818 4607 5629 4831
rect 11576 4599 12387 4823
rect 12624 4595 13435 4819
rect 15526 4601 16337 4825
rect 22541 4603 23352 4827
rect 23589 4599 24400 4823
rect 26491 4605 27302 4829
rect 33249 4597 34060 4821
rect 34297 4593 35108 4817
rect 37199 4599 38010 4823
rect 6616 4353 7427 4577
rect 9154 4350 9965 4574
rect 17324 4347 18135 4571
rect 19862 4344 20673 4568
rect 28289 4351 29100 4575
rect 30827 4348 31638 4572
rect 38997 4345 39808 4569
rect 41535 4342 42346 4566
rect 868 3926 1679 4150
rect 3363 3921 4174 4145
rect 11576 3920 12387 4144
rect 14071 3915 14882 4139
rect 22541 3924 23352 4148
rect 25036 3919 25847 4143
rect 33249 3918 34060 4142
rect 35744 3913 36555 4137
rect 8106 3675 8917 3899
rect 9154 3671 9965 3895
rect 18814 3669 19625 3893
rect 19862 3665 20673 3889
rect 29779 3673 30590 3897
rect 30827 3669 31638 3893
rect 40487 3667 41298 3891
rect 41535 3663 42346 3887
rect 868 3158 1679 3382
rect 1916 3154 2727 3378
rect 11576 3152 12387 3376
rect 12624 3148 13435 3372
rect 22541 3156 23352 3380
rect 23589 3152 24400 3376
rect 33249 3150 34060 3374
rect 34297 3146 35108 3370
rect 6659 2908 7470 3132
rect 9154 2903 9965 3127
rect 17367 2902 18178 3126
rect 19862 2897 20673 3121
rect 28332 2906 29143 3130
rect 30827 2901 31638 3125
rect 39040 2900 39851 3124
rect 41535 2895 42346 3119
rect 868 2479 1679 2703
rect 11576 2473 12387 2697
rect 22541 2477 23352 2701
rect 33249 2471 34060 2695
rect 8106 2228 8917 2452
rect 9154 2224 9965 2448
rect 18814 2222 19625 2446
rect 19862 2218 20673 2442
rect 29779 2226 30590 2450
rect 30827 2222 31638 2446
rect 40487 2220 41298 2444
rect 41535 2216 42346 2440
rect 10579 320 11390 544
rect 21216 307 22027 531
rect 32252 318 33063 542
<< nmos >>
rect 9223 13608 9273 13650
rect 9431 13608 9481 13650
rect 9639 13608 9689 13650
rect 9852 13608 9902 13650
rect 933 13479 983 13521
rect 1146 13479 1196 13521
rect 1354 13479 1404 13521
rect 1562 13479 1612 13521
rect 1981 13475 2031 13517
rect 2194 13475 2244 13517
rect 2402 13475 2452 13517
rect 2610 13475 2660 13517
rect 19931 13602 19981 13644
rect 20139 13602 20189 13644
rect 20347 13602 20397 13644
rect 20560 13602 20610 13644
rect 11641 13473 11691 13515
rect 11854 13473 11904 13515
rect 12062 13473 12112 13515
rect 12270 13473 12320 13515
rect 12689 13469 12739 13511
rect 12902 13469 12952 13511
rect 13110 13469 13160 13511
rect 13318 13469 13368 13511
rect 30896 13606 30946 13648
rect 31104 13606 31154 13648
rect 31312 13606 31362 13648
rect 31525 13606 31575 13648
rect 22606 13477 22656 13519
rect 22819 13477 22869 13519
rect 23027 13477 23077 13519
rect 23235 13477 23285 13519
rect 23654 13473 23704 13515
rect 23867 13473 23917 13515
rect 24075 13473 24125 13515
rect 24283 13473 24333 13515
rect 41604 13600 41654 13642
rect 41812 13600 41862 13642
rect 42020 13600 42070 13642
rect 42233 13600 42283 13642
rect 33314 13471 33364 13513
rect 33527 13471 33577 13513
rect 33735 13471 33785 13513
rect 33943 13471 33993 13513
rect 34362 13467 34412 13509
rect 34575 13467 34625 13509
rect 34783 13467 34833 13509
rect 34991 13467 35041 13509
rect 8175 12933 8225 12975
rect 8383 12933 8433 12975
rect 8591 12933 8641 12975
rect 8804 12933 8854 12975
rect 933 12800 983 12842
rect 1146 12800 1196 12842
rect 1354 12800 1404 12842
rect 1562 12800 1612 12842
rect 9223 12929 9273 12971
rect 9431 12929 9481 12971
rect 9639 12929 9689 12971
rect 9852 12929 9902 12971
rect 3428 12795 3478 12837
rect 3641 12795 3691 12837
rect 3849 12795 3899 12837
rect 4057 12795 4107 12837
rect 18883 12927 18933 12969
rect 19091 12927 19141 12969
rect 19299 12927 19349 12969
rect 19512 12927 19562 12969
rect 11641 12794 11691 12836
rect 11854 12794 11904 12836
rect 12062 12794 12112 12836
rect 12270 12794 12320 12836
rect 19931 12923 19981 12965
rect 20139 12923 20189 12965
rect 20347 12923 20397 12965
rect 20560 12923 20610 12965
rect 14136 12789 14186 12831
rect 14349 12789 14399 12831
rect 14557 12789 14607 12831
rect 14765 12789 14815 12831
rect 29848 12931 29898 12973
rect 30056 12931 30106 12973
rect 30264 12931 30314 12973
rect 30477 12931 30527 12973
rect 22606 12798 22656 12840
rect 22819 12798 22869 12840
rect 23027 12798 23077 12840
rect 23235 12798 23285 12840
rect 30896 12927 30946 12969
rect 31104 12927 31154 12969
rect 31312 12927 31362 12969
rect 31525 12927 31575 12969
rect 25101 12793 25151 12835
rect 25314 12793 25364 12835
rect 25522 12793 25572 12835
rect 25730 12793 25780 12835
rect 40556 12925 40606 12967
rect 40764 12925 40814 12967
rect 40972 12925 41022 12967
rect 41185 12925 41235 12967
rect 33314 12792 33364 12834
rect 33527 12792 33577 12834
rect 33735 12792 33785 12834
rect 33943 12792 33993 12834
rect 41604 12921 41654 12963
rect 41812 12921 41862 12963
rect 42020 12921 42070 12963
rect 42233 12921 42283 12963
rect 35809 12787 35859 12829
rect 36022 12787 36072 12829
rect 36230 12787 36280 12829
rect 36438 12787 36488 12829
rect 6728 12166 6778 12208
rect 6936 12166 6986 12208
rect 7144 12166 7194 12208
rect 7357 12166 7407 12208
rect 933 12032 983 12074
rect 1146 12032 1196 12074
rect 1354 12032 1404 12074
rect 1562 12032 1612 12074
rect 9223 12161 9273 12203
rect 9431 12161 9481 12203
rect 9639 12161 9689 12203
rect 9852 12161 9902 12203
rect 1981 12028 2031 12070
rect 2194 12028 2244 12070
rect 2402 12028 2452 12070
rect 2610 12028 2660 12070
rect 17436 12160 17486 12202
rect 17644 12160 17694 12202
rect 17852 12160 17902 12202
rect 18065 12160 18115 12202
rect 11641 12026 11691 12068
rect 11854 12026 11904 12068
rect 12062 12026 12112 12068
rect 12270 12026 12320 12068
rect 19931 12155 19981 12197
rect 20139 12155 20189 12197
rect 20347 12155 20397 12197
rect 20560 12155 20610 12197
rect 12689 12022 12739 12064
rect 12902 12022 12952 12064
rect 13110 12022 13160 12064
rect 13318 12022 13368 12064
rect 28401 12164 28451 12206
rect 28609 12164 28659 12206
rect 28817 12164 28867 12206
rect 29030 12164 29080 12206
rect 22606 12030 22656 12072
rect 22819 12030 22869 12072
rect 23027 12030 23077 12072
rect 23235 12030 23285 12072
rect 30896 12159 30946 12201
rect 31104 12159 31154 12201
rect 31312 12159 31362 12201
rect 31525 12159 31575 12201
rect 23654 12026 23704 12068
rect 23867 12026 23917 12068
rect 24075 12026 24125 12068
rect 24283 12026 24333 12068
rect 39109 12158 39159 12200
rect 39317 12158 39367 12200
rect 39525 12158 39575 12200
rect 39738 12158 39788 12200
rect 33314 12024 33364 12066
rect 33527 12024 33577 12066
rect 33735 12024 33785 12066
rect 33943 12024 33993 12066
rect 41604 12153 41654 12195
rect 41812 12153 41862 12195
rect 42020 12153 42070 12195
rect 42233 12153 42283 12195
rect 34362 12020 34412 12062
rect 34575 12020 34625 12062
rect 34783 12020 34833 12062
rect 34991 12020 35041 12062
rect 8175 11486 8225 11528
rect 8383 11486 8433 11528
rect 8591 11486 8641 11528
rect 8804 11486 8854 11528
rect 933 11353 983 11395
rect 1146 11353 1196 11395
rect 1354 11353 1404 11395
rect 1562 11353 1612 11395
rect 9223 11482 9273 11524
rect 9431 11482 9481 11524
rect 9639 11482 9689 11524
rect 9852 11482 9902 11524
rect 3471 11350 3521 11392
rect 3684 11350 3734 11392
rect 3892 11350 3942 11392
rect 4100 11350 4150 11392
rect 18883 11480 18933 11522
rect 19091 11480 19141 11522
rect 19299 11480 19349 11522
rect 19512 11480 19562 11522
rect 11641 11347 11691 11389
rect 11854 11347 11904 11389
rect 12062 11347 12112 11389
rect 12270 11347 12320 11389
rect 19931 11476 19981 11518
rect 20139 11476 20189 11518
rect 20347 11476 20397 11518
rect 20560 11476 20610 11518
rect 14179 11344 14229 11386
rect 14392 11344 14442 11386
rect 14600 11344 14650 11386
rect 14808 11344 14858 11386
rect 29848 11484 29898 11526
rect 30056 11484 30106 11526
rect 30264 11484 30314 11526
rect 30477 11484 30527 11526
rect 22606 11351 22656 11393
rect 22819 11351 22869 11393
rect 23027 11351 23077 11393
rect 23235 11351 23285 11393
rect 30896 11480 30946 11522
rect 31104 11480 31154 11522
rect 31312 11480 31362 11522
rect 31525 11480 31575 11522
rect 25144 11348 25194 11390
rect 25357 11348 25407 11390
rect 25565 11348 25615 11390
rect 25773 11348 25823 11390
rect 40556 11478 40606 11520
rect 40764 11478 40814 11520
rect 40972 11478 41022 11520
rect 41185 11478 41235 11520
rect 33314 11345 33364 11387
rect 33527 11345 33577 11387
rect 33735 11345 33785 11387
rect 33943 11345 33993 11387
rect 41604 11474 41654 11516
rect 41812 11474 41862 11516
rect 42020 11474 42070 11516
rect 42233 11474 42283 11516
rect 35852 11342 35902 11384
rect 36065 11342 36115 11384
rect 36273 11342 36323 11384
rect 36481 11342 36531 11384
rect 6686 10644 6736 10686
rect 6894 10644 6944 10686
rect 7102 10644 7152 10686
rect 7315 10644 7365 10686
rect 934 10512 984 10554
rect 1147 10512 1197 10554
rect 1355 10512 1405 10554
rect 1563 10512 1613 10554
rect 9224 10641 9274 10683
rect 9432 10641 9482 10683
rect 9640 10641 9690 10683
rect 9853 10641 9903 10683
rect 1982 10508 2032 10550
rect 2195 10508 2245 10550
rect 2403 10508 2453 10550
rect 2611 10508 2661 10550
rect 17394 10638 17444 10680
rect 17602 10638 17652 10680
rect 17810 10638 17860 10680
rect 18023 10638 18073 10680
rect 11642 10506 11692 10548
rect 11855 10506 11905 10548
rect 12063 10506 12113 10548
rect 12271 10506 12321 10548
rect 19932 10635 19982 10677
rect 20140 10635 20190 10677
rect 20348 10635 20398 10677
rect 20561 10635 20611 10677
rect 12690 10502 12740 10544
rect 12903 10502 12953 10544
rect 13111 10502 13161 10544
rect 13319 10502 13369 10544
rect 28359 10642 28409 10684
rect 28567 10642 28617 10684
rect 28775 10642 28825 10684
rect 28988 10642 29038 10684
rect 22607 10510 22657 10552
rect 22820 10510 22870 10552
rect 23028 10510 23078 10552
rect 23236 10510 23286 10552
rect 30897 10639 30947 10681
rect 31105 10639 31155 10681
rect 31313 10639 31363 10681
rect 31526 10639 31576 10681
rect 23655 10506 23705 10548
rect 23868 10506 23918 10548
rect 24076 10506 24126 10548
rect 24284 10506 24334 10548
rect 39067 10636 39117 10678
rect 39275 10636 39325 10678
rect 39483 10636 39533 10678
rect 39696 10636 39746 10678
rect 33315 10504 33365 10546
rect 33528 10504 33578 10546
rect 33736 10504 33786 10546
rect 33944 10504 33994 10546
rect 41605 10633 41655 10675
rect 41813 10633 41863 10675
rect 42021 10633 42071 10675
rect 42234 10633 42284 10675
rect 34363 10500 34413 10542
rect 34576 10500 34626 10542
rect 34784 10500 34834 10542
rect 34992 10500 35042 10542
rect 8176 9966 8226 10008
rect 8384 9966 8434 10008
rect 8592 9966 8642 10008
rect 8805 9966 8855 10008
rect 934 9833 984 9875
rect 1147 9833 1197 9875
rect 1355 9833 1405 9875
rect 1563 9833 1613 9875
rect 9224 9962 9274 10004
rect 9432 9962 9482 10004
rect 9640 9962 9690 10004
rect 9853 9962 9903 10004
rect 3429 9828 3479 9870
rect 3642 9828 3692 9870
rect 3850 9828 3900 9870
rect 4058 9828 4108 9870
rect 18884 9960 18934 10002
rect 19092 9960 19142 10002
rect 19300 9960 19350 10002
rect 19513 9960 19563 10002
rect 11642 9827 11692 9869
rect 11855 9827 11905 9869
rect 12063 9827 12113 9869
rect 12271 9827 12321 9869
rect 19932 9956 19982 9998
rect 20140 9956 20190 9998
rect 20348 9956 20398 9998
rect 20561 9956 20611 9998
rect 14137 9822 14187 9864
rect 14350 9822 14400 9864
rect 14558 9822 14608 9864
rect 14766 9822 14816 9864
rect 29849 9964 29899 10006
rect 30057 9964 30107 10006
rect 30265 9964 30315 10006
rect 30478 9964 30528 10006
rect 22607 9831 22657 9873
rect 22820 9831 22870 9873
rect 23028 9831 23078 9873
rect 23236 9831 23286 9873
rect 30897 9960 30947 10002
rect 31105 9960 31155 10002
rect 31313 9960 31363 10002
rect 31526 9960 31576 10002
rect 25102 9826 25152 9868
rect 25315 9826 25365 9868
rect 25523 9826 25573 9868
rect 25731 9826 25781 9868
rect 40557 9958 40607 10000
rect 40765 9958 40815 10000
rect 40973 9958 41023 10000
rect 41186 9958 41236 10000
rect 33315 9825 33365 9867
rect 33528 9825 33578 9867
rect 33736 9825 33786 9867
rect 33944 9825 33994 9867
rect 41605 9954 41655 9996
rect 41813 9954 41863 9996
rect 42021 9954 42071 9996
rect 42234 9954 42284 9996
rect 35810 9820 35860 9862
rect 36023 9820 36073 9862
rect 36231 9820 36281 9862
rect 36439 9820 36489 9862
rect 6729 9199 6779 9241
rect 6937 9199 6987 9241
rect 7145 9199 7195 9241
rect 7358 9199 7408 9241
rect 934 9065 984 9107
rect 1147 9065 1197 9107
rect 1355 9065 1405 9107
rect 1563 9065 1613 9107
rect 9224 9194 9274 9236
rect 9432 9194 9482 9236
rect 9640 9194 9690 9236
rect 9853 9194 9903 9236
rect 1982 9061 2032 9103
rect 2195 9061 2245 9103
rect 2403 9061 2453 9103
rect 2611 9061 2661 9103
rect 17437 9193 17487 9235
rect 17645 9193 17695 9235
rect 17853 9193 17903 9235
rect 18066 9193 18116 9235
rect 11642 9059 11692 9101
rect 11855 9059 11905 9101
rect 12063 9059 12113 9101
rect 12271 9059 12321 9101
rect 19932 9188 19982 9230
rect 20140 9188 20190 9230
rect 20348 9188 20398 9230
rect 20561 9188 20611 9230
rect 12690 9055 12740 9097
rect 12903 9055 12953 9097
rect 13111 9055 13161 9097
rect 13319 9055 13369 9097
rect 28402 9197 28452 9239
rect 28610 9197 28660 9239
rect 28818 9197 28868 9239
rect 29031 9197 29081 9239
rect 22607 9063 22657 9105
rect 22820 9063 22870 9105
rect 23028 9063 23078 9105
rect 23236 9063 23286 9105
rect 30897 9192 30947 9234
rect 31105 9192 31155 9234
rect 31313 9192 31363 9234
rect 31526 9192 31576 9234
rect 23655 9059 23705 9101
rect 23868 9059 23918 9101
rect 24076 9059 24126 9101
rect 24284 9059 24334 9101
rect 39110 9191 39160 9233
rect 39318 9191 39368 9233
rect 39526 9191 39576 9233
rect 39739 9191 39789 9233
rect 33315 9057 33365 9099
rect 33528 9057 33578 9099
rect 33736 9057 33786 9099
rect 33944 9057 33994 9099
rect 41605 9186 41655 9228
rect 41813 9186 41863 9228
rect 42021 9186 42071 9228
rect 42234 9186 42284 9228
rect 34363 9053 34413 9095
rect 34576 9053 34626 9095
rect 34784 9053 34834 9095
rect 34992 9053 35042 9095
rect 8176 8519 8226 8561
rect 8384 8519 8434 8561
rect 8592 8519 8642 8561
rect 8805 8519 8855 8561
rect 934 8386 984 8428
rect 1147 8386 1197 8428
rect 1355 8386 1405 8428
rect 1563 8386 1613 8428
rect 9224 8515 9274 8557
rect 9432 8515 9482 8557
rect 9640 8515 9690 8557
rect 9853 8515 9903 8557
rect 4537 8377 4587 8419
rect 4750 8377 4800 8419
rect 4958 8377 5008 8419
rect 5166 8377 5216 8419
rect 18884 8513 18934 8555
rect 19092 8513 19142 8555
rect 19300 8513 19350 8555
rect 19513 8513 19563 8555
rect 11642 8380 11692 8422
rect 11855 8380 11905 8422
rect 12063 8380 12113 8422
rect 12271 8380 12321 8422
rect 19932 8509 19982 8551
rect 20140 8509 20190 8551
rect 20348 8509 20398 8551
rect 20561 8509 20611 8551
rect 15245 8371 15295 8413
rect 15458 8371 15508 8413
rect 15666 8371 15716 8413
rect 15874 8371 15924 8413
rect 29849 8517 29899 8559
rect 30057 8517 30107 8559
rect 30265 8517 30315 8559
rect 30478 8517 30528 8559
rect 22607 8384 22657 8426
rect 22820 8384 22870 8426
rect 23028 8384 23078 8426
rect 23236 8384 23286 8426
rect 30897 8513 30947 8555
rect 31105 8513 31155 8555
rect 31313 8513 31363 8555
rect 31526 8513 31576 8555
rect 26210 8375 26260 8417
rect 26423 8375 26473 8417
rect 26631 8375 26681 8417
rect 26839 8375 26889 8417
rect 40557 8511 40607 8553
rect 40765 8511 40815 8553
rect 40973 8511 41023 8553
rect 41186 8511 41236 8553
rect 33315 8378 33365 8420
rect 33528 8378 33578 8420
rect 33736 8378 33786 8420
rect 33944 8378 33994 8420
rect 41605 8507 41655 8549
rect 41813 8507 41863 8549
rect 42021 8507 42071 8549
rect 42234 8507 42284 8549
rect 36918 8369 36968 8411
rect 37131 8369 37181 8411
rect 37339 8369 37389 8411
rect 37547 8369 37597 8411
rect 5618 7609 5668 7651
rect 5826 7609 5876 7651
rect 6034 7609 6084 7651
rect 6247 7609 6297 7651
rect 931 7471 981 7513
rect 1144 7471 1194 7513
rect 1352 7471 1402 7513
rect 1560 7471 1610 7513
rect 9221 7600 9271 7642
rect 9429 7600 9479 7642
rect 9637 7600 9687 7642
rect 9850 7600 9900 7642
rect 1979 7467 2029 7509
rect 2192 7467 2242 7509
rect 2400 7467 2450 7509
rect 2608 7467 2658 7509
rect 16326 7603 16376 7645
rect 16534 7603 16584 7645
rect 16742 7603 16792 7645
rect 16955 7603 17005 7645
rect 11639 7465 11689 7507
rect 11852 7465 11902 7507
rect 12060 7465 12110 7507
rect 12268 7465 12318 7507
rect 19929 7594 19979 7636
rect 20137 7594 20187 7636
rect 20345 7594 20395 7636
rect 20558 7594 20608 7636
rect 12687 7461 12737 7503
rect 12900 7461 12950 7503
rect 13108 7461 13158 7503
rect 13316 7461 13366 7503
rect 27291 7607 27341 7649
rect 27499 7607 27549 7649
rect 27707 7607 27757 7649
rect 27920 7607 27970 7649
rect 22604 7469 22654 7511
rect 22817 7469 22867 7511
rect 23025 7469 23075 7511
rect 23233 7469 23283 7511
rect 30894 7598 30944 7640
rect 31102 7598 31152 7640
rect 31310 7598 31360 7640
rect 31523 7598 31573 7640
rect 23652 7465 23702 7507
rect 23865 7465 23915 7507
rect 24073 7465 24123 7507
rect 24281 7465 24331 7507
rect 37999 7601 38049 7643
rect 38207 7601 38257 7643
rect 38415 7601 38465 7643
rect 38628 7601 38678 7643
rect 33312 7463 33362 7505
rect 33525 7463 33575 7505
rect 33733 7463 33783 7505
rect 33941 7463 33991 7505
rect 41602 7592 41652 7634
rect 41810 7592 41860 7634
rect 42018 7592 42068 7634
rect 42231 7592 42281 7634
rect 34360 7459 34410 7501
rect 34573 7459 34623 7501
rect 34781 7459 34831 7501
rect 34989 7459 35039 7501
rect 8173 6925 8223 6967
rect 8381 6925 8431 6967
rect 8589 6925 8639 6967
rect 8802 6925 8852 6967
rect 931 6792 981 6834
rect 1144 6792 1194 6834
rect 1352 6792 1402 6834
rect 1560 6792 1610 6834
rect 9221 6921 9271 6963
rect 9429 6921 9479 6963
rect 9637 6921 9687 6963
rect 9850 6921 9900 6963
rect 3426 6787 3476 6829
rect 3639 6787 3689 6829
rect 3847 6787 3897 6829
rect 4055 6787 4105 6829
rect 18881 6919 18931 6961
rect 19089 6919 19139 6961
rect 19297 6919 19347 6961
rect 19510 6919 19560 6961
rect 11639 6786 11689 6828
rect 11852 6786 11902 6828
rect 12060 6786 12110 6828
rect 12268 6786 12318 6828
rect 19929 6915 19979 6957
rect 20137 6915 20187 6957
rect 20345 6915 20395 6957
rect 20558 6915 20608 6957
rect 14134 6781 14184 6823
rect 14347 6781 14397 6823
rect 14555 6781 14605 6823
rect 14763 6781 14813 6823
rect 29846 6923 29896 6965
rect 30054 6923 30104 6965
rect 30262 6923 30312 6965
rect 30475 6923 30525 6965
rect 22604 6790 22654 6832
rect 22817 6790 22867 6832
rect 23025 6790 23075 6832
rect 23233 6790 23283 6832
rect 30894 6919 30944 6961
rect 31102 6919 31152 6961
rect 31310 6919 31360 6961
rect 31523 6919 31573 6961
rect 25099 6785 25149 6827
rect 25312 6785 25362 6827
rect 25520 6785 25570 6827
rect 25728 6785 25778 6827
rect 40554 6917 40604 6959
rect 40762 6917 40812 6959
rect 40970 6917 41020 6959
rect 41183 6917 41233 6959
rect 33312 6784 33362 6826
rect 33525 6784 33575 6826
rect 33733 6784 33783 6826
rect 33941 6784 33991 6826
rect 41602 6913 41652 6955
rect 41810 6913 41860 6955
rect 42018 6913 42068 6955
rect 42231 6913 42281 6955
rect 35807 6779 35857 6821
rect 36020 6779 36070 6821
rect 36228 6779 36278 6821
rect 36436 6779 36486 6821
rect 6726 6158 6776 6200
rect 6934 6158 6984 6200
rect 7142 6158 7192 6200
rect 7355 6158 7405 6200
rect 931 6024 981 6066
rect 1144 6024 1194 6066
rect 1352 6024 1402 6066
rect 1560 6024 1610 6066
rect 9221 6153 9271 6195
rect 9429 6153 9479 6195
rect 9637 6153 9687 6195
rect 9850 6153 9900 6195
rect 1979 6020 2029 6062
rect 2192 6020 2242 6062
rect 2400 6020 2450 6062
rect 2608 6020 2658 6062
rect 17434 6152 17484 6194
rect 17642 6152 17692 6194
rect 17850 6152 17900 6194
rect 18063 6152 18113 6194
rect 11639 6018 11689 6060
rect 11852 6018 11902 6060
rect 12060 6018 12110 6060
rect 12268 6018 12318 6060
rect 19929 6147 19979 6189
rect 20137 6147 20187 6189
rect 20345 6147 20395 6189
rect 20558 6147 20608 6189
rect 12687 6014 12737 6056
rect 12900 6014 12950 6056
rect 13108 6014 13158 6056
rect 13316 6014 13366 6056
rect 28399 6156 28449 6198
rect 28607 6156 28657 6198
rect 28815 6156 28865 6198
rect 29028 6156 29078 6198
rect 22604 6022 22654 6064
rect 22817 6022 22867 6064
rect 23025 6022 23075 6064
rect 23233 6022 23283 6064
rect 30894 6151 30944 6193
rect 31102 6151 31152 6193
rect 31310 6151 31360 6193
rect 31523 6151 31573 6193
rect 23652 6018 23702 6060
rect 23865 6018 23915 6060
rect 24073 6018 24123 6060
rect 24281 6018 24331 6060
rect 39107 6150 39157 6192
rect 39315 6150 39365 6192
rect 39523 6150 39573 6192
rect 39736 6150 39786 6192
rect 33312 6016 33362 6058
rect 33525 6016 33575 6058
rect 33733 6016 33783 6058
rect 33941 6016 33991 6058
rect 41602 6145 41652 6187
rect 41810 6145 41860 6187
rect 42018 6145 42068 6187
rect 42231 6145 42281 6187
rect 34360 6012 34410 6054
rect 34573 6012 34623 6054
rect 34781 6012 34831 6054
rect 34989 6012 35039 6054
rect 8173 5478 8223 5520
rect 8381 5478 8431 5520
rect 8589 5478 8639 5520
rect 8802 5478 8852 5520
rect 931 5345 981 5387
rect 1144 5345 1194 5387
rect 1352 5345 1402 5387
rect 1560 5345 1610 5387
rect 9221 5474 9271 5516
rect 9429 5474 9479 5516
rect 9637 5474 9687 5516
rect 9850 5474 9900 5516
rect 3469 5342 3519 5384
rect 3682 5342 3732 5384
rect 3890 5342 3940 5384
rect 4098 5342 4148 5384
rect 18881 5472 18931 5514
rect 19089 5472 19139 5514
rect 19297 5472 19347 5514
rect 19510 5472 19560 5514
rect 11639 5339 11689 5381
rect 11852 5339 11902 5381
rect 12060 5339 12110 5381
rect 12268 5339 12318 5381
rect 19929 5468 19979 5510
rect 20137 5468 20187 5510
rect 20345 5468 20395 5510
rect 20558 5468 20608 5510
rect 14177 5336 14227 5378
rect 14390 5336 14440 5378
rect 14598 5336 14648 5378
rect 14806 5336 14856 5378
rect 29846 5476 29896 5518
rect 30054 5476 30104 5518
rect 30262 5476 30312 5518
rect 30475 5476 30525 5518
rect 22604 5343 22654 5385
rect 22817 5343 22867 5385
rect 23025 5343 23075 5385
rect 23233 5343 23283 5385
rect 30894 5472 30944 5514
rect 31102 5472 31152 5514
rect 31310 5472 31360 5514
rect 31523 5472 31573 5514
rect 25142 5340 25192 5382
rect 25355 5340 25405 5382
rect 25563 5340 25613 5382
rect 25771 5340 25821 5382
rect 40554 5470 40604 5512
rect 40762 5470 40812 5512
rect 40970 5470 41020 5512
rect 41183 5470 41233 5512
rect 33312 5337 33362 5379
rect 33525 5337 33575 5379
rect 33733 5337 33783 5379
rect 33941 5337 33991 5379
rect 41602 5466 41652 5508
rect 41810 5466 41860 5508
rect 42018 5466 42068 5508
rect 42231 5466 42281 5508
rect 35850 5334 35900 5376
rect 36063 5334 36113 5376
rect 36271 5334 36321 5376
rect 36479 5334 36529 5376
rect 6684 4636 6734 4678
rect 6892 4636 6942 4678
rect 7100 4636 7150 4678
rect 7313 4636 7363 4678
rect 932 4504 982 4546
rect 1145 4504 1195 4546
rect 1353 4504 1403 4546
rect 1561 4504 1611 4546
rect 9222 4633 9272 4675
rect 9430 4633 9480 4675
rect 9638 4633 9688 4675
rect 9851 4633 9901 4675
rect 1980 4500 2030 4542
rect 2193 4500 2243 4542
rect 2401 4500 2451 4542
rect 2609 4500 2659 4542
rect 4882 4506 4932 4548
rect 5095 4506 5145 4548
rect 5303 4506 5353 4548
rect 5511 4506 5561 4548
rect 17392 4630 17442 4672
rect 17600 4630 17650 4672
rect 17808 4630 17858 4672
rect 18021 4630 18071 4672
rect 11640 4498 11690 4540
rect 11853 4498 11903 4540
rect 12061 4498 12111 4540
rect 12269 4498 12319 4540
rect 19930 4627 19980 4669
rect 20138 4627 20188 4669
rect 20346 4627 20396 4669
rect 20559 4627 20609 4669
rect 12688 4494 12738 4536
rect 12901 4494 12951 4536
rect 13109 4494 13159 4536
rect 13317 4494 13367 4536
rect 15590 4500 15640 4542
rect 15803 4500 15853 4542
rect 16011 4500 16061 4542
rect 16219 4500 16269 4542
rect 28357 4634 28407 4676
rect 28565 4634 28615 4676
rect 28773 4634 28823 4676
rect 28986 4634 29036 4676
rect 22605 4502 22655 4544
rect 22818 4502 22868 4544
rect 23026 4502 23076 4544
rect 23234 4502 23284 4544
rect 30895 4631 30945 4673
rect 31103 4631 31153 4673
rect 31311 4631 31361 4673
rect 31524 4631 31574 4673
rect 23653 4498 23703 4540
rect 23866 4498 23916 4540
rect 24074 4498 24124 4540
rect 24282 4498 24332 4540
rect 26555 4504 26605 4546
rect 26768 4504 26818 4546
rect 26976 4504 27026 4546
rect 27184 4504 27234 4546
rect 39065 4628 39115 4670
rect 39273 4628 39323 4670
rect 39481 4628 39531 4670
rect 39694 4628 39744 4670
rect 33313 4496 33363 4538
rect 33526 4496 33576 4538
rect 33734 4496 33784 4538
rect 33942 4496 33992 4538
rect 41603 4625 41653 4667
rect 41811 4625 41861 4667
rect 42019 4625 42069 4667
rect 42232 4625 42282 4667
rect 34361 4492 34411 4534
rect 34574 4492 34624 4534
rect 34782 4492 34832 4534
rect 34990 4492 35040 4534
rect 37263 4498 37313 4540
rect 37476 4498 37526 4540
rect 37684 4498 37734 4540
rect 37892 4498 37942 4540
rect 8174 3958 8224 4000
rect 8382 3958 8432 4000
rect 8590 3958 8640 4000
rect 8803 3958 8853 4000
rect 932 3825 982 3867
rect 1145 3825 1195 3867
rect 1353 3825 1403 3867
rect 1561 3825 1611 3867
rect 9222 3954 9272 3996
rect 9430 3954 9480 3996
rect 9638 3954 9688 3996
rect 9851 3954 9901 3996
rect 3427 3820 3477 3862
rect 3640 3820 3690 3862
rect 3848 3820 3898 3862
rect 4056 3820 4106 3862
rect 18882 3952 18932 3994
rect 19090 3952 19140 3994
rect 19298 3952 19348 3994
rect 19511 3952 19561 3994
rect 11640 3819 11690 3861
rect 11853 3819 11903 3861
rect 12061 3819 12111 3861
rect 12269 3819 12319 3861
rect 19930 3948 19980 3990
rect 20138 3948 20188 3990
rect 20346 3948 20396 3990
rect 20559 3948 20609 3990
rect 14135 3814 14185 3856
rect 14348 3814 14398 3856
rect 14556 3814 14606 3856
rect 14764 3814 14814 3856
rect 29847 3956 29897 3998
rect 30055 3956 30105 3998
rect 30263 3956 30313 3998
rect 30476 3956 30526 3998
rect 22605 3823 22655 3865
rect 22818 3823 22868 3865
rect 23026 3823 23076 3865
rect 23234 3823 23284 3865
rect 30895 3952 30945 3994
rect 31103 3952 31153 3994
rect 31311 3952 31361 3994
rect 31524 3952 31574 3994
rect 25100 3818 25150 3860
rect 25313 3818 25363 3860
rect 25521 3818 25571 3860
rect 25729 3818 25779 3860
rect 40555 3950 40605 3992
rect 40763 3950 40813 3992
rect 40971 3950 41021 3992
rect 41184 3950 41234 3992
rect 33313 3817 33363 3859
rect 33526 3817 33576 3859
rect 33734 3817 33784 3859
rect 33942 3817 33992 3859
rect 41603 3946 41653 3988
rect 41811 3946 41861 3988
rect 42019 3946 42069 3988
rect 42232 3946 42282 3988
rect 35808 3812 35858 3854
rect 36021 3812 36071 3854
rect 36229 3812 36279 3854
rect 36437 3812 36487 3854
rect 6727 3191 6777 3233
rect 6935 3191 6985 3233
rect 7143 3191 7193 3233
rect 7356 3191 7406 3233
rect 932 3057 982 3099
rect 1145 3057 1195 3099
rect 1353 3057 1403 3099
rect 1561 3057 1611 3099
rect 9222 3186 9272 3228
rect 9430 3186 9480 3228
rect 9638 3186 9688 3228
rect 9851 3186 9901 3228
rect 1980 3053 2030 3095
rect 2193 3053 2243 3095
rect 2401 3053 2451 3095
rect 2609 3053 2659 3095
rect 17435 3185 17485 3227
rect 17643 3185 17693 3227
rect 17851 3185 17901 3227
rect 18064 3185 18114 3227
rect 11640 3051 11690 3093
rect 11853 3051 11903 3093
rect 12061 3051 12111 3093
rect 12269 3051 12319 3093
rect 19930 3180 19980 3222
rect 20138 3180 20188 3222
rect 20346 3180 20396 3222
rect 20559 3180 20609 3222
rect 12688 3047 12738 3089
rect 12901 3047 12951 3089
rect 13109 3047 13159 3089
rect 13317 3047 13367 3089
rect 28400 3189 28450 3231
rect 28608 3189 28658 3231
rect 28816 3189 28866 3231
rect 29029 3189 29079 3231
rect 22605 3055 22655 3097
rect 22818 3055 22868 3097
rect 23026 3055 23076 3097
rect 23234 3055 23284 3097
rect 30895 3184 30945 3226
rect 31103 3184 31153 3226
rect 31311 3184 31361 3226
rect 31524 3184 31574 3226
rect 23653 3051 23703 3093
rect 23866 3051 23916 3093
rect 24074 3051 24124 3093
rect 24282 3051 24332 3093
rect 39108 3183 39158 3225
rect 39316 3183 39366 3225
rect 39524 3183 39574 3225
rect 39737 3183 39787 3225
rect 33313 3049 33363 3091
rect 33526 3049 33576 3091
rect 33734 3049 33784 3091
rect 33942 3049 33992 3091
rect 41603 3178 41653 3220
rect 41811 3178 41861 3220
rect 42019 3178 42069 3220
rect 42232 3178 42282 3220
rect 34361 3045 34411 3087
rect 34574 3045 34624 3087
rect 34782 3045 34832 3087
rect 34990 3045 35040 3087
rect 8174 2511 8224 2553
rect 8382 2511 8432 2553
rect 8590 2511 8640 2553
rect 8803 2511 8853 2553
rect 9222 2507 9272 2549
rect 9430 2507 9480 2549
rect 9638 2507 9688 2549
rect 9851 2507 9901 2549
rect 932 2378 982 2420
rect 1145 2378 1195 2420
rect 1353 2378 1403 2420
rect 1561 2378 1611 2420
rect 18882 2505 18932 2547
rect 19090 2505 19140 2547
rect 19298 2505 19348 2547
rect 19511 2505 19561 2547
rect 19930 2501 19980 2543
rect 20138 2501 20188 2543
rect 20346 2501 20396 2543
rect 20559 2501 20609 2543
rect 11640 2372 11690 2414
rect 11853 2372 11903 2414
rect 12061 2372 12111 2414
rect 12269 2372 12319 2414
rect 29847 2509 29897 2551
rect 30055 2509 30105 2551
rect 30263 2509 30313 2551
rect 30476 2509 30526 2551
rect 30895 2505 30945 2547
rect 31103 2505 31153 2547
rect 31311 2505 31361 2547
rect 31524 2505 31574 2547
rect 22605 2376 22655 2418
rect 22818 2376 22868 2418
rect 23026 2376 23076 2418
rect 23234 2376 23284 2418
rect 40555 2503 40605 2545
rect 40763 2503 40813 2545
rect 40971 2503 41021 2545
rect 41184 2503 41234 2545
rect 41603 2499 41653 2541
rect 41811 2499 41861 2541
rect 42019 2499 42069 2541
rect 42232 2499 42282 2541
rect 33313 2370 33363 2412
rect 33526 2370 33576 2412
rect 33734 2370 33784 2412
rect 33942 2370 33992 2412
rect 10643 219 10693 261
rect 10856 219 10906 261
rect 11064 219 11114 261
rect 11272 219 11322 261
rect 21280 206 21330 248
rect 21493 206 21543 248
rect 21701 206 21751 248
rect 21909 206 21959 248
rect 32316 217 32366 259
rect 32529 217 32579 259
rect 32737 217 32787 259
rect 32945 217 32995 259
<< pmos >>
rect 933 13598 983 13698
rect 1146 13598 1196 13698
rect 1354 13598 1404 13698
rect 1562 13598 1612 13698
rect 1981 13594 2031 13694
rect 2194 13594 2244 13694
rect 2402 13594 2452 13694
rect 2610 13594 2660 13694
rect 11641 13592 11691 13692
rect 11854 13592 11904 13692
rect 12062 13592 12112 13692
rect 12270 13592 12320 13692
rect 9223 13431 9273 13531
rect 9431 13431 9481 13531
rect 9639 13431 9689 13531
rect 9852 13431 9902 13531
rect 12689 13588 12739 13688
rect 12902 13588 12952 13688
rect 13110 13588 13160 13688
rect 13318 13588 13368 13688
rect 22606 13596 22656 13696
rect 22819 13596 22869 13696
rect 23027 13596 23077 13696
rect 23235 13596 23285 13696
rect 19931 13425 19981 13525
rect 20139 13425 20189 13525
rect 20347 13425 20397 13525
rect 20560 13425 20610 13525
rect 23654 13592 23704 13692
rect 23867 13592 23917 13692
rect 24075 13592 24125 13692
rect 24283 13592 24333 13692
rect 33314 13590 33364 13690
rect 33527 13590 33577 13690
rect 33735 13590 33785 13690
rect 33943 13590 33993 13690
rect 30896 13429 30946 13529
rect 31104 13429 31154 13529
rect 31312 13429 31362 13529
rect 31525 13429 31575 13529
rect 34362 13586 34412 13686
rect 34575 13586 34625 13686
rect 34783 13586 34833 13686
rect 34991 13586 35041 13686
rect 41604 13423 41654 13523
rect 41812 13423 41862 13523
rect 42020 13423 42070 13523
rect 42233 13423 42283 13523
rect 933 12919 983 13019
rect 1146 12919 1196 13019
rect 1354 12919 1404 13019
rect 1562 12919 1612 13019
rect 3428 12914 3478 13014
rect 3641 12914 3691 13014
rect 3849 12914 3899 13014
rect 4057 12914 4107 13014
rect 8175 12756 8225 12856
rect 8383 12756 8433 12856
rect 8591 12756 8641 12856
rect 8804 12756 8854 12856
rect 11641 12913 11691 13013
rect 11854 12913 11904 13013
rect 12062 12913 12112 13013
rect 12270 12913 12320 13013
rect 9223 12752 9273 12852
rect 9431 12752 9481 12852
rect 9639 12752 9689 12852
rect 9852 12752 9902 12852
rect 14136 12908 14186 13008
rect 14349 12908 14399 13008
rect 14557 12908 14607 13008
rect 14765 12908 14815 13008
rect 18883 12750 18933 12850
rect 19091 12750 19141 12850
rect 19299 12750 19349 12850
rect 19512 12750 19562 12850
rect 22606 12917 22656 13017
rect 22819 12917 22869 13017
rect 23027 12917 23077 13017
rect 23235 12917 23285 13017
rect 19931 12746 19981 12846
rect 20139 12746 20189 12846
rect 20347 12746 20397 12846
rect 20560 12746 20610 12846
rect 25101 12912 25151 13012
rect 25314 12912 25364 13012
rect 25522 12912 25572 13012
rect 25730 12912 25780 13012
rect 29848 12754 29898 12854
rect 30056 12754 30106 12854
rect 30264 12754 30314 12854
rect 30477 12754 30527 12854
rect 33314 12911 33364 13011
rect 33527 12911 33577 13011
rect 33735 12911 33785 13011
rect 33943 12911 33993 13011
rect 30896 12750 30946 12850
rect 31104 12750 31154 12850
rect 31312 12750 31362 12850
rect 31525 12750 31575 12850
rect 35809 12906 35859 13006
rect 36022 12906 36072 13006
rect 36230 12906 36280 13006
rect 36438 12906 36488 13006
rect 40556 12748 40606 12848
rect 40764 12748 40814 12848
rect 40972 12748 41022 12848
rect 41185 12748 41235 12848
rect 41604 12744 41654 12844
rect 41812 12744 41862 12844
rect 42020 12744 42070 12844
rect 42233 12744 42283 12844
rect 933 12151 983 12251
rect 1146 12151 1196 12251
rect 1354 12151 1404 12251
rect 1562 12151 1612 12251
rect 1981 12147 2031 12247
rect 2194 12147 2244 12247
rect 2402 12147 2452 12247
rect 2610 12147 2660 12247
rect 6728 11989 6778 12089
rect 6936 11989 6986 12089
rect 7144 11989 7194 12089
rect 7357 11989 7407 12089
rect 11641 12145 11691 12245
rect 11854 12145 11904 12245
rect 12062 12145 12112 12245
rect 12270 12145 12320 12245
rect 9223 11984 9273 12084
rect 9431 11984 9481 12084
rect 9639 11984 9689 12084
rect 9852 11984 9902 12084
rect 12689 12141 12739 12241
rect 12902 12141 12952 12241
rect 13110 12141 13160 12241
rect 13318 12141 13368 12241
rect 17436 11983 17486 12083
rect 17644 11983 17694 12083
rect 17852 11983 17902 12083
rect 18065 11983 18115 12083
rect 22606 12149 22656 12249
rect 22819 12149 22869 12249
rect 23027 12149 23077 12249
rect 23235 12149 23285 12249
rect 19931 11978 19981 12078
rect 20139 11978 20189 12078
rect 20347 11978 20397 12078
rect 20560 11978 20610 12078
rect 23654 12145 23704 12245
rect 23867 12145 23917 12245
rect 24075 12145 24125 12245
rect 24283 12145 24333 12245
rect 28401 11987 28451 12087
rect 28609 11987 28659 12087
rect 28817 11987 28867 12087
rect 29030 11987 29080 12087
rect 33314 12143 33364 12243
rect 33527 12143 33577 12243
rect 33735 12143 33785 12243
rect 33943 12143 33993 12243
rect 30896 11982 30946 12082
rect 31104 11982 31154 12082
rect 31312 11982 31362 12082
rect 31525 11982 31575 12082
rect 34362 12139 34412 12239
rect 34575 12139 34625 12239
rect 34783 12139 34833 12239
rect 34991 12139 35041 12239
rect 39109 11981 39159 12081
rect 39317 11981 39367 12081
rect 39525 11981 39575 12081
rect 39738 11981 39788 12081
rect 41604 11976 41654 12076
rect 41812 11976 41862 12076
rect 42020 11976 42070 12076
rect 42233 11976 42283 12076
rect 933 11472 983 11572
rect 1146 11472 1196 11572
rect 1354 11472 1404 11572
rect 1562 11472 1612 11572
rect 3471 11469 3521 11569
rect 3684 11469 3734 11569
rect 3892 11469 3942 11569
rect 4100 11469 4150 11569
rect 8175 11309 8225 11409
rect 8383 11309 8433 11409
rect 8591 11309 8641 11409
rect 8804 11309 8854 11409
rect 11641 11466 11691 11566
rect 11854 11466 11904 11566
rect 12062 11466 12112 11566
rect 12270 11466 12320 11566
rect 9223 11305 9273 11405
rect 9431 11305 9481 11405
rect 9639 11305 9689 11405
rect 9852 11305 9902 11405
rect 14179 11463 14229 11563
rect 14392 11463 14442 11563
rect 14600 11463 14650 11563
rect 14808 11463 14858 11563
rect 18883 11303 18933 11403
rect 19091 11303 19141 11403
rect 19299 11303 19349 11403
rect 19512 11303 19562 11403
rect 22606 11470 22656 11570
rect 22819 11470 22869 11570
rect 23027 11470 23077 11570
rect 23235 11470 23285 11570
rect 19931 11299 19981 11399
rect 20139 11299 20189 11399
rect 20347 11299 20397 11399
rect 20560 11299 20610 11399
rect 25144 11467 25194 11567
rect 25357 11467 25407 11567
rect 25565 11467 25615 11567
rect 25773 11467 25823 11567
rect 29848 11307 29898 11407
rect 30056 11307 30106 11407
rect 30264 11307 30314 11407
rect 30477 11307 30527 11407
rect 33314 11464 33364 11564
rect 33527 11464 33577 11564
rect 33735 11464 33785 11564
rect 33943 11464 33993 11564
rect 30896 11303 30946 11403
rect 31104 11303 31154 11403
rect 31312 11303 31362 11403
rect 31525 11303 31575 11403
rect 35852 11461 35902 11561
rect 36065 11461 36115 11561
rect 36273 11461 36323 11561
rect 36481 11461 36531 11561
rect 40556 11301 40606 11401
rect 40764 11301 40814 11401
rect 40972 11301 41022 11401
rect 41185 11301 41235 11401
rect 41604 11297 41654 11397
rect 41812 11297 41862 11397
rect 42020 11297 42070 11397
rect 42233 11297 42283 11397
rect 934 10631 984 10731
rect 1147 10631 1197 10731
rect 1355 10631 1405 10731
rect 1563 10631 1613 10731
rect 1982 10627 2032 10727
rect 2195 10627 2245 10727
rect 2403 10627 2453 10727
rect 2611 10627 2661 10727
rect 6686 10467 6736 10567
rect 6894 10467 6944 10567
rect 7102 10467 7152 10567
rect 7315 10467 7365 10567
rect 11642 10625 11692 10725
rect 11855 10625 11905 10725
rect 12063 10625 12113 10725
rect 12271 10625 12321 10725
rect 9224 10464 9274 10564
rect 9432 10464 9482 10564
rect 9640 10464 9690 10564
rect 9853 10464 9903 10564
rect 12690 10621 12740 10721
rect 12903 10621 12953 10721
rect 13111 10621 13161 10721
rect 13319 10621 13369 10721
rect 17394 10461 17444 10561
rect 17602 10461 17652 10561
rect 17810 10461 17860 10561
rect 18023 10461 18073 10561
rect 22607 10629 22657 10729
rect 22820 10629 22870 10729
rect 23028 10629 23078 10729
rect 23236 10629 23286 10729
rect 19932 10458 19982 10558
rect 20140 10458 20190 10558
rect 20348 10458 20398 10558
rect 20561 10458 20611 10558
rect 23655 10625 23705 10725
rect 23868 10625 23918 10725
rect 24076 10625 24126 10725
rect 24284 10625 24334 10725
rect 28359 10465 28409 10565
rect 28567 10465 28617 10565
rect 28775 10465 28825 10565
rect 28988 10465 29038 10565
rect 33315 10623 33365 10723
rect 33528 10623 33578 10723
rect 33736 10623 33786 10723
rect 33944 10623 33994 10723
rect 30897 10462 30947 10562
rect 31105 10462 31155 10562
rect 31313 10462 31363 10562
rect 31526 10462 31576 10562
rect 34363 10619 34413 10719
rect 34576 10619 34626 10719
rect 34784 10619 34834 10719
rect 34992 10619 35042 10719
rect 39067 10459 39117 10559
rect 39275 10459 39325 10559
rect 39483 10459 39533 10559
rect 39696 10459 39746 10559
rect 41605 10456 41655 10556
rect 41813 10456 41863 10556
rect 42021 10456 42071 10556
rect 42234 10456 42284 10556
rect 934 9952 984 10052
rect 1147 9952 1197 10052
rect 1355 9952 1405 10052
rect 1563 9952 1613 10052
rect 3429 9947 3479 10047
rect 3642 9947 3692 10047
rect 3850 9947 3900 10047
rect 4058 9947 4108 10047
rect 8176 9789 8226 9889
rect 8384 9789 8434 9889
rect 8592 9789 8642 9889
rect 8805 9789 8855 9889
rect 11642 9946 11692 10046
rect 11855 9946 11905 10046
rect 12063 9946 12113 10046
rect 12271 9946 12321 10046
rect 9224 9785 9274 9885
rect 9432 9785 9482 9885
rect 9640 9785 9690 9885
rect 9853 9785 9903 9885
rect 14137 9941 14187 10041
rect 14350 9941 14400 10041
rect 14558 9941 14608 10041
rect 14766 9941 14816 10041
rect 18884 9783 18934 9883
rect 19092 9783 19142 9883
rect 19300 9783 19350 9883
rect 19513 9783 19563 9883
rect 22607 9950 22657 10050
rect 22820 9950 22870 10050
rect 23028 9950 23078 10050
rect 23236 9950 23286 10050
rect 19932 9779 19982 9879
rect 20140 9779 20190 9879
rect 20348 9779 20398 9879
rect 20561 9779 20611 9879
rect 25102 9945 25152 10045
rect 25315 9945 25365 10045
rect 25523 9945 25573 10045
rect 25731 9945 25781 10045
rect 29849 9787 29899 9887
rect 30057 9787 30107 9887
rect 30265 9787 30315 9887
rect 30478 9787 30528 9887
rect 33315 9944 33365 10044
rect 33528 9944 33578 10044
rect 33736 9944 33786 10044
rect 33944 9944 33994 10044
rect 30897 9783 30947 9883
rect 31105 9783 31155 9883
rect 31313 9783 31363 9883
rect 31526 9783 31576 9883
rect 35810 9939 35860 10039
rect 36023 9939 36073 10039
rect 36231 9939 36281 10039
rect 36439 9939 36489 10039
rect 40557 9781 40607 9881
rect 40765 9781 40815 9881
rect 40973 9781 41023 9881
rect 41186 9781 41236 9881
rect 41605 9777 41655 9877
rect 41813 9777 41863 9877
rect 42021 9777 42071 9877
rect 42234 9777 42284 9877
rect 934 9184 984 9284
rect 1147 9184 1197 9284
rect 1355 9184 1405 9284
rect 1563 9184 1613 9284
rect 1982 9180 2032 9280
rect 2195 9180 2245 9280
rect 2403 9180 2453 9280
rect 2611 9180 2661 9280
rect 6729 9022 6779 9122
rect 6937 9022 6987 9122
rect 7145 9022 7195 9122
rect 7358 9022 7408 9122
rect 11642 9178 11692 9278
rect 11855 9178 11905 9278
rect 12063 9178 12113 9278
rect 12271 9178 12321 9278
rect 9224 9017 9274 9117
rect 9432 9017 9482 9117
rect 9640 9017 9690 9117
rect 9853 9017 9903 9117
rect 12690 9174 12740 9274
rect 12903 9174 12953 9274
rect 13111 9174 13161 9274
rect 13319 9174 13369 9274
rect 17437 9016 17487 9116
rect 17645 9016 17695 9116
rect 17853 9016 17903 9116
rect 18066 9016 18116 9116
rect 22607 9182 22657 9282
rect 22820 9182 22870 9282
rect 23028 9182 23078 9282
rect 23236 9182 23286 9282
rect 19932 9011 19982 9111
rect 20140 9011 20190 9111
rect 20348 9011 20398 9111
rect 20561 9011 20611 9111
rect 23655 9178 23705 9278
rect 23868 9178 23918 9278
rect 24076 9178 24126 9278
rect 24284 9178 24334 9278
rect 28402 9020 28452 9120
rect 28610 9020 28660 9120
rect 28818 9020 28868 9120
rect 29031 9020 29081 9120
rect 33315 9176 33365 9276
rect 33528 9176 33578 9276
rect 33736 9176 33786 9276
rect 33944 9176 33994 9276
rect 30897 9015 30947 9115
rect 31105 9015 31155 9115
rect 31313 9015 31363 9115
rect 31526 9015 31576 9115
rect 34363 9172 34413 9272
rect 34576 9172 34626 9272
rect 34784 9172 34834 9272
rect 34992 9172 35042 9272
rect 39110 9014 39160 9114
rect 39318 9014 39368 9114
rect 39526 9014 39576 9114
rect 39739 9014 39789 9114
rect 41605 9009 41655 9109
rect 41813 9009 41863 9109
rect 42021 9009 42071 9109
rect 42234 9009 42284 9109
rect 934 8505 984 8605
rect 1147 8505 1197 8605
rect 1355 8505 1405 8605
rect 1563 8505 1613 8605
rect 4537 8496 4587 8596
rect 4750 8496 4800 8596
rect 4958 8496 5008 8596
rect 5166 8496 5216 8596
rect 8176 8342 8226 8442
rect 8384 8342 8434 8442
rect 8592 8342 8642 8442
rect 8805 8342 8855 8442
rect 11642 8499 11692 8599
rect 11855 8499 11905 8599
rect 12063 8499 12113 8599
rect 12271 8499 12321 8599
rect 9224 8338 9274 8438
rect 9432 8338 9482 8438
rect 9640 8338 9690 8438
rect 9853 8338 9903 8438
rect 15245 8490 15295 8590
rect 15458 8490 15508 8590
rect 15666 8490 15716 8590
rect 15874 8490 15924 8590
rect 18884 8336 18934 8436
rect 19092 8336 19142 8436
rect 19300 8336 19350 8436
rect 19513 8336 19563 8436
rect 22607 8503 22657 8603
rect 22820 8503 22870 8603
rect 23028 8503 23078 8603
rect 23236 8503 23286 8603
rect 19932 8332 19982 8432
rect 20140 8332 20190 8432
rect 20348 8332 20398 8432
rect 20561 8332 20611 8432
rect 26210 8494 26260 8594
rect 26423 8494 26473 8594
rect 26631 8494 26681 8594
rect 26839 8494 26889 8594
rect 29849 8340 29899 8440
rect 30057 8340 30107 8440
rect 30265 8340 30315 8440
rect 30478 8340 30528 8440
rect 33315 8497 33365 8597
rect 33528 8497 33578 8597
rect 33736 8497 33786 8597
rect 33944 8497 33994 8597
rect 30897 8336 30947 8436
rect 31105 8336 31155 8436
rect 31313 8336 31363 8436
rect 31526 8336 31576 8436
rect 36918 8488 36968 8588
rect 37131 8488 37181 8588
rect 37339 8488 37389 8588
rect 37547 8488 37597 8588
rect 40557 8334 40607 8434
rect 40765 8334 40815 8434
rect 40973 8334 41023 8434
rect 41186 8334 41236 8434
rect 41605 8330 41655 8430
rect 41813 8330 41863 8430
rect 42021 8330 42071 8430
rect 42234 8330 42284 8430
rect 931 7590 981 7690
rect 1144 7590 1194 7690
rect 1352 7590 1402 7690
rect 1560 7590 1610 7690
rect 1979 7586 2029 7686
rect 2192 7586 2242 7686
rect 2400 7586 2450 7686
rect 2608 7586 2658 7686
rect 5618 7432 5668 7532
rect 5826 7432 5876 7532
rect 6034 7432 6084 7532
rect 6247 7432 6297 7532
rect 11639 7584 11689 7684
rect 11852 7584 11902 7684
rect 12060 7584 12110 7684
rect 12268 7584 12318 7684
rect 9221 7423 9271 7523
rect 9429 7423 9479 7523
rect 9637 7423 9687 7523
rect 9850 7423 9900 7523
rect 12687 7580 12737 7680
rect 12900 7580 12950 7680
rect 13108 7580 13158 7680
rect 13316 7580 13366 7680
rect 16326 7426 16376 7526
rect 16534 7426 16584 7526
rect 16742 7426 16792 7526
rect 16955 7426 17005 7526
rect 22604 7588 22654 7688
rect 22817 7588 22867 7688
rect 23025 7588 23075 7688
rect 23233 7588 23283 7688
rect 19929 7417 19979 7517
rect 20137 7417 20187 7517
rect 20345 7417 20395 7517
rect 20558 7417 20608 7517
rect 23652 7584 23702 7684
rect 23865 7584 23915 7684
rect 24073 7584 24123 7684
rect 24281 7584 24331 7684
rect 27291 7430 27341 7530
rect 27499 7430 27549 7530
rect 27707 7430 27757 7530
rect 27920 7430 27970 7530
rect 33312 7582 33362 7682
rect 33525 7582 33575 7682
rect 33733 7582 33783 7682
rect 33941 7582 33991 7682
rect 30894 7421 30944 7521
rect 31102 7421 31152 7521
rect 31310 7421 31360 7521
rect 31523 7421 31573 7521
rect 34360 7578 34410 7678
rect 34573 7578 34623 7678
rect 34781 7578 34831 7678
rect 34989 7578 35039 7678
rect 37999 7424 38049 7524
rect 38207 7424 38257 7524
rect 38415 7424 38465 7524
rect 38628 7424 38678 7524
rect 41602 7415 41652 7515
rect 41810 7415 41860 7515
rect 42018 7415 42068 7515
rect 42231 7415 42281 7515
rect 931 6911 981 7011
rect 1144 6911 1194 7011
rect 1352 6911 1402 7011
rect 1560 6911 1610 7011
rect 3426 6906 3476 7006
rect 3639 6906 3689 7006
rect 3847 6906 3897 7006
rect 4055 6906 4105 7006
rect 8173 6748 8223 6848
rect 8381 6748 8431 6848
rect 8589 6748 8639 6848
rect 8802 6748 8852 6848
rect 11639 6905 11689 7005
rect 11852 6905 11902 7005
rect 12060 6905 12110 7005
rect 12268 6905 12318 7005
rect 9221 6744 9271 6844
rect 9429 6744 9479 6844
rect 9637 6744 9687 6844
rect 9850 6744 9900 6844
rect 14134 6900 14184 7000
rect 14347 6900 14397 7000
rect 14555 6900 14605 7000
rect 14763 6900 14813 7000
rect 18881 6742 18931 6842
rect 19089 6742 19139 6842
rect 19297 6742 19347 6842
rect 19510 6742 19560 6842
rect 22604 6909 22654 7009
rect 22817 6909 22867 7009
rect 23025 6909 23075 7009
rect 23233 6909 23283 7009
rect 19929 6738 19979 6838
rect 20137 6738 20187 6838
rect 20345 6738 20395 6838
rect 20558 6738 20608 6838
rect 25099 6904 25149 7004
rect 25312 6904 25362 7004
rect 25520 6904 25570 7004
rect 25728 6904 25778 7004
rect 29846 6746 29896 6846
rect 30054 6746 30104 6846
rect 30262 6746 30312 6846
rect 30475 6746 30525 6846
rect 33312 6903 33362 7003
rect 33525 6903 33575 7003
rect 33733 6903 33783 7003
rect 33941 6903 33991 7003
rect 30894 6742 30944 6842
rect 31102 6742 31152 6842
rect 31310 6742 31360 6842
rect 31523 6742 31573 6842
rect 35807 6898 35857 6998
rect 36020 6898 36070 6998
rect 36228 6898 36278 6998
rect 36436 6898 36486 6998
rect 40554 6740 40604 6840
rect 40762 6740 40812 6840
rect 40970 6740 41020 6840
rect 41183 6740 41233 6840
rect 41602 6736 41652 6836
rect 41810 6736 41860 6836
rect 42018 6736 42068 6836
rect 42231 6736 42281 6836
rect 931 6143 981 6243
rect 1144 6143 1194 6243
rect 1352 6143 1402 6243
rect 1560 6143 1610 6243
rect 1979 6139 2029 6239
rect 2192 6139 2242 6239
rect 2400 6139 2450 6239
rect 2608 6139 2658 6239
rect 6726 5981 6776 6081
rect 6934 5981 6984 6081
rect 7142 5981 7192 6081
rect 7355 5981 7405 6081
rect 11639 6137 11689 6237
rect 11852 6137 11902 6237
rect 12060 6137 12110 6237
rect 12268 6137 12318 6237
rect 9221 5976 9271 6076
rect 9429 5976 9479 6076
rect 9637 5976 9687 6076
rect 9850 5976 9900 6076
rect 12687 6133 12737 6233
rect 12900 6133 12950 6233
rect 13108 6133 13158 6233
rect 13316 6133 13366 6233
rect 17434 5975 17484 6075
rect 17642 5975 17692 6075
rect 17850 5975 17900 6075
rect 18063 5975 18113 6075
rect 22604 6141 22654 6241
rect 22817 6141 22867 6241
rect 23025 6141 23075 6241
rect 23233 6141 23283 6241
rect 19929 5970 19979 6070
rect 20137 5970 20187 6070
rect 20345 5970 20395 6070
rect 20558 5970 20608 6070
rect 23652 6137 23702 6237
rect 23865 6137 23915 6237
rect 24073 6137 24123 6237
rect 24281 6137 24331 6237
rect 28399 5979 28449 6079
rect 28607 5979 28657 6079
rect 28815 5979 28865 6079
rect 29028 5979 29078 6079
rect 33312 6135 33362 6235
rect 33525 6135 33575 6235
rect 33733 6135 33783 6235
rect 33941 6135 33991 6235
rect 30894 5974 30944 6074
rect 31102 5974 31152 6074
rect 31310 5974 31360 6074
rect 31523 5974 31573 6074
rect 34360 6131 34410 6231
rect 34573 6131 34623 6231
rect 34781 6131 34831 6231
rect 34989 6131 35039 6231
rect 39107 5973 39157 6073
rect 39315 5973 39365 6073
rect 39523 5973 39573 6073
rect 39736 5973 39786 6073
rect 41602 5968 41652 6068
rect 41810 5968 41860 6068
rect 42018 5968 42068 6068
rect 42231 5968 42281 6068
rect 931 5464 981 5564
rect 1144 5464 1194 5564
rect 1352 5464 1402 5564
rect 1560 5464 1610 5564
rect 3469 5461 3519 5561
rect 3682 5461 3732 5561
rect 3890 5461 3940 5561
rect 4098 5461 4148 5561
rect 8173 5301 8223 5401
rect 8381 5301 8431 5401
rect 8589 5301 8639 5401
rect 8802 5301 8852 5401
rect 11639 5458 11689 5558
rect 11852 5458 11902 5558
rect 12060 5458 12110 5558
rect 12268 5458 12318 5558
rect 9221 5297 9271 5397
rect 9429 5297 9479 5397
rect 9637 5297 9687 5397
rect 9850 5297 9900 5397
rect 14177 5455 14227 5555
rect 14390 5455 14440 5555
rect 14598 5455 14648 5555
rect 14806 5455 14856 5555
rect 18881 5295 18931 5395
rect 19089 5295 19139 5395
rect 19297 5295 19347 5395
rect 19510 5295 19560 5395
rect 22604 5462 22654 5562
rect 22817 5462 22867 5562
rect 23025 5462 23075 5562
rect 23233 5462 23283 5562
rect 19929 5291 19979 5391
rect 20137 5291 20187 5391
rect 20345 5291 20395 5391
rect 20558 5291 20608 5391
rect 25142 5459 25192 5559
rect 25355 5459 25405 5559
rect 25563 5459 25613 5559
rect 25771 5459 25821 5559
rect 29846 5299 29896 5399
rect 30054 5299 30104 5399
rect 30262 5299 30312 5399
rect 30475 5299 30525 5399
rect 33312 5456 33362 5556
rect 33525 5456 33575 5556
rect 33733 5456 33783 5556
rect 33941 5456 33991 5556
rect 30894 5295 30944 5395
rect 31102 5295 31152 5395
rect 31310 5295 31360 5395
rect 31523 5295 31573 5395
rect 35850 5453 35900 5553
rect 36063 5453 36113 5553
rect 36271 5453 36321 5553
rect 36479 5453 36529 5553
rect 40554 5293 40604 5393
rect 40762 5293 40812 5393
rect 40970 5293 41020 5393
rect 41183 5293 41233 5393
rect 41602 5289 41652 5389
rect 41810 5289 41860 5389
rect 42018 5289 42068 5389
rect 42231 5289 42281 5389
rect 932 4623 982 4723
rect 1145 4623 1195 4723
rect 1353 4623 1403 4723
rect 1561 4623 1611 4723
rect 1980 4619 2030 4719
rect 2193 4619 2243 4719
rect 2401 4619 2451 4719
rect 2609 4619 2659 4719
rect 4882 4625 4932 4725
rect 5095 4625 5145 4725
rect 5303 4625 5353 4725
rect 5511 4625 5561 4725
rect 6684 4459 6734 4559
rect 6892 4459 6942 4559
rect 7100 4459 7150 4559
rect 7313 4459 7363 4559
rect 11640 4617 11690 4717
rect 11853 4617 11903 4717
rect 12061 4617 12111 4717
rect 12269 4617 12319 4717
rect 9222 4456 9272 4556
rect 9430 4456 9480 4556
rect 9638 4456 9688 4556
rect 9851 4456 9901 4556
rect 12688 4613 12738 4713
rect 12901 4613 12951 4713
rect 13109 4613 13159 4713
rect 13317 4613 13367 4713
rect 15590 4619 15640 4719
rect 15803 4619 15853 4719
rect 16011 4619 16061 4719
rect 16219 4619 16269 4719
rect 17392 4453 17442 4553
rect 17600 4453 17650 4553
rect 17808 4453 17858 4553
rect 18021 4453 18071 4553
rect 22605 4621 22655 4721
rect 22818 4621 22868 4721
rect 23026 4621 23076 4721
rect 23234 4621 23284 4721
rect 19930 4450 19980 4550
rect 20138 4450 20188 4550
rect 20346 4450 20396 4550
rect 20559 4450 20609 4550
rect 23653 4617 23703 4717
rect 23866 4617 23916 4717
rect 24074 4617 24124 4717
rect 24282 4617 24332 4717
rect 26555 4623 26605 4723
rect 26768 4623 26818 4723
rect 26976 4623 27026 4723
rect 27184 4623 27234 4723
rect 28357 4457 28407 4557
rect 28565 4457 28615 4557
rect 28773 4457 28823 4557
rect 28986 4457 29036 4557
rect 33313 4615 33363 4715
rect 33526 4615 33576 4715
rect 33734 4615 33784 4715
rect 33942 4615 33992 4715
rect 30895 4454 30945 4554
rect 31103 4454 31153 4554
rect 31311 4454 31361 4554
rect 31524 4454 31574 4554
rect 34361 4611 34411 4711
rect 34574 4611 34624 4711
rect 34782 4611 34832 4711
rect 34990 4611 35040 4711
rect 37263 4617 37313 4717
rect 37476 4617 37526 4717
rect 37684 4617 37734 4717
rect 37892 4617 37942 4717
rect 39065 4451 39115 4551
rect 39273 4451 39323 4551
rect 39481 4451 39531 4551
rect 39694 4451 39744 4551
rect 41603 4448 41653 4548
rect 41811 4448 41861 4548
rect 42019 4448 42069 4548
rect 42232 4448 42282 4548
rect 932 3944 982 4044
rect 1145 3944 1195 4044
rect 1353 3944 1403 4044
rect 1561 3944 1611 4044
rect 3427 3939 3477 4039
rect 3640 3939 3690 4039
rect 3848 3939 3898 4039
rect 4056 3939 4106 4039
rect 8174 3781 8224 3881
rect 8382 3781 8432 3881
rect 8590 3781 8640 3881
rect 8803 3781 8853 3881
rect 11640 3938 11690 4038
rect 11853 3938 11903 4038
rect 12061 3938 12111 4038
rect 12269 3938 12319 4038
rect 9222 3777 9272 3877
rect 9430 3777 9480 3877
rect 9638 3777 9688 3877
rect 9851 3777 9901 3877
rect 14135 3933 14185 4033
rect 14348 3933 14398 4033
rect 14556 3933 14606 4033
rect 14764 3933 14814 4033
rect 18882 3775 18932 3875
rect 19090 3775 19140 3875
rect 19298 3775 19348 3875
rect 19511 3775 19561 3875
rect 22605 3942 22655 4042
rect 22818 3942 22868 4042
rect 23026 3942 23076 4042
rect 23234 3942 23284 4042
rect 19930 3771 19980 3871
rect 20138 3771 20188 3871
rect 20346 3771 20396 3871
rect 20559 3771 20609 3871
rect 25100 3937 25150 4037
rect 25313 3937 25363 4037
rect 25521 3937 25571 4037
rect 25729 3937 25779 4037
rect 29847 3779 29897 3879
rect 30055 3779 30105 3879
rect 30263 3779 30313 3879
rect 30476 3779 30526 3879
rect 33313 3936 33363 4036
rect 33526 3936 33576 4036
rect 33734 3936 33784 4036
rect 33942 3936 33992 4036
rect 30895 3775 30945 3875
rect 31103 3775 31153 3875
rect 31311 3775 31361 3875
rect 31524 3775 31574 3875
rect 35808 3931 35858 4031
rect 36021 3931 36071 4031
rect 36229 3931 36279 4031
rect 36437 3931 36487 4031
rect 40555 3773 40605 3873
rect 40763 3773 40813 3873
rect 40971 3773 41021 3873
rect 41184 3773 41234 3873
rect 41603 3769 41653 3869
rect 41811 3769 41861 3869
rect 42019 3769 42069 3869
rect 42232 3769 42282 3869
rect 932 3176 982 3276
rect 1145 3176 1195 3276
rect 1353 3176 1403 3276
rect 1561 3176 1611 3276
rect 1980 3172 2030 3272
rect 2193 3172 2243 3272
rect 2401 3172 2451 3272
rect 2609 3172 2659 3272
rect 6727 3014 6777 3114
rect 6935 3014 6985 3114
rect 7143 3014 7193 3114
rect 7356 3014 7406 3114
rect 11640 3170 11690 3270
rect 11853 3170 11903 3270
rect 12061 3170 12111 3270
rect 12269 3170 12319 3270
rect 9222 3009 9272 3109
rect 9430 3009 9480 3109
rect 9638 3009 9688 3109
rect 9851 3009 9901 3109
rect 12688 3166 12738 3266
rect 12901 3166 12951 3266
rect 13109 3166 13159 3266
rect 13317 3166 13367 3266
rect 17435 3008 17485 3108
rect 17643 3008 17693 3108
rect 17851 3008 17901 3108
rect 18064 3008 18114 3108
rect 22605 3174 22655 3274
rect 22818 3174 22868 3274
rect 23026 3174 23076 3274
rect 23234 3174 23284 3274
rect 19930 3003 19980 3103
rect 20138 3003 20188 3103
rect 20346 3003 20396 3103
rect 20559 3003 20609 3103
rect 23653 3170 23703 3270
rect 23866 3170 23916 3270
rect 24074 3170 24124 3270
rect 24282 3170 24332 3270
rect 28400 3012 28450 3112
rect 28608 3012 28658 3112
rect 28816 3012 28866 3112
rect 29029 3012 29079 3112
rect 33313 3168 33363 3268
rect 33526 3168 33576 3268
rect 33734 3168 33784 3268
rect 33942 3168 33992 3268
rect 30895 3007 30945 3107
rect 31103 3007 31153 3107
rect 31311 3007 31361 3107
rect 31524 3007 31574 3107
rect 34361 3164 34411 3264
rect 34574 3164 34624 3264
rect 34782 3164 34832 3264
rect 34990 3164 35040 3264
rect 39108 3006 39158 3106
rect 39316 3006 39366 3106
rect 39524 3006 39574 3106
rect 39737 3006 39787 3106
rect 41603 3001 41653 3101
rect 41811 3001 41861 3101
rect 42019 3001 42069 3101
rect 42232 3001 42282 3101
rect 932 2497 982 2597
rect 1145 2497 1195 2597
rect 1353 2497 1403 2597
rect 1561 2497 1611 2597
rect 8174 2334 8224 2434
rect 8382 2334 8432 2434
rect 8590 2334 8640 2434
rect 8803 2334 8853 2434
rect 11640 2491 11690 2591
rect 11853 2491 11903 2591
rect 12061 2491 12111 2591
rect 12269 2491 12319 2591
rect 9222 2330 9272 2430
rect 9430 2330 9480 2430
rect 9638 2330 9688 2430
rect 9851 2330 9901 2430
rect 18882 2328 18932 2428
rect 19090 2328 19140 2428
rect 19298 2328 19348 2428
rect 19511 2328 19561 2428
rect 22605 2495 22655 2595
rect 22818 2495 22868 2595
rect 23026 2495 23076 2595
rect 23234 2495 23284 2595
rect 19930 2324 19980 2424
rect 20138 2324 20188 2424
rect 20346 2324 20396 2424
rect 20559 2324 20609 2424
rect 29847 2332 29897 2432
rect 30055 2332 30105 2432
rect 30263 2332 30313 2432
rect 30476 2332 30526 2432
rect 33313 2489 33363 2589
rect 33526 2489 33576 2589
rect 33734 2489 33784 2589
rect 33942 2489 33992 2589
rect 30895 2328 30945 2428
rect 31103 2328 31153 2428
rect 31311 2328 31361 2428
rect 31524 2328 31574 2428
rect 40555 2326 40605 2426
rect 40763 2326 40813 2426
rect 40971 2326 41021 2426
rect 41184 2326 41234 2426
rect 41603 2322 41653 2422
rect 41811 2322 41861 2422
rect 42019 2322 42069 2422
rect 42232 2322 42282 2422
rect 10643 338 10693 438
rect 10856 338 10906 438
rect 11064 338 11114 438
rect 11272 338 11322 438
rect 21280 325 21330 425
rect 21493 325 21543 425
rect 21701 325 21751 425
rect 21909 325 21959 425
rect 32316 336 32366 436
rect 32529 336 32579 436
rect 32737 336 32787 436
rect 32945 336 32995 436
<< ndiff >>
rect 9174 13638 9223 13650
rect 9174 13618 9185 13638
rect 9205 13618 9223 13638
rect 9174 13608 9223 13618
rect 9273 13634 9317 13650
rect 9273 13614 9288 13634
rect 9308 13614 9317 13634
rect 9273 13608 9317 13614
rect 9387 13634 9431 13650
rect 9387 13614 9396 13634
rect 9416 13614 9431 13634
rect 9387 13608 9431 13614
rect 9481 13638 9530 13650
rect 9481 13618 9499 13638
rect 9519 13618 9530 13638
rect 9481 13608 9530 13618
rect 9595 13634 9639 13650
rect 9595 13614 9604 13634
rect 9624 13614 9639 13634
rect 9595 13608 9639 13614
rect 9689 13638 9738 13650
rect 9689 13618 9707 13638
rect 9727 13618 9738 13638
rect 9689 13608 9738 13618
rect 9808 13634 9852 13650
rect 9808 13614 9817 13634
rect 9837 13614 9852 13634
rect 9808 13608 9852 13614
rect 9902 13638 9951 13650
rect 9902 13618 9920 13638
rect 9940 13618 9951 13638
rect 9902 13608 9951 13618
rect 884 13511 933 13521
rect 884 13491 895 13511
rect 915 13491 933 13511
rect 884 13479 933 13491
rect 983 13515 1027 13521
rect 983 13495 998 13515
rect 1018 13495 1027 13515
rect 983 13479 1027 13495
rect 1097 13511 1146 13521
rect 1097 13491 1108 13511
rect 1128 13491 1146 13511
rect 1097 13479 1146 13491
rect 1196 13515 1240 13521
rect 1196 13495 1211 13515
rect 1231 13495 1240 13515
rect 1196 13479 1240 13495
rect 1305 13511 1354 13521
rect 1305 13491 1316 13511
rect 1336 13491 1354 13511
rect 1305 13479 1354 13491
rect 1404 13515 1448 13521
rect 1404 13495 1419 13515
rect 1439 13495 1448 13515
rect 1404 13479 1448 13495
rect 1518 13515 1562 13521
rect 1518 13495 1527 13515
rect 1547 13495 1562 13515
rect 1518 13479 1562 13495
rect 1612 13511 1661 13521
rect 1612 13491 1630 13511
rect 1650 13491 1661 13511
rect 1612 13479 1661 13491
rect 1932 13507 1981 13517
rect 1932 13487 1943 13507
rect 1963 13487 1981 13507
rect 1932 13475 1981 13487
rect 2031 13511 2075 13517
rect 2031 13491 2046 13511
rect 2066 13491 2075 13511
rect 2031 13475 2075 13491
rect 2145 13507 2194 13517
rect 2145 13487 2156 13507
rect 2176 13487 2194 13507
rect 2145 13475 2194 13487
rect 2244 13511 2288 13517
rect 2244 13491 2259 13511
rect 2279 13491 2288 13511
rect 2244 13475 2288 13491
rect 2353 13507 2402 13517
rect 2353 13487 2364 13507
rect 2384 13487 2402 13507
rect 2353 13475 2402 13487
rect 2452 13511 2496 13517
rect 2452 13491 2467 13511
rect 2487 13491 2496 13511
rect 2452 13475 2496 13491
rect 2566 13511 2610 13517
rect 2566 13491 2575 13511
rect 2595 13491 2610 13511
rect 2566 13475 2610 13491
rect 2660 13507 2709 13517
rect 2660 13487 2678 13507
rect 2698 13487 2709 13507
rect 2660 13475 2709 13487
rect 19882 13632 19931 13644
rect 19882 13612 19893 13632
rect 19913 13612 19931 13632
rect 19882 13602 19931 13612
rect 19981 13628 20025 13644
rect 19981 13608 19996 13628
rect 20016 13608 20025 13628
rect 19981 13602 20025 13608
rect 20095 13628 20139 13644
rect 20095 13608 20104 13628
rect 20124 13608 20139 13628
rect 20095 13602 20139 13608
rect 20189 13632 20238 13644
rect 20189 13612 20207 13632
rect 20227 13612 20238 13632
rect 20189 13602 20238 13612
rect 20303 13628 20347 13644
rect 20303 13608 20312 13628
rect 20332 13608 20347 13628
rect 20303 13602 20347 13608
rect 20397 13632 20446 13644
rect 20397 13612 20415 13632
rect 20435 13612 20446 13632
rect 20397 13602 20446 13612
rect 20516 13628 20560 13644
rect 20516 13608 20525 13628
rect 20545 13608 20560 13628
rect 20516 13602 20560 13608
rect 20610 13632 20659 13644
rect 20610 13612 20628 13632
rect 20648 13612 20659 13632
rect 20610 13602 20659 13612
rect 11592 13505 11641 13515
rect 11592 13485 11603 13505
rect 11623 13485 11641 13505
rect 11592 13473 11641 13485
rect 11691 13509 11735 13515
rect 11691 13489 11706 13509
rect 11726 13489 11735 13509
rect 11691 13473 11735 13489
rect 11805 13505 11854 13515
rect 11805 13485 11816 13505
rect 11836 13485 11854 13505
rect 11805 13473 11854 13485
rect 11904 13509 11948 13515
rect 11904 13489 11919 13509
rect 11939 13489 11948 13509
rect 11904 13473 11948 13489
rect 12013 13505 12062 13515
rect 12013 13485 12024 13505
rect 12044 13485 12062 13505
rect 12013 13473 12062 13485
rect 12112 13509 12156 13515
rect 12112 13489 12127 13509
rect 12147 13489 12156 13509
rect 12112 13473 12156 13489
rect 12226 13509 12270 13515
rect 12226 13489 12235 13509
rect 12255 13489 12270 13509
rect 12226 13473 12270 13489
rect 12320 13505 12369 13515
rect 12320 13485 12338 13505
rect 12358 13485 12369 13505
rect 12320 13473 12369 13485
rect 12640 13501 12689 13511
rect 12640 13481 12651 13501
rect 12671 13481 12689 13501
rect 12640 13469 12689 13481
rect 12739 13505 12783 13511
rect 12739 13485 12754 13505
rect 12774 13485 12783 13505
rect 12739 13469 12783 13485
rect 12853 13501 12902 13511
rect 12853 13481 12864 13501
rect 12884 13481 12902 13501
rect 12853 13469 12902 13481
rect 12952 13505 12996 13511
rect 12952 13485 12967 13505
rect 12987 13485 12996 13505
rect 12952 13469 12996 13485
rect 13061 13501 13110 13511
rect 13061 13481 13072 13501
rect 13092 13481 13110 13501
rect 13061 13469 13110 13481
rect 13160 13505 13204 13511
rect 13160 13485 13175 13505
rect 13195 13485 13204 13505
rect 13160 13469 13204 13485
rect 13274 13505 13318 13511
rect 13274 13485 13283 13505
rect 13303 13485 13318 13505
rect 13274 13469 13318 13485
rect 13368 13501 13417 13511
rect 13368 13481 13386 13501
rect 13406 13481 13417 13501
rect 13368 13469 13417 13481
rect 30847 13636 30896 13648
rect 30847 13616 30858 13636
rect 30878 13616 30896 13636
rect 30847 13606 30896 13616
rect 30946 13632 30990 13648
rect 30946 13612 30961 13632
rect 30981 13612 30990 13632
rect 30946 13606 30990 13612
rect 31060 13632 31104 13648
rect 31060 13612 31069 13632
rect 31089 13612 31104 13632
rect 31060 13606 31104 13612
rect 31154 13636 31203 13648
rect 31154 13616 31172 13636
rect 31192 13616 31203 13636
rect 31154 13606 31203 13616
rect 31268 13632 31312 13648
rect 31268 13612 31277 13632
rect 31297 13612 31312 13632
rect 31268 13606 31312 13612
rect 31362 13636 31411 13648
rect 31362 13616 31380 13636
rect 31400 13616 31411 13636
rect 31362 13606 31411 13616
rect 31481 13632 31525 13648
rect 31481 13612 31490 13632
rect 31510 13612 31525 13632
rect 31481 13606 31525 13612
rect 31575 13636 31624 13648
rect 31575 13616 31593 13636
rect 31613 13616 31624 13636
rect 31575 13606 31624 13616
rect 22557 13509 22606 13519
rect 22557 13489 22568 13509
rect 22588 13489 22606 13509
rect 22557 13477 22606 13489
rect 22656 13513 22700 13519
rect 22656 13493 22671 13513
rect 22691 13493 22700 13513
rect 22656 13477 22700 13493
rect 22770 13509 22819 13519
rect 22770 13489 22781 13509
rect 22801 13489 22819 13509
rect 22770 13477 22819 13489
rect 22869 13513 22913 13519
rect 22869 13493 22884 13513
rect 22904 13493 22913 13513
rect 22869 13477 22913 13493
rect 22978 13509 23027 13519
rect 22978 13489 22989 13509
rect 23009 13489 23027 13509
rect 22978 13477 23027 13489
rect 23077 13513 23121 13519
rect 23077 13493 23092 13513
rect 23112 13493 23121 13513
rect 23077 13477 23121 13493
rect 23191 13513 23235 13519
rect 23191 13493 23200 13513
rect 23220 13493 23235 13513
rect 23191 13477 23235 13493
rect 23285 13509 23334 13519
rect 23285 13489 23303 13509
rect 23323 13489 23334 13509
rect 23285 13477 23334 13489
rect 23605 13505 23654 13515
rect 23605 13485 23616 13505
rect 23636 13485 23654 13505
rect 23605 13473 23654 13485
rect 23704 13509 23748 13515
rect 23704 13489 23719 13509
rect 23739 13489 23748 13509
rect 23704 13473 23748 13489
rect 23818 13505 23867 13515
rect 23818 13485 23829 13505
rect 23849 13485 23867 13505
rect 23818 13473 23867 13485
rect 23917 13509 23961 13515
rect 23917 13489 23932 13509
rect 23952 13489 23961 13509
rect 23917 13473 23961 13489
rect 24026 13505 24075 13515
rect 24026 13485 24037 13505
rect 24057 13485 24075 13505
rect 24026 13473 24075 13485
rect 24125 13509 24169 13515
rect 24125 13489 24140 13509
rect 24160 13489 24169 13509
rect 24125 13473 24169 13489
rect 24239 13509 24283 13515
rect 24239 13489 24248 13509
rect 24268 13489 24283 13509
rect 24239 13473 24283 13489
rect 24333 13505 24382 13515
rect 24333 13485 24351 13505
rect 24371 13485 24382 13505
rect 24333 13473 24382 13485
rect 41555 13630 41604 13642
rect 41555 13610 41566 13630
rect 41586 13610 41604 13630
rect 41555 13600 41604 13610
rect 41654 13626 41698 13642
rect 41654 13606 41669 13626
rect 41689 13606 41698 13626
rect 41654 13600 41698 13606
rect 41768 13626 41812 13642
rect 41768 13606 41777 13626
rect 41797 13606 41812 13626
rect 41768 13600 41812 13606
rect 41862 13630 41911 13642
rect 41862 13610 41880 13630
rect 41900 13610 41911 13630
rect 41862 13600 41911 13610
rect 41976 13626 42020 13642
rect 41976 13606 41985 13626
rect 42005 13606 42020 13626
rect 41976 13600 42020 13606
rect 42070 13630 42119 13642
rect 42070 13610 42088 13630
rect 42108 13610 42119 13630
rect 42070 13600 42119 13610
rect 42189 13626 42233 13642
rect 42189 13606 42198 13626
rect 42218 13606 42233 13626
rect 42189 13600 42233 13606
rect 42283 13630 42332 13642
rect 42283 13610 42301 13630
rect 42321 13610 42332 13630
rect 42283 13600 42332 13610
rect 33265 13503 33314 13513
rect 33265 13483 33276 13503
rect 33296 13483 33314 13503
rect 33265 13471 33314 13483
rect 33364 13507 33408 13513
rect 33364 13487 33379 13507
rect 33399 13487 33408 13507
rect 33364 13471 33408 13487
rect 33478 13503 33527 13513
rect 33478 13483 33489 13503
rect 33509 13483 33527 13503
rect 33478 13471 33527 13483
rect 33577 13507 33621 13513
rect 33577 13487 33592 13507
rect 33612 13487 33621 13507
rect 33577 13471 33621 13487
rect 33686 13503 33735 13513
rect 33686 13483 33697 13503
rect 33717 13483 33735 13503
rect 33686 13471 33735 13483
rect 33785 13507 33829 13513
rect 33785 13487 33800 13507
rect 33820 13487 33829 13507
rect 33785 13471 33829 13487
rect 33899 13507 33943 13513
rect 33899 13487 33908 13507
rect 33928 13487 33943 13507
rect 33899 13471 33943 13487
rect 33993 13503 34042 13513
rect 33993 13483 34011 13503
rect 34031 13483 34042 13503
rect 33993 13471 34042 13483
rect 34313 13499 34362 13509
rect 34313 13479 34324 13499
rect 34344 13479 34362 13499
rect 34313 13467 34362 13479
rect 34412 13503 34456 13509
rect 34412 13483 34427 13503
rect 34447 13483 34456 13503
rect 34412 13467 34456 13483
rect 34526 13499 34575 13509
rect 34526 13479 34537 13499
rect 34557 13479 34575 13499
rect 34526 13467 34575 13479
rect 34625 13503 34669 13509
rect 34625 13483 34640 13503
rect 34660 13483 34669 13503
rect 34625 13467 34669 13483
rect 34734 13499 34783 13509
rect 34734 13479 34745 13499
rect 34765 13479 34783 13499
rect 34734 13467 34783 13479
rect 34833 13503 34877 13509
rect 34833 13483 34848 13503
rect 34868 13483 34877 13503
rect 34833 13467 34877 13483
rect 34947 13503 34991 13509
rect 34947 13483 34956 13503
rect 34976 13483 34991 13503
rect 34947 13467 34991 13483
rect 35041 13499 35090 13509
rect 35041 13479 35059 13499
rect 35079 13479 35090 13499
rect 35041 13467 35090 13479
rect 8126 12963 8175 12975
rect 8126 12943 8137 12963
rect 8157 12943 8175 12963
rect 8126 12933 8175 12943
rect 8225 12959 8269 12975
rect 8225 12939 8240 12959
rect 8260 12939 8269 12959
rect 8225 12933 8269 12939
rect 8339 12959 8383 12975
rect 8339 12939 8348 12959
rect 8368 12939 8383 12959
rect 8339 12933 8383 12939
rect 8433 12963 8482 12975
rect 8433 12943 8451 12963
rect 8471 12943 8482 12963
rect 8433 12933 8482 12943
rect 8547 12959 8591 12975
rect 8547 12939 8556 12959
rect 8576 12939 8591 12959
rect 8547 12933 8591 12939
rect 8641 12963 8690 12975
rect 8641 12943 8659 12963
rect 8679 12943 8690 12963
rect 8641 12933 8690 12943
rect 8760 12959 8804 12975
rect 8760 12939 8769 12959
rect 8789 12939 8804 12959
rect 8760 12933 8804 12939
rect 8854 12963 8903 12975
rect 8854 12943 8872 12963
rect 8892 12943 8903 12963
rect 8854 12933 8903 12943
rect 9174 12959 9223 12971
rect 9174 12939 9185 12959
rect 9205 12939 9223 12959
rect 884 12832 933 12842
rect 884 12812 895 12832
rect 915 12812 933 12832
rect 884 12800 933 12812
rect 983 12836 1027 12842
rect 983 12816 998 12836
rect 1018 12816 1027 12836
rect 983 12800 1027 12816
rect 1097 12832 1146 12842
rect 1097 12812 1108 12832
rect 1128 12812 1146 12832
rect 1097 12800 1146 12812
rect 1196 12836 1240 12842
rect 1196 12816 1211 12836
rect 1231 12816 1240 12836
rect 1196 12800 1240 12816
rect 1305 12832 1354 12842
rect 1305 12812 1316 12832
rect 1336 12812 1354 12832
rect 1305 12800 1354 12812
rect 1404 12836 1448 12842
rect 1404 12816 1419 12836
rect 1439 12816 1448 12836
rect 1404 12800 1448 12816
rect 1518 12836 1562 12842
rect 1518 12816 1527 12836
rect 1547 12816 1562 12836
rect 1518 12800 1562 12816
rect 1612 12832 1661 12842
rect 9174 12929 9223 12939
rect 9273 12955 9317 12971
rect 9273 12935 9288 12955
rect 9308 12935 9317 12955
rect 9273 12929 9317 12935
rect 9387 12955 9431 12971
rect 9387 12935 9396 12955
rect 9416 12935 9431 12955
rect 9387 12929 9431 12935
rect 9481 12959 9530 12971
rect 9481 12939 9499 12959
rect 9519 12939 9530 12959
rect 9481 12929 9530 12939
rect 9595 12955 9639 12971
rect 9595 12935 9604 12955
rect 9624 12935 9639 12955
rect 9595 12929 9639 12935
rect 9689 12959 9738 12971
rect 9689 12939 9707 12959
rect 9727 12939 9738 12959
rect 9689 12929 9738 12939
rect 9808 12955 9852 12971
rect 9808 12935 9817 12955
rect 9837 12935 9852 12955
rect 9808 12929 9852 12935
rect 9902 12959 9951 12971
rect 9902 12939 9920 12959
rect 9940 12939 9951 12959
rect 9902 12929 9951 12939
rect 1612 12812 1630 12832
rect 1650 12812 1661 12832
rect 1612 12800 1661 12812
rect 3379 12827 3428 12837
rect 3379 12807 3390 12827
rect 3410 12807 3428 12827
rect 3379 12795 3428 12807
rect 3478 12831 3522 12837
rect 3478 12811 3493 12831
rect 3513 12811 3522 12831
rect 3478 12795 3522 12811
rect 3592 12827 3641 12837
rect 3592 12807 3603 12827
rect 3623 12807 3641 12827
rect 3592 12795 3641 12807
rect 3691 12831 3735 12837
rect 3691 12811 3706 12831
rect 3726 12811 3735 12831
rect 3691 12795 3735 12811
rect 3800 12827 3849 12837
rect 3800 12807 3811 12827
rect 3831 12807 3849 12827
rect 3800 12795 3849 12807
rect 3899 12831 3943 12837
rect 3899 12811 3914 12831
rect 3934 12811 3943 12831
rect 3899 12795 3943 12811
rect 4013 12831 4057 12837
rect 4013 12811 4022 12831
rect 4042 12811 4057 12831
rect 4013 12795 4057 12811
rect 4107 12827 4156 12837
rect 4107 12807 4125 12827
rect 4145 12807 4156 12827
rect 4107 12795 4156 12807
rect 18834 12957 18883 12969
rect 18834 12937 18845 12957
rect 18865 12937 18883 12957
rect 18834 12927 18883 12937
rect 18933 12953 18977 12969
rect 18933 12933 18948 12953
rect 18968 12933 18977 12953
rect 18933 12927 18977 12933
rect 19047 12953 19091 12969
rect 19047 12933 19056 12953
rect 19076 12933 19091 12953
rect 19047 12927 19091 12933
rect 19141 12957 19190 12969
rect 19141 12937 19159 12957
rect 19179 12937 19190 12957
rect 19141 12927 19190 12937
rect 19255 12953 19299 12969
rect 19255 12933 19264 12953
rect 19284 12933 19299 12953
rect 19255 12927 19299 12933
rect 19349 12957 19398 12969
rect 19349 12937 19367 12957
rect 19387 12937 19398 12957
rect 19349 12927 19398 12937
rect 19468 12953 19512 12969
rect 19468 12933 19477 12953
rect 19497 12933 19512 12953
rect 19468 12927 19512 12933
rect 19562 12957 19611 12969
rect 19562 12937 19580 12957
rect 19600 12937 19611 12957
rect 19562 12927 19611 12937
rect 19882 12953 19931 12965
rect 19882 12933 19893 12953
rect 19913 12933 19931 12953
rect 11592 12826 11641 12836
rect 11592 12806 11603 12826
rect 11623 12806 11641 12826
rect 11592 12794 11641 12806
rect 11691 12830 11735 12836
rect 11691 12810 11706 12830
rect 11726 12810 11735 12830
rect 11691 12794 11735 12810
rect 11805 12826 11854 12836
rect 11805 12806 11816 12826
rect 11836 12806 11854 12826
rect 11805 12794 11854 12806
rect 11904 12830 11948 12836
rect 11904 12810 11919 12830
rect 11939 12810 11948 12830
rect 11904 12794 11948 12810
rect 12013 12826 12062 12836
rect 12013 12806 12024 12826
rect 12044 12806 12062 12826
rect 12013 12794 12062 12806
rect 12112 12830 12156 12836
rect 12112 12810 12127 12830
rect 12147 12810 12156 12830
rect 12112 12794 12156 12810
rect 12226 12830 12270 12836
rect 12226 12810 12235 12830
rect 12255 12810 12270 12830
rect 12226 12794 12270 12810
rect 12320 12826 12369 12836
rect 19882 12923 19931 12933
rect 19981 12949 20025 12965
rect 19981 12929 19996 12949
rect 20016 12929 20025 12949
rect 19981 12923 20025 12929
rect 20095 12949 20139 12965
rect 20095 12929 20104 12949
rect 20124 12929 20139 12949
rect 20095 12923 20139 12929
rect 20189 12953 20238 12965
rect 20189 12933 20207 12953
rect 20227 12933 20238 12953
rect 20189 12923 20238 12933
rect 20303 12949 20347 12965
rect 20303 12929 20312 12949
rect 20332 12929 20347 12949
rect 20303 12923 20347 12929
rect 20397 12953 20446 12965
rect 20397 12933 20415 12953
rect 20435 12933 20446 12953
rect 20397 12923 20446 12933
rect 20516 12949 20560 12965
rect 20516 12929 20525 12949
rect 20545 12929 20560 12949
rect 20516 12923 20560 12929
rect 20610 12953 20659 12965
rect 20610 12933 20628 12953
rect 20648 12933 20659 12953
rect 20610 12923 20659 12933
rect 12320 12806 12338 12826
rect 12358 12806 12369 12826
rect 12320 12794 12369 12806
rect 14087 12821 14136 12831
rect 14087 12801 14098 12821
rect 14118 12801 14136 12821
rect 14087 12789 14136 12801
rect 14186 12825 14230 12831
rect 14186 12805 14201 12825
rect 14221 12805 14230 12825
rect 14186 12789 14230 12805
rect 14300 12821 14349 12831
rect 14300 12801 14311 12821
rect 14331 12801 14349 12821
rect 14300 12789 14349 12801
rect 14399 12825 14443 12831
rect 14399 12805 14414 12825
rect 14434 12805 14443 12825
rect 14399 12789 14443 12805
rect 14508 12821 14557 12831
rect 14508 12801 14519 12821
rect 14539 12801 14557 12821
rect 14508 12789 14557 12801
rect 14607 12825 14651 12831
rect 14607 12805 14622 12825
rect 14642 12805 14651 12825
rect 14607 12789 14651 12805
rect 14721 12825 14765 12831
rect 14721 12805 14730 12825
rect 14750 12805 14765 12825
rect 14721 12789 14765 12805
rect 14815 12821 14864 12831
rect 14815 12801 14833 12821
rect 14853 12801 14864 12821
rect 14815 12789 14864 12801
rect 29799 12961 29848 12973
rect 29799 12941 29810 12961
rect 29830 12941 29848 12961
rect 29799 12931 29848 12941
rect 29898 12957 29942 12973
rect 29898 12937 29913 12957
rect 29933 12937 29942 12957
rect 29898 12931 29942 12937
rect 30012 12957 30056 12973
rect 30012 12937 30021 12957
rect 30041 12937 30056 12957
rect 30012 12931 30056 12937
rect 30106 12961 30155 12973
rect 30106 12941 30124 12961
rect 30144 12941 30155 12961
rect 30106 12931 30155 12941
rect 30220 12957 30264 12973
rect 30220 12937 30229 12957
rect 30249 12937 30264 12957
rect 30220 12931 30264 12937
rect 30314 12961 30363 12973
rect 30314 12941 30332 12961
rect 30352 12941 30363 12961
rect 30314 12931 30363 12941
rect 30433 12957 30477 12973
rect 30433 12937 30442 12957
rect 30462 12937 30477 12957
rect 30433 12931 30477 12937
rect 30527 12961 30576 12973
rect 30527 12941 30545 12961
rect 30565 12941 30576 12961
rect 30527 12931 30576 12941
rect 30847 12957 30896 12969
rect 30847 12937 30858 12957
rect 30878 12937 30896 12957
rect 22557 12830 22606 12840
rect 22557 12810 22568 12830
rect 22588 12810 22606 12830
rect 22557 12798 22606 12810
rect 22656 12834 22700 12840
rect 22656 12814 22671 12834
rect 22691 12814 22700 12834
rect 22656 12798 22700 12814
rect 22770 12830 22819 12840
rect 22770 12810 22781 12830
rect 22801 12810 22819 12830
rect 22770 12798 22819 12810
rect 22869 12834 22913 12840
rect 22869 12814 22884 12834
rect 22904 12814 22913 12834
rect 22869 12798 22913 12814
rect 22978 12830 23027 12840
rect 22978 12810 22989 12830
rect 23009 12810 23027 12830
rect 22978 12798 23027 12810
rect 23077 12834 23121 12840
rect 23077 12814 23092 12834
rect 23112 12814 23121 12834
rect 23077 12798 23121 12814
rect 23191 12834 23235 12840
rect 23191 12814 23200 12834
rect 23220 12814 23235 12834
rect 23191 12798 23235 12814
rect 23285 12830 23334 12840
rect 30847 12927 30896 12937
rect 30946 12953 30990 12969
rect 30946 12933 30961 12953
rect 30981 12933 30990 12953
rect 30946 12927 30990 12933
rect 31060 12953 31104 12969
rect 31060 12933 31069 12953
rect 31089 12933 31104 12953
rect 31060 12927 31104 12933
rect 31154 12957 31203 12969
rect 31154 12937 31172 12957
rect 31192 12937 31203 12957
rect 31154 12927 31203 12937
rect 31268 12953 31312 12969
rect 31268 12933 31277 12953
rect 31297 12933 31312 12953
rect 31268 12927 31312 12933
rect 31362 12957 31411 12969
rect 31362 12937 31380 12957
rect 31400 12937 31411 12957
rect 31362 12927 31411 12937
rect 31481 12953 31525 12969
rect 31481 12933 31490 12953
rect 31510 12933 31525 12953
rect 31481 12927 31525 12933
rect 31575 12957 31624 12969
rect 31575 12937 31593 12957
rect 31613 12937 31624 12957
rect 31575 12927 31624 12937
rect 23285 12810 23303 12830
rect 23323 12810 23334 12830
rect 23285 12798 23334 12810
rect 25052 12825 25101 12835
rect 25052 12805 25063 12825
rect 25083 12805 25101 12825
rect 25052 12793 25101 12805
rect 25151 12829 25195 12835
rect 25151 12809 25166 12829
rect 25186 12809 25195 12829
rect 25151 12793 25195 12809
rect 25265 12825 25314 12835
rect 25265 12805 25276 12825
rect 25296 12805 25314 12825
rect 25265 12793 25314 12805
rect 25364 12829 25408 12835
rect 25364 12809 25379 12829
rect 25399 12809 25408 12829
rect 25364 12793 25408 12809
rect 25473 12825 25522 12835
rect 25473 12805 25484 12825
rect 25504 12805 25522 12825
rect 25473 12793 25522 12805
rect 25572 12829 25616 12835
rect 25572 12809 25587 12829
rect 25607 12809 25616 12829
rect 25572 12793 25616 12809
rect 25686 12829 25730 12835
rect 25686 12809 25695 12829
rect 25715 12809 25730 12829
rect 25686 12793 25730 12809
rect 25780 12825 25829 12835
rect 25780 12805 25798 12825
rect 25818 12805 25829 12825
rect 25780 12793 25829 12805
rect 40507 12955 40556 12967
rect 40507 12935 40518 12955
rect 40538 12935 40556 12955
rect 40507 12925 40556 12935
rect 40606 12951 40650 12967
rect 40606 12931 40621 12951
rect 40641 12931 40650 12951
rect 40606 12925 40650 12931
rect 40720 12951 40764 12967
rect 40720 12931 40729 12951
rect 40749 12931 40764 12951
rect 40720 12925 40764 12931
rect 40814 12955 40863 12967
rect 40814 12935 40832 12955
rect 40852 12935 40863 12955
rect 40814 12925 40863 12935
rect 40928 12951 40972 12967
rect 40928 12931 40937 12951
rect 40957 12931 40972 12951
rect 40928 12925 40972 12931
rect 41022 12955 41071 12967
rect 41022 12935 41040 12955
rect 41060 12935 41071 12955
rect 41022 12925 41071 12935
rect 41141 12951 41185 12967
rect 41141 12931 41150 12951
rect 41170 12931 41185 12951
rect 41141 12925 41185 12931
rect 41235 12955 41284 12967
rect 41235 12935 41253 12955
rect 41273 12935 41284 12955
rect 41235 12925 41284 12935
rect 41555 12951 41604 12963
rect 41555 12931 41566 12951
rect 41586 12931 41604 12951
rect 33265 12824 33314 12834
rect 33265 12804 33276 12824
rect 33296 12804 33314 12824
rect 33265 12792 33314 12804
rect 33364 12828 33408 12834
rect 33364 12808 33379 12828
rect 33399 12808 33408 12828
rect 33364 12792 33408 12808
rect 33478 12824 33527 12834
rect 33478 12804 33489 12824
rect 33509 12804 33527 12824
rect 33478 12792 33527 12804
rect 33577 12828 33621 12834
rect 33577 12808 33592 12828
rect 33612 12808 33621 12828
rect 33577 12792 33621 12808
rect 33686 12824 33735 12834
rect 33686 12804 33697 12824
rect 33717 12804 33735 12824
rect 33686 12792 33735 12804
rect 33785 12828 33829 12834
rect 33785 12808 33800 12828
rect 33820 12808 33829 12828
rect 33785 12792 33829 12808
rect 33899 12828 33943 12834
rect 33899 12808 33908 12828
rect 33928 12808 33943 12828
rect 33899 12792 33943 12808
rect 33993 12824 34042 12834
rect 41555 12921 41604 12931
rect 41654 12947 41698 12963
rect 41654 12927 41669 12947
rect 41689 12927 41698 12947
rect 41654 12921 41698 12927
rect 41768 12947 41812 12963
rect 41768 12927 41777 12947
rect 41797 12927 41812 12947
rect 41768 12921 41812 12927
rect 41862 12951 41911 12963
rect 41862 12931 41880 12951
rect 41900 12931 41911 12951
rect 41862 12921 41911 12931
rect 41976 12947 42020 12963
rect 41976 12927 41985 12947
rect 42005 12927 42020 12947
rect 41976 12921 42020 12927
rect 42070 12951 42119 12963
rect 42070 12931 42088 12951
rect 42108 12931 42119 12951
rect 42070 12921 42119 12931
rect 42189 12947 42233 12963
rect 42189 12927 42198 12947
rect 42218 12927 42233 12947
rect 42189 12921 42233 12927
rect 42283 12951 42332 12963
rect 42283 12931 42301 12951
rect 42321 12931 42332 12951
rect 42283 12921 42332 12931
rect 33993 12804 34011 12824
rect 34031 12804 34042 12824
rect 33993 12792 34042 12804
rect 35760 12819 35809 12829
rect 35760 12799 35771 12819
rect 35791 12799 35809 12819
rect 35760 12787 35809 12799
rect 35859 12823 35903 12829
rect 35859 12803 35874 12823
rect 35894 12803 35903 12823
rect 35859 12787 35903 12803
rect 35973 12819 36022 12829
rect 35973 12799 35984 12819
rect 36004 12799 36022 12819
rect 35973 12787 36022 12799
rect 36072 12823 36116 12829
rect 36072 12803 36087 12823
rect 36107 12803 36116 12823
rect 36072 12787 36116 12803
rect 36181 12819 36230 12829
rect 36181 12799 36192 12819
rect 36212 12799 36230 12819
rect 36181 12787 36230 12799
rect 36280 12823 36324 12829
rect 36280 12803 36295 12823
rect 36315 12803 36324 12823
rect 36280 12787 36324 12803
rect 36394 12823 36438 12829
rect 36394 12803 36403 12823
rect 36423 12803 36438 12823
rect 36394 12787 36438 12803
rect 36488 12819 36537 12829
rect 36488 12799 36506 12819
rect 36526 12799 36537 12819
rect 36488 12787 36537 12799
rect 6679 12196 6728 12208
rect 6679 12176 6690 12196
rect 6710 12176 6728 12196
rect 6679 12166 6728 12176
rect 6778 12192 6822 12208
rect 6778 12172 6793 12192
rect 6813 12172 6822 12192
rect 6778 12166 6822 12172
rect 6892 12192 6936 12208
rect 6892 12172 6901 12192
rect 6921 12172 6936 12192
rect 6892 12166 6936 12172
rect 6986 12196 7035 12208
rect 6986 12176 7004 12196
rect 7024 12176 7035 12196
rect 6986 12166 7035 12176
rect 7100 12192 7144 12208
rect 7100 12172 7109 12192
rect 7129 12172 7144 12192
rect 7100 12166 7144 12172
rect 7194 12196 7243 12208
rect 7194 12176 7212 12196
rect 7232 12176 7243 12196
rect 7194 12166 7243 12176
rect 7313 12192 7357 12208
rect 7313 12172 7322 12192
rect 7342 12172 7357 12192
rect 7313 12166 7357 12172
rect 7407 12196 7456 12208
rect 7407 12176 7425 12196
rect 7445 12176 7456 12196
rect 7407 12166 7456 12176
rect 9174 12191 9223 12203
rect 9174 12171 9185 12191
rect 9205 12171 9223 12191
rect 884 12064 933 12074
rect 884 12044 895 12064
rect 915 12044 933 12064
rect 884 12032 933 12044
rect 983 12068 1027 12074
rect 983 12048 998 12068
rect 1018 12048 1027 12068
rect 983 12032 1027 12048
rect 1097 12064 1146 12074
rect 1097 12044 1108 12064
rect 1128 12044 1146 12064
rect 1097 12032 1146 12044
rect 1196 12068 1240 12074
rect 1196 12048 1211 12068
rect 1231 12048 1240 12068
rect 1196 12032 1240 12048
rect 1305 12064 1354 12074
rect 1305 12044 1316 12064
rect 1336 12044 1354 12064
rect 1305 12032 1354 12044
rect 1404 12068 1448 12074
rect 1404 12048 1419 12068
rect 1439 12048 1448 12068
rect 1404 12032 1448 12048
rect 1518 12068 1562 12074
rect 1518 12048 1527 12068
rect 1547 12048 1562 12068
rect 1518 12032 1562 12048
rect 1612 12064 1661 12074
rect 9174 12161 9223 12171
rect 9273 12187 9317 12203
rect 9273 12167 9288 12187
rect 9308 12167 9317 12187
rect 9273 12161 9317 12167
rect 9387 12187 9431 12203
rect 9387 12167 9396 12187
rect 9416 12167 9431 12187
rect 9387 12161 9431 12167
rect 9481 12191 9530 12203
rect 9481 12171 9499 12191
rect 9519 12171 9530 12191
rect 9481 12161 9530 12171
rect 9595 12187 9639 12203
rect 9595 12167 9604 12187
rect 9624 12167 9639 12187
rect 9595 12161 9639 12167
rect 9689 12191 9738 12203
rect 9689 12171 9707 12191
rect 9727 12171 9738 12191
rect 9689 12161 9738 12171
rect 9808 12187 9852 12203
rect 9808 12167 9817 12187
rect 9837 12167 9852 12187
rect 9808 12161 9852 12167
rect 9902 12191 9951 12203
rect 9902 12171 9920 12191
rect 9940 12171 9951 12191
rect 9902 12161 9951 12171
rect 1612 12044 1630 12064
rect 1650 12044 1661 12064
rect 1612 12032 1661 12044
rect 1932 12060 1981 12070
rect 1932 12040 1943 12060
rect 1963 12040 1981 12060
rect 1932 12028 1981 12040
rect 2031 12064 2075 12070
rect 2031 12044 2046 12064
rect 2066 12044 2075 12064
rect 2031 12028 2075 12044
rect 2145 12060 2194 12070
rect 2145 12040 2156 12060
rect 2176 12040 2194 12060
rect 2145 12028 2194 12040
rect 2244 12064 2288 12070
rect 2244 12044 2259 12064
rect 2279 12044 2288 12064
rect 2244 12028 2288 12044
rect 2353 12060 2402 12070
rect 2353 12040 2364 12060
rect 2384 12040 2402 12060
rect 2353 12028 2402 12040
rect 2452 12064 2496 12070
rect 2452 12044 2467 12064
rect 2487 12044 2496 12064
rect 2452 12028 2496 12044
rect 2566 12064 2610 12070
rect 2566 12044 2575 12064
rect 2595 12044 2610 12064
rect 2566 12028 2610 12044
rect 2660 12060 2709 12070
rect 2660 12040 2678 12060
rect 2698 12040 2709 12060
rect 2660 12028 2709 12040
rect 17387 12190 17436 12202
rect 17387 12170 17398 12190
rect 17418 12170 17436 12190
rect 17387 12160 17436 12170
rect 17486 12186 17530 12202
rect 17486 12166 17501 12186
rect 17521 12166 17530 12186
rect 17486 12160 17530 12166
rect 17600 12186 17644 12202
rect 17600 12166 17609 12186
rect 17629 12166 17644 12186
rect 17600 12160 17644 12166
rect 17694 12190 17743 12202
rect 17694 12170 17712 12190
rect 17732 12170 17743 12190
rect 17694 12160 17743 12170
rect 17808 12186 17852 12202
rect 17808 12166 17817 12186
rect 17837 12166 17852 12186
rect 17808 12160 17852 12166
rect 17902 12190 17951 12202
rect 17902 12170 17920 12190
rect 17940 12170 17951 12190
rect 17902 12160 17951 12170
rect 18021 12186 18065 12202
rect 18021 12166 18030 12186
rect 18050 12166 18065 12186
rect 18021 12160 18065 12166
rect 18115 12190 18164 12202
rect 18115 12170 18133 12190
rect 18153 12170 18164 12190
rect 18115 12160 18164 12170
rect 19882 12185 19931 12197
rect 19882 12165 19893 12185
rect 19913 12165 19931 12185
rect 11592 12058 11641 12068
rect 11592 12038 11603 12058
rect 11623 12038 11641 12058
rect 11592 12026 11641 12038
rect 11691 12062 11735 12068
rect 11691 12042 11706 12062
rect 11726 12042 11735 12062
rect 11691 12026 11735 12042
rect 11805 12058 11854 12068
rect 11805 12038 11816 12058
rect 11836 12038 11854 12058
rect 11805 12026 11854 12038
rect 11904 12062 11948 12068
rect 11904 12042 11919 12062
rect 11939 12042 11948 12062
rect 11904 12026 11948 12042
rect 12013 12058 12062 12068
rect 12013 12038 12024 12058
rect 12044 12038 12062 12058
rect 12013 12026 12062 12038
rect 12112 12062 12156 12068
rect 12112 12042 12127 12062
rect 12147 12042 12156 12062
rect 12112 12026 12156 12042
rect 12226 12062 12270 12068
rect 12226 12042 12235 12062
rect 12255 12042 12270 12062
rect 12226 12026 12270 12042
rect 12320 12058 12369 12068
rect 19882 12155 19931 12165
rect 19981 12181 20025 12197
rect 19981 12161 19996 12181
rect 20016 12161 20025 12181
rect 19981 12155 20025 12161
rect 20095 12181 20139 12197
rect 20095 12161 20104 12181
rect 20124 12161 20139 12181
rect 20095 12155 20139 12161
rect 20189 12185 20238 12197
rect 20189 12165 20207 12185
rect 20227 12165 20238 12185
rect 20189 12155 20238 12165
rect 20303 12181 20347 12197
rect 20303 12161 20312 12181
rect 20332 12161 20347 12181
rect 20303 12155 20347 12161
rect 20397 12185 20446 12197
rect 20397 12165 20415 12185
rect 20435 12165 20446 12185
rect 20397 12155 20446 12165
rect 20516 12181 20560 12197
rect 20516 12161 20525 12181
rect 20545 12161 20560 12181
rect 20516 12155 20560 12161
rect 20610 12185 20659 12197
rect 20610 12165 20628 12185
rect 20648 12165 20659 12185
rect 20610 12155 20659 12165
rect 12320 12038 12338 12058
rect 12358 12038 12369 12058
rect 12320 12026 12369 12038
rect 12640 12054 12689 12064
rect 12640 12034 12651 12054
rect 12671 12034 12689 12054
rect 12640 12022 12689 12034
rect 12739 12058 12783 12064
rect 12739 12038 12754 12058
rect 12774 12038 12783 12058
rect 12739 12022 12783 12038
rect 12853 12054 12902 12064
rect 12853 12034 12864 12054
rect 12884 12034 12902 12054
rect 12853 12022 12902 12034
rect 12952 12058 12996 12064
rect 12952 12038 12967 12058
rect 12987 12038 12996 12058
rect 12952 12022 12996 12038
rect 13061 12054 13110 12064
rect 13061 12034 13072 12054
rect 13092 12034 13110 12054
rect 13061 12022 13110 12034
rect 13160 12058 13204 12064
rect 13160 12038 13175 12058
rect 13195 12038 13204 12058
rect 13160 12022 13204 12038
rect 13274 12058 13318 12064
rect 13274 12038 13283 12058
rect 13303 12038 13318 12058
rect 13274 12022 13318 12038
rect 13368 12054 13417 12064
rect 13368 12034 13386 12054
rect 13406 12034 13417 12054
rect 13368 12022 13417 12034
rect 28352 12194 28401 12206
rect 28352 12174 28363 12194
rect 28383 12174 28401 12194
rect 28352 12164 28401 12174
rect 28451 12190 28495 12206
rect 28451 12170 28466 12190
rect 28486 12170 28495 12190
rect 28451 12164 28495 12170
rect 28565 12190 28609 12206
rect 28565 12170 28574 12190
rect 28594 12170 28609 12190
rect 28565 12164 28609 12170
rect 28659 12194 28708 12206
rect 28659 12174 28677 12194
rect 28697 12174 28708 12194
rect 28659 12164 28708 12174
rect 28773 12190 28817 12206
rect 28773 12170 28782 12190
rect 28802 12170 28817 12190
rect 28773 12164 28817 12170
rect 28867 12194 28916 12206
rect 28867 12174 28885 12194
rect 28905 12174 28916 12194
rect 28867 12164 28916 12174
rect 28986 12190 29030 12206
rect 28986 12170 28995 12190
rect 29015 12170 29030 12190
rect 28986 12164 29030 12170
rect 29080 12194 29129 12206
rect 29080 12174 29098 12194
rect 29118 12174 29129 12194
rect 29080 12164 29129 12174
rect 30847 12189 30896 12201
rect 30847 12169 30858 12189
rect 30878 12169 30896 12189
rect 22557 12062 22606 12072
rect 22557 12042 22568 12062
rect 22588 12042 22606 12062
rect 22557 12030 22606 12042
rect 22656 12066 22700 12072
rect 22656 12046 22671 12066
rect 22691 12046 22700 12066
rect 22656 12030 22700 12046
rect 22770 12062 22819 12072
rect 22770 12042 22781 12062
rect 22801 12042 22819 12062
rect 22770 12030 22819 12042
rect 22869 12066 22913 12072
rect 22869 12046 22884 12066
rect 22904 12046 22913 12066
rect 22869 12030 22913 12046
rect 22978 12062 23027 12072
rect 22978 12042 22989 12062
rect 23009 12042 23027 12062
rect 22978 12030 23027 12042
rect 23077 12066 23121 12072
rect 23077 12046 23092 12066
rect 23112 12046 23121 12066
rect 23077 12030 23121 12046
rect 23191 12066 23235 12072
rect 23191 12046 23200 12066
rect 23220 12046 23235 12066
rect 23191 12030 23235 12046
rect 23285 12062 23334 12072
rect 30847 12159 30896 12169
rect 30946 12185 30990 12201
rect 30946 12165 30961 12185
rect 30981 12165 30990 12185
rect 30946 12159 30990 12165
rect 31060 12185 31104 12201
rect 31060 12165 31069 12185
rect 31089 12165 31104 12185
rect 31060 12159 31104 12165
rect 31154 12189 31203 12201
rect 31154 12169 31172 12189
rect 31192 12169 31203 12189
rect 31154 12159 31203 12169
rect 31268 12185 31312 12201
rect 31268 12165 31277 12185
rect 31297 12165 31312 12185
rect 31268 12159 31312 12165
rect 31362 12189 31411 12201
rect 31362 12169 31380 12189
rect 31400 12169 31411 12189
rect 31362 12159 31411 12169
rect 31481 12185 31525 12201
rect 31481 12165 31490 12185
rect 31510 12165 31525 12185
rect 31481 12159 31525 12165
rect 31575 12189 31624 12201
rect 31575 12169 31593 12189
rect 31613 12169 31624 12189
rect 31575 12159 31624 12169
rect 23285 12042 23303 12062
rect 23323 12042 23334 12062
rect 23285 12030 23334 12042
rect 23605 12058 23654 12068
rect 23605 12038 23616 12058
rect 23636 12038 23654 12058
rect 23605 12026 23654 12038
rect 23704 12062 23748 12068
rect 23704 12042 23719 12062
rect 23739 12042 23748 12062
rect 23704 12026 23748 12042
rect 23818 12058 23867 12068
rect 23818 12038 23829 12058
rect 23849 12038 23867 12058
rect 23818 12026 23867 12038
rect 23917 12062 23961 12068
rect 23917 12042 23932 12062
rect 23952 12042 23961 12062
rect 23917 12026 23961 12042
rect 24026 12058 24075 12068
rect 24026 12038 24037 12058
rect 24057 12038 24075 12058
rect 24026 12026 24075 12038
rect 24125 12062 24169 12068
rect 24125 12042 24140 12062
rect 24160 12042 24169 12062
rect 24125 12026 24169 12042
rect 24239 12062 24283 12068
rect 24239 12042 24248 12062
rect 24268 12042 24283 12062
rect 24239 12026 24283 12042
rect 24333 12058 24382 12068
rect 24333 12038 24351 12058
rect 24371 12038 24382 12058
rect 24333 12026 24382 12038
rect 39060 12188 39109 12200
rect 39060 12168 39071 12188
rect 39091 12168 39109 12188
rect 39060 12158 39109 12168
rect 39159 12184 39203 12200
rect 39159 12164 39174 12184
rect 39194 12164 39203 12184
rect 39159 12158 39203 12164
rect 39273 12184 39317 12200
rect 39273 12164 39282 12184
rect 39302 12164 39317 12184
rect 39273 12158 39317 12164
rect 39367 12188 39416 12200
rect 39367 12168 39385 12188
rect 39405 12168 39416 12188
rect 39367 12158 39416 12168
rect 39481 12184 39525 12200
rect 39481 12164 39490 12184
rect 39510 12164 39525 12184
rect 39481 12158 39525 12164
rect 39575 12188 39624 12200
rect 39575 12168 39593 12188
rect 39613 12168 39624 12188
rect 39575 12158 39624 12168
rect 39694 12184 39738 12200
rect 39694 12164 39703 12184
rect 39723 12164 39738 12184
rect 39694 12158 39738 12164
rect 39788 12188 39837 12200
rect 39788 12168 39806 12188
rect 39826 12168 39837 12188
rect 39788 12158 39837 12168
rect 41555 12183 41604 12195
rect 41555 12163 41566 12183
rect 41586 12163 41604 12183
rect 33265 12056 33314 12066
rect 33265 12036 33276 12056
rect 33296 12036 33314 12056
rect 33265 12024 33314 12036
rect 33364 12060 33408 12066
rect 33364 12040 33379 12060
rect 33399 12040 33408 12060
rect 33364 12024 33408 12040
rect 33478 12056 33527 12066
rect 33478 12036 33489 12056
rect 33509 12036 33527 12056
rect 33478 12024 33527 12036
rect 33577 12060 33621 12066
rect 33577 12040 33592 12060
rect 33612 12040 33621 12060
rect 33577 12024 33621 12040
rect 33686 12056 33735 12066
rect 33686 12036 33697 12056
rect 33717 12036 33735 12056
rect 33686 12024 33735 12036
rect 33785 12060 33829 12066
rect 33785 12040 33800 12060
rect 33820 12040 33829 12060
rect 33785 12024 33829 12040
rect 33899 12060 33943 12066
rect 33899 12040 33908 12060
rect 33928 12040 33943 12060
rect 33899 12024 33943 12040
rect 33993 12056 34042 12066
rect 41555 12153 41604 12163
rect 41654 12179 41698 12195
rect 41654 12159 41669 12179
rect 41689 12159 41698 12179
rect 41654 12153 41698 12159
rect 41768 12179 41812 12195
rect 41768 12159 41777 12179
rect 41797 12159 41812 12179
rect 41768 12153 41812 12159
rect 41862 12183 41911 12195
rect 41862 12163 41880 12183
rect 41900 12163 41911 12183
rect 41862 12153 41911 12163
rect 41976 12179 42020 12195
rect 41976 12159 41985 12179
rect 42005 12159 42020 12179
rect 41976 12153 42020 12159
rect 42070 12183 42119 12195
rect 42070 12163 42088 12183
rect 42108 12163 42119 12183
rect 42070 12153 42119 12163
rect 42189 12179 42233 12195
rect 42189 12159 42198 12179
rect 42218 12159 42233 12179
rect 42189 12153 42233 12159
rect 42283 12183 42332 12195
rect 42283 12163 42301 12183
rect 42321 12163 42332 12183
rect 42283 12153 42332 12163
rect 33993 12036 34011 12056
rect 34031 12036 34042 12056
rect 33993 12024 34042 12036
rect 34313 12052 34362 12062
rect 34313 12032 34324 12052
rect 34344 12032 34362 12052
rect 34313 12020 34362 12032
rect 34412 12056 34456 12062
rect 34412 12036 34427 12056
rect 34447 12036 34456 12056
rect 34412 12020 34456 12036
rect 34526 12052 34575 12062
rect 34526 12032 34537 12052
rect 34557 12032 34575 12052
rect 34526 12020 34575 12032
rect 34625 12056 34669 12062
rect 34625 12036 34640 12056
rect 34660 12036 34669 12056
rect 34625 12020 34669 12036
rect 34734 12052 34783 12062
rect 34734 12032 34745 12052
rect 34765 12032 34783 12052
rect 34734 12020 34783 12032
rect 34833 12056 34877 12062
rect 34833 12036 34848 12056
rect 34868 12036 34877 12056
rect 34833 12020 34877 12036
rect 34947 12056 34991 12062
rect 34947 12036 34956 12056
rect 34976 12036 34991 12056
rect 34947 12020 34991 12036
rect 35041 12052 35090 12062
rect 35041 12032 35059 12052
rect 35079 12032 35090 12052
rect 35041 12020 35090 12032
rect 8126 11516 8175 11528
rect 8126 11496 8137 11516
rect 8157 11496 8175 11516
rect 8126 11486 8175 11496
rect 8225 11512 8269 11528
rect 8225 11492 8240 11512
rect 8260 11492 8269 11512
rect 8225 11486 8269 11492
rect 8339 11512 8383 11528
rect 8339 11492 8348 11512
rect 8368 11492 8383 11512
rect 8339 11486 8383 11492
rect 8433 11516 8482 11528
rect 8433 11496 8451 11516
rect 8471 11496 8482 11516
rect 8433 11486 8482 11496
rect 8547 11512 8591 11528
rect 8547 11492 8556 11512
rect 8576 11492 8591 11512
rect 8547 11486 8591 11492
rect 8641 11516 8690 11528
rect 8641 11496 8659 11516
rect 8679 11496 8690 11516
rect 8641 11486 8690 11496
rect 8760 11512 8804 11528
rect 8760 11492 8769 11512
rect 8789 11492 8804 11512
rect 8760 11486 8804 11492
rect 8854 11516 8903 11528
rect 8854 11496 8872 11516
rect 8892 11496 8903 11516
rect 8854 11486 8903 11496
rect 9174 11512 9223 11524
rect 9174 11492 9185 11512
rect 9205 11492 9223 11512
rect 884 11385 933 11395
rect 884 11365 895 11385
rect 915 11365 933 11385
rect 884 11353 933 11365
rect 983 11389 1027 11395
rect 983 11369 998 11389
rect 1018 11369 1027 11389
rect 983 11353 1027 11369
rect 1097 11385 1146 11395
rect 1097 11365 1108 11385
rect 1128 11365 1146 11385
rect 1097 11353 1146 11365
rect 1196 11389 1240 11395
rect 1196 11369 1211 11389
rect 1231 11369 1240 11389
rect 1196 11353 1240 11369
rect 1305 11385 1354 11395
rect 1305 11365 1316 11385
rect 1336 11365 1354 11385
rect 1305 11353 1354 11365
rect 1404 11389 1448 11395
rect 1404 11369 1419 11389
rect 1439 11369 1448 11389
rect 1404 11353 1448 11369
rect 1518 11389 1562 11395
rect 1518 11369 1527 11389
rect 1547 11369 1562 11389
rect 1518 11353 1562 11369
rect 1612 11385 1661 11395
rect 9174 11482 9223 11492
rect 9273 11508 9317 11524
rect 9273 11488 9288 11508
rect 9308 11488 9317 11508
rect 9273 11482 9317 11488
rect 9387 11508 9431 11524
rect 9387 11488 9396 11508
rect 9416 11488 9431 11508
rect 9387 11482 9431 11488
rect 9481 11512 9530 11524
rect 9481 11492 9499 11512
rect 9519 11492 9530 11512
rect 9481 11482 9530 11492
rect 9595 11508 9639 11524
rect 9595 11488 9604 11508
rect 9624 11488 9639 11508
rect 9595 11482 9639 11488
rect 9689 11512 9738 11524
rect 9689 11492 9707 11512
rect 9727 11492 9738 11512
rect 9689 11482 9738 11492
rect 9808 11508 9852 11524
rect 9808 11488 9817 11508
rect 9837 11488 9852 11508
rect 9808 11482 9852 11488
rect 9902 11512 9951 11524
rect 9902 11492 9920 11512
rect 9940 11492 9951 11512
rect 9902 11482 9951 11492
rect 1612 11365 1630 11385
rect 1650 11365 1661 11385
rect 1612 11353 1661 11365
rect 3422 11382 3471 11392
rect 3422 11362 3433 11382
rect 3453 11362 3471 11382
rect 3422 11350 3471 11362
rect 3521 11386 3565 11392
rect 3521 11366 3536 11386
rect 3556 11366 3565 11386
rect 3521 11350 3565 11366
rect 3635 11382 3684 11392
rect 3635 11362 3646 11382
rect 3666 11362 3684 11382
rect 3635 11350 3684 11362
rect 3734 11386 3778 11392
rect 3734 11366 3749 11386
rect 3769 11366 3778 11386
rect 3734 11350 3778 11366
rect 3843 11382 3892 11392
rect 3843 11362 3854 11382
rect 3874 11362 3892 11382
rect 3843 11350 3892 11362
rect 3942 11386 3986 11392
rect 3942 11366 3957 11386
rect 3977 11366 3986 11386
rect 3942 11350 3986 11366
rect 4056 11386 4100 11392
rect 4056 11366 4065 11386
rect 4085 11366 4100 11386
rect 4056 11350 4100 11366
rect 4150 11382 4199 11392
rect 4150 11362 4168 11382
rect 4188 11362 4199 11382
rect 4150 11350 4199 11362
rect 18834 11510 18883 11522
rect 18834 11490 18845 11510
rect 18865 11490 18883 11510
rect 18834 11480 18883 11490
rect 18933 11506 18977 11522
rect 18933 11486 18948 11506
rect 18968 11486 18977 11506
rect 18933 11480 18977 11486
rect 19047 11506 19091 11522
rect 19047 11486 19056 11506
rect 19076 11486 19091 11506
rect 19047 11480 19091 11486
rect 19141 11510 19190 11522
rect 19141 11490 19159 11510
rect 19179 11490 19190 11510
rect 19141 11480 19190 11490
rect 19255 11506 19299 11522
rect 19255 11486 19264 11506
rect 19284 11486 19299 11506
rect 19255 11480 19299 11486
rect 19349 11510 19398 11522
rect 19349 11490 19367 11510
rect 19387 11490 19398 11510
rect 19349 11480 19398 11490
rect 19468 11506 19512 11522
rect 19468 11486 19477 11506
rect 19497 11486 19512 11506
rect 19468 11480 19512 11486
rect 19562 11510 19611 11522
rect 19562 11490 19580 11510
rect 19600 11490 19611 11510
rect 19562 11480 19611 11490
rect 19882 11506 19931 11518
rect 19882 11486 19893 11506
rect 19913 11486 19931 11506
rect 11592 11379 11641 11389
rect 11592 11359 11603 11379
rect 11623 11359 11641 11379
rect 11592 11347 11641 11359
rect 11691 11383 11735 11389
rect 11691 11363 11706 11383
rect 11726 11363 11735 11383
rect 11691 11347 11735 11363
rect 11805 11379 11854 11389
rect 11805 11359 11816 11379
rect 11836 11359 11854 11379
rect 11805 11347 11854 11359
rect 11904 11383 11948 11389
rect 11904 11363 11919 11383
rect 11939 11363 11948 11383
rect 11904 11347 11948 11363
rect 12013 11379 12062 11389
rect 12013 11359 12024 11379
rect 12044 11359 12062 11379
rect 12013 11347 12062 11359
rect 12112 11383 12156 11389
rect 12112 11363 12127 11383
rect 12147 11363 12156 11383
rect 12112 11347 12156 11363
rect 12226 11383 12270 11389
rect 12226 11363 12235 11383
rect 12255 11363 12270 11383
rect 12226 11347 12270 11363
rect 12320 11379 12369 11389
rect 19882 11476 19931 11486
rect 19981 11502 20025 11518
rect 19981 11482 19996 11502
rect 20016 11482 20025 11502
rect 19981 11476 20025 11482
rect 20095 11502 20139 11518
rect 20095 11482 20104 11502
rect 20124 11482 20139 11502
rect 20095 11476 20139 11482
rect 20189 11506 20238 11518
rect 20189 11486 20207 11506
rect 20227 11486 20238 11506
rect 20189 11476 20238 11486
rect 20303 11502 20347 11518
rect 20303 11482 20312 11502
rect 20332 11482 20347 11502
rect 20303 11476 20347 11482
rect 20397 11506 20446 11518
rect 20397 11486 20415 11506
rect 20435 11486 20446 11506
rect 20397 11476 20446 11486
rect 20516 11502 20560 11518
rect 20516 11482 20525 11502
rect 20545 11482 20560 11502
rect 20516 11476 20560 11482
rect 20610 11506 20659 11518
rect 20610 11486 20628 11506
rect 20648 11486 20659 11506
rect 20610 11476 20659 11486
rect 12320 11359 12338 11379
rect 12358 11359 12369 11379
rect 12320 11347 12369 11359
rect 14130 11376 14179 11386
rect 14130 11356 14141 11376
rect 14161 11356 14179 11376
rect 14130 11344 14179 11356
rect 14229 11380 14273 11386
rect 14229 11360 14244 11380
rect 14264 11360 14273 11380
rect 14229 11344 14273 11360
rect 14343 11376 14392 11386
rect 14343 11356 14354 11376
rect 14374 11356 14392 11376
rect 14343 11344 14392 11356
rect 14442 11380 14486 11386
rect 14442 11360 14457 11380
rect 14477 11360 14486 11380
rect 14442 11344 14486 11360
rect 14551 11376 14600 11386
rect 14551 11356 14562 11376
rect 14582 11356 14600 11376
rect 14551 11344 14600 11356
rect 14650 11380 14694 11386
rect 14650 11360 14665 11380
rect 14685 11360 14694 11380
rect 14650 11344 14694 11360
rect 14764 11380 14808 11386
rect 14764 11360 14773 11380
rect 14793 11360 14808 11380
rect 14764 11344 14808 11360
rect 14858 11376 14907 11386
rect 14858 11356 14876 11376
rect 14896 11356 14907 11376
rect 14858 11344 14907 11356
rect 29799 11514 29848 11526
rect 29799 11494 29810 11514
rect 29830 11494 29848 11514
rect 29799 11484 29848 11494
rect 29898 11510 29942 11526
rect 29898 11490 29913 11510
rect 29933 11490 29942 11510
rect 29898 11484 29942 11490
rect 30012 11510 30056 11526
rect 30012 11490 30021 11510
rect 30041 11490 30056 11510
rect 30012 11484 30056 11490
rect 30106 11514 30155 11526
rect 30106 11494 30124 11514
rect 30144 11494 30155 11514
rect 30106 11484 30155 11494
rect 30220 11510 30264 11526
rect 30220 11490 30229 11510
rect 30249 11490 30264 11510
rect 30220 11484 30264 11490
rect 30314 11514 30363 11526
rect 30314 11494 30332 11514
rect 30352 11494 30363 11514
rect 30314 11484 30363 11494
rect 30433 11510 30477 11526
rect 30433 11490 30442 11510
rect 30462 11490 30477 11510
rect 30433 11484 30477 11490
rect 30527 11514 30576 11526
rect 30527 11494 30545 11514
rect 30565 11494 30576 11514
rect 30527 11484 30576 11494
rect 30847 11510 30896 11522
rect 30847 11490 30858 11510
rect 30878 11490 30896 11510
rect 22557 11383 22606 11393
rect 22557 11363 22568 11383
rect 22588 11363 22606 11383
rect 22557 11351 22606 11363
rect 22656 11387 22700 11393
rect 22656 11367 22671 11387
rect 22691 11367 22700 11387
rect 22656 11351 22700 11367
rect 22770 11383 22819 11393
rect 22770 11363 22781 11383
rect 22801 11363 22819 11383
rect 22770 11351 22819 11363
rect 22869 11387 22913 11393
rect 22869 11367 22884 11387
rect 22904 11367 22913 11387
rect 22869 11351 22913 11367
rect 22978 11383 23027 11393
rect 22978 11363 22989 11383
rect 23009 11363 23027 11383
rect 22978 11351 23027 11363
rect 23077 11387 23121 11393
rect 23077 11367 23092 11387
rect 23112 11367 23121 11387
rect 23077 11351 23121 11367
rect 23191 11387 23235 11393
rect 23191 11367 23200 11387
rect 23220 11367 23235 11387
rect 23191 11351 23235 11367
rect 23285 11383 23334 11393
rect 30847 11480 30896 11490
rect 30946 11506 30990 11522
rect 30946 11486 30961 11506
rect 30981 11486 30990 11506
rect 30946 11480 30990 11486
rect 31060 11506 31104 11522
rect 31060 11486 31069 11506
rect 31089 11486 31104 11506
rect 31060 11480 31104 11486
rect 31154 11510 31203 11522
rect 31154 11490 31172 11510
rect 31192 11490 31203 11510
rect 31154 11480 31203 11490
rect 31268 11506 31312 11522
rect 31268 11486 31277 11506
rect 31297 11486 31312 11506
rect 31268 11480 31312 11486
rect 31362 11510 31411 11522
rect 31362 11490 31380 11510
rect 31400 11490 31411 11510
rect 31362 11480 31411 11490
rect 31481 11506 31525 11522
rect 31481 11486 31490 11506
rect 31510 11486 31525 11506
rect 31481 11480 31525 11486
rect 31575 11510 31624 11522
rect 31575 11490 31593 11510
rect 31613 11490 31624 11510
rect 31575 11480 31624 11490
rect 23285 11363 23303 11383
rect 23323 11363 23334 11383
rect 23285 11351 23334 11363
rect 25095 11380 25144 11390
rect 25095 11360 25106 11380
rect 25126 11360 25144 11380
rect 25095 11348 25144 11360
rect 25194 11384 25238 11390
rect 25194 11364 25209 11384
rect 25229 11364 25238 11384
rect 25194 11348 25238 11364
rect 25308 11380 25357 11390
rect 25308 11360 25319 11380
rect 25339 11360 25357 11380
rect 25308 11348 25357 11360
rect 25407 11384 25451 11390
rect 25407 11364 25422 11384
rect 25442 11364 25451 11384
rect 25407 11348 25451 11364
rect 25516 11380 25565 11390
rect 25516 11360 25527 11380
rect 25547 11360 25565 11380
rect 25516 11348 25565 11360
rect 25615 11384 25659 11390
rect 25615 11364 25630 11384
rect 25650 11364 25659 11384
rect 25615 11348 25659 11364
rect 25729 11384 25773 11390
rect 25729 11364 25738 11384
rect 25758 11364 25773 11384
rect 25729 11348 25773 11364
rect 25823 11380 25872 11390
rect 25823 11360 25841 11380
rect 25861 11360 25872 11380
rect 25823 11348 25872 11360
rect 40507 11508 40556 11520
rect 40507 11488 40518 11508
rect 40538 11488 40556 11508
rect 40507 11478 40556 11488
rect 40606 11504 40650 11520
rect 40606 11484 40621 11504
rect 40641 11484 40650 11504
rect 40606 11478 40650 11484
rect 40720 11504 40764 11520
rect 40720 11484 40729 11504
rect 40749 11484 40764 11504
rect 40720 11478 40764 11484
rect 40814 11508 40863 11520
rect 40814 11488 40832 11508
rect 40852 11488 40863 11508
rect 40814 11478 40863 11488
rect 40928 11504 40972 11520
rect 40928 11484 40937 11504
rect 40957 11484 40972 11504
rect 40928 11478 40972 11484
rect 41022 11508 41071 11520
rect 41022 11488 41040 11508
rect 41060 11488 41071 11508
rect 41022 11478 41071 11488
rect 41141 11504 41185 11520
rect 41141 11484 41150 11504
rect 41170 11484 41185 11504
rect 41141 11478 41185 11484
rect 41235 11508 41284 11520
rect 41235 11488 41253 11508
rect 41273 11488 41284 11508
rect 41235 11478 41284 11488
rect 41555 11504 41604 11516
rect 41555 11484 41566 11504
rect 41586 11484 41604 11504
rect 33265 11377 33314 11387
rect 33265 11357 33276 11377
rect 33296 11357 33314 11377
rect 33265 11345 33314 11357
rect 33364 11381 33408 11387
rect 33364 11361 33379 11381
rect 33399 11361 33408 11381
rect 33364 11345 33408 11361
rect 33478 11377 33527 11387
rect 33478 11357 33489 11377
rect 33509 11357 33527 11377
rect 33478 11345 33527 11357
rect 33577 11381 33621 11387
rect 33577 11361 33592 11381
rect 33612 11361 33621 11381
rect 33577 11345 33621 11361
rect 33686 11377 33735 11387
rect 33686 11357 33697 11377
rect 33717 11357 33735 11377
rect 33686 11345 33735 11357
rect 33785 11381 33829 11387
rect 33785 11361 33800 11381
rect 33820 11361 33829 11381
rect 33785 11345 33829 11361
rect 33899 11381 33943 11387
rect 33899 11361 33908 11381
rect 33928 11361 33943 11381
rect 33899 11345 33943 11361
rect 33993 11377 34042 11387
rect 41555 11474 41604 11484
rect 41654 11500 41698 11516
rect 41654 11480 41669 11500
rect 41689 11480 41698 11500
rect 41654 11474 41698 11480
rect 41768 11500 41812 11516
rect 41768 11480 41777 11500
rect 41797 11480 41812 11500
rect 41768 11474 41812 11480
rect 41862 11504 41911 11516
rect 41862 11484 41880 11504
rect 41900 11484 41911 11504
rect 41862 11474 41911 11484
rect 41976 11500 42020 11516
rect 41976 11480 41985 11500
rect 42005 11480 42020 11500
rect 41976 11474 42020 11480
rect 42070 11504 42119 11516
rect 42070 11484 42088 11504
rect 42108 11484 42119 11504
rect 42070 11474 42119 11484
rect 42189 11500 42233 11516
rect 42189 11480 42198 11500
rect 42218 11480 42233 11500
rect 42189 11474 42233 11480
rect 42283 11504 42332 11516
rect 42283 11484 42301 11504
rect 42321 11484 42332 11504
rect 42283 11474 42332 11484
rect 33993 11357 34011 11377
rect 34031 11357 34042 11377
rect 33993 11345 34042 11357
rect 35803 11374 35852 11384
rect 35803 11354 35814 11374
rect 35834 11354 35852 11374
rect 35803 11342 35852 11354
rect 35902 11378 35946 11384
rect 35902 11358 35917 11378
rect 35937 11358 35946 11378
rect 35902 11342 35946 11358
rect 36016 11374 36065 11384
rect 36016 11354 36027 11374
rect 36047 11354 36065 11374
rect 36016 11342 36065 11354
rect 36115 11378 36159 11384
rect 36115 11358 36130 11378
rect 36150 11358 36159 11378
rect 36115 11342 36159 11358
rect 36224 11374 36273 11384
rect 36224 11354 36235 11374
rect 36255 11354 36273 11374
rect 36224 11342 36273 11354
rect 36323 11378 36367 11384
rect 36323 11358 36338 11378
rect 36358 11358 36367 11378
rect 36323 11342 36367 11358
rect 36437 11378 36481 11384
rect 36437 11358 36446 11378
rect 36466 11358 36481 11378
rect 36437 11342 36481 11358
rect 36531 11374 36580 11384
rect 36531 11354 36549 11374
rect 36569 11354 36580 11374
rect 36531 11342 36580 11354
rect 6637 10674 6686 10686
rect 6637 10654 6648 10674
rect 6668 10654 6686 10674
rect 6637 10644 6686 10654
rect 6736 10670 6780 10686
rect 6736 10650 6751 10670
rect 6771 10650 6780 10670
rect 6736 10644 6780 10650
rect 6850 10670 6894 10686
rect 6850 10650 6859 10670
rect 6879 10650 6894 10670
rect 6850 10644 6894 10650
rect 6944 10674 6993 10686
rect 6944 10654 6962 10674
rect 6982 10654 6993 10674
rect 6944 10644 6993 10654
rect 7058 10670 7102 10686
rect 7058 10650 7067 10670
rect 7087 10650 7102 10670
rect 7058 10644 7102 10650
rect 7152 10674 7201 10686
rect 7152 10654 7170 10674
rect 7190 10654 7201 10674
rect 7152 10644 7201 10654
rect 7271 10670 7315 10686
rect 7271 10650 7280 10670
rect 7300 10650 7315 10670
rect 7271 10644 7315 10650
rect 7365 10674 7414 10686
rect 7365 10654 7383 10674
rect 7403 10654 7414 10674
rect 7365 10644 7414 10654
rect 9175 10671 9224 10683
rect 9175 10651 9186 10671
rect 9206 10651 9224 10671
rect 885 10544 934 10554
rect 885 10524 896 10544
rect 916 10524 934 10544
rect 885 10512 934 10524
rect 984 10548 1028 10554
rect 984 10528 999 10548
rect 1019 10528 1028 10548
rect 984 10512 1028 10528
rect 1098 10544 1147 10554
rect 1098 10524 1109 10544
rect 1129 10524 1147 10544
rect 1098 10512 1147 10524
rect 1197 10548 1241 10554
rect 1197 10528 1212 10548
rect 1232 10528 1241 10548
rect 1197 10512 1241 10528
rect 1306 10544 1355 10554
rect 1306 10524 1317 10544
rect 1337 10524 1355 10544
rect 1306 10512 1355 10524
rect 1405 10548 1449 10554
rect 1405 10528 1420 10548
rect 1440 10528 1449 10548
rect 1405 10512 1449 10528
rect 1519 10548 1563 10554
rect 1519 10528 1528 10548
rect 1548 10528 1563 10548
rect 1519 10512 1563 10528
rect 1613 10544 1662 10554
rect 9175 10641 9224 10651
rect 9274 10667 9318 10683
rect 9274 10647 9289 10667
rect 9309 10647 9318 10667
rect 9274 10641 9318 10647
rect 9388 10667 9432 10683
rect 9388 10647 9397 10667
rect 9417 10647 9432 10667
rect 9388 10641 9432 10647
rect 9482 10671 9531 10683
rect 9482 10651 9500 10671
rect 9520 10651 9531 10671
rect 9482 10641 9531 10651
rect 9596 10667 9640 10683
rect 9596 10647 9605 10667
rect 9625 10647 9640 10667
rect 9596 10641 9640 10647
rect 9690 10671 9739 10683
rect 9690 10651 9708 10671
rect 9728 10651 9739 10671
rect 9690 10641 9739 10651
rect 9809 10667 9853 10683
rect 9809 10647 9818 10667
rect 9838 10647 9853 10667
rect 9809 10641 9853 10647
rect 9903 10671 9952 10683
rect 9903 10651 9921 10671
rect 9941 10651 9952 10671
rect 9903 10641 9952 10651
rect 1613 10524 1631 10544
rect 1651 10524 1662 10544
rect 1613 10512 1662 10524
rect 1933 10540 1982 10550
rect 1933 10520 1944 10540
rect 1964 10520 1982 10540
rect 1933 10508 1982 10520
rect 2032 10544 2076 10550
rect 2032 10524 2047 10544
rect 2067 10524 2076 10544
rect 2032 10508 2076 10524
rect 2146 10540 2195 10550
rect 2146 10520 2157 10540
rect 2177 10520 2195 10540
rect 2146 10508 2195 10520
rect 2245 10544 2289 10550
rect 2245 10524 2260 10544
rect 2280 10524 2289 10544
rect 2245 10508 2289 10524
rect 2354 10540 2403 10550
rect 2354 10520 2365 10540
rect 2385 10520 2403 10540
rect 2354 10508 2403 10520
rect 2453 10544 2497 10550
rect 2453 10524 2468 10544
rect 2488 10524 2497 10544
rect 2453 10508 2497 10524
rect 2567 10544 2611 10550
rect 2567 10524 2576 10544
rect 2596 10524 2611 10544
rect 2567 10508 2611 10524
rect 2661 10540 2710 10550
rect 2661 10520 2679 10540
rect 2699 10520 2710 10540
rect 2661 10508 2710 10520
rect 17345 10668 17394 10680
rect 17345 10648 17356 10668
rect 17376 10648 17394 10668
rect 17345 10638 17394 10648
rect 17444 10664 17488 10680
rect 17444 10644 17459 10664
rect 17479 10644 17488 10664
rect 17444 10638 17488 10644
rect 17558 10664 17602 10680
rect 17558 10644 17567 10664
rect 17587 10644 17602 10664
rect 17558 10638 17602 10644
rect 17652 10668 17701 10680
rect 17652 10648 17670 10668
rect 17690 10648 17701 10668
rect 17652 10638 17701 10648
rect 17766 10664 17810 10680
rect 17766 10644 17775 10664
rect 17795 10644 17810 10664
rect 17766 10638 17810 10644
rect 17860 10668 17909 10680
rect 17860 10648 17878 10668
rect 17898 10648 17909 10668
rect 17860 10638 17909 10648
rect 17979 10664 18023 10680
rect 17979 10644 17988 10664
rect 18008 10644 18023 10664
rect 17979 10638 18023 10644
rect 18073 10668 18122 10680
rect 18073 10648 18091 10668
rect 18111 10648 18122 10668
rect 18073 10638 18122 10648
rect 19883 10665 19932 10677
rect 19883 10645 19894 10665
rect 19914 10645 19932 10665
rect 11593 10538 11642 10548
rect 11593 10518 11604 10538
rect 11624 10518 11642 10538
rect 11593 10506 11642 10518
rect 11692 10542 11736 10548
rect 11692 10522 11707 10542
rect 11727 10522 11736 10542
rect 11692 10506 11736 10522
rect 11806 10538 11855 10548
rect 11806 10518 11817 10538
rect 11837 10518 11855 10538
rect 11806 10506 11855 10518
rect 11905 10542 11949 10548
rect 11905 10522 11920 10542
rect 11940 10522 11949 10542
rect 11905 10506 11949 10522
rect 12014 10538 12063 10548
rect 12014 10518 12025 10538
rect 12045 10518 12063 10538
rect 12014 10506 12063 10518
rect 12113 10542 12157 10548
rect 12113 10522 12128 10542
rect 12148 10522 12157 10542
rect 12113 10506 12157 10522
rect 12227 10542 12271 10548
rect 12227 10522 12236 10542
rect 12256 10522 12271 10542
rect 12227 10506 12271 10522
rect 12321 10538 12370 10548
rect 19883 10635 19932 10645
rect 19982 10661 20026 10677
rect 19982 10641 19997 10661
rect 20017 10641 20026 10661
rect 19982 10635 20026 10641
rect 20096 10661 20140 10677
rect 20096 10641 20105 10661
rect 20125 10641 20140 10661
rect 20096 10635 20140 10641
rect 20190 10665 20239 10677
rect 20190 10645 20208 10665
rect 20228 10645 20239 10665
rect 20190 10635 20239 10645
rect 20304 10661 20348 10677
rect 20304 10641 20313 10661
rect 20333 10641 20348 10661
rect 20304 10635 20348 10641
rect 20398 10665 20447 10677
rect 20398 10645 20416 10665
rect 20436 10645 20447 10665
rect 20398 10635 20447 10645
rect 20517 10661 20561 10677
rect 20517 10641 20526 10661
rect 20546 10641 20561 10661
rect 20517 10635 20561 10641
rect 20611 10665 20660 10677
rect 20611 10645 20629 10665
rect 20649 10645 20660 10665
rect 20611 10635 20660 10645
rect 12321 10518 12339 10538
rect 12359 10518 12370 10538
rect 12321 10506 12370 10518
rect 12641 10534 12690 10544
rect 12641 10514 12652 10534
rect 12672 10514 12690 10534
rect 12641 10502 12690 10514
rect 12740 10538 12784 10544
rect 12740 10518 12755 10538
rect 12775 10518 12784 10538
rect 12740 10502 12784 10518
rect 12854 10534 12903 10544
rect 12854 10514 12865 10534
rect 12885 10514 12903 10534
rect 12854 10502 12903 10514
rect 12953 10538 12997 10544
rect 12953 10518 12968 10538
rect 12988 10518 12997 10538
rect 12953 10502 12997 10518
rect 13062 10534 13111 10544
rect 13062 10514 13073 10534
rect 13093 10514 13111 10534
rect 13062 10502 13111 10514
rect 13161 10538 13205 10544
rect 13161 10518 13176 10538
rect 13196 10518 13205 10538
rect 13161 10502 13205 10518
rect 13275 10538 13319 10544
rect 13275 10518 13284 10538
rect 13304 10518 13319 10538
rect 13275 10502 13319 10518
rect 13369 10534 13418 10544
rect 13369 10514 13387 10534
rect 13407 10514 13418 10534
rect 13369 10502 13418 10514
rect 28310 10672 28359 10684
rect 28310 10652 28321 10672
rect 28341 10652 28359 10672
rect 28310 10642 28359 10652
rect 28409 10668 28453 10684
rect 28409 10648 28424 10668
rect 28444 10648 28453 10668
rect 28409 10642 28453 10648
rect 28523 10668 28567 10684
rect 28523 10648 28532 10668
rect 28552 10648 28567 10668
rect 28523 10642 28567 10648
rect 28617 10672 28666 10684
rect 28617 10652 28635 10672
rect 28655 10652 28666 10672
rect 28617 10642 28666 10652
rect 28731 10668 28775 10684
rect 28731 10648 28740 10668
rect 28760 10648 28775 10668
rect 28731 10642 28775 10648
rect 28825 10672 28874 10684
rect 28825 10652 28843 10672
rect 28863 10652 28874 10672
rect 28825 10642 28874 10652
rect 28944 10668 28988 10684
rect 28944 10648 28953 10668
rect 28973 10648 28988 10668
rect 28944 10642 28988 10648
rect 29038 10672 29087 10684
rect 29038 10652 29056 10672
rect 29076 10652 29087 10672
rect 29038 10642 29087 10652
rect 30848 10669 30897 10681
rect 30848 10649 30859 10669
rect 30879 10649 30897 10669
rect 22558 10542 22607 10552
rect 22558 10522 22569 10542
rect 22589 10522 22607 10542
rect 22558 10510 22607 10522
rect 22657 10546 22701 10552
rect 22657 10526 22672 10546
rect 22692 10526 22701 10546
rect 22657 10510 22701 10526
rect 22771 10542 22820 10552
rect 22771 10522 22782 10542
rect 22802 10522 22820 10542
rect 22771 10510 22820 10522
rect 22870 10546 22914 10552
rect 22870 10526 22885 10546
rect 22905 10526 22914 10546
rect 22870 10510 22914 10526
rect 22979 10542 23028 10552
rect 22979 10522 22990 10542
rect 23010 10522 23028 10542
rect 22979 10510 23028 10522
rect 23078 10546 23122 10552
rect 23078 10526 23093 10546
rect 23113 10526 23122 10546
rect 23078 10510 23122 10526
rect 23192 10546 23236 10552
rect 23192 10526 23201 10546
rect 23221 10526 23236 10546
rect 23192 10510 23236 10526
rect 23286 10542 23335 10552
rect 30848 10639 30897 10649
rect 30947 10665 30991 10681
rect 30947 10645 30962 10665
rect 30982 10645 30991 10665
rect 30947 10639 30991 10645
rect 31061 10665 31105 10681
rect 31061 10645 31070 10665
rect 31090 10645 31105 10665
rect 31061 10639 31105 10645
rect 31155 10669 31204 10681
rect 31155 10649 31173 10669
rect 31193 10649 31204 10669
rect 31155 10639 31204 10649
rect 31269 10665 31313 10681
rect 31269 10645 31278 10665
rect 31298 10645 31313 10665
rect 31269 10639 31313 10645
rect 31363 10669 31412 10681
rect 31363 10649 31381 10669
rect 31401 10649 31412 10669
rect 31363 10639 31412 10649
rect 31482 10665 31526 10681
rect 31482 10645 31491 10665
rect 31511 10645 31526 10665
rect 31482 10639 31526 10645
rect 31576 10669 31625 10681
rect 31576 10649 31594 10669
rect 31614 10649 31625 10669
rect 31576 10639 31625 10649
rect 23286 10522 23304 10542
rect 23324 10522 23335 10542
rect 23286 10510 23335 10522
rect 23606 10538 23655 10548
rect 23606 10518 23617 10538
rect 23637 10518 23655 10538
rect 23606 10506 23655 10518
rect 23705 10542 23749 10548
rect 23705 10522 23720 10542
rect 23740 10522 23749 10542
rect 23705 10506 23749 10522
rect 23819 10538 23868 10548
rect 23819 10518 23830 10538
rect 23850 10518 23868 10538
rect 23819 10506 23868 10518
rect 23918 10542 23962 10548
rect 23918 10522 23933 10542
rect 23953 10522 23962 10542
rect 23918 10506 23962 10522
rect 24027 10538 24076 10548
rect 24027 10518 24038 10538
rect 24058 10518 24076 10538
rect 24027 10506 24076 10518
rect 24126 10542 24170 10548
rect 24126 10522 24141 10542
rect 24161 10522 24170 10542
rect 24126 10506 24170 10522
rect 24240 10542 24284 10548
rect 24240 10522 24249 10542
rect 24269 10522 24284 10542
rect 24240 10506 24284 10522
rect 24334 10538 24383 10548
rect 24334 10518 24352 10538
rect 24372 10518 24383 10538
rect 24334 10506 24383 10518
rect 39018 10666 39067 10678
rect 39018 10646 39029 10666
rect 39049 10646 39067 10666
rect 39018 10636 39067 10646
rect 39117 10662 39161 10678
rect 39117 10642 39132 10662
rect 39152 10642 39161 10662
rect 39117 10636 39161 10642
rect 39231 10662 39275 10678
rect 39231 10642 39240 10662
rect 39260 10642 39275 10662
rect 39231 10636 39275 10642
rect 39325 10666 39374 10678
rect 39325 10646 39343 10666
rect 39363 10646 39374 10666
rect 39325 10636 39374 10646
rect 39439 10662 39483 10678
rect 39439 10642 39448 10662
rect 39468 10642 39483 10662
rect 39439 10636 39483 10642
rect 39533 10666 39582 10678
rect 39533 10646 39551 10666
rect 39571 10646 39582 10666
rect 39533 10636 39582 10646
rect 39652 10662 39696 10678
rect 39652 10642 39661 10662
rect 39681 10642 39696 10662
rect 39652 10636 39696 10642
rect 39746 10666 39795 10678
rect 39746 10646 39764 10666
rect 39784 10646 39795 10666
rect 39746 10636 39795 10646
rect 41556 10663 41605 10675
rect 41556 10643 41567 10663
rect 41587 10643 41605 10663
rect 33266 10536 33315 10546
rect 33266 10516 33277 10536
rect 33297 10516 33315 10536
rect 33266 10504 33315 10516
rect 33365 10540 33409 10546
rect 33365 10520 33380 10540
rect 33400 10520 33409 10540
rect 33365 10504 33409 10520
rect 33479 10536 33528 10546
rect 33479 10516 33490 10536
rect 33510 10516 33528 10536
rect 33479 10504 33528 10516
rect 33578 10540 33622 10546
rect 33578 10520 33593 10540
rect 33613 10520 33622 10540
rect 33578 10504 33622 10520
rect 33687 10536 33736 10546
rect 33687 10516 33698 10536
rect 33718 10516 33736 10536
rect 33687 10504 33736 10516
rect 33786 10540 33830 10546
rect 33786 10520 33801 10540
rect 33821 10520 33830 10540
rect 33786 10504 33830 10520
rect 33900 10540 33944 10546
rect 33900 10520 33909 10540
rect 33929 10520 33944 10540
rect 33900 10504 33944 10520
rect 33994 10536 34043 10546
rect 41556 10633 41605 10643
rect 41655 10659 41699 10675
rect 41655 10639 41670 10659
rect 41690 10639 41699 10659
rect 41655 10633 41699 10639
rect 41769 10659 41813 10675
rect 41769 10639 41778 10659
rect 41798 10639 41813 10659
rect 41769 10633 41813 10639
rect 41863 10663 41912 10675
rect 41863 10643 41881 10663
rect 41901 10643 41912 10663
rect 41863 10633 41912 10643
rect 41977 10659 42021 10675
rect 41977 10639 41986 10659
rect 42006 10639 42021 10659
rect 41977 10633 42021 10639
rect 42071 10663 42120 10675
rect 42071 10643 42089 10663
rect 42109 10643 42120 10663
rect 42071 10633 42120 10643
rect 42190 10659 42234 10675
rect 42190 10639 42199 10659
rect 42219 10639 42234 10659
rect 42190 10633 42234 10639
rect 42284 10663 42333 10675
rect 42284 10643 42302 10663
rect 42322 10643 42333 10663
rect 42284 10633 42333 10643
rect 33994 10516 34012 10536
rect 34032 10516 34043 10536
rect 33994 10504 34043 10516
rect 34314 10532 34363 10542
rect 34314 10512 34325 10532
rect 34345 10512 34363 10532
rect 34314 10500 34363 10512
rect 34413 10536 34457 10542
rect 34413 10516 34428 10536
rect 34448 10516 34457 10536
rect 34413 10500 34457 10516
rect 34527 10532 34576 10542
rect 34527 10512 34538 10532
rect 34558 10512 34576 10532
rect 34527 10500 34576 10512
rect 34626 10536 34670 10542
rect 34626 10516 34641 10536
rect 34661 10516 34670 10536
rect 34626 10500 34670 10516
rect 34735 10532 34784 10542
rect 34735 10512 34746 10532
rect 34766 10512 34784 10532
rect 34735 10500 34784 10512
rect 34834 10536 34878 10542
rect 34834 10516 34849 10536
rect 34869 10516 34878 10536
rect 34834 10500 34878 10516
rect 34948 10536 34992 10542
rect 34948 10516 34957 10536
rect 34977 10516 34992 10536
rect 34948 10500 34992 10516
rect 35042 10532 35091 10542
rect 35042 10512 35060 10532
rect 35080 10512 35091 10532
rect 35042 10500 35091 10512
rect 8127 9996 8176 10008
rect 8127 9976 8138 9996
rect 8158 9976 8176 9996
rect 8127 9966 8176 9976
rect 8226 9992 8270 10008
rect 8226 9972 8241 9992
rect 8261 9972 8270 9992
rect 8226 9966 8270 9972
rect 8340 9992 8384 10008
rect 8340 9972 8349 9992
rect 8369 9972 8384 9992
rect 8340 9966 8384 9972
rect 8434 9996 8483 10008
rect 8434 9976 8452 9996
rect 8472 9976 8483 9996
rect 8434 9966 8483 9976
rect 8548 9992 8592 10008
rect 8548 9972 8557 9992
rect 8577 9972 8592 9992
rect 8548 9966 8592 9972
rect 8642 9996 8691 10008
rect 8642 9976 8660 9996
rect 8680 9976 8691 9996
rect 8642 9966 8691 9976
rect 8761 9992 8805 10008
rect 8761 9972 8770 9992
rect 8790 9972 8805 9992
rect 8761 9966 8805 9972
rect 8855 9996 8904 10008
rect 8855 9976 8873 9996
rect 8893 9976 8904 9996
rect 8855 9966 8904 9976
rect 9175 9992 9224 10004
rect 9175 9972 9186 9992
rect 9206 9972 9224 9992
rect 885 9865 934 9875
rect 885 9845 896 9865
rect 916 9845 934 9865
rect 885 9833 934 9845
rect 984 9869 1028 9875
rect 984 9849 999 9869
rect 1019 9849 1028 9869
rect 984 9833 1028 9849
rect 1098 9865 1147 9875
rect 1098 9845 1109 9865
rect 1129 9845 1147 9865
rect 1098 9833 1147 9845
rect 1197 9869 1241 9875
rect 1197 9849 1212 9869
rect 1232 9849 1241 9869
rect 1197 9833 1241 9849
rect 1306 9865 1355 9875
rect 1306 9845 1317 9865
rect 1337 9845 1355 9865
rect 1306 9833 1355 9845
rect 1405 9869 1449 9875
rect 1405 9849 1420 9869
rect 1440 9849 1449 9869
rect 1405 9833 1449 9849
rect 1519 9869 1563 9875
rect 1519 9849 1528 9869
rect 1548 9849 1563 9869
rect 1519 9833 1563 9849
rect 1613 9865 1662 9875
rect 9175 9962 9224 9972
rect 9274 9988 9318 10004
rect 9274 9968 9289 9988
rect 9309 9968 9318 9988
rect 9274 9962 9318 9968
rect 9388 9988 9432 10004
rect 9388 9968 9397 9988
rect 9417 9968 9432 9988
rect 9388 9962 9432 9968
rect 9482 9992 9531 10004
rect 9482 9972 9500 9992
rect 9520 9972 9531 9992
rect 9482 9962 9531 9972
rect 9596 9988 9640 10004
rect 9596 9968 9605 9988
rect 9625 9968 9640 9988
rect 9596 9962 9640 9968
rect 9690 9992 9739 10004
rect 9690 9972 9708 9992
rect 9728 9972 9739 9992
rect 9690 9962 9739 9972
rect 9809 9988 9853 10004
rect 9809 9968 9818 9988
rect 9838 9968 9853 9988
rect 9809 9962 9853 9968
rect 9903 9992 9952 10004
rect 9903 9972 9921 9992
rect 9941 9972 9952 9992
rect 9903 9962 9952 9972
rect 1613 9845 1631 9865
rect 1651 9845 1662 9865
rect 1613 9833 1662 9845
rect 3380 9860 3429 9870
rect 3380 9840 3391 9860
rect 3411 9840 3429 9860
rect 3380 9828 3429 9840
rect 3479 9864 3523 9870
rect 3479 9844 3494 9864
rect 3514 9844 3523 9864
rect 3479 9828 3523 9844
rect 3593 9860 3642 9870
rect 3593 9840 3604 9860
rect 3624 9840 3642 9860
rect 3593 9828 3642 9840
rect 3692 9864 3736 9870
rect 3692 9844 3707 9864
rect 3727 9844 3736 9864
rect 3692 9828 3736 9844
rect 3801 9860 3850 9870
rect 3801 9840 3812 9860
rect 3832 9840 3850 9860
rect 3801 9828 3850 9840
rect 3900 9864 3944 9870
rect 3900 9844 3915 9864
rect 3935 9844 3944 9864
rect 3900 9828 3944 9844
rect 4014 9864 4058 9870
rect 4014 9844 4023 9864
rect 4043 9844 4058 9864
rect 4014 9828 4058 9844
rect 4108 9860 4157 9870
rect 4108 9840 4126 9860
rect 4146 9840 4157 9860
rect 4108 9828 4157 9840
rect 18835 9990 18884 10002
rect 18835 9970 18846 9990
rect 18866 9970 18884 9990
rect 18835 9960 18884 9970
rect 18934 9986 18978 10002
rect 18934 9966 18949 9986
rect 18969 9966 18978 9986
rect 18934 9960 18978 9966
rect 19048 9986 19092 10002
rect 19048 9966 19057 9986
rect 19077 9966 19092 9986
rect 19048 9960 19092 9966
rect 19142 9990 19191 10002
rect 19142 9970 19160 9990
rect 19180 9970 19191 9990
rect 19142 9960 19191 9970
rect 19256 9986 19300 10002
rect 19256 9966 19265 9986
rect 19285 9966 19300 9986
rect 19256 9960 19300 9966
rect 19350 9990 19399 10002
rect 19350 9970 19368 9990
rect 19388 9970 19399 9990
rect 19350 9960 19399 9970
rect 19469 9986 19513 10002
rect 19469 9966 19478 9986
rect 19498 9966 19513 9986
rect 19469 9960 19513 9966
rect 19563 9990 19612 10002
rect 19563 9970 19581 9990
rect 19601 9970 19612 9990
rect 19563 9960 19612 9970
rect 19883 9986 19932 9998
rect 19883 9966 19894 9986
rect 19914 9966 19932 9986
rect 11593 9859 11642 9869
rect 11593 9839 11604 9859
rect 11624 9839 11642 9859
rect 11593 9827 11642 9839
rect 11692 9863 11736 9869
rect 11692 9843 11707 9863
rect 11727 9843 11736 9863
rect 11692 9827 11736 9843
rect 11806 9859 11855 9869
rect 11806 9839 11817 9859
rect 11837 9839 11855 9859
rect 11806 9827 11855 9839
rect 11905 9863 11949 9869
rect 11905 9843 11920 9863
rect 11940 9843 11949 9863
rect 11905 9827 11949 9843
rect 12014 9859 12063 9869
rect 12014 9839 12025 9859
rect 12045 9839 12063 9859
rect 12014 9827 12063 9839
rect 12113 9863 12157 9869
rect 12113 9843 12128 9863
rect 12148 9843 12157 9863
rect 12113 9827 12157 9843
rect 12227 9863 12271 9869
rect 12227 9843 12236 9863
rect 12256 9843 12271 9863
rect 12227 9827 12271 9843
rect 12321 9859 12370 9869
rect 19883 9956 19932 9966
rect 19982 9982 20026 9998
rect 19982 9962 19997 9982
rect 20017 9962 20026 9982
rect 19982 9956 20026 9962
rect 20096 9982 20140 9998
rect 20096 9962 20105 9982
rect 20125 9962 20140 9982
rect 20096 9956 20140 9962
rect 20190 9986 20239 9998
rect 20190 9966 20208 9986
rect 20228 9966 20239 9986
rect 20190 9956 20239 9966
rect 20304 9982 20348 9998
rect 20304 9962 20313 9982
rect 20333 9962 20348 9982
rect 20304 9956 20348 9962
rect 20398 9986 20447 9998
rect 20398 9966 20416 9986
rect 20436 9966 20447 9986
rect 20398 9956 20447 9966
rect 20517 9982 20561 9998
rect 20517 9962 20526 9982
rect 20546 9962 20561 9982
rect 20517 9956 20561 9962
rect 20611 9986 20660 9998
rect 20611 9966 20629 9986
rect 20649 9966 20660 9986
rect 20611 9956 20660 9966
rect 12321 9839 12339 9859
rect 12359 9839 12370 9859
rect 12321 9827 12370 9839
rect 14088 9854 14137 9864
rect 14088 9834 14099 9854
rect 14119 9834 14137 9854
rect 14088 9822 14137 9834
rect 14187 9858 14231 9864
rect 14187 9838 14202 9858
rect 14222 9838 14231 9858
rect 14187 9822 14231 9838
rect 14301 9854 14350 9864
rect 14301 9834 14312 9854
rect 14332 9834 14350 9854
rect 14301 9822 14350 9834
rect 14400 9858 14444 9864
rect 14400 9838 14415 9858
rect 14435 9838 14444 9858
rect 14400 9822 14444 9838
rect 14509 9854 14558 9864
rect 14509 9834 14520 9854
rect 14540 9834 14558 9854
rect 14509 9822 14558 9834
rect 14608 9858 14652 9864
rect 14608 9838 14623 9858
rect 14643 9838 14652 9858
rect 14608 9822 14652 9838
rect 14722 9858 14766 9864
rect 14722 9838 14731 9858
rect 14751 9838 14766 9858
rect 14722 9822 14766 9838
rect 14816 9854 14865 9864
rect 14816 9834 14834 9854
rect 14854 9834 14865 9854
rect 14816 9822 14865 9834
rect 29800 9994 29849 10006
rect 29800 9974 29811 9994
rect 29831 9974 29849 9994
rect 29800 9964 29849 9974
rect 29899 9990 29943 10006
rect 29899 9970 29914 9990
rect 29934 9970 29943 9990
rect 29899 9964 29943 9970
rect 30013 9990 30057 10006
rect 30013 9970 30022 9990
rect 30042 9970 30057 9990
rect 30013 9964 30057 9970
rect 30107 9994 30156 10006
rect 30107 9974 30125 9994
rect 30145 9974 30156 9994
rect 30107 9964 30156 9974
rect 30221 9990 30265 10006
rect 30221 9970 30230 9990
rect 30250 9970 30265 9990
rect 30221 9964 30265 9970
rect 30315 9994 30364 10006
rect 30315 9974 30333 9994
rect 30353 9974 30364 9994
rect 30315 9964 30364 9974
rect 30434 9990 30478 10006
rect 30434 9970 30443 9990
rect 30463 9970 30478 9990
rect 30434 9964 30478 9970
rect 30528 9994 30577 10006
rect 30528 9974 30546 9994
rect 30566 9974 30577 9994
rect 30528 9964 30577 9974
rect 30848 9990 30897 10002
rect 30848 9970 30859 9990
rect 30879 9970 30897 9990
rect 22558 9863 22607 9873
rect 22558 9843 22569 9863
rect 22589 9843 22607 9863
rect 22558 9831 22607 9843
rect 22657 9867 22701 9873
rect 22657 9847 22672 9867
rect 22692 9847 22701 9867
rect 22657 9831 22701 9847
rect 22771 9863 22820 9873
rect 22771 9843 22782 9863
rect 22802 9843 22820 9863
rect 22771 9831 22820 9843
rect 22870 9867 22914 9873
rect 22870 9847 22885 9867
rect 22905 9847 22914 9867
rect 22870 9831 22914 9847
rect 22979 9863 23028 9873
rect 22979 9843 22990 9863
rect 23010 9843 23028 9863
rect 22979 9831 23028 9843
rect 23078 9867 23122 9873
rect 23078 9847 23093 9867
rect 23113 9847 23122 9867
rect 23078 9831 23122 9847
rect 23192 9867 23236 9873
rect 23192 9847 23201 9867
rect 23221 9847 23236 9867
rect 23192 9831 23236 9847
rect 23286 9863 23335 9873
rect 30848 9960 30897 9970
rect 30947 9986 30991 10002
rect 30947 9966 30962 9986
rect 30982 9966 30991 9986
rect 30947 9960 30991 9966
rect 31061 9986 31105 10002
rect 31061 9966 31070 9986
rect 31090 9966 31105 9986
rect 31061 9960 31105 9966
rect 31155 9990 31204 10002
rect 31155 9970 31173 9990
rect 31193 9970 31204 9990
rect 31155 9960 31204 9970
rect 31269 9986 31313 10002
rect 31269 9966 31278 9986
rect 31298 9966 31313 9986
rect 31269 9960 31313 9966
rect 31363 9990 31412 10002
rect 31363 9970 31381 9990
rect 31401 9970 31412 9990
rect 31363 9960 31412 9970
rect 31482 9986 31526 10002
rect 31482 9966 31491 9986
rect 31511 9966 31526 9986
rect 31482 9960 31526 9966
rect 31576 9990 31625 10002
rect 31576 9970 31594 9990
rect 31614 9970 31625 9990
rect 31576 9960 31625 9970
rect 23286 9843 23304 9863
rect 23324 9843 23335 9863
rect 23286 9831 23335 9843
rect 25053 9858 25102 9868
rect 25053 9838 25064 9858
rect 25084 9838 25102 9858
rect 25053 9826 25102 9838
rect 25152 9862 25196 9868
rect 25152 9842 25167 9862
rect 25187 9842 25196 9862
rect 25152 9826 25196 9842
rect 25266 9858 25315 9868
rect 25266 9838 25277 9858
rect 25297 9838 25315 9858
rect 25266 9826 25315 9838
rect 25365 9862 25409 9868
rect 25365 9842 25380 9862
rect 25400 9842 25409 9862
rect 25365 9826 25409 9842
rect 25474 9858 25523 9868
rect 25474 9838 25485 9858
rect 25505 9838 25523 9858
rect 25474 9826 25523 9838
rect 25573 9862 25617 9868
rect 25573 9842 25588 9862
rect 25608 9842 25617 9862
rect 25573 9826 25617 9842
rect 25687 9862 25731 9868
rect 25687 9842 25696 9862
rect 25716 9842 25731 9862
rect 25687 9826 25731 9842
rect 25781 9858 25830 9868
rect 25781 9838 25799 9858
rect 25819 9838 25830 9858
rect 25781 9826 25830 9838
rect 40508 9988 40557 10000
rect 40508 9968 40519 9988
rect 40539 9968 40557 9988
rect 40508 9958 40557 9968
rect 40607 9984 40651 10000
rect 40607 9964 40622 9984
rect 40642 9964 40651 9984
rect 40607 9958 40651 9964
rect 40721 9984 40765 10000
rect 40721 9964 40730 9984
rect 40750 9964 40765 9984
rect 40721 9958 40765 9964
rect 40815 9988 40864 10000
rect 40815 9968 40833 9988
rect 40853 9968 40864 9988
rect 40815 9958 40864 9968
rect 40929 9984 40973 10000
rect 40929 9964 40938 9984
rect 40958 9964 40973 9984
rect 40929 9958 40973 9964
rect 41023 9988 41072 10000
rect 41023 9968 41041 9988
rect 41061 9968 41072 9988
rect 41023 9958 41072 9968
rect 41142 9984 41186 10000
rect 41142 9964 41151 9984
rect 41171 9964 41186 9984
rect 41142 9958 41186 9964
rect 41236 9988 41285 10000
rect 41236 9968 41254 9988
rect 41274 9968 41285 9988
rect 41236 9958 41285 9968
rect 41556 9984 41605 9996
rect 41556 9964 41567 9984
rect 41587 9964 41605 9984
rect 33266 9857 33315 9867
rect 33266 9837 33277 9857
rect 33297 9837 33315 9857
rect 33266 9825 33315 9837
rect 33365 9861 33409 9867
rect 33365 9841 33380 9861
rect 33400 9841 33409 9861
rect 33365 9825 33409 9841
rect 33479 9857 33528 9867
rect 33479 9837 33490 9857
rect 33510 9837 33528 9857
rect 33479 9825 33528 9837
rect 33578 9861 33622 9867
rect 33578 9841 33593 9861
rect 33613 9841 33622 9861
rect 33578 9825 33622 9841
rect 33687 9857 33736 9867
rect 33687 9837 33698 9857
rect 33718 9837 33736 9857
rect 33687 9825 33736 9837
rect 33786 9861 33830 9867
rect 33786 9841 33801 9861
rect 33821 9841 33830 9861
rect 33786 9825 33830 9841
rect 33900 9861 33944 9867
rect 33900 9841 33909 9861
rect 33929 9841 33944 9861
rect 33900 9825 33944 9841
rect 33994 9857 34043 9867
rect 41556 9954 41605 9964
rect 41655 9980 41699 9996
rect 41655 9960 41670 9980
rect 41690 9960 41699 9980
rect 41655 9954 41699 9960
rect 41769 9980 41813 9996
rect 41769 9960 41778 9980
rect 41798 9960 41813 9980
rect 41769 9954 41813 9960
rect 41863 9984 41912 9996
rect 41863 9964 41881 9984
rect 41901 9964 41912 9984
rect 41863 9954 41912 9964
rect 41977 9980 42021 9996
rect 41977 9960 41986 9980
rect 42006 9960 42021 9980
rect 41977 9954 42021 9960
rect 42071 9984 42120 9996
rect 42071 9964 42089 9984
rect 42109 9964 42120 9984
rect 42071 9954 42120 9964
rect 42190 9980 42234 9996
rect 42190 9960 42199 9980
rect 42219 9960 42234 9980
rect 42190 9954 42234 9960
rect 42284 9984 42333 9996
rect 42284 9964 42302 9984
rect 42322 9964 42333 9984
rect 42284 9954 42333 9964
rect 33994 9837 34012 9857
rect 34032 9837 34043 9857
rect 33994 9825 34043 9837
rect 35761 9852 35810 9862
rect 35761 9832 35772 9852
rect 35792 9832 35810 9852
rect 35761 9820 35810 9832
rect 35860 9856 35904 9862
rect 35860 9836 35875 9856
rect 35895 9836 35904 9856
rect 35860 9820 35904 9836
rect 35974 9852 36023 9862
rect 35974 9832 35985 9852
rect 36005 9832 36023 9852
rect 35974 9820 36023 9832
rect 36073 9856 36117 9862
rect 36073 9836 36088 9856
rect 36108 9836 36117 9856
rect 36073 9820 36117 9836
rect 36182 9852 36231 9862
rect 36182 9832 36193 9852
rect 36213 9832 36231 9852
rect 36182 9820 36231 9832
rect 36281 9856 36325 9862
rect 36281 9836 36296 9856
rect 36316 9836 36325 9856
rect 36281 9820 36325 9836
rect 36395 9856 36439 9862
rect 36395 9836 36404 9856
rect 36424 9836 36439 9856
rect 36395 9820 36439 9836
rect 36489 9852 36538 9862
rect 36489 9832 36507 9852
rect 36527 9832 36538 9852
rect 36489 9820 36538 9832
rect 6680 9229 6729 9241
rect 6680 9209 6691 9229
rect 6711 9209 6729 9229
rect 6680 9199 6729 9209
rect 6779 9225 6823 9241
rect 6779 9205 6794 9225
rect 6814 9205 6823 9225
rect 6779 9199 6823 9205
rect 6893 9225 6937 9241
rect 6893 9205 6902 9225
rect 6922 9205 6937 9225
rect 6893 9199 6937 9205
rect 6987 9229 7036 9241
rect 6987 9209 7005 9229
rect 7025 9209 7036 9229
rect 6987 9199 7036 9209
rect 7101 9225 7145 9241
rect 7101 9205 7110 9225
rect 7130 9205 7145 9225
rect 7101 9199 7145 9205
rect 7195 9229 7244 9241
rect 7195 9209 7213 9229
rect 7233 9209 7244 9229
rect 7195 9199 7244 9209
rect 7314 9225 7358 9241
rect 7314 9205 7323 9225
rect 7343 9205 7358 9225
rect 7314 9199 7358 9205
rect 7408 9229 7457 9241
rect 7408 9209 7426 9229
rect 7446 9209 7457 9229
rect 7408 9199 7457 9209
rect 9175 9224 9224 9236
rect 9175 9204 9186 9224
rect 9206 9204 9224 9224
rect 885 9097 934 9107
rect 885 9077 896 9097
rect 916 9077 934 9097
rect 885 9065 934 9077
rect 984 9101 1028 9107
rect 984 9081 999 9101
rect 1019 9081 1028 9101
rect 984 9065 1028 9081
rect 1098 9097 1147 9107
rect 1098 9077 1109 9097
rect 1129 9077 1147 9097
rect 1098 9065 1147 9077
rect 1197 9101 1241 9107
rect 1197 9081 1212 9101
rect 1232 9081 1241 9101
rect 1197 9065 1241 9081
rect 1306 9097 1355 9107
rect 1306 9077 1317 9097
rect 1337 9077 1355 9097
rect 1306 9065 1355 9077
rect 1405 9101 1449 9107
rect 1405 9081 1420 9101
rect 1440 9081 1449 9101
rect 1405 9065 1449 9081
rect 1519 9101 1563 9107
rect 1519 9081 1528 9101
rect 1548 9081 1563 9101
rect 1519 9065 1563 9081
rect 1613 9097 1662 9107
rect 9175 9194 9224 9204
rect 9274 9220 9318 9236
rect 9274 9200 9289 9220
rect 9309 9200 9318 9220
rect 9274 9194 9318 9200
rect 9388 9220 9432 9236
rect 9388 9200 9397 9220
rect 9417 9200 9432 9220
rect 9388 9194 9432 9200
rect 9482 9224 9531 9236
rect 9482 9204 9500 9224
rect 9520 9204 9531 9224
rect 9482 9194 9531 9204
rect 9596 9220 9640 9236
rect 9596 9200 9605 9220
rect 9625 9200 9640 9220
rect 9596 9194 9640 9200
rect 9690 9224 9739 9236
rect 9690 9204 9708 9224
rect 9728 9204 9739 9224
rect 9690 9194 9739 9204
rect 9809 9220 9853 9236
rect 9809 9200 9818 9220
rect 9838 9200 9853 9220
rect 9809 9194 9853 9200
rect 9903 9224 9952 9236
rect 9903 9204 9921 9224
rect 9941 9204 9952 9224
rect 9903 9194 9952 9204
rect 1613 9077 1631 9097
rect 1651 9077 1662 9097
rect 1613 9065 1662 9077
rect 1933 9093 1982 9103
rect 1933 9073 1944 9093
rect 1964 9073 1982 9093
rect 1933 9061 1982 9073
rect 2032 9097 2076 9103
rect 2032 9077 2047 9097
rect 2067 9077 2076 9097
rect 2032 9061 2076 9077
rect 2146 9093 2195 9103
rect 2146 9073 2157 9093
rect 2177 9073 2195 9093
rect 2146 9061 2195 9073
rect 2245 9097 2289 9103
rect 2245 9077 2260 9097
rect 2280 9077 2289 9097
rect 2245 9061 2289 9077
rect 2354 9093 2403 9103
rect 2354 9073 2365 9093
rect 2385 9073 2403 9093
rect 2354 9061 2403 9073
rect 2453 9097 2497 9103
rect 2453 9077 2468 9097
rect 2488 9077 2497 9097
rect 2453 9061 2497 9077
rect 2567 9097 2611 9103
rect 2567 9077 2576 9097
rect 2596 9077 2611 9097
rect 2567 9061 2611 9077
rect 2661 9093 2710 9103
rect 2661 9073 2679 9093
rect 2699 9073 2710 9093
rect 2661 9061 2710 9073
rect 17388 9223 17437 9235
rect 17388 9203 17399 9223
rect 17419 9203 17437 9223
rect 17388 9193 17437 9203
rect 17487 9219 17531 9235
rect 17487 9199 17502 9219
rect 17522 9199 17531 9219
rect 17487 9193 17531 9199
rect 17601 9219 17645 9235
rect 17601 9199 17610 9219
rect 17630 9199 17645 9219
rect 17601 9193 17645 9199
rect 17695 9223 17744 9235
rect 17695 9203 17713 9223
rect 17733 9203 17744 9223
rect 17695 9193 17744 9203
rect 17809 9219 17853 9235
rect 17809 9199 17818 9219
rect 17838 9199 17853 9219
rect 17809 9193 17853 9199
rect 17903 9223 17952 9235
rect 17903 9203 17921 9223
rect 17941 9203 17952 9223
rect 17903 9193 17952 9203
rect 18022 9219 18066 9235
rect 18022 9199 18031 9219
rect 18051 9199 18066 9219
rect 18022 9193 18066 9199
rect 18116 9223 18165 9235
rect 18116 9203 18134 9223
rect 18154 9203 18165 9223
rect 18116 9193 18165 9203
rect 19883 9218 19932 9230
rect 19883 9198 19894 9218
rect 19914 9198 19932 9218
rect 11593 9091 11642 9101
rect 11593 9071 11604 9091
rect 11624 9071 11642 9091
rect 11593 9059 11642 9071
rect 11692 9095 11736 9101
rect 11692 9075 11707 9095
rect 11727 9075 11736 9095
rect 11692 9059 11736 9075
rect 11806 9091 11855 9101
rect 11806 9071 11817 9091
rect 11837 9071 11855 9091
rect 11806 9059 11855 9071
rect 11905 9095 11949 9101
rect 11905 9075 11920 9095
rect 11940 9075 11949 9095
rect 11905 9059 11949 9075
rect 12014 9091 12063 9101
rect 12014 9071 12025 9091
rect 12045 9071 12063 9091
rect 12014 9059 12063 9071
rect 12113 9095 12157 9101
rect 12113 9075 12128 9095
rect 12148 9075 12157 9095
rect 12113 9059 12157 9075
rect 12227 9095 12271 9101
rect 12227 9075 12236 9095
rect 12256 9075 12271 9095
rect 12227 9059 12271 9075
rect 12321 9091 12370 9101
rect 19883 9188 19932 9198
rect 19982 9214 20026 9230
rect 19982 9194 19997 9214
rect 20017 9194 20026 9214
rect 19982 9188 20026 9194
rect 20096 9214 20140 9230
rect 20096 9194 20105 9214
rect 20125 9194 20140 9214
rect 20096 9188 20140 9194
rect 20190 9218 20239 9230
rect 20190 9198 20208 9218
rect 20228 9198 20239 9218
rect 20190 9188 20239 9198
rect 20304 9214 20348 9230
rect 20304 9194 20313 9214
rect 20333 9194 20348 9214
rect 20304 9188 20348 9194
rect 20398 9218 20447 9230
rect 20398 9198 20416 9218
rect 20436 9198 20447 9218
rect 20398 9188 20447 9198
rect 20517 9214 20561 9230
rect 20517 9194 20526 9214
rect 20546 9194 20561 9214
rect 20517 9188 20561 9194
rect 20611 9218 20660 9230
rect 20611 9198 20629 9218
rect 20649 9198 20660 9218
rect 20611 9188 20660 9198
rect 12321 9071 12339 9091
rect 12359 9071 12370 9091
rect 12321 9059 12370 9071
rect 12641 9087 12690 9097
rect 12641 9067 12652 9087
rect 12672 9067 12690 9087
rect 12641 9055 12690 9067
rect 12740 9091 12784 9097
rect 12740 9071 12755 9091
rect 12775 9071 12784 9091
rect 12740 9055 12784 9071
rect 12854 9087 12903 9097
rect 12854 9067 12865 9087
rect 12885 9067 12903 9087
rect 12854 9055 12903 9067
rect 12953 9091 12997 9097
rect 12953 9071 12968 9091
rect 12988 9071 12997 9091
rect 12953 9055 12997 9071
rect 13062 9087 13111 9097
rect 13062 9067 13073 9087
rect 13093 9067 13111 9087
rect 13062 9055 13111 9067
rect 13161 9091 13205 9097
rect 13161 9071 13176 9091
rect 13196 9071 13205 9091
rect 13161 9055 13205 9071
rect 13275 9091 13319 9097
rect 13275 9071 13284 9091
rect 13304 9071 13319 9091
rect 13275 9055 13319 9071
rect 13369 9087 13418 9097
rect 13369 9067 13387 9087
rect 13407 9067 13418 9087
rect 13369 9055 13418 9067
rect 28353 9227 28402 9239
rect 28353 9207 28364 9227
rect 28384 9207 28402 9227
rect 28353 9197 28402 9207
rect 28452 9223 28496 9239
rect 28452 9203 28467 9223
rect 28487 9203 28496 9223
rect 28452 9197 28496 9203
rect 28566 9223 28610 9239
rect 28566 9203 28575 9223
rect 28595 9203 28610 9223
rect 28566 9197 28610 9203
rect 28660 9227 28709 9239
rect 28660 9207 28678 9227
rect 28698 9207 28709 9227
rect 28660 9197 28709 9207
rect 28774 9223 28818 9239
rect 28774 9203 28783 9223
rect 28803 9203 28818 9223
rect 28774 9197 28818 9203
rect 28868 9227 28917 9239
rect 28868 9207 28886 9227
rect 28906 9207 28917 9227
rect 28868 9197 28917 9207
rect 28987 9223 29031 9239
rect 28987 9203 28996 9223
rect 29016 9203 29031 9223
rect 28987 9197 29031 9203
rect 29081 9227 29130 9239
rect 29081 9207 29099 9227
rect 29119 9207 29130 9227
rect 29081 9197 29130 9207
rect 30848 9222 30897 9234
rect 30848 9202 30859 9222
rect 30879 9202 30897 9222
rect 22558 9095 22607 9105
rect 22558 9075 22569 9095
rect 22589 9075 22607 9095
rect 22558 9063 22607 9075
rect 22657 9099 22701 9105
rect 22657 9079 22672 9099
rect 22692 9079 22701 9099
rect 22657 9063 22701 9079
rect 22771 9095 22820 9105
rect 22771 9075 22782 9095
rect 22802 9075 22820 9095
rect 22771 9063 22820 9075
rect 22870 9099 22914 9105
rect 22870 9079 22885 9099
rect 22905 9079 22914 9099
rect 22870 9063 22914 9079
rect 22979 9095 23028 9105
rect 22979 9075 22990 9095
rect 23010 9075 23028 9095
rect 22979 9063 23028 9075
rect 23078 9099 23122 9105
rect 23078 9079 23093 9099
rect 23113 9079 23122 9099
rect 23078 9063 23122 9079
rect 23192 9099 23236 9105
rect 23192 9079 23201 9099
rect 23221 9079 23236 9099
rect 23192 9063 23236 9079
rect 23286 9095 23335 9105
rect 30848 9192 30897 9202
rect 30947 9218 30991 9234
rect 30947 9198 30962 9218
rect 30982 9198 30991 9218
rect 30947 9192 30991 9198
rect 31061 9218 31105 9234
rect 31061 9198 31070 9218
rect 31090 9198 31105 9218
rect 31061 9192 31105 9198
rect 31155 9222 31204 9234
rect 31155 9202 31173 9222
rect 31193 9202 31204 9222
rect 31155 9192 31204 9202
rect 31269 9218 31313 9234
rect 31269 9198 31278 9218
rect 31298 9198 31313 9218
rect 31269 9192 31313 9198
rect 31363 9222 31412 9234
rect 31363 9202 31381 9222
rect 31401 9202 31412 9222
rect 31363 9192 31412 9202
rect 31482 9218 31526 9234
rect 31482 9198 31491 9218
rect 31511 9198 31526 9218
rect 31482 9192 31526 9198
rect 31576 9222 31625 9234
rect 31576 9202 31594 9222
rect 31614 9202 31625 9222
rect 31576 9192 31625 9202
rect 23286 9075 23304 9095
rect 23324 9075 23335 9095
rect 23286 9063 23335 9075
rect 23606 9091 23655 9101
rect 23606 9071 23617 9091
rect 23637 9071 23655 9091
rect 23606 9059 23655 9071
rect 23705 9095 23749 9101
rect 23705 9075 23720 9095
rect 23740 9075 23749 9095
rect 23705 9059 23749 9075
rect 23819 9091 23868 9101
rect 23819 9071 23830 9091
rect 23850 9071 23868 9091
rect 23819 9059 23868 9071
rect 23918 9095 23962 9101
rect 23918 9075 23933 9095
rect 23953 9075 23962 9095
rect 23918 9059 23962 9075
rect 24027 9091 24076 9101
rect 24027 9071 24038 9091
rect 24058 9071 24076 9091
rect 24027 9059 24076 9071
rect 24126 9095 24170 9101
rect 24126 9075 24141 9095
rect 24161 9075 24170 9095
rect 24126 9059 24170 9075
rect 24240 9095 24284 9101
rect 24240 9075 24249 9095
rect 24269 9075 24284 9095
rect 24240 9059 24284 9075
rect 24334 9091 24383 9101
rect 24334 9071 24352 9091
rect 24372 9071 24383 9091
rect 24334 9059 24383 9071
rect 39061 9221 39110 9233
rect 39061 9201 39072 9221
rect 39092 9201 39110 9221
rect 39061 9191 39110 9201
rect 39160 9217 39204 9233
rect 39160 9197 39175 9217
rect 39195 9197 39204 9217
rect 39160 9191 39204 9197
rect 39274 9217 39318 9233
rect 39274 9197 39283 9217
rect 39303 9197 39318 9217
rect 39274 9191 39318 9197
rect 39368 9221 39417 9233
rect 39368 9201 39386 9221
rect 39406 9201 39417 9221
rect 39368 9191 39417 9201
rect 39482 9217 39526 9233
rect 39482 9197 39491 9217
rect 39511 9197 39526 9217
rect 39482 9191 39526 9197
rect 39576 9221 39625 9233
rect 39576 9201 39594 9221
rect 39614 9201 39625 9221
rect 39576 9191 39625 9201
rect 39695 9217 39739 9233
rect 39695 9197 39704 9217
rect 39724 9197 39739 9217
rect 39695 9191 39739 9197
rect 39789 9221 39838 9233
rect 39789 9201 39807 9221
rect 39827 9201 39838 9221
rect 39789 9191 39838 9201
rect 41556 9216 41605 9228
rect 41556 9196 41567 9216
rect 41587 9196 41605 9216
rect 33266 9089 33315 9099
rect 33266 9069 33277 9089
rect 33297 9069 33315 9089
rect 33266 9057 33315 9069
rect 33365 9093 33409 9099
rect 33365 9073 33380 9093
rect 33400 9073 33409 9093
rect 33365 9057 33409 9073
rect 33479 9089 33528 9099
rect 33479 9069 33490 9089
rect 33510 9069 33528 9089
rect 33479 9057 33528 9069
rect 33578 9093 33622 9099
rect 33578 9073 33593 9093
rect 33613 9073 33622 9093
rect 33578 9057 33622 9073
rect 33687 9089 33736 9099
rect 33687 9069 33698 9089
rect 33718 9069 33736 9089
rect 33687 9057 33736 9069
rect 33786 9093 33830 9099
rect 33786 9073 33801 9093
rect 33821 9073 33830 9093
rect 33786 9057 33830 9073
rect 33900 9093 33944 9099
rect 33900 9073 33909 9093
rect 33929 9073 33944 9093
rect 33900 9057 33944 9073
rect 33994 9089 34043 9099
rect 41556 9186 41605 9196
rect 41655 9212 41699 9228
rect 41655 9192 41670 9212
rect 41690 9192 41699 9212
rect 41655 9186 41699 9192
rect 41769 9212 41813 9228
rect 41769 9192 41778 9212
rect 41798 9192 41813 9212
rect 41769 9186 41813 9192
rect 41863 9216 41912 9228
rect 41863 9196 41881 9216
rect 41901 9196 41912 9216
rect 41863 9186 41912 9196
rect 41977 9212 42021 9228
rect 41977 9192 41986 9212
rect 42006 9192 42021 9212
rect 41977 9186 42021 9192
rect 42071 9216 42120 9228
rect 42071 9196 42089 9216
rect 42109 9196 42120 9216
rect 42071 9186 42120 9196
rect 42190 9212 42234 9228
rect 42190 9192 42199 9212
rect 42219 9192 42234 9212
rect 42190 9186 42234 9192
rect 42284 9216 42333 9228
rect 42284 9196 42302 9216
rect 42322 9196 42333 9216
rect 42284 9186 42333 9196
rect 33994 9069 34012 9089
rect 34032 9069 34043 9089
rect 33994 9057 34043 9069
rect 34314 9085 34363 9095
rect 34314 9065 34325 9085
rect 34345 9065 34363 9085
rect 34314 9053 34363 9065
rect 34413 9089 34457 9095
rect 34413 9069 34428 9089
rect 34448 9069 34457 9089
rect 34413 9053 34457 9069
rect 34527 9085 34576 9095
rect 34527 9065 34538 9085
rect 34558 9065 34576 9085
rect 34527 9053 34576 9065
rect 34626 9089 34670 9095
rect 34626 9069 34641 9089
rect 34661 9069 34670 9089
rect 34626 9053 34670 9069
rect 34735 9085 34784 9095
rect 34735 9065 34746 9085
rect 34766 9065 34784 9085
rect 34735 9053 34784 9065
rect 34834 9089 34878 9095
rect 34834 9069 34849 9089
rect 34869 9069 34878 9089
rect 34834 9053 34878 9069
rect 34948 9089 34992 9095
rect 34948 9069 34957 9089
rect 34977 9069 34992 9089
rect 34948 9053 34992 9069
rect 35042 9085 35091 9095
rect 35042 9065 35060 9085
rect 35080 9065 35091 9085
rect 35042 9053 35091 9065
rect 8127 8549 8176 8561
rect 8127 8529 8138 8549
rect 8158 8529 8176 8549
rect 8127 8519 8176 8529
rect 8226 8545 8270 8561
rect 8226 8525 8241 8545
rect 8261 8525 8270 8545
rect 8226 8519 8270 8525
rect 8340 8545 8384 8561
rect 8340 8525 8349 8545
rect 8369 8525 8384 8545
rect 8340 8519 8384 8525
rect 8434 8549 8483 8561
rect 8434 8529 8452 8549
rect 8472 8529 8483 8549
rect 8434 8519 8483 8529
rect 8548 8545 8592 8561
rect 8548 8525 8557 8545
rect 8577 8525 8592 8545
rect 8548 8519 8592 8525
rect 8642 8549 8691 8561
rect 8642 8529 8660 8549
rect 8680 8529 8691 8549
rect 8642 8519 8691 8529
rect 8761 8545 8805 8561
rect 8761 8525 8770 8545
rect 8790 8525 8805 8545
rect 8761 8519 8805 8525
rect 8855 8549 8904 8561
rect 8855 8529 8873 8549
rect 8893 8529 8904 8549
rect 8855 8519 8904 8529
rect 9175 8545 9224 8557
rect 9175 8525 9186 8545
rect 9206 8525 9224 8545
rect 885 8418 934 8428
rect 885 8398 896 8418
rect 916 8398 934 8418
rect 885 8386 934 8398
rect 984 8422 1028 8428
rect 984 8402 999 8422
rect 1019 8402 1028 8422
rect 984 8386 1028 8402
rect 1098 8418 1147 8428
rect 1098 8398 1109 8418
rect 1129 8398 1147 8418
rect 1098 8386 1147 8398
rect 1197 8422 1241 8428
rect 1197 8402 1212 8422
rect 1232 8402 1241 8422
rect 1197 8386 1241 8402
rect 1306 8418 1355 8428
rect 1306 8398 1317 8418
rect 1337 8398 1355 8418
rect 1306 8386 1355 8398
rect 1405 8422 1449 8428
rect 1405 8402 1420 8422
rect 1440 8402 1449 8422
rect 1405 8386 1449 8402
rect 1519 8422 1563 8428
rect 1519 8402 1528 8422
rect 1548 8402 1563 8422
rect 1519 8386 1563 8402
rect 1613 8418 1662 8428
rect 9175 8515 9224 8525
rect 9274 8541 9318 8557
rect 9274 8521 9289 8541
rect 9309 8521 9318 8541
rect 9274 8515 9318 8521
rect 9388 8541 9432 8557
rect 9388 8521 9397 8541
rect 9417 8521 9432 8541
rect 9388 8515 9432 8521
rect 9482 8545 9531 8557
rect 9482 8525 9500 8545
rect 9520 8525 9531 8545
rect 9482 8515 9531 8525
rect 9596 8541 9640 8557
rect 9596 8521 9605 8541
rect 9625 8521 9640 8541
rect 9596 8515 9640 8521
rect 9690 8545 9739 8557
rect 9690 8525 9708 8545
rect 9728 8525 9739 8545
rect 9690 8515 9739 8525
rect 9809 8541 9853 8557
rect 9809 8521 9818 8541
rect 9838 8521 9853 8541
rect 9809 8515 9853 8521
rect 9903 8545 9952 8557
rect 9903 8525 9921 8545
rect 9941 8525 9952 8545
rect 9903 8515 9952 8525
rect 1613 8398 1631 8418
rect 1651 8398 1662 8418
rect 1613 8386 1662 8398
rect 4488 8409 4537 8419
rect 4488 8389 4499 8409
rect 4519 8389 4537 8409
rect 4488 8377 4537 8389
rect 4587 8413 4631 8419
rect 4587 8393 4602 8413
rect 4622 8393 4631 8413
rect 4587 8377 4631 8393
rect 4701 8409 4750 8419
rect 4701 8389 4712 8409
rect 4732 8389 4750 8409
rect 4701 8377 4750 8389
rect 4800 8413 4844 8419
rect 4800 8393 4815 8413
rect 4835 8393 4844 8413
rect 4800 8377 4844 8393
rect 4909 8409 4958 8419
rect 4909 8389 4920 8409
rect 4940 8389 4958 8409
rect 4909 8377 4958 8389
rect 5008 8413 5052 8419
rect 5008 8393 5023 8413
rect 5043 8393 5052 8413
rect 5008 8377 5052 8393
rect 5122 8413 5166 8419
rect 5122 8393 5131 8413
rect 5151 8393 5166 8413
rect 5122 8377 5166 8393
rect 5216 8409 5265 8419
rect 5216 8389 5234 8409
rect 5254 8389 5265 8409
rect 5216 8377 5265 8389
rect 18835 8543 18884 8555
rect 18835 8523 18846 8543
rect 18866 8523 18884 8543
rect 18835 8513 18884 8523
rect 18934 8539 18978 8555
rect 18934 8519 18949 8539
rect 18969 8519 18978 8539
rect 18934 8513 18978 8519
rect 19048 8539 19092 8555
rect 19048 8519 19057 8539
rect 19077 8519 19092 8539
rect 19048 8513 19092 8519
rect 19142 8543 19191 8555
rect 19142 8523 19160 8543
rect 19180 8523 19191 8543
rect 19142 8513 19191 8523
rect 19256 8539 19300 8555
rect 19256 8519 19265 8539
rect 19285 8519 19300 8539
rect 19256 8513 19300 8519
rect 19350 8543 19399 8555
rect 19350 8523 19368 8543
rect 19388 8523 19399 8543
rect 19350 8513 19399 8523
rect 19469 8539 19513 8555
rect 19469 8519 19478 8539
rect 19498 8519 19513 8539
rect 19469 8513 19513 8519
rect 19563 8543 19612 8555
rect 19563 8523 19581 8543
rect 19601 8523 19612 8543
rect 19563 8513 19612 8523
rect 19883 8539 19932 8551
rect 19883 8519 19894 8539
rect 19914 8519 19932 8539
rect 11593 8412 11642 8422
rect 11593 8392 11604 8412
rect 11624 8392 11642 8412
rect 11593 8380 11642 8392
rect 11692 8416 11736 8422
rect 11692 8396 11707 8416
rect 11727 8396 11736 8416
rect 11692 8380 11736 8396
rect 11806 8412 11855 8422
rect 11806 8392 11817 8412
rect 11837 8392 11855 8412
rect 11806 8380 11855 8392
rect 11905 8416 11949 8422
rect 11905 8396 11920 8416
rect 11940 8396 11949 8416
rect 11905 8380 11949 8396
rect 12014 8412 12063 8422
rect 12014 8392 12025 8412
rect 12045 8392 12063 8412
rect 12014 8380 12063 8392
rect 12113 8416 12157 8422
rect 12113 8396 12128 8416
rect 12148 8396 12157 8416
rect 12113 8380 12157 8396
rect 12227 8416 12271 8422
rect 12227 8396 12236 8416
rect 12256 8396 12271 8416
rect 12227 8380 12271 8396
rect 12321 8412 12370 8422
rect 19883 8509 19932 8519
rect 19982 8535 20026 8551
rect 19982 8515 19997 8535
rect 20017 8515 20026 8535
rect 19982 8509 20026 8515
rect 20096 8535 20140 8551
rect 20096 8515 20105 8535
rect 20125 8515 20140 8535
rect 20096 8509 20140 8515
rect 20190 8539 20239 8551
rect 20190 8519 20208 8539
rect 20228 8519 20239 8539
rect 20190 8509 20239 8519
rect 20304 8535 20348 8551
rect 20304 8515 20313 8535
rect 20333 8515 20348 8535
rect 20304 8509 20348 8515
rect 20398 8539 20447 8551
rect 20398 8519 20416 8539
rect 20436 8519 20447 8539
rect 20398 8509 20447 8519
rect 20517 8535 20561 8551
rect 20517 8515 20526 8535
rect 20546 8515 20561 8535
rect 20517 8509 20561 8515
rect 20611 8539 20660 8551
rect 20611 8519 20629 8539
rect 20649 8519 20660 8539
rect 20611 8509 20660 8519
rect 12321 8392 12339 8412
rect 12359 8392 12370 8412
rect 12321 8380 12370 8392
rect 15196 8403 15245 8413
rect 15196 8383 15207 8403
rect 15227 8383 15245 8403
rect 15196 8371 15245 8383
rect 15295 8407 15339 8413
rect 15295 8387 15310 8407
rect 15330 8387 15339 8407
rect 15295 8371 15339 8387
rect 15409 8403 15458 8413
rect 15409 8383 15420 8403
rect 15440 8383 15458 8403
rect 15409 8371 15458 8383
rect 15508 8407 15552 8413
rect 15508 8387 15523 8407
rect 15543 8387 15552 8407
rect 15508 8371 15552 8387
rect 15617 8403 15666 8413
rect 15617 8383 15628 8403
rect 15648 8383 15666 8403
rect 15617 8371 15666 8383
rect 15716 8407 15760 8413
rect 15716 8387 15731 8407
rect 15751 8387 15760 8407
rect 15716 8371 15760 8387
rect 15830 8407 15874 8413
rect 15830 8387 15839 8407
rect 15859 8387 15874 8407
rect 15830 8371 15874 8387
rect 15924 8403 15973 8413
rect 15924 8383 15942 8403
rect 15962 8383 15973 8403
rect 15924 8371 15973 8383
rect 29800 8547 29849 8559
rect 29800 8527 29811 8547
rect 29831 8527 29849 8547
rect 29800 8517 29849 8527
rect 29899 8543 29943 8559
rect 29899 8523 29914 8543
rect 29934 8523 29943 8543
rect 29899 8517 29943 8523
rect 30013 8543 30057 8559
rect 30013 8523 30022 8543
rect 30042 8523 30057 8543
rect 30013 8517 30057 8523
rect 30107 8547 30156 8559
rect 30107 8527 30125 8547
rect 30145 8527 30156 8547
rect 30107 8517 30156 8527
rect 30221 8543 30265 8559
rect 30221 8523 30230 8543
rect 30250 8523 30265 8543
rect 30221 8517 30265 8523
rect 30315 8547 30364 8559
rect 30315 8527 30333 8547
rect 30353 8527 30364 8547
rect 30315 8517 30364 8527
rect 30434 8543 30478 8559
rect 30434 8523 30443 8543
rect 30463 8523 30478 8543
rect 30434 8517 30478 8523
rect 30528 8547 30577 8559
rect 30528 8527 30546 8547
rect 30566 8527 30577 8547
rect 30528 8517 30577 8527
rect 30848 8543 30897 8555
rect 30848 8523 30859 8543
rect 30879 8523 30897 8543
rect 22558 8416 22607 8426
rect 22558 8396 22569 8416
rect 22589 8396 22607 8416
rect 22558 8384 22607 8396
rect 22657 8420 22701 8426
rect 22657 8400 22672 8420
rect 22692 8400 22701 8420
rect 22657 8384 22701 8400
rect 22771 8416 22820 8426
rect 22771 8396 22782 8416
rect 22802 8396 22820 8416
rect 22771 8384 22820 8396
rect 22870 8420 22914 8426
rect 22870 8400 22885 8420
rect 22905 8400 22914 8420
rect 22870 8384 22914 8400
rect 22979 8416 23028 8426
rect 22979 8396 22990 8416
rect 23010 8396 23028 8416
rect 22979 8384 23028 8396
rect 23078 8420 23122 8426
rect 23078 8400 23093 8420
rect 23113 8400 23122 8420
rect 23078 8384 23122 8400
rect 23192 8420 23236 8426
rect 23192 8400 23201 8420
rect 23221 8400 23236 8420
rect 23192 8384 23236 8400
rect 23286 8416 23335 8426
rect 30848 8513 30897 8523
rect 30947 8539 30991 8555
rect 30947 8519 30962 8539
rect 30982 8519 30991 8539
rect 30947 8513 30991 8519
rect 31061 8539 31105 8555
rect 31061 8519 31070 8539
rect 31090 8519 31105 8539
rect 31061 8513 31105 8519
rect 31155 8543 31204 8555
rect 31155 8523 31173 8543
rect 31193 8523 31204 8543
rect 31155 8513 31204 8523
rect 31269 8539 31313 8555
rect 31269 8519 31278 8539
rect 31298 8519 31313 8539
rect 31269 8513 31313 8519
rect 31363 8543 31412 8555
rect 31363 8523 31381 8543
rect 31401 8523 31412 8543
rect 31363 8513 31412 8523
rect 31482 8539 31526 8555
rect 31482 8519 31491 8539
rect 31511 8519 31526 8539
rect 31482 8513 31526 8519
rect 31576 8543 31625 8555
rect 31576 8523 31594 8543
rect 31614 8523 31625 8543
rect 31576 8513 31625 8523
rect 23286 8396 23304 8416
rect 23324 8396 23335 8416
rect 23286 8384 23335 8396
rect 26161 8407 26210 8417
rect 26161 8387 26172 8407
rect 26192 8387 26210 8407
rect 26161 8375 26210 8387
rect 26260 8411 26304 8417
rect 26260 8391 26275 8411
rect 26295 8391 26304 8411
rect 26260 8375 26304 8391
rect 26374 8407 26423 8417
rect 26374 8387 26385 8407
rect 26405 8387 26423 8407
rect 26374 8375 26423 8387
rect 26473 8411 26517 8417
rect 26473 8391 26488 8411
rect 26508 8391 26517 8411
rect 26473 8375 26517 8391
rect 26582 8407 26631 8417
rect 26582 8387 26593 8407
rect 26613 8387 26631 8407
rect 26582 8375 26631 8387
rect 26681 8411 26725 8417
rect 26681 8391 26696 8411
rect 26716 8391 26725 8411
rect 26681 8375 26725 8391
rect 26795 8411 26839 8417
rect 26795 8391 26804 8411
rect 26824 8391 26839 8411
rect 26795 8375 26839 8391
rect 26889 8407 26938 8417
rect 26889 8387 26907 8407
rect 26927 8387 26938 8407
rect 26889 8375 26938 8387
rect 40508 8541 40557 8553
rect 40508 8521 40519 8541
rect 40539 8521 40557 8541
rect 40508 8511 40557 8521
rect 40607 8537 40651 8553
rect 40607 8517 40622 8537
rect 40642 8517 40651 8537
rect 40607 8511 40651 8517
rect 40721 8537 40765 8553
rect 40721 8517 40730 8537
rect 40750 8517 40765 8537
rect 40721 8511 40765 8517
rect 40815 8541 40864 8553
rect 40815 8521 40833 8541
rect 40853 8521 40864 8541
rect 40815 8511 40864 8521
rect 40929 8537 40973 8553
rect 40929 8517 40938 8537
rect 40958 8517 40973 8537
rect 40929 8511 40973 8517
rect 41023 8541 41072 8553
rect 41023 8521 41041 8541
rect 41061 8521 41072 8541
rect 41023 8511 41072 8521
rect 41142 8537 41186 8553
rect 41142 8517 41151 8537
rect 41171 8517 41186 8537
rect 41142 8511 41186 8517
rect 41236 8541 41285 8553
rect 41236 8521 41254 8541
rect 41274 8521 41285 8541
rect 41236 8511 41285 8521
rect 41556 8537 41605 8549
rect 41556 8517 41567 8537
rect 41587 8517 41605 8537
rect 33266 8410 33315 8420
rect 33266 8390 33277 8410
rect 33297 8390 33315 8410
rect 33266 8378 33315 8390
rect 33365 8414 33409 8420
rect 33365 8394 33380 8414
rect 33400 8394 33409 8414
rect 33365 8378 33409 8394
rect 33479 8410 33528 8420
rect 33479 8390 33490 8410
rect 33510 8390 33528 8410
rect 33479 8378 33528 8390
rect 33578 8414 33622 8420
rect 33578 8394 33593 8414
rect 33613 8394 33622 8414
rect 33578 8378 33622 8394
rect 33687 8410 33736 8420
rect 33687 8390 33698 8410
rect 33718 8390 33736 8410
rect 33687 8378 33736 8390
rect 33786 8414 33830 8420
rect 33786 8394 33801 8414
rect 33821 8394 33830 8414
rect 33786 8378 33830 8394
rect 33900 8414 33944 8420
rect 33900 8394 33909 8414
rect 33929 8394 33944 8414
rect 33900 8378 33944 8394
rect 33994 8410 34043 8420
rect 41556 8507 41605 8517
rect 41655 8533 41699 8549
rect 41655 8513 41670 8533
rect 41690 8513 41699 8533
rect 41655 8507 41699 8513
rect 41769 8533 41813 8549
rect 41769 8513 41778 8533
rect 41798 8513 41813 8533
rect 41769 8507 41813 8513
rect 41863 8537 41912 8549
rect 41863 8517 41881 8537
rect 41901 8517 41912 8537
rect 41863 8507 41912 8517
rect 41977 8533 42021 8549
rect 41977 8513 41986 8533
rect 42006 8513 42021 8533
rect 41977 8507 42021 8513
rect 42071 8537 42120 8549
rect 42071 8517 42089 8537
rect 42109 8517 42120 8537
rect 42071 8507 42120 8517
rect 42190 8533 42234 8549
rect 42190 8513 42199 8533
rect 42219 8513 42234 8533
rect 42190 8507 42234 8513
rect 42284 8537 42333 8549
rect 42284 8517 42302 8537
rect 42322 8517 42333 8537
rect 42284 8507 42333 8517
rect 33994 8390 34012 8410
rect 34032 8390 34043 8410
rect 33994 8378 34043 8390
rect 36869 8401 36918 8411
rect 36869 8381 36880 8401
rect 36900 8381 36918 8401
rect 36869 8369 36918 8381
rect 36968 8405 37012 8411
rect 36968 8385 36983 8405
rect 37003 8385 37012 8405
rect 36968 8369 37012 8385
rect 37082 8401 37131 8411
rect 37082 8381 37093 8401
rect 37113 8381 37131 8401
rect 37082 8369 37131 8381
rect 37181 8405 37225 8411
rect 37181 8385 37196 8405
rect 37216 8385 37225 8405
rect 37181 8369 37225 8385
rect 37290 8401 37339 8411
rect 37290 8381 37301 8401
rect 37321 8381 37339 8401
rect 37290 8369 37339 8381
rect 37389 8405 37433 8411
rect 37389 8385 37404 8405
rect 37424 8385 37433 8405
rect 37389 8369 37433 8385
rect 37503 8405 37547 8411
rect 37503 8385 37512 8405
rect 37532 8385 37547 8405
rect 37503 8369 37547 8385
rect 37597 8401 37646 8411
rect 37597 8381 37615 8401
rect 37635 8381 37646 8401
rect 37597 8369 37646 8381
rect 5569 7639 5618 7651
rect 5569 7619 5580 7639
rect 5600 7619 5618 7639
rect 5569 7609 5618 7619
rect 5668 7635 5712 7651
rect 5668 7615 5683 7635
rect 5703 7615 5712 7635
rect 5668 7609 5712 7615
rect 5782 7635 5826 7651
rect 5782 7615 5791 7635
rect 5811 7615 5826 7635
rect 5782 7609 5826 7615
rect 5876 7639 5925 7651
rect 5876 7619 5894 7639
rect 5914 7619 5925 7639
rect 5876 7609 5925 7619
rect 5990 7635 6034 7651
rect 5990 7615 5999 7635
rect 6019 7615 6034 7635
rect 5990 7609 6034 7615
rect 6084 7639 6133 7651
rect 6084 7619 6102 7639
rect 6122 7619 6133 7639
rect 6084 7609 6133 7619
rect 6203 7635 6247 7651
rect 6203 7615 6212 7635
rect 6232 7615 6247 7635
rect 6203 7609 6247 7615
rect 6297 7639 6346 7651
rect 6297 7619 6315 7639
rect 6335 7619 6346 7639
rect 6297 7609 6346 7619
rect 9172 7630 9221 7642
rect 9172 7610 9183 7630
rect 9203 7610 9221 7630
rect 882 7503 931 7513
rect 882 7483 893 7503
rect 913 7483 931 7503
rect 882 7471 931 7483
rect 981 7507 1025 7513
rect 981 7487 996 7507
rect 1016 7487 1025 7507
rect 981 7471 1025 7487
rect 1095 7503 1144 7513
rect 1095 7483 1106 7503
rect 1126 7483 1144 7503
rect 1095 7471 1144 7483
rect 1194 7507 1238 7513
rect 1194 7487 1209 7507
rect 1229 7487 1238 7507
rect 1194 7471 1238 7487
rect 1303 7503 1352 7513
rect 1303 7483 1314 7503
rect 1334 7483 1352 7503
rect 1303 7471 1352 7483
rect 1402 7507 1446 7513
rect 1402 7487 1417 7507
rect 1437 7487 1446 7507
rect 1402 7471 1446 7487
rect 1516 7507 1560 7513
rect 1516 7487 1525 7507
rect 1545 7487 1560 7507
rect 1516 7471 1560 7487
rect 1610 7503 1659 7513
rect 9172 7600 9221 7610
rect 9271 7626 9315 7642
rect 9271 7606 9286 7626
rect 9306 7606 9315 7626
rect 9271 7600 9315 7606
rect 9385 7626 9429 7642
rect 9385 7606 9394 7626
rect 9414 7606 9429 7626
rect 9385 7600 9429 7606
rect 9479 7630 9528 7642
rect 9479 7610 9497 7630
rect 9517 7610 9528 7630
rect 9479 7600 9528 7610
rect 9593 7626 9637 7642
rect 9593 7606 9602 7626
rect 9622 7606 9637 7626
rect 9593 7600 9637 7606
rect 9687 7630 9736 7642
rect 9687 7610 9705 7630
rect 9725 7610 9736 7630
rect 9687 7600 9736 7610
rect 9806 7626 9850 7642
rect 9806 7606 9815 7626
rect 9835 7606 9850 7626
rect 9806 7600 9850 7606
rect 9900 7630 9949 7642
rect 9900 7610 9918 7630
rect 9938 7610 9949 7630
rect 9900 7600 9949 7610
rect 1610 7483 1628 7503
rect 1648 7483 1659 7503
rect 1610 7471 1659 7483
rect 1930 7499 1979 7509
rect 1930 7479 1941 7499
rect 1961 7479 1979 7499
rect 1930 7467 1979 7479
rect 2029 7503 2073 7509
rect 2029 7483 2044 7503
rect 2064 7483 2073 7503
rect 2029 7467 2073 7483
rect 2143 7499 2192 7509
rect 2143 7479 2154 7499
rect 2174 7479 2192 7499
rect 2143 7467 2192 7479
rect 2242 7503 2286 7509
rect 2242 7483 2257 7503
rect 2277 7483 2286 7503
rect 2242 7467 2286 7483
rect 2351 7499 2400 7509
rect 2351 7479 2362 7499
rect 2382 7479 2400 7499
rect 2351 7467 2400 7479
rect 2450 7503 2494 7509
rect 2450 7483 2465 7503
rect 2485 7483 2494 7503
rect 2450 7467 2494 7483
rect 2564 7503 2608 7509
rect 2564 7483 2573 7503
rect 2593 7483 2608 7503
rect 2564 7467 2608 7483
rect 2658 7499 2707 7509
rect 2658 7479 2676 7499
rect 2696 7479 2707 7499
rect 2658 7467 2707 7479
rect 16277 7633 16326 7645
rect 16277 7613 16288 7633
rect 16308 7613 16326 7633
rect 16277 7603 16326 7613
rect 16376 7629 16420 7645
rect 16376 7609 16391 7629
rect 16411 7609 16420 7629
rect 16376 7603 16420 7609
rect 16490 7629 16534 7645
rect 16490 7609 16499 7629
rect 16519 7609 16534 7629
rect 16490 7603 16534 7609
rect 16584 7633 16633 7645
rect 16584 7613 16602 7633
rect 16622 7613 16633 7633
rect 16584 7603 16633 7613
rect 16698 7629 16742 7645
rect 16698 7609 16707 7629
rect 16727 7609 16742 7629
rect 16698 7603 16742 7609
rect 16792 7633 16841 7645
rect 16792 7613 16810 7633
rect 16830 7613 16841 7633
rect 16792 7603 16841 7613
rect 16911 7629 16955 7645
rect 16911 7609 16920 7629
rect 16940 7609 16955 7629
rect 16911 7603 16955 7609
rect 17005 7633 17054 7645
rect 17005 7613 17023 7633
rect 17043 7613 17054 7633
rect 17005 7603 17054 7613
rect 19880 7624 19929 7636
rect 19880 7604 19891 7624
rect 19911 7604 19929 7624
rect 11590 7497 11639 7507
rect 11590 7477 11601 7497
rect 11621 7477 11639 7497
rect 11590 7465 11639 7477
rect 11689 7501 11733 7507
rect 11689 7481 11704 7501
rect 11724 7481 11733 7501
rect 11689 7465 11733 7481
rect 11803 7497 11852 7507
rect 11803 7477 11814 7497
rect 11834 7477 11852 7497
rect 11803 7465 11852 7477
rect 11902 7501 11946 7507
rect 11902 7481 11917 7501
rect 11937 7481 11946 7501
rect 11902 7465 11946 7481
rect 12011 7497 12060 7507
rect 12011 7477 12022 7497
rect 12042 7477 12060 7497
rect 12011 7465 12060 7477
rect 12110 7501 12154 7507
rect 12110 7481 12125 7501
rect 12145 7481 12154 7501
rect 12110 7465 12154 7481
rect 12224 7501 12268 7507
rect 12224 7481 12233 7501
rect 12253 7481 12268 7501
rect 12224 7465 12268 7481
rect 12318 7497 12367 7507
rect 19880 7594 19929 7604
rect 19979 7620 20023 7636
rect 19979 7600 19994 7620
rect 20014 7600 20023 7620
rect 19979 7594 20023 7600
rect 20093 7620 20137 7636
rect 20093 7600 20102 7620
rect 20122 7600 20137 7620
rect 20093 7594 20137 7600
rect 20187 7624 20236 7636
rect 20187 7604 20205 7624
rect 20225 7604 20236 7624
rect 20187 7594 20236 7604
rect 20301 7620 20345 7636
rect 20301 7600 20310 7620
rect 20330 7600 20345 7620
rect 20301 7594 20345 7600
rect 20395 7624 20444 7636
rect 20395 7604 20413 7624
rect 20433 7604 20444 7624
rect 20395 7594 20444 7604
rect 20514 7620 20558 7636
rect 20514 7600 20523 7620
rect 20543 7600 20558 7620
rect 20514 7594 20558 7600
rect 20608 7624 20657 7636
rect 20608 7604 20626 7624
rect 20646 7604 20657 7624
rect 20608 7594 20657 7604
rect 12318 7477 12336 7497
rect 12356 7477 12367 7497
rect 12318 7465 12367 7477
rect 12638 7493 12687 7503
rect 12638 7473 12649 7493
rect 12669 7473 12687 7493
rect 12638 7461 12687 7473
rect 12737 7497 12781 7503
rect 12737 7477 12752 7497
rect 12772 7477 12781 7497
rect 12737 7461 12781 7477
rect 12851 7493 12900 7503
rect 12851 7473 12862 7493
rect 12882 7473 12900 7493
rect 12851 7461 12900 7473
rect 12950 7497 12994 7503
rect 12950 7477 12965 7497
rect 12985 7477 12994 7497
rect 12950 7461 12994 7477
rect 13059 7493 13108 7503
rect 13059 7473 13070 7493
rect 13090 7473 13108 7493
rect 13059 7461 13108 7473
rect 13158 7497 13202 7503
rect 13158 7477 13173 7497
rect 13193 7477 13202 7497
rect 13158 7461 13202 7477
rect 13272 7497 13316 7503
rect 13272 7477 13281 7497
rect 13301 7477 13316 7497
rect 13272 7461 13316 7477
rect 13366 7493 13415 7503
rect 13366 7473 13384 7493
rect 13404 7473 13415 7493
rect 13366 7461 13415 7473
rect 27242 7637 27291 7649
rect 27242 7617 27253 7637
rect 27273 7617 27291 7637
rect 27242 7607 27291 7617
rect 27341 7633 27385 7649
rect 27341 7613 27356 7633
rect 27376 7613 27385 7633
rect 27341 7607 27385 7613
rect 27455 7633 27499 7649
rect 27455 7613 27464 7633
rect 27484 7613 27499 7633
rect 27455 7607 27499 7613
rect 27549 7637 27598 7649
rect 27549 7617 27567 7637
rect 27587 7617 27598 7637
rect 27549 7607 27598 7617
rect 27663 7633 27707 7649
rect 27663 7613 27672 7633
rect 27692 7613 27707 7633
rect 27663 7607 27707 7613
rect 27757 7637 27806 7649
rect 27757 7617 27775 7637
rect 27795 7617 27806 7637
rect 27757 7607 27806 7617
rect 27876 7633 27920 7649
rect 27876 7613 27885 7633
rect 27905 7613 27920 7633
rect 27876 7607 27920 7613
rect 27970 7637 28019 7649
rect 27970 7617 27988 7637
rect 28008 7617 28019 7637
rect 27970 7607 28019 7617
rect 30845 7628 30894 7640
rect 30845 7608 30856 7628
rect 30876 7608 30894 7628
rect 22555 7501 22604 7511
rect 22555 7481 22566 7501
rect 22586 7481 22604 7501
rect 22555 7469 22604 7481
rect 22654 7505 22698 7511
rect 22654 7485 22669 7505
rect 22689 7485 22698 7505
rect 22654 7469 22698 7485
rect 22768 7501 22817 7511
rect 22768 7481 22779 7501
rect 22799 7481 22817 7501
rect 22768 7469 22817 7481
rect 22867 7505 22911 7511
rect 22867 7485 22882 7505
rect 22902 7485 22911 7505
rect 22867 7469 22911 7485
rect 22976 7501 23025 7511
rect 22976 7481 22987 7501
rect 23007 7481 23025 7501
rect 22976 7469 23025 7481
rect 23075 7505 23119 7511
rect 23075 7485 23090 7505
rect 23110 7485 23119 7505
rect 23075 7469 23119 7485
rect 23189 7505 23233 7511
rect 23189 7485 23198 7505
rect 23218 7485 23233 7505
rect 23189 7469 23233 7485
rect 23283 7501 23332 7511
rect 30845 7598 30894 7608
rect 30944 7624 30988 7640
rect 30944 7604 30959 7624
rect 30979 7604 30988 7624
rect 30944 7598 30988 7604
rect 31058 7624 31102 7640
rect 31058 7604 31067 7624
rect 31087 7604 31102 7624
rect 31058 7598 31102 7604
rect 31152 7628 31201 7640
rect 31152 7608 31170 7628
rect 31190 7608 31201 7628
rect 31152 7598 31201 7608
rect 31266 7624 31310 7640
rect 31266 7604 31275 7624
rect 31295 7604 31310 7624
rect 31266 7598 31310 7604
rect 31360 7628 31409 7640
rect 31360 7608 31378 7628
rect 31398 7608 31409 7628
rect 31360 7598 31409 7608
rect 31479 7624 31523 7640
rect 31479 7604 31488 7624
rect 31508 7604 31523 7624
rect 31479 7598 31523 7604
rect 31573 7628 31622 7640
rect 31573 7608 31591 7628
rect 31611 7608 31622 7628
rect 31573 7598 31622 7608
rect 23283 7481 23301 7501
rect 23321 7481 23332 7501
rect 23283 7469 23332 7481
rect 23603 7497 23652 7507
rect 23603 7477 23614 7497
rect 23634 7477 23652 7497
rect 23603 7465 23652 7477
rect 23702 7501 23746 7507
rect 23702 7481 23717 7501
rect 23737 7481 23746 7501
rect 23702 7465 23746 7481
rect 23816 7497 23865 7507
rect 23816 7477 23827 7497
rect 23847 7477 23865 7497
rect 23816 7465 23865 7477
rect 23915 7501 23959 7507
rect 23915 7481 23930 7501
rect 23950 7481 23959 7501
rect 23915 7465 23959 7481
rect 24024 7497 24073 7507
rect 24024 7477 24035 7497
rect 24055 7477 24073 7497
rect 24024 7465 24073 7477
rect 24123 7501 24167 7507
rect 24123 7481 24138 7501
rect 24158 7481 24167 7501
rect 24123 7465 24167 7481
rect 24237 7501 24281 7507
rect 24237 7481 24246 7501
rect 24266 7481 24281 7501
rect 24237 7465 24281 7481
rect 24331 7497 24380 7507
rect 24331 7477 24349 7497
rect 24369 7477 24380 7497
rect 24331 7465 24380 7477
rect 37950 7631 37999 7643
rect 37950 7611 37961 7631
rect 37981 7611 37999 7631
rect 37950 7601 37999 7611
rect 38049 7627 38093 7643
rect 38049 7607 38064 7627
rect 38084 7607 38093 7627
rect 38049 7601 38093 7607
rect 38163 7627 38207 7643
rect 38163 7607 38172 7627
rect 38192 7607 38207 7627
rect 38163 7601 38207 7607
rect 38257 7631 38306 7643
rect 38257 7611 38275 7631
rect 38295 7611 38306 7631
rect 38257 7601 38306 7611
rect 38371 7627 38415 7643
rect 38371 7607 38380 7627
rect 38400 7607 38415 7627
rect 38371 7601 38415 7607
rect 38465 7631 38514 7643
rect 38465 7611 38483 7631
rect 38503 7611 38514 7631
rect 38465 7601 38514 7611
rect 38584 7627 38628 7643
rect 38584 7607 38593 7627
rect 38613 7607 38628 7627
rect 38584 7601 38628 7607
rect 38678 7631 38727 7643
rect 38678 7611 38696 7631
rect 38716 7611 38727 7631
rect 38678 7601 38727 7611
rect 41553 7622 41602 7634
rect 41553 7602 41564 7622
rect 41584 7602 41602 7622
rect 33263 7495 33312 7505
rect 33263 7475 33274 7495
rect 33294 7475 33312 7495
rect 33263 7463 33312 7475
rect 33362 7499 33406 7505
rect 33362 7479 33377 7499
rect 33397 7479 33406 7499
rect 33362 7463 33406 7479
rect 33476 7495 33525 7505
rect 33476 7475 33487 7495
rect 33507 7475 33525 7495
rect 33476 7463 33525 7475
rect 33575 7499 33619 7505
rect 33575 7479 33590 7499
rect 33610 7479 33619 7499
rect 33575 7463 33619 7479
rect 33684 7495 33733 7505
rect 33684 7475 33695 7495
rect 33715 7475 33733 7495
rect 33684 7463 33733 7475
rect 33783 7499 33827 7505
rect 33783 7479 33798 7499
rect 33818 7479 33827 7499
rect 33783 7463 33827 7479
rect 33897 7499 33941 7505
rect 33897 7479 33906 7499
rect 33926 7479 33941 7499
rect 33897 7463 33941 7479
rect 33991 7495 34040 7505
rect 41553 7592 41602 7602
rect 41652 7618 41696 7634
rect 41652 7598 41667 7618
rect 41687 7598 41696 7618
rect 41652 7592 41696 7598
rect 41766 7618 41810 7634
rect 41766 7598 41775 7618
rect 41795 7598 41810 7618
rect 41766 7592 41810 7598
rect 41860 7622 41909 7634
rect 41860 7602 41878 7622
rect 41898 7602 41909 7622
rect 41860 7592 41909 7602
rect 41974 7618 42018 7634
rect 41974 7598 41983 7618
rect 42003 7598 42018 7618
rect 41974 7592 42018 7598
rect 42068 7622 42117 7634
rect 42068 7602 42086 7622
rect 42106 7602 42117 7622
rect 42068 7592 42117 7602
rect 42187 7618 42231 7634
rect 42187 7598 42196 7618
rect 42216 7598 42231 7618
rect 42187 7592 42231 7598
rect 42281 7622 42330 7634
rect 42281 7602 42299 7622
rect 42319 7602 42330 7622
rect 42281 7592 42330 7602
rect 33991 7475 34009 7495
rect 34029 7475 34040 7495
rect 33991 7463 34040 7475
rect 34311 7491 34360 7501
rect 34311 7471 34322 7491
rect 34342 7471 34360 7491
rect 34311 7459 34360 7471
rect 34410 7495 34454 7501
rect 34410 7475 34425 7495
rect 34445 7475 34454 7495
rect 34410 7459 34454 7475
rect 34524 7491 34573 7501
rect 34524 7471 34535 7491
rect 34555 7471 34573 7491
rect 34524 7459 34573 7471
rect 34623 7495 34667 7501
rect 34623 7475 34638 7495
rect 34658 7475 34667 7495
rect 34623 7459 34667 7475
rect 34732 7491 34781 7501
rect 34732 7471 34743 7491
rect 34763 7471 34781 7491
rect 34732 7459 34781 7471
rect 34831 7495 34875 7501
rect 34831 7475 34846 7495
rect 34866 7475 34875 7495
rect 34831 7459 34875 7475
rect 34945 7495 34989 7501
rect 34945 7475 34954 7495
rect 34974 7475 34989 7495
rect 34945 7459 34989 7475
rect 35039 7491 35088 7501
rect 35039 7471 35057 7491
rect 35077 7471 35088 7491
rect 35039 7459 35088 7471
rect 8124 6955 8173 6967
rect 8124 6935 8135 6955
rect 8155 6935 8173 6955
rect 8124 6925 8173 6935
rect 8223 6951 8267 6967
rect 8223 6931 8238 6951
rect 8258 6931 8267 6951
rect 8223 6925 8267 6931
rect 8337 6951 8381 6967
rect 8337 6931 8346 6951
rect 8366 6931 8381 6951
rect 8337 6925 8381 6931
rect 8431 6955 8480 6967
rect 8431 6935 8449 6955
rect 8469 6935 8480 6955
rect 8431 6925 8480 6935
rect 8545 6951 8589 6967
rect 8545 6931 8554 6951
rect 8574 6931 8589 6951
rect 8545 6925 8589 6931
rect 8639 6955 8688 6967
rect 8639 6935 8657 6955
rect 8677 6935 8688 6955
rect 8639 6925 8688 6935
rect 8758 6951 8802 6967
rect 8758 6931 8767 6951
rect 8787 6931 8802 6951
rect 8758 6925 8802 6931
rect 8852 6955 8901 6967
rect 8852 6935 8870 6955
rect 8890 6935 8901 6955
rect 8852 6925 8901 6935
rect 9172 6951 9221 6963
rect 9172 6931 9183 6951
rect 9203 6931 9221 6951
rect 882 6824 931 6834
rect 882 6804 893 6824
rect 913 6804 931 6824
rect 882 6792 931 6804
rect 981 6828 1025 6834
rect 981 6808 996 6828
rect 1016 6808 1025 6828
rect 981 6792 1025 6808
rect 1095 6824 1144 6834
rect 1095 6804 1106 6824
rect 1126 6804 1144 6824
rect 1095 6792 1144 6804
rect 1194 6828 1238 6834
rect 1194 6808 1209 6828
rect 1229 6808 1238 6828
rect 1194 6792 1238 6808
rect 1303 6824 1352 6834
rect 1303 6804 1314 6824
rect 1334 6804 1352 6824
rect 1303 6792 1352 6804
rect 1402 6828 1446 6834
rect 1402 6808 1417 6828
rect 1437 6808 1446 6828
rect 1402 6792 1446 6808
rect 1516 6828 1560 6834
rect 1516 6808 1525 6828
rect 1545 6808 1560 6828
rect 1516 6792 1560 6808
rect 1610 6824 1659 6834
rect 9172 6921 9221 6931
rect 9271 6947 9315 6963
rect 9271 6927 9286 6947
rect 9306 6927 9315 6947
rect 9271 6921 9315 6927
rect 9385 6947 9429 6963
rect 9385 6927 9394 6947
rect 9414 6927 9429 6947
rect 9385 6921 9429 6927
rect 9479 6951 9528 6963
rect 9479 6931 9497 6951
rect 9517 6931 9528 6951
rect 9479 6921 9528 6931
rect 9593 6947 9637 6963
rect 9593 6927 9602 6947
rect 9622 6927 9637 6947
rect 9593 6921 9637 6927
rect 9687 6951 9736 6963
rect 9687 6931 9705 6951
rect 9725 6931 9736 6951
rect 9687 6921 9736 6931
rect 9806 6947 9850 6963
rect 9806 6927 9815 6947
rect 9835 6927 9850 6947
rect 9806 6921 9850 6927
rect 9900 6951 9949 6963
rect 9900 6931 9918 6951
rect 9938 6931 9949 6951
rect 9900 6921 9949 6931
rect 1610 6804 1628 6824
rect 1648 6804 1659 6824
rect 1610 6792 1659 6804
rect 3377 6819 3426 6829
rect 3377 6799 3388 6819
rect 3408 6799 3426 6819
rect 3377 6787 3426 6799
rect 3476 6823 3520 6829
rect 3476 6803 3491 6823
rect 3511 6803 3520 6823
rect 3476 6787 3520 6803
rect 3590 6819 3639 6829
rect 3590 6799 3601 6819
rect 3621 6799 3639 6819
rect 3590 6787 3639 6799
rect 3689 6823 3733 6829
rect 3689 6803 3704 6823
rect 3724 6803 3733 6823
rect 3689 6787 3733 6803
rect 3798 6819 3847 6829
rect 3798 6799 3809 6819
rect 3829 6799 3847 6819
rect 3798 6787 3847 6799
rect 3897 6823 3941 6829
rect 3897 6803 3912 6823
rect 3932 6803 3941 6823
rect 3897 6787 3941 6803
rect 4011 6823 4055 6829
rect 4011 6803 4020 6823
rect 4040 6803 4055 6823
rect 4011 6787 4055 6803
rect 4105 6819 4154 6829
rect 4105 6799 4123 6819
rect 4143 6799 4154 6819
rect 4105 6787 4154 6799
rect 18832 6949 18881 6961
rect 18832 6929 18843 6949
rect 18863 6929 18881 6949
rect 18832 6919 18881 6929
rect 18931 6945 18975 6961
rect 18931 6925 18946 6945
rect 18966 6925 18975 6945
rect 18931 6919 18975 6925
rect 19045 6945 19089 6961
rect 19045 6925 19054 6945
rect 19074 6925 19089 6945
rect 19045 6919 19089 6925
rect 19139 6949 19188 6961
rect 19139 6929 19157 6949
rect 19177 6929 19188 6949
rect 19139 6919 19188 6929
rect 19253 6945 19297 6961
rect 19253 6925 19262 6945
rect 19282 6925 19297 6945
rect 19253 6919 19297 6925
rect 19347 6949 19396 6961
rect 19347 6929 19365 6949
rect 19385 6929 19396 6949
rect 19347 6919 19396 6929
rect 19466 6945 19510 6961
rect 19466 6925 19475 6945
rect 19495 6925 19510 6945
rect 19466 6919 19510 6925
rect 19560 6949 19609 6961
rect 19560 6929 19578 6949
rect 19598 6929 19609 6949
rect 19560 6919 19609 6929
rect 19880 6945 19929 6957
rect 19880 6925 19891 6945
rect 19911 6925 19929 6945
rect 11590 6818 11639 6828
rect 11590 6798 11601 6818
rect 11621 6798 11639 6818
rect 11590 6786 11639 6798
rect 11689 6822 11733 6828
rect 11689 6802 11704 6822
rect 11724 6802 11733 6822
rect 11689 6786 11733 6802
rect 11803 6818 11852 6828
rect 11803 6798 11814 6818
rect 11834 6798 11852 6818
rect 11803 6786 11852 6798
rect 11902 6822 11946 6828
rect 11902 6802 11917 6822
rect 11937 6802 11946 6822
rect 11902 6786 11946 6802
rect 12011 6818 12060 6828
rect 12011 6798 12022 6818
rect 12042 6798 12060 6818
rect 12011 6786 12060 6798
rect 12110 6822 12154 6828
rect 12110 6802 12125 6822
rect 12145 6802 12154 6822
rect 12110 6786 12154 6802
rect 12224 6822 12268 6828
rect 12224 6802 12233 6822
rect 12253 6802 12268 6822
rect 12224 6786 12268 6802
rect 12318 6818 12367 6828
rect 19880 6915 19929 6925
rect 19979 6941 20023 6957
rect 19979 6921 19994 6941
rect 20014 6921 20023 6941
rect 19979 6915 20023 6921
rect 20093 6941 20137 6957
rect 20093 6921 20102 6941
rect 20122 6921 20137 6941
rect 20093 6915 20137 6921
rect 20187 6945 20236 6957
rect 20187 6925 20205 6945
rect 20225 6925 20236 6945
rect 20187 6915 20236 6925
rect 20301 6941 20345 6957
rect 20301 6921 20310 6941
rect 20330 6921 20345 6941
rect 20301 6915 20345 6921
rect 20395 6945 20444 6957
rect 20395 6925 20413 6945
rect 20433 6925 20444 6945
rect 20395 6915 20444 6925
rect 20514 6941 20558 6957
rect 20514 6921 20523 6941
rect 20543 6921 20558 6941
rect 20514 6915 20558 6921
rect 20608 6945 20657 6957
rect 20608 6925 20626 6945
rect 20646 6925 20657 6945
rect 20608 6915 20657 6925
rect 12318 6798 12336 6818
rect 12356 6798 12367 6818
rect 12318 6786 12367 6798
rect 14085 6813 14134 6823
rect 14085 6793 14096 6813
rect 14116 6793 14134 6813
rect 14085 6781 14134 6793
rect 14184 6817 14228 6823
rect 14184 6797 14199 6817
rect 14219 6797 14228 6817
rect 14184 6781 14228 6797
rect 14298 6813 14347 6823
rect 14298 6793 14309 6813
rect 14329 6793 14347 6813
rect 14298 6781 14347 6793
rect 14397 6817 14441 6823
rect 14397 6797 14412 6817
rect 14432 6797 14441 6817
rect 14397 6781 14441 6797
rect 14506 6813 14555 6823
rect 14506 6793 14517 6813
rect 14537 6793 14555 6813
rect 14506 6781 14555 6793
rect 14605 6817 14649 6823
rect 14605 6797 14620 6817
rect 14640 6797 14649 6817
rect 14605 6781 14649 6797
rect 14719 6817 14763 6823
rect 14719 6797 14728 6817
rect 14748 6797 14763 6817
rect 14719 6781 14763 6797
rect 14813 6813 14862 6823
rect 14813 6793 14831 6813
rect 14851 6793 14862 6813
rect 14813 6781 14862 6793
rect 29797 6953 29846 6965
rect 29797 6933 29808 6953
rect 29828 6933 29846 6953
rect 29797 6923 29846 6933
rect 29896 6949 29940 6965
rect 29896 6929 29911 6949
rect 29931 6929 29940 6949
rect 29896 6923 29940 6929
rect 30010 6949 30054 6965
rect 30010 6929 30019 6949
rect 30039 6929 30054 6949
rect 30010 6923 30054 6929
rect 30104 6953 30153 6965
rect 30104 6933 30122 6953
rect 30142 6933 30153 6953
rect 30104 6923 30153 6933
rect 30218 6949 30262 6965
rect 30218 6929 30227 6949
rect 30247 6929 30262 6949
rect 30218 6923 30262 6929
rect 30312 6953 30361 6965
rect 30312 6933 30330 6953
rect 30350 6933 30361 6953
rect 30312 6923 30361 6933
rect 30431 6949 30475 6965
rect 30431 6929 30440 6949
rect 30460 6929 30475 6949
rect 30431 6923 30475 6929
rect 30525 6953 30574 6965
rect 30525 6933 30543 6953
rect 30563 6933 30574 6953
rect 30525 6923 30574 6933
rect 30845 6949 30894 6961
rect 30845 6929 30856 6949
rect 30876 6929 30894 6949
rect 22555 6822 22604 6832
rect 22555 6802 22566 6822
rect 22586 6802 22604 6822
rect 22555 6790 22604 6802
rect 22654 6826 22698 6832
rect 22654 6806 22669 6826
rect 22689 6806 22698 6826
rect 22654 6790 22698 6806
rect 22768 6822 22817 6832
rect 22768 6802 22779 6822
rect 22799 6802 22817 6822
rect 22768 6790 22817 6802
rect 22867 6826 22911 6832
rect 22867 6806 22882 6826
rect 22902 6806 22911 6826
rect 22867 6790 22911 6806
rect 22976 6822 23025 6832
rect 22976 6802 22987 6822
rect 23007 6802 23025 6822
rect 22976 6790 23025 6802
rect 23075 6826 23119 6832
rect 23075 6806 23090 6826
rect 23110 6806 23119 6826
rect 23075 6790 23119 6806
rect 23189 6826 23233 6832
rect 23189 6806 23198 6826
rect 23218 6806 23233 6826
rect 23189 6790 23233 6806
rect 23283 6822 23332 6832
rect 30845 6919 30894 6929
rect 30944 6945 30988 6961
rect 30944 6925 30959 6945
rect 30979 6925 30988 6945
rect 30944 6919 30988 6925
rect 31058 6945 31102 6961
rect 31058 6925 31067 6945
rect 31087 6925 31102 6945
rect 31058 6919 31102 6925
rect 31152 6949 31201 6961
rect 31152 6929 31170 6949
rect 31190 6929 31201 6949
rect 31152 6919 31201 6929
rect 31266 6945 31310 6961
rect 31266 6925 31275 6945
rect 31295 6925 31310 6945
rect 31266 6919 31310 6925
rect 31360 6949 31409 6961
rect 31360 6929 31378 6949
rect 31398 6929 31409 6949
rect 31360 6919 31409 6929
rect 31479 6945 31523 6961
rect 31479 6925 31488 6945
rect 31508 6925 31523 6945
rect 31479 6919 31523 6925
rect 31573 6949 31622 6961
rect 31573 6929 31591 6949
rect 31611 6929 31622 6949
rect 31573 6919 31622 6929
rect 23283 6802 23301 6822
rect 23321 6802 23332 6822
rect 23283 6790 23332 6802
rect 25050 6817 25099 6827
rect 25050 6797 25061 6817
rect 25081 6797 25099 6817
rect 25050 6785 25099 6797
rect 25149 6821 25193 6827
rect 25149 6801 25164 6821
rect 25184 6801 25193 6821
rect 25149 6785 25193 6801
rect 25263 6817 25312 6827
rect 25263 6797 25274 6817
rect 25294 6797 25312 6817
rect 25263 6785 25312 6797
rect 25362 6821 25406 6827
rect 25362 6801 25377 6821
rect 25397 6801 25406 6821
rect 25362 6785 25406 6801
rect 25471 6817 25520 6827
rect 25471 6797 25482 6817
rect 25502 6797 25520 6817
rect 25471 6785 25520 6797
rect 25570 6821 25614 6827
rect 25570 6801 25585 6821
rect 25605 6801 25614 6821
rect 25570 6785 25614 6801
rect 25684 6821 25728 6827
rect 25684 6801 25693 6821
rect 25713 6801 25728 6821
rect 25684 6785 25728 6801
rect 25778 6817 25827 6827
rect 25778 6797 25796 6817
rect 25816 6797 25827 6817
rect 25778 6785 25827 6797
rect 40505 6947 40554 6959
rect 40505 6927 40516 6947
rect 40536 6927 40554 6947
rect 40505 6917 40554 6927
rect 40604 6943 40648 6959
rect 40604 6923 40619 6943
rect 40639 6923 40648 6943
rect 40604 6917 40648 6923
rect 40718 6943 40762 6959
rect 40718 6923 40727 6943
rect 40747 6923 40762 6943
rect 40718 6917 40762 6923
rect 40812 6947 40861 6959
rect 40812 6927 40830 6947
rect 40850 6927 40861 6947
rect 40812 6917 40861 6927
rect 40926 6943 40970 6959
rect 40926 6923 40935 6943
rect 40955 6923 40970 6943
rect 40926 6917 40970 6923
rect 41020 6947 41069 6959
rect 41020 6927 41038 6947
rect 41058 6927 41069 6947
rect 41020 6917 41069 6927
rect 41139 6943 41183 6959
rect 41139 6923 41148 6943
rect 41168 6923 41183 6943
rect 41139 6917 41183 6923
rect 41233 6947 41282 6959
rect 41233 6927 41251 6947
rect 41271 6927 41282 6947
rect 41233 6917 41282 6927
rect 41553 6943 41602 6955
rect 41553 6923 41564 6943
rect 41584 6923 41602 6943
rect 33263 6816 33312 6826
rect 33263 6796 33274 6816
rect 33294 6796 33312 6816
rect 33263 6784 33312 6796
rect 33362 6820 33406 6826
rect 33362 6800 33377 6820
rect 33397 6800 33406 6820
rect 33362 6784 33406 6800
rect 33476 6816 33525 6826
rect 33476 6796 33487 6816
rect 33507 6796 33525 6816
rect 33476 6784 33525 6796
rect 33575 6820 33619 6826
rect 33575 6800 33590 6820
rect 33610 6800 33619 6820
rect 33575 6784 33619 6800
rect 33684 6816 33733 6826
rect 33684 6796 33695 6816
rect 33715 6796 33733 6816
rect 33684 6784 33733 6796
rect 33783 6820 33827 6826
rect 33783 6800 33798 6820
rect 33818 6800 33827 6820
rect 33783 6784 33827 6800
rect 33897 6820 33941 6826
rect 33897 6800 33906 6820
rect 33926 6800 33941 6820
rect 33897 6784 33941 6800
rect 33991 6816 34040 6826
rect 41553 6913 41602 6923
rect 41652 6939 41696 6955
rect 41652 6919 41667 6939
rect 41687 6919 41696 6939
rect 41652 6913 41696 6919
rect 41766 6939 41810 6955
rect 41766 6919 41775 6939
rect 41795 6919 41810 6939
rect 41766 6913 41810 6919
rect 41860 6943 41909 6955
rect 41860 6923 41878 6943
rect 41898 6923 41909 6943
rect 41860 6913 41909 6923
rect 41974 6939 42018 6955
rect 41974 6919 41983 6939
rect 42003 6919 42018 6939
rect 41974 6913 42018 6919
rect 42068 6943 42117 6955
rect 42068 6923 42086 6943
rect 42106 6923 42117 6943
rect 42068 6913 42117 6923
rect 42187 6939 42231 6955
rect 42187 6919 42196 6939
rect 42216 6919 42231 6939
rect 42187 6913 42231 6919
rect 42281 6943 42330 6955
rect 42281 6923 42299 6943
rect 42319 6923 42330 6943
rect 42281 6913 42330 6923
rect 33991 6796 34009 6816
rect 34029 6796 34040 6816
rect 33991 6784 34040 6796
rect 35758 6811 35807 6821
rect 35758 6791 35769 6811
rect 35789 6791 35807 6811
rect 35758 6779 35807 6791
rect 35857 6815 35901 6821
rect 35857 6795 35872 6815
rect 35892 6795 35901 6815
rect 35857 6779 35901 6795
rect 35971 6811 36020 6821
rect 35971 6791 35982 6811
rect 36002 6791 36020 6811
rect 35971 6779 36020 6791
rect 36070 6815 36114 6821
rect 36070 6795 36085 6815
rect 36105 6795 36114 6815
rect 36070 6779 36114 6795
rect 36179 6811 36228 6821
rect 36179 6791 36190 6811
rect 36210 6791 36228 6811
rect 36179 6779 36228 6791
rect 36278 6815 36322 6821
rect 36278 6795 36293 6815
rect 36313 6795 36322 6815
rect 36278 6779 36322 6795
rect 36392 6815 36436 6821
rect 36392 6795 36401 6815
rect 36421 6795 36436 6815
rect 36392 6779 36436 6795
rect 36486 6811 36535 6821
rect 36486 6791 36504 6811
rect 36524 6791 36535 6811
rect 36486 6779 36535 6791
rect 6677 6188 6726 6200
rect 6677 6168 6688 6188
rect 6708 6168 6726 6188
rect 6677 6158 6726 6168
rect 6776 6184 6820 6200
rect 6776 6164 6791 6184
rect 6811 6164 6820 6184
rect 6776 6158 6820 6164
rect 6890 6184 6934 6200
rect 6890 6164 6899 6184
rect 6919 6164 6934 6184
rect 6890 6158 6934 6164
rect 6984 6188 7033 6200
rect 6984 6168 7002 6188
rect 7022 6168 7033 6188
rect 6984 6158 7033 6168
rect 7098 6184 7142 6200
rect 7098 6164 7107 6184
rect 7127 6164 7142 6184
rect 7098 6158 7142 6164
rect 7192 6188 7241 6200
rect 7192 6168 7210 6188
rect 7230 6168 7241 6188
rect 7192 6158 7241 6168
rect 7311 6184 7355 6200
rect 7311 6164 7320 6184
rect 7340 6164 7355 6184
rect 7311 6158 7355 6164
rect 7405 6188 7454 6200
rect 7405 6168 7423 6188
rect 7443 6168 7454 6188
rect 7405 6158 7454 6168
rect 9172 6183 9221 6195
rect 9172 6163 9183 6183
rect 9203 6163 9221 6183
rect 882 6056 931 6066
rect 882 6036 893 6056
rect 913 6036 931 6056
rect 882 6024 931 6036
rect 981 6060 1025 6066
rect 981 6040 996 6060
rect 1016 6040 1025 6060
rect 981 6024 1025 6040
rect 1095 6056 1144 6066
rect 1095 6036 1106 6056
rect 1126 6036 1144 6056
rect 1095 6024 1144 6036
rect 1194 6060 1238 6066
rect 1194 6040 1209 6060
rect 1229 6040 1238 6060
rect 1194 6024 1238 6040
rect 1303 6056 1352 6066
rect 1303 6036 1314 6056
rect 1334 6036 1352 6056
rect 1303 6024 1352 6036
rect 1402 6060 1446 6066
rect 1402 6040 1417 6060
rect 1437 6040 1446 6060
rect 1402 6024 1446 6040
rect 1516 6060 1560 6066
rect 1516 6040 1525 6060
rect 1545 6040 1560 6060
rect 1516 6024 1560 6040
rect 1610 6056 1659 6066
rect 9172 6153 9221 6163
rect 9271 6179 9315 6195
rect 9271 6159 9286 6179
rect 9306 6159 9315 6179
rect 9271 6153 9315 6159
rect 9385 6179 9429 6195
rect 9385 6159 9394 6179
rect 9414 6159 9429 6179
rect 9385 6153 9429 6159
rect 9479 6183 9528 6195
rect 9479 6163 9497 6183
rect 9517 6163 9528 6183
rect 9479 6153 9528 6163
rect 9593 6179 9637 6195
rect 9593 6159 9602 6179
rect 9622 6159 9637 6179
rect 9593 6153 9637 6159
rect 9687 6183 9736 6195
rect 9687 6163 9705 6183
rect 9725 6163 9736 6183
rect 9687 6153 9736 6163
rect 9806 6179 9850 6195
rect 9806 6159 9815 6179
rect 9835 6159 9850 6179
rect 9806 6153 9850 6159
rect 9900 6183 9949 6195
rect 9900 6163 9918 6183
rect 9938 6163 9949 6183
rect 9900 6153 9949 6163
rect 1610 6036 1628 6056
rect 1648 6036 1659 6056
rect 1610 6024 1659 6036
rect 1930 6052 1979 6062
rect 1930 6032 1941 6052
rect 1961 6032 1979 6052
rect 1930 6020 1979 6032
rect 2029 6056 2073 6062
rect 2029 6036 2044 6056
rect 2064 6036 2073 6056
rect 2029 6020 2073 6036
rect 2143 6052 2192 6062
rect 2143 6032 2154 6052
rect 2174 6032 2192 6052
rect 2143 6020 2192 6032
rect 2242 6056 2286 6062
rect 2242 6036 2257 6056
rect 2277 6036 2286 6056
rect 2242 6020 2286 6036
rect 2351 6052 2400 6062
rect 2351 6032 2362 6052
rect 2382 6032 2400 6052
rect 2351 6020 2400 6032
rect 2450 6056 2494 6062
rect 2450 6036 2465 6056
rect 2485 6036 2494 6056
rect 2450 6020 2494 6036
rect 2564 6056 2608 6062
rect 2564 6036 2573 6056
rect 2593 6036 2608 6056
rect 2564 6020 2608 6036
rect 2658 6052 2707 6062
rect 2658 6032 2676 6052
rect 2696 6032 2707 6052
rect 2658 6020 2707 6032
rect 17385 6182 17434 6194
rect 17385 6162 17396 6182
rect 17416 6162 17434 6182
rect 17385 6152 17434 6162
rect 17484 6178 17528 6194
rect 17484 6158 17499 6178
rect 17519 6158 17528 6178
rect 17484 6152 17528 6158
rect 17598 6178 17642 6194
rect 17598 6158 17607 6178
rect 17627 6158 17642 6178
rect 17598 6152 17642 6158
rect 17692 6182 17741 6194
rect 17692 6162 17710 6182
rect 17730 6162 17741 6182
rect 17692 6152 17741 6162
rect 17806 6178 17850 6194
rect 17806 6158 17815 6178
rect 17835 6158 17850 6178
rect 17806 6152 17850 6158
rect 17900 6182 17949 6194
rect 17900 6162 17918 6182
rect 17938 6162 17949 6182
rect 17900 6152 17949 6162
rect 18019 6178 18063 6194
rect 18019 6158 18028 6178
rect 18048 6158 18063 6178
rect 18019 6152 18063 6158
rect 18113 6182 18162 6194
rect 18113 6162 18131 6182
rect 18151 6162 18162 6182
rect 18113 6152 18162 6162
rect 19880 6177 19929 6189
rect 19880 6157 19891 6177
rect 19911 6157 19929 6177
rect 11590 6050 11639 6060
rect 11590 6030 11601 6050
rect 11621 6030 11639 6050
rect 11590 6018 11639 6030
rect 11689 6054 11733 6060
rect 11689 6034 11704 6054
rect 11724 6034 11733 6054
rect 11689 6018 11733 6034
rect 11803 6050 11852 6060
rect 11803 6030 11814 6050
rect 11834 6030 11852 6050
rect 11803 6018 11852 6030
rect 11902 6054 11946 6060
rect 11902 6034 11917 6054
rect 11937 6034 11946 6054
rect 11902 6018 11946 6034
rect 12011 6050 12060 6060
rect 12011 6030 12022 6050
rect 12042 6030 12060 6050
rect 12011 6018 12060 6030
rect 12110 6054 12154 6060
rect 12110 6034 12125 6054
rect 12145 6034 12154 6054
rect 12110 6018 12154 6034
rect 12224 6054 12268 6060
rect 12224 6034 12233 6054
rect 12253 6034 12268 6054
rect 12224 6018 12268 6034
rect 12318 6050 12367 6060
rect 19880 6147 19929 6157
rect 19979 6173 20023 6189
rect 19979 6153 19994 6173
rect 20014 6153 20023 6173
rect 19979 6147 20023 6153
rect 20093 6173 20137 6189
rect 20093 6153 20102 6173
rect 20122 6153 20137 6173
rect 20093 6147 20137 6153
rect 20187 6177 20236 6189
rect 20187 6157 20205 6177
rect 20225 6157 20236 6177
rect 20187 6147 20236 6157
rect 20301 6173 20345 6189
rect 20301 6153 20310 6173
rect 20330 6153 20345 6173
rect 20301 6147 20345 6153
rect 20395 6177 20444 6189
rect 20395 6157 20413 6177
rect 20433 6157 20444 6177
rect 20395 6147 20444 6157
rect 20514 6173 20558 6189
rect 20514 6153 20523 6173
rect 20543 6153 20558 6173
rect 20514 6147 20558 6153
rect 20608 6177 20657 6189
rect 20608 6157 20626 6177
rect 20646 6157 20657 6177
rect 20608 6147 20657 6157
rect 12318 6030 12336 6050
rect 12356 6030 12367 6050
rect 12318 6018 12367 6030
rect 12638 6046 12687 6056
rect 12638 6026 12649 6046
rect 12669 6026 12687 6046
rect 12638 6014 12687 6026
rect 12737 6050 12781 6056
rect 12737 6030 12752 6050
rect 12772 6030 12781 6050
rect 12737 6014 12781 6030
rect 12851 6046 12900 6056
rect 12851 6026 12862 6046
rect 12882 6026 12900 6046
rect 12851 6014 12900 6026
rect 12950 6050 12994 6056
rect 12950 6030 12965 6050
rect 12985 6030 12994 6050
rect 12950 6014 12994 6030
rect 13059 6046 13108 6056
rect 13059 6026 13070 6046
rect 13090 6026 13108 6046
rect 13059 6014 13108 6026
rect 13158 6050 13202 6056
rect 13158 6030 13173 6050
rect 13193 6030 13202 6050
rect 13158 6014 13202 6030
rect 13272 6050 13316 6056
rect 13272 6030 13281 6050
rect 13301 6030 13316 6050
rect 13272 6014 13316 6030
rect 13366 6046 13415 6056
rect 13366 6026 13384 6046
rect 13404 6026 13415 6046
rect 13366 6014 13415 6026
rect 28350 6186 28399 6198
rect 28350 6166 28361 6186
rect 28381 6166 28399 6186
rect 28350 6156 28399 6166
rect 28449 6182 28493 6198
rect 28449 6162 28464 6182
rect 28484 6162 28493 6182
rect 28449 6156 28493 6162
rect 28563 6182 28607 6198
rect 28563 6162 28572 6182
rect 28592 6162 28607 6182
rect 28563 6156 28607 6162
rect 28657 6186 28706 6198
rect 28657 6166 28675 6186
rect 28695 6166 28706 6186
rect 28657 6156 28706 6166
rect 28771 6182 28815 6198
rect 28771 6162 28780 6182
rect 28800 6162 28815 6182
rect 28771 6156 28815 6162
rect 28865 6186 28914 6198
rect 28865 6166 28883 6186
rect 28903 6166 28914 6186
rect 28865 6156 28914 6166
rect 28984 6182 29028 6198
rect 28984 6162 28993 6182
rect 29013 6162 29028 6182
rect 28984 6156 29028 6162
rect 29078 6186 29127 6198
rect 29078 6166 29096 6186
rect 29116 6166 29127 6186
rect 29078 6156 29127 6166
rect 30845 6181 30894 6193
rect 30845 6161 30856 6181
rect 30876 6161 30894 6181
rect 22555 6054 22604 6064
rect 22555 6034 22566 6054
rect 22586 6034 22604 6054
rect 22555 6022 22604 6034
rect 22654 6058 22698 6064
rect 22654 6038 22669 6058
rect 22689 6038 22698 6058
rect 22654 6022 22698 6038
rect 22768 6054 22817 6064
rect 22768 6034 22779 6054
rect 22799 6034 22817 6054
rect 22768 6022 22817 6034
rect 22867 6058 22911 6064
rect 22867 6038 22882 6058
rect 22902 6038 22911 6058
rect 22867 6022 22911 6038
rect 22976 6054 23025 6064
rect 22976 6034 22987 6054
rect 23007 6034 23025 6054
rect 22976 6022 23025 6034
rect 23075 6058 23119 6064
rect 23075 6038 23090 6058
rect 23110 6038 23119 6058
rect 23075 6022 23119 6038
rect 23189 6058 23233 6064
rect 23189 6038 23198 6058
rect 23218 6038 23233 6058
rect 23189 6022 23233 6038
rect 23283 6054 23332 6064
rect 30845 6151 30894 6161
rect 30944 6177 30988 6193
rect 30944 6157 30959 6177
rect 30979 6157 30988 6177
rect 30944 6151 30988 6157
rect 31058 6177 31102 6193
rect 31058 6157 31067 6177
rect 31087 6157 31102 6177
rect 31058 6151 31102 6157
rect 31152 6181 31201 6193
rect 31152 6161 31170 6181
rect 31190 6161 31201 6181
rect 31152 6151 31201 6161
rect 31266 6177 31310 6193
rect 31266 6157 31275 6177
rect 31295 6157 31310 6177
rect 31266 6151 31310 6157
rect 31360 6181 31409 6193
rect 31360 6161 31378 6181
rect 31398 6161 31409 6181
rect 31360 6151 31409 6161
rect 31479 6177 31523 6193
rect 31479 6157 31488 6177
rect 31508 6157 31523 6177
rect 31479 6151 31523 6157
rect 31573 6181 31622 6193
rect 31573 6161 31591 6181
rect 31611 6161 31622 6181
rect 31573 6151 31622 6161
rect 23283 6034 23301 6054
rect 23321 6034 23332 6054
rect 23283 6022 23332 6034
rect 23603 6050 23652 6060
rect 23603 6030 23614 6050
rect 23634 6030 23652 6050
rect 23603 6018 23652 6030
rect 23702 6054 23746 6060
rect 23702 6034 23717 6054
rect 23737 6034 23746 6054
rect 23702 6018 23746 6034
rect 23816 6050 23865 6060
rect 23816 6030 23827 6050
rect 23847 6030 23865 6050
rect 23816 6018 23865 6030
rect 23915 6054 23959 6060
rect 23915 6034 23930 6054
rect 23950 6034 23959 6054
rect 23915 6018 23959 6034
rect 24024 6050 24073 6060
rect 24024 6030 24035 6050
rect 24055 6030 24073 6050
rect 24024 6018 24073 6030
rect 24123 6054 24167 6060
rect 24123 6034 24138 6054
rect 24158 6034 24167 6054
rect 24123 6018 24167 6034
rect 24237 6054 24281 6060
rect 24237 6034 24246 6054
rect 24266 6034 24281 6054
rect 24237 6018 24281 6034
rect 24331 6050 24380 6060
rect 24331 6030 24349 6050
rect 24369 6030 24380 6050
rect 24331 6018 24380 6030
rect 39058 6180 39107 6192
rect 39058 6160 39069 6180
rect 39089 6160 39107 6180
rect 39058 6150 39107 6160
rect 39157 6176 39201 6192
rect 39157 6156 39172 6176
rect 39192 6156 39201 6176
rect 39157 6150 39201 6156
rect 39271 6176 39315 6192
rect 39271 6156 39280 6176
rect 39300 6156 39315 6176
rect 39271 6150 39315 6156
rect 39365 6180 39414 6192
rect 39365 6160 39383 6180
rect 39403 6160 39414 6180
rect 39365 6150 39414 6160
rect 39479 6176 39523 6192
rect 39479 6156 39488 6176
rect 39508 6156 39523 6176
rect 39479 6150 39523 6156
rect 39573 6180 39622 6192
rect 39573 6160 39591 6180
rect 39611 6160 39622 6180
rect 39573 6150 39622 6160
rect 39692 6176 39736 6192
rect 39692 6156 39701 6176
rect 39721 6156 39736 6176
rect 39692 6150 39736 6156
rect 39786 6180 39835 6192
rect 39786 6160 39804 6180
rect 39824 6160 39835 6180
rect 39786 6150 39835 6160
rect 41553 6175 41602 6187
rect 41553 6155 41564 6175
rect 41584 6155 41602 6175
rect 33263 6048 33312 6058
rect 33263 6028 33274 6048
rect 33294 6028 33312 6048
rect 33263 6016 33312 6028
rect 33362 6052 33406 6058
rect 33362 6032 33377 6052
rect 33397 6032 33406 6052
rect 33362 6016 33406 6032
rect 33476 6048 33525 6058
rect 33476 6028 33487 6048
rect 33507 6028 33525 6048
rect 33476 6016 33525 6028
rect 33575 6052 33619 6058
rect 33575 6032 33590 6052
rect 33610 6032 33619 6052
rect 33575 6016 33619 6032
rect 33684 6048 33733 6058
rect 33684 6028 33695 6048
rect 33715 6028 33733 6048
rect 33684 6016 33733 6028
rect 33783 6052 33827 6058
rect 33783 6032 33798 6052
rect 33818 6032 33827 6052
rect 33783 6016 33827 6032
rect 33897 6052 33941 6058
rect 33897 6032 33906 6052
rect 33926 6032 33941 6052
rect 33897 6016 33941 6032
rect 33991 6048 34040 6058
rect 41553 6145 41602 6155
rect 41652 6171 41696 6187
rect 41652 6151 41667 6171
rect 41687 6151 41696 6171
rect 41652 6145 41696 6151
rect 41766 6171 41810 6187
rect 41766 6151 41775 6171
rect 41795 6151 41810 6171
rect 41766 6145 41810 6151
rect 41860 6175 41909 6187
rect 41860 6155 41878 6175
rect 41898 6155 41909 6175
rect 41860 6145 41909 6155
rect 41974 6171 42018 6187
rect 41974 6151 41983 6171
rect 42003 6151 42018 6171
rect 41974 6145 42018 6151
rect 42068 6175 42117 6187
rect 42068 6155 42086 6175
rect 42106 6155 42117 6175
rect 42068 6145 42117 6155
rect 42187 6171 42231 6187
rect 42187 6151 42196 6171
rect 42216 6151 42231 6171
rect 42187 6145 42231 6151
rect 42281 6175 42330 6187
rect 42281 6155 42299 6175
rect 42319 6155 42330 6175
rect 42281 6145 42330 6155
rect 33991 6028 34009 6048
rect 34029 6028 34040 6048
rect 33991 6016 34040 6028
rect 34311 6044 34360 6054
rect 34311 6024 34322 6044
rect 34342 6024 34360 6044
rect 34311 6012 34360 6024
rect 34410 6048 34454 6054
rect 34410 6028 34425 6048
rect 34445 6028 34454 6048
rect 34410 6012 34454 6028
rect 34524 6044 34573 6054
rect 34524 6024 34535 6044
rect 34555 6024 34573 6044
rect 34524 6012 34573 6024
rect 34623 6048 34667 6054
rect 34623 6028 34638 6048
rect 34658 6028 34667 6048
rect 34623 6012 34667 6028
rect 34732 6044 34781 6054
rect 34732 6024 34743 6044
rect 34763 6024 34781 6044
rect 34732 6012 34781 6024
rect 34831 6048 34875 6054
rect 34831 6028 34846 6048
rect 34866 6028 34875 6048
rect 34831 6012 34875 6028
rect 34945 6048 34989 6054
rect 34945 6028 34954 6048
rect 34974 6028 34989 6048
rect 34945 6012 34989 6028
rect 35039 6044 35088 6054
rect 35039 6024 35057 6044
rect 35077 6024 35088 6044
rect 35039 6012 35088 6024
rect 8124 5508 8173 5520
rect 8124 5488 8135 5508
rect 8155 5488 8173 5508
rect 8124 5478 8173 5488
rect 8223 5504 8267 5520
rect 8223 5484 8238 5504
rect 8258 5484 8267 5504
rect 8223 5478 8267 5484
rect 8337 5504 8381 5520
rect 8337 5484 8346 5504
rect 8366 5484 8381 5504
rect 8337 5478 8381 5484
rect 8431 5508 8480 5520
rect 8431 5488 8449 5508
rect 8469 5488 8480 5508
rect 8431 5478 8480 5488
rect 8545 5504 8589 5520
rect 8545 5484 8554 5504
rect 8574 5484 8589 5504
rect 8545 5478 8589 5484
rect 8639 5508 8688 5520
rect 8639 5488 8657 5508
rect 8677 5488 8688 5508
rect 8639 5478 8688 5488
rect 8758 5504 8802 5520
rect 8758 5484 8767 5504
rect 8787 5484 8802 5504
rect 8758 5478 8802 5484
rect 8852 5508 8901 5520
rect 8852 5488 8870 5508
rect 8890 5488 8901 5508
rect 8852 5478 8901 5488
rect 9172 5504 9221 5516
rect 9172 5484 9183 5504
rect 9203 5484 9221 5504
rect 882 5377 931 5387
rect 882 5357 893 5377
rect 913 5357 931 5377
rect 882 5345 931 5357
rect 981 5381 1025 5387
rect 981 5361 996 5381
rect 1016 5361 1025 5381
rect 981 5345 1025 5361
rect 1095 5377 1144 5387
rect 1095 5357 1106 5377
rect 1126 5357 1144 5377
rect 1095 5345 1144 5357
rect 1194 5381 1238 5387
rect 1194 5361 1209 5381
rect 1229 5361 1238 5381
rect 1194 5345 1238 5361
rect 1303 5377 1352 5387
rect 1303 5357 1314 5377
rect 1334 5357 1352 5377
rect 1303 5345 1352 5357
rect 1402 5381 1446 5387
rect 1402 5361 1417 5381
rect 1437 5361 1446 5381
rect 1402 5345 1446 5361
rect 1516 5381 1560 5387
rect 1516 5361 1525 5381
rect 1545 5361 1560 5381
rect 1516 5345 1560 5361
rect 1610 5377 1659 5387
rect 9172 5474 9221 5484
rect 9271 5500 9315 5516
rect 9271 5480 9286 5500
rect 9306 5480 9315 5500
rect 9271 5474 9315 5480
rect 9385 5500 9429 5516
rect 9385 5480 9394 5500
rect 9414 5480 9429 5500
rect 9385 5474 9429 5480
rect 9479 5504 9528 5516
rect 9479 5484 9497 5504
rect 9517 5484 9528 5504
rect 9479 5474 9528 5484
rect 9593 5500 9637 5516
rect 9593 5480 9602 5500
rect 9622 5480 9637 5500
rect 9593 5474 9637 5480
rect 9687 5504 9736 5516
rect 9687 5484 9705 5504
rect 9725 5484 9736 5504
rect 9687 5474 9736 5484
rect 9806 5500 9850 5516
rect 9806 5480 9815 5500
rect 9835 5480 9850 5500
rect 9806 5474 9850 5480
rect 9900 5504 9949 5516
rect 9900 5484 9918 5504
rect 9938 5484 9949 5504
rect 9900 5474 9949 5484
rect 1610 5357 1628 5377
rect 1648 5357 1659 5377
rect 1610 5345 1659 5357
rect 3420 5374 3469 5384
rect 3420 5354 3431 5374
rect 3451 5354 3469 5374
rect 3420 5342 3469 5354
rect 3519 5378 3563 5384
rect 3519 5358 3534 5378
rect 3554 5358 3563 5378
rect 3519 5342 3563 5358
rect 3633 5374 3682 5384
rect 3633 5354 3644 5374
rect 3664 5354 3682 5374
rect 3633 5342 3682 5354
rect 3732 5378 3776 5384
rect 3732 5358 3747 5378
rect 3767 5358 3776 5378
rect 3732 5342 3776 5358
rect 3841 5374 3890 5384
rect 3841 5354 3852 5374
rect 3872 5354 3890 5374
rect 3841 5342 3890 5354
rect 3940 5378 3984 5384
rect 3940 5358 3955 5378
rect 3975 5358 3984 5378
rect 3940 5342 3984 5358
rect 4054 5378 4098 5384
rect 4054 5358 4063 5378
rect 4083 5358 4098 5378
rect 4054 5342 4098 5358
rect 4148 5374 4197 5384
rect 4148 5354 4166 5374
rect 4186 5354 4197 5374
rect 4148 5342 4197 5354
rect 18832 5502 18881 5514
rect 18832 5482 18843 5502
rect 18863 5482 18881 5502
rect 18832 5472 18881 5482
rect 18931 5498 18975 5514
rect 18931 5478 18946 5498
rect 18966 5478 18975 5498
rect 18931 5472 18975 5478
rect 19045 5498 19089 5514
rect 19045 5478 19054 5498
rect 19074 5478 19089 5498
rect 19045 5472 19089 5478
rect 19139 5502 19188 5514
rect 19139 5482 19157 5502
rect 19177 5482 19188 5502
rect 19139 5472 19188 5482
rect 19253 5498 19297 5514
rect 19253 5478 19262 5498
rect 19282 5478 19297 5498
rect 19253 5472 19297 5478
rect 19347 5502 19396 5514
rect 19347 5482 19365 5502
rect 19385 5482 19396 5502
rect 19347 5472 19396 5482
rect 19466 5498 19510 5514
rect 19466 5478 19475 5498
rect 19495 5478 19510 5498
rect 19466 5472 19510 5478
rect 19560 5502 19609 5514
rect 19560 5482 19578 5502
rect 19598 5482 19609 5502
rect 19560 5472 19609 5482
rect 19880 5498 19929 5510
rect 19880 5478 19891 5498
rect 19911 5478 19929 5498
rect 11590 5371 11639 5381
rect 11590 5351 11601 5371
rect 11621 5351 11639 5371
rect 11590 5339 11639 5351
rect 11689 5375 11733 5381
rect 11689 5355 11704 5375
rect 11724 5355 11733 5375
rect 11689 5339 11733 5355
rect 11803 5371 11852 5381
rect 11803 5351 11814 5371
rect 11834 5351 11852 5371
rect 11803 5339 11852 5351
rect 11902 5375 11946 5381
rect 11902 5355 11917 5375
rect 11937 5355 11946 5375
rect 11902 5339 11946 5355
rect 12011 5371 12060 5381
rect 12011 5351 12022 5371
rect 12042 5351 12060 5371
rect 12011 5339 12060 5351
rect 12110 5375 12154 5381
rect 12110 5355 12125 5375
rect 12145 5355 12154 5375
rect 12110 5339 12154 5355
rect 12224 5375 12268 5381
rect 12224 5355 12233 5375
rect 12253 5355 12268 5375
rect 12224 5339 12268 5355
rect 12318 5371 12367 5381
rect 19880 5468 19929 5478
rect 19979 5494 20023 5510
rect 19979 5474 19994 5494
rect 20014 5474 20023 5494
rect 19979 5468 20023 5474
rect 20093 5494 20137 5510
rect 20093 5474 20102 5494
rect 20122 5474 20137 5494
rect 20093 5468 20137 5474
rect 20187 5498 20236 5510
rect 20187 5478 20205 5498
rect 20225 5478 20236 5498
rect 20187 5468 20236 5478
rect 20301 5494 20345 5510
rect 20301 5474 20310 5494
rect 20330 5474 20345 5494
rect 20301 5468 20345 5474
rect 20395 5498 20444 5510
rect 20395 5478 20413 5498
rect 20433 5478 20444 5498
rect 20395 5468 20444 5478
rect 20514 5494 20558 5510
rect 20514 5474 20523 5494
rect 20543 5474 20558 5494
rect 20514 5468 20558 5474
rect 20608 5498 20657 5510
rect 20608 5478 20626 5498
rect 20646 5478 20657 5498
rect 20608 5468 20657 5478
rect 12318 5351 12336 5371
rect 12356 5351 12367 5371
rect 12318 5339 12367 5351
rect 14128 5368 14177 5378
rect 14128 5348 14139 5368
rect 14159 5348 14177 5368
rect 14128 5336 14177 5348
rect 14227 5372 14271 5378
rect 14227 5352 14242 5372
rect 14262 5352 14271 5372
rect 14227 5336 14271 5352
rect 14341 5368 14390 5378
rect 14341 5348 14352 5368
rect 14372 5348 14390 5368
rect 14341 5336 14390 5348
rect 14440 5372 14484 5378
rect 14440 5352 14455 5372
rect 14475 5352 14484 5372
rect 14440 5336 14484 5352
rect 14549 5368 14598 5378
rect 14549 5348 14560 5368
rect 14580 5348 14598 5368
rect 14549 5336 14598 5348
rect 14648 5372 14692 5378
rect 14648 5352 14663 5372
rect 14683 5352 14692 5372
rect 14648 5336 14692 5352
rect 14762 5372 14806 5378
rect 14762 5352 14771 5372
rect 14791 5352 14806 5372
rect 14762 5336 14806 5352
rect 14856 5368 14905 5378
rect 14856 5348 14874 5368
rect 14894 5348 14905 5368
rect 14856 5336 14905 5348
rect 29797 5506 29846 5518
rect 29797 5486 29808 5506
rect 29828 5486 29846 5506
rect 29797 5476 29846 5486
rect 29896 5502 29940 5518
rect 29896 5482 29911 5502
rect 29931 5482 29940 5502
rect 29896 5476 29940 5482
rect 30010 5502 30054 5518
rect 30010 5482 30019 5502
rect 30039 5482 30054 5502
rect 30010 5476 30054 5482
rect 30104 5506 30153 5518
rect 30104 5486 30122 5506
rect 30142 5486 30153 5506
rect 30104 5476 30153 5486
rect 30218 5502 30262 5518
rect 30218 5482 30227 5502
rect 30247 5482 30262 5502
rect 30218 5476 30262 5482
rect 30312 5506 30361 5518
rect 30312 5486 30330 5506
rect 30350 5486 30361 5506
rect 30312 5476 30361 5486
rect 30431 5502 30475 5518
rect 30431 5482 30440 5502
rect 30460 5482 30475 5502
rect 30431 5476 30475 5482
rect 30525 5506 30574 5518
rect 30525 5486 30543 5506
rect 30563 5486 30574 5506
rect 30525 5476 30574 5486
rect 30845 5502 30894 5514
rect 30845 5482 30856 5502
rect 30876 5482 30894 5502
rect 22555 5375 22604 5385
rect 22555 5355 22566 5375
rect 22586 5355 22604 5375
rect 22555 5343 22604 5355
rect 22654 5379 22698 5385
rect 22654 5359 22669 5379
rect 22689 5359 22698 5379
rect 22654 5343 22698 5359
rect 22768 5375 22817 5385
rect 22768 5355 22779 5375
rect 22799 5355 22817 5375
rect 22768 5343 22817 5355
rect 22867 5379 22911 5385
rect 22867 5359 22882 5379
rect 22902 5359 22911 5379
rect 22867 5343 22911 5359
rect 22976 5375 23025 5385
rect 22976 5355 22987 5375
rect 23007 5355 23025 5375
rect 22976 5343 23025 5355
rect 23075 5379 23119 5385
rect 23075 5359 23090 5379
rect 23110 5359 23119 5379
rect 23075 5343 23119 5359
rect 23189 5379 23233 5385
rect 23189 5359 23198 5379
rect 23218 5359 23233 5379
rect 23189 5343 23233 5359
rect 23283 5375 23332 5385
rect 30845 5472 30894 5482
rect 30944 5498 30988 5514
rect 30944 5478 30959 5498
rect 30979 5478 30988 5498
rect 30944 5472 30988 5478
rect 31058 5498 31102 5514
rect 31058 5478 31067 5498
rect 31087 5478 31102 5498
rect 31058 5472 31102 5478
rect 31152 5502 31201 5514
rect 31152 5482 31170 5502
rect 31190 5482 31201 5502
rect 31152 5472 31201 5482
rect 31266 5498 31310 5514
rect 31266 5478 31275 5498
rect 31295 5478 31310 5498
rect 31266 5472 31310 5478
rect 31360 5502 31409 5514
rect 31360 5482 31378 5502
rect 31398 5482 31409 5502
rect 31360 5472 31409 5482
rect 31479 5498 31523 5514
rect 31479 5478 31488 5498
rect 31508 5478 31523 5498
rect 31479 5472 31523 5478
rect 31573 5502 31622 5514
rect 31573 5482 31591 5502
rect 31611 5482 31622 5502
rect 31573 5472 31622 5482
rect 23283 5355 23301 5375
rect 23321 5355 23332 5375
rect 23283 5343 23332 5355
rect 25093 5372 25142 5382
rect 25093 5352 25104 5372
rect 25124 5352 25142 5372
rect 25093 5340 25142 5352
rect 25192 5376 25236 5382
rect 25192 5356 25207 5376
rect 25227 5356 25236 5376
rect 25192 5340 25236 5356
rect 25306 5372 25355 5382
rect 25306 5352 25317 5372
rect 25337 5352 25355 5372
rect 25306 5340 25355 5352
rect 25405 5376 25449 5382
rect 25405 5356 25420 5376
rect 25440 5356 25449 5376
rect 25405 5340 25449 5356
rect 25514 5372 25563 5382
rect 25514 5352 25525 5372
rect 25545 5352 25563 5372
rect 25514 5340 25563 5352
rect 25613 5376 25657 5382
rect 25613 5356 25628 5376
rect 25648 5356 25657 5376
rect 25613 5340 25657 5356
rect 25727 5376 25771 5382
rect 25727 5356 25736 5376
rect 25756 5356 25771 5376
rect 25727 5340 25771 5356
rect 25821 5372 25870 5382
rect 25821 5352 25839 5372
rect 25859 5352 25870 5372
rect 25821 5340 25870 5352
rect 40505 5500 40554 5512
rect 40505 5480 40516 5500
rect 40536 5480 40554 5500
rect 40505 5470 40554 5480
rect 40604 5496 40648 5512
rect 40604 5476 40619 5496
rect 40639 5476 40648 5496
rect 40604 5470 40648 5476
rect 40718 5496 40762 5512
rect 40718 5476 40727 5496
rect 40747 5476 40762 5496
rect 40718 5470 40762 5476
rect 40812 5500 40861 5512
rect 40812 5480 40830 5500
rect 40850 5480 40861 5500
rect 40812 5470 40861 5480
rect 40926 5496 40970 5512
rect 40926 5476 40935 5496
rect 40955 5476 40970 5496
rect 40926 5470 40970 5476
rect 41020 5500 41069 5512
rect 41020 5480 41038 5500
rect 41058 5480 41069 5500
rect 41020 5470 41069 5480
rect 41139 5496 41183 5512
rect 41139 5476 41148 5496
rect 41168 5476 41183 5496
rect 41139 5470 41183 5476
rect 41233 5500 41282 5512
rect 41233 5480 41251 5500
rect 41271 5480 41282 5500
rect 41233 5470 41282 5480
rect 41553 5496 41602 5508
rect 41553 5476 41564 5496
rect 41584 5476 41602 5496
rect 33263 5369 33312 5379
rect 33263 5349 33274 5369
rect 33294 5349 33312 5369
rect 33263 5337 33312 5349
rect 33362 5373 33406 5379
rect 33362 5353 33377 5373
rect 33397 5353 33406 5373
rect 33362 5337 33406 5353
rect 33476 5369 33525 5379
rect 33476 5349 33487 5369
rect 33507 5349 33525 5369
rect 33476 5337 33525 5349
rect 33575 5373 33619 5379
rect 33575 5353 33590 5373
rect 33610 5353 33619 5373
rect 33575 5337 33619 5353
rect 33684 5369 33733 5379
rect 33684 5349 33695 5369
rect 33715 5349 33733 5369
rect 33684 5337 33733 5349
rect 33783 5373 33827 5379
rect 33783 5353 33798 5373
rect 33818 5353 33827 5373
rect 33783 5337 33827 5353
rect 33897 5373 33941 5379
rect 33897 5353 33906 5373
rect 33926 5353 33941 5373
rect 33897 5337 33941 5353
rect 33991 5369 34040 5379
rect 41553 5466 41602 5476
rect 41652 5492 41696 5508
rect 41652 5472 41667 5492
rect 41687 5472 41696 5492
rect 41652 5466 41696 5472
rect 41766 5492 41810 5508
rect 41766 5472 41775 5492
rect 41795 5472 41810 5492
rect 41766 5466 41810 5472
rect 41860 5496 41909 5508
rect 41860 5476 41878 5496
rect 41898 5476 41909 5496
rect 41860 5466 41909 5476
rect 41974 5492 42018 5508
rect 41974 5472 41983 5492
rect 42003 5472 42018 5492
rect 41974 5466 42018 5472
rect 42068 5496 42117 5508
rect 42068 5476 42086 5496
rect 42106 5476 42117 5496
rect 42068 5466 42117 5476
rect 42187 5492 42231 5508
rect 42187 5472 42196 5492
rect 42216 5472 42231 5492
rect 42187 5466 42231 5472
rect 42281 5496 42330 5508
rect 42281 5476 42299 5496
rect 42319 5476 42330 5496
rect 42281 5466 42330 5476
rect 33991 5349 34009 5369
rect 34029 5349 34040 5369
rect 33991 5337 34040 5349
rect 35801 5366 35850 5376
rect 35801 5346 35812 5366
rect 35832 5346 35850 5366
rect 35801 5334 35850 5346
rect 35900 5370 35944 5376
rect 35900 5350 35915 5370
rect 35935 5350 35944 5370
rect 35900 5334 35944 5350
rect 36014 5366 36063 5376
rect 36014 5346 36025 5366
rect 36045 5346 36063 5366
rect 36014 5334 36063 5346
rect 36113 5370 36157 5376
rect 36113 5350 36128 5370
rect 36148 5350 36157 5370
rect 36113 5334 36157 5350
rect 36222 5366 36271 5376
rect 36222 5346 36233 5366
rect 36253 5346 36271 5366
rect 36222 5334 36271 5346
rect 36321 5370 36365 5376
rect 36321 5350 36336 5370
rect 36356 5350 36365 5370
rect 36321 5334 36365 5350
rect 36435 5370 36479 5376
rect 36435 5350 36444 5370
rect 36464 5350 36479 5370
rect 36435 5334 36479 5350
rect 36529 5366 36578 5376
rect 36529 5346 36547 5366
rect 36567 5346 36578 5366
rect 36529 5334 36578 5346
rect 6635 4666 6684 4678
rect 6635 4646 6646 4666
rect 6666 4646 6684 4666
rect 6635 4636 6684 4646
rect 6734 4662 6778 4678
rect 6734 4642 6749 4662
rect 6769 4642 6778 4662
rect 6734 4636 6778 4642
rect 6848 4662 6892 4678
rect 6848 4642 6857 4662
rect 6877 4642 6892 4662
rect 6848 4636 6892 4642
rect 6942 4666 6991 4678
rect 6942 4646 6960 4666
rect 6980 4646 6991 4666
rect 6942 4636 6991 4646
rect 7056 4662 7100 4678
rect 7056 4642 7065 4662
rect 7085 4642 7100 4662
rect 7056 4636 7100 4642
rect 7150 4666 7199 4678
rect 7150 4646 7168 4666
rect 7188 4646 7199 4666
rect 7150 4636 7199 4646
rect 7269 4662 7313 4678
rect 7269 4642 7278 4662
rect 7298 4642 7313 4662
rect 7269 4636 7313 4642
rect 7363 4666 7412 4678
rect 7363 4646 7381 4666
rect 7401 4646 7412 4666
rect 7363 4636 7412 4646
rect 9173 4663 9222 4675
rect 9173 4643 9184 4663
rect 9204 4643 9222 4663
rect 883 4536 932 4546
rect 883 4516 894 4536
rect 914 4516 932 4536
rect 883 4504 932 4516
rect 982 4540 1026 4546
rect 982 4520 997 4540
rect 1017 4520 1026 4540
rect 982 4504 1026 4520
rect 1096 4536 1145 4546
rect 1096 4516 1107 4536
rect 1127 4516 1145 4536
rect 1096 4504 1145 4516
rect 1195 4540 1239 4546
rect 1195 4520 1210 4540
rect 1230 4520 1239 4540
rect 1195 4504 1239 4520
rect 1304 4536 1353 4546
rect 1304 4516 1315 4536
rect 1335 4516 1353 4536
rect 1304 4504 1353 4516
rect 1403 4540 1447 4546
rect 1403 4520 1418 4540
rect 1438 4520 1447 4540
rect 1403 4504 1447 4520
rect 1517 4540 1561 4546
rect 1517 4520 1526 4540
rect 1546 4520 1561 4540
rect 1517 4504 1561 4520
rect 1611 4536 1660 4546
rect 9173 4633 9222 4643
rect 9272 4659 9316 4675
rect 9272 4639 9287 4659
rect 9307 4639 9316 4659
rect 9272 4633 9316 4639
rect 9386 4659 9430 4675
rect 9386 4639 9395 4659
rect 9415 4639 9430 4659
rect 9386 4633 9430 4639
rect 9480 4663 9529 4675
rect 9480 4643 9498 4663
rect 9518 4643 9529 4663
rect 9480 4633 9529 4643
rect 9594 4659 9638 4675
rect 9594 4639 9603 4659
rect 9623 4639 9638 4659
rect 9594 4633 9638 4639
rect 9688 4663 9737 4675
rect 9688 4643 9706 4663
rect 9726 4643 9737 4663
rect 9688 4633 9737 4643
rect 9807 4659 9851 4675
rect 9807 4639 9816 4659
rect 9836 4639 9851 4659
rect 9807 4633 9851 4639
rect 9901 4663 9950 4675
rect 9901 4643 9919 4663
rect 9939 4643 9950 4663
rect 9901 4633 9950 4643
rect 1611 4516 1629 4536
rect 1649 4516 1660 4536
rect 1611 4504 1660 4516
rect 1931 4532 1980 4542
rect 1931 4512 1942 4532
rect 1962 4512 1980 4532
rect 1931 4500 1980 4512
rect 2030 4536 2074 4542
rect 2030 4516 2045 4536
rect 2065 4516 2074 4536
rect 2030 4500 2074 4516
rect 2144 4532 2193 4542
rect 2144 4512 2155 4532
rect 2175 4512 2193 4532
rect 2144 4500 2193 4512
rect 2243 4536 2287 4542
rect 2243 4516 2258 4536
rect 2278 4516 2287 4536
rect 2243 4500 2287 4516
rect 2352 4532 2401 4542
rect 2352 4512 2363 4532
rect 2383 4512 2401 4532
rect 2352 4500 2401 4512
rect 2451 4536 2495 4542
rect 2451 4516 2466 4536
rect 2486 4516 2495 4536
rect 2451 4500 2495 4516
rect 2565 4536 2609 4542
rect 2565 4516 2574 4536
rect 2594 4516 2609 4536
rect 2565 4500 2609 4516
rect 2659 4532 2708 4542
rect 2659 4512 2677 4532
rect 2697 4512 2708 4532
rect 2659 4500 2708 4512
rect 4833 4538 4882 4548
rect 4833 4518 4844 4538
rect 4864 4518 4882 4538
rect 4833 4506 4882 4518
rect 4932 4542 4976 4548
rect 4932 4522 4947 4542
rect 4967 4522 4976 4542
rect 4932 4506 4976 4522
rect 5046 4538 5095 4548
rect 5046 4518 5057 4538
rect 5077 4518 5095 4538
rect 5046 4506 5095 4518
rect 5145 4542 5189 4548
rect 5145 4522 5160 4542
rect 5180 4522 5189 4542
rect 5145 4506 5189 4522
rect 5254 4538 5303 4548
rect 5254 4518 5265 4538
rect 5285 4518 5303 4538
rect 5254 4506 5303 4518
rect 5353 4542 5397 4548
rect 5353 4522 5368 4542
rect 5388 4522 5397 4542
rect 5353 4506 5397 4522
rect 5467 4542 5511 4548
rect 5467 4522 5476 4542
rect 5496 4522 5511 4542
rect 5467 4506 5511 4522
rect 5561 4538 5610 4548
rect 5561 4518 5579 4538
rect 5599 4518 5610 4538
rect 5561 4506 5610 4518
rect 17343 4660 17392 4672
rect 17343 4640 17354 4660
rect 17374 4640 17392 4660
rect 17343 4630 17392 4640
rect 17442 4656 17486 4672
rect 17442 4636 17457 4656
rect 17477 4636 17486 4656
rect 17442 4630 17486 4636
rect 17556 4656 17600 4672
rect 17556 4636 17565 4656
rect 17585 4636 17600 4656
rect 17556 4630 17600 4636
rect 17650 4660 17699 4672
rect 17650 4640 17668 4660
rect 17688 4640 17699 4660
rect 17650 4630 17699 4640
rect 17764 4656 17808 4672
rect 17764 4636 17773 4656
rect 17793 4636 17808 4656
rect 17764 4630 17808 4636
rect 17858 4660 17907 4672
rect 17858 4640 17876 4660
rect 17896 4640 17907 4660
rect 17858 4630 17907 4640
rect 17977 4656 18021 4672
rect 17977 4636 17986 4656
rect 18006 4636 18021 4656
rect 17977 4630 18021 4636
rect 18071 4660 18120 4672
rect 18071 4640 18089 4660
rect 18109 4640 18120 4660
rect 18071 4630 18120 4640
rect 19881 4657 19930 4669
rect 19881 4637 19892 4657
rect 19912 4637 19930 4657
rect 11591 4530 11640 4540
rect 11591 4510 11602 4530
rect 11622 4510 11640 4530
rect 11591 4498 11640 4510
rect 11690 4534 11734 4540
rect 11690 4514 11705 4534
rect 11725 4514 11734 4534
rect 11690 4498 11734 4514
rect 11804 4530 11853 4540
rect 11804 4510 11815 4530
rect 11835 4510 11853 4530
rect 11804 4498 11853 4510
rect 11903 4534 11947 4540
rect 11903 4514 11918 4534
rect 11938 4514 11947 4534
rect 11903 4498 11947 4514
rect 12012 4530 12061 4540
rect 12012 4510 12023 4530
rect 12043 4510 12061 4530
rect 12012 4498 12061 4510
rect 12111 4534 12155 4540
rect 12111 4514 12126 4534
rect 12146 4514 12155 4534
rect 12111 4498 12155 4514
rect 12225 4534 12269 4540
rect 12225 4514 12234 4534
rect 12254 4514 12269 4534
rect 12225 4498 12269 4514
rect 12319 4530 12368 4540
rect 19881 4627 19930 4637
rect 19980 4653 20024 4669
rect 19980 4633 19995 4653
rect 20015 4633 20024 4653
rect 19980 4627 20024 4633
rect 20094 4653 20138 4669
rect 20094 4633 20103 4653
rect 20123 4633 20138 4653
rect 20094 4627 20138 4633
rect 20188 4657 20237 4669
rect 20188 4637 20206 4657
rect 20226 4637 20237 4657
rect 20188 4627 20237 4637
rect 20302 4653 20346 4669
rect 20302 4633 20311 4653
rect 20331 4633 20346 4653
rect 20302 4627 20346 4633
rect 20396 4657 20445 4669
rect 20396 4637 20414 4657
rect 20434 4637 20445 4657
rect 20396 4627 20445 4637
rect 20515 4653 20559 4669
rect 20515 4633 20524 4653
rect 20544 4633 20559 4653
rect 20515 4627 20559 4633
rect 20609 4657 20658 4669
rect 20609 4637 20627 4657
rect 20647 4637 20658 4657
rect 20609 4627 20658 4637
rect 12319 4510 12337 4530
rect 12357 4510 12368 4530
rect 12319 4498 12368 4510
rect 12639 4526 12688 4536
rect 12639 4506 12650 4526
rect 12670 4506 12688 4526
rect 12639 4494 12688 4506
rect 12738 4530 12782 4536
rect 12738 4510 12753 4530
rect 12773 4510 12782 4530
rect 12738 4494 12782 4510
rect 12852 4526 12901 4536
rect 12852 4506 12863 4526
rect 12883 4506 12901 4526
rect 12852 4494 12901 4506
rect 12951 4530 12995 4536
rect 12951 4510 12966 4530
rect 12986 4510 12995 4530
rect 12951 4494 12995 4510
rect 13060 4526 13109 4536
rect 13060 4506 13071 4526
rect 13091 4506 13109 4526
rect 13060 4494 13109 4506
rect 13159 4530 13203 4536
rect 13159 4510 13174 4530
rect 13194 4510 13203 4530
rect 13159 4494 13203 4510
rect 13273 4530 13317 4536
rect 13273 4510 13282 4530
rect 13302 4510 13317 4530
rect 13273 4494 13317 4510
rect 13367 4526 13416 4536
rect 13367 4506 13385 4526
rect 13405 4506 13416 4526
rect 13367 4494 13416 4506
rect 15541 4532 15590 4542
rect 15541 4512 15552 4532
rect 15572 4512 15590 4532
rect 15541 4500 15590 4512
rect 15640 4536 15684 4542
rect 15640 4516 15655 4536
rect 15675 4516 15684 4536
rect 15640 4500 15684 4516
rect 15754 4532 15803 4542
rect 15754 4512 15765 4532
rect 15785 4512 15803 4532
rect 15754 4500 15803 4512
rect 15853 4536 15897 4542
rect 15853 4516 15868 4536
rect 15888 4516 15897 4536
rect 15853 4500 15897 4516
rect 15962 4532 16011 4542
rect 15962 4512 15973 4532
rect 15993 4512 16011 4532
rect 15962 4500 16011 4512
rect 16061 4536 16105 4542
rect 16061 4516 16076 4536
rect 16096 4516 16105 4536
rect 16061 4500 16105 4516
rect 16175 4536 16219 4542
rect 16175 4516 16184 4536
rect 16204 4516 16219 4536
rect 16175 4500 16219 4516
rect 16269 4532 16318 4542
rect 16269 4512 16287 4532
rect 16307 4512 16318 4532
rect 16269 4500 16318 4512
rect 28308 4664 28357 4676
rect 28308 4644 28319 4664
rect 28339 4644 28357 4664
rect 28308 4634 28357 4644
rect 28407 4660 28451 4676
rect 28407 4640 28422 4660
rect 28442 4640 28451 4660
rect 28407 4634 28451 4640
rect 28521 4660 28565 4676
rect 28521 4640 28530 4660
rect 28550 4640 28565 4660
rect 28521 4634 28565 4640
rect 28615 4664 28664 4676
rect 28615 4644 28633 4664
rect 28653 4644 28664 4664
rect 28615 4634 28664 4644
rect 28729 4660 28773 4676
rect 28729 4640 28738 4660
rect 28758 4640 28773 4660
rect 28729 4634 28773 4640
rect 28823 4664 28872 4676
rect 28823 4644 28841 4664
rect 28861 4644 28872 4664
rect 28823 4634 28872 4644
rect 28942 4660 28986 4676
rect 28942 4640 28951 4660
rect 28971 4640 28986 4660
rect 28942 4634 28986 4640
rect 29036 4664 29085 4676
rect 29036 4644 29054 4664
rect 29074 4644 29085 4664
rect 29036 4634 29085 4644
rect 30846 4661 30895 4673
rect 30846 4641 30857 4661
rect 30877 4641 30895 4661
rect 22556 4534 22605 4544
rect 22556 4514 22567 4534
rect 22587 4514 22605 4534
rect 22556 4502 22605 4514
rect 22655 4538 22699 4544
rect 22655 4518 22670 4538
rect 22690 4518 22699 4538
rect 22655 4502 22699 4518
rect 22769 4534 22818 4544
rect 22769 4514 22780 4534
rect 22800 4514 22818 4534
rect 22769 4502 22818 4514
rect 22868 4538 22912 4544
rect 22868 4518 22883 4538
rect 22903 4518 22912 4538
rect 22868 4502 22912 4518
rect 22977 4534 23026 4544
rect 22977 4514 22988 4534
rect 23008 4514 23026 4534
rect 22977 4502 23026 4514
rect 23076 4538 23120 4544
rect 23076 4518 23091 4538
rect 23111 4518 23120 4538
rect 23076 4502 23120 4518
rect 23190 4538 23234 4544
rect 23190 4518 23199 4538
rect 23219 4518 23234 4538
rect 23190 4502 23234 4518
rect 23284 4534 23333 4544
rect 30846 4631 30895 4641
rect 30945 4657 30989 4673
rect 30945 4637 30960 4657
rect 30980 4637 30989 4657
rect 30945 4631 30989 4637
rect 31059 4657 31103 4673
rect 31059 4637 31068 4657
rect 31088 4637 31103 4657
rect 31059 4631 31103 4637
rect 31153 4661 31202 4673
rect 31153 4641 31171 4661
rect 31191 4641 31202 4661
rect 31153 4631 31202 4641
rect 31267 4657 31311 4673
rect 31267 4637 31276 4657
rect 31296 4637 31311 4657
rect 31267 4631 31311 4637
rect 31361 4661 31410 4673
rect 31361 4641 31379 4661
rect 31399 4641 31410 4661
rect 31361 4631 31410 4641
rect 31480 4657 31524 4673
rect 31480 4637 31489 4657
rect 31509 4637 31524 4657
rect 31480 4631 31524 4637
rect 31574 4661 31623 4673
rect 31574 4641 31592 4661
rect 31612 4641 31623 4661
rect 31574 4631 31623 4641
rect 23284 4514 23302 4534
rect 23322 4514 23333 4534
rect 23284 4502 23333 4514
rect 23604 4530 23653 4540
rect 23604 4510 23615 4530
rect 23635 4510 23653 4530
rect 23604 4498 23653 4510
rect 23703 4534 23747 4540
rect 23703 4514 23718 4534
rect 23738 4514 23747 4534
rect 23703 4498 23747 4514
rect 23817 4530 23866 4540
rect 23817 4510 23828 4530
rect 23848 4510 23866 4530
rect 23817 4498 23866 4510
rect 23916 4534 23960 4540
rect 23916 4514 23931 4534
rect 23951 4514 23960 4534
rect 23916 4498 23960 4514
rect 24025 4530 24074 4540
rect 24025 4510 24036 4530
rect 24056 4510 24074 4530
rect 24025 4498 24074 4510
rect 24124 4534 24168 4540
rect 24124 4514 24139 4534
rect 24159 4514 24168 4534
rect 24124 4498 24168 4514
rect 24238 4534 24282 4540
rect 24238 4514 24247 4534
rect 24267 4514 24282 4534
rect 24238 4498 24282 4514
rect 24332 4530 24381 4540
rect 24332 4510 24350 4530
rect 24370 4510 24381 4530
rect 24332 4498 24381 4510
rect 26506 4536 26555 4546
rect 26506 4516 26517 4536
rect 26537 4516 26555 4536
rect 26506 4504 26555 4516
rect 26605 4540 26649 4546
rect 26605 4520 26620 4540
rect 26640 4520 26649 4540
rect 26605 4504 26649 4520
rect 26719 4536 26768 4546
rect 26719 4516 26730 4536
rect 26750 4516 26768 4536
rect 26719 4504 26768 4516
rect 26818 4540 26862 4546
rect 26818 4520 26833 4540
rect 26853 4520 26862 4540
rect 26818 4504 26862 4520
rect 26927 4536 26976 4546
rect 26927 4516 26938 4536
rect 26958 4516 26976 4536
rect 26927 4504 26976 4516
rect 27026 4540 27070 4546
rect 27026 4520 27041 4540
rect 27061 4520 27070 4540
rect 27026 4504 27070 4520
rect 27140 4540 27184 4546
rect 27140 4520 27149 4540
rect 27169 4520 27184 4540
rect 27140 4504 27184 4520
rect 27234 4536 27283 4546
rect 27234 4516 27252 4536
rect 27272 4516 27283 4536
rect 27234 4504 27283 4516
rect 39016 4658 39065 4670
rect 39016 4638 39027 4658
rect 39047 4638 39065 4658
rect 39016 4628 39065 4638
rect 39115 4654 39159 4670
rect 39115 4634 39130 4654
rect 39150 4634 39159 4654
rect 39115 4628 39159 4634
rect 39229 4654 39273 4670
rect 39229 4634 39238 4654
rect 39258 4634 39273 4654
rect 39229 4628 39273 4634
rect 39323 4658 39372 4670
rect 39323 4638 39341 4658
rect 39361 4638 39372 4658
rect 39323 4628 39372 4638
rect 39437 4654 39481 4670
rect 39437 4634 39446 4654
rect 39466 4634 39481 4654
rect 39437 4628 39481 4634
rect 39531 4658 39580 4670
rect 39531 4638 39549 4658
rect 39569 4638 39580 4658
rect 39531 4628 39580 4638
rect 39650 4654 39694 4670
rect 39650 4634 39659 4654
rect 39679 4634 39694 4654
rect 39650 4628 39694 4634
rect 39744 4658 39793 4670
rect 39744 4638 39762 4658
rect 39782 4638 39793 4658
rect 39744 4628 39793 4638
rect 41554 4655 41603 4667
rect 41554 4635 41565 4655
rect 41585 4635 41603 4655
rect 33264 4528 33313 4538
rect 33264 4508 33275 4528
rect 33295 4508 33313 4528
rect 33264 4496 33313 4508
rect 33363 4532 33407 4538
rect 33363 4512 33378 4532
rect 33398 4512 33407 4532
rect 33363 4496 33407 4512
rect 33477 4528 33526 4538
rect 33477 4508 33488 4528
rect 33508 4508 33526 4528
rect 33477 4496 33526 4508
rect 33576 4532 33620 4538
rect 33576 4512 33591 4532
rect 33611 4512 33620 4532
rect 33576 4496 33620 4512
rect 33685 4528 33734 4538
rect 33685 4508 33696 4528
rect 33716 4508 33734 4528
rect 33685 4496 33734 4508
rect 33784 4532 33828 4538
rect 33784 4512 33799 4532
rect 33819 4512 33828 4532
rect 33784 4496 33828 4512
rect 33898 4532 33942 4538
rect 33898 4512 33907 4532
rect 33927 4512 33942 4532
rect 33898 4496 33942 4512
rect 33992 4528 34041 4538
rect 41554 4625 41603 4635
rect 41653 4651 41697 4667
rect 41653 4631 41668 4651
rect 41688 4631 41697 4651
rect 41653 4625 41697 4631
rect 41767 4651 41811 4667
rect 41767 4631 41776 4651
rect 41796 4631 41811 4651
rect 41767 4625 41811 4631
rect 41861 4655 41910 4667
rect 41861 4635 41879 4655
rect 41899 4635 41910 4655
rect 41861 4625 41910 4635
rect 41975 4651 42019 4667
rect 41975 4631 41984 4651
rect 42004 4631 42019 4651
rect 41975 4625 42019 4631
rect 42069 4655 42118 4667
rect 42069 4635 42087 4655
rect 42107 4635 42118 4655
rect 42069 4625 42118 4635
rect 42188 4651 42232 4667
rect 42188 4631 42197 4651
rect 42217 4631 42232 4651
rect 42188 4625 42232 4631
rect 42282 4655 42331 4667
rect 42282 4635 42300 4655
rect 42320 4635 42331 4655
rect 42282 4625 42331 4635
rect 33992 4508 34010 4528
rect 34030 4508 34041 4528
rect 33992 4496 34041 4508
rect 34312 4524 34361 4534
rect 34312 4504 34323 4524
rect 34343 4504 34361 4524
rect 34312 4492 34361 4504
rect 34411 4528 34455 4534
rect 34411 4508 34426 4528
rect 34446 4508 34455 4528
rect 34411 4492 34455 4508
rect 34525 4524 34574 4534
rect 34525 4504 34536 4524
rect 34556 4504 34574 4524
rect 34525 4492 34574 4504
rect 34624 4528 34668 4534
rect 34624 4508 34639 4528
rect 34659 4508 34668 4528
rect 34624 4492 34668 4508
rect 34733 4524 34782 4534
rect 34733 4504 34744 4524
rect 34764 4504 34782 4524
rect 34733 4492 34782 4504
rect 34832 4528 34876 4534
rect 34832 4508 34847 4528
rect 34867 4508 34876 4528
rect 34832 4492 34876 4508
rect 34946 4528 34990 4534
rect 34946 4508 34955 4528
rect 34975 4508 34990 4528
rect 34946 4492 34990 4508
rect 35040 4524 35089 4534
rect 35040 4504 35058 4524
rect 35078 4504 35089 4524
rect 35040 4492 35089 4504
rect 37214 4530 37263 4540
rect 37214 4510 37225 4530
rect 37245 4510 37263 4530
rect 37214 4498 37263 4510
rect 37313 4534 37357 4540
rect 37313 4514 37328 4534
rect 37348 4514 37357 4534
rect 37313 4498 37357 4514
rect 37427 4530 37476 4540
rect 37427 4510 37438 4530
rect 37458 4510 37476 4530
rect 37427 4498 37476 4510
rect 37526 4534 37570 4540
rect 37526 4514 37541 4534
rect 37561 4514 37570 4534
rect 37526 4498 37570 4514
rect 37635 4530 37684 4540
rect 37635 4510 37646 4530
rect 37666 4510 37684 4530
rect 37635 4498 37684 4510
rect 37734 4534 37778 4540
rect 37734 4514 37749 4534
rect 37769 4514 37778 4534
rect 37734 4498 37778 4514
rect 37848 4534 37892 4540
rect 37848 4514 37857 4534
rect 37877 4514 37892 4534
rect 37848 4498 37892 4514
rect 37942 4530 37991 4540
rect 37942 4510 37960 4530
rect 37980 4510 37991 4530
rect 37942 4498 37991 4510
rect 8125 3988 8174 4000
rect 8125 3968 8136 3988
rect 8156 3968 8174 3988
rect 8125 3958 8174 3968
rect 8224 3984 8268 4000
rect 8224 3964 8239 3984
rect 8259 3964 8268 3984
rect 8224 3958 8268 3964
rect 8338 3984 8382 4000
rect 8338 3964 8347 3984
rect 8367 3964 8382 3984
rect 8338 3958 8382 3964
rect 8432 3988 8481 4000
rect 8432 3968 8450 3988
rect 8470 3968 8481 3988
rect 8432 3958 8481 3968
rect 8546 3984 8590 4000
rect 8546 3964 8555 3984
rect 8575 3964 8590 3984
rect 8546 3958 8590 3964
rect 8640 3988 8689 4000
rect 8640 3968 8658 3988
rect 8678 3968 8689 3988
rect 8640 3958 8689 3968
rect 8759 3984 8803 4000
rect 8759 3964 8768 3984
rect 8788 3964 8803 3984
rect 8759 3958 8803 3964
rect 8853 3988 8902 4000
rect 8853 3968 8871 3988
rect 8891 3968 8902 3988
rect 8853 3958 8902 3968
rect 9173 3984 9222 3996
rect 9173 3964 9184 3984
rect 9204 3964 9222 3984
rect 883 3857 932 3867
rect 883 3837 894 3857
rect 914 3837 932 3857
rect 883 3825 932 3837
rect 982 3861 1026 3867
rect 982 3841 997 3861
rect 1017 3841 1026 3861
rect 982 3825 1026 3841
rect 1096 3857 1145 3867
rect 1096 3837 1107 3857
rect 1127 3837 1145 3857
rect 1096 3825 1145 3837
rect 1195 3861 1239 3867
rect 1195 3841 1210 3861
rect 1230 3841 1239 3861
rect 1195 3825 1239 3841
rect 1304 3857 1353 3867
rect 1304 3837 1315 3857
rect 1335 3837 1353 3857
rect 1304 3825 1353 3837
rect 1403 3861 1447 3867
rect 1403 3841 1418 3861
rect 1438 3841 1447 3861
rect 1403 3825 1447 3841
rect 1517 3861 1561 3867
rect 1517 3841 1526 3861
rect 1546 3841 1561 3861
rect 1517 3825 1561 3841
rect 1611 3857 1660 3867
rect 9173 3954 9222 3964
rect 9272 3980 9316 3996
rect 9272 3960 9287 3980
rect 9307 3960 9316 3980
rect 9272 3954 9316 3960
rect 9386 3980 9430 3996
rect 9386 3960 9395 3980
rect 9415 3960 9430 3980
rect 9386 3954 9430 3960
rect 9480 3984 9529 3996
rect 9480 3964 9498 3984
rect 9518 3964 9529 3984
rect 9480 3954 9529 3964
rect 9594 3980 9638 3996
rect 9594 3960 9603 3980
rect 9623 3960 9638 3980
rect 9594 3954 9638 3960
rect 9688 3984 9737 3996
rect 9688 3964 9706 3984
rect 9726 3964 9737 3984
rect 9688 3954 9737 3964
rect 9807 3980 9851 3996
rect 9807 3960 9816 3980
rect 9836 3960 9851 3980
rect 9807 3954 9851 3960
rect 9901 3984 9950 3996
rect 9901 3964 9919 3984
rect 9939 3964 9950 3984
rect 9901 3954 9950 3964
rect 1611 3837 1629 3857
rect 1649 3837 1660 3857
rect 1611 3825 1660 3837
rect 3378 3852 3427 3862
rect 3378 3832 3389 3852
rect 3409 3832 3427 3852
rect 3378 3820 3427 3832
rect 3477 3856 3521 3862
rect 3477 3836 3492 3856
rect 3512 3836 3521 3856
rect 3477 3820 3521 3836
rect 3591 3852 3640 3862
rect 3591 3832 3602 3852
rect 3622 3832 3640 3852
rect 3591 3820 3640 3832
rect 3690 3856 3734 3862
rect 3690 3836 3705 3856
rect 3725 3836 3734 3856
rect 3690 3820 3734 3836
rect 3799 3852 3848 3862
rect 3799 3832 3810 3852
rect 3830 3832 3848 3852
rect 3799 3820 3848 3832
rect 3898 3856 3942 3862
rect 3898 3836 3913 3856
rect 3933 3836 3942 3856
rect 3898 3820 3942 3836
rect 4012 3856 4056 3862
rect 4012 3836 4021 3856
rect 4041 3836 4056 3856
rect 4012 3820 4056 3836
rect 4106 3852 4155 3862
rect 4106 3832 4124 3852
rect 4144 3832 4155 3852
rect 4106 3820 4155 3832
rect 18833 3982 18882 3994
rect 18833 3962 18844 3982
rect 18864 3962 18882 3982
rect 18833 3952 18882 3962
rect 18932 3978 18976 3994
rect 18932 3958 18947 3978
rect 18967 3958 18976 3978
rect 18932 3952 18976 3958
rect 19046 3978 19090 3994
rect 19046 3958 19055 3978
rect 19075 3958 19090 3978
rect 19046 3952 19090 3958
rect 19140 3982 19189 3994
rect 19140 3962 19158 3982
rect 19178 3962 19189 3982
rect 19140 3952 19189 3962
rect 19254 3978 19298 3994
rect 19254 3958 19263 3978
rect 19283 3958 19298 3978
rect 19254 3952 19298 3958
rect 19348 3982 19397 3994
rect 19348 3962 19366 3982
rect 19386 3962 19397 3982
rect 19348 3952 19397 3962
rect 19467 3978 19511 3994
rect 19467 3958 19476 3978
rect 19496 3958 19511 3978
rect 19467 3952 19511 3958
rect 19561 3982 19610 3994
rect 19561 3962 19579 3982
rect 19599 3962 19610 3982
rect 19561 3952 19610 3962
rect 19881 3978 19930 3990
rect 19881 3958 19892 3978
rect 19912 3958 19930 3978
rect 11591 3851 11640 3861
rect 11591 3831 11602 3851
rect 11622 3831 11640 3851
rect 11591 3819 11640 3831
rect 11690 3855 11734 3861
rect 11690 3835 11705 3855
rect 11725 3835 11734 3855
rect 11690 3819 11734 3835
rect 11804 3851 11853 3861
rect 11804 3831 11815 3851
rect 11835 3831 11853 3851
rect 11804 3819 11853 3831
rect 11903 3855 11947 3861
rect 11903 3835 11918 3855
rect 11938 3835 11947 3855
rect 11903 3819 11947 3835
rect 12012 3851 12061 3861
rect 12012 3831 12023 3851
rect 12043 3831 12061 3851
rect 12012 3819 12061 3831
rect 12111 3855 12155 3861
rect 12111 3835 12126 3855
rect 12146 3835 12155 3855
rect 12111 3819 12155 3835
rect 12225 3855 12269 3861
rect 12225 3835 12234 3855
rect 12254 3835 12269 3855
rect 12225 3819 12269 3835
rect 12319 3851 12368 3861
rect 19881 3948 19930 3958
rect 19980 3974 20024 3990
rect 19980 3954 19995 3974
rect 20015 3954 20024 3974
rect 19980 3948 20024 3954
rect 20094 3974 20138 3990
rect 20094 3954 20103 3974
rect 20123 3954 20138 3974
rect 20094 3948 20138 3954
rect 20188 3978 20237 3990
rect 20188 3958 20206 3978
rect 20226 3958 20237 3978
rect 20188 3948 20237 3958
rect 20302 3974 20346 3990
rect 20302 3954 20311 3974
rect 20331 3954 20346 3974
rect 20302 3948 20346 3954
rect 20396 3978 20445 3990
rect 20396 3958 20414 3978
rect 20434 3958 20445 3978
rect 20396 3948 20445 3958
rect 20515 3974 20559 3990
rect 20515 3954 20524 3974
rect 20544 3954 20559 3974
rect 20515 3948 20559 3954
rect 20609 3978 20658 3990
rect 20609 3958 20627 3978
rect 20647 3958 20658 3978
rect 20609 3948 20658 3958
rect 12319 3831 12337 3851
rect 12357 3831 12368 3851
rect 12319 3819 12368 3831
rect 14086 3846 14135 3856
rect 14086 3826 14097 3846
rect 14117 3826 14135 3846
rect 14086 3814 14135 3826
rect 14185 3850 14229 3856
rect 14185 3830 14200 3850
rect 14220 3830 14229 3850
rect 14185 3814 14229 3830
rect 14299 3846 14348 3856
rect 14299 3826 14310 3846
rect 14330 3826 14348 3846
rect 14299 3814 14348 3826
rect 14398 3850 14442 3856
rect 14398 3830 14413 3850
rect 14433 3830 14442 3850
rect 14398 3814 14442 3830
rect 14507 3846 14556 3856
rect 14507 3826 14518 3846
rect 14538 3826 14556 3846
rect 14507 3814 14556 3826
rect 14606 3850 14650 3856
rect 14606 3830 14621 3850
rect 14641 3830 14650 3850
rect 14606 3814 14650 3830
rect 14720 3850 14764 3856
rect 14720 3830 14729 3850
rect 14749 3830 14764 3850
rect 14720 3814 14764 3830
rect 14814 3846 14863 3856
rect 14814 3826 14832 3846
rect 14852 3826 14863 3846
rect 14814 3814 14863 3826
rect 29798 3986 29847 3998
rect 29798 3966 29809 3986
rect 29829 3966 29847 3986
rect 29798 3956 29847 3966
rect 29897 3982 29941 3998
rect 29897 3962 29912 3982
rect 29932 3962 29941 3982
rect 29897 3956 29941 3962
rect 30011 3982 30055 3998
rect 30011 3962 30020 3982
rect 30040 3962 30055 3982
rect 30011 3956 30055 3962
rect 30105 3986 30154 3998
rect 30105 3966 30123 3986
rect 30143 3966 30154 3986
rect 30105 3956 30154 3966
rect 30219 3982 30263 3998
rect 30219 3962 30228 3982
rect 30248 3962 30263 3982
rect 30219 3956 30263 3962
rect 30313 3986 30362 3998
rect 30313 3966 30331 3986
rect 30351 3966 30362 3986
rect 30313 3956 30362 3966
rect 30432 3982 30476 3998
rect 30432 3962 30441 3982
rect 30461 3962 30476 3982
rect 30432 3956 30476 3962
rect 30526 3986 30575 3998
rect 30526 3966 30544 3986
rect 30564 3966 30575 3986
rect 30526 3956 30575 3966
rect 30846 3982 30895 3994
rect 30846 3962 30857 3982
rect 30877 3962 30895 3982
rect 22556 3855 22605 3865
rect 22556 3835 22567 3855
rect 22587 3835 22605 3855
rect 22556 3823 22605 3835
rect 22655 3859 22699 3865
rect 22655 3839 22670 3859
rect 22690 3839 22699 3859
rect 22655 3823 22699 3839
rect 22769 3855 22818 3865
rect 22769 3835 22780 3855
rect 22800 3835 22818 3855
rect 22769 3823 22818 3835
rect 22868 3859 22912 3865
rect 22868 3839 22883 3859
rect 22903 3839 22912 3859
rect 22868 3823 22912 3839
rect 22977 3855 23026 3865
rect 22977 3835 22988 3855
rect 23008 3835 23026 3855
rect 22977 3823 23026 3835
rect 23076 3859 23120 3865
rect 23076 3839 23091 3859
rect 23111 3839 23120 3859
rect 23076 3823 23120 3839
rect 23190 3859 23234 3865
rect 23190 3839 23199 3859
rect 23219 3839 23234 3859
rect 23190 3823 23234 3839
rect 23284 3855 23333 3865
rect 30846 3952 30895 3962
rect 30945 3978 30989 3994
rect 30945 3958 30960 3978
rect 30980 3958 30989 3978
rect 30945 3952 30989 3958
rect 31059 3978 31103 3994
rect 31059 3958 31068 3978
rect 31088 3958 31103 3978
rect 31059 3952 31103 3958
rect 31153 3982 31202 3994
rect 31153 3962 31171 3982
rect 31191 3962 31202 3982
rect 31153 3952 31202 3962
rect 31267 3978 31311 3994
rect 31267 3958 31276 3978
rect 31296 3958 31311 3978
rect 31267 3952 31311 3958
rect 31361 3982 31410 3994
rect 31361 3962 31379 3982
rect 31399 3962 31410 3982
rect 31361 3952 31410 3962
rect 31480 3978 31524 3994
rect 31480 3958 31489 3978
rect 31509 3958 31524 3978
rect 31480 3952 31524 3958
rect 31574 3982 31623 3994
rect 31574 3962 31592 3982
rect 31612 3962 31623 3982
rect 31574 3952 31623 3962
rect 23284 3835 23302 3855
rect 23322 3835 23333 3855
rect 23284 3823 23333 3835
rect 25051 3850 25100 3860
rect 25051 3830 25062 3850
rect 25082 3830 25100 3850
rect 25051 3818 25100 3830
rect 25150 3854 25194 3860
rect 25150 3834 25165 3854
rect 25185 3834 25194 3854
rect 25150 3818 25194 3834
rect 25264 3850 25313 3860
rect 25264 3830 25275 3850
rect 25295 3830 25313 3850
rect 25264 3818 25313 3830
rect 25363 3854 25407 3860
rect 25363 3834 25378 3854
rect 25398 3834 25407 3854
rect 25363 3818 25407 3834
rect 25472 3850 25521 3860
rect 25472 3830 25483 3850
rect 25503 3830 25521 3850
rect 25472 3818 25521 3830
rect 25571 3854 25615 3860
rect 25571 3834 25586 3854
rect 25606 3834 25615 3854
rect 25571 3818 25615 3834
rect 25685 3854 25729 3860
rect 25685 3834 25694 3854
rect 25714 3834 25729 3854
rect 25685 3818 25729 3834
rect 25779 3850 25828 3860
rect 25779 3830 25797 3850
rect 25817 3830 25828 3850
rect 25779 3818 25828 3830
rect 40506 3980 40555 3992
rect 40506 3960 40517 3980
rect 40537 3960 40555 3980
rect 40506 3950 40555 3960
rect 40605 3976 40649 3992
rect 40605 3956 40620 3976
rect 40640 3956 40649 3976
rect 40605 3950 40649 3956
rect 40719 3976 40763 3992
rect 40719 3956 40728 3976
rect 40748 3956 40763 3976
rect 40719 3950 40763 3956
rect 40813 3980 40862 3992
rect 40813 3960 40831 3980
rect 40851 3960 40862 3980
rect 40813 3950 40862 3960
rect 40927 3976 40971 3992
rect 40927 3956 40936 3976
rect 40956 3956 40971 3976
rect 40927 3950 40971 3956
rect 41021 3980 41070 3992
rect 41021 3960 41039 3980
rect 41059 3960 41070 3980
rect 41021 3950 41070 3960
rect 41140 3976 41184 3992
rect 41140 3956 41149 3976
rect 41169 3956 41184 3976
rect 41140 3950 41184 3956
rect 41234 3980 41283 3992
rect 41234 3960 41252 3980
rect 41272 3960 41283 3980
rect 41234 3950 41283 3960
rect 41554 3976 41603 3988
rect 41554 3956 41565 3976
rect 41585 3956 41603 3976
rect 33264 3849 33313 3859
rect 33264 3829 33275 3849
rect 33295 3829 33313 3849
rect 33264 3817 33313 3829
rect 33363 3853 33407 3859
rect 33363 3833 33378 3853
rect 33398 3833 33407 3853
rect 33363 3817 33407 3833
rect 33477 3849 33526 3859
rect 33477 3829 33488 3849
rect 33508 3829 33526 3849
rect 33477 3817 33526 3829
rect 33576 3853 33620 3859
rect 33576 3833 33591 3853
rect 33611 3833 33620 3853
rect 33576 3817 33620 3833
rect 33685 3849 33734 3859
rect 33685 3829 33696 3849
rect 33716 3829 33734 3849
rect 33685 3817 33734 3829
rect 33784 3853 33828 3859
rect 33784 3833 33799 3853
rect 33819 3833 33828 3853
rect 33784 3817 33828 3833
rect 33898 3853 33942 3859
rect 33898 3833 33907 3853
rect 33927 3833 33942 3853
rect 33898 3817 33942 3833
rect 33992 3849 34041 3859
rect 41554 3946 41603 3956
rect 41653 3972 41697 3988
rect 41653 3952 41668 3972
rect 41688 3952 41697 3972
rect 41653 3946 41697 3952
rect 41767 3972 41811 3988
rect 41767 3952 41776 3972
rect 41796 3952 41811 3972
rect 41767 3946 41811 3952
rect 41861 3976 41910 3988
rect 41861 3956 41879 3976
rect 41899 3956 41910 3976
rect 41861 3946 41910 3956
rect 41975 3972 42019 3988
rect 41975 3952 41984 3972
rect 42004 3952 42019 3972
rect 41975 3946 42019 3952
rect 42069 3976 42118 3988
rect 42069 3956 42087 3976
rect 42107 3956 42118 3976
rect 42069 3946 42118 3956
rect 42188 3972 42232 3988
rect 42188 3952 42197 3972
rect 42217 3952 42232 3972
rect 42188 3946 42232 3952
rect 42282 3976 42331 3988
rect 42282 3956 42300 3976
rect 42320 3956 42331 3976
rect 42282 3946 42331 3956
rect 33992 3829 34010 3849
rect 34030 3829 34041 3849
rect 33992 3817 34041 3829
rect 35759 3844 35808 3854
rect 35759 3824 35770 3844
rect 35790 3824 35808 3844
rect 35759 3812 35808 3824
rect 35858 3848 35902 3854
rect 35858 3828 35873 3848
rect 35893 3828 35902 3848
rect 35858 3812 35902 3828
rect 35972 3844 36021 3854
rect 35972 3824 35983 3844
rect 36003 3824 36021 3844
rect 35972 3812 36021 3824
rect 36071 3848 36115 3854
rect 36071 3828 36086 3848
rect 36106 3828 36115 3848
rect 36071 3812 36115 3828
rect 36180 3844 36229 3854
rect 36180 3824 36191 3844
rect 36211 3824 36229 3844
rect 36180 3812 36229 3824
rect 36279 3848 36323 3854
rect 36279 3828 36294 3848
rect 36314 3828 36323 3848
rect 36279 3812 36323 3828
rect 36393 3848 36437 3854
rect 36393 3828 36402 3848
rect 36422 3828 36437 3848
rect 36393 3812 36437 3828
rect 36487 3844 36536 3854
rect 36487 3824 36505 3844
rect 36525 3824 36536 3844
rect 36487 3812 36536 3824
rect 6678 3221 6727 3233
rect 6678 3201 6689 3221
rect 6709 3201 6727 3221
rect 6678 3191 6727 3201
rect 6777 3217 6821 3233
rect 6777 3197 6792 3217
rect 6812 3197 6821 3217
rect 6777 3191 6821 3197
rect 6891 3217 6935 3233
rect 6891 3197 6900 3217
rect 6920 3197 6935 3217
rect 6891 3191 6935 3197
rect 6985 3221 7034 3233
rect 6985 3201 7003 3221
rect 7023 3201 7034 3221
rect 6985 3191 7034 3201
rect 7099 3217 7143 3233
rect 7099 3197 7108 3217
rect 7128 3197 7143 3217
rect 7099 3191 7143 3197
rect 7193 3221 7242 3233
rect 7193 3201 7211 3221
rect 7231 3201 7242 3221
rect 7193 3191 7242 3201
rect 7312 3217 7356 3233
rect 7312 3197 7321 3217
rect 7341 3197 7356 3217
rect 7312 3191 7356 3197
rect 7406 3221 7455 3233
rect 7406 3201 7424 3221
rect 7444 3201 7455 3221
rect 7406 3191 7455 3201
rect 9173 3216 9222 3228
rect 9173 3196 9184 3216
rect 9204 3196 9222 3216
rect 883 3089 932 3099
rect 883 3069 894 3089
rect 914 3069 932 3089
rect 883 3057 932 3069
rect 982 3093 1026 3099
rect 982 3073 997 3093
rect 1017 3073 1026 3093
rect 982 3057 1026 3073
rect 1096 3089 1145 3099
rect 1096 3069 1107 3089
rect 1127 3069 1145 3089
rect 1096 3057 1145 3069
rect 1195 3093 1239 3099
rect 1195 3073 1210 3093
rect 1230 3073 1239 3093
rect 1195 3057 1239 3073
rect 1304 3089 1353 3099
rect 1304 3069 1315 3089
rect 1335 3069 1353 3089
rect 1304 3057 1353 3069
rect 1403 3093 1447 3099
rect 1403 3073 1418 3093
rect 1438 3073 1447 3093
rect 1403 3057 1447 3073
rect 1517 3093 1561 3099
rect 1517 3073 1526 3093
rect 1546 3073 1561 3093
rect 1517 3057 1561 3073
rect 1611 3089 1660 3099
rect 9173 3186 9222 3196
rect 9272 3212 9316 3228
rect 9272 3192 9287 3212
rect 9307 3192 9316 3212
rect 9272 3186 9316 3192
rect 9386 3212 9430 3228
rect 9386 3192 9395 3212
rect 9415 3192 9430 3212
rect 9386 3186 9430 3192
rect 9480 3216 9529 3228
rect 9480 3196 9498 3216
rect 9518 3196 9529 3216
rect 9480 3186 9529 3196
rect 9594 3212 9638 3228
rect 9594 3192 9603 3212
rect 9623 3192 9638 3212
rect 9594 3186 9638 3192
rect 9688 3216 9737 3228
rect 9688 3196 9706 3216
rect 9726 3196 9737 3216
rect 9688 3186 9737 3196
rect 9807 3212 9851 3228
rect 9807 3192 9816 3212
rect 9836 3192 9851 3212
rect 9807 3186 9851 3192
rect 9901 3216 9950 3228
rect 9901 3196 9919 3216
rect 9939 3196 9950 3216
rect 9901 3186 9950 3196
rect 1611 3069 1629 3089
rect 1649 3069 1660 3089
rect 1611 3057 1660 3069
rect 1931 3085 1980 3095
rect 1931 3065 1942 3085
rect 1962 3065 1980 3085
rect 1931 3053 1980 3065
rect 2030 3089 2074 3095
rect 2030 3069 2045 3089
rect 2065 3069 2074 3089
rect 2030 3053 2074 3069
rect 2144 3085 2193 3095
rect 2144 3065 2155 3085
rect 2175 3065 2193 3085
rect 2144 3053 2193 3065
rect 2243 3089 2287 3095
rect 2243 3069 2258 3089
rect 2278 3069 2287 3089
rect 2243 3053 2287 3069
rect 2352 3085 2401 3095
rect 2352 3065 2363 3085
rect 2383 3065 2401 3085
rect 2352 3053 2401 3065
rect 2451 3089 2495 3095
rect 2451 3069 2466 3089
rect 2486 3069 2495 3089
rect 2451 3053 2495 3069
rect 2565 3089 2609 3095
rect 2565 3069 2574 3089
rect 2594 3069 2609 3089
rect 2565 3053 2609 3069
rect 2659 3085 2708 3095
rect 2659 3065 2677 3085
rect 2697 3065 2708 3085
rect 2659 3053 2708 3065
rect 17386 3215 17435 3227
rect 17386 3195 17397 3215
rect 17417 3195 17435 3215
rect 17386 3185 17435 3195
rect 17485 3211 17529 3227
rect 17485 3191 17500 3211
rect 17520 3191 17529 3211
rect 17485 3185 17529 3191
rect 17599 3211 17643 3227
rect 17599 3191 17608 3211
rect 17628 3191 17643 3211
rect 17599 3185 17643 3191
rect 17693 3215 17742 3227
rect 17693 3195 17711 3215
rect 17731 3195 17742 3215
rect 17693 3185 17742 3195
rect 17807 3211 17851 3227
rect 17807 3191 17816 3211
rect 17836 3191 17851 3211
rect 17807 3185 17851 3191
rect 17901 3215 17950 3227
rect 17901 3195 17919 3215
rect 17939 3195 17950 3215
rect 17901 3185 17950 3195
rect 18020 3211 18064 3227
rect 18020 3191 18029 3211
rect 18049 3191 18064 3211
rect 18020 3185 18064 3191
rect 18114 3215 18163 3227
rect 18114 3195 18132 3215
rect 18152 3195 18163 3215
rect 18114 3185 18163 3195
rect 19881 3210 19930 3222
rect 19881 3190 19892 3210
rect 19912 3190 19930 3210
rect 11591 3083 11640 3093
rect 11591 3063 11602 3083
rect 11622 3063 11640 3083
rect 11591 3051 11640 3063
rect 11690 3087 11734 3093
rect 11690 3067 11705 3087
rect 11725 3067 11734 3087
rect 11690 3051 11734 3067
rect 11804 3083 11853 3093
rect 11804 3063 11815 3083
rect 11835 3063 11853 3083
rect 11804 3051 11853 3063
rect 11903 3087 11947 3093
rect 11903 3067 11918 3087
rect 11938 3067 11947 3087
rect 11903 3051 11947 3067
rect 12012 3083 12061 3093
rect 12012 3063 12023 3083
rect 12043 3063 12061 3083
rect 12012 3051 12061 3063
rect 12111 3087 12155 3093
rect 12111 3067 12126 3087
rect 12146 3067 12155 3087
rect 12111 3051 12155 3067
rect 12225 3087 12269 3093
rect 12225 3067 12234 3087
rect 12254 3067 12269 3087
rect 12225 3051 12269 3067
rect 12319 3083 12368 3093
rect 19881 3180 19930 3190
rect 19980 3206 20024 3222
rect 19980 3186 19995 3206
rect 20015 3186 20024 3206
rect 19980 3180 20024 3186
rect 20094 3206 20138 3222
rect 20094 3186 20103 3206
rect 20123 3186 20138 3206
rect 20094 3180 20138 3186
rect 20188 3210 20237 3222
rect 20188 3190 20206 3210
rect 20226 3190 20237 3210
rect 20188 3180 20237 3190
rect 20302 3206 20346 3222
rect 20302 3186 20311 3206
rect 20331 3186 20346 3206
rect 20302 3180 20346 3186
rect 20396 3210 20445 3222
rect 20396 3190 20414 3210
rect 20434 3190 20445 3210
rect 20396 3180 20445 3190
rect 20515 3206 20559 3222
rect 20515 3186 20524 3206
rect 20544 3186 20559 3206
rect 20515 3180 20559 3186
rect 20609 3210 20658 3222
rect 20609 3190 20627 3210
rect 20647 3190 20658 3210
rect 20609 3180 20658 3190
rect 12319 3063 12337 3083
rect 12357 3063 12368 3083
rect 12319 3051 12368 3063
rect 12639 3079 12688 3089
rect 12639 3059 12650 3079
rect 12670 3059 12688 3079
rect 12639 3047 12688 3059
rect 12738 3083 12782 3089
rect 12738 3063 12753 3083
rect 12773 3063 12782 3083
rect 12738 3047 12782 3063
rect 12852 3079 12901 3089
rect 12852 3059 12863 3079
rect 12883 3059 12901 3079
rect 12852 3047 12901 3059
rect 12951 3083 12995 3089
rect 12951 3063 12966 3083
rect 12986 3063 12995 3083
rect 12951 3047 12995 3063
rect 13060 3079 13109 3089
rect 13060 3059 13071 3079
rect 13091 3059 13109 3079
rect 13060 3047 13109 3059
rect 13159 3083 13203 3089
rect 13159 3063 13174 3083
rect 13194 3063 13203 3083
rect 13159 3047 13203 3063
rect 13273 3083 13317 3089
rect 13273 3063 13282 3083
rect 13302 3063 13317 3083
rect 13273 3047 13317 3063
rect 13367 3079 13416 3089
rect 13367 3059 13385 3079
rect 13405 3059 13416 3079
rect 13367 3047 13416 3059
rect 28351 3219 28400 3231
rect 28351 3199 28362 3219
rect 28382 3199 28400 3219
rect 28351 3189 28400 3199
rect 28450 3215 28494 3231
rect 28450 3195 28465 3215
rect 28485 3195 28494 3215
rect 28450 3189 28494 3195
rect 28564 3215 28608 3231
rect 28564 3195 28573 3215
rect 28593 3195 28608 3215
rect 28564 3189 28608 3195
rect 28658 3219 28707 3231
rect 28658 3199 28676 3219
rect 28696 3199 28707 3219
rect 28658 3189 28707 3199
rect 28772 3215 28816 3231
rect 28772 3195 28781 3215
rect 28801 3195 28816 3215
rect 28772 3189 28816 3195
rect 28866 3219 28915 3231
rect 28866 3199 28884 3219
rect 28904 3199 28915 3219
rect 28866 3189 28915 3199
rect 28985 3215 29029 3231
rect 28985 3195 28994 3215
rect 29014 3195 29029 3215
rect 28985 3189 29029 3195
rect 29079 3219 29128 3231
rect 29079 3199 29097 3219
rect 29117 3199 29128 3219
rect 29079 3189 29128 3199
rect 30846 3214 30895 3226
rect 30846 3194 30857 3214
rect 30877 3194 30895 3214
rect 22556 3087 22605 3097
rect 22556 3067 22567 3087
rect 22587 3067 22605 3087
rect 22556 3055 22605 3067
rect 22655 3091 22699 3097
rect 22655 3071 22670 3091
rect 22690 3071 22699 3091
rect 22655 3055 22699 3071
rect 22769 3087 22818 3097
rect 22769 3067 22780 3087
rect 22800 3067 22818 3087
rect 22769 3055 22818 3067
rect 22868 3091 22912 3097
rect 22868 3071 22883 3091
rect 22903 3071 22912 3091
rect 22868 3055 22912 3071
rect 22977 3087 23026 3097
rect 22977 3067 22988 3087
rect 23008 3067 23026 3087
rect 22977 3055 23026 3067
rect 23076 3091 23120 3097
rect 23076 3071 23091 3091
rect 23111 3071 23120 3091
rect 23076 3055 23120 3071
rect 23190 3091 23234 3097
rect 23190 3071 23199 3091
rect 23219 3071 23234 3091
rect 23190 3055 23234 3071
rect 23284 3087 23333 3097
rect 30846 3184 30895 3194
rect 30945 3210 30989 3226
rect 30945 3190 30960 3210
rect 30980 3190 30989 3210
rect 30945 3184 30989 3190
rect 31059 3210 31103 3226
rect 31059 3190 31068 3210
rect 31088 3190 31103 3210
rect 31059 3184 31103 3190
rect 31153 3214 31202 3226
rect 31153 3194 31171 3214
rect 31191 3194 31202 3214
rect 31153 3184 31202 3194
rect 31267 3210 31311 3226
rect 31267 3190 31276 3210
rect 31296 3190 31311 3210
rect 31267 3184 31311 3190
rect 31361 3214 31410 3226
rect 31361 3194 31379 3214
rect 31399 3194 31410 3214
rect 31361 3184 31410 3194
rect 31480 3210 31524 3226
rect 31480 3190 31489 3210
rect 31509 3190 31524 3210
rect 31480 3184 31524 3190
rect 31574 3214 31623 3226
rect 31574 3194 31592 3214
rect 31612 3194 31623 3214
rect 31574 3184 31623 3194
rect 23284 3067 23302 3087
rect 23322 3067 23333 3087
rect 23284 3055 23333 3067
rect 23604 3083 23653 3093
rect 23604 3063 23615 3083
rect 23635 3063 23653 3083
rect 23604 3051 23653 3063
rect 23703 3087 23747 3093
rect 23703 3067 23718 3087
rect 23738 3067 23747 3087
rect 23703 3051 23747 3067
rect 23817 3083 23866 3093
rect 23817 3063 23828 3083
rect 23848 3063 23866 3083
rect 23817 3051 23866 3063
rect 23916 3087 23960 3093
rect 23916 3067 23931 3087
rect 23951 3067 23960 3087
rect 23916 3051 23960 3067
rect 24025 3083 24074 3093
rect 24025 3063 24036 3083
rect 24056 3063 24074 3083
rect 24025 3051 24074 3063
rect 24124 3087 24168 3093
rect 24124 3067 24139 3087
rect 24159 3067 24168 3087
rect 24124 3051 24168 3067
rect 24238 3087 24282 3093
rect 24238 3067 24247 3087
rect 24267 3067 24282 3087
rect 24238 3051 24282 3067
rect 24332 3083 24381 3093
rect 24332 3063 24350 3083
rect 24370 3063 24381 3083
rect 24332 3051 24381 3063
rect 39059 3213 39108 3225
rect 39059 3193 39070 3213
rect 39090 3193 39108 3213
rect 39059 3183 39108 3193
rect 39158 3209 39202 3225
rect 39158 3189 39173 3209
rect 39193 3189 39202 3209
rect 39158 3183 39202 3189
rect 39272 3209 39316 3225
rect 39272 3189 39281 3209
rect 39301 3189 39316 3209
rect 39272 3183 39316 3189
rect 39366 3213 39415 3225
rect 39366 3193 39384 3213
rect 39404 3193 39415 3213
rect 39366 3183 39415 3193
rect 39480 3209 39524 3225
rect 39480 3189 39489 3209
rect 39509 3189 39524 3209
rect 39480 3183 39524 3189
rect 39574 3213 39623 3225
rect 39574 3193 39592 3213
rect 39612 3193 39623 3213
rect 39574 3183 39623 3193
rect 39693 3209 39737 3225
rect 39693 3189 39702 3209
rect 39722 3189 39737 3209
rect 39693 3183 39737 3189
rect 39787 3213 39836 3225
rect 39787 3193 39805 3213
rect 39825 3193 39836 3213
rect 39787 3183 39836 3193
rect 41554 3208 41603 3220
rect 41554 3188 41565 3208
rect 41585 3188 41603 3208
rect 33264 3081 33313 3091
rect 33264 3061 33275 3081
rect 33295 3061 33313 3081
rect 33264 3049 33313 3061
rect 33363 3085 33407 3091
rect 33363 3065 33378 3085
rect 33398 3065 33407 3085
rect 33363 3049 33407 3065
rect 33477 3081 33526 3091
rect 33477 3061 33488 3081
rect 33508 3061 33526 3081
rect 33477 3049 33526 3061
rect 33576 3085 33620 3091
rect 33576 3065 33591 3085
rect 33611 3065 33620 3085
rect 33576 3049 33620 3065
rect 33685 3081 33734 3091
rect 33685 3061 33696 3081
rect 33716 3061 33734 3081
rect 33685 3049 33734 3061
rect 33784 3085 33828 3091
rect 33784 3065 33799 3085
rect 33819 3065 33828 3085
rect 33784 3049 33828 3065
rect 33898 3085 33942 3091
rect 33898 3065 33907 3085
rect 33927 3065 33942 3085
rect 33898 3049 33942 3065
rect 33992 3081 34041 3091
rect 41554 3178 41603 3188
rect 41653 3204 41697 3220
rect 41653 3184 41668 3204
rect 41688 3184 41697 3204
rect 41653 3178 41697 3184
rect 41767 3204 41811 3220
rect 41767 3184 41776 3204
rect 41796 3184 41811 3204
rect 41767 3178 41811 3184
rect 41861 3208 41910 3220
rect 41861 3188 41879 3208
rect 41899 3188 41910 3208
rect 41861 3178 41910 3188
rect 41975 3204 42019 3220
rect 41975 3184 41984 3204
rect 42004 3184 42019 3204
rect 41975 3178 42019 3184
rect 42069 3208 42118 3220
rect 42069 3188 42087 3208
rect 42107 3188 42118 3208
rect 42069 3178 42118 3188
rect 42188 3204 42232 3220
rect 42188 3184 42197 3204
rect 42217 3184 42232 3204
rect 42188 3178 42232 3184
rect 42282 3208 42331 3220
rect 42282 3188 42300 3208
rect 42320 3188 42331 3208
rect 42282 3178 42331 3188
rect 33992 3061 34010 3081
rect 34030 3061 34041 3081
rect 33992 3049 34041 3061
rect 34312 3077 34361 3087
rect 34312 3057 34323 3077
rect 34343 3057 34361 3077
rect 34312 3045 34361 3057
rect 34411 3081 34455 3087
rect 34411 3061 34426 3081
rect 34446 3061 34455 3081
rect 34411 3045 34455 3061
rect 34525 3077 34574 3087
rect 34525 3057 34536 3077
rect 34556 3057 34574 3077
rect 34525 3045 34574 3057
rect 34624 3081 34668 3087
rect 34624 3061 34639 3081
rect 34659 3061 34668 3081
rect 34624 3045 34668 3061
rect 34733 3077 34782 3087
rect 34733 3057 34744 3077
rect 34764 3057 34782 3077
rect 34733 3045 34782 3057
rect 34832 3081 34876 3087
rect 34832 3061 34847 3081
rect 34867 3061 34876 3081
rect 34832 3045 34876 3061
rect 34946 3081 34990 3087
rect 34946 3061 34955 3081
rect 34975 3061 34990 3081
rect 34946 3045 34990 3061
rect 35040 3077 35089 3087
rect 35040 3057 35058 3077
rect 35078 3057 35089 3077
rect 35040 3045 35089 3057
rect 8125 2541 8174 2553
rect 8125 2521 8136 2541
rect 8156 2521 8174 2541
rect 8125 2511 8174 2521
rect 8224 2537 8268 2553
rect 8224 2517 8239 2537
rect 8259 2517 8268 2537
rect 8224 2511 8268 2517
rect 8338 2537 8382 2553
rect 8338 2517 8347 2537
rect 8367 2517 8382 2537
rect 8338 2511 8382 2517
rect 8432 2541 8481 2553
rect 8432 2521 8450 2541
rect 8470 2521 8481 2541
rect 8432 2511 8481 2521
rect 8546 2537 8590 2553
rect 8546 2517 8555 2537
rect 8575 2517 8590 2537
rect 8546 2511 8590 2517
rect 8640 2541 8689 2553
rect 8640 2521 8658 2541
rect 8678 2521 8689 2541
rect 8640 2511 8689 2521
rect 8759 2537 8803 2553
rect 8759 2517 8768 2537
rect 8788 2517 8803 2537
rect 8759 2511 8803 2517
rect 8853 2541 8902 2553
rect 8853 2521 8871 2541
rect 8891 2521 8902 2541
rect 8853 2511 8902 2521
rect 9173 2537 9222 2549
rect 9173 2517 9184 2537
rect 9204 2517 9222 2537
rect 9173 2507 9222 2517
rect 9272 2533 9316 2549
rect 9272 2513 9287 2533
rect 9307 2513 9316 2533
rect 9272 2507 9316 2513
rect 9386 2533 9430 2549
rect 9386 2513 9395 2533
rect 9415 2513 9430 2533
rect 9386 2507 9430 2513
rect 9480 2537 9529 2549
rect 9480 2517 9498 2537
rect 9518 2517 9529 2537
rect 9480 2507 9529 2517
rect 9594 2533 9638 2549
rect 9594 2513 9603 2533
rect 9623 2513 9638 2533
rect 9594 2507 9638 2513
rect 9688 2537 9737 2549
rect 9688 2517 9706 2537
rect 9726 2517 9737 2537
rect 9688 2507 9737 2517
rect 9807 2533 9851 2549
rect 9807 2513 9816 2533
rect 9836 2513 9851 2533
rect 9807 2507 9851 2513
rect 9901 2537 9950 2549
rect 9901 2517 9919 2537
rect 9939 2517 9950 2537
rect 9901 2507 9950 2517
rect 883 2410 932 2420
rect 883 2390 894 2410
rect 914 2390 932 2410
rect 883 2378 932 2390
rect 982 2414 1026 2420
rect 982 2394 997 2414
rect 1017 2394 1026 2414
rect 982 2378 1026 2394
rect 1096 2410 1145 2420
rect 1096 2390 1107 2410
rect 1127 2390 1145 2410
rect 1096 2378 1145 2390
rect 1195 2414 1239 2420
rect 1195 2394 1210 2414
rect 1230 2394 1239 2414
rect 1195 2378 1239 2394
rect 1304 2410 1353 2420
rect 1304 2390 1315 2410
rect 1335 2390 1353 2410
rect 1304 2378 1353 2390
rect 1403 2414 1447 2420
rect 1403 2394 1418 2414
rect 1438 2394 1447 2414
rect 1403 2378 1447 2394
rect 1517 2414 1561 2420
rect 1517 2394 1526 2414
rect 1546 2394 1561 2414
rect 1517 2378 1561 2394
rect 1611 2410 1660 2420
rect 1611 2390 1629 2410
rect 1649 2390 1660 2410
rect 1611 2378 1660 2390
rect 18833 2535 18882 2547
rect 18833 2515 18844 2535
rect 18864 2515 18882 2535
rect 18833 2505 18882 2515
rect 18932 2531 18976 2547
rect 18932 2511 18947 2531
rect 18967 2511 18976 2531
rect 18932 2505 18976 2511
rect 19046 2531 19090 2547
rect 19046 2511 19055 2531
rect 19075 2511 19090 2531
rect 19046 2505 19090 2511
rect 19140 2535 19189 2547
rect 19140 2515 19158 2535
rect 19178 2515 19189 2535
rect 19140 2505 19189 2515
rect 19254 2531 19298 2547
rect 19254 2511 19263 2531
rect 19283 2511 19298 2531
rect 19254 2505 19298 2511
rect 19348 2535 19397 2547
rect 19348 2515 19366 2535
rect 19386 2515 19397 2535
rect 19348 2505 19397 2515
rect 19467 2531 19511 2547
rect 19467 2511 19476 2531
rect 19496 2511 19511 2531
rect 19467 2505 19511 2511
rect 19561 2535 19610 2547
rect 19561 2515 19579 2535
rect 19599 2515 19610 2535
rect 19561 2505 19610 2515
rect 19881 2531 19930 2543
rect 19881 2511 19892 2531
rect 19912 2511 19930 2531
rect 19881 2501 19930 2511
rect 19980 2527 20024 2543
rect 19980 2507 19995 2527
rect 20015 2507 20024 2527
rect 19980 2501 20024 2507
rect 20094 2527 20138 2543
rect 20094 2507 20103 2527
rect 20123 2507 20138 2527
rect 20094 2501 20138 2507
rect 20188 2531 20237 2543
rect 20188 2511 20206 2531
rect 20226 2511 20237 2531
rect 20188 2501 20237 2511
rect 20302 2527 20346 2543
rect 20302 2507 20311 2527
rect 20331 2507 20346 2527
rect 20302 2501 20346 2507
rect 20396 2531 20445 2543
rect 20396 2511 20414 2531
rect 20434 2511 20445 2531
rect 20396 2501 20445 2511
rect 20515 2527 20559 2543
rect 20515 2507 20524 2527
rect 20544 2507 20559 2527
rect 20515 2501 20559 2507
rect 20609 2531 20658 2543
rect 20609 2511 20627 2531
rect 20647 2511 20658 2531
rect 20609 2501 20658 2511
rect 11591 2404 11640 2414
rect 11591 2384 11602 2404
rect 11622 2384 11640 2404
rect 11591 2372 11640 2384
rect 11690 2408 11734 2414
rect 11690 2388 11705 2408
rect 11725 2388 11734 2408
rect 11690 2372 11734 2388
rect 11804 2404 11853 2414
rect 11804 2384 11815 2404
rect 11835 2384 11853 2404
rect 11804 2372 11853 2384
rect 11903 2408 11947 2414
rect 11903 2388 11918 2408
rect 11938 2388 11947 2408
rect 11903 2372 11947 2388
rect 12012 2404 12061 2414
rect 12012 2384 12023 2404
rect 12043 2384 12061 2404
rect 12012 2372 12061 2384
rect 12111 2408 12155 2414
rect 12111 2388 12126 2408
rect 12146 2388 12155 2408
rect 12111 2372 12155 2388
rect 12225 2408 12269 2414
rect 12225 2388 12234 2408
rect 12254 2388 12269 2408
rect 12225 2372 12269 2388
rect 12319 2404 12368 2414
rect 12319 2384 12337 2404
rect 12357 2384 12368 2404
rect 12319 2372 12368 2384
rect 29798 2539 29847 2551
rect 29798 2519 29809 2539
rect 29829 2519 29847 2539
rect 29798 2509 29847 2519
rect 29897 2535 29941 2551
rect 29897 2515 29912 2535
rect 29932 2515 29941 2535
rect 29897 2509 29941 2515
rect 30011 2535 30055 2551
rect 30011 2515 30020 2535
rect 30040 2515 30055 2535
rect 30011 2509 30055 2515
rect 30105 2539 30154 2551
rect 30105 2519 30123 2539
rect 30143 2519 30154 2539
rect 30105 2509 30154 2519
rect 30219 2535 30263 2551
rect 30219 2515 30228 2535
rect 30248 2515 30263 2535
rect 30219 2509 30263 2515
rect 30313 2539 30362 2551
rect 30313 2519 30331 2539
rect 30351 2519 30362 2539
rect 30313 2509 30362 2519
rect 30432 2535 30476 2551
rect 30432 2515 30441 2535
rect 30461 2515 30476 2535
rect 30432 2509 30476 2515
rect 30526 2539 30575 2551
rect 30526 2519 30544 2539
rect 30564 2519 30575 2539
rect 30526 2509 30575 2519
rect 30846 2535 30895 2547
rect 30846 2515 30857 2535
rect 30877 2515 30895 2535
rect 30846 2505 30895 2515
rect 30945 2531 30989 2547
rect 30945 2511 30960 2531
rect 30980 2511 30989 2531
rect 30945 2505 30989 2511
rect 31059 2531 31103 2547
rect 31059 2511 31068 2531
rect 31088 2511 31103 2531
rect 31059 2505 31103 2511
rect 31153 2535 31202 2547
rect 31153 2515 31171 2535
rect 31191 2515 31202 2535
rect 31153 2505 31202 2515
rect 31267 2531 31311 2547
rect 31267 2511 31276 2531
rect 31296 2511 31311 2531
rect 31267 2505 31311 2511
rect 31361 2535 31410 2547
rect 31361 2515 31379 2535
rect 31399 2515 31410 2535
rect 31361 2505 31410 2515
rect 31480 2531 31524 2547
rect 31480 2511 31489 2531
rect 31509 2511 31524 2531
rect 31480 2505 31524 2511
rect 31574 2535 31623 2547
rect 31574 2515 31592 2535
rect 31612 2515 31623 2535
rect 31574 2505 31623 2515
rect 22556 2408 22605 2418
rect 22556 2388 22567 2408
rect 22587 2388 22605 2408
rect 22556 2376 22605 2388
rect 22655 2412 22699 2418
rect 22655 2392 22670 2412
rect 22690 2392 22699 2412
rect 22655 2376 22699 2392
rect 22769 2408 22818 2418
rect 22769 2388 22780 2408
rect 22800 2388 22818 2408
rect 22769 2376 22818 2388
rect 22868 2412 22912 2418
rect 22868 2392 22883 2412
rect 22903 2392 22912 2412
rect 22868 2376 22912 2392
rect 22977 2408 23026 2418
rect 22977 2388 22988 2408
rect 23008 2388 23026 2408
rect 22977 2376 23026 2388
rect 23076 2412 23120 2418
rect 23076 2392 23091 2412
rect 23111 2392 23120 2412
rect 23076 2376 23120 2392
rect 23190 2412 23234 2418
rect 23190 2392 23199 2412
rect 23219 2392 23234 2412
rect 23190 2376 23234 2392
rect 23284 2408 23333 2418
rect 23284 2388 23302 2408
rect 23322 2388 23333 2408
rect 23284 2376 23333 2388
rect 40506 2533 40555 2545
rect 40506 2513 40517 2533
rect 40537 2513 40555 2533
rect 40506 2503 40555 2513
rect 40605 2529 40649 2545
rect 40605 2509 40620 2529
rect 40640 2509 40649 2529
rect 40605 2503 40649 2509
rect 40719 2529 40763 2545
rect 40719 2509 40728 2529
rect 40748 2509 40763 2529
rect 40719 2503 40763 2509
rect 40813 2533 40862 2545
rect 40813 2513 40831 2533
rect 40851 2513 40862 2533
rect 40813 2503 40862 2513
rect 40927 2529 40971 2545
rect 40927 2509 40936 2529
rect 40956 2509 40971 2529
rect 40927 2503 40971 2509
rect 41021 2533 41070 2545
rect 41021 2513 41039 2533
rect 41059 2513 41070 2533
rect 41021 2503 41070 2513
rect 41140 2529 41184 2545
rect 41140 2509 41149 2529
rect 41169 2509 41184 2529
rect 41140 2503 41184 2509
rect 41234 2533 41283 2545
rect 41234 2513 41252 2533
rect 41272 2513 41283 2533
rect 41234 2503 41283 2513
rect 41554 2529 41603 2541
rect 41554 2509 41565 2529
rect 41585 2509 41603 2529
rect 41554 2499 41603 2509
rect 41653 2525 41697 2541
rect 41653 2505 41668 2525
rect 41688 2505 41697 2525
rect 41653 2499 41697 2505
rect 41767 2525 41811 2541
rect 41767 2505 41776 2525
rect 41796 2505 41811 2525
rect 41767 2499 41811 2505
rect 41861 2529 41910 2541
rect 41861 2509 41879 2529
rect 41899 2509 41910 2529
rect 41861 2499 41910 2509
rect 41975 2525 42019 2541
rect 41975 2505 41984 2525
rect 42004 2505 42019 2525
rect 41975 2499 42019 2505
rect 42069 2529 42118 2541
rect 42069 2509 42087 2529
rect 42107 2509 42118 2529
rect 42069 2499 42118 2509
rect 42188 2525 42232 2541
rect 42188 2505 42197 2525
rect 42217 2505 42232 2525
rect 42188 2499 42232 2505
rect 42282 2529 42331 2541
rect 42282 2509 42300 2529
rect 42320 2509 42331 2529
rect 42282 2499 42331 2509
rect 33264 2402 33313 2412
rect 33264 2382 33275 2402
rect 33295 2382 33313 2402
rect 33264 2370 33313 2382
rect 33363 2406 33407 2412
rect 33363 2386 33378 2406
rect 33398 2386 33407 2406
rect 33363 2370 33407 2386
rect 33477 2402 33526 2412
rect 33477 2382 33488 2402
rect 33508 2382 33526 2402
rect 33477 2370 33526 2382
rect 33576 2406 33620 2412
rect 33576 2386 33591 2406
rect 33611 2386 33620 2406
rect 33576 2370 33620 2386
rect 33685 2402 33734 2412
rect 33685 2382 33696 2402
rect 33716 2382 33734 2402
rect 33685 2370 33734 2382
rect 33784 2406 33828 2412
rect 33784 2386 33799 2406
rect 33819 2386 33828 2406
rect 33784 2370 33828 2386
rect 33898 2406 33942 2412
rect 33898 2386 33907 2406
rect 33927 2386 33942 2406
rect 33898 2370 33942 2386
rect 33992 2402 34041 2412
rect 33992 2382 34010 2402
rect 34030 2382 34041 2402
rect 33992 2370 34041 2382
rect 10594 251 10643 261
rect 10594 231 10605 251
rect 10625 231 10643 251
rect 10594 219 10643 231
rect 10693 255 10737 261
rect 10693 235 10708 255
rect 10728 235 10737 255
rect 10693 219 10737 235
rect 10807 251 10856 261
rect 10807 231 10818 251
rect 10838 231 10856 251
rect 10807 219 10856 231
rect 10906 255 10950 261
rect 10906 235 10921 255
rect 10941 235 10950 255
rect 10906 219 10950 235
rect 11015 251 11064 261
rect 11015 231 11026 251
rect 11046 231 11064 251
rect 11015 219 11064 231
rect 11114 255 11158 261
rect 11114 235 11129 255
rect 11149 235 11158 255
rect 11114 219 11158 235
rect 11228 255 11272 261
rect 11228 235 11237 255
rect 11257 235 11272 255
rect 11228 219 11272 235
rect 11322 251 11371 261
rect 11322 231 11340 251
rect 11360 231 11371 251
rect 32267 249 32316 259
rect 11322 219 11371 231
rect 21231 238 21280 248
rect 21231 218 21242 238
rect 21262 218 21280 238
rect 21231 206 21280 218
rect 21330 242 21374 248
rect 21330 222 21345 242
rect 21365 222 21374 242
rect 21330 206 21374 222
rect 21444 238 21493 248
rect 21444 218 21455 238
rect 21475 218 21493 238
rect 21444 206 21493 218
rect 21543 242 21587 248
rect 21543 222 21558 242
rect 21578 222 21587 242
rect 21543 206 21587 222
rect 21652 238 21701 248
rect 21652 218 21663 238
rect 21683 218 21701 238
rect 21652 206 21701 218
rect 21751 242 21795 248
rect 21751 222 21766 242
rect 21786 222 21795 242
rect 21751 206 21795 222
rect 21865 242 21909 248
rect 21865 222 21874 242
rect 21894 222 21909 242
rect 21865 206 21909 222
rect 21959 238 22008 248
rect 21959 218 21977 238
rect 21997 218 22008 238
rect 21959 206 22008 218
rect 32267 229 32278 249
rect 32298 229 32316 249
rect 32267 217 32316 229
rect 32366 253 32410 259
rect 32366 233 32381 253
rect 32401 233 32410 253
rect 32366 217 32410 233
rect 32480 249 32529 259
rect 32480 229 32491 249
rect 32511 229 32529 249
rect 32480 217 32529 229
rect 32579 253 32623 259
rect 32579 233 32594 253
rect 32614 233 32623 253
rect 32579 217 32623 233
rect 32688 249 32737 259
rect 32688 229 32699 249
rect 32719 229 32737 249
rect 32688 217 32737 229
rect 32787 253 32831 259
rect 32787 233 32802 253
rect 32822 233 32831 253
rect 32787 217 32831 233
rect 32901 253 32945 259
rect 32901 233 32910 253
rect 32930 233 32945 253
rect 32901 217 32945 233
rect 32995 249 33044 259
rect 32995 229 33013 249
rect 33033 229 33044 249
rect 32995 217 33044 229
<< pdiff >>
rect 889 13660 933 13698
rect 889 13640 901 13660
rect 921 13640 933 13660
rect 889 13598 933 13640
rect 983 13660 1025 13698
rect 983 13640 997 13660
rect 1017 13640 1025 13660
rect 983 13598 1025 13640
rect 1102 13660 1146 13698
rect 1102 13640 1114 13660
rect 1134 13640 1146 13660
rect 1102 13598 1146 13640
rect 1196 13660 1238 13698
rect 1196 13640 1210 13660
rect 1230 13640 1238 13660
rect 1196 13598 1238 13640
rect 1310 13660 1354 13698
rect 1310 13640 1322 13660
rect 1342 13640 1354 13660
rect 1310 13598 1354 13640
rect 1404 13660 1446 13698
rect 1404 13640 1418 13660
rect 1438 13640 1446 13660
rect 1404 13598 1446 13640
rect 1520 13660 1562 13698
rect 1520 13640 1528 13660
rect 1548 13640 1562 13660
rect 1520 13598 1562 13640
rect 1612 13667 1657 13698
rect 1612 13660 1656 13667
rect 1612 13640 1624 13660
rect 1644 13640 1656 13660
rect 1612 13598 1656 13640
rect 1937 13656 1981 13694
rect 1937 13636 1949 13656
rect 1969 13636 1981 13656
rect 1937 13594 1981 13636
rect 2031 13656 2073 13694
rect 2031 13636 2045 13656
rect 2065 13636 2073 13656
rect 2031 13594 2073 13636
rect 2150 13656 2194 13694
rect 2150 13636 2162 13656
rect 2182 13636 2194 13656
rect 2150 13594 2194 13636
rect 2244 13656 2286 13694
rect 2244 13636 2258 13656
rect 2278 13636 2286 13656
rect 2244 13594 2286 13636
rect 2358 13656 2402 13694
rect 2358 13636 2370 13656
rect 2390 13636 2402 13656
rect 2358 13594 2402 13636
rect 2452 13656 2494 13694
rect 2452 13636 2466 13656
rect 2486 13636 2494 13656
rect 2452 13594 2494 13636
rect 2568 13656 2610 13694
rect 2568 13636 2576 13656
rect 2596 13636 2610 13656
rect 2568 13594 2610 13636
rect 2660 13663 2705 13694
rect 2660 13656 2704 13663
rect 2660 13636 2672 13656
rect 2692 13636 2704 13656
rect 2660 13594 2704 13636
rect 11597 13654 11641 13692
rect 11597 13634 11609 13654
rect 11629 13634 11641 13654
rect 11597 13592 11641 13634
rect 11691 13654 11733 13692
rect 11691 13634 11705 13654
rect 11725 13634 11733 13654
rect 11691 13592 11733 13634
rect 11810 13654 11854 13692
rect 11810 13634 11822 13654
rect 11842 13634 11854 13654
rect 11810 13592 11854 13634
rect 11904 13654 11946 13692
rect 11904 13634 11918 13654
rect 11938 13634 11946 13654
rect 11904 13592 11946 13634
rect 12018 13654 12062 13692
rect 12018 13634 12030 13654
rect 12050 13634 12062 13654
rect 12018 13592 12062 13634
rect 12112 13654 12154 13692
rect 12112 13634 12126 13654
rect 12146 13634 12154 13654
rect 12112 13592 12154 13634
rect 12228 13654 12270 13692
rect 12228 13634 12236 13654
rect 12256 13634 12270 13654
rect 12228 13592 12270 13634
rect 12320 13661 12365 13692
rect 12320 13654 12364 13661
rect 12320 13634 12332 13654
rect 12352 13634 12364 13654
rect 12320 13592 12364 13634
rect 12645 13650 12689 13688
rect 12645 13630 12657 13650
rect 12677 13630 12689 13650
rect 9179 13489 9223 13531
rect 9179 13469 9191 13489
rect 9211 13469 9223 13489
rect 9179 13462 9223 13469
rect 9178 13431 9223 13462
rect 9273 13489 9315 13531
rect 9273 13469 9287 13489
rect 9307 13469 9315 13489
rect 9273 13431 9315 13469
rect 9389 13489 9431 13531
rect 9389 13469 9397 13489
rect 9417 13469 9431 13489
rect 9389 13431 9431 13469
rect 9481 13489 9525 13531
rect 9481 13469 9493 13489
rect 9513 13469 9525 13489
rect 9481 13431 9525 13469
rect 9597 13489 9639 13531
rect 9597 13469 9605 13489
rect 9625 13469 9639 13489
rect 9597 13431 9639 13469
rect 9689 13489 9733 13531
rect 9689 13469 9701 13489
rect 9721 13469 9733 13489
rect 9689 13431 9733 13469
rect 9810 13489 9852 13531
rect 9810 13469 9818 13489
rect 9838 13469 9852 13489
rect 9810 13431 9852 13469
rect 9902 13489 9946 13531
rect 12645 13588 12689 13630
rect 12739 13650 12781 13688
rect 12739 13630 12753 13650
rect 12773 13630 12781 13650
rect 12739 13588 12781 13630
rect 12858 13650 12902 13688
rect 12858 13630 12870 13650
rect 12890 13630 12902 13650
rect 12858 13588 12902 13630
rect 12952 13650 12994 13688
rect 12952 13630 12966 13650
rect 12986 13630 12994 13650
rect 12952 13588 12994 13630
rect 13066 13650 13110 13688
rect 13066 13630 13078 13650
rect 13098 13630 13110 13650
rect 13066 13588 13110 13630
rect 13160 13650 13202 13688
rect 13160 13630 13174 13650
rect 13194 13630 13202 13650
rect 13160 13588 13202 13630
rect 13276 13650 13318 13688
rect 13276 13630 13284 13650
rect 13304 13630 13318 13650
rect 13276 13588 13318 13630
rect 13368 13657 13413 13688
rect 13368 13650 13412 13657
rect 13368 13630 13380 13650
rect 13400 13630 13412 13650
rect 22562 13658 22606 13696
rect 13368 13588 13412 13630
rect 9902 13469 9914 13489
rect 9934 13469 9946 13489
rect 9902 13431 9946 13469
rect 22562 13638 22574 13658
rect 22594 13638 22606 13658
rect 22562 13596 22606 13638
rect 22656 13658 22698 13696
rect 22656 13638 22670 13658
rect 22690 13638 22698 13658
rect 22656 13596 22698 13638
rect 22775 13658 22819 13696
rect 22775 13638 22787 13658
rect 22807 13638 22819 13658
rect 22775 13596 22819 13638
rect 22869 13658 22911 13696
rect 22869 13638 22883 13658
rect 22903 13638 22911 13658
rect 22869 13596 22911 13638
rect 22983 13658 23027 13696
rect 22983 13638 22995 13658
rect 23015 13638 23027 13658
rect 22983 13596 23027 13638
rect 23077 13658 23119 13696
rect 23077 13638 23091 13658
rect 23111 13638 23119 13658
rect 23077 13596 23119 13638
rect 23193 13658 23235 13696
rect 23193 13638 23201 13658
rect 23221 13638 23235 13658
rect 23193 13596 23235 13638
rect 23285 13665 23330 13696
rect 23285 13658 23329 13665
rect 23285 13638 23297 13658
rect 23317 13638 23329 13658
rect 23285 13596 23329 13638
rect 23610 13654 23654 13692
rect 23610 13634 23622 13654
rect 23642 13634 23654 13654
rect 19887 13483 19931 13525
rect 19887 13463 19899 13483
rect 19919 13463 19931 13483
rect 19887 13456 19931 13463
rect 19886 13425 19931 13456
rect 19981 13483 20023 13525
rect 19981 13463 19995 13483
rect 20015 13463 20023 13483
rect 19981 13425 20023 13463
rect 20097 13483 20139 13525
rect 20097 13463 20105 13483
rect 20125 13463 20139 13483
rect 20097 13425 20139 13463
rect 20189 13483 20233 13525
rect 20189 13463 20201 13483
rect 20221 13463 20233 13483
rect 20189 13425 20233 13463
rect 20305 13483 20347 13525
rect 20305 13463 20313 13483
rect 20333 13463 20347 13483
rect 20305 13425 20347 13463
rect 20397 13483 20441 13525
rect 20397 13463 20409 13483
rect 20429 13463 20441 13483
rect 20397 13425 20441 13463
rect 20518 13483 20560 13525
rect 20518 13463 20526 13483
rect 20546 13463 20560 13483
rect 20518 13425 20560 13463
rect 20610 13483 20654 13525
rect 23610 13592 23654 13634
rect 23704 13654 23746 13692
rect 23704 13634 23718 13654
rect 23738 13634 23746 13654
rect 23704 13592 23746 13634
rect 23823 13654 23867 13692
rect 23823 13634 23835 13654
rect 23855 13634 23867 13654
rect 23823 13592 23867 13634
rect 23917 13654 23959 13692
rect 23917 13634 23931 13654
rect 23951 13634 23959 13654
rect 23917 13592 23959 13634
rect 24031 13654 24075 13692
rect 24031 13634 24043 13654
rect 24063 13634 24075 13654
rect 24031 13592 24075 13634
rect 24125 13654 24167 13692
rect 24125 13634 24139 13654
rect 24159 13634 24167 13654
rect 24125 13592 24167 13634
rect 24241 13654 24283 13692
rect 24241 13634 24249 13654
rect 24269 13634 24283 13654
rect 24241 13592 24283 13634
rect 24333 13661 24378 13692
rect 24333 13654 24377 13661
rect 24333 13634 24345 13654
rect 24365 13634 24377 13654
rect 24333 13592 24377 13634
rect 33270 13652 33314 13690
rect 20610 13463 20622 13483
rect 20642 13463 20654 13483
rect 20610 13425 20654 13463
rect 33270 13632 33282 13652
rect 33302 13632 33314 13652
rect 33270 13590 33314 13632
rect 33364 13652 33406 13690
rect 33364 13632 33378 13652
rect 33398 13632 33406 13652
rect 33364 13590 33406 13632
rect 33483 13652 33527 13690
rect 33483 13632 33495 13652
rect 33515 13632 33527 13652
rect 33483 13590 33527 13632
rect 33577 13652 33619 13690
rect 33577 13632 33591 13652
rect 33611 13632 33619 13652
rect 33577 13590 33619 13632
rect 33691 13652 33735 13690
rect 33691 13632 33703 13652
rect 33723 13632 33735 13652
rect 33691 13590 33735 13632
rect 33785 13652 33827 13690
rect 33785 13632 33799 13652
rect 33819 13632 33827 13652
rect 33785 13590 33827 13632
rect 33901 13652 33943 13690
rect 33901 13632 33909 13652
rect 33929 13632 33943 13652
rect 33901 13590 33943 13632
rect 33993 13659 34038 13690
rect 33993 13652 34037 13659
rect 33993 13632 34005 13652
rect 34025 13632 34037 13652
rect 33993 13590 34037 13632
rect 34318 13648 34362 13686
rect 34318 13628 34330 13648
rect 34350 13628 34362 13648
rect 30852 13487 30896 13529
rect 30852 13467 30864 13487
rect 30884 13467 30896 13487
rect 30852 13460 30896 13467
rect 30851 13429 30896 13460
rect 30946 13487 30988 13529
rect 30946 13467 30960 13487
rect 30980 13467 30988 13487
rect 30946 13429 30988 13467
rect 31062 13487 31104 13529
rect 31062 13467 31070 13487
rect 31090 13467 31104 13487
rect 31062 13429 31104 13467
rect 31154 13487 31198 13529
rect 31154 13467 31166 13487
rect 31186 13467 31198 13487
rect 31154 13429 31198 13467
rect 31270 13487 31312 13529
rect 31270 13467 31278 13487
rect 31298 13467 31312 13487
rect 31270 13429 31312 13467
rect 31362 13487 31406 13529
rect 31362 13467 31374 13487
rect 31394 13467 31406 13487
rect 31362 13429 31406 13467
rect 31483 13487 31525 13529
rect 31483 13467 31491 13487
rect 31511 13467 31525 13487
rect 31483 13429 31525 13467
rect 31575 13487 31619 13529
rect 34318 13586 34362 13628
rect 34412 13648 34454 13686
rect 34412 13628 34426 13648
rect 34446 13628 34454 13648
rect 34412 13586 34454 13628
rect 34531 13648 34575 13686
rect 34531 13628 34543 13648
rect 34563 13628 34575 13648
rect 34531 13586 34575 13628
rect 34625 13648 34667 13686
rect 34625 13628 34639 13648
rect 34659 13628 34667 13648
rect 34625 13586 34667 13628
rect 34739 13648 34783 13686
rect 34739 13628 34751 13648
rect 34771 13628 34783 13648
rect 34739 13586 34783 13628
rect 34833 13648 34875 13686
rect 34833 13628 34847 13648
rect 34867 13628 34875 13648
rect 34833 13586 34875 13628
rect 34949 13648 34991 13686
rect 34949 13628 34957 13648
rect 34977 13628 34991 13648
rect 34949 13586 34991 13628
rect 35041 13655 35086 13686
rect 35041 13648 35085 13655
rect 35041 13628 35053 13648
rect 35073 13628 35085 13648
rect 35041 13586 35085 13628
rect 31575 13467 31587 13487
rect 31607 13467 31619 13487
rect 31575 13429 31619 13467
rect 41560 13481 41604 13523
rect 41560 13461 41572 13481
rect 41592 13461 41604 13481
rect 41560 13454 41604 13461
rect 41559 13423 41604 13454
rect 41654 13481 41696 13523
rect 41654 13461 41668 13481
rect 41688 13461 41696 13481
rect 41654 13423 41696 13461
rect 41770 13481 41812 13523
rect 41770 13461 41778 13481
rect 41798 13461 41812 13481
rect 41770 13423 41812 13461
rect 41862 13481 41906 13523
rect 41862 13461 41874 13481
rect 41894 13461 41906 13481
rect 41862 13423 41906 13461
rect 41978 13481 42020 13523
rect 41978 13461 41986 13481
rect 42006 13461 42020 13481
rect 41978 13423 42020 13461
rect 42070 13481 42114 13523
rect 42070 13461 42082 13481
rect 42102 13461 42114 13481
rect 42070 13423 42114 13461
rect 42191 13481 42233 13523
rect 42191 13461 42199 13481
rect 42219 13461 42233 13481
rect 42191 13423 42233 13461
rect 42283 13481 42327 13523
rect 42283 13461 42295 13481
rect 42315 13461 42327 13481
rect 42283 13423 42327 13461
rect 889 12981 933 13019
rect 889 12961 901 12981
rect 921 12961 933 12981
rect 889 12919 933 12961
rect 983 12981 1025 13019
rect 983 12961 997 12981
rect 1017 12961 1025 12981
rect 983 12919 1025 12961
rect 1102 12981 1146 13019
rect 1102 12961 1114 12981
rect 1134 12961 1146 12981
rect 1102 12919 1146 12961
rect 1196 12981 1238 13019
rect 1196 12961 1210 12981
rect 1230 12961 1238 12981
rect 1196 12919 1238 12961
rect 1310 12981 1354 13019
rect 1310 12961 1322 12981
rect 1342 12961 1354 12981
rect 1310 12919 1354 12961
rect 1404 12981 1446 13019
rect 1404 12961 1418 12981
rect 1438 12961 1446 12981
rect 1404 12919 1446 12961
rect 1520 12981 1562 13019
rect 1520 12961 1528 12981
rect 1548 12961 1562 12981
rect 1520 12919 1562 12961
rect 1612 12988 1657 13019
rect 1612 12981 1656 12988
rect 1612 12961 1624 12981
rect 1644 12961 1656 12981
rect 1612 12919 1656 12961
rect 3384 12976 3428 13014
rect 3384 12956 3396 12976
rect 3416 12956 3428 12976
rect 3384 12914 3428 12956
rect 3478 12976 3520 13014
rect 3478 12956 3492 12976
rect 3512 12956 3520 12976
rect 3478 12914 3520 12956
rect 3597 12976 3641 13014
rect 3597 12956 3609 12976
rect 3629 12956 3641 12976
rect 3597 12914 3641 12956
rect 3691 12976 3733 13014
rect 3691 12956 3705 12976
rect 3725 12956 3733 12976
rect 3691 12914 3733 12956
rect 3805 12976 3849 13014
rect 3805 12956 3817 12976
rect 3837 12956 3849 12976
rect 3805 12914 3849 12956
rect 3899 12976 3941 13014
rect 3899 12956 3913 12976
rect 3933 12956 3941 12976
rect 3899 12914 3941 12956
rect 4015 12976 4057 13014
rect 4015 12956 4023 12976
rect 4043 12956 4057 12976
rect 4015 12914 4057 12956
rect 4107 12983 4152 13014
rect 4107 12976 4151 12983
rect 4107 12956 4119 12976
rect 4139 12956 4151 12976
rect 4107 12914 4151 12956
rect 11597 12975 11641 13013
rect 11597 12955 11609 12975
rect 11629 12955 11641 12975
rect 8131 12814 8175 12856
rect 8131 12794 8143 12814
rect 8163 12794 8175 12814
rect 8131 12787 8175 12794
rect 8130 12756 8175 12787
rect 8225 12814 8267 12856
rect 8225 12794 8239 12814
rect 8259 12794 8267 12814
rect 8225 12756 8267 12794
rect 8341 12814 8383 12856
rect 8341 12794 8349 12814
rect 8369 12794 8383 12814
rect 8341 12756 8383 12794
rect 8433 12814 8477 12856
rect 8433 12794 8445 12814
rect 8465 12794 8477 12814
rect 8433 12756 8477 12794
rect 8549 12814 8591 12856
rect 8549 12794 8557 12814
rect 8577 12794 8591 12814
rect 8549 12756 8591 12794
rect 8641 12814 8685 12856
rect 8641 12794 8653 12814
rect 8673 12794 8685 12814
rect 8641 12756 8685 12794
rect 8762 12814 8804 12856
rect 8762 12794 8770 12814
rect 8790 12794 8804 12814
rect 8762 12756 8804 12794
rect 8854 12814 8898 12856
rect 11597 12913 11641 12955
rect 11691 12975 11733 13013
rect 11691 12955 11705 12975
rect 11725 12955 11733 12975
rect 11691 12913 11733 12955
rect 11810 12975 11854 13013
rect 11810 12955 11822 12975
rect 11842 12955 11854 12975
rect 11810 12913 11854 12955
rect 11904 12975 11946 13013
rect 11904 12955 11918 12975
rect 11938 12955 11946 12975
rect 11904 12913 11946 12955
rect 12018 12975 12062 13013
rect 12018 12955 12030 12975
rect 12050 12955 12062 12975
rect 12018 12913 12062 12955
rect 12112 12975 12154 13013
rect 12112 12955 12126 12975
rect 12146 12955 12154 12975
rect 12112 12913 12154 12955
rect 12228 12975 12270 13013
rect 12228 12955 12236 12975
rect 12256 12955 12270 12975
rect 12228 12913 12270 12955
rect 12320 12982 12365 13013
rect 12320 12975 12364 12982
rect 12320 12955 12332 12975
rect 12352 12955 12364 12975
rect 12320 12913 12364 12955
rect 14092 12970 14136 13008
rect 14092 12950 14104 12970
rect 14124 12950 14136 12970
rect 8854 12794 8866 12814
rect 8886 12794 8898 12814
rect 8854 12756 8898 12794
rect 9179 12810 9223 12852
rect 9179 12790 9191 12810
rect 9211 12790 9223 12810
rect 9179 12783 9223 12790
rect 9178 12752 9223 12783
rect 9273 12810 9315 12852
rect 9273 12790 9287 12810
rect 9307 12790 9315 12810
rect 9273 12752 9315 12790
rect 9389 12810 9431 12852
rect 9389 12790 9397 12810
rect 9417 12790 9431 12810
rect 9389 12752 9431 12790
rect 9481 12810 9525 12852
rect 9481 12790 9493 12810
rect 9513 12790 9525 12810
rect 9481 12752 9525 12790
rect 9597 12810 9639 12852
rect 9597 12790 9605 12810
rect 9625 12790 9639 12810
rect 9597 12752 9639 12790
rect 9689 12810 9733 12852
rect 9689 12790 9701 12810
rect 9721 12790 9733 12810
rect 9689 12752 9733 12790
rect 9810 12810 9852 12852
rect 9810 12790 9818 12810
rect 9838 12790 9852 12810
rect 9810 12752 9852 12790
rect 9902 12810 9946 12852
rect 9902 12790 9914 12810
rect 9934 12790 9946 12810
rect 14092 12908 14136 12950
rect 14186 12970 14228 13008
rect 14186 12950 14200 12970
rect 14220 12950 14228 12970
rect 14186 12908 14228 12950
rect 14305 12970 14349 13008
rect 14305 12950 14317 12970
rect 14337 12950 14349 12970
rect 14305 12908 14349 12950
rect 14399 12970 14441 13008
rect 14399 12950 14413 12970
rect 14433 12950 14441 12970
rect 14399 12908 14441 12950
rect 14513 12970 14557 13008
rect 14513 12950 14525 12970
rect 14545 12950 14557 12970
rect 14513 12908 14557 12950
rect 14607 12970 14649 13008
rect 14607 12950 14621 12970
rect 14641 12950 14649 12970
rect 14607 12908 14649 12950
rect 14723 12970 14765 13008
rect 14723 12950 14731 12970
rect 14751 12950 14765 12970
rect 14723 12908 14765 12950
rect 14815 12977 14860 13008
rect 14815 12970 14859 12977
rect 14815 12950 14827 12970
rect 14847 12950 14859 12970
rect 14815 12908 14859 12950
rect 9902 12752 9946 12790
rect 22562 12979 22606 13017
rect 22562 12959 22574 12979
rect 22594 12959 22606 12979
rect 18839 12808 18883 12850
rect 18839 12788 18851 12808
rect 18871 12788 18883 12808
rect 18839 12781 18883 12788
rect 18838 12750 18883 12781
rect 18933 12808 18975 12850
rect 18933 12788 18947 12808
rect 18967 12788 18975 12808
rect 18933 12750 18975 12788
rect 19049 12808 19091 12850
rect 19049 12788 19057 12808
rect 19077 12788 19091 12808
rect 19049 12750 19091 12788
rect 19141 12808 19185 12850
rect 19141 12788 19153 12808
rect 19173 12788 19185 12808
rect 19141 12750 19185 12788
rect 19257 12808 19299 12850
rect 19257 12788 19265 12808
rect 19285 12788 19299 12808
rect 19257 12750 19299 12788
rect 19349 12808 19393 12850
rect 19349 12788 19361 12808
rect 19381 12788 19393 12808
rect 19349 12750 19393 12788
rect 19470 12808 19512 12850
rect 19470 12788 19478 12808
rect 19498 12788 19512 12808
rect 19470 12750 19512 12788
rect 19562 12808 19606 12850
rect 22562 12917 22606 12959
rect 22656 12979 22698 13017
rect 22656 12959 22670 12979
rect 22690 12959 22698 12979
rect 22656 12917 22698 12959
rect 22775 12979 22819 13017
rect 22775 12959 22787 12979
rect 22807 12959 22819 12979
rect 22775 12917 22819 12959
rect 22869 12979 22911 13017
rect 22869 12959 22883 12979
rect 22903 12959 22911 12979
rect 22869 12917 22911 12959
rect 22983 12979 23027 13017
rect 22983 12959 22995 12979
rect 23015 12959 23027 12979
rect 22983 12917 23027 12959
rect 23077 12979 23119 13017
rect 23077 12959 23091 12979
rect 23111 12959 23119 12979
rect 23077 12917 23119 12959
rect 23193 12979 23235 13017
rect 23193 12959 23201 12979
rect 23221 12959 23235 12979
rect 23193 12917 23235 12959
rect 23285 12986 23330 13017
rect 23285 12979 23329 12986
rect 23285 12959 23297 12979
rect 23317 12959 23329 12979
rect 23285 12917 23329 12959
rect 25057 12974 25101 13012
rect 25057 12954 25069 12974
rect 25089 12954 25101 12974
rect 19562 12788 19574 12808
rect 19594 12788 19606 12808
rect 19562 12750 19606 12788
rect 19887 12804 19931 12846
rect 19887 12784 19899 12804
rect 19919 12784 19931 12804
rect 19887 12777 19931 12784
rect 19886 12746 19931 12777
rect 19981 12804 20023 12846
rect 19981 12784 19995 12804
rect 20015 12784 20023 12804
rect 19981 12746 20023 12784
rect 20097 12804 20139 12846
rect 20097 12784 20105 12804
rect 20125 12784 20139 12804
rect 20097 12746 20139 12784
rect 20189 12804 20233 12846
rect 20189 12784 20201 12804
rect 20221 12784 20233 12804
rect 20189 12746 20233 12784
rect 20305 12804 20347 12846
rect 20305 12784 20313 12804
rect 20333 12784 20347 12804
rect 20305 12746 20347 12784
rect 20397 12804 20441 12846
rect 20397 12784 20409 12804
rect 20429 12784 20441 12804
rect 20397 12746 20441 12784
rect 20518 12804 20560 12846
rect 20518 12784 20526 12804
rect 20546 12784 20560 12804
rect 20518 12746 20560 12784
rect 20610 12804 20654 12846
rect 20610 12784 20622 12804
rect 20642 12784 20654 12804
rect 25057 12912 25101 12954
rect 25151 12974 25193 13012
rect 25151 12954 25165 12974
rect 25185 12954 25193 12974
rect 25151 12912 25193 12954
rect 25270 12974 25314 13012
rect 25270 12954 25282 12974
rect 25302 12954 25314 12974
rect 25270 12912 25314 12954
rect 25364 12974 25406 13012
rect 25364 12954 25378 12974
rect 25398 12954 25406 12974
rect 25364 12912 25406 12954
rect 25478 12974 25522 13012
rect 25478 12954 25490 12974
rect 25510 12954 25522 12974
rect 25478 12912 25522 12954
rect 25572 12974 25614 13012
rect 25572 12954 25586 12974
rect 25606 12954 25614 12974
rect 25572 12912 25614 12954
rect 25688 12974 25730 13012
rect 25688 12954 25696 12974
rect 25716 12954 25730 12974
rect 25688 12912 25730 12954
rect 25780 12981 25825 13012
rect 25780 12974 25824 12981
rect 25780 12954 25792 12974
rect 25812 12954 25824 12974
rect 25780 12912 25824 12954
rect 33270 12973 33314 13011
rect 33270 12953 33282 12973
rect 33302 12953 33314 12973
rect 20610 12746 20654 12784
rect 29804 12812 29848 12854
rect 29804 12792 29816 12812
rect 29836 12792 29848 12812
rect 29804 12785 29848 12792
rect 29803 12754 29848 12785
rect 29898 12812 29940 12854
rect 29898 12792 29912 12812
rect 29932 12792 29940 12812
rect 29898 12754 29940 12792
rect 30014 12812 30056 12854
rect 30014 12792 30022 12812
rect 30042 12792 30056 12812
rect 30014 12754 30056 12792
rect 30106 12812 30150 12854
rect 30106 12792 30118 12812
rect 30138 12792 30150 12812
rect 30106 12754 30150 12792
rect 30222 12812 30264 12854
rect 30222 12792 30230 12812
rect 30250 12792 30264 12812
rect 30222 12754 30264 12792
rect 30314 12812 30358 12854
rect 30314 12792 30326 12812
rect 30346 12792 30358 12812
rect 30314 12754 30358 12792
rect 30435 12812 30477 12854
rect 30435 12792 30443 12812
rect 30463 12792 30477 12812
rect 30435 12754 30477 12792
rect 30527 12812 30571 12854
rect 33270 12911 33314 12953
rect 33364 12973 33406 13011
rect 33364 12953 33378 12973
rect 33398 12953 33406 12973
rect 33364 12911 33406 12953
rect 33483 12973 33527 13011
rect 33483 12953 33495 12973
rect 33515 12953 33527 12973
rect 33483 12911 33527 12953
rect 33577 12973 33619 13011
rect 33577 12953 33591 12973
rect 33611 12953 33619 12973
rect 33577 12911 33619 12953
rect 33691 12973 33735 13011
rect 33691 12953 33703 12973
rect 33723 12953 33735 12973
rect 33691 12911 33735 12953
rect 33785 12973 33827 13011
rect 33785 12953 33799 12973
rect 33819 12953 33827 12973
rect 33785 12911 33827 12953
rect 33901 12973 33943 13011
rect 33901 12953 33909 12973
rect 33929 12953 33943 12973
rect 33901 12911 33943 12953
rect 33993 12980 34038 13011
rect 33993 12973 34037 12980
rect 33993 12953 34005 12973
rect 34025 12953 34037 12973
rect 33993 12911 34037 12953
rect 35765 12968 35809 13006
rect 35765 12948 35777 12968
rect 35797 12948 35809 12968
rect 30527 12792 30539 12812
rect 30559 12792 30571 12812
rect 30527 12754 30571 12792
rect 30852 12808 30896 12850
rect 30852 12788 30864 12808
rect 30884 12788 30896 12808
rect 30852 12781 30896 12788
rect 30851 12750 30896 12781
rect 30946 12808 30988 12850
rect 30946 12788 30960 12808
rect 30980 12788 30988 12808
rect 30946 12750 30988 12788
rect 31062 12808 31104 12850
rect 31062 12788 31070 12808
rect 31090 12788 31104 12808
rect 31062 12750 31104 12788
rect 31154 12808 31198 12850
rect 31154 12788 31166 12808
rect 31186 12788 31198 12808
rect 31154 12750 31198 12788
rect 31270 12808 31312 12850
rect 31270 12788 31278 12808
rect 31298 12788 31312 12808
rect 31270 12750 31312 12788
rect 31362 12808 31406 12850
rect 31362 12788 31374 12808
rect 31394 12788 31406 12808
rect 31362 12750 31406 12788
rect 31483 12808 31525 12850
rect 31483 12788 31491 12808
rect 31511 12788 31525 12808
rect 31483 12750 31525 12788
rect 31575 12808 31619 12850
rect 31575 12788 31587 12808
rect 31607 12788 31619 12808
rect 35765 12906 35809 12948
rect 35859 12968 35901 13006
rect 35859 12948 35873 12968
rect 35893 12948 35901 12968
rect 35859 12906 35901 12948
rect 35978 12968 36022 13006
rect 35978 12948 35990 12968
rect 36010 12948 36022 12968
rect 35978 12906 36022 12948
rect 36072 12968 36114 13006
rect 36072 12948 36086 12968
rect 36106 12948 36114 12968
rect 36072 12906 36114 12948
rect 36186 12968 36230 13006
rect 36186 12948 36198 12968
rect 36218 12948 36230 12968
rect 36186 12906 36230 12948
rect 36280 12968 36322 13006
rect 36280 12948 36294 12968
rect 36314 12948 36322 12968
rect 36280 12906 36322 12948
rect 36396 12968 36438 13006
rect 36396 12948 36404 12968
rect 36424 12948 36438 12968
rect 36396 12906 36438 12948
rect 36488 12975 36533 13006
rect 36488 12968 36532 12975
rect 36488 12948 36500 12968
rect 36520 12948 36532 12968
rect 36488 12906 36532 12948
rect 31575 12750 31619 12788
rect 40512 12806 40556 12848
rect 40512 12786 40524 12806
rect 40544 12786 40556 12806
rect 40512 12779 40556 12786
rect 40511 12748 40556 12779
rect 40606 12806 40648 12848
rect 40606 12786 40620 12806
rect 40640 12786 40648 12806
rect 40606 12748 40648 12786
rect 40722 12806 40764 12848
rect 40722 12786 40730 12806
rect 40750 12786 40764 12806
rect 40722 12748 40764 12786
rect 40814 12806 40858 12848
rect 40814 12786 40826 12806
rect 40846 12786 40858 12806
rect 40814 12748 40858 12786
rect 40930 12806 40972 12848
rect 40930 12786 40938 12806
rect 40958 12786 40972 12806
rect 40930 12748 40972 12786
rect 41022 12806 41066 12848
rect 41022 12786 41034 12806
rect 41054 12786 41066 12806
rect 41022 12748 41066 12786
rect 41143 12806 41185 12848
rect 41143 12786 41151 12806
rect 41171 12786 41185 12806
rect 41143 12748 41185 12786
rect 41235 12806 41279 12848
rect 41235 12786 41247 12806
rect 41267 12786 41279 12806
rect 41235 12748 41279 12786
rect 41560 12802 41604 12844
rect 41560 12782 41572 12802
rect 41592 12782 41604 12802
rect 41560 12775 41604 12782
rect 41559 12744 41604 12775
rect 41654 12802 41696 12844
rect 41654 12782 41668 12802
rect 41688 12782 41696 12802
rect 41654 12744 41696 12782
rect 41770 12802 41812 12844
rect 41770 12782 41778 12802
rect 41798 12782 41812 12802
rect 41770 12744 41812 12782
rect 41862 12802 41906 12844
rect 41862 12782 41874 12802
rect 41894 12782 41906 12802
rect 41862 12744 41906 12782
rect 41978 12802 42020 12844
rect 41978 12782 41986 12802
rect 42006 12782 42020 12802
rect 41978 12744 42020 12782
rect 42070 12802 42114 12844
rect 42070 12782 42082 12802
rect 42102 12782 42114 12802
rect 42070 12744 42114 12782
rect 42191 12802 42233 12844
rect 42191 12782 42199 12802
rect 42219 12782 42233 12802
rect 42191 12744 42233 12782
rect 42283 12802 42327 12844
rect 42283 12782 42295 12802
rect 42315 12782 42327 12802
rect 42283 12744 42327 12782
rect 889 12213 933 12251
rect 889 12193 901 12213
rect 921 12193 933 12213
rect 889 12151 933 12193
rect 983 12213 1025 12251
rect 983 12193 997 12213
rect 1017 12193 1025 12213
rect 983 12151 1025 12193
rect 1102 12213 1146 12251
rect 1102 12193 1114 12213
rect 1134 12193 1146 12213
rect 1102 12151 1146 12193
rect 1196 12213 1238 12251
rect 1196 12193 1210 12213
rect 1230 12193 1238 12213
rect 1196 12151 1238 12193
rect 1310 12213 1354 12251
rect 1310 12193 1322 12213
rect 1342 12193 1354 12213
rect 1310 12151 1354 12193
rect 1404 12213 1446 12251
rect 1404 12193 1418 12213
rect 1438 12193 1446 12213
rect 1404 12151 1446 12193
rect 1520 12213 1562 12251
rect 1520 12193 1528 12213
rect 1548 12193 1562 12213
rect 1520 12151 1562 12193
rect 1612 12220 1657 12251
rect 1612 12213 1656 12220
rect 1612 12193 1624 12213
rect 1644 12193 1656 12213
rect 1612 12151 1656 12193
rect 1937 12209 1981 12247
rect 1937 12189 1949 12209
rect 1969 12189 1981 12209
rect 1937 12147 1981 12189
rect 2031 12209 2073 12247
rect 2031 12189 2045 12209
rect 2065 12189 2073 12209
rect 2031 12147 2073 12189
rect 2150 12209 2194 12247
rect 2150 12189 2162 12209
rect 2182 12189 2194 12209
rect 2150 12147 2194 12189
rect 2244 12209 2286 12247
rect 2244 12189 2258 12209
rect 2278 12189 2286 12209
rect 2244 12147 2286 12189
rect 2358 12209 2402 12247
rect 2358 12189 2370 12209
rect 2390 12189 2402 12209
rect 2358 12147 2402 12189
rect 2452 12209 2494 12247
rect 2452 12189 2466 12209
rect 2486 12189 2494 12209
rect 2452 12147 2494 12189
rect 2568 12209 2610 12247
rect 2568 12189 2576 12209
rect 2596 12189 2610 12209
rect 2568 12147 2610 12189
rect 2660 12216 2705 12247
rect 2660 12209 2704 12216
rect 2660 12189 2672 12209
rect 2692 12189 2704 12209
rect 2660 12147 2704 12189
rect 11597 12207 11641 12245
rect 6684 12047 6728 12089
rect 6684 12027 6696 12047
rect 6716 12027 6728 12047
rect 6684 12020 6728 12027
rect 6683 11989 6728 12020
rect 6778 12047 6820 12089
rect 6778 12027 6792 12047
rect 6812 12027 6820 12047
rect 6778 11989 6820 12027
rect 6894 12047 6936 12089
rect 6894 12027 6902 12047
rect 6922 12027 6936 12047
rect 6894 11989 6936 12027
rect 6986 12047 7030 12089
rect 6986 12027 6998 12047
rect 7018 12027 7030 12047
rect 6986 11989 7030 12027
rect 7102 12047 7144 12089
rect 7102 12027 7110 12047
rect 7130 12027 7144 12047
rect 7102 11989 7144 12027
rect 7194 12047 7238 12089
rect 7194 12027 7206 12047
rect 7226 12027 7238 12047
rect 7194 11989 7238 12027
rect 7315 12047 7357 12089
rect 7315 12027 7323 12047
rect 7343 12027 7357 12047
rect 7315 11989 7357 12027
rect 7407 12047 7451 12089
rect 11597 12187 11609 12207
rect 11629 12187 11641 12207
rect 11597 12145 11641 12187
rect 11691 12207 11733 12245
rect 11691 12187 11705 12207
rect 11725 12187 11733 12207
rect 11691 12145 11733 12187
rect 11810 12207 11854 12245
rect 11810 12187 11822 12207
rect 11842 12187 11854 12207
rect 11810 12145 11854 12187
rect 11904 12207 11946 12245
rect 11904 12187 11918 12207
rect 11938 12187 11946 12207
rect 11904 12145 11946 12187
rect 12018 12207 12062 12245
rect 12018 12187 12030 12207
rect 12050 12187 12062 12207
rect 12018 12145 12062 12187
rect 12112 12207 12154 12245
rect 12112 12187 12126 12207
rect 12146 12187 12154 12207
rect 12112 12145 12154 12187
rect 12228 12207 12270 12245
rect 12228 12187 12236 12207
rect 12256 12187 12270 12207
rect 12228 12145 12270 12187
rect 12320 12214 12365 12245
rect 12320 12207 12364 12214
rect 12320 12187 12332 12207
rect 12352 12187 12364 12207
rect 12320 12145 12364 12187
rect 12645 12203 12689 12241
rect 12645 12183 12657 12203
rect 12677 12183 12689 12203
rect 7407 12027 7419 12047
rect 7439 12027 7451 12047
rect 7407 11989 7451 12027
rect 9179 12042 9223 12084
rect 9179 12022 9191 12042
rect 9211 12022 9223 12042
rect 9179 12015 9223 12022
rect 9178 11984 9223 12015
rect 9273 12042 9315 12084
rect 9273 12022 9287 12042
rect 9307 12022 9315 12042
rect 9273 11984 9315 12022
rect 9389 12042 9431 12084
rect 9389 12022 9397 12042
rect 9417 12022 9431 12042
rect 9389 11984 9431 12022
rect 9481 12042 9525 12084
rect 9481 12022 9493 12042
rect 9513 12022 9525 12042
rect 9481 11984 9525 12022
rect 9597 12042 9639 12084
rect 9597 12022 9605 12042
rect 9625 12022 9639 12042
rect 9597 11984 9639 12022
rect 9689 12042 9733 12084
rect 9689 12022 9701 12042
rect 9721 12022 9733 12042
rect 9689 11984 9733 12022
rect 9810 12042 9852 12084
rect 9810 12022 9818 12042
rect 9838 12022 9852 12042
rect 9810 11984 9852 12022
rect 9902 12042 9946 12084
rect 12645 12141 12689 12183
rect 12739 12203 12781 12241
rect 12739 12183 12753 12203
rect 12773 12183 12781 12203
rect 12739 12141 12781 12183
rect 12858 12203 12902 12241
rect 12858 12183 12870 12203
rect 12890 12183 12902 12203
rect 12858 12141 12902 12183
rect 12952 12203 12994 12241
rect 12952 12183 12966 12203
rect 12986 12183 12994 12203
rect 12952 12141 12994 12183
rect 13066 12203 13110 12241
rect 13066 12183 13078 12203
rect 13098 12183 13110 12203
rect 13066 12141 13110 12183
rect 13160 12203 13202 12241
rect 13160 12183 13174 12203
rect 13194 12183 13202 12203
rect 13160 12141 13202 12183
rect 13276 12203 13318 12241
rect 13276 12183 13284 12203
rect 13304 12183 13318 12203
rect 13276 12141 13318 12183
rect 13368 12210 13413 12241
rect 13368 12203 13412 12210
rect 13368 12183 13380 12203
rect 13400 12183 13412 12203
rect 13368 12141 13412 12183
rect 22562 12211 22606 12249
rect 9902 12022 9914 12042
rect 9934 12022 9946 12042
rect 9902 11984 9946 12022
rect 17392 12041 17436 12083
rect 17392 12021 17404 12041
rect 17424 12021 17436 12041
rect 17392 12014 17436 12021
rect 17391 11983 17436 12014
rect 17486 12041 17528 12083
rect 17486 12021 17500 12041
rect 17520 12021 17528 12041
rect 17486 11983 17528 12021
rect 17602 12041 17644 12083
rect 17602 12021 17610 12041
rect 17630 12021 17644 12041
rect 17602 11983 17644 12021
rect 17694 12041 17738 12083
rect 17694 12021 17706 12041
rect 17726 12021 17738 12041
rect 17694 11983 17738 12021
rect 17810 12041 17852 12083
rect 17810 12021 17818 12041
rect 17838 12021 17852 12041
rect 17810 11983 17852 12021
rect 17902 12041 17946 12083
rect 17902 12021 17914 12041
rect 17934 12021 17946 12041
rect 17902 11983 17946 12021
rect 18023 12041 18065 12083
rect 18023 12021 18031 12041
rect 18051 12021 18065 12041
rect 18023 11983 18065 12021
rect 18115 12041 18159 12083
rect 22562 12191 22574 12211
rect 22594 12191 22606 12211
rect 22562 12149 22606 12191
rect 22656 12211 22698 12249
rect 22656 12191 22670 12211
rect 22690 12191 22698 12211
rect 22656 12149 22698 12191
rect 22775 12211 22819 12249
rect 22775 12191 22787 12211
rect 22807 12191 22819 12211
rect 22775 12149 22819 12191
rect 22869 12211 22911 12249
rect 22869 12191 22883 12211
rect 22903 12191 22911 12211
rect 22869 12149 22911 12191
rect 22983 12211 23027 12249
rect 22983 12191 22995 12211
rect 23015 12191 23027 12211
rect 22983 12149 23027 12191
rect 23077 12211 23119 12249
rect 23077 12191 23091 12211
rect 23111 12191 23119 12211
rect 23077 12149 23119 12191
rect 23193 12211 23235 12249
rect 23193 12191 23201 12211
rect 23221 12191 23235 12211
rect 23193 12149 23235 12191
rect 23285 12218 23330 12249
rect 23285 12211 23329 12218
rect 23285 12191 23297 12211
rect 23317 12191 23329 12211
rect 23285 12149 23329 12191
rect 23610 12207 23654 12245
rect 23610 12187 23622 12207
rect 23642 12187 23654 12207
rect 18115 12021 18127 12041
rect 18147 12021 18159 12041
rect 18115 11983 18159 12021
rect 19887 12036 19931 12078
rect 19887 12016 19899 12036
rect 19919 12016 19931 12036
rect 19887 12009 19931 12016
rect 19886 11978 19931 12009
rect 19981 12036 20023 12078
rect 19981 12016 19995 12036
rect 20015 12016 20023 12036
rect 19981 11978 20023 12016
rect 20097 12036 20139 12078
rect 20097 12016 20105 12036
rect 20125 12016 20139 12036
rect 20097 11978 20139 12016
rect 20189 12036 20233 12078
rect 20189 12016 20201 12036
rect 20221 12016 20233 12036
rect 20189 11978 20233 12016
rect 20305 12036 20347 12078
rect 20305 12016 20313 12036
rect 20333 12016 20347 12036
rect 20305 11978 20347 12016
rect 20397 12036 20441 12078
rect 20397 12016 20409 12036
rect 20429 12016 20441 12036
rect 20397 11978 20441 12016
rect 20518 12036 20560 12078
rect 20518 12016 20526 12036
rect 20546 12016 20560 12036
rect 20518 11978 20560 12016
rect 20610 12036 20654 12078
rect 23610 12145 23654 12187
rect 23704 12207 23746 12245
rect 23704 12187 23718 12207
rect 23738 12187 23746 12207
rect 23704 12145 23746 12187
rect 23823 12207 23867 12245
rect 23823 12187 23835 12207
rect 23855 12187 23867 12207
rect 23823 12145 23867 12187
rect 23917 12207 23959 12245
rect 23917 12187 23931 12207
rect 23951 12187 23959 12207
rect 23917 12145 23959 12187
rect 24031 12207 24075 12245
rect 24031 12187 24043 12207
rect 24063 12187 24075 12207
rect 24031 12145 24075 12187
rect 24125 12207 24167 12245
rect 24125 12187 24139 12207
rect 24159 12187 24167 12207
rect 24125 12145 24167 12187
rect 24241 12207 24283 12245
rect 24241 12187 24249 12207
rect 24269 12187 24283 12207
rect 24241 12145 24283 12187
rect 24333 12214 24378 12245
rect 24333 12207 24377 12214
rect 24333 12187 24345 12207
rect 24365 12187 24377 12207
rect 24333 12145 24377 12187
rect 20610 12016 20622 12036
rect 20642 12016 20654 12036
rect 20610 11978 20654 12016
rect 33270 12205 33314 12243
rect 28357 12045 28401 12087
rect 28357 12025 28369 12045
rect 28389 12025 28401 12045
rect 28357 12018 28401 12025
rect 28356 11987 28401 12018
rect 28451 12045 28493 12087
rect 28451 12025 28465 12045
rect 28485 12025 28493 12045
rect 28451 11987 28493 12025
rect 28567 12045 28609 12087
rect 28567 12025 28575 12045
rect 28595 12025 28609 12045
rect 28567 11987 28609 12025
rect 28659 12045 28703 12087
rect 28659 12025 28671 12045
rect 28691 12025 28703 12045
rect 28659 11987 28703 12025
rect 28775 12045 28817 12087
rect 28775 12025 28783 12045
rect 28803 12025 28817 12045
rect 28775 11987 28817 12025
rect 28867 12045 28911 12087
rect 28867 12025 28879 12045
rect 28899 12025 28911 12045
rect 28867 11987 28911 12025
rect 28988 12045 29030 12087
rect 28988 12025 28996 12045
rect 29016 12025 29030 12045
rect 28988 11987 29030 12025
rect 29080 12045 29124 12087
rect 33270 12185 33282 12205
rect 33302 12185 33314 12205
rect 33270 12143 33314 12185
rect 33364 12205 33406 12243
rect 33364 12185 33378 12205
rect 33398 12185 33406 12205
rect 33364 12143 33406 12185
rect 33483 12205 33527 12243
rect 33483 12185 33495 12205
rect 33515 12185 33527 12205
rect 33483 12143 33527 12185
rect 33577 12205 33619 12243
rect 33577 12185 33591 12205
rect 33611 12185 33619 12205
rect 33577 12143 33619 12185
rect 33691 12205 33735 12243
rect 33691 12185 33703 12205
rect 33723 12185 33735 12205
rect 33691 12143 33735 12185
rect 33785 12205 33827 12243
rect 33785 12185 33799 12205
rect 33819 12185 33827 12205
rect 33785 12143 33827 12185
rect 33901 12205 33943 12243
rect 33901 12185 33909 12205
rect 33929 12185 33943 12205
rect 33901 12143 33943 12185
rect 33993 12212 34038 12243
rect 33993 12205 34037 12212
rect 33993 12185 34005 12205
rect 34025 12185 34037 12205
rect 33993 12143 34037 12185
rect 34318 12201 34362 12239
rect 34318 12181 34330 12201
rect 34350 12181 34362 12201
rect 29080 12025 29092 12045
rect 29112 12025 29124 12045
rect 29080 11987 29124 12025
rect 30852 12040 30896 12082
rect 30852 12020 30864 12040
rect 30884 12020 30896 12040
rect 30852 12013 30896 12020
rect 30851 11982 30896 12013
rect 30946 12040 30988 12082
rect 30946 12020 30960 12040
rect 30980 12020 30988 12040
rect 30946 11982 30988 12020
rect 31062 12040 31104 12082
rect 31062 12020 31070 12040
rect 31090 12020 31104 12040
rect 31062 11982 31104 12020
rect 31154 12040 31198 12082
rect 31154 12020 31166 12040
rect 31186 12020 31198 12040
rect 31154 11982 31198 12020
rect 31270 12040 31312 12082
rect 31270 12020 31278 12040
rect 31298 12020 31312 12040
rect 31270 11982 31312 12020
rect 31362 12040 31406 12082
rect 31362 12020 31374 12040
rect 31394 12020 31406 12040
rect 31362 11982 31406 12020
rect 31483 12040 31525 12082
rect 31483 12020 31491 12040
rect 31511 12020 31525 12040
rect 31483 11982 31525 12020
rect 31575 12040 31619 12082
rect 34318 12139 34362 12181
rect 34412 12201 34454 12239
rect 34412 12181 34426 12201
rect 34446 12181 34454 12201
rect 34412 12139 34454 12181
rect 34531 12201 34575 12239
rect 34531 12181 34543 12201
rect 34563 12181 34575 12201
rect 34531 12139 34575 12181
rect 34625 12201 34667 12239
rect 34625 12181 34639 12201
rect 34659 12181 34667 12201
rect 34625 12139 34667 12181
rect 34739 12201 34783 12239
rect 34739 12181 34751 12201
rect 34771 12181 34783 12201
rect 34739 12139 34783 12181
rect 34833 12201 34875 12239
rect 34833 12181 34847 12201
rect 34867 12181 34875 12201
rect 34833 12139 34875 12181
rect 34949 12201 34991 12239
rect 34949 12181 34957 12201
rect 34977 12181 34991 12201
rect 34949 12139 34991 12181
rect 35041 12208 35086 12239
rect 35041 12201 35085 12208
rect 35041 12181 35053 12201
rect 35073 12181 35085 12201
rect 35041 12139 35085 12181
rect 31575 12020 31587 12040
rect 31607 12020 31619 12040
rect 31575 11982 31619 12020
rect 39065 12039 39109 12081
rect 39065 12019 39077 12039
rect 39097 12019 39109 12039
rect 39065 12012 39109 12019
rect 39064 11981 39109 12012
rect 39159 12039 39201 12081
rect 39159 12019 39173 12039
rect 39193 12019 39201 12039
rect 39159 11981 39201 12019
rect 39275 12039 39317 12081
rect 39275 12019 39283 12039
rect 39303 12019 39317 12039
rect 39275 11981 39317 12019
rect 39367 12039 39411 12081
rect 39367 12019 39379 12039
rect 39399 12019 39411 12039
rect 39367 11981 39411 12019
rect 39483 12039 39525 12081
rect 39483 12019 39491 12039
rect 39511 12019 39525 12039
rect 39483 11981 39525 12019
rect 39575 12039 39619 12081
rect 39575 12019 39587 12039
rect 39607 12019 39619 12039
rect 39575 11981 39619 12019
rect 39696 12039 39738 12081
rect 39696 12019 39704 12039
rect 39724 12019 39738 12039
rect 39696 11981 39738 12019
rect 39788 12039 39832 12081
rect 39788 12019 39800 12039
rect 39820 12019 39832 12039
rect 39788 11981 39832 12019
rect 41560 12034 41604 12076
rect 41560 12014 41572 12034
rect 41592 12014 41604 12034
rect 41560 12007 41604 12014
rect 41559 11976 41604 12007
rect 41654 12034 41696 12076
rect 41654 12014 41668 12034
rect 41688 12014 41696 12034
rect 41654 11976 41696 12014
rect 41770 12034 41812 12076
rect 41770 12014 41778 12034
rect 41798 12014 41812 12034
rect 41770 11976 41812 12014
rect 41862 12034 41906 12076
rect 41862 12014 41874 12034
rect 41894 12014 41906 12034
rect 41862 11976 41906 12014
rect 41978 12034 42020 12076
rect 41978 12014 41986 12034
rect 42006 12014 42020 12034
rect 41978 11976 42020 12014
rect 42070 12034 42114 12076
rect 42070 12014 42082 12034
rect 42102 12014 42114 12034
rect 42070 11976 42114 12014
rect 42191 12034 42233 12076
rect 42191 12014 42199 12034
rect 42219 12014 42233 12034
rect 42191 11976 42233 12014
rect 42283 12034 42327 12076
rect 42283 12014 42295 12034
rect 42315 12014 42327 12034
rect 42283 11976 42327 12014
rect 889 11534 933 11572
rect 889 11514 901 11534
rect 921 11514 933 11534
rect 889 11472 933 11514
rect 983 11534 1025 11572
rect 983 11514 997 11534
rect 1017 11514 1025 11534
rect 983 11472 1025 11514
rect 1102 11534 1146 11572
rect 1102 11514 1114 11534
rect 1134 11514 1146 11534
rect 1102 11472 1146 11514
rect 1196 11534 1238 11572
rect 1196 11514 1210 11534
rect 1230 11514 1238 11534
rect 1196 11472 1238 11514
rect 1310 11534 1354 11572
rect 1310 11514 1322 11534
rect 1342 11514 1354 11534
rect 1310 11472 1354 11514
rect 1404 11534 1446 11572
rect 1404 11514 1418 11534
rect 1438 11514 1446 11534
rect 1404 11472 1446 11514
rect 1520 11534 1562 11572
rect 1520 11514 1528 11534
rect 1548 11514 1562 11534
rect 1520 11472 1562 11514
rect 1612 11541 1657 11572
rect 1612 11534 1656 11541
rect 1612 11514 1624 11534
rect 1644 11514 1656 11534
rect 1612 11472 1656 11514
rect 3427 11531 3471 11569
rect 3427 11511 3439 11531
rect 3459 11511 3471 11531
rect 3427 11469 3471 11511
rect 3521 11531 3563 11569
rect 3521 11511 3535 11531
rect 3555 11511 3563 11531
rect 3521 11469 3563 11511
rect 3640 11531 3684 11569
rect 3640 11511 3652 11531
rect 3672 11511 3684 11531
rect 3640 11469 3684 11511
rect 3734 11531 3776 11569
rect 3734 11511 3748 11531
rect 3768 11511 3776 11531
rect 3734 11469 3776 11511
rect 3848 11531 3892 11569
rect 3848 11511 3860 11531
rect 3880 11511 3892 11531
rect 3848 11469 3892 11511
rect 3942 11531 3984 11569
rect 3942 11511 3956 11531
rect 3976 11511 3984 11531
rect 3942 11469 3984 11511
rect 4058 11531 4100 11569
rect 4058 11511 4066 11531
rect 4086 11511 4100 11531
rect 4058 11469 4100 11511
rect 4150 11538 4195 11569
rect 4150 11531 4194 11538
rect 4150 11511 4162 11531
rect 4182 11511 4194 11531
rect 4150 11469 4194 11511
rect 11597 11528 11641 11566
rect 11597 11508 11609 11528
rect 11629 11508 11641 11528
rect 8131 11367 8175 11409
rect 8131 11347 8143 11367
rect 8163 11347 8175 11367
rect 8131 11340 8175 11347
rect 8130 11309 8175 11340
rect 8225 11367 8267 11409
rect 8225 11347 8239 11367
rect 8259 11347 8267 11367
rect 8225 11309 8267 11347
rect 8341 11367 8383 11409
rect 8341 11347 8349 11367
rect 8369 11347 8383 11367
rect 8341 11309 8383 11347
rect 8433 11367 8477 11409
rect 8433 11347 8445 11367
rect 8465 11347 8477 11367
rect 8433 11309 8477 11347
rect 8549 11367 8591 11409
rect 8549 11347 8557 11367
rect 8577 11347 8591 11367
rect 8549 11309 8591 11347
rect 8641 11367 8685 11409
rect 8641 11347 8653 11367
rect 8673 11347 8685 11367
rect 8641 11309 8685 11347
rect 8762 11367 8804 11409
rect 8762 11347 8770 11367
rect 8790 11347 8804 11367
rect 8762 11309 8804 11347
rect 8854 11367 8898 11409
rect 11597 11466 11641 11508
rect 11691 11528 11733 11566
rect 11691 11508 11705 11528
rect 11725 11508 11733 11528
rect 11691 11466 11733 11508
rect 11810 11528 11854 11566
rect 11810 11508 11822 11528
rect 11842 11508 11854 11528
rect 11810 11466 11854 11508
rect 11904 11528 11946 11566
rect 11904 11508 11918 11528
rect 11938 11508 11946 11528
rect 11904 11466 11946 11508
rect 12018 11528 12062 11566
rect 12018 11508 12030 11528
rect 12050 11508 12062 11528
rect 12018 11466 12062 11508
rect 12112 11528 12154 11566
rect 12112 11508 12126 11528
rect 12146 11508 12154 11528
rect 12112 11466 12154 11508
rect 12228 11528 12270 11566
rect 12228 11508 12236 11528
rect 12256 11508 12270 11528
rect 12228 11466 12270 11508
rect 12320 11535 12365 11566
rect 12320 11528 12364 11535
rect 12320 11508 12332 11528
rect 12352 11508 12364 11528
rect 12320 11466 12364 11508
rect 14135 11525 14179 11563
rect 14135 11505 14147 11525
rect 14167 11505 14179 11525
rect 8854 11347 8866 11367
rect 8886 11347 8898 11367
rect 8854 11309 8898 11347
rect 9179 11363 9223 11405
rect 9179 11343 9191 11363
rect 9211 11343 9223 11363
rect 9179 11336 9223 11343
rect 9178 11305 9223 11336
rect 9273 11363 9315 11405
rect 9273 11343 9287 11363
rect 9307 11343 9315 11363
rect 9273 11305 9315 11343
rect 9389 11363 9431 11405
rect 9389 11343 9397 11363
rect 9417 11343 9431 11363
rect 9389 11305 9431 11343
rect 9481 11363 9525 11405
rect 9481 11343 9493 11363
rect 9513 11343 9525 11363
rect 9481 11305 9525 11343
rect 9597 11363 9639 11405
rect 9597 11343 9605 11363
rect 9625 11343 9639 11363
rect 9597 11305 9639 11343
rect 9689 11363 9733 11405
rect 9689 11343 9701 11363
rect 9721 11343 9733 11363
rect 9689 11305 9733 11343
rect 9810 11363 9852 11405
rect 9810 11343 9818 11363
rect 9838 11343 9852 11363
rect 9810 11305 9852 11343
rect 9902 11363 9946 11405
rect 9902 11343 9914 11363
rect 9934 11343 9946 11363
rect 14135 11463 14179 11505
rect 14229 11525 14271 11563
rect 14229 11505 14243 11525
rect 14263 11505 14271 11525
rect 14229 11463 14271 11505
rect 14348 11525 14392 11563
rect 14348 11505 14360 11525
rect 14380 11505 14392 11525
rect 14348 11463 14392 11505
rect 14442 11525 14484 11563
rect 14442 11505 14456 11525
rect 14476 11505 14484 11525
rect 14442 11463 14484 11505
rect 14556 11525 14600 11563
rect 14556 11505 14568 11525
rect 14588 11505 14600 11525
rect 14556 11463 14600 11505
rect 14650 11525 14692 11563
rect 14650 11505 14664 11525
rect 14684 11505 14692 11525
rect 14650 11463 14692 11505
rect 14766 11525 14808 11563
rect 14766 11505 14774 11525
rect 14794 11505 14808 11525
rect 14766 11463 14808 11505
rect 14858 11532 14903 11563
rect 14858 11525 14902 11532
rect 14858 11505 14870 11525
rect 14890 11505 14902 11525
rect 14858 11463 14902 11505
rect 9902 11305 9946 11343
rect 22562 11532 22606 11570
rect 22562 11512 22574 11532
rect 22594 11512 22606 11532
rect 18839 11361 18883 11403
rect 18839 11341 18851 11361
rect 18871 11341 18883 11361
rect 18839 11334 18883 11341
rect 18838 11303 18883 11334
rect 18933 11361 18975 11403
rect 18933 11341 18947 11361
rect 18967 11341 18975 11361
rect 18933 11303 18975 11341
rect 19049 11361 19091 11403
rect 19049 11341 19057 11361
rect 19077 11341 19091 11361
rect 19049 11303 19091 11341
rect 19141 11361 19185 11403
rect 19141 11341 19153 11361
rect 19173 11341 19185 11361
rect 19141 11303 19185 11341
rect 19257 11361 19299 11403
rect 19257 11341 19265 11361
rect 19285 11341 19299 11361
rect 19257 11303 19299 11341
rect 19349 11361 19393 11403
rect 19349 11341 19361 11361
rect 19381 11341 19393 11361
rect 19349 11303 19393 11341
rect 19470 11361 19512 11403
rect 19470 11341 19478 11361
rect 19498 11341 19512 11361
rect 19470 11303 19512 11341
rect 19562 11361 19606 11403
rect 22562 11470 22606 11512
rect 22656 11532 22698 11570
rect 22656 11512 22670 11532
rect 22690 11512 22698 11532
rect 22656 11470 22698 11512
rect 22775 11532 22819 11570
rect 22775 11512 22787 11532
rect 22807 11512 22819 11532
rect 22775 11470 22819 11512
rect 22869 11532 22911 11570
rect 22869 11512 22883 11532
rect 22903 11512 22911 11532
rect 22869 11470 22911 11512
rect 22983 11532 23027 11570
rect 22983 11512 22995 11532
rect 23015 11512 23027 11532
rect 22983 11470 23027 11512
rect 23077 11532 23119 11570
rect 23077 11512 23091 11532
rect 23111 11512 23119 11532
rect 23077 11470 23119 11512
rect 23193 11532 23235 11570
rect 23193 11512 23201 11532
rect 23221 11512 23235 11532
rect 23193 11470 23235 11512
rect 23285 11539 23330 11570
rect 23285 11532 23329 11539
rect 23285 11512 23297 11532
rect 23317 11512 23329 11532
rect 23285 11470 23329 11512
rect 25100 11529 25144 11567
rect 25100 11509 25112 11529
rect 25132 11509 25144 11529
rect 19562 11341 19574 11361
rect 19594 11341 19606 11361
rect 19562 11303 19606 11341
rect 19887 11357 19931 11399
rect 19887 11337 19899 11357
rect 19919 11337 19931 11357
rect 19887 11330 19931 11337
rect 19886 11299 19931 11330
rect 19981 11357 20023 11399
rect 19981 11337 19995 11357
rect 20015 11337 20023 11357
rect 19981 11299 20023 11337
rect 20097 11357 20139 11399
rect 20097 11337 20105 11357
rect 20125 11337 20139 11357
rect 20097 11299 20139 11337
rect 20189 11357 20233 11399
rect 20189 11337 20201 11357
rect 20221 11337 20233 11357
rect 20189 11299 20233 11337
rect 20305 11357 20347 11399
rect 20305 11337 20313 11357
rect 20333 11337 20347 11357
rect 20305 11299 20347 11337
rect 20397 11357 20441 11399
rect 20397 11337 20409 11357
rect 20429 11337 20441 11357
rect 20397 11299 20441 11337
rect 20518 11357 20560 11399
rect 20518 11337 20526 11357
rect 20546 11337 20560 11357
rect 20518 11299 20560 11337
rect 20610 11357 20654 11399
rect 20610 11337 20622 11357
rect 20642 11337 20654 11357
rect 25100 11467 25144 11509
rect 25194 11529 25236 11567
rect 25194 11509 25208 11529
rect 25228 11509 25236 11529
rect 25194 11467 25236 11509
rect 25313 11529 25357 11567
rect 25313 11509 25325 11529
rect 25345 11509 25357 11529
rect 25313 11467 25357 11509
rect 25407 11529 25449 11567
rect 25407 11509 25421 11529
rect 25441 11509 25449 11529
rect 25407 11467 25449 11509
rect 25521 11529 25565 11567
rect 25521 11509 25533 11529
rect 25553 11509 25565 11529
rect 25521 11467 25565 11509
rect 25615 11529 25657 11567
rect 25615 11509 25629 11529
rect 25649 11509 25657 11529
rect 25615 11467 25657 11509
rect 25731 11529 25773 11567
rect 25731 11509 25739 11529
rect 25759 11509 25773 11529
rect 25731 11467 25773 11509
rect 25823 11536 25868 11567
rect 25823 11529 25867 11536
rect 25823 11509 25835 11529
rect 25855 11509 25867 11529
rect 25823 11467 25867 11509
rect 33270 11526 33314 11564
rect 33270 11506 33282 11526
rect 33302 11506 33314 11526
rect 20610 11299 20654 11337
rect 29804 11365 29848 11407
rect 29804 11345 29816 11365
rect 29836 11345 29848 11365
rect 29804 11338 29848 11345
rect 29803 11307 29848 11338
rect 29898 11365 29940 11407
rect 29898 11345 29912 11365
rect 29932 11345 29940 11365
rect 29898 11307 29940 11345
rect 30014 11365 30056 11407
rect 30014 11345 30022 11365
rect 30042 11345 30056 11365
rect 30014 11307 30056 11345
rect 30106 11365 30150 11407
rect 30106 11345 30118 11365
rect 30138 11345 30150 11365
rect 30106 11307 30150 11345
rect 30222 11365 30264 11407
rect 30222 11345 30230 11365
rect 30250 11345 30264 11365
rect 30222 11307 30264 11345
rect 30314 11365 30358 11407
rect 30314 11345 30326 11365
rect 30346 11345 30358 11365
rect 30314 11307 30358 11345
rect 30435 11365 30477 11407
rect 30435 11345 30443 11365
rect 30463 11345 30477 11365
rect 30435 11307 30477 11345
rect 30527 11365 30571 11407
rect 33270 11464 33314 11506
rect 33364 11526 33406 11564
rect 33364 11506 33378 11526
rect 33398 11506 33406 11526
rect 33364 11464 33406 11506
rect 33483 11526 33527 11564
rect 33483 11506 33495 11526
rect 33515 11506 33527 11526
rect 33483 11464 33527 11506
rect 33577 11526 33619 11564
rect 33577 11506 33591 11526
rect 33611 11506 33619 11526
rect 33577 11464 33619 11506
rect 33691 11526 33735 11564
rect 33691 11506 33703 11526
rect 33723 11506 33735 11526
rect 33691 11464 33735 11506
rect 33785 11526 33827 11564
rect 33785 11506 33799 11526
rect 33819 11506 33827 11526
rect 33785 11464 33827 11506
rect 33901 11526 33943 11564
rect 33901 11506 33909 11526
rect 33929 11506 33943 11526
rect 33901 11464 33943 11506
rect 33993 11533 34038 11564
rect 33993 11526 34037 11533
rect 33993 11506 34005 11526
rect 34025 11506 34037 11526
rect 33993 11464 34037 11506
rect 35808 11523 35852 11561
rect 35808 11503 35820 11523
rect 35840 11503 35852 11523
rect 30527 11345 30539 11365
rect 30559 11345 30571 11365
rect 30527 11307 30571 11345
rect 30852 11361 30896 11403
rect 30852 11341 30864 11361
rect 30884 11341 30896 11361
rect 30852 11334 30896 11341
rect 30851 11303 30896 11334
rect 30946 11361 30988 11403
rect 30946 11341 30960 11361
rect 30980 11341 30988 11361
rect 30946 11303 30988 11341
rect 31062 11361 31104 11403
rect 31062 11341 31070 11361
rect 31090 11341 31104 11361
rect 31062 11303 31104 11341
rect 31154 11361 31198 11403
rect 31154 11341 31166 11361
rect 31186 11341 31198 11361
rect 31154 11303 31198 11341
rect 31270 11361 31312 11403
rect 31270 11341 31278 11361
rect 31298 11341 31312 11361
rect 31270 11303 31312 11341
rect 31362 11361 31406 11403
rect 31362 11341 31374 11361
rect 31394 11341 31406 11361
rect 31362 11303 31406 11341
rect 31483 11361 31525 11403
rect 31483 11341 31491 11361
rect 31511 11341 31525 11361
rect 31483 11303 31525 11341
rect 31575 11361 31619 11403
rect 31575 11341 31587 11361
rect 31607 11341 31619 11361
rect 35808 11461 35852 11503
rect 35902 11523 35944 11561
rect 35902 11503 35916 11523
rect 35936 11503 35944 11523
rect 35902 11461 35944 11503
rect 36021 11523 36065 11561
rect 36021 11503 36033 11523
rect 36053 11503 36065 11523
rect 36021 11461 36065 11503
rect 36115 11523 36157 11561
rect 36115 11503 36129 11523
rect 36149 11503 36157 11523
rect 36115 11461 36157 11503
rect 36229 11523 36273 11561
rect 36229 11503 36241 11523
rect 36261 11503 36273 11523
rect 36229 11461 36273 11503
rect 36323 11523 36365 11561
rect 36323 11503 36337 11523
rect 36357 11503 36365 11523
rect 36323 11461 36365 11503
rect 36439 11523 36481 11561
rect 36439 11503 36447 11523
rect 36467 11503 36481 11523
rect 36439 11461 36481 11503
rect 36531 11530 36576 11561
rect 36531 11523 36575 11530
rect 36531 11503 36543 11523
rect 36563 11503 36575 11523
rect 36531 11461 36575 11503
rect 31575 11303 31619 11341
rect 40512 11359 40556 11401
rect 40512 11339 40524 11359
rect 40544 11339 40556 11359
rect 40512 11332 40556 11339
rect 40511 11301 40556 11332
rect 40606 11359 40648 11401
rect 40606 11339 40620 11359
rect 40640 11339 40648 11359
rect 40606 11301 40648 11339
rect 40722 11359 40764 11401
rect 40722 11339 40730 11359
rect 40750 11339 40764 11359
rect 40722 11301 40764 11339
rect 40814 11359 40858 11401
rect 40814 11339 40826 11359
rect 40846 11339 40858 11359
rect 40814 11301 40858 11339
rect 40930 11359 40972 11401
rect 40930 11339 40938 11359
rect 40958 11339 40972 11359
rect 40930 11301 40972 11339
rect 41022 11359 41066 11401
rect 41022 11339 41034 11359
rect 41054 11339 41066 11359
rect 41022 11301 41066 11339
rect 41143 11359 41185 11401
rect 41143 11339 41151 11359
rect 41171 11339 41185 11359
rect 41143 11301 41185 11339
rect 41235 11359 41279 11401
rect 41235 11339 41247 11359
rect 41267 11339 41279 11359
rect 41235 11301 41279 11339
rect 41560 11355 41604 11397
rect 41560 11335 41572 11355
rect 41592 11335 41604 11355
rect 41560 11328 41604 11335
rect 41559 11297 41604 11328
rect 41654 11355 41696 11397
rect 41654 11335 41668 11355
rect 41688 11335 41696 11355
rect 41654 11297 41696 11335
rect 41770 11355 41812 11397
rect 41770 11335 41778 11355
rect 41798 11335 41812 11355
rect 41770 11297 41812 11335
rect 41862 11355 41906 11397
rect 41862 11335 41874 11355
rect 41894 11335 41906 11355
rect 41862 11297 41906 11335
rect 41978 11355 42020 11397
rect 41978 11335 41986 11355
rect 42006 11335 42020 11355
rect 41978 11297 42020 11335
rect 42070 11355 42114 11397
rect 42070 11335 42082 11355
rect 42102 11335 42114 11355
rect 42070 11297 42114 11335
rect 42191 11355 42233 11397
rect 42191 11335 42199 11355
rect 42219 11335 42233 11355
rect 42191 11297 42233 11335
rect 42283 11355 42327 11397
rect 42283 11335 42295 11355
rect 42315 11335 42327 11355
rect 42283 11297 42327 11335
rect 890 10693 934 10731
rect 890 10673 902 10693
rect 922 10673 934 10693
rect 890 10631 934 10673
rect 984 10693 1026 10731
rect 984 10673 998 10693
rect 1018 10673 1026 10693
rect 984 10631 1026 10673
rect 1103 10693 1147 10731
rect 1103 10673 1115 10693
rect 1135 10673 1147 10693
rect 1103 10631 1147 10673
rect 1197 10693 1239 10731
rect 1197 10673 1211 10693
rect 1231 10673 1239 10693
rect 1197 10631 1239 10673
rect 1311 10693 1355 10731
rect 1311 10673 1323 10693
rect 1343 10673 1355 10693
rect 1311 10631 1355 10673
rect 1405 10693 1447 10731
rect 1405 10673 1419 10693
rect 1439 10673 1447 10693
rect 1405 10631 1447 10673
rect 1521 10693 1563 10731
rect 1521 10673 1529 10693
rect 1549 10673 1563 10693
rect 1521 10631 1563 10673
rect 1613 10700 1658 10731
rect 1613 10693 1657 10700
rect 1613 10673 1625 10693
rect 1645 10673 1657 10693
rect 1613 10631 1657 10673
rect 1938 10689 1982 10727
rect 1938 10669 1950 10689
rect 1970 10669 1982 10689
rect 1938 10627 1982 10669
rect 2032 10689 2074 10727
rect 2032 10669 2046 10689
rect 2066 10669 2074 10689
rect 2032 10627 2074 10669
rect 2151 10689 2195 10727
rect 2151 10669 2163 10689
rect 2183 10669 2195 10689
rect 2151 10627 2195 10669
rect 2245 10689 2287 10727
rect 2245 10669 2259 10689
rect 2279 10669 2287 10689
rect 2245 10627 2287 10669
rect 2359 10689 2403 10727
rect 2359 10669 2371 10689
rect 2391 10669 2403 10689
rect 2359 10627 2403 10669
rect 2453 10689 2495 10727
rect 2453 10669 2467 10689
rect 2487 10669 2495 10689
rect 2453 10627 2495 10669
rect 2569 10689 2611 10727
rect 2569 10669 2577 10689
rect 2597 10669 2611 10689
rect 2569 10627 2611 10669
rect 2661 10696 2706 10727
rect 2661 10689 2705 10696
rect 2661 10669 2673 10689
rect 2693 10669 2705 10689
rect 2661 10627 2705 10669
rect 11598 10687 11642 10725
rect 6642 10525 6686 10567
rect 6642 10505 6654 10525
rect 6674 10505 6686 10525
rect 6642 10498 6686 10505
rect 6641 10467 6686 10498
rect 6736 10525 6778 10567
rect 6736 10505 6750 10525
rect 6770 10505 6778 10525
rect 6736 10467 6778 10505
rect 6852 10525 6894 10567
rect 6852 10505 6860 10525
rect 6880 10505 6894 10525
rect 6852 10467 6894 10505
rect 6944 10525 6988 10567
rect 6944 10505 6956 10525
rect 6976 10505 6988 10525
rect 6944 10467 6988 10505
rect 7060 10525 7102 10567
rect 7060 10505 7068 10525
rect 7088 10505 7102 10525
rect 7060 10467 7102 10505
rect 7152 10525 7196 10567
rect 7152 10505 7164 10525
rect 7184 10505 7196 10525
rect 7152 10467 7196 10505
rect 7273 10525 7315 10567
rect 7273 10505 7281 10525
rect 7301 10505 7315 10525
rect 7273 10467 7315 10505
rect 7365 10525 7409 10567
rect 11598 10667 11610 10687
rect 11630 10667 11642 10687
rect 11598 10625 11642 10667
rect 11692 10687 11734 10725
rect 11692 10667 11706 10687
rect 11726 10667 11734 10687
rect 11692 10625 11734 10667
rect 11811 10687 11855 10725
rect 11811 10667 11823 10687
rect 11843 10667 11855 10687
rect 11811 10625 11855 10667
rect 11905 10687 11947 10725
rect 11905 10667 11919 10687
rect 11939 10667 11947 10687
rect 11905 10625 11947 10667
rect 12019 10687 12063 10725
rect 12019 10667 12031 10687
rect 12051 10667 12063 10687
rect 12019 10625 12063 10667
rect 12113 10687 12155 10725
rect 12113 10667 12127 10687
rect 12147 10667 12155 10687
rect 12113 10625 12155 10667
rect 12229 10687 12271 10725
rect 12229 10667 12237 10687
rect 12257 10667 12271 10687
rect 12229 10625 12271 10667
rect 12321 10694 12366 10725
rect 12321 10687 12365 10694
rect 12321 10667 12333 10687
rect 12353 10667 12365 10687
rect 12321 10625 12365 10667
rect 12646 10683 12690 10721
rect 12646 10663 12658 10683
rect 12678 10663 12690 10683
rect 7365 10505 7377 10525
rect 7397 10505 7409 10525
rect 7365 10467 7409 10505
rect 9180 10522 9224 10564
rect 9180 10502 9192 10522
rect 9212 10502 9224 10522
rect 9180 10495 9224 10502
rect 9179 10464 9224 10495
rect 9274 10522 9316 10564
rect 9274 10502 9288 10522
rect 9308 10502 9316 10522
rect 9274 10464 9316 10502
rect 9390 10522 9432 10564
rect 9390 10502 9398 10522
rect 9418 10502 9432 10522
rect 9390 10464 9432 10502
rect 9482 10522 9526 10564
rect 9482 10502 9494 10522
rect 9514 10502 9526 10522
rect 9482 10464 9526 10502
rect 9598 10522 9640 10564
rect 9598 10502 9606 10522
rect 9626 10502 9640 10522
rect 9598 10464 9640 10502
rect 9690 10522 9734 10564
rect 9690 10502 9702 10522
rect 9722 10502 9734 10522
rect 9690 10464 9734 10502
rect 9811 10522 9853 10564
rect 9811 10502 9819 10522
rect 9839 10502 9853 10522
rect 9811 10464 9853 10502
rect 9903 10522 9947 10564
rect 12646 10621 12690 10663
rect 12740 10683 12782 10721
rect 12740 10663 12754 10683
rect 12774 10663 12782 10683
rect 12740 10621 12782 10663
rect 12859 10683 12903 10721
rect 12859 10663 12871 10683
rect 12891 10663 12903 10683
rect 12859 10621 12903 10663
rect 12953 10683 12995 10721
rect 12953 10663 12967 10683
rect 12987 10663 12995 10683
rect 12953 10621 12995 10663
rect 13067 10683 13111 10721
rect 13067 10663 13079 10683
rect 13099 10663 13111 10683
rect 13067 10621 13111 10663
rect 13161 10683 13203 10721
rect 13161 10663 13175 10683
rect 13195 10663 13203 10683
rect 13161 10621 13203 10663
rect 13277 10683 13319 10721
rect 13277 10663 13285 10683
rect 13305 10663 13319 10683
rect 13277 10621 13319 10663
rect 13369 10690 13414 10721
rect 13369 10683 13413 10690
rect 13369 10663 13381 10683
rect 13401 10663 13413 10683
rect 13369 10621 13413 10663
rect 22563 10691 22607 10729
rect 9903 10502 9915 10522
rect 9935 10502 9947 10522
rect 9903 10464 9947 10502
rect 17350 10519 17394 10561
rect 17350 10499 17362 10519
rect 17382 10499 17394 10519
rect 17350 10492 17394 10499
rect 17349 10461 17394 10492
rect 17444 10519 17486 10561
rect 17444 10499 17458 10519
rect 17478 10499 17486 10519
rect 17444 10461 17486 10499
rect 17560 10519 17602 10561
rect 17560 10499 17568 10519
rect 17588 10499 17602 10519
rect 17560 10461 17602 10499
rect 17652 10519 17696 10561
rect 17652 10499 17664 10519
rect 17684 10499 17696 10519
rect 17652 10461 17696 10499
rect 17768 10519 17810 10561
rect 17768 10499 17776 10519
rect 17796 10499 17810 10519
rect 17768 10461 17810 10499
rect 17860 10519 17904 10561
rect 17860 10499 17872 10519
rect 17892 10499 17904 10519
rect 17860 10461 17904 10499
rect 17981 10519 18023 10561
rect 17981 10499 17989 10519
rect 18009 10499 18023 10519
rect 17981 10461 18023 10499
rect 18073 10519 18117 10561
rect 22563 10671 22575 10691
rect 22595 10671 22607 10691
rect 22563 10629 22607 10671
rect 22657 10691 22699 10729
rect 22657 10671 22671 10691
rect 22691 10671 22699 10691
rect 22657 10629 22699 10671
rect 22776 10691 22820 10729
rect 22776 10671 22788 10691
rect 22808 10671 22820 10691
rect 22776 10629 22820 10671
rect 22870 10691 22912 10729
rect 22870 10671 22884 10691
rect 22904 10671 22912 10691
rect 22870 10629 22912 10671
rect 22984 10691 23028 10729
rect 22984 10671 22996 10691
rect 23016 10671 23028 10691
rect 22984 10629 23028 10671
rect 23078 10691 23120 10729
rect 23078 10671 23092 10691
rect 23112 10671 23120 10691
rect 23078 10629 23120 10671
rect 23194 10691 23236 10729
rect 23194 10671 23202 10691
rect 23222 10671 23236 10691
rect 23194 10629 23236 10671
rect 23286 10698 23331 10729
rect 23286 10691 23330 10698
rect 23286 10671 23298 10691
rect 23318 10671 23330 10691
rect 23286 10629 23330 10671
rect 23611 10687 23655 10725
rect 23611 10667 23623 10687
rect 23643 10667 23655 10687
rect 18073 10499 18085 10519
rect 18105 10499 18117 10519
rect 18073 10461 18117 10499
rect 19888 10516 19932 10558
rect 19888 10496 19900 10516
rect 19920 10496 19932 10516
rect 19888 10489 19932 10496
rect 19887 10458 19932 10489
rect 19982 10516 20024 10558
rect 19982 10496 19996 10516
rect 20016 10496 20024 10516
rect 19982 10458 20024 10496
rect 20098 10516 20140 10558
rect 20098 10496 20106 10516
rect 20126 10496 20140 10516
rect 20098 10458 20140 10496
rect 20190 10516 20234 10558
rect 20190 10496 20202 10516
rect 20222 10496 20234 10516
rect 20190 10458 20234 10496
rect 20306 10516 20348 10558
rect 20306 10496 20314 10516
rect 20334 10496 20348 10516
rect 20306 10458 20348 10496
rect 20398 10516 20442 10558
rect 20398 10496 20410 10516
rect 20430 10496 20442 10516
rect 20398 10458 20442 10496
rect 20519 10516 20561 10558
rect 20519 10496 20527 10516
rect 20547 10496 20561 10516
rect 20519 10458 20561 10496
rect 20611 10516 20655 10558
rect 23611 10625 23655 10667
rect 23705 10687 23747 10725
rect 23705 10667 23719 10687
rect 23739 10667 23747 10687
rect 23705 10625 23747 10667
rect 23824 10687 23868 10725
rect 23824 10667 23836 10687
rect 23856 10667 23868 10687
rect 23824 10625 23868 10667
rect 23918 10687 23960 10725
rect 23918 10667 23932 10687
rect 23952 10667 23960 10687
rect 23918 10625 23960 10667
rect 24032 10687 24076 10725
rect 24032 10667 24044 10687
rect 24064 10667 24076 10687
rect 24032 10625 24076 10667
rect 24126 10687 24168 10725
rect 24126 10667 24140 10687
rect 24160 10667 24168 10687
rect 24126 10625 24168 10667
rect 24242 10687 24284 10725
rect 24242 10667 24250 10687
rect 24270 10667 24284 10687
rect 24242 10625 24284 10667
rect 24334 10694 24379 10725
rect 24334 10687 24378 10694
rect 24334 10667 24346 10687
rect 24366 10667 24378 10687
rect 24334 10625 24378 10667
rect 20611 10496 20623 10516
rect 20643 10496 20655 10516
rect 20611 10458 20655 10496
rect 33271 10685 33315 10723
rect 28315 10523 28359 10565
rect 28315 10503 28327 10523
rect 28347 10503 28359 10523
rect 28315 10496 28359 10503
rect 28314 10465 28359 10496
rect 28409 10523 28451 10565
rect 28409 10503 28423 10523
rect 28443 10503 28451 10523
rect 28409 10465 28451 10503
rect 28525 10523 28567 10565
rect 28525 10503 28533 10523
rect 28553 10503 28567 10523
rect 28525 10465 28567 10503
rect 28617 10523 28661 10565
rect 28617 10503 28629 10523
rect 28649 10503 28661 10523
rect 28617 10465 28661 10503
rect 28733 10523 28775 10565
rect 28733 10503 28741 10523
rect 28761 10503 28775 10523
rect 28733 10465 28775 10503
rect 28825 10523 28869 10565
rect 28825 10503 28837 10523
rect 28857 10503 28869 10523
rect 28825 10465 28869 10503
rect 28946 10523 28988 10565
rect 28946 10503 28954 10523
rect 28974 10503 28988 10523
rect 28946 10465 28988 10503
rect 29038 10523 29082 10565
rect 33271 10665 33283 10685
rect 33303 10665 33315 10685
rect 33271 10623 33315 10665
rect 33365 10685 33407 10723
rect 33365 10665 33379 10685
rect 33399 10665 33407 10685
rect 33365 10623 33407 10665
rect 33484 10685 33528 10723
rect 33484 10665 33496 10685
rect 33516 10665 33528 10685
rect 33484 10623 33528 10665
rect 33578 10685 33620 10723
rect 33578 10665 33592 10685
rect 33612 10665 33620 10685
rect 33578 10623 33620 10665
rect 33692 10685 33736 10723
rect 33692 10665 33704 10685
rect 33724 10665 33736 10685
rect 33692 10623 33736 10665
rect 33786 10685 33828 10723
rect 33786 10665 33800 10685
rect 33820 10665 33828 10685
rect 33786 10623 33828 10665
rect 33902 10685 33944 10723
rect 33902 10665 33910 10685
rect 33930 10665 33944 10685
rect 33902 10623 33944 10665
rect 33994 10692 34039 10723
rect 33994 10685 34038 10692
rect 33994 10665 34006 10685
rect 34026 10665 34038 10685
rect 33994 10623 34038 10665
rect 34319 10681 34363 10719
rect 34319 10661 34331 10681
rect 34351 10661 34363 10681
rect 29038 10503 29050 10523
rect 29070 10503 29082 10523
rect 29038 10465 29082 10503
rect 30853 10520 30897 10562
rect 30853 10500 30865 10520
rect 30885 10500 30897 10520
rect 30853 10493 30897 10500
rect 30852 10462 30897 10493
rect 30947 10520 30989 10562
rect 30947 10500 30961 10520
rect 30981 10500 30989 10520
rect 30947 10462 30989 10500
rect 31063 10520 31105 10562
rect 31063 10500 31071 10520
rect 31091 10500 31105 10520
rect 31063 10462 31105 10500
rect 31155 10520 31199 10562
rect 31155 10500 31167 10520
rect 31187 10500 31199 10520
rect 31155 10462 31199 10500
rect 31271 10520 31313 10562
rect 31271 10500 31279 10520
rect 31299 10500 31313 10520
rect 31271 10462 31313 10500
rect 31363 10520 31407 10562
rect 31363 10500 31375 10520
rect 31395 10500 31407 10520
rect 31363 10462 31407 10500
rect 31484 10520 31526 10562
rect 31484 10500 31492 10520
rect 31512 10500 31526 10520
rect 31484 10462 31526 10500
rect 31576 10520 31620 10562
rect 34319 10619 34363 10661
rect 34413 10681 34455 10719
rect 34413 10661 34427 10681
rect 34447 10661 34455 10681
rect 34413 10619 34455 10661
rect 34532 10681 34576 10719
rect 34532 10661 34544 10681
rect 34564 10661 34576 10681
rect 34532 10619 34576 10661
rect 34626 10681 34668 10719
rect 34626 10661 34640 10681
rect 34660 10661 34668 10681
rect 34626 10619 34668 10661
rect 34740 10681 34784 10719
rect 34740 10661 34752 10681
rect 34772 10661 34784 10681
rect 34740 10619 34784 10661
rect 34834 10681 34876 10719
rect 34834 10661 34848 10681
rect 34868 10661 34876 10681
rect 34834 10619 34876 10661
rect 34950 10681 34992 10719
rect 34950 10661 34958 10681
rect 34978 10661 34992 10681
rect 34950 10619 34992 10661
rect 35042 10688 35087 10719
rect 35042 10681 35086 10688
rect 35042 10661 35054 10681
rect 35074 10661 35086 10681
rect 35042 10619 35086 10661
rect 31576 10500 31588 10520
rect 31608 10500 31620 10520
rect 31576 10462 31620 10500
rect 39023 10517 39067 10559
rect 39023 10497 39035 10517
rect 39055 10497 39067 10517
rect 39023 10490 39067 10497
rect 39022 10459 39067 10490
rect 39117 10517 39159 10559
rect 39117 10497 39131 10517
rect 39151 10497 39159 10517
rect 39117 10459 39159 10497
rect 39233 10517 39275 10559
rect 39233 10497 39241 10517
rect 39261 10497 39275 10517
rect 39233 10459 39275 10497
rect 39325 10517 39369 10559
rect 39325 10497 39337 10517
rect 39357 10497 39369 10517
rect 39325 10459 39369 10497
rect 39441 10517 39483 10559
rect 39441 10497 39449 10517
rect 39469 10497 39483 10517
rect 39441 10459 39483 10497
rect 39533 10517 39577 10559
rect 39533 10497 39545 10517
rect 39565 10497 39577 10517
rect 39533 10459 39577 10497
rect 39654 10517 39696 10559
rect 39654 10497 39662 10517
rect 39682 10497 39696 10517
rect 39654 10459 39696 10497
rect 39746 10517 39790 10559
rect 39746 10497 39758 10517
rect 39778 10497 39790 10517
rect 39746 10459 39790 10497
rect 41561 10514 41605 10556
rect 41561 10494 41573 10514
rect 41593 10494 41605 10514
rect 41561 10487 41605 10494
rect 41560 10456 41605 10487
rect 41655 10514 41697 10556
rect 41655 10494 41669 10514
rect 41689 10494 41697 10514
rect 41655 10456 41697 10494
rect 41771 10514 41813 10556
rect 41771 10494 41779 10514
rect 41799 10494 41813 10514
rect 41771 10456 41813 10494
rect 41863 10514 41907 10556
rect 41863 10494 41875 10514
rect 41895 10494 41907 10514
rect 41863 10456 41907 10494
rect 41979 10514 42021 10556
rect 41979 10494 41987 10514
rect 42007 10494 42021 10514
rect 41979 10456 42021 10494
rect 42071 10514 42115 10556
rect 42071 10494 42083 10514
rect 42103 10494 42115 10514
rect 42071 10456 42115 10494
rect 42192 10514 42234 10556
rect 42192 10494 42200 10514
rect 42220 10494 42234 10514
rect 42192 10456 42234 10494
rect 42284 10514 42328 10556
rect 42284 10494 42296 10514
rect 42316 10494 42328 10514
rect 42284 10456 42328 10494
rect 890 10014 934 10052
rect 890 9994 902 10014
rect 922 9994 934 10014
rect 890 9952 934 9994
rect 984 10014 1026 10052
rect 984 9994 998 10014
rect 1018 9994 1026 10014
rect 984 9952 1026 9994
rect 1103 10014 1147 10052
rect 1103 9994 1115 10014
rect 1135 9994 1147 10014
rect 1103 9952 1147 9994
rect 1197 10014 1239 10052
rect 1197 9994 1211 10014
rect 1231 9994 1239 10014
rect 1197 9952 1239 9994
rect 1311 10014 1355 10052
rect 1311 9994 1323 10014
rect 1343 9994 1355 10014
rect 1311 9952 1355 9994
rect 1405 10014 1447 10052
rect 1405 9994 1419 10014
rect 1439 9994 1447 10014
rect 1405 9952 1447 9994
rect 1521 10014 1563 10052
rect 1521 9994 1529 10014
rect 1549 9994 1563 10014
rect 1521 9952 1563 9994
rect 1613 10021 1658 10052
rect 1613 10014 1657 10021
rect 1613 9994 1625 10014
rect 1645 9994 1657 10014
rect 1613 9952 1657 9994
rect 3385 10009 3429 10047
rect 3385 9989 3397 10009
rect 3417 9989 3429 10009
rect 3385 9947 3429 9989
rect 3479 10009 3521 10047
rect 3479 9989 3493 10009
rect 3513 9989 3521 10009
rect 3479 9947 3521 9989
rect 3598 10009 3642 10047
rect 3598 9989 3610 10009
rect 3630 9989 3642 10009
rect 3598 9947 3642 9989
rect 3692 10009 3734 10047
rect 3692 9989 3706 10009
rect 3726 9989 3734 10009
rect 3692 9947 3734 9989
rect 3806 10009 3850 10047
rect 3806 9989 3818 10009
rect 3838 9989 3850 10009
rect 3806 9947 3850 9989
rect 3900 10009 3942 10047
rect 3900 9989 3914 10009
rect 3934 9989 3942 10009
rect 3900 9947 3942 9989
rect 4016 10009 4058 10047
rect 4016 9989 4024 10009
rect 4044 9989 4058 10009
rect 4016 9947 4058 9989
rect 4108 10016 4153 10047
rect 4108 10009 4152 10016
rect 4108 9989 4120 10009
rect 4140 9989 4152 10009
rect 4108 9947 4152 9989
rect 11598 10008 11642 10046
rect 11598 9988 11610 10008
rect 11630 9988 11642 10008
rect 8132 9847 8176 9889
rect 8132 9827 8144 9847
rect 8164 9827 8176 9847
rect 8132 9820 8176 9827
rect 8131 9789 8176 9820
rect 8226 9847 8268 9889
rect 8226 9827 8240 9847
rect 8260 9827 8268 9847
rect 8226 9789 8268 9827
rect 8342 9847 8384 9889
rect 8342 9827 8350 9847
rect 8370 9827 8384 9847
rect 8342 9789 8384 9827
rect 8434 9847 8478 9889
rect 8434 9827 8446 9847
rect 8466 9827 8478 9847
rect 8434 9789 8478 9827
rect 8550 9847 8592 9889
rect 8550 9827 8558 9847
rect 8578 9827 8592 9847
rect 8550 9789 8592 9827
rect 8642 9847 8686 9889
rect 8642 9827 8654 9847
rect 8674 9827 8686 9847
rect 8642 9789 8686 9827
rect 8763 9847 8805 9889
rect 8763 9827 8771 9847
rect 8791 9827 8805 9847
rect 8763 9789 8805 9827
rect 8855 9847 8899 9889
rect 11598 9946 11642 9988
rect 11692 10008 11734 10046
rect 11692 9988 11706 10008
rect 11726 9988 11734 10008
rect 11692 9946 11734 9988
rect 11811 10008 11855 10046
rect 11811 9988 11823 10008
rect 11843 9988 11855 10008
rect 11811 9946 11855 9988
rect 11905 10008 11947 10046
rect 11905 9988 11919 10008
rect 11939 9988 11947 10008
rect 11905 9946 11947 9988
rect 12019 10008 12063 10046
rect 12019 9988 12031 10008
rect 12051 9988 12063 10008
rect 12019 9946 12063 9988
rect 12113 10008 12155 10046
rect 12113 9988 12127 10008
rect 12147 9988 12155 10008
rect 12113 9946 12155 9988
rect 12229 10008 12271 10046
rect 12229 9988 12237 10008
rect 12257 9988 12271 10008
rect 12229 9946 12271 9988
rect 12321 10015 12366 10046
rect 12321 10008 12365 10015
rect 12321 9988 12333 10008
rect 12353 9988 12365 10008
rect 12321 9946 12365 9988
rect 14093 10003 14137 10041
rect 14093 9983 14105 10003
rect 14125 9983 14137 10003
rect 8855 9827 8867 9847
rect 8887 9827 8899 9847
rect 8855 9789 8899 9827
rect 9180 9843 9224 9885
rect 9180 9823 9192 9843
rect 9212 9823 9224 9843
rect 9180 9816 9224 9823
rect 9179 9785 9224 9816
rect 9274 9843 9316 9885
rect 9274 9823 9288 9843
rect 9308 9823 9316 9843
rect 9274 9785 9316 9823
rect 9390 9843 9432 9885
rect 9390 9823 9398 9843
rect 9418 9823 9432 9843
rect 9390 9785 9432 9823
rect 9482 9843 9526 9885
rect 9482 9823 9494 9843
rect 9514 9823 9526 9843
rect 9482 9785 9526 9823
rect 9598 9843 9640 9885
rect 9598 9823 9606 9843
rect 9626 9823 9640 9843
rect 9598 9785 9640 9823
rect 9690 9843 9734 9885
rect 9690 9823 9702 9843
rect 9722 9823 9734 9843
rect 9690 9785 9734 9823
rect 9811 9843 9853 9885
rect 9811 9823 9819 9843
rect 9839 9823 9853 9843
rect 9811 9785 9853 9823
rect 9903 9843 9947 9885
rect 9903 9823 9915 9843
rect 9935 9823 9947 9843
rect 14093 9941 14137 9983
rect 14187 10003 14229 10041
rect 14187 9983 14201 10003
rect 14221 9983 14229 10003
rect 14187 9941 14229 9983
rect 14306 10003 14350 10041
rect 14306 9983 14318 10003
rect 14338 9983 14350 10003
rect 14306 9941 14350 9983
rect 14400 10003 14442 10041
rect 14400 9983 14414 10003
rect 14434 9983 14442 10003
rect 14400 9941 14442 9983
rect 14514 10003 14558 10041
rect 14514 9983 14526 10003
rect 14546 9983 14558 10003
rect 14514 9941 14558 9983
rect 14608 10003 14650 10041
rect 14608 9983 14622 10003
rect 14642 9983 14650 10003
rect 14608 9941 14650 9983
rect 14724 10003 14766 10041
rect 14724 9983 14732 10003
rect 14752 9983 14766 10003
rect 14724 9941 14766 9983
rect 14816 10010 14861 10041
rect 14816 10003 14860 10010
rect 14816 9983 14828 10003
rect 14848 9983 14860 10003
rect 14816 9941 14860 9983
rect 9903 9785 9947 9823
rect 22563 10012 22607 10050
rect 22563 9992 22575 10012
rect 22595 9992 22607 10012
rect 18840 9841 18884 9883
rect 18840 9821 18852 9841
rect 18872 9821 18884 9841
rect 18840 9814 18884 9821
rect 18839 9783 18884 9814
rect 18934 9841 18976 9883
rect 18934 9821 18948 9841
rect 18968 9821 18976 9841
rect 18934 9783 18976 9821
rect 19050 9841 19092 9883
rect 19050 9821 19058 9841
rect 19078 9821 19092 9841
rect 19050 9783 19092 9821
rect 19142 9841 19186 9883
rect 19142 9821 19154 9841
rect 19174 9821 19186 9841
rect 19142 9783 19186 9821
rect 19258 9841 19300 9883
rect 19258 9821 19266 9841
rect 19286 9821 19300 9841
rect 19258 9783 19300 9821
rect 19350 9841 19394 9883
rect 19350 9821 19362 9841
rect 19382 9821 19394 9841
rect 19350 9783 19394 9821
rect 19471 9841 19513 9883
rect 19471 9821 19479 9841
rect 19499 9821 19513 9841
rect 19471 9783 19513 9821
rect 19563 9841 19607 9883
rect 22563 9950 22607 9992
rect 22657 10012 22699 10050
rect 22657 9992 22671 10012
rect 22691 9992 22699 10012
rect 22657 9950 22699 9992
rect 22776 10012 22820 10050
rect 22776 9992 22788 10012
rect 22808 9992 22820 10012
rect 22776 9950 22820 9992
rect 22870 10012 22912 10050
rect 22870 9992 22884 10012
rect 22904 9992 22912 10012
rect 22870 9950 22912 9992
rect 22984 10012 23028 10050
rect 22984 9992 22996 10012
rect 23016 9992 23028 10012
rect 22984 9950 23028 9992
rect 23078 10012 23120 10050
rect 23078 9992 23092 10012
rect 23112 9992 23120 10012
rect 23078 9950 23120 9992
rect 23194 10012 23236 10050
rect 23194 9992 23202 10012
rect 23222 9992 23236 10012
rect 23194 9950 23236 9992
rect 23286 10019 23331 10050
rect 23286 10012 23330 10019
rect 23286 9992 23298 10012
rect 23318 9992 23330 10012
rect 23286 9950 23330 9992
rect 25058 10007 25102 10045
rect 25058 9987 25070 10007
rect 25090 9987 25102 10007
rect 19563 9821 19575 9841
rect 19595 9821 19607 9841
rect 19563 9783 19607 9821
rect 19888 9837 19932 9879
rect 19888 9817 19900 9837
rect 19920 9817 19932 9837
rect 19888 9810 19932 9817
rect 19887 9779 19932 9810
rect 19982 9837 20024 9879
rect 19982 9817 19996 9837
rect 20016 9817 20024 9837
rect 19982 9779 20024 9817
rect 20098 9837 20140 9879
rect 20098 9817 20106 9837
rect 20126 9817 20140 9837
rect 20098 9779 20140 9817
rect 20190 9837 20234 9879
rect 20190 9817 20202 9837
rect 20222 9817 20234 9837
rect 20190 9779 20234 9817
rect 20306 9837 20348 9879
rect 20306 9817 20314 9837
rect 20334 9817 20348 9837
rect 20306 9779 20348 9817
rect 20398 9837 20442 9879
rect 20398 9817 20410 9837
rect 20430 9817 20442 9837
rect 20398 9779 20442 9817
rect 20519 9837 20561 9879
rect 20519 9817 20527 9837
rect 20547 9817 20561 9837
rect 20519 9779 20561 9817
rect 20611 9837 20655 9879
rect 20611 9817 20623 9837
rect 20643 9817 20655 9837
rect 25058 9945 25102 9987
rect 25152 10007 25194 10045
rect 25152 9987 25166 10007
rect 25186 9987 25194 10007
rect 25152 9945 25194 9987
rect 25271 10007 25315 10045
rect 25271 9987 25283 10007
rect 25303 9987 25315 10007
rect 25271 9945 25315 9987
rect 25365 10007 25407 10045
rect 25365 9987 25379 10007
rect 25399 9987 25407 10007
rect 25365 9945 25407 9987
rect 25479 10007 25523 10045
rect 25479 9987 25491 10007
rect 25511 9987 25523 10007
rect 25479 9945 25523 9987
rect 25573 10007 25615 10045
rect 25573 9987 25587 10007
rect 25607 9987 25615 10007
rect 25573 9945 25615 9987
rect 25689 10007 25731 10045
rect 25689 9987 25697 10007
rect 25717 9987 25731 10007
rect 25689 9945 25731 9987
rect 25781 10014 25826 10045
rect 25781 10007 25825 10014
rect 25781 9987 25793 10007
rect 25813 9987 25825 10007
rect 25781 9945 25825 9987
rect 33271 10006 33315 10044
rect 33271 9986 33283 10006
rect 33303 9986 33315 10006
rect 20611 9779 20655 9817
rect 29805 9845 29849 9887
rect 29805 9825 29817 9845
rect 29837 9825 29849 9845
rect 29805 9818 29849 9825
rect 29804 9787 29849 9818
rect 29899 9845 29941 9887
rect 29899 9825 29913 9845
rect 29933 9825 29941 9845
rect 29899 9787 29941 9825
rect 30015 9845 30057 9887
rect 30015 9825 30023 9845
rect 30043 9825 30057 9845
rect 30015 9787 30057 9825
rect 30107 9845 30151 9887
rect 30107 9825 30119 9845
rect 30139 9825 30151 9845
rect 30107 9787 30151 9825
rect 30223 9845 30265 9887
rect 30223 9825 30231 9845
rect 30251 9825 30265 9845
rect 30223 9787 30265 9825
rect 30315 9845 30359 9887
rect 30315 9825 30327 9845
rect 30347 9825 30359 9845
rect 30315 9787 30359 9825
rect 30436 9845 30478 9887
rect 30436 9825 30444 9845
rect 30464 9825 30478 9845
rect 30436 9787 30478 9825
rect 30528 9845 30572 9887
rect 33271 9944 33315 9986
rect 33365 10006 33407 10044
rect 33365 9986 33379 10006
rect 33399 9986 33407 10006
rect 33365 9944 33407 9986
rect 33484 10006 33528 10044
rect 33484 9986 33496 10006
rect 33516 9986 33528 10006
rect 33484 9944 33528 9986
rect 33578 10006 33620 10044
rect 33578 9986 33592 10006
rect 33612 9986 33620 10006
rect 33578 9944 33620 9986
rect 33692 10006 33736 10044
rect 33692 9986 33704 10006
rect 33724 9986 33736 10006
rect 33692 9944 33736 9986
rect 33786 10006 33828 10044
rect 33786 9986 33800 10006
rect 33820 9986 33828 10006
rect 33786 9944 33828 9986
rect 33902 10006 33944 10044
rect 33902 9986 33910 10006
rect 33930 9986 33944 10006
rect 33902 9944 33944 9986
rect 33994 10013 34039 10044
rect 33994 10006 34038 10013
rect 33994 9986 34006 10006
rect 34026 9986 34038 10006
rect 33994 9944 34038 9986
rect 35766 10001 35810 10039
rect 35766 9981 35778 10001
rect 35798 9981 35810 10001
rect 30528 9825 30540 9845
rect 30560 9825 30572 9845
rect 30528 9787 30572 9825
rect 30853 9841 30897 9883
rect 30853 9821 30865 9841
rect 30885 9821 30897 9841
rect 30853 9814 30897 9821
rect 30852 9783 30897 9814
rect 30947 9841 30989 9883
rect 30947 9821 30961 9841
rect 30981 9821 30989 9841
rect 30947 9783 30989 9821
rect 31063 9841 31105 9883
rect 31063 9821 31071 9841
rect 31091 9821 31105 9841
rect 31063 9783 31105 9821
rect 31155 9841 31199 9883
rect 31155 9821 31167 9841
rect 31187 9821 31199 9841
rect 31155 9783 31199 9821
rect 31271 9841 31313 9883
rect 31271 9821 31279 9841
rect 31299 9821 31313 9841
rect 31271 9783 31313 9821
rect 31363 9841 31407 9883
rect 31363 9821 31375 9841
rect 31395 9821 31407 9841
rect 31363 9783 31407 9821
rect 31484 9841 31526 9883
rect 31484 9821 31492 9841
rect 31512 9821 31526 9841
rect 31484 9783 31526 9821
rect 31576 9841 31620 9883
rect 31576 9821 31588 9841
rect 31608 9821 31620 9841
rect 35766 9939 35810 9981
rect 35860 10001 35902 10039
rect 35860 9981 35874 10001
rect 35894 9981 35902 10001
rect 35860 9939 35902 9981
rect 35979 10001 36023 10039
rect 35979 9981 35991 10001
rect 36011 9981 36023 10001
rect 35979 9939 36023 9981
rect 36073 10001 36115 10039
rect 36073 9981 36087 10001
rect 36107 9981 36115 10001
rect 36073 9939 36115 9981
rect 36187 10001 36231 10039
rect 36187 9981 36199 10001
rect 36219 9981 36231 10001
rect 36187 9939 36231 9981
rect 36281 10001 36323 10039
rect 36281 9981 36295 10001
rect 36315 9981 36323 10001
rect 36281 9939 36323 9981
rect 36397 10001 36439 10039
rect 36397 9981 36405 10001
rect 36425 9981 36439 10001
rect 36397 9939 36439 9981
rect 36489 10008 36534 10039
rect 36489 10001 36533 10008
rect 36489 9981 36501 10001
rect 36521 9981 36533 10001
rect 36489 9939 36533 9981
rect 31576 9783 31620 9821
rect 40513 9839 40557 9881
rect 40513 9819 40525 9839
rect 40545 9819 40557 9839
rect 40513 9812 40557 9819
rect 40512 9781 40557 9812
rect 40607 9839 40649 9881
rect 40607 9819 40621 9839
rect 40641 9819 40649 9839
rect 40607 9781 40649 9819
rect 40723 9839 40765 9881
rect 40723 9819 40731 9839
rect 40751 9819 40765 9839
rect 40723 9781 40765 9819
rect 40815 9839 40859 9881
rect 40815 9819 40827 9839
rect 40847 9819 40859 9839
rect 40815 9781 40859 9819
rect 40931 9839 40973 9881
rect 40931 9819 40939 9839
rect 40959 9819 40973 9839
rect 40931 9781 40973 9819
rect 41023 9839 41067 9881
rect 41023 9819 41035 9839
rect 41055 9819 41067 9839
rect 41023 9781 41067 9819
rect 41144 9839 41186 9881
rect 41144 9819 41152 9839
rect 41172 9819 41186 9839
rect 41144 9781 41186 9819
rect 41236 9839 41280 9881
rect 41236 9819 41248 9839
rect 41268 9819 41280 9839
rect 41236 9781 41280 9819
rect 41561 9835 41605 9877
rect 41561 9815 41573 9835
rect 41593 9815 41605 9835
rect 41561 9808 41605 9815
rect 41560 9777 41605 9808
rect 41655 9835 41697 9877
rect 41655 9815 41669 9835
rect 41689 9815 41697 9835
rect 41655 9777 41697 9815
rect 41771 9835 41813 9877
rect 41771 9815 41779 9835
rect 41799 9815 41813 9835
rect 41771 9777 41813 9815
rect 41863 9835 41907 9877
rect 41863 9815 41875 9835
rect 41895 9815 41907 9835
rect 41863 9777 41907 9815
rect 41979 9835 42021 9877
rect 41979 9815 41987 9835
rect 42007 9815 42021 9835
rect 41979 9777 42021 9815
rect 42071 9835 42115 9877
rect 42071 9815 42083 9835
rect 42103 9815 42115 9835
rect 42071 9777 42115 9815
rect 42192 9835 42234 9877
rect 42192 9815 42200 9835
rect 42220 9815 42234 9835
rect 42192 9777 42234 9815
rect 42284 9835 42328 9877
rect 42284 9815 42296 9835
rect 42316 9815 42328 9835
rect 42284 9777 42328 9815
rect 890 9246 934 9284
rect 890 9226 902 9246
rect 922 9226 934 9246
rect 890 9184 934 9226
rect 984 9246 1026 9284
rect 984 9226 998 9246
rect 1018 9226 1026 9246
rect 984 9184 1026 9226
rect 1103 9246 1147 9284
rect 1103 9226 1115 9246
rect 1135 9226 1147 9246
rect 1103 9184 1147 9226
rect 1197 9246 1239 9284
rect 1197 9226 1211 9246
rect 1231 9226 1239 9246
rect 1197 9184 1239 9226
rect 1311 9246 1355 9284
rect 1311 9226 1323 9246
rect 1343 9226 1355 9246
rect 1311 9184 1355 9226
rect 1405 9246 1447 9284
rect 1405 9226 1419 9246
rect 1439 9226 1447 9246
rect 1405 9184 1447 9226
rect 1521 9246 1563 9284
rect 1521 9226 1529 9246
rect 1549 9226 1563 9246
rect 1521 9184 1563 9226
rect 1613 9253 1658 9284
rect 1613 9246 1657 9253
rect 1613 9226 1625 9246
rect 1645 9226 1657 9246
rect 1613 9184 1657 9226
rect 1938 9242 1982 9280
rect 1938 9222 1950 9242
rect 1970 9222 1982 9242
rect 1938 9180 1982 9222
rect 2032 9242 2074 9280
rect 2032 9222 2046 9242
rect 2066 9222 2074 9242
rect 2032 9180 2074 9222
rect 2151 9242 2195 9280
rect 2151 9222 2163 9242
rect 2183 9222 2195 9242
rect 2151 9180 2195 9222
rect 2245 9242 2287 9280
rect 2245 9222 2259 9242
rect 2279 9222 2287 9242
rect 2245 9180 2287 9222
rect 2359 9242 2403 9280
rect 2359 9222 2371 9242
rect 2391 9222 2403 9242
rect 2359 9180 2403 9222
rect 2453 9242 2495 9280
rect 2453 9222 2467 9242
rect 2487 9222 2495 9242
rect 2453 9180 2495 9222
rect 2569 9242 2611 9280
rect 2569 9222 2577 9242
rect 2597 9222 2611 9242
rect 2569 9180 2611 9222
rect 2661 9249 2706 9280
rect 2661 9242 2705 9249
rect 2661 9222 2673 9242
rect 2693 9222 2705 9242
rect 2661 9180 2705 9222
rect 11598 9240 11642 9278
rect 6685 9080 6729 9122
rect 6685 9060 6697 9080
rect 6717 9060 6729 9080
rect 6685 9053 6729 9060
rect 6684 9022 6729 9053
rect 6779 9080 6821 9122
rect 6779 9060 6793 9080
rect 6813 9060 6821 9080
rect 6779 9022 6821 9060
rect 6895 9080 6937 9122
rect 6895 9060 6903 9080
rect 6923 9060 6937 9080
rect 6895 9022 6937 9060
rect 6987 9080 7031 9122
rect 6987 9060 6999 9080
rect 7019 9060 7031 9080
rect 6987 9022 7031 9060
rect 7103 9080 7145 9122
rect 7103 9060 7111 9080
rect 7131 9060 7145 9080
rect 7103 9022 7145 9060
rect 7195 9080 7239 9122
rect 7195 9060 7207 9080
rect 7227 9060 7239 9080
rect 7195 9022 7239 9060
rect 7316 9080 7358 9122
rect 7316 9060 7324 9080
rect 7344 9060 7358 9080
rect 7316 9022 7358 9060
rect 7408 9080 7452 9122
rect 11598 9220 11610 9240
rect 11630 9220 11642 9240
rect 11598 9178 11642 9220
rect 11692 9240 11734 9278
rect 11692 9220 11706 9240
rect 11726 9220 11734 9240
rect 11692 9178 11734 9220
rect 11811 9240 11855 9278
rect 11811 9220 11823 9240
rect 11843 9220 11855 9240
rect 11811 9178 11855 9220
rect 11905 9240 11947 9278
rect 11905 9220 11919 9240
rect 11939 9220 11947 9240
rect 11905 9178 11947 9220
rect 12019 9240 12063 9278
rect 12019 9220 12031 9240
rect 12051 9220 12063 9240
rect 12019 9178 12063 9220
rect 12113 9240 12155 9278
rect 12113 9220 12127 9240
rect 12147 9220 12155 9240
rect 12113 9178 12155 9220
rect 12229 9240 12271 9278
rect 12229 9220 12237 9240
rect 12257 9220 12271 9240
rect 12229 9178 12271 9220
rect 12321 9247 12366 9278
rect 12321 9240 12365 9247
rect 12321 9220 12333 9240
rect 12353 9220 12365 9240
rect 12321 9178 12365 9220
rect 12646 9236 12690 9274
rect 12646 9216 12658 9236
rect 12678 9216 12690 9236
rect 7408 9060 7420 9080
rect 7440 9060 7452 9080
rect 7408 9022 7452 9060
rect 9180 9075 9224 9117
rect 9180 9055 9192 9075
rect 9212 9055 9224 9075
rect 9180 9048 9224 9055
rect 9179 9017 9224 9048
rect 9274 9075 9316 9117
rect 9274 9055 9288 9075
rect 9308 9055 9316 9075
rect 9274 9017 9316 9055
rect 9390 9075 9432 9117
rect 9390 9055 9398 9075
rect 9418 9055 9432 9075
rect 9390 9017 9432 9055
rect 9482 9075 9526 9117
rect 9482 9055 9494 9075
rect 9514 9055 9526 9075
rect 9482 9017 9526 9055
rect 9598 9075 9640 9117
rect 9598 9055 9606 9075
rect 9626 9055 9640 9075
rect 9598 9017 9640 9055
rect 9690 9075 9734 9117
rect 9690 9055 9702 9075
rect 9722 9055 9734 9075
rect 9690 9017 9734 9055
rect 9811 9075 9853 9117
rect 9811 9055 9819 9075
rect 9839 9055 9853 9075
rect 9811 9017 9853 9055
rect 9903 9075 9947 9117
rect 12646 9174 12690 9216
rect 12740 9236 12782 9274
rect 12740 9216 12754 9236
rect 12774 9216 12782 9236
rect 12740 9174 12782 9216
rect 12859 9236 12903 9274
rect 12859 9216 12871 9236
rect 12891 9216 12903 9236
rect 12859 9174 12903 9216
rect 12953 9236 12995 9274
rect 12953 9216 12967 9236
rect 12987 9216 12995 9236
rect 12953 9174 12995 9216
rect 13067 9236 13111 9274
rect 13067 9216 13079 9236
rect 13099 9216 13111 9236
rect 13067 9174 13111 9216
rect 13161 9236 13203 9274
rect 13161 9216 13175 9236
rect 13195 9216 13203 9236
rect 13161 9174 13203 9216
rect 13277 9236 13319 9274
rect 13277 9216 13285 9236
rect 13305 9216 13319 9236
rect 13277 9174 13319 9216
rect 13369 9243 13414 9274
rect 13369 9236 13413 9243
rect 13369 9216 13381 9236
rect 13401 9216 13413 9236
rect 13369 9174 13413 9216
rect 22563 9244 22607 9282
rect 9903 9055 9915 9075
rect 9935 9055 9947 9075
rect 9903 9017 9947 9055
rect 17393 9074 17437 9116
rect 17393 9054 17405 9074
rect 17425 9054 17437 9074
rect 17393 9047 17437 9054
rect 17392 9016 17437 9047
rect 17487 9074 17529 9116
rect 17487 9054 17501 9074
rect 17521 9054 17529 9074
rect 17487 9016 17529 9054
rect 17603 9074 17645 9116
rect 17603 9054 17611 9074
rect 17631 9054 17645 9074
rect 17603 9016 17645 9054
rect 17695 9074 17739 9116
rect 17695 9054 17707 9074
rect 17727 9054 17739 9074
rect 17695 9016 17739 9054
rect 17811 9074 17853 9116
rect 17811 9054 17819 9074
rect 17839 9054 17853 9074
rect 17811 9016 17853 9054
rect 17903 9074 17947 9116
rect 17903 9054 17915 9074
rect 17935 9054 17947 9074
rect 17903 9016 17947 9054
rect 18024 9074 18066 9116
rect 18024 9054 18032 9074
rect 18052 9054 18066 9074
rect 18024 9016 18066 9054
rect 18116 9074 18160 9116
rect 22563 9224 22575 9244
rect 22595 9224 22607 9244
rect 22563 9182 22607 9224
rect 22657 9244 22699 9282
rect 22657 9224 22671 9244
rect 22691 9224 22699 9244
rect 22657 9182 22699 9224
rect 22776 9244 22820 9282
rect 22776 9224 22788 9244
rect 22808 9224 22820 9244
rect 22776 9182 22820 9224
rect 22870 9244 22912 9282
rect 22870 9224 22884 9244
rect 22904 9224 22912 9244
rect 22870 9182 22912 9224
rect 22984 9244 23028 9282
rect 22984 9224 22996 9244
rect 23016 9224 23028 9244
rect 22984 9182 23028 9224
rect 23078 9244 23120 9282
rect 23078 9224 23092 9244
rect 23112 9224 23120 9244
rect 23078 9182 23120 9224
rect 23194 9244 23236 9282
rect 23194 9224 23202 9244
rect 23222 9224 23236 9244
rect 23194 9182 23236 9224
rect 23286 9251 23331 9282
rect 23286 9244 23330 9251
rect 23286 9224 23298 9244
rect 23318 9224 23330 9244
rect 23286 9182 23330 9224
rect 23611 9240 23655 9278
rect 23611 9220 23623 9240
rect 23643 9220 23655 9240
rect 18116 9054 18128 9074
rect 18148 9054 18160 9074
rect 18116 9016 18160 9054
rect 19888 9069 19932 9111
rect 19888 9049 19900 9069
rect 19920 9049 19932 9069
rect 19888 9042 19932 9049
rect 19887 9011 19932 9042
rect 19982 9069 20024 9111
rect 19982 9049 19996 9069
rect 20016 9049 20024 9069
rect 19982 9011 20024 9049
rect 20098 9069 20140 9111
rect 20098 9049 20106 9069
rect 20126 9049 20140 9069
rect 20098 9011 20140 9049
rect 20190 9069 20234 9111
rect 20190 9049 20202 9069
rect 20222 9049 20234 9069
rect 20190 9011 20234 9049
rect 20306 9069 20348 9111
rect 20306 9049 20314 9069
rect 20334 9049 20348 9069
rect 20306 9011 20348 9049
rect 20398 9069 20442 9111
rect 20398 9049 20410 9069
rect 20430 9049 20442 9069
rect 20398 9011 20442 9049
rect 20519 9069 20561 9111
rect 20519 9049 20527 9069
rect 20547 9049 20561 9069
rect 20519 9011 20561 9049
rect 20611 9069 20655 9111
rect 23611 9178 23655 9220
rect 23705 9240 23747 9278
rect 23705 9220 23719 9240
rect 23739 9220 23747 9240
rect 23705 9178 23747 9220
rect 23824 9240 23868 9278
rect 23824 9220 23836 9240
rect 23856 9220 23868 9240
rect 23824 9178 23868 9220
rect 23918 9240 23960 9278
rect 23918 9220 23932 9240
rect 23952 9220 23960 9240
rect 23918 9178 23960 9220
rect 24032 9240 24076 9278
rect 24032 9220 24044 9240
rect 24064 9220 24076 9240
rect 24032 9178 24076 9220
rect 24126 9240 24168 9278
rect 24126 9220 24140 9240
rect 24160 9220 24168 9240
rect 24126 9178 24168 9220
rect 24242 9240 24284 9278
rect 24242 9220 24250 9240
rect 24270 9220 24284 9240
rect 24242 9178 24284 9220
rect 24334 9247 24379 9278
rect 24334 9240 24378 9247
rect 24334 9220 24346 9240
rect 24366 9220 24378 9240
rect 24334 9178 24378 9220
rect 20611 9049 20623 9069
rect 20643 9049 20655 9069
rect 20611 9011 20655 9049
rect 33271 9238 33315 9276
rect 28358 9078 28402 9120
rect 28358 9058 28370 9078
rect 28390 9058 28402 9078
rect 28358 9051 28402 9058
rect 28357 9020 28402 9051
rect 28452 9078 28494 9120
rect 28452 9058 28466 9078
rect 28486 9058 28494 9078
rect 28452 9020 28494 9058
rect 28568 9078 28610 9120
rect 28568 9058 28576 9078
rect 28596 9058 28610 9078
rect 28568 9020 28610 9058
rect 28660 9078 28704 9120
rect 28660 9058 28672 9078
rect 28692 9058 28704 9078
rect 28660 9020 28704 9058
rect 28776 9078 28818 9120
rect 28776 9058 28784 9078
rect 28804 9058 28818 9078
rect 28776 9020 28818 9058
rect 28868 9078 28912 9120
rect 28868 9058 28880 9078
rect 28900 9058 28912 9078
rect 28868 9020 28912 9058
rect 28989 9078 29031 9120
rect 28989 9058 28997 9078
rect 29017 9058 29031 9078
rect 28989 9020 29031 9058
rect 29081 9078 29125 9120
rect 33271 9218 33283 9238
rect 33303 9218 33315 9238
rect 33271 9176 33315 9218
rect 33365 9238 33407 9276
rect 33365 9218 33379 9238
rect 33399 9218 33407 9238
rect 33365 9176 33407 9218
rect 33484 9238 33528 9276
rect 33484 9218 33496 9238
rect 33516 9218 33528 9238
rect 33484 9176 33528 9218
rect 33578 9238 33620 9276
rect 33578 9218 33592 9238
rect 33612 9218 33620 9238
rect 33578 9176 33620 9218
rect 33692 9238 33736 9276
rect 33692 9218 33704 9238
rect 33724 9218 33736 9238
rect 33692 9176 33736 9218
rect 33786 9238 33828 9276
rect 33786 9218 33800 9238
rect 33820 9218 33828 9238
rect 33786 9176 33828 9218
rect 33902 9238 33944 9276
rect 33902 9218 33910 9238
rect 33930 9218 33944 9238
rect 33902 9176 33944 9218
rect 33994 9245 34039 9276
rect 33994 9238 34038 9245
rect 33994 9218 34006 9238
rect 34026 9218 34038 9238
rect 33994 9176 34038 9218
rect 34319 9234 34363 9272
rect 34319 9214 34331 9234
rect 34351 9214 34363 9234
rect 29081 9058 29093 9078
rect 29113 9058 29125 9078
rect 29081 9020 29125 9058
rect 30853 9073 30897 9115
rect 30853 9053 30865 9073
rect 30885 9053 30897 9073
rect 30853 9046 30897 9053
rect 30852 9015 30897 9046
rect 30947 9073 30989 9115
rect 30947 9053 30961 9073
rect 30981 9053 30989 9073
rect 30947 9015 30989 9053
rect 31063 9073 31105 9115
rect 31063 9053 31071 9073
rect 31091 9053 31105 9073
rect 31063 9015 31105 9053
rect 31155 9073 31199 9115
rect 31155 9053 31167 9073
rect 31187 9053 31199 9073
rect 31155 9015 31199 9053
rect 31271 9073 31313 9115
rect 31271 9053 31279 9073
rect 31299 9053 31313 9073
rect 31271 9015 31313 9053
rect 31363 9073 31407 9115
rect 31363 9053 31375 9073
rect 31395 9053 31407 9073
rect 31363 9015 31407 9053
rect 31484 9073 31526 9115
rect 31484 9053 31492 9073
rect 31512 9053 31526 9073
rect 31484 9015 31526 9053
rect 31576 9073 31620 9115
rect 34319 9172 34363 9214
rect 34413 9234 34455 9272
rect 34413 9214 34427 9234
rect 34447 9214 34455 9234
rect 34413 9172 34455 9214
rect 34532 9234 34576 9272
rect 34532 9214 34544 9234
rect 34564 9214 34576 9234
rect 34532 9172 34576 9214
rect 34626 9234 34668 9272
rect 34626 9214 34640 9234
rect 34660 9214 34668 9234
rect 34626 9172 34668 9214
rect 34740 9234 34784 9272
rect 34740 9214 34752 9234
rect 34772 9214 34784 9234
rect 34740 9172 34784 9214
rect 34834 9234 34876 9272
rect 34834 9214 34848 9234
rect 34868 9214 34876 9234
rect 34834 9172 34876 9214
rect 34950 9234 34992 9272
rect 34950 9214 34958 9234
rect 34978 9214 34992 9234
rect 34950 9172 34992 9214
rect 35042 9241 35087 9272
rect 35042 9234 35086 9241
rect 35042 9214 35054 9234
rect 35074 9214 35086 9234
rect 35042 9172 35086 9214
rect 31576 9053 31588 9073
rect 31608 9053 31620 9073
rect 31576 9015 31620 9053
rect 39066 9072 39110 9114
rect 39066 9052 39078 9072
rect 39098 9052 39110 9072
rect 39066 9045 39110 9052
rect 39065 9014 39110 9045
rect 39160 9072 39202 9114
rect 39160 9052 39174 9072
rect 39194 9052 39202 9072
rect 39160 9014 39202 9052
rect 39276 9072 39318 9114
rect 39276 9052 39284 9072
rect 39304 9052 39318 9072
rect 39276 9014 39318 9052
rect 39368 9072 39412 9114
rect 39368 9052 39380 9072
rect 39400 9052 39412 9072
rect 39368 9014 39412 9052
rect 39484 9072 39526 9114
rect 39484 9052 39492 9072
rect 39512 9052 39526 9072
rect 39484 9014 39526 9052
rect 39576 9072 39620 9114
rect 39576 9052 39588 9072
rect 39608 9052 39620 9072
rect 39576 9014 39620 9052
rect 39697 9072 39739 9114
rect 39697 9052 39705 9072
rect 39725 9052 39739 9072
rect 39697 9014 39739 9052
rect 39789 9072 39833 9114
rect 39789 9052 39801 9072
rect 39821 9052 39833 9072
rect 39789 9014 39833 9052
rect 41561 9067 41605 9109
rect 41561 9047 41573 9067
rect 41593 9047 41605 9067
rect 41561 9040 41605 9047
rect 41560 9009 41605 9040
rect 41655 9067 41697 9109
rect 41655 9047 41669 9067
rect 41689 9047 41697 9067
rect 41655 9009 41697 9047
rect 41771 9067 41813 9109
rect 41771 9047 41779 9067
rect 41799 9047 41813 9067
rect 41771 9009 41813 9047
rect 41863 9067 41907 9109
rect 41863 9047 41875 9067
rect 41895 9047 41907 9067
rect 41863 9009 41907 9047
rect 41979 9067 42021 9109
rect 41979 9047 41987 9067
rect 42007 9047 42021 9067
rect 41979 9009 42021 9047
rect 42071 9067 42115 9109
rect 42071 9047 42083 9067
rect 42103 9047 42115 9067
rect 42071 9009 42115 9047
rect 42192 9067 42234 9109
rect 42192 9047 42200 9067
rect 42220 9047 42234 9067
rect 42192 9009 42234 9047
rect 42284 9067 42328 9109
rect 42284 9047 42296 9067
rect 42316 9047 42328 9067
rect 42284 9009 42328 9047
rect 890 8567 934 8605
rect 890 8547 902 8567
rect 922 8547 934 8567
rect 890 8505 934 8547
rect 984 8567 1026 8605
rect 984 8547 998 8567
rect 1018 8547 1026 8567
rect 984 8505 1026 8547
rect 1103 8567 1147 8605
rect 1103 8547 1115 8567
rect 1135 8547 1147 8567
rect 1103 8505 1147 8547
rect 1197 8567 1239 8605
rect 1197 8547 1211 8567
rect 1231 8547 1239 8567
rect 1197 8505 1239 8547
rect 1311 8567 1355 8605
rect 1311 8547 1323 8567
rect 1343 8547 1355 8567
rect 1311 8505 1355 8547
rect 1405 8567 1447 8605
rect 1405 8547 1419 8567
rect 1439 8547 1447 8567
rect 1405 8505 1447 8547
rect 1521 8567 1563 8605
rect 1521 8547 1529 8567
rect 1549 8547 1563 8567
rect 1521 8505 1563 8547
rect 1613 8574 1658 8605
rect 1613 8567 1657 8574
rect 1613 8547 1625 8567
rect 1645 8547 1657 8567
rect 1613 8505 1657 8547
rect 4493 8558 4537 8596
rect 4493 8538 4505 8558
rect 4525 8538 4537 8558
rect 4493 8496 4537 8538
rect 4587 8558 4629 8596
rect 4587 8538 4601 8558
rect 4621 8538 4629 8558
rect 4587 8496 4629 8538
rect 4706 8558 4750 8596
rect 4706 8538 4718 8558
rect 4738 8538 4750 8558
rect 4706 8496 4750 8538
rect 4800 8558 4842 8596
rect 4800 8538 4814 8558
rect 4834 8538 4842 8558
rect 4800 8496 4842 8538
rect 4914 8558 4958 8596
rect 4914 8538 4926 8558
rect 4946 8538 4958 8558
rect 4914 8496 4958 8538
rect 5008 8558 5050 8596
rect 5008 8538 5022 8558
rect 5042 8538 5050 8558
rect 5008 8496 5050 8538
rect 5124 8558 5166 8596
rect 5124 8538 5132 8558
rect 5152 8538 5166 8558
rect 5124 8496 5166 8538
rect 5216 8565 5261 8596
rect 5216 8558 5260 8565
rect 5216 8538 5228 8558
rect 5248 8538 5260 8558
rect 5216 8496 5260 8538
rect 11598 8561 11642 8599
rect 11598 8541 11610 8561
rect 11630 8541 11642 8561
rect 8132 8400 8176 8442
rect 8132 8380 8144 8400
rect 8164 8380 8176 8400
rect 8132 8373 8176 8380
rect 8131 8342 8176 8373
rect 8226 8400 8268 8442
rect 8226 8380 8240 8400
rect 8260 8380 8268 8400
rect 8226 8342 8268 8380
rect 8342 8400 8384 8442
rect 8342 8380 8350 8400
rect 8370 8380 8384 8400
rect 8342 8342 8384 8380
rect 8434 8400 8478 8442
rect 8434 8380 8446 8400
rect 8466 8380 8478 8400
rect 8434 8342 8478 8380
rect 8550 8400 8592 8442
rect 8550 8380 8558 8400
rect 8578 8380 8592 8400
rect 8550 8342 8592 8380
rect 8642 8400 8686 8442
rect 8642 8380 8654 8400
rect 8674 8380 8686 8400
rect 8642 8342 8686 8380
rect 8763 8400 8805 8442
rect 8763 8380 8771 8400
rect 8791 8380 8805 8400
rect 8763 8342 8805 8380
rect 8855 8400 8899 8442
rect 11598 8499 11642 8541
rect 11692 8561 11734 8599
rect 11692 8541 11706 8561
rect 11726 8541 11734 8561
rect 11692 8499 11734 8541
rect 11811 8561 11855 8599
rect 11811 8541 11823 8561
rect 11843 8541 11855 8561
rect 11811 8499 11855 8541
rect 11905 8561 11947 8599
rect 11905 8541 11919 8561
rect 11939 8541 11947 8561
rect 11905 8499 11947 8541
rect 12019 8561 12063 8599
rect 12019 8541 12031 8561
rect 12051 8541 12063 8561
rect 12019 8499 12063 8541
rect 12113 8561 12155 8599
rect 12113 8541 12127 8561
rect 12147 8541 12155 8561
rect 12113 8499 12155 8541
rect 12229 8561 12271 8599
rect 12229 8541 12237 8561
rect 12257 8541 12271 8561
rect 12229 8499 12271 8541
rect 12321 8568 12366 8599
rect 12321 8561 12365 8568
rect 12321 8541 12333 8561
rect 12353 8541 12365 8561
rect 12321 8499 12365 8541
rect 15201 8552 15245 8590
rect 15201 8532 15213 8552
rect 15233 8532 15245 8552
rect 8855 8380 8867 8400
rect 8887 8380 8899 8400
rect 8855 8342 8899 8380
rect 9180 8396 9224 8438
rect 9180 8376 9192 8396
rect 9212 8376 9224 8396
rect 9180 8369 9224 8376
rect 9179 8338 9224 8369
rect 9274 8396 9316 8438
rect 9274 8376 9288 8396
rect 9308 8376 9316 8396
rect 9274 8338 9316 8376
rect 9390 8396 9432 8438
rect 9390 8376 9398 8396
rect 9418 8376 9432 8396
rect 9390 8338 9432 8376
rect 9482 8396 9526 8438
rect 9482 8376 9494 8396
rect 9514 8376 9526 8396
rect 9482 8338 9526 8376
rect 9598 8396 9640 8438
rect 9598 8376 9606 8396
rect 9626 8376 9640 8396
rect 9598 8338 9640 8376
rect 9690 8396 9734 8438
rect 9690 8376 9702 8396
rect 9722 8376 9734 8396
rect 9690 8338 9734 8376
rect 9811 8396 9853 8438
rect 9811 8376 9819 8396
rect 9839 8376 9853 8396
rect 9811 8338 9853 8376
rect 9903 8396 9947 8438
rect 9903 8376 9915 8396
rect 9935 8376 9947 8396
rect 15201 8490 15245 8532
rect 15295 8552 15337 8590
rect 15295 8532 15309 8552
rect 15329 8532 15337 8552
rect 15295 8490 15337 8532
rect 15414 8552 15458 8590
rect 15414 8532 15426 8552
rect 15446 8532 15458 8552
rect 15414 8490 15458 8532
rect 15508 8552 15550 8590
rect 15508 8532 15522 8552
rect 15542 8532 15550 8552
rect 15508 8490 15550 8532
rect 15622 8552 15666 8590
rect 15622 8532 15634 8552
rect 15654 8532 15666 8552
rect 15622 8490 15666 8532
rect 15716 8552 15758 8590
rect 15716 8532 15730 8552
rect 15750 8532 15758 8552
rect 15716 8490 15758 8532
rect 15832 8552 15874 8590
rect 15832 8532 15840 8552
rect 15860 8532 15874 8552
rect 15832 8490 15874 8532
rect 15924 8559 15969 8590
rect 15924 8552 15968 8559
rect 15924 8532 15936 8552
rect 15956 8532 15968 8552
rect 15924 8490 15968 8532
rect 9903 8338 9947 8376
rect 22563 8565 22607 8603
rect 22563 8545 22575 8565
rect 22595 8545 22607 8565
rect 18840 8394 18884 8436
rect 18840 8374 18852 8394
rect 18872 8374 18884 8394
rect 18840 8367 18884 8374
rect 18839 8336 18884 8367
rect 18934 8394 18976 8436
rect 18934 8374 18948 8394
rect 18968 8374 18976 8394
rect 18934 8336 18976 8374
rect 19050 8394 19092 8436
rect 19050 8374 19058 8394
rect 19078 8374 19092 8394
rect 19050 8336 19092 8374
rect 19142 8394 19186 8436
rect 19142 8374 19154 8394
rect 19174 8374 19186 8394
rect 19142 8336 19186 8374
rect 19258 8394 19300 8436
rect 19258 8374 19266 8394
rect 19286 8374 19300 8394
rect 19258 8336 19300 8374
rect 19350 8394 19394 8436
rect 19350 8374 19362 8394
rect 19382 8374 19394 8394
rect 19350 8336 19394 8374
rect 19471 8394 19513 8436
rect 19471 8374 19479 8394
rect 19499 8374 19513 8394
rect 19471 8336 19513 8374
rect 19563 8394 19607 8436
rect 22563 8503 22607 8545
rect 22657 8565 22699 8603
rect 22657 8545 22671 8565
rect 22691 8545 22699 8565
rect 22657 8503 22699 8545
rect 22776 8565 22820 8603
rect 22776 8545 22788 8565
rect 22808 8545 22820 8565
rect 22776 8503 22820 8545
rect 22870 8565 22912 8603
rect 22870 8545 22884 8565
rect 22904 8545 22912 8565
rect 22870 8503 22912 8545
rect 22984 8565 23028 8603
rect 22984 8545 22996 8565
rect 23016 8545 23028 8565
rect 22984 8503 23028 8545
rect 23078 8565 23120 8603
rect 23078 8545 23092 8565
rect 23112 8545 23120 8565
rect 23078 8503 23120 8545
rect 23194 8565 23236 8603
rect 23194 8545 23202 8565
rect 23222 8545 23236 8565
rect 23194 8503 23236 8545
rect 23286 8572 23331 8603
rect 23286 8565 23330 8572
rect 23286 8545 23298 8565
rect 23318 8545 23330 8565
rect 23286 8503 23330 8545
rect 26166 8556 26210 8594
rect 26166 8536 26178 8556
rect 26198 8536 26210 8556
rect 19563 8374 19575 8394
rect 19595 8374 19607 8394
rect 19563 8336 19607 8374
rect 19888 8390 19932 8432
rect 19888 8370 19900 8390
rect 19920 8370 19932 8390
rect 19888 8363 19932 8370
rect 19887 8332 19932 8363
rect 19982 8390 20024 8432
rect 19982 8370 19996 8390
rect 20016 8370 20024 8390
rect 19982 8332 20024 8370
rect 20098 8390 20140 8432
rect 20098 8370 20106 8390
rect 20126 8370 20140 8390
rect 20098 8332 20140 8370
rect 20190 8390 20234 8432
rect 20190 8370 20202 8390
rect 20222 8370 20234 8390
rect 20190 8332 20234 8370
rect 20306 8390 20348 8432
rect 20306 8370 20314 8390
rect 20334 8370 20348 8390
rect 20306 8332 20348 8370
rect 20398 8390 20442 8432
rect 20398 8370 20410 8390
rect 20430 8370 20442 8390
rect 20398 8332 20442 8370
rect 20519 8390 20561 8432
rect 20519 8370 20527 8390
rect 20547 8370 20561 8390
rect 20519 8332 20561 8370
rect 20611 8390 20655 8432
rect 20611 8370 20623 8390
rect 20643 8370 20655 8390
rect 26166 8494 26210 8536
rect 26260 8556 26302 8594
rect 26260 8536 26274 8556
rect 26294 8536 26302 8556
rect 26260 8494 26302 8536
rect 26379 8556 26423 8594
rect 26379 8536 26391 8556
rect 26411 8536 26423 8556
rect 26379 8494 26423 8536
rect 26473 8556 26515 8594
rect 26473 8536 26487 8556
rect 26507 8536 26515 8556
rect 26473 8494 26515 8536
rect 26587 8556 26631 8594
rect 26587 8536 26599 8556
rect 26619 8536 26631 8556
rect 26587 8494 26631 8536
rect 26681 8556 26723 8594
rect 26681 8536 26695 8556
rect 26715 8536 26723 8556
rect 26681 8494 26723 8536
rect 26797 8556 26839 8594
rect 26797 8536 26805 8556
rect 26825 8536 26839 8556
rect 26797 8494 26839 8536
rect 26889 8563 26934 8594
rect 26889 8556 26933 8563
rect 26889 8536 26901 8556
rect 26921 8536 26933 8556
rect 26889 8494 26933 8536
rect 33271 8559 33315 8597
rect 33271 8539 33283 8559
rect 33303 8539 33315 8559
rect 20611 8332 20655 8370
rect 29805 8398 29849 8440
rect 29805 8378 29817 8398
rect 29837 8378 29849 8398
rect 29805 8371 29849 8378
rect 29804 8340 29849 8371
rect 29899 8398 29941 8440
rect 29899 8378 29913 8398
rect 29933 8378 29941 8398
rect 29899 8340 29941 8378
rect 30015 8398 30057 8440
rect 30015 8378 30023 8398
rect 30043 8378 30057 8398
rect 30015 8340 30057 8378
rect 30107 8398 30151 8440
rect 30107 8378 30119 8398
rect 30139 8378 30151 8398
rect 30107 8340 30151 8378
rect 30223 8398 30265 8440
rect 30223 8378 30231 8398
rect 30251 8378 30265 8398
rect 30223 8340 30265 8378
rect 30315 8398 30359 8440
rect 30315 8378 30327 8398
rect 30347 8378 30359 8398
rect 30315 8340 30359 8378
rect 30436 8398 30478 8440
rect 30436 8378 30444 8398
rect 30464 8378 30478 8398
rect 30436 8340 30478 8378
rect 30528 8398 30572 8440
rect 33271 8497 33315 8539
rect 33365 8559 33407 8597
rect 33365 8539 33379 8559
rect 33399 8539 33407 8559
rect 33365 8497 33407 8539
rect 33484 8559 33528 8597
rect 33484 8539 33496 8559
rect 33516 8539 33528 8559
rect 33484 8497 33528 8539
rect 33578 8559 33620 8597
rect 33578 8539 33592 8559
rect 33612 8539 33620 8559
rect 33578 8497 33620 8539
rect 33692 8559 33736 8597
rect 33692 8539 33704 8559
rect 33724 8539 33736 8559
rect 33692 8497 33736 8539
rect 33786 8559 33828 8597
rect 33786 8539 33800 8559
rect 33820 8539 33828 8559
rect 33786 8497 33828 8539
rect 33902 8559 33944 8597
rect 33902 8539 33910 8559
rect 33930 8539 33944 8559
rect 33902 8497 33944 8539
rect 33994 8566 34039 8597
rect 33994 8559 34038 8566
rect 33994 8539 34006 8559
rect 34026 8539 34038 8559
rect 33994 8497 34038 8539
rect 36874 8550 36918 8588
rect 36874 8530 36886 8550
rect 36906 8530 36918 8550
rect 30528 8378 30540 8398
rect 30560 8378 30572 8398
rect 30528 8340 30572 8378
rect 30853 8394 30897 8436
rect 30853 8374 30865 8394
rect 30885 8374 30897 8394
rect 30853 8367 30897 8374
rect 30852 8336 30897 8367
rect 30947 8394 30989 8436
rect 30947 8374 30961 8394
rect 30981 8374 30989 8394
rect 30947 8336 30989 8374
rect 31063 8394 31105 8436
rect 31063 8374 31071 8394
rect 31091 8374 31105 8394
rect 31063 8336 31105 8374
rect 31155 8394 31199 8436
rect 31155 8374 31167 8394
rect 31187 8374 31199 8394
rect 31155 8336 31199 8374
rect 31271 8394 31313 8436
rect 31271 8374 31279 8394
rect 31299 8374 31313 8394
rect 31271 8336 31313 8374
rect 31363 8394 31407 8436
rect 31363 8374 31375 8394
rect 31395 8374 31407 8394
rect 31363 8336 31407 8374
rect 31484 8394 31526 8436
rect 31484 8374 31492 8394
rect 31512 8374 31526 8394
rect 31484 8336 31526 8374
rect 31576 8394 31620 8436
rect 31576 8374 31588 8394
rect 31608 8374 31620 8394
rect 36874 8488 36918 8530
rect 36968 8550 37010 8588
rect 36968 8530 36982 8550
rect 37002 8530 37010 8550
rect 36968 8488 37010 8530
rect 37087 8550 37131 8588
rect 37087 8530 37099 8550
rect 37119 8530 37131 8550
rect 37087 8488 37131 8530
rect 37181 8550 37223 8588
rect 37181 8530 37195 8550
rect 37215 8530 37223 8550
rect 37181 8488 37223 8530
rect 37295 8550 37339 8588
rect 37295 8530 37307 8550
rect 37327 8530 37339 8550
rect 37295 8488 37339 8530
rect 37389 8550 37431 8588
rect 37389 8530 37403 8550
rect 37423 8530 37431 8550
rect 37389 8488 37431 8530
rect 37505 8550 37547 8588
rect 37505 8530 37513 8550
rect 37533 8530 37547 8550
rect 37505 8488 37547 8530
rect 37597 8557 37642 8588
rect 37597 8550 37641 8557
rect 37597 8530 37609 8550
rect 37629 8530 37641 8550
rect 37597 8488 37641 8530
rect 31576 8336 31620 8374
rect 40513 8392 40557 8434
rect 40513 8372 40525 8392
rect 40545 8372 40557 8392
rect 40513 8365 40557 8372
rect 40512 8334 40557 8365
rect 40607 8392 40649 8434
rect 40607 8372 40621 8392
rect 40641 8372 40649 8392
rect 40607 8334 40649 8372
rect 40723 8392 40765 8434
rect 40723 8372 40731 8392
rect 40751 8372 40765 8392
rect 40723 8334 40765 8372
rect 40815 8392 40859 8434
rect 40815 8372 40827 8392
rect 40847 8372 40859 8392
rect 40815 8334 40859 8372
rect 40931 8392 40973 8434
rect 40931 8372 40939 8392
rect 40959 8372 40973 8392
rect 40931 8334 40973 8372
rect 41023 8392 41067 8434
rect 41023 8372 41035 8392
rect 41055 8372 41067 8392
rect 41023 8334 41067 8372
rect 41144 8392 41186 8434
rect 41144 8372 41152 8392
rect 41172 8372 41186 8392
rect 41144 8334 41186 8372
rect 41236 8392 41280 8434
rect 41236 8372 41248 8392
rect 41268 8372 41280 8392
rect 41236 8334 41280 8372
rect 41561 8388 41605 8430
rect 41561 8368 41573 8388
rect 41593 8368 41605 8388
rect 41561 8361 41605 8368
rect 41560 8330 41605 8361
rect 41655 8388 41697 8430
rect 41655 8368 41669 8388
rect 41689 8368 41697 8388
rect 41655 8330 41697 8368
rect 41771 8388 41813 8430
rect 41771 8368 41779 8388
rect 41799 8368 41813 8388
rect 41771 8330 41813 8368
rect 41863 8388 41907 8430
rect 41863 8368 41875 8388
rect 41895 8368 41907 8388
rect 41863 8330 41907 8368
rect 41979 8388 42021 8430
rect 41979 8368 41987 8388
rect 42007 8368 42021 8388
rect 41979 8330 42021 8368
rect 42071 8388 42115 8430
rect 42071 8368 42083 8388
rect 42103 8368 42115 8388
rect 42071 8330 42115 8368
rect 42192 8388 42234 8430
rect 42192 8368 42200 8388
rect 42220 8368 42234 8388
rect 42192 8330 42234 8368
rect 42284 8388 42328 8430
rect 42284 8368 42296 8388
rect 42316 8368 42328 8388
rect 42284 8330 42328 8368
rect 887 7652 931 7690
rect 887 7632 899 7652
rect 919 7632 931 7652
rect 887 7590 931 7632
rect 981 7652 1023 7690
rect 981 7632 995 7652
rect 1015 7632 1023 7652
rect 981 7590 1023 7632
rect 1100 7652 1144 7690
rect 1100 7632 1112 7652
rect 1132 7632 1144 7652
rect 1100 7590 1144 7632
rect 1194 7652 1236 7690
rect 1194 7632 1208 7652
rect 1228 7632 1236 7652
rect 1194 7590 1236 7632
rect 1308 7652 1352 7690
rect 1308 7632 1320 7652
rect 1340 7632 1352 7652
rect 1308 7590 1352 7632
rect 1402 7652 1444 7690
rect 1402 7632 1416 7652
rect 1436 7632 1444 7652
rect 1402 7590 1444 7632
rect 1518 7652 1560 7690
rect 1518 7632 1526 7652
rect 1546 7632 1560 7652
rect 1518 7590 1560 7632
rect 1610 7659 1655 7690
rect 1610 7652 1654 7659
rect 1610 7632 1622 7652
rect 1642 7632 1654 7652
rect 1610 7590 1654 7632
rect 1935 7648 1979 7686
rect 1935 7628 1947 7648
rect 1967 7628 1979 7648
rect 1935 7586 1979 7628
rect 2029 7648 2071 7686
rect 2029 7628 2043 7648
rect 2063 7628 2071 7648
rect 2029 7586 2071 7628
rect 2148 7648 2192 7686
rect 2148 7628 2160 7648
rect 2180 7628 2192 7648
rect 2148 7586 2192 7628
rect 2242 7648 2284 7686
rect 2242 7628 2256 7648
rect 2276 7628 2284 7648
rect 2242 7586 2284 7628
rect 2356 7648 2400 7686
rect 2356 7628 2368 7648
rect 2388 7628 2400 7648
rect 2356 7586 2400 7628
rect 2450 7648 2492 7686
rect 2450 7628 2464 7648
rect 2484 7628 2492 7648
rect 2450 7586 2492 7628
rect 2566 7648 2608 7686
rect 2566 7628 2574 7648
rect 2594 7628 2608 7648
rect 2566 7586 2608 7628
rect 2658 7655 2703 7686
rect 2658 7648 2702 7655
rect 2658 7628 2670 7648
rect 2690 7628 2702 7648
rect 2658 7586 2702 7628
rect 11595 7646 11639 7684
rect 5574 7490 5618 7532
rect 5574 7470 5586 7490
rect 5606 7470 5618 7490
rect 5574 7463 5618 7470
rect 5573 7432 5618 7463
rect 5668 7490 5710 7532
rect 5668 7470 5682 7490
rect 5702 7470 5710 7490
rect 5668 7432 5710 7470
rect 5784 7490 5826 7532
rect 5784 7470 5792 7490
rect 5812 7470 5826 7490
rect 5784 7432 5826 7470
rect 5876 7490 5920 7532
rect 5876 7470 5888 7490
rect 5908 7470 5920 7490
rect 5876 7432 5920 7470
rect 5992 7490 6034 7532
rect 5992 7470 6000 7490
rect 6020 7470 6034 7490
rect 5992 7432 6034 7470
rect 6084 7490 6128 7532
rect 6084 7470 6096 7490
rect 6116 7470 6128 7490
rect 6084 7432 6128 7470
rect 6205 7490 6247 7532
rect 6205 7470 6213 7490
rect 6233 7470 6247 7490
rect 6205 7432 6247 7470
rect 6297 7490 6341 7532
rect 11595 7626 11607 7646
rect 11627 7626 11639 7646
rect 11595 7584 11639 7626
rect 11689 7646 11731 7684
rect 11689 7626 11703 7646
rect 11723 7626 11731 7646
rect 11689 7584 11731 7626
rect 11808 7646 11852 7684
rect 11808 7626 11820 7646
rect 11840 7626 11852 7646
rect 11808 7584 11852 7626
rect 11902 7646 11944 7684
rect 11902 7626 11916 7646
rect 11936 7626 11944 7646
rect 11902 7584 11944 7626
rect 12016 7646 12060 7684
rect 12016 7626 12028 7646
rect 12048 7626 12060 7646
rect 12016 7584 12060 7626
rect 12110 7646 12152 7684
rect 12110 7626 12124 7646
rect 12144 7626 12152 7646
rect 12110 7584 12152 7626
rect 12226 7646 12268 7684
rect 12226 7626 12234 7646
rect 12254 7626 12268 7646
rect 12226 7584 12268 7626
rect 12318 7653 12363 7684
rect 12318 7646 12362 7653
rect 12318 7626 12330 7646
rect 12350 7626 12362 7646
rect 12318 7584 12362 7626
rect 12643 7642 12687 7680
rect 12643 7622 12655 7642
rect 12675 7622 12687 7642
rect 6297 7470 6309 7490
rect 6329 7470 6341 7490
rect 6297 7432 6341 7470
rect 9177 7481 9221 7523
rect 9177 7461 9189 7481
rect 9209 7461 9221 7481
rect 9177 7454 9221 7461
rect 9176 7423 9221 7454
rect 9271 7481 9313 7523
rect 9271 7461 9285 7481
rect 9305 7461 9313 7481
rect 9271 7423 9313 7461
rect 9387 7481 9429 7523
rect 9387 7461 9395 7481
rect 9415 7461 9429 7481
rect 9387 7423 9429 7461
rect 9479 7481 9523 7523
rect 9479 7461 9491 7481
rect 9511 7461 9523 7481
rect 9479 7423 9523 7461
rect 9595 7481 9637 7523
rect 9595 7461 9603 7481
rect 9623 7461 9637 7481
rect 9595 7423 9637 7461
rect 9687 7481 9731 7523
rect 9687 7461 9699 7481
rect 9719 7461 9731 7481
rect 9687 7423 9731 7461
rect 9808 7481 9850 7523
rect 9808 7461 9816 7481
rect 9836 7461 9850 7481
rect 9808 7423 9850 7461
rect 9900 7481 9944 7523
rect 12643 7580 12687 7622
rect 12737 7642 12779 7680
rect 12737 7622 12751 7642
rect 12771 7622 12779 7642
rect 12737 7580 12779 7622
rect 12856 7642 12900 7680
rect 12856 7622 12868 7642
rect 12888 7622 12900 7642
rect 12856 7580 12900 7622
rect 12950 7642 12992 7680
rect 12950 7622 12964 7642
rect 12984 7622 12992 7642
rect 12950 7580 12992 7622
rect 13064 7642 13108 7680
rect 13064 7622 13076 7642
rect 13096 7622 13108 7642
rect 13064 7580 13108 7622
rect 13158 7642 13200 7680
rect 13158 7622 13172 7642
rect 13192 7622 13200 7642
rect 13158 7580 13200 7622
rect 13274 7642 13316 7680
rect 13274 7622 13282 7642
rect 13302 7622 13316 7642
rect 13274 7580 13316 7622
rect 13366 7649 13411 7680
rect 13366 7642 13410 7649
rect 13366 7622 13378 7642
rect 13398 7622 13410 7642
rect 13366 7580 13410 7622
rect 22560 7650 22604 7688
rect 9900 7461 9912 7481
rect 9932 7461 9944 7481
rect 9900 7423 9944 7461
rect 16282 7484 16326 7526
rect 16282 7464 16294 7484
rect 16314 7464 16326 7484
rect 16282 7457 16326 7464
rect 16281 7426 16326 7457
rect 16376 7484 16418 7526
rect 16376 7464 16390 7484
rect 16410 7464 16418 7484
rect 16376 7426 16418 7464
rect 16492 7484 16534 7526
rect 16492 7464 16500 7484
rect 16520 7464 16534 7484
rect 16492 7426 16534 7464
rect 16584 7484 16628 7526
rect 16584 7464 16596 7484
rect 16616 7464 16628 7484
rect 16584 7426 16628 7464
rect 16700 7484 16742 7526
rect 16700 7464 16708 7484
rect 16728 7464 16742 7484
rect 16700 7426 16742 7464
rect 16792 7484 16836 7526
rect 16792 7464 16804 7484
rect 16824 7464 16836 7484
rect 16792 7426 16836 7464
rect 16913 7484 16955 7526
rect 16913 7464 16921 7484
rect 16941 7464 16955 7484
rect 16913 7426 16955 7464
rect 17005 7484 17049 7526
rect 22560 7630 22572 7650
rect 22592 7630 22604 7650
rect 22560 7588 22604 7630
rect 22654 7650 22696 7688
rect 22654 7630 22668 7650
rect 22688 7630 22696 7650
rect 22654 7588 22696 7630
rect 22773 7650 22817 7688
rect 22773 7630 22785 7650
rect 22805 7630 22817 7650
rect 22773 7588 22817 7630
rect 22867 7650 22909 7688
rect 22867 7630 22881 7650
rect 22901 7630 22909 7650
rect 22867 7588 22909 7630
rect 22981 7650 23025 7688
rect 22981 7630 22993 7650
rect 23013 7630 23025 7650
rect 22981 7588 23025 7630
rect 23075 7650 23117 7688
rect 23075 7630 23089 7650
rect 23109 7630 23117 7650
rect 23075 7588 23117 7630
rect 23191 7650 23233 7688
rect 23191 7630 23199 7650
rect 23219 7630 23233 7650
rect 23191 7588 23233 7630
rect 23283 7657 23328 7688
rect 23283 7650 23327 7657
rect 23283 7630 23295 7650
rect 23315 7630 23327 7650
rect 23283 7588 23327 7630
rect 23608 7646 23652 7684
rect 23608 7626 23620 7646
rect 23640 7626 23652 7646
rect 17005 7464 17017 7484
rect 17037 7464 17049 7484
rect 17005 7426 17049 7464
rect 19885 7475 19929 7517
rect 19885 7455 19897 7475
rect 19917 7455 19929 7475
rect 19885 7448 19929 7455
rect 19884 7417 19929 7448
rect 19979 7475 20021 7517
rect 19979 7455 19993 7475
rect 20013 7455 20021 7475
rect 19979 7417 20021 7455
rect 20095 7475 20137 7517
rect 20095 7455 20103 7475
rect 20123 7455 20137 7475
rect 20095 7417 20137 7455
rect 20187 7475 20231 7517
rect 20187 7455 20199 7475
rect 20219 7455 20231 7475
rect 20187 7417 20231 7455
rect 20303 7475 20345 7517
rect 20303 7455 20311 7475
rect 20331 7455 20345 7475
rect 20303 7417 20345 7455
rect 20395 7475 20439 7517
rect 20395 7455 20407 7475
rect 20427 7455 20439 7475
rect 20395 7417 20439 7455
rect 20516 7475 20558 7517
rect 20516 7455 20524 7475
rect 20544 7455 20558 7475
rect 20516 7417 20558 7455
rect 20608 7475 20652 7517
rect 23608 7584 23652 7626
rect 23702 7646 23744 7684
rect 23702 7626 23716 7646
rect 23736 7626 23744 7646
rect 23702 7584 23744 7626
rect 23821 7646 23865 7684
rect 23821 7626 23833 7646
rect 23853 7626 23865 7646
rect 23821 7584 23865 7626
rect 23915 7646 23957 7684
rect 23915 7626 23929 7646
rect 23949 7626 23957 7646
rect 23915 7584 23957 7626
rect 24029 7646 24073 7684
rect 24029 7626 24041 7646
rect 24061 7626 24073 7646
rect 24029 7584 24073 7626
rect 24123 7646 24165 7684
rect 24123 7626 24137 7646
rect 24157 7626 24165 7646
rect 24123 7584 24165 7626
rect 24239 7646 24281 7684
rect 24239 7626 24247 7646
rect 24267 7626 24281 7646
rect 24239 7584 24281 7626
rect 24331 7653 24376 7684
rect 24331 7646 24375 7653
rect 24331 7626 24343 7646
rect 24363 7626 24375 7646
rect 24331 7584 24375 7626
rect 20608 7455 20620 7475
rect 20640 7455 20652 7475
rect 20608 7417 20652 7455
rect 33268 7644 33312 7682
rect 27247 7488 27291 7530
rect 27247 7468 27259 7488
rect 27279 7468 27291 7488
rect 27247 7461 27291 7468
rect 27246 7430 27291 7461
rect 27341 7488 27383 7530
rect 27341 7468 27355 7488
rect 27375 7468 27383 7488
rect 27341 7430 27383 7468
rect 27457 7488 27499 7530
rect 27457 7468 27465 7488
rect 27485 7468 27499 7488
rect 27457 7430 27499 7468
rect 27549 7488 27593 7530
rect 27549 7468 27561 7488
rect 27581 7468 27593 7488
rect 27549 7430 27593 7468
rect 27665 7488 27707 7530
rect 27665 7468 27673 7488
rect 27693 7468 27707 7488
rect 27665 7430 27707 7468
rect 27757 7488 27801 7530
rect 27757 7468 27769 7488
rect 27789 7468 27801 7488
rect 27757 7430 27801 7468
rect 27878 7488 27920 7530
rect 27878 7468 27886 7488
rect 27906 7468 27920 7488
rect 27878 7430 27920 7468
rect 27970 7488 28014 7530
rect 33268 7624 33280 7644
rect 33300 7624 33312 7644
rect 33268 7582 33312 7624
rect 33362 7644 33404 7682
rect 33362 7624 33376 7644
rect 33396 7624 33404 7644
rect 33362 7582 33404 7624
rect 33481 7644 33525 7682
rect 33481 7624 33493 7644
rect 33513 7624 33525 7644
rect 33481 7582 33525 7624
rect 33575 7644 33617 7682
rect 33575 7624 33589 7644
rect 33609 7624 33617 7644
rect 33575 7582 33617 7624
rect 33689 7644 33733 7682
rect 33689 7624 33701 7644
rect 33721 7624 33733 7644
rect 33689 7582 33733 7624
rect 33783 7644 33825 7682
rect 33783 7624 33797 7644
rect 33817 7624 33825 7644
rect 33783 7582 33825 7624
rect 33899 7644 33941 7682
rect 33899 7624 33907 7644
rect 33927 7624 33941 7644
rect 33899 7582 33941 7624
rect 33991 7651 34036 7682
rect 33991 7644 34035 7651
rect 33991 7624 34003 7644
rect 34023 7624 34035 7644
rect 33991 7582 34035 7624
rect 34316 7640 34360 7678
rect 34316 7620 34328 7640
rect 34348 7620 34360 7640
rect 27970 7468 27982 7488
rect 28002 7468 28014 7488
rect 27970 7430 28014 7468
rect 30850 7479 30894 7521
rect 30850 7459 30862 7479
rect 30882 7459 30894 7479
rect 30850 7452 30894 7459
rect 30849 7421 30894 7452
rect 30944 7479 30986 7521
rect 30944 7459 30958 7479
rect 30978 7459 30986 7479
rect 30944 7421 30986 7459
rect 31060 7479 31102 7521
rect 31060 7459 31068 7479
rect 31088 7459 31102 7479
rect 31060 7421 31102 7459
rect 31152 7479 31196 7521
rect 31152 7459 31164 7479
rect 31184 7459 31196 7479
rect 31152 7421 31196 7459
rect 31268 7479 31310 7521
rect 31268 7459 31276 7479
rect 31296 7459 31310 7479
rect 31268 7421 31310 7459
rect 31360 7479 31404 7521
rect 31360 7459 31372 7479
rect 31392 7459 31404 7479
rect 31360 7421 31404 7459
rect 31481 7479 31523 7521
rect 31481 7459 31489 7479
rect 31509 7459 31523 7479
rect 31481 7421 31523 7459
rect 31573 7479 31617 7521
rect 34316 7578 34360 7620
rect 34410 7640 34452 7678
rect 34410 7620 34424 7640
rect 34444 7620 34452 7640
rect 34410 7578 34452 7620
rect 34529 7640 34573 7678
rect 34529 7620 34541 7640
rect 34561 7620 34573 7640
rect 34529 7578 34573 7620
rect 34623 7640 34665 7678
rect 34623 7620 34637 7640
rect 34657 7620 34665 7640
rect 34623 7578 34665 7620
rect 34737 7640 34781 7678
rect 34737 7620 34749 7640
rect 34769 7620 34781 7640
rect 34737 7578 34781 7620
rect 34831 7640 34873 7678
rect 34831 7620 34845 7640
rect 34865 7620 34873 7640
rect 34831 7578 34873 7620
rect 34947 7640 34989 7678
rect 34947 7620 34955 7640
rect 34975 7620 34989 7640
rect 34947 7578 34989 7620
rect 35039 7647 35084 7678
rect 35039 7640 35083 7647
rect 35039 7620 35051 7640
rect 35071 7620 35083 7640
rect 35039 7578 35083 7620
rect 31573 7459 31585 7479
rect 31605 7459 31617 7479
rect 31573 7421 31617 7459
rect 37955 7482 37999 7524
rect 37955 7462 37967 7482
rect 37987 7462 37999 7482
rect 37955 7455 37999 7462
rect 37954 7424 37999 7455
rect 38049 7482 38091 7524
rect 38049 7462 38063 7482
rect 38083 7462 38091 7482
rect 38049 7424 38091 7462
rect 38165 7482 38207 7524
rect 38165 7462 38173 7482
rect 38193 7462 38207 7482
rect 38165 7424 38207 7462
rect 38257 7482 38301 7524
rect 38257 7462 38269 7482
rect 38289 7462 38301 7482
rect 38257 7424 38301 7462
rect 38373 7482 38415 7524
rect 38373 7462 38381 7482
rect 38401 7462 38415 7482
rect 38373 7424 38415 7462
rect 38465 7482 38509 7524
rect 38465 7462 38477 7482
rect 38497 7462 38509 7482
rect 38465 7424 38509 7462
rect 38586 7482 38628 7524
rect 38586 7462 38594 7482
rect 38614 7462 38628 7482
rect 38586 7424 38628 7462
rect 38678 7482 38722 7524
rect 38678 7462 38690 7482
rect 38710 7462 38722 7482
rect 38678 7424 38722 7462
rect 41558 7473 41602 7515
rect 41558 7453 41570 7473
rect 41590 7453 41602 7473
rect 41558 7446 41602 7453
rect 41557 7415 41602 7446
rect 41652 7473 41694 7515
rect 41652 7453 41666 7473
rect 41686 7453 41694 7473
rect 41652 7415 41694 7453
rect 41768 7473 41810 7515
rect 41768 7453 41776 7473
rect 41796 7453 41810 7473
rect 41768 7415 41810 7453
rect 41860 7473 41904 7515
rect 41860 7453 41872 7473
rect 41892 7453 41904 7473
rect 41860 7415 41904 7453
rect 41976 7473 42018 7515
rect 41976 7453 41984 7473
rect 42004 7453 42018 7473
rect 41976 7415 42018 7453
rect 42068 7473 42112 7515
rect 42068 7453 42080 7473
rect 42100 7453 42112 7473
rect 42068 7415 42112 7453
rect 42189 7473 42231 7515
rect 42189 7453 42197 7473
rect 42217 7453 42231 7473
rect 42189 7415 42231 7453
rect 42281 7473 42325 7515
rect 42281 7453 42293 7473
rect 42313 7453 42325 7473
rect 42281 7415 42325 7453
rect 887 6973 931 7011
rect 887 6953 899 6973
rect 919 6953 931 6973
rect 887 6911 931 6953
rect 981 6973 1023 7011
rect 981 6953 995 6973
rect 1015 6953 1023 6973
rect 981 6911 1023 6953
rect 1100 6973 1144 7011
rect 1100 6953 1112 6973
rect 1132 6953 1144 6973
rect 1100 6911 1144 6953
rect 1194 6973 1236 7011
rect 1194 6953 1208 6973
rect 1228 6953 1236 6973
rect 1194 6911 1236 6953
rect 1308 6973 1352 7011
rect 1308 6953 1320 6973
rect 1340 6953 1352 6973
rect 1308 6911 1352 6953
rect 1402 6973 1444 7011
rect 1402 6953 1416 6973
rect 1436 6953 1444 6973
rect 1402 6911 1444 6953
rect 1518 6973 1560 7011
rect 1518 6953 1526 6973
rect 1546 6953 1560 6973
rect 1518 6911 1560 6953
rect 1610 6980 1655 7011
rect 1610 6973 1654 6980
rect 1610 6953 1622 6973
rect 1642 6953 1654 6973
rect 1610 6911 1654 6953
rect 3382 6968 3426 7006
rect 3382 6948 3394 6968
rect 3414 6948 3426 6968
rect 3382 6906 3426 6948
rect 3476 6968 3518 7006
rect 3476 6948 3490 6968
rect 3510 6948 3518 6968
rect 3476 6906 3518 6948
rect 3595 6968 3639 7006
rect 3595 6948 3607 6968
rect 3627 6948 3639 6968
rect 3595 6906 3639 6948
rect 3689 6968 3731 7006
rect 3689 6948 3703 6968
rect 3723 6948 3731 6968
rect 3689 6906 3731 6948
rect 3803 6968 3847 7006
rect 3803 6948 3815 6968
rect 3835 6948 3847 6968
rect 3803 6906 3847 6948
rect 3897 6968 3939 7006
rect 3897 6948 3911 6968
rect 3931 6948 3939 6968
rect 3897 6906 3939 6948
rect 4013 6968 4055 7006
rect 4013 6948 4021 6968
rect 4041 6948 4055 6968
rect 4013 6906 4055 6948
rect 4105 6975 4150 7006
rect 4105 6968 4149 6975
rect 4105 6948 4117 6968
rect 4137 6948 4149 6968
rect 4105 6906 4149 6948
rect 11595 6967 11639 7005
rect 11595 6947 11607 6967
rect 11627 6947 11639 6967
rect 8129 6806 8173 6848
rect 8129 6786 8141 6806
rect 8161 6786 8173 6806
rect 8129 6779 8173 6786
rect 8128 6748 8173 6779
rect 8223 6806 8265 6848
rect 8223 6786 8237 6806
rect 8257 6786 8265 6806
rect 8223 6748 8265 6786
rect 8339 6806 8381 6848
rect 8339 6786 8347 6806
rect 8367 6786 8381 6806
rect 8339 6748 8381 6786
rect 8431 6806 8475 6848
rect 8431 6786 8443 6806
rect 8463 6786 8475 6806
rect 8431 6748 8475 6786
rect 8547 6806 8589 6848
rect 8547 6786 8555 6806
rect 8575 6786 8589 6806
rect 8547 6748 8589 6786
rect 8639 6806 8683 6848
rect 8639 6786 8651 6806
rect 8671 6786 8683 6806
rect 8639 6748 8683 6786
rect 8760 6806 8802 6848
rect 8760 6786 8768 6806
rect 8788 6786 8802 6806
rect 8760 6748 8802 6786
rect 8852 6806 8896 6848
rect 11595 6905 11639 6947
rect 11689 6967 11731 7005
rect 11689 6947 11703 6967
rect 11723 6947 11731 6967
rect 11689 6905 11731 6947
rect 11808 6967 11852 7005
rect 11808 6947 11820 6967
rect 11840 6947 11852 6967
rect 11808 6905 11852 6947
rect 11902 6967 11944 7005
rect 11902 6947 11916 6967
rect 11936 6947 11944 6967
rect 11902 6905 11944 6947
rect 12016 6967 12060 7005
rect 12016 6947 12028 6967
rect 12048 6947 12060 6967
rect 12016 6905 12060 6947
rect 12110 6967 12152 7005
rect 12110 6947 12124 6967
rect 12144 6947 12152 6967
rect 12110 6905 12152 6947
rect 12226 6967 12268 7005
rect 12226 6947 12234 6967
rect 12254 6947 12268 6967
rect 12226 6905 12268 6947
rect 12318 6974 12363 7005
rect 12318 6967 12362 6974
rect 12318 6947 12330 6967
rect 12350 6947 12362 6967
rect 12318 6905 12362 6947
rect 14090 6962 14134 7000
rect 14090 6942 14102 6962
rect 14122 6942 14134 6962
rect 8852 6786 8864 6806
rect 8884 6786 8896 6806
rect 8852 6748 8896 6786
rect 9177 6802 9221 6844
rect 9177 6782 9189 6802
rect 9209 6782 9221 6802
rect 9177 6775 9221 6782
rect 9176 6744 9221 6775
rect 9271 6802 9313 6844
rect 9271 6782 9285 6802
rect 9305 6782 9313 6802
rect 9271 6744 9313 6782
rect 9387 6802 9429 6844
rect 9387 6782 9395 6802
rect 9415 6782 9429 6802
rect 9387 6744 9429 6782
rect 9479 6802 9523 6844
rect 9479 6782 9491 6802
rect 9511 6782 9523 6802
rect 9479 6744 9523 6782
rect 9595 6802 9637 6844
rect 9595 6782 9603 6802
rect 9623 6782 9637 6802
rect 9595 6744 9637 6782
rect 9687 6802 9731 6844
rect 9687 6782 9699 6802
rect 9719 6782 9731 6802
rect 9687 6744 9731 6782
rect 9808 6802 9850 6844
rect 9808 6782 9816 6802
rect 9836 6782 9850 6802
rect 9808 6744 9850 6782
rect 9900 6802 9944 6844
rect 9900 6782 9912 6802
rect 9932 6782 9944 6802
rect 14090 6900 14134 6942
rect 14184 6962 14226 7000
rect 14184 6942 14198 6962
rect 14218 6942 14226 6962
rect 14184 6900 14226 6942
rect 14303 6962 14347 7000
rect 14303 6942 14315 6962
rect 14335 6942 14347 6962
rect 14303 6900 14347 6942
rect 14397 6962 14439 7000
rect 14397 6942 14411 6962
rect 14431 6942 14439 6962
rect 14397 6900 14439 6942
rect 14511 6962 14555 7000
rect 14511 6942 14523 6962
rect 14543 6942 14555 6962
rect 14511 6900 14555 6942
rect 14605 6962 14647 7000
rect 14605 6942 14619 6962
rect 14639 6942 14647 6962
rect 14605 6900 14647 6942
rect 14721 6962 14763 7000
rect 14721 6942 14729 6962
rect 14749 6942 14763 6962
rect 14721 6900 14763 6942
rect 14813 6969 14858 7000
rect 14813 6962 14857 6969
rect 14813 6942 14825 6962
rect 14845 6942 14857 6962
rect 14813 6900 14857 6942
rect 9900 6744 9944 6782
rect 22560 6971 22604 7009
rect 22560 6951 22572 6971
rect 22592 6951 22604 6971
rect 18837 6800 18881 6842
rect 18837 6780 18849 6800
rect 18869 6780 18881 6800
rect 18837 6773 18881 6780
rect 18836 6742 18881 6773
rect 18931 6800 18973 6842
rect 18931 6780 18945 6800
rect 18965 6780 18973 6800
rect 18931 6742 18973 6780
rect 19047 6800 19089 6842
rect 19047 6780 19055 6800
rect 19075 6780 19089 6800
rect 19047 6742 19089 6780
rect 19139 6800 19183 6842
rect 19139 6780 19151 6800
rect 19171 6780 19183 6800
rect 19139 6742 19183 6780
rect 19255 6800 19297 6842
rect 19255 6780 19263 6800
rect 19283 6780 19297 6800
rect 19255 6742 19297 6780
rect 19347 6800 19391 6842
rect 19347 6780 19359 6800
rect 19379 6780 19391 6800
rect 19347 6742 19391 6780
rect 19468 6800 19510 6842
rect 19468 6780 19476 6800
rect 19496 6780 19510 6800
rect 19468 6742 19510 6780
rect 19560 6800 19604 6842
rect 22560 6909 22604 6951
rect 22654 6971 22696 7009
rect 22654 6951 22668 6971
rect 22688 6951 22696 6971
rect 22654 6909 22696 6951
rect 22773 6971 22817 7009
rect 22773 6951 22785 6971
rect 22805 6951 22817 6971
rect 22773 6909 22817 6951
rect 22867 6971 22909 7009
rect 22867 6951 22881 6971
rect 22901 6951 22909 6971
rect 22867 6909 22909 6951
rect 22981 6971 23025 7009
rect 22981 6951 22993 6971
rect 23013 6951 23025 6971
rect 22981 6909 23025 6951
rect 23075 6971 23117 7009
rect 23075 6951 23089 6971
rect 23109 6951 23117 6971
rect 23075 6909 23117 6951
rect 23191 6971 23233 7009
rect 23191 6951 23199 6971
rect 23219 6951 23233 6971
rect 23191 6909 23233 6951
rect 23283 6978 23328 7009
rect 23283 6971 23327 6978
rect 23283 6951 23295 6971
rect 23315 6951 23327 6971
rect 23283 6909 23327 6951
rect 25055 6966 25099 7004
rect 25055 6946 25067 6966
rect 25087 6946 25099 6966
rect 19560 6780 19572 6800
rect 19592 6780 19604 6800
rect 19560 6742 19604 6780
rect 19885 6796 19929 6838
rect 19885 6776 19897 6796
rect 19917 6776 19929 6796
rect 19885 6769 19929 6776
rect 19884 6738 19929 6769
rect 19979 6796 20021 6838
rect 19979 6776 19993 6796
rect 20013 6776 20021 6796
rect 19979 6738 20021 6776
rect 20095 6796 20137 6838
rect 20095 6776 20103 6796
rect 20123 6776 20137 6796
rect 20095 6738 20137 6776
rect 20187 6796 20231 6838
rect 20187 6776 20199 6796
rect 20219 6776 20231 6796
rect 20187 6738 20231 6776
rect 20303 6796 20345 6838
rect 20303 6776 20311 6796
rect 20331 6776 20345 6796
rect 20303 6738 20345 6776
rect 20395 6796 20439 6838
rect 20395 6776 20407 6796
rect 20427 6776 20439 6796
rect 20395 6738 20439 6776
rect 20516 6796 20558 6838
rect 20516 6776 20524 6796
rect 20544 6776 20558 6796
rect 20516 6738 20558 6776
rect 20608 6796 20652 6838
rect 20608 6776 20620 6796
rect 20640 6776 20652 6796
rect 25055 6904 25099 6946
rect 25149 6966 25191 7004
rect 25149 6946 25163 6966
rect 25183 6946 25191 6966
rect 25149 6904 25191 6946
rect 25268 6966 25312 7004
rect 25268 6946 25280 6966
rect 25300 6946 25312 6966
rect 25268 6904 25312 6946
rect 25362 6966 25404 7004
rect 25362 6946 25376 6966
rect 25396 6946 25404 6966
rect 25362 6904 25404 6946
rect 25476 6966 25520 7004
rect 25476 6946 25488 6966
rect 25508 6946 25520 6966
rect 25476 6904 25520 6946
rect 25570 6966 25612 7004
rect 25570 6946 25584 6966
rect 25604 6946 25612 6966
rect 25570 6904 25612 6946
rect 25686 6966 25728 7004
rect 25686 6946 25694 6966
rect 25714 6946 25728 6966
rect 25686 6904 25728 6946
rect 25778 6973 25823 7004
rect 25778 6966 25822 6973
rect 25778 6946 25790 6966
rect 25810 6946 25822 6966
rect 25778 6904 25822 6946
rect 33268 6965 33312 7003
rect 33268 6945 33280 6965
rect 33300 6945 33312 6965
rect 20608 6738 20652 6776
rect 29802 6804 29846 6846
rect 29802 6784 29814 6804
rect 29834 6784 29846 6804
rect 29802 6777 29846 6784
rect 29801 6746 29846 6777
rect 29896 6804 29938 6846
rect 29896 6784 29910 6804
rect 29930 6784 29938 6804
rect 29896 6746 29938 6784
rect 30012 6804 30054 6846
rect 30012 6784 30020 6804
rect 30040 6784 30054 6804
rect 30012 6746 30054 6784
rect 30104 6804 30148 6846
rect 30104 6784 30116 6804
rect 30136 6784 30148 6804
rect 30104 6746 30148 6784
rect 30220 6804 30262 6846
rect 30220 6784 30228 6804
rect 30248 6784 30262 6804
rect 30220 6746 30262 6784
rect 30312 6804 30356 6846
rect 30312 6784 30324 6804
rect 30344 6784 30356 6804
rect 30312 6746 30356 6784
rect 30433 6804 30475 6846
rect 30433 6784 30441 6804
rect 30461 6784 30475 6804
rect 30433 6746 30475 6784
rect 30525 6804 30569 6846
rect 33268 6903 33312 6945
rect 33362 6965 33404 7003
rect 33362 6945 33376 6965
rect 33396 6945 33404 6965
rect 33362 6903 33404 6945
rect 33481 6965 33525 7003
rect 33481 6945 33493 6965
rect 33513 6945 33525 6965
rect 33481 6903 33525 6945
rect 33575 6965 33617 7003
rect 33575 6945 33589 6965
rect 33609 6945 33617 6965
rect 33575 6903 33617 6945
rect 33689 6965 33733 7003
rect 33689 6945 33701 6965
rect 33721 6945 33733 6965
rect 33689 6903 33733 6945
rect 33783 6965 33825 7003
rect 33783 6945 33797 6965
rect 33817 6945 33825 6965
rect 33783 6903 33825 6945
rect 33899 6965 33941 7003
rect 33899 6945 33907 6965
rect 33927 6945 33941 6965
rect 33899 6903 33941 6945
rect 33991 6972 34036 7003
rect 33991 6965 34035 6972
rect 33991 6945 34003 6965
rect 34023 6945 34035 6965
rect 33991 6903 34035 6945
rect 35763 6960 35807 6998
rect 35763 6940 35775 6960
rect 35795 6940 35807 6960
rect 30525 6784 30537 6804
rect 30557 6784 30569 6804
rect 30525 6746 30569 6784
rect 30850 6800 30894 6842
rect 30850 6780 30862 6800
rect 30882 6780 30894 6800
rect 30850 6773 30894 6780
rect 30849 6742 30894 6773
rect 30944 6800 30986 6842
rect 30944 6780 30958 6800
rect 30978 6780 30986 6800
rect 30944 6742 30986 6780
rect 31060 6800 31102 6842
rect 31060 6780 31068 6800
rect 31088 6780 31102 6800
rect 31060 6742 31102 6780
rect 31152 6800 31196 6842
rect 31152 6780 31164 6800
rect 31184 6780 31196 6800
rect 31152 6742 31196 6780
rect 31268 6800 31310 6842
rect 31268 6780 31276 6800
rect 31296 6780 31310 6800
rect 31268 6742 31310 6780
rect 31360 6800 31404 6842
rect 31360 6780 31372 6800
rect 31392 6780 31404 6800
rect 31360 6742 31404 6780
rect 31481 6800 31523 6842
rect 31481 6780 31489 6800
rect 31509 6780 31523 6800
rect 31481 6742 31523 6780
rect 31573 6800 31617 6842
rect 31573 6780 31585 6800
rect 31605 6780 31617 6800
rect 35763 6898 35807 6940
rect 35857 6960 35899 6998
rect 35857 6940 35871 6960
rect 35891 6940 35899 6960
rect 35857 6898 35899 6940
rect 35976 6960 36020 6998
rect 35976 6940 35988 6960
rect 36008 6940 36020 6960
rect 35976 6898 36020 6940
rect 36070 6960 36112 6998
rect 36070 6940 36084 6960
rect 36104 6940 36112 6960
rect 36070 6898 36112 6940
rect 36184 6960 36228 6998
rect 36184 6940 36196 6960
rect 36216 6940 36228 6960
rect 36184 6898 36228 6940
rect 36278 6960 36320 6998
rect 36278 6940 36292 6960
rect 36312 6940 36320 6960
rect 36278 6898 36320 6940
rect 36394 6960 36436 6998
rect 36394 6940 36402 6960
rect 36422 6940 36436 6960
rect 36394 6898 36436 6940
rect 36486 6967 36531 6998
rect 36486 6960 36530 6967
rect 36486 6940 36498 6960
rect 36518 6940 36530 6960
rect 36486 6898 36530 6940
rect 31573 6742 31617 6780
rect 40510 6798 40554 6840
rect 40510 6778 40522 6798
rect 40542 6778 40554 6798
rect 40510 6771 40554 6778
rect 40509 6740 40554 6771
rect 40604 6798 40646 6840
rect 40604 6778 40618 6798
rect 40638 6778 40646 6798
rect 40604 6740 40646 6778
rect 40720 6798 40762 6840
rect 40720 6778 40728 6798
rect 40748 6778 40762 6798
rect 40720 6740 40762 6778
rect 40812 6798 40856 6840
rect 40812 6778 40824 6798
rect 40844 6778 40856 6798
rect 40812 6740 40856 6778
rect 40928 6798 40970 6840
rect 40928 6778 40936 6798
rect 40956 6778 40970 6798
rect 40928 6740 40970 6778
rect 41020 6798 41064 6840
rect 41020 6778 41032 6798
rect 41052 6778 41064 6798
rect 41020 6740 41064 6778
rect 41141 6798 41183 6840
rect 41141 6778 41149 6798
rect 41169 6778 41183 6798
rect 41141 6740 41183 6778
rect 41233 6798 41277 6840
rect 41233 6778 41245 6798
rect 41265 6778 41277 6798
rect 41233 6740 41277 6778
rect 41558 6794 41602 6836
rect 41558 6774 41570 6794
rect 41590 6774 41602 6794
rect 41558 6767 41602 6774
rect 41557 6736 41602 6767
rect 41652 6794 41694 6836
rect 41652 6774 41666 6794
rect 41686 6774 41694 6794
rect 41652 6736 41694 6774
rect 41768 6794 41810 6836
rect 41768 6774 41776 6794
rect 41796 6774 41810 6794
rect 41768 6736 41810 6774
rect 41860 6794 41904 6836
rect 41860 6774 41872 6794
rect 41892 6774 41904 6794
rect 41860 6736 41904 6774
rect 41976 6794 42018 6836
rect 41976 6774 41984 6794
rect 42004 6774 42018 6794
rect 41976 6736 42018 6774
rect 42068 6794 42112 6836
rect 42068 6774 42080 6794
rect 42100 6774 42112 6794
rect 42068 6736 42112 6774
rect 42189 6794 42231 6836
rect 42189 6774 42197 6794
rect 42217 6774 42231 6794
rect 42189 6736 42231 6774
rect 42281 6794 42325 6836
rect 42281 6774 42293 6794
rect 42313 6774 42325 6794
rect 42281 6736 42325 6774
rect 887 6205 931 6243
rect 887 6185 899 6205
rect 919 6185 931 6205
rect 887 6143 931 6185
rect 981 6205 1023 6243
rect 981 6185 995 6205
rect 1015 6185 1023 6205
rect 981 6143 1023 6185
rect 1100 6205 1144 6243
rect 1100 6185 1112 6205
rect 1132 6185 1144 6205
rect 1100 6143 1144 6185
rect 1194 6205 1236 6243
rect 1194 6185 1208 6205
rect 1228 6185 1236 6205
rect 1194 6143 1236 6185
rect 1308 6205 1352 6243
rect 1308 6185 1320 6205
rect 1340 6185 1352 6205
rect 1308 6143 1352 6185
rect 1402 6205 1444 6243
rect 1402 6185 1416 6205
rect 1436 6185 1444 6205
rect 1402 6143 1444 6185
rect 1518 6205 1560 6243
rect 1518 6185 1526 6205
rect 1546 6185 1560 6205
rect 1518 6143 1560 6185
rect 1610 6212 1655 6243
rect 1610 6205 1654 6212
rect 1610 6185 1622 6205
rect 1642 6185 1654 6205
rect 1610 6143 1654 6185
rect 1935 6201 1979 6239
rect 1935 6181 1947 6201
rect 1967 6181 1979 6201
rect 1935 6139 1979 6181
rect 2029 6201 2071 6239
rect 2029 6181 2043 6201
rect 2063 6181 2071 6201
rect 2029 6139 2071 6181
rect 2148 6201 2192 6239
rect 2148 6181 2160 6201
rect 2180 6181 2192 6201
rect 2148 6139 2192 6181
rect 2242 6201 2284 6239
rect 2242 6181 2256 6201
rect 2276 6181 2284 6201
rect 2242 6139 2284 6181
rect 2356 6201 2400 6239
rect 2356 6181 2368 6201
rect 2388 6181 2400 6201
rect 2356 6139 2400 6181
rect 2450 6201 2492 6239
rect 2450 6181 2464 6201
rect 2484 6181 2492 6201
rect 2450 6139 2492 6181
rect 2566 6201 2608 6239
rect 2566 6181 2574 6201
rect 2594 6181 2608 6201
rect 2566 6139 2608 6181
rect 2658 6208 2703 6239
rect 2658 6201 2702 6208
rect 2658 6181 2670 6201
rect 2690 6181 2702 6201
rect 2658 6139 2702 6181
rect 11595 6199 11639 6237
rect 6682 6039 6726 6081
rect 6682 6019 6694 6039
rect 6714 6019 6726 6039
rect 6682 6012 6726 6019
rect 6681 5981 6726 6012
rect 6776 6039 6818 6081
rect 6776 6019 6790 6039
rect 6810 6019 6818 6039
rect 6776 5981 6818 6019
rect 6892 6039 6934 6081
rect 6892 6019 6900 6039
rect 6920 6019 6934 6039
rect 6892 5981 6934 6019
rect 6984 6039 7028 6081
rect 6984 6019 6996 6039
rect 7016 6019 7028 6039
rect 6984 5981 7028 6019
rect 7100 6039 7142 6081
rect 7100 6019 7108 6039
rect 7128 6019 7142 6039
rect 7100 5981 7142 6019
rect 7192 6039 7236 6081
rect 7192 6019 7204 6039
rect 7224 6019 7236 6039
rect 7192 5981 7236 6019
rect 7313 6039 7355 6081
rect 7313 6019 7321 6039
rect 7341 6019 7355 6039
rect 7313 5981 7355 6019
rect 7405 6039 7449 6081
rect 11595 6179 11607 6199
rect 11627 6179 11639 6199
rect 11595 6137 11639 6179
rect 11689 6199 11731 6237
rect 11689 6179 11703 6199
rect 11723 6179 11731 6199
rect 11689 6137 11731 6179
rect 11808 6199 11852 6237
rect 11808 6179 11820 6199
rect 11840 6179 11852 6199
rect 11808 6137 11852 6179
rect 11902 6199 11944 6237
rect 11902 6179 11916 6199
rect 11936 6179 11944 6199
rect 11902 6137 11944 6179
rect 12016 6199 12060 6237
rect 12016 6179 12028 6199
rect 12048 6179 12060 6199
rect 12016 6137 12060 6179
rect 12110 6199 12152 6237
rect 12110 6179 12124 6199
rect 12144 6179 12152 6199
rect 12110 6137 12152 6179
rect 12226 6199 12268 6237
rect 12226 6179 12234 6199
rect 12254 6179 12268 6199
rect 12226 6137 12268 6179
rect 12318 6206 12363 6237
rect 12318 6199 12362 6206
rect 12318 6179 12330 6199
rect 12350 6179 12362 6199
rect 12318 6137 12362 6179
rect 12643 6195 12687 6233
rect 12643 6175 12655 6195
rect 12675 6175 12687 6195
rect 7405 6019 7417 6039
rect 7437 6019 7449 6039
rect 7405 5981 7449 6019
rect 9177 6034 9221 6076
rect 9177 6014 9189 6034
rect 9209 6014 9221 6034
rect 9177 6007 9221 6014
rect 9176 5976 9221 6007
rect 9271 6034 9313 6076
rect 9271 6014 9285 6034
rect 9305 6014 9313 6034
rect 9271 5976 9313 6014
rect 9387 6034 9429 6076
rect 9387 6014 9395 6034
rect 9415 6014 9429 6034
rect 9387 5976 9429 6014
rect 9479 6034 9523 6076
rect 9479 6014 9491 6034
rect 9511 6014 9523 6034
rect 9479 5976 9523 6014
rect 9595 6034 9637 6076
rect 9595 6014 9603 6034
rect 9623 6014 9637 6034
rect 9595 5976 9637 6014
rect 9687 6034 9731 6076
rect 9687 6014 9699 6034
rect 9719 6014 9731 6034
rect 9687 5976 9731 6014
rect 9808 6034 9850 6076
rect 9808 6014 9816 6034
rect 9836 6014 9850 6034
rect 9808 5976 9850 6014
rect 9900 6034 9944 6076
rect 12643 6133 12687 6175
rect 12737 6195 12779 6233
rect 12737 6175 12751 6195
rect 12771 6175 12779 6195
rect 12737 6133 12779 6175
rect 12856 6195 12900 6233
rect 12856 6175 12868 6195
rect 12888 6175 12900 6195
rect 12856 6133 12900 6175
rect 12950 6195 12992 6233
rect 12950 6175 12964 6195
rect 12984 6175 12992 6195
rect 12950 6133 12992 6175
rect 13064 6195 13108 6233
rect 13064 6175 13076 6195
rect 13096 6175 13108 6195
rect 13064 6133 13108 6175
rect 13158 6195 13200 6233
rect 13158 6175 13172 6195
rect 13192 6175 13200 6195
rect 13158 6133 13200 6175
rect 13274 6195 13316 6233
rect 13274 6175 13282 6195
rect 13302 6175 13316 6195
rect 13274 6133 13316 6175
rect 13366 6202 13411 6233
rect 13366 6195 13410 6202
rect 13366 6175 13378 6195
rect 13398 6175 13410 6195
rect 13366 6133 13410 6175
rect 22560 6203 22604 6241
rect 9900 6014 9912 6034
rect 9932 6014 9944 6034
rect 9900 5976 9944 6014
rect 17390 6033 17434 6075
rect 17390 6013 17402 6033
rect 17422 6013 17434 6033
rect 17390 6006 17434 6013
rect 17389 5975 17434 6006
rect 17484 6033 17526 6075
rect 17484 6013 17498 6033
rect 17518 6013 17526 6033
rect 17484 5975 17526 6013
rect 17600 6033 17642 6075
rect 17600 6013 17608 6033
rect 17628 6013 17642 6033
rect 17600 5975 17642 6013
rect 17692 6033 17736 6075
rect 17692 6013 17704 6033
rect 17724 6013 17736 6033
rect 17692 5975 17736 6013
rect 17808 6033 17850 6075
rect 17808 6013 17816 6033
rect 17836 6013 17850 6033
rect 17808 5975 17850 6013
rect 17900 6033 17944 6075
rect 17900 6013 17912 6033
rect 17932 6013 17944 6033
rect 17900 5975 17944 6013
rect 18021 6033 18063 6075
rect 18021 6013 18029 6033
rect 18049 6013 18063 6033
rect 18021 5975 18063 6013
rect 18113 6033 18157 6075
rect 22560 6183 22572 6203
rect 22592 6183 22604 6203
rect 22560 6141 22604 6183
rect 22654 6203 22696 6241
rect 22654 6183 22668 6203
rect 22688 6183 22696 6203
rect 22654 6141 22696 6183
rect 22773 6203 22817 6241
rect 22773 6183 22785 6203
rect 22805 6183 22817 6203
rect 22773 6141 22817 6183
rect 22867 6203 22909 6241
rect 22867 6183 22881 6203
rect 22901 6183 22909 6203
rect 22867 6141 22909 6183
rect 22981 6203 23025 6241
rect 22981 6183 22993 6203
rect 23013 6183 23025 6203
rect 22981 6141 23025 6183
rect 23075 6203 23117 6241
rect 23075 6183 23089 6203
rect 23109 6183 23117 6203
rect 23075 6141 23117 6183
rect 23191 6203 23233 6241
rect 23191 6183 23199 6203
rect 23219 6183 23233 6203
rect 23191 6141 23233 6183
rect 23283 6210 23328 6241
rect 23283 6203 23327 6210
rect 23283 6183 23295 6203
rect 23315 6183 23327 6203
rect 23283 6141 23327 6183
rect 23608 6199 23652 6237
rect 23608 6179 23620 6199
rect 23640 6179 23652 6199
rect 18113 6013 18125 6033
rect 18145 6013 18157 6033
rect 18113 5975 18157 6013
rect 19885 6028 19929 6070
rect 19885 6008 19897 6028
rect 19917 6008 19929 6028
rect 19885 6001 19929 6008
rect 19884 5970 19929 6001
rect 19979 6028 20021 6070
rect 19979 6008 19993 6028
rect 20013 6008 20021 6028
rect 19979 5970 20021 6008
rect 20095 6028 20137 6070
rect 20095 6008 20103 6028
rect 20123 6008 20137 6028
rect 20095 5970 20137 6008
rect 20187 6028 20231 6070
rect 20187 6008 20199 6028
rect 20219 6008 20231 6028
rect 20187 5970 20231 6008
rect 20303 6028 20345 6070
rect 20303 6008 20311 6028
rect 20331 6008 20345 6028
rect 20303 5970 20345 6008
rect 20395 6028 20439 6070
rect 20395 6008 20407 6028
rect 20427 6008 20439 6028
rect 20395 5970 20439 6008
rect 20516 6028 20558 6070
rect 20516 6008 20524 6028
rect 20544 6008 20558 6028
rect 20516 5970 20558 6008
rect 20608 6028 20652 6070
rect 23608 6137 23652 6179
rect 23702 6199 23744 6237
rect 23702 6179 23716 6199
rect 23736 6179 23744 6199
rect 23702 6137 23744 6179
rect 23821 6199 23865 6237
rect 23821 6179 23833 6199
rect 23853 6179 23865 6199
rect 23821 6137 23865 6179
rect 23915 6199 23957 6237
rect 23915 6179 23929 6199
rect 23949 6179 23957 6199
rect 23915 6137 23957 6179
rect 24029 6199 24073 6237
rect 24029 6179 24041 6199
rect 24061 6179 24073 6199
rect 24029 6137 24073 6179
rect 24123 6199 24165 6237
rect 24123 6179 24137 6199
rect 24157 6179 24165 6199
rect 24123 6137 24165 6179
rect 24239 6199 24281 6237
rect 24239 6179 24247 6199
rect 24267 6179 24281 6199
rect 24239 6137 24281 6179
rect 24331 6206 24376 6237
rect 24331 6199 24375 6206
rect 24331 6179 24343 6199
rect 24363 6179 24375 6199
rect 24331 6137 24375 6179
rect 20608 6008 20620 6028
rect 20640 6008 20652 6028
rect 20608 5970 20652 6008
rect 33268 6197 33312 6235
rect 28355 6037 28399 6079
rect 28355 6017 28367 6037
rect 28387 6017 28399 6037
rect 28355 6010 28399 6017
rect 28354 5979 28399 6010
rect 28449 6037 28491 6079
rect 28449 6017 28463 6037
rect 28483 6017 28491 6037
rect 28449 5979 28491 6017
rect 28565 6037 28607 6079
rect 28565 6017 28573 6037
rect 28593 6017 28607 6037
rect 28565 5979 28607 6017
rect 28657 6037 28701 6079
rect 28657 6017 28669 6037
rect 28689 6017 28701 6037
rect 28657 5979 28701 6017
rect 28773 6037 28815 6079
rect 28773 6017 28781 6037
rect 28801 6017 28815 6037
rect 28773 5979 28815 6017
rect 28865 6037 28909 6079
rect 28865 6017 28877 6037
rect 28897 6017 28909 6037
rect 28865 5979 28909 6017
rect 28986 6037 29028 6079
rect 28986 6017 28994 6037
rect 29014 6017 29028 6037
rect 28986 5979 29028 6017
rect 29078 6037 29122 6079
rect 33268 6177 33280 6197
rect 33300 6177 33312 6197
rect 33268 6135 33312 6177
rect 33362 6197 33404 6235
rect 33362 6177 33376 6197
rect 33396 6177 33404 6197
rect 33362 6135 33404 6177
rect 33481 6197 33525 6235
rect 33481 6177 33493 6197
rect 33513 6177 33525 6197
rect 33481 6135 33525 6177
rect 33575 6197 33617 6235
rect 33575 6177 33589 6197
rect 33609 6177 33617 6197
rect 33575 6135 33617 6177
rect 33689 6197 33733 6235
rect 33689 6177 33701 6197
rect 33721 6177 33733 6197
rect 33689 6135 33733 6177
rect 33783 6197 33825 6235
rect 33783 6177 33797 6197
rect 33817 6177 33825 6197
rect 33783 6135 33825 6177
rect 33899 6197 33941 6235
rect 33899 6177 33907 6197
rect 33927 6177 33941 6197
rect 33899 6135 33941 6177
rect 33991 6204 34036 6235
rect 33991 6197 34035 6204
rect 33991 6177 34003 6197
rect 34023 6177 34035 6197
rect 33991 6135 34035 6177
rect 34316 6193 34360 6231
rect 34316 6173 34328 6193
rect 34348 6173 34360 6193
rect 29078 6017 29090 6037
rect 29110 6017 29122 6037
rect 29078 5979 29122 6017
rect 30850 6032 30894 6074
rect 30850 6012 30862 6032
rect 30882 6012 30894 6032
rect 30850 6005 30894 6012
rect 30849 5974 30894 6005
rect 30944 6032 30986 6074
rect 30944 6012 30958 6032
rect 30978 6012 30986 6032
rect 30944 5974 30986 6012
rect 31060 6032 31102 6074
rect 31060 6012 31068 6032
rect 31088 6012 31102 6032
rect 31060 5974 31102 6012
rect 31152 6032 31196 6074
rect 31152 6012 31164 6032
rect 31184 6012 31196 6032
rect 31152 5974 31196 6012
rect 31268 6032 31310 6074
rect 31268 6012 31276 6032
rect 31296 6012 31310 6032
rect 31268 5974 31310 6012
rect 31360 6032 31404 6074
rect 31360 6012 31372 6032
rect 31392 6012 31404 6032
rect 31360 5974 31404 6012
rect 31481 6032 31523 6074
rect 31481 6012 31489 6032
rect 31509 6012 31523 6032
rect 31481 5974 31523 6012
rect 31573 6032 31617 6074
rect 34316 6131 34360 6173
rect 34410 6193 34452 6231
rect 34410 6173 34424 6193
rect 34444 6173 34452 6193
rect 34410 6131 34452 6173
rect 34529 6193 34573 6231
rect 34529 6173 34541 6193
rect 34561 6173 34573 6193
rect 34529 6131 34573 6173
rect 34623 6193 34665 6231
rect 34623 6173 34637 6193
rect 34657 6173 34665 6193
rect 34623 6131 34665 6173
rect 34737 6193 34781 6231
rect 34737 6173 34749 6193
rect 34769 6173 34781 6193
rect 34737 6131 34781 6173
rect 34831 6193 34873 6231
rect 34831 6173 34845 6193
rect 34865 6173 34873 6193
rect 34831 6131 34873 6173
rect 34947 6193 34989 6231
rect 34947 6173 34955 6193
rect 34975 6173 34989 6193
rect 34947 6131 34989 6173
rect 35039 6200 35084 6231
rect 35039 6193 35083 6200
rect 35039 6173 35051 6193
rect 35071 6173 35083 6193
rect 35039 6131 35083 6173
rect 31573 6012 31585 6032
rect 31605 6012 31617 6032
rect 31573 5974 31617 6012
rect 39063 6031 39107 6073
rect 39063 6011 39075 6031
rect 39095 6011 39107 6031
rect 39063 6004 39107 6011
rect 39062 5973 39107 6004
rect 39157 6031 39199 6073
rect 39157 6011 39171 6031
rect 39191 6011 39199 6031
rect 39157 5973 39199 6011
rect 39273 6031 39315 6073
rect 39273 6011 39281 6031
rect 39301 6011 39315 6031
rect 39273 5973 39315 6011
rect 39365 6031 39409 6073
rect 39365 6011 39377 6031
rect 39397 6011 39409 6031
rect 39365 5973 39409 6011
rect 39481 6031 39523 6073
rect 39481 6011 39489 6031
rect 39509 6011 39523 6031
rect 39481 5973 39523 6011
rect 39573 6031 39617 6073
rect 39573 6011 39585 6031
rect 39605 6011 39617 6031
rect 39573 5973 39617 6011
rect 39694 6031 39736 6073
rect 39694 6011 39702 6031
rect 39722 6011 39736 6031
rect 39694 5973 39736 6011
rect 39786 6031 39830 6073
rect 39786 6011 39798 6031
rect 39818 6011 39830 6031
rect 39786 5973 39830 6011
rect 41558 6026 41602 6068
rect 41558 6006 41570 6026
rect 41590 6006 41602 6026
rect 41558 5999 41602 6006
rect 41557 5968 41602 5999
rect 41652 6026 41694 6068
rect 41652 6006 41666 6026
rect 41686 6006 41694 6026
rect 41652 5968 41694 6006
rect 41768 6026 41810 6068
rect 41768 6006 41776 6026
rect 41796 6006 41810 6026
rect 41768 5968 41810 6006
rect 41860 6026 41904 6068
rect 41860 6006 41872 6026
rect 41892 6006 41904 6026
rect 41860 5968 41904 6006
rect 41976 6026 42018 6068
rect 41976 6006 41984 6026
rect 42004 6006 42018 6026
rect 41976 5968 42018 6006
rect 42068 6026 42112 6068
rect 42068 6006 42080 6026
rect 42100 6006 42112 6026
rect 42068 5968 42112 6006
rect 42189 6026 42231 6068
rect 42189 6006 42197 6026
rect 42217 6006 42231 6026
rect 42189 5968 42231 6006
rect 42281 6026 42325 6068
rect 42281 6006 42293 6026
rect 42313 6006 42325 6026
rect 42281 5968 42325 6006
rect 887 5526 931 5564
rect 887 5506 899 5526
rect 919 5506 931 5526
rect 887 5464 931 5506
rect 981 5526 1023 5564
rect 981 5506 995 5526
rect 1015 5506 1023 5526
rect 981 5464 1023 5506
rect 1100 5526 1144 5564
rect 1100 5506 1112 5526
rect 1132 5506 1144 5526
rect 1100 5464 1144 5506
rect 1194 5526 1236 5564
rect 1194 5506 1208 5526
rect 1228 5506 1236 5526
rect 1194 5464 1236 5506
rect 1308 5526 1352 5564
rect 1308 5506 1320 5526
rect 1340 5506 1352 5526
rect 1308 5464 1352 5506
rect 1402 5526 1444 5564
rect 1402 5506 1416 5526
rect 1436 5506 1444 5526
rect 1402 5464 1444 5506
rect 1518 5526 1560 5564
rect 1518 5506 1526 5526
rect 1546 5506 1560 5526
rect 1518 5464 1560 5506
rect 1610 5533 1655 5564
rect 1610 5526 1654 5533
rect 1610 5506 1622 5526
rect 1642 5506 1654 5526
rect 1610 5464 1654 5506
rect 3425 5523 3469 5561
rect 3425 5503 3437 5523
rect 3457 5503 3469 5523
rect 3425 5461 3469 5503
rect 3519 5523 3561 5561
rect 3519 5503 3533 5523
rect 3553 5503 3561 5523
rect 3519 5461 3561 5503
rect 3638 5523 3682 5561
rect 3638 5503 3650 5523
rect 3670 5503 3682 5523
rect 3638 5461 3682 5503
rect 3732 5523 3774 5561
rect 3732 5503 3746 5523
rect 3766 5503 3774 5523
rect 3732 5461 3774 5503
rect 3846 5523 3890 5561
rect 3846 5503 3858 5523
rect 3878 5503 3890 5523
rect 3846 5461 3890 5503
rect 3940 5523 3982 5561
rect 3940 5503 3954 5523
rect 3974 5503 3982 5523
rect 3940 5461 3982 5503
rect 4056 5523 4098 5561
rect 4056 5503 4064 5523
rect 4084 5503 4098 5523
rect 4056 5461 4098 5503
rect 4148 5530 4193 5561
rect 4148 5523 4192 5530
rect 4148 5503 4160 5523
rect 4180 5503 4192 5523
rect 4148 5461 4192 5503
rect 11595 5520 11639 5558
rect 11595 5500 11607 5520
rect 11627 5500 11639 5520
rect 8129 5359 8173 5401
rect 8129 5339 8141 5359
rect 8161 5339 8173 5359
rect 8129 5332 8173 5339
rect 8128 5301 8173 5332
rect 8223 5359 8265 5401
rect 8223 5339 8237 5359
rect 8257 5339 8265 5359
rect 8223 5301 8265 5339
rect 8339 5359 8381 5401
rect 8339 5339 8347 5359
rect 8367 5339 8381 5359
rect 8339 5301 8381 5339
rect 8431 5359 8475 5401
rect 8431 5339 8443 5359
rect 8463 5339 8475 5359
rect 8431 5301 8475 5339
rect 8547 5359 8589 5401
rect 8547 5339 8555 5359
rect 8575 5339 8589 5359
rect 8547 5301 8589 5339
rect 8639 5359 8683 5401
rect 8639 5339 8651 5359
rect 8671 5339 8683 5359
rect 8639 5301 8683 5339
rect 8760 5359 8802 5401
rect 8760 5339 8768 5359
rect 8788 5339 8802 5359
rect 8760 5301 8802 5339
rect 8852 5359 8896 5401
rect 11595 5458 11639 5500
rect 11689 5520 11731 5558
rect 11689 5500 11703 5520
rect 11723 5500 11731 5520
rect 11689 5458 11731 5500
rect 11808 5520 11852 5558
rect 11808 5500 11820 5520
rect 11840 5500 11852 5520
rect 11808 5458 11852 5500
rect 11902 5520 11944 5558
rect 11902 5500 11916 5520
rect 11936 5500 11944 5520
rect 11902 5458 11944 5500
rect 12016 5520 12060 5558
rect 12016 5500 12028 5520
rect 12048 5500 12060 5520
rect 12016 5458 12060 5500
rect 12110 5520 12152 5558
rect 12110 5500 12124 5520
rect 12144 5500 12152 5520
rect 12110 5458 12152 5500
rect 12226 5520 12268 5558
rect 12226 5500 12234 5520
rect 12254 5500 12268 5520
rect 12226 5458 12268 5500
rect 12318 5527 12363 5558
rect 12318 5520 12362 5527
rect 12318 5500 12330 5520
rect 12350 5500 12362 5520
rect 12318 5458 12362 5500
rect 14133 5517 14177 5555
rect 14133 5497 14145 5517
rect 14165 5497 14177 5517
rect 8852 5339 8864 5359
rect 8884 5339 8896 5359
rect 8852 5301 8896 5339
rect 9177 5355 9221 5397
rect 9177 5335 9189 5355
rect 9209 5335 9221 5355
rect 9177 5328 9221 5335
rect 9176 5297 9221 5328
rect 9271 5355 9313 5397
rect 9271 5335 9285 5355
rect 9305 5335 9313 5355
rect 9271 5297 9313 5335
rect 9387 5355 9429 5397
rect 9387 5335 9395 5355
rect 9415 5335 9429 5355
rect 9387 5297 9429 5335
rect 9479 5355 9523 5397
rect 9479 5335 9491 5355
rect 9511 5335 9523 5355
rect 9479 5297 9523 5335
rect 9595 5355 9637 5397
rect 9595 5335 9603 5355
rect 9623 5335 9637 5355
rect 9595 5297 9637 5335
rect 9687 5355 9731 5397
rect 9687 5335 9699 5355
rect 9719 5335 9731 5355
rect 9687 5297 9731 5335
rect 9808 5355 9850 5397
rect 9808 5335 9816 5355
rect 9836 5335 9850 5355
rect 9808 5297 9850 5335
rect 9900 5355 9944 5397
rect 9900 5335 9912 5355
rect 9932 5335 9944 5355
rect 14133 5455 14177 5497
rect 14227 5517 14269 5555
rect 14227 5497 14241 5517
rect 14261 5497 14269 5517
rect 14227 5455 14269 5497
rect 14346 5517 14390 5555
rect 14346 5497 14358 5517
rect 14378 5497 14390 5517
rect 14346 5455 14390 5497
rect 14440 5517 14482 5555
rect 14440 5497 14454 5517
rect 14474 5497 14482 5517
rect 14440 5455 14482 5497
rect 14554 5517 14598 5555
rect 14554 5497 14566 5517
rect 14586 5497 14598 5517
rect 14554 5455 14598 5497
rect 14648 5517 14690 5555
rect 14648 5497 14662 5517
rect 14682 5497 14690 5517
rect 14648 5455 14690 5497
rect 14764 5517 14806 5555
rect 14764 5497 14772 5517
rect 14792 5497 14806 5517
rect 14764 5455 14806 5497
rect 14856 5524 14901 5555
rect 14856 5517 14900 5524
rect 14856 5497 14868 5517
rect 14888 5497 14900 5517
rect 14856 5455 14900 5497
rect 9900 5297 9944 5335
rect 22560 5524 22604 5562
rect 22560 5504 22572 5524
rect 22592 5504 22604 5524
rect 18837 5353 18881 5395
rect 18837 5333 18849 5353
rect 18869 5333 18881 5353
rect 18837 5326 18881 5333
rect 18836 5295 18881 5326
rect 18931 5353 18973 5395
rect 18931 5333 18945 5353
rect 18965 5333 18973 5353
rect 18931 5295 18973 5333
rect 19047 5353 19089 5395
rect 19047 5333 19055 5353
rect 19075 5333 19089 5353
rect 19047 5295 19089 5333
rect 19139 5353 19183 5395
rect 19139 5333 19151 5353
rect 19171 5333 19183 5353
rect 19139 5295 19183 5333
rect 19255 5353 19297 5395
rect 19255 5333 19263 5353
rect 19283 5333 19297 5353
rect 19255 5295 19297 5333
rect 19347 5353 19391 5395
rect 19347 5333 19359 5353
rect 19379 5333 19391 5353
rect 19347 5295 19391 5333
rect 19468 5353 19510 5395
rect 19468 5333 19476 5353
rect 19496 5333 19510 5353
rect 19468 5295 19510 5333
rect 19560 5353 19604 5395
rect 22560 5462 22604 5504
rect 22654 5524 22696 5562
rect 22654 5504 22668 5524
rect 22688 5504 22696 5524
rect 22654 5462 22696 5504
rect 22773 5524 22817 5562
rect 22773 5504 22785 5524
rect 22805 5504 22817 5524
rect 22773 5462 22817 5504
rect 22867 5524 22909 5562
rect 22867 5504 22881 5524
rect 22901 5504 22909 5524
rect 22867 5462 22909 5504
rect 22981 5524 23025 5562
rect 22981 5504 22993 5524
rect 23013 5504 23025 5524
rect 22981 5462 23025 5504
rect 23075 5524 23117 5562
rect 23075 5504 23089 5524
rect 23109 5504 23117 5524
rect 23075 5462 23117 5504
rect 23191 5524 23233 5562
rect 23191 5504 23199 5524
rect 23219 5504 23233 5524
rect 23191 5462 23233 5504
rect 23283 5531 23328 5562
rect 23283 5524 23327 5531
rect 23283 5504 23295 5524
rect 23315 5504 23327 5524
rect 23283 5462 23327 5504
rect 25098 5521 25142 5559
rect 25098 5501 25110 5521
rect 25130 5501 25142 5521
rect 19560 5333 19572 5353
rect 19592 5333 19604 5353
rect 19560 5295 19604 5333
rect 19885 5349 19929 5391
rect 19885 5329 19897 5349
rect 19917 5329 19929 5349
rect 19885 5322 19929 5329
rect 19884 5291 19929 5322
rect 19979 5349 20021 5391
rect 19979 5329 19993 5349
rect 20013 5329 20021 5349
rect 19979 5291 20021 5329
rect 20095 5349 20137 5391
rect 20095 5329 20103 5349
rect 20123 5329 20137 5349
rect 20095 5291 20137 5329
rect 20187 5349 20231 5391
rect 20187 5329 20199 5349
rect 20219 5329 20231 5349
rect 20187 5291 20231 5329
rect 20303 5349 20345 5391
rect 20303 5329 20311 5349
rect 20331 5329 20345 5349
rect 20303 5291 20345 5329
rect 20395 5349 20439 5391
rect 20395 5329 20407 5349
rect 20427 5329 20439 5349
rect 20395 5291 20439 5329
rect 20516 5349 20558 5391
rect 20516 5329 20524 5349
rect 20544 5329 20558 5349
rect 20516 5291 20558 5329
rect 20608 5349 20652 5391
rect 20608 5329 20620 5349
rect 20640 5329 20652 5349
rect 25098 5459 25142 5501
rect 25192 5521 25234 5559
rect 25192 5501 25206 5521
rect 25226 5501 25234 5521
rect 25192 5459 25234 5501
rect 25311 5521 25355 5559
rect 25311 5501 25323 5521
rect 25343 5501 25355 5521
rect 25311 5459 25355 5501
rect 25405 5521 25447 5559
rect 25405 5501 25419 5521
rect 25439 5501 25447 5521
rect 25405 5459 25447 5501
rect 25519 5521 25563 5559
rect 25519 5501 25531 5521
rect 25551 5501 25563 5521
rect 25519 5459 25563 5501
rect 25613 5521 25655 5559
rect 25613 5501 25627 5521
rect 25647 5501 25655 5521
rect 25613 5459 25655 5501
rect 25729 5521 25771 5559
rect 25729 5501 25737 5521
rect 25757 5501 25771 5521
rect 25729 5459 25771 5501
rect 25821 5528 25866 5559
rect 25821 5521 25865 5528
rect 25821 5501 25833 5521
rect 25853 5501 25865 5521
rect 25821 5459 25865 5501
rect 33268 5518 33312 5556
rect 33268 5498 33280 5518
rect 33300 5498 33312 5518
rect 20608 5291 20652 5329
rect 29802 5357 29846 5399
rect 29802 5337 29814 5357
rect 29834 5337 29846 5357
rect 29802 5330 29846 5337
rect 29801 5299 29846 5330
rect 29896 5357 29938 5399
rect 29896 5337 29910 5357
rect 29930 5337 29938 5357
rect 29896 5299 29938 5337
rect 30012 5357 30054 5399
rect 30012 5337 30020 5357
rect 30040 5337 30054 5357
rect 30012 5299 30054 5337
rect 30104 5357 30148 5399
rect 30104 5337 30116 5357
rect 30136 5337 30148 5357
rect 30104 5299 30148 5337
rect 30220 5357 30262 5399
rect 30220 5337 30228 5357
rect 30248 5337 30262 5357
rect 30220 5299 30262 5337
rect 30312 5357 30356 5399
rect 30312 5337 30324 5357
rect 30344 5337 30356 5357
rect 30312 5299 30356 5337
rect 30433 5357 30475 5399
rect 30433 5337 30441 5357
rect 30461 5337 30475 5357
rect 30433 5299 30475 5337
rect 30525 5357 30569 5399
rect 33268 5456 33312 5498
rect 33362 5518 33404 5556
rect 33362 5498 33376 5518
rect 33396 5498 33404 5518
rect 33362 5456 33404 5498
rect 33481 5518 33525 5556
rect 33481 5498 33493 5518
rect 33513 5498 33525 5518
rect 33481 5456 33525 5498
rect 33575 5518 33617 5556
rect 33575 5498 33589 5518
rect 33609 5498 33617 5518
rect 33575 5456 33617 5498
rect 33689 5518 33733 5556
rect 33689 5498 33701 5518
rect 33721 5498 33733 5518
rect 33689 5456 33733 5498
rect 33783 5518 33825 5556
rect 33783 5498 33797 5518
rect 33817 5498 33825 5518
rect 33783 5456 33825 5498
rect 33899 5518 33941 5556
rect 33899 5498 33907 5518
rect 33927 5498 33941 5518
rect 33899 5456 33941 5498
rect 33991 5525 34036 5556
rect 33991 5518 34035 5525
rect 33991 5498 34003 5518
rect 34023 5498 34035 5518
rect 33991 5456 34035 5498
rect 35806 5515 35850 5553
rect 35806 5495 35818 5515
rect 35838 5495 35850 5515
rect 30525 5337 30537 5357
rect 30557 5337 30569 5357
rect 30525 5299 30569 5337
rect 30850 5353 30894 5395
rect 30850 5333 30862 5353
rect 30882 5333 30894 5353
rect 30850 5326 30894 5333
rect 30849 5295 30894 5326
rect 30944 5353 30986 5395
rect 30944 5333 30958 5353
rect 30978 5333 30986 5353
rect 30944 5295 30986 5333
rect 31060 5353 31102 5395
rect 31060 5333 31068 5353
rect 31088 5333 31102 5353
rect 31060 5295 31102 5333
rect 31152 5353 31196 5395
rect 31152 5333 31164 5353
rect 31184 5333 31196 5353
rect 31152 5295 31196 5333
rect 31268 5353 31310 5395
rect 31268 5333 31276 5353
rect 31296 5333 31310 5353
rect 31268 5295 31310 5333
rect 31360 5353 31404 5395
rect 31360 5333 31372 5353
rect 31392 5333 31404 5353
rect 31360 5295 31404 5333
rect 31481 5353 31523 5395
rect 31481 5333 31489 5353
rect 31509 5333 31523 5353
rect 31481 5295 31523 5333
rect 31573 5353 31617 5395
rect 31573 5333 31585 5353
rect 31605 5333 31617 5353
rect 35806 5453 35850 5495
rect 35900 5515 35942 5553
rect 35900 5495 35914 5515
rect 35934 5495 35942 5515
rect 35900 5453 35942 5495
rect 36019 5515 36063 5553
rect 36019 5495 36031 5515
rect 36051 5495 36063 5515
rect 36019 5453 36063 5495
rect 36113 5515 36155 5553
rect 36113 5495 36127 5515
rect 36147 5495 36155 5515
rect 36113 5453 36155 5495
rect 36227 5515 36271 5553
rect 36227 5495 36239 5515
rect 36259 5495 36271 5515
rect 36227 5453 36271 5495
rect 36321 5515 36363 5553
rect 36321 5495 36335 5515
rect 36355 5495 36363 5515
rect 36321 5453 36363 5495
rect 36437 5515 36479 5553
rect 36437 5495 36445 5515
rect 36465 5495 36479 5515
rect 36437 5453 36479 5495
rect 36529 5522 36574 5553
rect 36529 5515 36573 5522
rect 36529 5495 36541 5515
rect 36561 5495 36573 5515
rect 36529 5453 36573 5495
rect 31573 5295 31617 5333
rect 40510 5351 40554 5393
rect 40510 5331 40522 5351
rect 40542 5331 40554 5351
rect 40510 5324 40554 5331
rect 40509 5293 40554 5324
rect 40604 5351 40646 5393
rect 40604 5331 40618 5351
rect 40638 5331 40646 5351
rect 40604 5293 40646 5331
rect 40720 5351 40762 5393
rect 40720 5331 40728 5351
rect 40748 5331 40762 5351
rect 40720 5293 40762 5331
rect 40812 5351 40856 5393
rect 40812 5331 40824 5351
rect 40844 5331 40856 5351
rect 40812 5293 40856 5331
rect 40928 5351 40970 5393
rect 40928 5331 40936 5351
rect 40956 5331 40970 5351
rect 40928 5293 40970 5331
rect 41020 5351 41064 5393
rect 41020 5331 41032 5351
rect 41052 5331 41064 5351
rect 41020 5293 41064 5331
rect 41141 5351 41183 5393
rect 41141 5331 41149 5351
rect 41169 5331 41183 5351
rect 41141 5293 41183 5331
rect 41233 5351 41277 5393
rect 41233 5331 41245 5351
rect 41265 5331 41277 5351
rect 41233 5293 41277 5331
rect 41558 5347 41602 5389
rect 41558 5327 41570 5347
rect 41590 5327 41602 5347
rect 41558 5320 41602 5327
rect 41557 5289 41602 5320
rect 41652 5347 41694 5389
rect 41652 5327 41666 5347
rect 41686 5327 41694 5347
rect 41652 5289 41694 5327
rect 41768 5347 41810 5389
rect 41768 5327 41776 5347
rect 41796 5327 41810 5347
rect 41768 5289 41810 5327
rect 41860 5347 41904 5389
rect 41860 5327 41872 5347
rect 41892 5327 41904 5347
rect 41860 5289 41904 5327
rect 41976 5347 42018 5389
rect 41976 5327 41984 5347
rect 42004 5327 42018 5347
rect 41976 5289 42018 5327
rect 42068 5347 42112 5389
rect 42068 5327 42080 5347
rect 42100 5327 42112 5347
rect 42068 5289 42112 5327
rect 42189 5347 42231 5389
rect 42189 5327 42197 5347
rect 42217 5327 42231 5347
rect 42189 5289 42231 5327
rect 42281 5347 42325 5389
rect 42281 5327 42293 5347
rect 42313 5327 42325 5347
rect 42281 5289 42325 5327
rect 888 4685 932 4723
rect 888 4665 900 4685
rect 920 4665 932 4685
rect 888 4623 932 4665
rect 982 4685 1024 4723
rect 982 4665 996 4685
rect 1016 4665 1024 4685
rect 982 4623 1024 4665
rect 1101 4685 1145 4723
rect 1101 4665 1113 4685
rect 1133 4665 1145 4685
rect 1101 4623 1145 4665
rect 1195 4685 1237 4723
rect 1195 4665 1209 4685
rect 1229 4665 1237 4685
rect 1195 4623 1237 4665
rect 1309 4685 1353 4723
rect 1309 4665 1321 4685
rect 1341 4665 1353 4685
rect 1309 4623 1353 4665
rect 1403 4685 1445 4723
rect 1403 4665 1417 4685
rect 1437 4665 1445 4685
rect 1403 4623 1445 4665
rect 1519 4685 1561 4723
rect 1519 4665 1527 4685
rect 1547 4665 1561 4685
rect 1519 4623 1561 4665
rect 1611 4692 1656 4723
rect 1611 4685 1655 4692
rect 1611 4665 1623 4685
rect 1643 4665 1655 4685
rect 1611 4623 1655 4665
rect 1936 4681 1980 4719
rect 1936 4661 1948 4681
rect 1968 4661 1980 4681
rect 1936 4619 1980 4661
rect 2030 4681 2072 4719
rect 2030 4661 2044 4681
rect 2064 4661 2072 4681
rect 2030 4619 2072 4661
rect 2149 4681 2193 4719
rect 2149 4661 2161 4681
rect 2181 4661 2193 4681
rect 2149 4619 2193 4661
rect 2243 4681 2285 4719
rect 2243 4661 2257 4681
rect 2277 4661 2285 4681
rect 2243 4619 2285 4661
rect 2357 4681 2401 4719
rect 2357 4661 2369 4681
rect 2389 4661 2401 4681
rect 2357 4619 2401 4661
rect 2451 4681 2493 4719
rect 2451 4661 2465 4681
rect 2485 4661 2493 4681
rect 2451 4619 2493 4661
rect 2567 4681 2609 4719
rect 2567 4661 2575 4681
rect 2595 4661 2609 4681
rect 2567 4619 2609 4661
rect 2659 4688 2704 4719
rect 2659 4681 2703 4688
rect 2659 4661 2671 4681
rect 2691 4661 2703 4681
rect 2659 4619 2703 4661
rect 4838 4687 4882 4725
rect 4838 4667 4850 4687
rect 4870 4667 4882 4687
rect 4838 4625 4882 4667
rect 4932 4687 4974 4725
rect 4932 4667 4946 4687
rect 4966 4667 4974 4687
rect 4932 4625 4974 4667
rect 5051 4687 5095 4725
rect 5051 4667 5063 4687
rect 5083 4667 5095 4687
rect 5051 4625 5095 4667
rect 5145 4687 5187 4725
rect 5145 4667 5159 4687
rect 5179 4667 5187 4687
rect 5145 4625 5187 4667
rect 5259 4687 5303 4725
rect 5259 4667 5271 4687
rect 5291 4667 5303 4687
rect 5259 4625 5303 4667
rect 5353 4687 5395 4725
rect 5353 4667 5367 4687
rect 5387 4667 5395 4687
rect 5353 4625 5395 4667
rect 5469 4687 5511 4725
rect 5469 4667 5477 4687
rect 5497 4667 5511 4687
rect 5469 4625 5511 4667
rect 5561 4694 5606 4725
rect 5561 4687 5605 4694
rect 5561 4667 5573 4687
rect 5593 4667 5605 4687
rect 5561 4625 5605 4667
rect 11596 4679 11640 4717
rect 6640 4517 6684 4559
rect 6640 4497 6652 4517
rect 6672 4497 6684 4517
rect 6640 4490 6684 4497
rect 6639 4459 6684 4490
rect 6734 4517 6776 4559
rect 6734 4497 6748 4517
rect 6768 4497 6776 4517
rect 6734 4459 6776 4497
rect 6850 4517 6892 4559
rect 6850 4497 6858 4517
rect 6878 4497 6892 4517
rect 6850 4459 6892 4497
rect 6942 4517 6986 4559
rect 6942 4497 6954 4517
rect 6974 4497 6986 4517
rect 6942 4459 6986 4497
rect 7058 4517 7100 4559
rect 7058 4497 7066 4517
rect 7086 4497 7100 4517
rect 7058 4459 7100 4497
rect 7150 4517 7194 4559
rect 7150 4497 7162 4517
rect 7182 4497 7194 4517
rect 7150 4459 7194 4497
rect 7271 4517 7313 4559
rect 7271 4497 7279 4517
rect 7299 4497 7313 4517
rect 7271 4459 7313 4497
rect 7363 4517 7407 4559
rect 11596 4659 11608 4679
rect 11628 4659 11640 4679
rect 11596 4617 11640 4659
rect 11690 4679 11732 4717
rect 11690 4659 11704 4679
rect 11724 4659 11732 4679
rect 11690 4617 11732 4659
rect 11809 4679 11853 4717
rect 11809 4659 11821 4679
rect 11841 4659 11853 4679
rect 11809 4617 11853 4659
rect 11903 4679 11945 4717
rect 11903 4659 11917 4679
rect 11937 4659 11945 4679
rect 11903 4617 11945 4659
rect 12017 4679 12061 4717
rect 12017 4659 12029 4679
rect 12049 4659 12061 4679
rect 12017 4617 12061 4659
rect 12111 4679 12153 4717
rect 12111 4659 12125 4679
rect 12145 4659 12153 4679
rect 12111 4617 12153 4659
rect 12227 4679 12269 4717
rect 12227 4659 12235 4679
rect 12255 4659 12269 4679
rect 12227 4617 12269 4659
rect 12319 4686 12364 4717
rect 12319 4679 12363 4686
rect 12319 4659 12331 4679
rect 12351 4659 12363 4679
rect 12319 4617 12363 4659
rect 12644 4675 12688 4713
rect 12644 4655 12656 4675
rect 12676 4655 12688 4675
rect 7363 4497 7375 4517
rect 7395 4497 7407 4517
rect 7363 4459 7407 4497
rect 9178 4514 9222 4556
rect 9178 4494 9190 4514
rect 9210 4494 9222 4514
rect 9178 4487 9222 4494
rect 9177 4456 9222 4487
rect 9272 4514 9314 4556
rect 9272 4494 9286 4514
rect 9306 4494 9314 4514
rect 9272 4456 9314 4494
rect 9388 4514 9430 4556
rect 9388 4494 9396 4514
rect 9416 4494 9430 4514
rect 9388 4456 9430 4494
rect 9480 4514 9524 4556
rect 9480 4494 9492 4514
rect 9512 4494 9524 4514
rect 9480 4456 9524 4494
rect 9596 4514 9638 4556
rect 9596 4494 9604 4514
rect 9624 4494 9638 4514
rect 9596 4456 9638 4494
rect 9688 4514 9732 4556
rect 9688 4494 9700 4514
rect 9720 4494 9732 4514
rect 9688 4456 9732 4494
rect 9809 4514 9851 4556
rect 9809 4494 9817 4514
rect 9837 4494 9851 4514
rect 9809 4456 9851 4494
rect 9901 4514 9945 4556
rect 12644 4613 12688 4655
rect 12738 4675 12780 4713
rect 12738 4655 12752 4675
rect 12772 4655 12780 4675
rect 12738 4613 12780 4655
rect 12857 4675 12901 4713
rect 12857 4655 12869 4675
rect 12889 4655 12901 4675
rect 12857 4613 12901 4655
rect 12951 4675 12993 4713
rect 12951 4655 12965 4675
rect 12985 4655 12993 4675
rect 12951 4613 12993 4655
rect 13065 4675 13109 4713
rect 13065 4655 13077 4675
rect 13097 4655 13109 4675
rect 13065 4613 13109 4655
rect 13159 4675 13201 4713
rect 13159 4655 13173 4675
rect 13193 4655 13201 4675
rect 13159 4613 13201 4655
rect 13275 4675 13317 4713
rect 13275 4655 13283 4675
rect 13303 4655 13317 4675
rect 13275 4613 13317 4655
rect 13367 4682 13412 4713
rect 13367 4675 13411 4682
rect 13367 4655 13379 4675
rect 13399 4655 13411 4675
rect 13367 4613 13411 4655
rect 15546 4681 15590 4719
rect 15546 4661 15558 4681
rect 15578 4661 15590 4681
rect 15546 4619 15590 4661
rect 15640 4681 15682 4719
rect 15640 4661 15654 4681
rect 15674 4661 15682 4681
rect 15640 4619 15682 4661
rect 15759 4681 15803 4719
rect 15759 4661 15771 4681
rect 15791 4661 15803 4681
rect 15759 4619 15803 4661
rect 15853 4681 15895 4719
rect 15853 4661 15867 4681
rect 15887 4661 15895 4681
rect 15853 4619 15895 4661
rect 15967 4681 16011 4719
rect 15967 4661 15979 4681
rect 15999 4661 16011 4681
rect 15967 4619 16011 4661
rect 16061 4681 16103 4719
rect 16061 4661 16075 4681
rect 16095 4661 16103 4681
rect 16061 4619 16103 4661
rect 16177 4681 16219 4719
rect 16177 4661 16185 4681
rect 16205 4661 16219 4681
rect 16177 4619 16219 4661
rect 16269 4688 16314 4719
rect 16269 4681 16313 4688
rect 16269 4661 16281 4681
rect 16301 4661 16313 4681
rect 16269 4619 16313 4661
rect 22561 4683 22605 4721
rect 9901 4494 9913 4514
rect 9933 4494 9945 4514
rect 9901 4456 9945 4494
rect 17348 4511 17392 4553
rect 17348 4491 17360 4511
rect 17380 4491 17392 4511
rect 17348 4484 17392 4491
rect 17347 4453 17392 4484
rect 17442 4511 17484 4553
rect 17442 4491 17456 4511
rect 17476 4491 17484 4511
rect 17442 4453 17484 4491
rect 17558 4511 17600 4553
rect 17558 4491 17566 4511
rect 17586 4491 17600 4511
rect 17558 4453 17600 4491
rect 17650 4511 17694 4553
rect 17650 4491 17662 4511
rect 17682 4491 17694 4511
rect 17650 4453 17694 4491
rect 17766 4511 17808 4553
rect 17766 4491 17774 4511
rect 17794 4491 17808 4511
rect 17766 4453 17808 4491
rect 17858 4511 17902 4553
rect 17858 4491 17870 4511
rect 17890 4491 17902 4511
rect 17858 4453 17902 4491
rect 17979 4511 18021 4553
rect 17979 4491 17987 4511
rect 18007 4491 18021 4511
rect 17979 4453 18021 4491
rect 18071 4511 18115 4553
rect 22561 4663 22573 4683
rect 22593 4663 22605 4683
rect 22561 4621 22605 4663
rect 22655 4683 22697 4721
rect 22655 4663 22669 4683
rect 22689 4663 22697 4683
rect 22655 4621 22697 4663
rect 22774 4683 22818 4721
rect 22774 4663 22786 4683
rect 22806 4663 22818 4683
rect 22774 4621 22818 4663
rect 22868 4683 22910 4721
rect 22868 4663 22882 4683
rect 22902 4663 22910 4683
rect 22868 4621 22910 4663
rect 22982 4683 23026 4721
rect 22982 4663 22994 4683
rect 23014 4663 23026 4683
rect 22982 4621 23026 4663
rect 23076 4683 23118 4721
rect 23076 4663 23090 4683
rect 23110 4663 23118 4683
rect 23076 4621 23118 4663
rect 23192 4683 23234 4721
rect 23192 4663 23200 4683
rect 23220 4663 23234 4683
rect 23192 4621 23234 4663
rect 23284 4690 23329 4721
rect 23284 4683 23328 4690
rect 23284 4663 23296 4683
rect 23316 4663 23328 4683
rect 23284 4621 23328 4663
rect 23609 4679 23653 4717
rect 23609 4659 23621 4679
rect 23641 4659 23653 4679
rect 18071 4491 18083 4511
rect 18103 4491 18115 4511
rect 18071 4453 18115 4491
rect 19886 4508 19930 4550
rect 19886 4488 19898 4508
rect 19918 4488 19930 4508
rect 19886 4481 19930 4488
rect 19885 4450 19930 4481
rect 19980 4508 20022 4550
rect 19980 4488 19994 4508
rect 20014 4488 20022 4508
rect 19980 4450 20022 4488
rect 20096 4508 20138 4550
rect 20096 4488 20104 4508
rect 20124 4488 20138 4508
rect 20096 4450 20138 4488
rect 20188 4508 20232 4550
rect 20188 4488 20200 4508
rect 20220 4488 20232 4508
rect 20188 4450 20232 4488
rect 20304 4508 20346 4550
rect 20304 4488 20312 4508
rect 20332 4488 20346 4508
rect 20304 4450 20346 4488
rect 20396 4508 20440 4550
rect 20396 4488 20408 4508
rect 20428 4488 20440 4508
rect 20396 4450 20440 4488
rect 20517 4508 20559 4550
rect 20517 4488 20525 4508
rect 20545 4488 20559 4508
rect 20517 4450 20559 4488
rect 20609 4508 20653 4550
rect 23609 4617 23653 4659
rect 23703 4679 23745 4717
rect 23703 4659 23717 4679
rect 23737 4659 23745 4679
rect 23703 4617 23745 4659
rect 23822 4679 23866 4717
rect 23822 4659 23834 4679
rect 23854 4659 23866 4679
rect 23822 4617 23866 4659
rect 23916 4679 23958 4717
rect 23916 4659 23930 4679
rect 23950 4659 23958 4679
rect 23916 4617 23958 4659
rect 24030 4679 24074 4717
rect 24030 4659 24042 4679
rect 24062 4659 24074 4679
rect 24030 4617 24074 4659
rect 24124 4679 24166 4717
rect 24124 4659 24138 4679
rect 24158 4659 24166 4679
rect 24124 4617 24166 4659
rect 24240 4679 24282 4717
rect 24240 4659 24248 4679
rect 24268 4659 24282 4679
rect 24240 4617 24282 4659
rect 24332 4686 24377 4717
rect 24332 4679 24376 4686
rect 24332 4659 24344 4679
rect 24364 4659 24376 4679
rect 24332 4617 24376 4659
rect 26511 4685 26555 4723
rect 26511 4665 26523 4685
rect 26543 4665 26555 4685
rect 26511 4623 26555 4665
rect 26605 4685 26647 4723
rect 26605 4665 26619 4685
rect 26639 4665 26647 4685
rect 26605 4623 26647 4665
rect 26724 4685 26768 4723
rect 26724 4665 26736 4685
rect 26756 4665 26768 4685
rect 26724 4623 26768 4665
rect 26818 4685 26860 4723
rect 26818 4665 26832 4685
rect 26852 4665 26860 4685
rect 26818 4623 26860 4665
rect 26932 4685 26976 4723
rect 26932 4665 26944 4685
rect 26964 4665 26976 4685
rect 26932 4623 26976 4665
rect 27026 4685 27068 4723
rect 27026 4665 27040 4685
rect 27060 4665 27068 4685
rect 27026 4623 27068 4665
rect 27142 4685 27184 4723
rect 27142 4665 27150 4685
rect 27170 4665 27184 4685
rect 27142 4623 27184 4665
rect 27234 4692 27279 4723
rect 27234 4685 27278 4692
rect 27234 4665 27246 4685
rect 27266 4665 27278 4685
rect 27234 4623 27278 4665
rect 20609 4488 20621 4508
rect 20641 4488 20653 4508
rect 20609 4450 20653 4488
rect 33269 4677 33313 4715
rect 28313 4515 28357 4557
rect 28313 4495 28325 4515
rect 28345 4495 28357 4515
rect 28313 4488 28357 4495
rect 28312 4457 28357 4488
rect 28407 4515 28449 4557
rect 28407 4495 28421 4515
rect 28441 4495 28449 4515
rect 28407 4457 28449 4495
rect 28523 4515 28565 4557
rect 28523 4495 28531 4515
rect 28551 4495 28565 4515
rect 28523 4457 28565 4495
rect 28615 4515 28659 4557
rect 28615 4495 28627 4515
rect 28647 4495 28659 4515
rect 28615 4457 28659 4495
rect 28731 4515 28773 4557
rect 28731 4495 28739 4515
rect 28759 4495 28773 4515
rect 28731 4457 28773 4495
rect 28823 4515 28867 4557
rect 28823 4495 28835 4515
rect 28855 4495 28867 4515
rect 28823 4457 28867 4495
rect 28944 4515 28986 4557
rect 28944 4495 28952 4515
rect 28972 4495 28986 4515
rect 28944 4457 28986 4495
rect 29036 4515 29080 4557
rect 33269 4657 33281 4677
rect 33301 4657 33313 4677
rect 33269 4615 33313 4657
rect 33363 4677 33405 4715
rect 33363 4657 33377 4677
rect 33397 4657 33405 4677
rect 33363 4615 33405 4657
rect 33482 4677 33526 4715
rect 33482 4657 33494 4677
rect 33514 4657 33526 4677
rect 33482 4615 33526 4657
rect 33576 4677 33618 4715
rect 33576 4657 33590 4677
rect 33610 4657 33618 4677
rect 33576 4615 33618 4657
rect 33690 4677 33734 4715
rect 33690 4657 33702 4677
rect 33722 4657 33734 4677
rect 33690 4615 33734 4657
rect 33784 4677 33826 4715
rect 33784 4657 33798 4677
rect 33818 4657 33826 4677
rect 33784 4615 33826 4657
rect 33900 4677 33942 4715
rect 33900 4657 33908 4677
rect 33928 4657 33942 4677
rect 33900 4615 33942 4657
rect 33992 4684 34037 4715
rect 33992 4677 34036 4684
rect 33992 4657 34004 4677
rect 34024 4657 34036 4677
rect 33992 4615 34036 4657
rect 34317 4673 34361 4711
rect 34317 4653 34329 4673
rect 34349 4653 34361 4673
rect 29036 4495 29048 4515
rect 29068 4495 29080 4515
rect 29036 4457 29080 4495
rect 30851 4512 30895 4554
rect 30851 4492 30863 4512
rect 30883 4492 30895 4512
rect 30851 4485 30895 4492
rect 30850 4454 30895 4485
rect 30945 4512 30987 4554
rect 30945 4492 30959 4512
rect 30979 4492 30987 4512
rect 30945 4454 30987 4492
rect 31061 4512 31103 4554
rect 31061 4492 31069 4512
rect 31089 4492 31103 4512
rect 31061 4454 31103 4492
rect 31153 4512 31197 4554
rect 31153 4492 31165 4512
rect 31185 4492 31197 4512
rect 31153 4454 31197 4492
rect 31269 4512 31311 4554
rect 31269 4492 31277 4512
rect 31297 4492 31311 4512
rect 31269 4454 31311 4492
rect 31361 4512 31405 4554
rect 31361 4492 31373 4512
rect 31393 4492 31405 4512
rect 31361 4454 31405 4492
rect 31482 4512 31524 4554
rect 31482 4492 31490 4512
rect 31510 4492 31524 4512
rect 31482 4454 31524 4492
rect 31574 4512 31618 4554
rect 34317 4611 34361 4653
rect 34411 4673 34453 4711
rect 34411 4653 34425 4673
rect 34445 4653 34453 4673
rect 34411 4611 34453 4653
rect 34530 4673 34574 4711
rect 34530 4653 34542 4673
rect 34562 4653 34574 4673
rect 34530 4611 34574 4653
rect 34624 4673 34666 4711
rect 34624 4653 34638 4673
rect 34658 4653 34666 4673
rect 34624 4611 34666 4653
rect 34738 4673 34782 4711
rect 34738 4653 34750 4673
rect 34770 4653 34782 4673
rect 34738 4611 34782 4653
rect 34832 4673 34874 4711
rect 34832 4653 34846 4673
rect 34866 4653 34874 4673
rect 34832 4611 34874 4653
rect 34948 4673 34990 4711
rect 34948 4653 34956 4673
rect 34976 4653 34990 4673
rect 34948 4611 34990 4653
rect 35040 4680 35085 4711
rect 35040 4673 35084 4680
rect 35040 4653 35052 4673
rect 35072 4653 35084 4673
rect 35040 4611 35084 4653
rect 37219 4679 37263 4717
rect 37219 4659 37231 4679
rect 37251 4659 37263 4679
rect 37219 4617 37263 4659
rect 37313 4679 37355 4717
rect 37313 4659 37327 4679
rect 37347 4659 37355 4679
rect 37313 4617 37355 4659
rect 37432 4679 37476 4717
rect 37432 4659 37444 4679
rect 37464 4659 37476 4679
rect 37432 4617 37476 4659
rect 37526 4679 37568 4717
rect 37526 4659 37540 4679
rect 37560 4659 37568 4679
rect 37526 4617 37568 4659
rect 37640 4679 37684 4717
rect 37640 4659 37652 4679
rect 37672 4659 37684 4679
rect 37640 4617 37684 4659
rect 37734 4679 37776 4717
rect 37734 4659 37748 4679
rect 37768 4659 37776 4679
rect 37734 4617 37776 4659
rect 37850 4679 37892 4717
rect 37850 4659 37858 4679
rect 37878 4659 37892 4679
rect 37850 4617 37892 4659
rect 37942 4686 37987 4717
rect 37942 4679 37986 4686
rect 37942 4659 37954 4679
rect 37974 4659 37986 4679
rect 37942 4617 37986 4659
rect 31574 4492 31586 4512
rect 31606 4492 31618 4512
rect 31574 4454 31618 4492
rect 39021 4509 39065 4551
rect 39021 4489 39033 4509
rect 39053 4489 39065 4509
rect 39021 4482 39065 4489
rect 39020 4451 39065 4482
rect 39115 4509 39157 4551
rect 39115 4489 39129 4509
rect 39149 4489 39157 4509
rect 39115 4451 39157 4489
rect 39231 4509 39273 4551
rect 39231 4489 39239 4509
rect 39259 4489 39273 4509
rect 39231 4451 39273 4489
rect 39323 4509 39367 4551
rect 39323 4489 39335 4509
rect 39355 4489 39367 4509
rect 39323 4451 39367 4489
rect 39439 4509 39481 4551
rect 39439 4489 39447 4509
rect 39467 4489 39481 4509
rect 39439 4451 39481 4489
rect 39531 4509 39575 4551
rect 39531 4489 39543 4509
rect 39563 4489 39575 4509
rect 39531 4451 39575 4489
rect 39652 4509 39694 4551
rect 39652 4489 39660 4509
rect 39680 4489 39694 4509
rect 39652 4451 39694 4489
rect 39744 4509 39788 4551
rect 39744 4489 39756 4509
rect 39776 4489 39788 4509
rect 39744 4451 39788 4489
rect 41559 4506 41603 4548
rect 41559 4486 41571 4506
rect 41591 4486 41603 4506
rect 41559 4479 41603 4486
rect 41558 4448 41603 4479
rect 41653 4506 41695 4548
rect 41653 4486 41667 4506
rect 41687 4486 41695 4506
rect 41653 4448 41695 4486
rect 41769 4506 41811 4548
rect 41769 4486 41777 4506
rect 41797 4486 41811 4506
rect 41769 4448 41811 4486
rect 41861 4506 41905 4548
rect 41861 4486 41873 4506
rect 41893 4486 41905 4506
rect 41861 4448 41905 4486
rect 41977 4506 42019 4548
rect 41977 4486 41985 4506
rect 42005 4486 42019 4506
rect 41977 4448 42019 4486
rect 42069 4506 42113 4548
rect 42069 4486 42081 4506
rect 42101 4486 42113 4506
rect 42069 4448 42113 4486
rect 42190 4506 42232 4548
rect 42190 4486 42198 4506
rect 42218 4486 42232 4506
rect 42190 4448 42232 4486
rect 42282 4506 42326 4548
rect 42282 4486 42294 4506
rect 42314 4486 42326 4506
rect 42282 4448 42326 4486
rect 888 4006 932 4044
rect 888 3986 900 4006
rect 920 3986 932 4006
rect 888 3944 932 3986
rect 982 4006 1024 4044
rect 982 3986 996 4006
rect 1016 3986 1024 4006
rect 982 3944 1024 3986
rect 1101 4006 1145 4044
rect 1101 3986 1113 4006
rect 1133 3986 1145 4006
rect 1101 3944 1145 3986
rect 1195 4006 1237 4044
rect 1195 3986 1209 4006
rect 1229 3986 1237 4006
rect 1195 3944 1237 3986
rect 1309 4006 1353 4044
rect 1309 3986 1321 4006
rect 1341 3986 1353 4006
rect 1309 3944 1353 3986
rect 1403 4006 1445 4044
rect 1403 3986 1417 4006
rect 1437 3986 1445 4006
rect 1403 3944 1445 3986
rect 1519 4006 1561 4044
rect 1519 3986 1527 4006
rect 1547 3986 1561 4006
rect 1519 3944 1561 3986
rect 1611 4013 1656 4044
rect 1611 4006 1655 4013
rect 1611 3986 1623 4006
rect 1643 3986 1655 4006
rect 1611 3944 1655 3986
rect 3383 4001 3427 4039
rect 3383 3981 3395 4001
rect 3415 3981 3427 4001
rect 3383 3939 3427 3981
rect 3477 4001 3519 4039
rect 3477 3981 3491 4001
rect 3511 3981 3519 4001
rect 3477 3939 3519 3981
rect 3596 4001 3640 4039
rect 3596 3981 3608 4001
rect 3628 3981 3640 4001
rect 3596 3939 3640 3981
rect 3690 4001 3732 4039
rect 3690 3981 3704 4001
rect 3724 3981 3732 4001
rect 3690 3939 3732 3981
rect 3804 4001 3848 4039
rect 3804 3981 3816 4001
rect 3836 3981 3848 4001
rect 3804 3939 3848 3981
rect 3898 4001 3940 4039
rect 3898 3981 3912 4001
rect 3932 3981 3940 4001
rect 3898 3939 3940 3981
rect 4014 4001 4056 4039
rect 4014 3981 4022 4001
rect 4042 3981 4056 4001
rect 4014 3939 4056 3981
rect 4106 4008 4151 4039
rect 4106 4001 4150 4008
rect 4106 3981 4118 4001
rect 4138 3981 4150 4001
rect 4106 3939 4150 3981
rect 11596 4000 11640 4038
rect 11596 3980 11608 4000
rect 11628 3980 11640 4000
rect 8130 3839 8174 3881
rect 8130 3819 8142 3839
rect 8162 3819 8174 3839
rect 8130 3812 8174 3819
rect 8129 3781 8174 3812
rect 8224 3839 8266 3881
rect 8224 3819 8238 3839
rect 8258 3819 8266 3839
rect 8224 3781 8266 3819
rect 8340 3839 8382 3881
rect 8340 3819 8348 3839
rect 8368 3819 8382 3839
rect 8340 3781 8382 3819
rect 8432 3839 8476 3881
rect 8432 3819 8444 3839
rect 8464 3819 8476 3839
rect 8432 3781 8476 3819
rect 8548 3839 8590 3881
rect 8548 3819 8556 3839
rect 8576 3819 8590 3839
rect 8548 3781 8590 3819
rect 8640 3839 8684 3881
rect 8640 3819 8652 3839
rect 8672 3819 8684 3839
rect 8640 3781 8684 3819
rect 8761 3839 8803 3881
rect 8761 3819 8769 3839
rect 8789 3819 8803 3839
rect 8761 3781 8803 3819
rect 8853 3839 8897 3881
rect 11596 3938 11640 3980
rect 11690 4000 11732 4038
rect 11690 3980 11704 4000
rect 11724 3980 11732 4000
rect 11690 3938 11732 3980
rect 11809 4000 11853 4038
rect 11809 3980 11821 4000
rect 11841 3980 11853 4000
rect 11809 3938 11853 3980
rect 11903 4000 11945 4038
rect 11903 3980 11917 4000
rect 11937 3980 11945 4000
rect 11903 3938 11945 3980
rect 12017 4000 12061 4038
rect 12017 3980 12029 4000
rect 12049 3980 12061 4000
rect 12017 3938 12061 3980
rect 12111 4000 12153 4038
rect 12111 3980 12125 4000
rect 12145 3980 12153 4000
rect 12111 3938 12153 3980
rect 12227 4000 12269 4038
rect 12227 3980 12235 4000
rect 12255 3980 12269 4000
rect 12227 3938 12269 3980
rect 12319 4007 12364 4038
rect 12319 4000 12363 4007
rect 12319 3980 12331 4000
rect 12351 3980 12363 4000
rect 12319 3938 12363 3980
rect 14091 3995 14135 4033
rect 14091 3975 14103 3995
rect 14123 3975 14135 3995
rect 8853 3819 8865 3839
rect 8885 3819 8897 3839
rect 8853 3781 8897 3819
rect 9178 3835 9222 3877
rect 9178 3815 9190 3835
rect 9210 3815 9222 3835
rect 9178 3808 9222 3815
rect 9177 3777 9222 3808
rect 9272 3835 9314 3877
rect 9272 3815 9286 3835
rect 9306 3815 9314 3835
rect 9272 3777 9314 3815
rect 9388 3835 9430 3877
rect 9388 3815 9396 3835
rect 9416 3815 9430 3835
rect 9388 3777 9430 3815
rect 9480 3835 9524 3877
rect 9480 3815 9492 3835
rect 9512 3815 9524 3835
rect 9480 3777 9524 3815
rect 9596 3835 9638 3877
rect 9596 3815 9604 3835
rect 9624 3815 9638 3835
rect 9596 3777 9638 3815
rect 9688 3835 9732 3877
rect 9688 3815 9700 3835
rect 9720 3815 9732 3835
rect 9688 3777 9732 3815
rect 9809 3835 9851 3877
rect 9809 3815 9817 3835
rect 9837 3815 9851 3835
rect 9809 3777 9851 3815
rect 9901 3835 9945 3877
rect 9901 3815 9913 3835
rect 9933 3815 9945 3835
rect 14091 3933 14135 3975
rect 14185 3995 14227 4033
rect 14185 3975 14199 3995
rect 14219 3975 14227 3995
rect 14185 3933 14227 3975
rect 14304 3995 14348 4033
rect 14304 3975 14316 3995
rect 14336 3975 14348 3995
rect 14304 3933 14348 3975
rect 14398 3995 14440 4033
rect 14398 3975 14412 3995
rect 14432 3975 14440 3995
rect 14398 3933 14440 3975
rect 14512 3995 14556 4033
rect 14512 3975 14524 3995
rect 14544 3975 14556 3995
rect 14512 3933 14556 3975
rect 14606 3995 14648 4033
rect 14606 3975 14620 3995
rect 14640 3975 14648 3995
rect 14606 3933 14648 3975
rect 14722 3995 14764 4033
rect 14722 3975 14730 3995
rect 14750 3975 14764 3995
rect 14722 3933 14764 3975
rect 14814 4002 14859 4033
rect 14814 3995 14858 4002
rect 14814 3975 14826 3995
rect 14846 3975 14858 3995
rect 14814 3933 14858 3975
rect 9901 3777 9945 3815
rect 22561 4004 22605 4042
rect 22561 3984 22573 4004
rect 22593 3984 22605 4004
rect 18838 3833 18882 3875
rect 18838 3813 18850 3833
rect 18870 3813 18882 3833
rect 18838 3806 18882 3813
rect 18837 3775 18882 3806
rect 18932 3833 18974 3875
rect 18932 3813 18946 3833
rect 18966 3813 18974 3833
rect 18932 3775 18974 3813
rect 19048 3833 19090 3875
rect 19048 3813 19056 3833
rect 19076 3813 19090 3833
rect 19048 3775 19090 3813
rect 19140 3833 19184 3875
rect 19140 3813 19152 3833
rect 19172 3813 19184 3833
rect 19140 3775 19184 3813
rect 19256 3833 19298 3875
rect 19256 3813 19264 3833
rect 19284 3813 19298 3833
rect 19256 3775 19298 3813
rect 19348 3833 19392 3875
rect 19348 3813 19360 3833
rect 19380 3813 19392 3833
rect 19348 3775 19392 3813
rect 19469 3833 19511 3875
rect 19469 3813 19477 3833
rect 19497 3813 19511 3833
rect 19469 3775 19511 3813
rect 19561 3833 19605 3875
rect 22561 3942 22605 3984
rect 22655 4004 22697 4042
rect 22655 3984 22669 4004
rect 22689 3984 22697 4004
rect 22655 3942 22697 3984
rect 22774 4004 22818 4042
rect 22774 3984 22786 4004
rect 22806 3984 22818 4004
rect 22774 3942 22818 3984
rect 22868 4004 22910 4042
rect 22868 3984 22882 4004
rect 22902 3984 22910 4004
rect 22868 3942 22910 3984
rect 22982 4004 23026 4042
rect 22982 3984 22994 4004
rect 23014 3984 23026 4004
rect 22982 3942 23026 3984
rect 23076 4004 23118 4042
rect 23076 3984 23090 4004
rect 23110 3984 23118 4004
rect 23076 3942 23118 3984
rect 23192 4004 23234 4042
rect 23192 3984 23200 4004
rect 23220 3984 23234 4004
rect 23192 3942 23234 3984
rect 23284 4011 23329 4042
rect 23284 4004 23328 4011
rect 23284 3984 23296 4004
rect 23316 3984 23328 4004
rect 23284 3942 23328 3984
rect 25056 3999 25100 4037
rect 25056 3979 25068 3999
rect 25088 3979 25100 3999
rect 19561 3813 19573 3833
rect 19593 3813 19605 3833
rect 19561 3775 19605 3813
rect 19886 3829 19930 3871
rect 19886 3809 19898 3829
rect 19918 3809 19930 3829
rect 19886 3802 19930 3809
rect 19885 3771 19930 3802
rect 19980 3829 20022 3871
rect 19980 3809 19994 3829
rect 20014 3809 20022 3829
rect 19980 3771 20022 3809
rect 20096 3829 20138 3871
rect 20096 3809 20104 3829
rect 20124 3809 20138 3829
rect 20096 3771 20138 3809
rect 20188 3829 20232 3871
rect 20188 3809 20200 3829
rect 20220 3809 20232 3829
rect 20188 3771 20232 3809
rect 20304 3829 20346 3871
rect 20304 3809 20312 3829
rect 20332 3809 20346 3829
rect 20304 3771 20346 3809
rect 20396 3829 20440 3871
rect 20396 3809 20408 3829
rect 20428 3809 20440 3829
rect 20396 3771 20440 3809
rect 20517 3829 20559 3871
rect 20517 3809 20525 3829
rect 20545 3809 20559 3829
rect 20517 3771 20559 3809
rect 20609 3829 20653 3871
rect 20609 3809 20621 3829
rect 20641 3809 20653 3829
rect 25056 3937 25100 3979
rect 25150 3999 25192 4037
rect 25150 3979 25164 3999
rect 25184 3979 25192 3999
rect 25150 3937 25192 3979
rect 25269 3999 25313 4037
rect 25269 3979 25281 3999
rect 25301 3979 25313 3999
rect 25269 3937 25313 3979
rect 25363 3999 25405 4037
rect 25363 3979 25377 3999
rect 25397 3979 25405 3999
rect 25363 3937 25405 3979
rect 25477 3999 25521 4037
rect 25477 3979 25489 3999
rect 25509 3979 25521 3999
rect 25477 3937 25521 3979
rect 25571 3999 25613 4037
rect 25571 3979 25585 3999
rect 25605 3979 25613 3999
rect 25571 3937 25613 3979
rect 25687 3999 25729 4037
rect 25687 3979 25695 3999
rect 25715 3979 25729 3999
rect 25687 3937 25729 3979
rect 25779 4006 25824 4037
rect 25779 3999 25823 4006
rect 25779 3979 25791 3999
rect 25811 3979 25823 3999
rect 25779 3937 25823 3979
rect 33269 3998 33313 4036
rect 33269 3978 33281 3998
rect 33301 3978 33313 3998
rect 20609 3771 20653 3809
rect 29803 3837 29847 3879
rect 29803 3817 29815 3837
rect 29835 3817 29847 3837
rect 29803 3810 29847 3817
rect 29802 3779 29847 3810
rect 29897 3837 29939 3879
rect 29897 3817 29911 3837
rect 29931 3817 29939 3837
rect 29897 3779 29939 3817
rect 30013 3837 30055 3879
rect 30013 3817 30021 3837
rect 30041 3817 30055 3837
rect 30013 3779 30055 3817
rect 30105 3837 30149 3879
rect 30105 3817 30117 3837
rect 30137 3817 30149 3837
rect 30105 3779 30149 3817
rect 30221 3837 30263 3879
rect 30221 3817 30229 3837
rect 30249 3817 30263 3837
rect 30221 3779 30263 3817
rect 30313 3837 30357 3879
rect 30313 3817 30325 3837
rect 30345 3817 30357 3837
rect 30313 3779 30357 3817
rect 30434 3837 30476 3879
rect 30434 3817 30442 3837
rect 30462 3817 30476 3837
rect 30434 3779 30476 3817
rect 30526 3837 30570 3879
rect 33269 3936 33313 3978
rect 33363 3998 33405 4036
rect 33363 3978 33377 3998
rect 33397 3978 33405 3998
rect 33363 3936 33405 3978
rect 33482 3998 33526 4036
rect 33482 3978 33494 3998
rect 33514 3978 33526 3998
rect 33482 3936 33526 3978
rect 33576 3998 33618 4036
rect 33576 3978 33590 3998
rect 33610 3978 33618 3998
rect 33576 3936 33618 3978
rect 33690 3998 33734 4036
rect 33690 3978 33702 3998
rect 33722 3978 33734 3998
rect 33690 3936 33734 3978
rect 33784 3998 33826 4036
rect 33784 3978 33798 3998
rect 33818 3978 33826 3998
rect 33784 3936 33826 3978
rect 33900 3998 33942 4036
rect 33900 3978 33908 3998
rect 33928 3978 33942 3998
rect 33900 3936 33942 3978
rect 33992 4005 34037 4036
rect 33992 3998 34036 4005
rect 33992 3978 34004 3998
rect 34024 3978 34036 3998
rect 33992 3936 34036 3978
rect 35764 3993 35808 4031
rect 35764 3973 35776 3993
rect 35796 3973 35808 3993
rect 30526 3817 30538 3837
rect 30558 3817 30570 3837
rect 30526 3779 30570 3817
rect 30851 3833 30895 3875
rect 30851 3813 30863 3833
rect 30883 3813 30895 3833
rect 30851 3806 30895 3813
rect 30850 3775 30895 3806
rect 30945 3833 30987 3875
rect 30945 3813 30959 3833
rect 30979 3813 30987 3833
rect 30945 3775 30987 3813
rect 31061 3833 31103 3875
rect 31061 3813 31069 3833
rect 31089 3813 31103 3833
rect 31061 3775 31103 3813
rect 31153 3833 31197 3875
rect 31153 3813 31165 3833
rect 31185 3813 31197 3833
rect 31153 3775 31197 3813
rect 31269 3833 31311 3875
rect 31269 3813 31277 3833
rect 31297 3813 31311 3833
rect 31269 3775 31311 3813
rect 31361 3833 31405 3875
rect 31361 3813 31373 3833
rect 31393 3813 31405 3833
rect 31361 3775 31405 3813
rect 31482 3833 31524 3875
rect 31482 3813 31490 3833
rect 31510 3813 31524 3833
rect 31482 3775 31524 3813
rect 31574 3833 31618 3875
rect 31574 3813 31586 3833
rect 31606 3813 31618 3833
rect 35764 3931 35808 3973
rect 35858 3993 35900 4031
rect 35858 3973 35872 3993
rect 35892 3973 35900 3993
rect 35858 3931 35900 3973
rect 35977 3993 36021 4031
rect 35977 3973 35989 3993
rect 36009 3973 36021 3993
rect 35977 3931 36021 3973
rect 36071 3993 36113 4031
rect 36071 3973 36085 3993
rect 36105 3973 36113 3993
rect 36071 3931 36113 3973
rect 36185 3993 36229 4031
rect 36185 3973 36197 3993
rect 36217 3973 36229 3993
rect 36185 3931 36229 3973
rect 36279 3993 36321 4031
rect 36279 3973 36293 3993
rect 36313 3973 36321 3993
rect 36279 3931 36321 3973
rect 36395 3993 36437 4031
rect 36395 3973 36403 3993
rect 36423 3973 36437 3993
rect 36395 3931 36437 3973
rect 36487 4000 36532 4031
rect 36487 3993 36531 4000
rect 36487 3973 36499 3993
rect 36519 3973 36531 3993
rect 36487 3931 36531 3973
rect 31574 3775 31618 3813
rect 40511 3831 40555 3873
rect 40511 3811 40523 3831
rect 40543 3811 40555 3831
rect 40511 3804 40555 3811
rect 40510 3773 40555 3804
rect 40605 3831 40647 3873
rect 40605 3811 40619 3831
rect 40639 3811 40647 3831
rect 40605 3773 40647 3811
rect 40721 3831 40763 3873
rect 40721 3811 40729 3831
rect 40749 3811 40763 3831
rect 40721 3773 40763 3811
rect 40813 3831 40857 3873
rect 40813 3811 40825 3831
rect 40845 3811 40857 3831
rect 40813 3773 40857 3811
rect 40929 3831 40971 3873
rect 40929 3811 40937 3831
rect 40957 3811 40971 3831
rect 40929 3773 40971 3811
rect 41021 3831 41065 3873
rect 41021 3811 41033 3831
rect 41053 3811 41065 3831
rect 41021 3773 41065 3811
rect 41142 3831 41184 3873
rect 41142 3811 41150 3831
rect 41170 3811 41184 3831
rect 41142 3773 41184 3811
rect 41234 3831 41278 3873
rect 41234 3811 41246 3831
rect 41266 3811 41278 3831
rect 41234 3773 41278 3811
rect 41559 3827 41603 3869
rect 41559 3807 41571 3827
rect 41591 3807 41603 3827
rect 41559 3800 41603 3807
rect 41558 3769 41603 3800
rect 41653 3827 41695 3869
rect 41653 3807 41667 3827
rect 41687 3807 41695 3827
rect 41653 3769 41695 3807
rect 41769 3827 41811 3869
rect 41769 3807 41777 3827
rect 41797 3807 41811 3827
rect 41769 3769 41811 3807
rect 41861 3827 41905 3869
rect 41861 3807 41873 3827
rect 41893 3807 41905 3827
rect 41861 3769 41905 3807
rect 41977 3827 42019 3869
rect 41977 3807 41985 3827
rect 42005 3807 42019 3827
rect 41977 3769 42019 3807
rect 42069 3827 42113 3869
rect 42069 3807 42081 3827
rect 42101 3807 42113 3827
rect 42069 3769 42113 3807
rect 42190 3827 42232 3869
rect 42190 3807 42198 3827
rect 42218 3807 42232 3827
rect 42190 3769 42232 3807
rect 42282 3827 42326 3869
rect 42282 3807 42294 3827
rect 42314 3807 42326 3827
rect 42282 3769 42326 3807
rect 888 3238 932 3276
rect 888 3218 900 3238
rect 920 3218 932 3238
rect 888 3176 932 3218
rect 982 3238 1024 3276
rect 982 3218 996 3238
rect 1016 3218 1024 3238
rect 982 3176 1024 3218
rect 1101 3238 1145 3276
rect 1101 3218 1113 3238
rect 1133 3218 1145 3238
rect 1101 3176 1145 3218
rect 1195 3238 1237 3276
rect 1195 3218 1209 3238
rect 1229 3218 1237 3238
rect 1195 3176 1237 3218
rect 1309 3238 1353 3276
rect 1309 3218 1321 3238
rect 1341 3218 1353 3238
rect 1309 3176 1353 3218
rect 1403 3238 1445 3276
rect 1403 3218 1417 3238
rect 1437 3218 1445 3238
rect 1403 3176 1445 3218
rect 1519 3238 1561 3276
rect 1519 3218 1527 3238
rect 1547 3218 1561 3238
rect 1519 3176 1561 3218
rect 1611 3245 1656 3276
rect 1611 3238 1655 3245
rect 1611 3218 1623 3238
rect 1643 3218 1655 3238
rect 1611 3176 1655 3218
rect 1936 3234 1980 3272
rect 1936 3214 1948 3234
rect 1968 3214 1980 3234
rect 1936 3172 1980 3214
rect 2030 3234 2072 3272
rect 2030 3214 2044 3234
rect 2064 3214 2072 3234
rect 2030 3172 2072 3214
rect 2149 3234 2193 3272
rect 2149 3214 2161 3234
rect 2181 3214 2193 3234
rect 2149 3172 2193 3214
rect 2243 3234 2285 3272
rect 2243 3214 2257 3234
rect 2277 3214 2285 3234
rect 2243 3172 2285 3214
rect 2357 3234 2401 3272
rect 2357 3214 2369 3234
rect 2389 3214 2401 3234
rect 2357 3172 2401 3214
rect 2451 3234 2493 3272
rect 2451 3214 2465 3234
rect 2485 3214 2493 3234
rect 2451 3172 2493 3214
rect 2567 3234 2609 3272
rect 2567 3214 2575 3234
rect 2595 3214 2609 3234
rect 2567 3172 2609 3214
rect 2659 3241 2704 3272
rect 2659 3234 2703 3241
rect 2659 3214 2671 3234
rect 2691 3214 2703 3234
rect 2659 3172 2703 3214
rect 11596 3232 11640 3270
rect 6683 3072 6727 3114
rect 6683 3052 6695 3072
rect 6715 3052 6727 3072
rect 6683 3045 6727 3052
rect 6682 3014 6727 3045
rect 6777 3072 6819 3114
rect 6777 3052 6791 3072
rect 6811 3052 6819 3072
rect 6777 3014 6819 3052
rect 6893 3072 6935 3114
rect 6893 3052 6901 3072
rect 6921 3052 6935 3072
rect 6893 3014 6935 3052
rect 6985 3072 7029 3114
rect 6985 3052 6997 3072
rect 7017 3052 7029 3072
rect 6985 3014 7029 3052
rect 7101 3072 7143 3114
rect 7101 3052 7109 3072
rect 7129 3052 7143 3072
rect 7101 3014 7143 3052
rect 7193 3072 7237 3114
rect 7193 3052 7205 3072
rect 7225 3052 7237 3072
rect 7193 3014 7237 3052
rect 7314 3072 7356 3114
rect 7314 3052 7322 3072
rect 7342 3052 7356 3072
rect 7314 3014 7356 3052
rect 7406 3072 7450 3114
rect 11596 3212 11608 3232
rect 11628 3212 11640 3232
rect 11596 3170 11640 3212
rect 11690 3232 11732 3270
rect 11690 3212 11704 3232
rect 11724 3212 11732 3232
rect 11690 3170 11732 3212
rect 11809 3232 11853 3270
rect 11809 3212 11821 3232
rect 11841 3212 11853 3232
rect 11809 3170 11853 3212
rect 11903 3232 11945 3270
rect 11903 3212 11917 3232
rect 11937 3212 11945 3232
rect 11903 3170 11945 3212
rect 12017 3232 12061 3270
rect 12017 3212 12029 3232
rect 12049 3212 12061 3232
rect 12017 3170 12061 3212
rect 12111 3232 12153 3270
rect 12111 3212 12125 3232
rect 12145 3212 12153 3232
rect 12111 3170 12153 3212
rect 12227 3232 12269 3270
rect 12227 3212 12235 3232
rect 12255 3212 12269 3232
rect 12227 3170 12269 3212
rect 12319 3239 12364 3270
rect 12319 3232 12363 3239
rect 12319 3212 12331 3232
rect 12351 3212 12363 3232
rect 12319 3170 12363 3212
rect 12644 3228 12688 3266
rect 12644 3208 12656 3228
rect 12676 3208 12688 3228
rect 7406 3052 7418 3072
rect 7438 3052 7450 3072
rect 7406 3014 7450 3052
rect 9178 3067 9222 3109
rect 9178 3047 9190 3067
rect 9210 3047 9222 3067
rect 9178 3040 9222 3047
rect 9177 3009 9222 3040
rect 9272 3067 9314 3109
rect 9272 3047 9286 3067
rect 9306 3047 9314 3067
rect 9272 3009 9314 3047
rect 9388 3067 9430 3109
rect 9388 3047 9396 3067
rect 9416 3047 9430 3067
rect 9388 3009 9430 3047
rect 9480 3067 9524 3109
rect 9480 3047 9492 3067
rect 9512 3047 9524 3067
rect 9480 3009 9524 3047
rect 9596 3067 9638 3109
rect 9596 3047 9604 3067
rect 9624 3047 9638 3067
rect 9596 3009 9638 3047
rect 9688 3067 9732 3109
rect 9688 3047 9700 3067
rect 9720 3047 9732 3067
rect 9688 3009 9732 3047
rect 9809 3067 9851 3109
rect 9809 3047 9817 3067
rect 9837 3047 9851 3067
rect 9809 3009 9851 3047
rect 9901 3067 9945 3109
rect 12644 3166 12688 3208
rect 12738 3228 12780 3266
rect 12738 3208 12752 3228
rect 12772 3208 12780 3228
rect 12738 3166 12780 3208
rect 12857 3228 12901 3266
rect 12857 3208 12869 3228
rect 12889 3208 12901 3228
rect 12857 3166 12901 3208
rect 12951 3228 12993 3266
rect 12951 3208 12965 3228
rect 12985 3208 12993 3228
rect 12951 3166 12993 3208
rect 13065 3228 13109 3266
rect 13065 3208 13077 3228
rect 13097 3208 13109 3228
rect 13065 3166 13109 3208
rect 13159 3228 13201 3266
rect 13159 3208 13173 3228
rect 13193 3208 13201 3228
rect 13159 3166 13201 3208
rect 13275 3228 13317 3266
rect 13275 3208 13283 3228
rect 13303 3208 13317 3228
rect 13275 3166 13317 3208
rect 13367 3235 13412 3266
rect 13367 3228 13411 3235
rect 13367 3208 13379 3228
rect 13399 3208 13411 3228
rect 13367 3166 13411 3208
rect 22561 3236 22605 3274
rect 9901 3047 9913 3067
rect 9933 3047 9945 3067
rect 9901 3009 9945 3047
rect 17391 3066 17435 3108
rect 17391 3046 17403 3066
rect 17423 3046 17435 3066
rect 17391 3039 17435 3046
rect 17390 3008 17435 3039
rect 17485 3066 17527 3108
rect 17485 3046 17499 3066
rect 17519 3046 17527 3066
rect 17485 3008 17527 3046
rect 17601 3066 17643 3108
rect 17601 3046 17609 3066
rect 17629 3046 17643 3066
rect 17601 3008 17643 3046
rect 17693 3066 17737 3108
rect 17693 3046 17705 3066
rect 17725 3046 17737 3066
rect 17693 3008 17737 3046
rect 17809 3066 17851 3108
rect 17809 3046 17817 3066
rect 17837 3046 17851 3066
rect 17809 3008 17851 3046
rect 17901 3066 17945 3108
rect 17901 3046 17913 3066
rect 17933 3046 17945 3066
rect 17901 3008 17945 3046
rect 18022 3066 18064 3108
rect 18022 3046 18030 3066
rect 18050 3046 18064 3066
rect 18022 3008 18064 3046
rect 18114 3066 18158 3108
rect 22561 3216 22573 3236
rect 22593 3216 22605 3236
rect 22561 3174 22605 3216
rect 22655 3236 22697 3274
rect 22655 3216 22669 3236
rect 22689 3216 22697 3236
rect 22655 3174 22697 3216
rect 22774 3236 22818 3274
rect 22774 3216 22786 3236
rect 22806 3216 22818 3236
rect 22774 3174 22818 3216
rect 22868 3236 22910 3274
rect 22868 3216 22882 3236
rect 22902 3216 22910 3236
rect 22868 3174 22910 3216
rect 22982 3236 23026 3274
rect 22982 3216 22994 3236
rect 23014 3216 23026 3236
rect 22982 3174 23026 3216
rect 23076 3236 23118 3274
rect 23076 3216 23090 3236
rect 23110 3216 23118 3236
rect 23076 3174 23118 3216
rect 23192 3236 23234 3274
rect 23192 3216 23200 3236
rect 23220 3216 23234 3236
rect 23192 3174 23234 3216
rect 23284 3243 23329 3274
rect 23284 3236 23328 3243
rect 23284 3216 23296 3236
rect 23316 3216 23328 3236
rect 23284 3174 23328 3216
rect 23609 3232 23653 3270
rect 23609 3212 23621 3232
rect 23641 3212 23653 3232
rect 18114 3046 18126 3066
rect 18146 3046 18158 3066
rect 18114 3008 18158 3046
rect 19886 3061 19930 3103
rect 19886 3041 19898 3061
rect 19918 3041 19930 3061
rect 19886 3034 19930 3041
rect 19885 3003 19930 3034
rect 19980 3061 20022 3103
rect 19980 3041 19994 3061
rect 20014 3041 20022 3061
rect 19980 3003 20022 3041
rect 20096 3061 20138 3103
rect 20096 3041 20104 3061
rect 20124 3041 20138 3061
rect 20096 3003 20138 3041
rect 20188 3061 20232 3103
rect 20188 3041 20200 3061
rect 20220 3041 20232 3061
rect 20188 3003 20232 3041
rect 20304 3061 20346 3103
rect 20304 3041 20312 3061
rect 20332 3041 20346 3061
rect 20304 3003 20346 3041
rect 20396 3061 20440 3103
rect 20396 3041 20408 3061
rect 20428 3041 20440 3061
rect 20396 3003 20440 3041
rect 20517 3061 20559 3103
rect 20517 3041 20525 3061
rect 20545 3041 20559 3061
rect 20517 3003 20559 3041
rect 20609 3061 20653 3103
rect 23609 3170 23653 3212
rect 23703 3232 23745 3270
rect 23703 3212 23717 3232
rect 23737 3212 23745 3232
rect 23703 3170 23745 3212
rect 23822 3232 23866 3270
rect 23822 3212 23834 3232
rect 23854 3212 23866 3232
rect 23822 3170 23866 3212
rect 23916 3232 23958 3270
rect 23916 3212 23930 3232
rect 23950 3212 23958 3232
rect 23916 3170 23958 3212
rect 24030 3232 24074 3270
rect 24030 3212 24042 3232
rect 24062 3212 24074 3232
rect 24030 3170 24074 3212
rect 24124 3232 24166 3270
rect 24124 3212 24138 3232
rect 24158 3212 24166 3232
rect 24124 3170 24166 3212
rect 24240 3232 24282 3270
rect 24240 3212 24248 3232
rect 24268 3212 24282 3232
rect 24240 3170 24282 3212
rect 24332 3239 24377 3270
rect 24332 3232 24376 3239
rect 24332 3212 24344 3232
rect 24364 3212 24376 3232
rect 24332 3170 24376 3212
rect 20609 3041 20621 3061
rect 20641 3041 20653 3061
rect 20609 3003 20653 3041
rect 33269 3230 33313 3268
rect 28356 3070 28400 3112
rect 28356 3050 28368 3070
rect 28388 3050 28400 3070
rect 28356 3043 28400 3050
rect 28355 3012 28400 3043
rect 28450 3070 28492 3112
rect 28450 3050 28464 3070
rect 28484 3050 28492 3070
rect 28450 3012 28492 3050
rect 28566 3070 28608 3112
rect 28566 3050 28574 3070
rect 28594 3050 28608 3070
rect 28566 3012 28608 3050
rect 28658 3070 28702 3112
rect 28658 3050 28670 3070
rect 28690 3050 28702 3070
rect 28658 3012 28702 3050
rect 28774 3070 28816 3112
rect 28774 3050 28782 3070
rect 28802 3050 28816 3070
rect 28774 3012 28816 3050
rect 28866 3070 28910 3112
rect 28866 3050 28878 3070
rect 28898 3050 28910 3070
rect 28866 3012 28910 3050
rect 28987 3070 29029 3112
rect 28987 3050 28995 3070
rect 29015 3050 29029 3070
rect 28987 3012 29029 3050
rect 29079 3070 29123 3112
rect 33269 3210 33281 3230
rect 33301 3210 33313 3230
rect 33269 3168 33313 3210
rect 33363 3230 33405 3268
rect 33363 3210 33377 3230
rect 33397 3210 33405 3230
rect 33363 3168 33405 3210
rect 33482 3230 33526 3268
rect 33482 3210 33494 3230
rect 33514 3210 33526 3230
rect 33482 3168 33526 3210
rect 33576 3230 33618 3268
rect 33576 3210 33590 3230
rect 33610 3210 33618 3230
rect 33576 3168 33618 3210
rect 33690 3230 33734 3268
rect 33690 3210 33702 3230
rect 33722 3210 33734 3230
rect 33690 3168 33734 3210
rect 33784 3230 33826 3268
rect 33784 3210 33798 3230
rect 33818 3210 33826 3230
rect 33784 3168 33826 3210
rect 33900 3230 33942 3268
rect 33900 3210 33908 3230
rect 33928 3210 33942 3230
rect 33900 3168 33942 3210
rect 33992 3237 34037 3268
rect 33992 3230 34036 3237
rect 33992 3210 34004 3230
rect 34024 3210 34036 3230
rect 33992 3168 34036 3210
rect 34317 3226 34361 3264
rect 34317 3206 34329 3226
rect 34349 3206 34361 3226
rect 29079 3050 29091 3070
rect 29111 3050 29123 3070
rect 29079 3012 29123 3050
rect 30851 3065 30895 3107
rect 30851 3045 30863 3065
rect 30883 3045 30895 3065
rect 30851 3038 30895 3045
rect 30850 3007 30895 3038
rect 30945 3065 30987 3107
rect 30945 3045 30959 3065
rect 30979 3045 30987 3065
rect 30945 3007 30987 3045
rect 31061 3065 31103 3107
rect 31061 3045 31069 3065
rect 31089 3045 31103 3065
rect 31061 3007 31103 3045
rect 31153 3065 31197 3107
rect 31153 3045 31165 3065
rect 31185 3045 31197 3065
rect 31153 3007 31197 3045
rect 31269 3065 31311 3107
rect 31269 3045 31277 3065
rect 31297 3045 31311 3065
rect 31269 3007 31311 3045
rect 31361 3065 31405 3107
rect 31361 3045 31373 3065
rect 31393 3045 31405 3065
rect 31361 3007 31405 3045
rect 31482 3065 31524 3107
rect 31482 3045 31490 3065
rect 31510 3045 31524 3065
rect 31482 3007 31524 3045
rect 31574 3065 31618 3107
rect 34317 3164 34361 3206
rect 34411 3226 34453 3264
rect 34411 3206 34425 3226
rect 34445 3206 34453 3226
rect 34411 3164 34453 3206
rect 34530 3226 34574 3264
rect 34530 3206 34542 3226
rect 34562 3206 34574 3226
rect 34530 3164 34574 3206
rect 34624 3226 34666 3264
rect 34624 3206 34638 3226
rect 34658 3206 34666 3226
rect 34624 3164 34666 3206
rect 34738 3226 34782 3264
rect 34738 3206 34750 3226
rect 34770 3206 34782 3226
rect 34738 3164 34782 3206
rect 34832 3226 34874 3264
rect 34832 3206 34846 3226
rect 34866 3206 34874 3226
rect 34832 3164 34874 3206
rect 34948 3226 34990 3264
rect 34948 3206 34956 3226
rect 34976 3206 34990 3226
rect 34948 3164 34990 3206
rect 35040 3233 35085 3264
rect 35040 3226 35084 3233
rect 35040 3206 35052 3226
rect 35072 3206 35084 3226
rect 35040 3164 35084 3206
rect 31574 3045 31586 3065
rect 31606 3045 31618 3065
rect 31574 3007 31618 3045
rect 39064 3064 39108 3106
rect 39064 3044 39076 3064
rect 39096 3044 39108 3064
rect 39064 3037 39108 3044
rect 39063 3006 39108 3037
rect 39158 3064 39200 3106
rect 39158 3044 39172 3064
rect 39192 3044 39200 3064
rect 39158 3006 39200 3044
rect 39274 3064 39316 3106
rect 39274 3044 39282 3064
rect 39302 3044 39316 3064
rect 39274 3006 39316 3044
rect 39366 3064 39410 3106
rect 39366 3044 39378 3064
rect 39398 3044 39410 3064
rect 39366 3006 39410 3044
rect 39482 3064 39524 3106
rect 39482 3044 39490 3064
rect 39510 3044 39524 3064
rect 39482 3006 39524 3044
rect 39574 3064 39618 3106
rect 39574 3044 39586 3064
rect 39606 3044 39618 3064
rect 39574 3006 39618 3044
rect 39695 3064 39737 3106
rect 39695 3044 39703 3064
rect 39723 3044 39737 3064
rect 39695 3006 39737 3044
rect 39787 3064 39831 3106
rect 39787 3044 39799 3064
rect 39819 3044 39831 3064
rect 39787 3006 39831 3044
rect 41559 3059 41603 3101
rect 41559 3039 41571 3059
rect 41591 3039 41603 3059
rect 41559 3032 41603 3039
rect 41558 3001 41603 3032
rect 41653 3059 41695 3101
rect 41653 3039 41667 3059
rect 41687 3039 41695 3059
rect 41653 3001 41695 3039
rect 41769 3059 41811 3101
rect 41769 3039 41777 3059
rect 41797 3039 41811 3059
rect 41769 3001 41811 3039
rect 41861 3059 41905 3101
rect 41861 3039 41873 3059
rect 41893 3039 41905 3059
rect 41861 3001 41905 3039
rect 41977 3059 42019 3101
rect 41977 3039 41985 3059
rect 42005 3039 42019 3059
rect 41977 3001 42019 3039
rect 42069 3059 42113 3101
rect 42069 3039 42081 3059
rect 42101 3039 42113 3059
rect 42069 3001 42113 3039
rect 42190 3059 42232 3101
rect 42190 3039 42198 3059
rect 42218 3039 42232 3059
rect 42190 3001 42232 3039
rect 42282 3059 42326 3101
rect 42282 3039 42294 3059
rect 42314 3039 42326 3059
rect 42282 3001 42326 3039
rect 888 2559 932 2597
rect 888 2539 900 2559
rect 920 2539 932 2559
rect 888 2497 932 2539
rect 982 2559 1024 2597
rect 982 2539 996 2559
rect 1016 2539 1024 2559
rect 982 2497 1024 2539
rect 1101 2559 1145 2597
rect 1101 2539 1113 2559
rect 1133 2539 1145 2559
rect 1101 2497 1145 2539
rect 1195 2559 1237 2597
rect 1195 2539 1209 2559
rect 1229 2539 1237 2559
rect 1195 2497 1237 2539
rect 1309 2559 1353 2597
rect 1309 2539 1321 2559
rect 1341 2539 1353 2559
rect 1309 2497 1353 2539
rect 1403 2559 1445 2597
rect 1403 2539 1417 2559
rect 1437 2539 1445 2559
rect 1403 2497 1445 2539
rect 1519 2559 1561 2597
rect 1519 2539 1527 2559
rect 1547 2539 1561 2559
rect 1519 2497 1561 2539
rect 1611 2566 1656 2597
rect 1611 2559 1655 2566
rect 1611 2539 1623 2559
rect 1643 2539 1655 2559
rect 1611 2497 1655 2539
rect 11596 2553 11640 2591
rect 11596 2533 11608 2553
rect 11628 2533 11640 2553
rect 8130 2392 8174 2434
rect 8130 2372 8142 2392
rect 8162 2372 8174 2392
rect 8130 2365 8174 2372
rect 8129 2334 8174 2365
rect 8224 2392 8266 2434
rect 8224 2372 8238 2392
rect 8258 2372 8266 2392
rect 8224 2334 8266 2372
rect 8340 2392 8382 2434
rect 8340 2372 8348 2392
rect 8368 2372 8382 2392
rect 8340 2334 8382 2372
rect 8432 2392 8476 2434
rect 8432 2372 8444 2392
rect 8464 2372 8476 2392
rect 8432 2334 8476 2372
rect 8548 2392 8590 2434
rect 8548 2372 8556 2392
rect 8576 2372 8590 2392
rect 8548 2334 8590 2372
rect 8640 2392 8684 2434
rect 8640 2372 8652 2392
rect 8672 2372 8684 2392
rect 8640 2334 8684 2372
rect 8761 2392 8803 2434
rect 8761 2372 8769 2392
rect 8789 2372 8803 2392
rect 8761 2334 8803 2372
rect 8853 2392 8897 2434
rect 11596 2491 11640 2533
rect 11690 2553 11732 2591
rect 11690 2533 11704 2553
rect 11724 2533 11732 2553
rect 11690 2491 11732 2533
rect 11809 2553 11853 2591
rect 11809 2533 11821 2553
rect 11841 2533 11853 2553
rect 11809 2491 11853 2533
rect 11903 2553 11945 2591
rect 11903 2533 11917 2553
rect 11937 2533 11945 2553
rect 11903 2491 11945 2533
rect 12017 2553 12061 2591
rect 12017 2533 12029 2553
rect 12049 2533 12061 2553
rect 12017 2491 12061 2533
rect 12111 2553 12153 2591
rect 12111 2533 12125 2553
rect 12145 2533 12153 2553
rect 12111 2491 12153 2533
rect 12227 2553 12269 2591
rect 12227 2533 12235 2553
rect 12255 2533 12269 2553
rect 12227 2491 12269 2533
rect 12319 2560 12364 2591
rect 12319 2553 12363 2560
rect 12319 2533 12331 2553
rect 12351 2533 12363 2553
rect 12319 2491 12363 2533
rect 8853 2372 8865 2392
rect 8885 2372 8897 2392
rect 8853 2334 8897 2372
rect 9178 2388 9222 2430
rect 9178 2368 9190 2388
rect 9210 2368 9222 2388
rect 9178 2361 9222 2368
rect 9177 2330 9222 2361
rect 9272 2388 9314 2430
rect 9272 2368 9286 2388
rect 9306 2368 9314 2388
rect 9272 2330 9314 2368
rect 9388 2388 9430 2430
rect 9388 2368 9396 2388
rect 9416 2368 9430 2388
rect 9388 2330 9430 2368
rect 9480 2388 9524 2430
rect 9480 2368 9492 2388
rect 9512 2368 9524 2388
rect 9480 2330 9524 2368
rect 9596 2388 9638 2430
rect 9596 2368 9604 2388
rect 9624 2368 9638 2388
rect 9596 2330 9638 2368
rect 9688 2388 9732 2430
rect 9688 2368 9700 2388
rect 9720 2368 9732 2388
rect 9688 2330 9732 2368
rect 9809 2388 9851 2430
rect 9809 2368 9817 2388
rect 9837 2368 9851 2388
rect 9809 2330 9851 2368
rect 9901 2388 9945 2430
rect 9901 2368 9913 2388
rect 9933 2368 9945 2388
rect 22561 2557 22605 2595
rect 22561 2537 22573 2557
rect 22593 2537 22605 2557
rect 9901 2330 9945 2368
rect 18838 2386 18882 2428
rect 18838 2366 18850 2386
rect 18870 2366 18882 2386
rect 18838 2359 18882 2366
rect 18837 2328 18882 2359
rect 18932 2386 18974 2428
rect 18932 2366 18946 2386
rect 18966 2366 18974 2386
rect 18932 2328 18974 2366
rect 19048 2386 19090 2428
rect 19048 2366 19056 2386
rect 19076 2366 19090 2386
rect 19048 2328 19090 2366
rect 19140 2386 19184 2428
rect 19140 2366 19152 2386
rect 19172 2366 19184 2386
rect 19140 2328 19184 2366
rect 19256 2386 19298 2428
rect 19256 2366 19264 2386
rect 19284 2366 19298 2386
rect 19256 2328 19298 2366
rect 19348 2386 19392 2428
rect 19348 2366 19360 2386
rect 19380 2366 19392 2386
rect 19348 2328 19392 2366
rect 19469 2386 19511 2428
rect 19469 2366 19477 2386
rect 19497 2366 19511 2386
rect 19469 2328 19511 2366
rect 19561 2386 19605 2428
rect 22561 2495 22605 2537
rect 22655 2557 22697 2595
rect 22655 2537 22669 2557
rect 22689 2537 22697 2557
rect 22655 2495 22697 2537
rect 22774 2557 22818 2595
rect 22774 2537 22786 2557
rect 22806 2537 22818 2557
rect 22774 2495 22818 2537
rect 22868 2557 22910 2595
rect 22868 2537 22882 2557
rect 22902 2537 22910 2557
rect 22868 2495 22910 2537
rect 22982 2557 23026 2595
rect 22982 2537 22994 2557
rect 23014 2537 23026 2557
rect 22982 2495 23026 2537
rect 23076 2557 23118 2595
rect 23076 2537 23090 2557
rect 23110 2537 23118 2557
rect 23076 2495 23118 2537
rect 23192 2557 23234 2595
rect 23192 2537 23200 2557
rect 23220 2537 23234 2557
rect 23192 2495 23234 2537
rect 23284 2564 23329 2595
rect 23284 2557 23328 2564
rect 23284 2537 23296 2557
rect 23316 2537 23328 2557
rect 23284 2495 23328 2537
rect 19561 2366 19573 2386
rect 19593 2366 19605 2386
rect 19561 2328 19605 2366
rect 19886 2382 19930 2424
rect 19886 2362 19898 2382
rect 19918 2362 19930 2382
rect 19886 2355 19930 2362
rect 19885 2324 19930 2355
rect 19980 2382 20022 2424
rect 19980 2362 19994 2382
rect 20014 2362 20022 2382
rect 19980 2324 20022 2362
rect 20096 2382 20138 2424
rect 20096 2362 20104 2382
rect 20124 2362 20138 2382
rect 20096 2324 20138 2362
rect 20188 2382 20232 2424
rect 20188 2362 20200 2382
rect 20220 2362 20232 2382
rect 20188 2324 20232 2362
rect 20304 2382 20346 2424
rect 20304 2362 20312 2382
rect 20332 2362 20346 2382
rect 20304 2324 20346 2362
rect 20396 2382 20440 2424
rect 20396 2362 20408 2382
rect 20428 2362 20440 2382
rect 20396 2324 20440 2362
rect 20517 2382 20559 2424
rect 20517 2362 20525 2382
rect 20545 2362 20559 2382
rect 20517 2324 20559 2362
rect 20609 2382 20653 2424
rect 20609 2362 20621 2382
rect 20641 2362 20653 2382
rect 33269 2551 33313 2589
rect 33269 2531 33281 2551
rect 33301 2531 33313 2551
rect 29803 2390 29847 2432
rect 20609 2324 20653 2362
rect 29803 2370 29815 2390
rect 29835 2370 29847 2390
rect 29803 2363 29847 2370
rect 29802 2332 29847 2363
rect 29897 2390 29939 2432
rect 29897 2370 29911 2390
rect 29931 2370 29939 2390
rect 29897 2332 29939 2370
rect 30013 2390 30055 2432
rect 30013 2370 30021 2390
rect 30041 2370 30055 2390
rect 30013 2332 30055 2370
rect 30105 2390 30149 2432
rect 30105 2370 30117 2390
rect 30137 2370 30149 2390
rect 30105 2332 30149 2370
rect 30221 2390 30263 2432
rect 30221 2370 30229 2390
rect 30249 2370 30263 2390
rect 30221 2332 30263 2370
rect 30313 2390 30357 2432
rect 30313 2370 30325 2390
rect 30345 2370 30357 2390
rect 30313 2332 30357 2370
rect 30434 2390 30476 2432
rect 30434 2370 30442 2390
rect 30462 2370 30476 2390
rect 30434 2332 30476 2370
rect 30526 2390 30570 2432
rect 33269 2489 33313 2531
rect 33363 2551 33405 2589
rect 33363 2531 33377 2551
rect 33397 2531 33405 2551
rect 33363 2489 33405 2531
rect 33482 2551 33526 2589
rect 33482 2531 33494 2551
rect 33514 2531 33526 2551
rect 33482 2489 33526 2531
rect 33576 2551 33618 2589
rect 33576 2531 33590 2551
rect 33610 2531 33618 2551
rect 33576 2489 33618 2531
rect 33690 2551 33734 2589
rect 33690 2531 33702 2551
rect 33722 2531 33734 2551
rect 33690 2489 33734 2531
rect 33784 2551 33826 2589
rect 33784 2531 33798 2551
rect 33818 2531 33826 2551
rect 33784 2489 33826 2531
rect 33900 2551 33942 2589
rect 33900 2531 33908 2551
rect 33928 2531 33942 2551
rect 33900 2489 33942 2531
rect 33992 2558 34037 2589
rect 33992 2551 34036 2558
rect 33992 2531 34004 2551
rect 34024 2531 34036 2551
rect 33992 2489 34036 2531
rect 30526 2370 30538 2390
rect 30558 2370 30570 2390
rect 30526 2332 30570 2370
rect 30851 2386 30895 2428
rect 30851 2366 30863 2386
rect 30883 2366 30895 2386
rect 30851 2359 30895 2366
rect 30850 2328 30895 2359
rect 30945 2386 30987 2428
rect 30945 2366 30959 2386
rect 30979 2366 30987 2386
rect 30945 2328 30987 2366
rect 31061 2386 31103 2428
rect 31061 2366 31069 2386
rect 31089 2366 31103 2386
rect 31061 2328 31103 2366
rect 31153 2386 31197 2428
rect 31153 2366 31165 2386
rect 31185 2366 31197 2386
rect 31153 2328 31197 2366
rect 31269 2386 31311 2428
rect 31269 2366 31277 2386
rect 31297 2366 31311 2386
rect 31269 2328 31311 2366
rect 31361 2386 31405 2428
rect 31361 2366 31373 2386
rect 31393 2366 31405 2386
rect 31361 2328 31405 2366
rect 31482 2386 31524 2428
rect 31482 2366 31490 2386
rect 31510 2366 31524 2386
rect 31482 2328 31524 2366
rect 31574 2386 31618 2428
rect 31574 2366 31586 2386
rect 31606 2366 31618 2386
rect 31574 2328 31618 2366
rect 40511 2384 40555 2426
rect 40511 2364 40523 2384
rect 40543 2364 40555 2384
rect 40511 2357 40555 2364
rect 40510 2326 40555 2357
rect 40605 2384 40647 2426
rect 40605 2364 40619 2384
rect 40639 2364 40647 2384
rect 40605 2326 40647 2364
rect 40721 2384 40763 2426
rect 40721 2364 40729 2384
rect 40749 2364 40763 2384
rect 40721 2326 40763 2364
rect 40813 2384 40857 2426
rect 40813 2364 40825 2384
rect 40845 2364 40857 2384
rect 40813 2326 40857 2364
rect 40929 2384 40971 2426
rect 40929 2364 40937 2384
rect 40957 2364 40971 2384
rect 40929 2326 40971 2364
rect 41021 2384 41065 2426
rect 41021 2364 41033 2384
rect 41053 2364 41065 2384
rect 41021 2326 41065 2364
rect 41142 2384 41184 2426
rect 41142 2364 41150 2384
rect 41170 2364 41184 2384
rect 41142 2326 41184 2364
rect 41234 2384 41278 2426
rect 41234 2364 41246 2384
rect 41266 2364 41278 2384
rect 41234 2326 41278 2364
rect 41559 2380 41603 2422
rect 41559 2360 41571 2380
rect 41591 2360 41603 2380
rect 41559 2353 41603 2360
rect 41558 2322 41603 2353
rect 41653 2380 41695 2422
rect 41653 2360 41667 2380
rect 41687 2360 41695 2380
rect 41653 2322 41695 2360
rect 41769 2380 41811 2422
rect 41769 2360 41777 2380
rect 41797 2360 41811 2380
rect 41769 2322 41811 2360
rect 41861 2380 41905 2422
rect 41861 2360 41873 2380
rect 41893 2360 41905 2380
rect 41861 2322 41905 2360
rect 41977 2380 42019 2422
rect 41977 2360 41985 2380
rect 42005 2360 42019 2380
rect 41977 2322 42019 2360
rect 42069 2380 42113 2422
rect 42069 2360 42081 2380
rect 42101 2360 42113 2380
rect 42069 2322 42113 2360
rect 42190 2380 42232 2422
rect 42190 2360 42198 2380
rect 42218 2360 42232 2380
rect 42190 2322 42232 2360
rect 42282 2380 42326 2422
rect 42282 2360 42294 2380
rect 42314 2360 42326 2380
rect 42282 2322 42326 2360
rect 10599 400 10643 438
rect 10599 380 10611 400
rect 10631 380 10643 400
rect 10599 338 10643 380
rect 10693 400 10735 438
rect 10693 380 10707 400
rect 10727 380 10735 400
rect 10693 338 10735 380
rect 10812 400 10856 438
rect 10812 380 10824 400
rect 10844 380 10856 400
rect 10812 338 10856 380
rect 10906 400 10948 438
rect 10906 380 10920 400
rect 10940 380 10948 400
rect 10906 338 10948 380
rect 11020 400 11064 438
rect 11020 380 11032 400
rect 11052 380 11064 400
rect 11020 338 11064 380
rect 11114 400 11156 438
rect 11114 380 11128 400
rect 11148 380 11156 400
rect 11114 338 11156 380
rect 11230 400 11272 438
rect 11230 380 11238 400
rect 11258 380 11272 400
rect 11230 338 11272 380
rect 11322 407 11367 438
rect 11322 400 11366 407
rect 11322 380 11334 400
rect 11354 380 11366 400
rect 11322 338 11366 380
rect 21236 387 21280 425
rect 21236 367 21248 387
rect 21268 367 21280 387
rect 21236 325 21280 367
rect 21330 387 21372 425
rect 21330 367 21344 387
rect 21364 367 21372 387
rect 21330 325 21372 367
rect 21449 387 21493 425
rect 21449 367 21461 387
rect 21481 367 21493 387
rect 21449 325 21493 367
rect 21543 387 21585 425
rect 21543 367 21557 387
rect 21577 367 21585 387
rect 21543 325 21585 367
rect 21657 387 21701 425
rect 21657 367 21669 387
rect 21689 367 21701 387
rect 21657 325 21701 367
rect 21751 387 21793 425
rect 21751 367 21765 387
rect 21785 367 21793 387
rect 21751 325 21793 367
rect 21867 387 21909 425
rect 21867 367 21875 387
rect 21895 367 21909 387
rect 21867 325 21909 367
rect 21959 394 22004 425
rect 32272 398 32316 436
rect 21959 387 22003 394
rect 21959 367 21971 387
rect 21991 367 22003 387
rect 21959 325 22003 367
rect 32272 378 32284 398
rect 32304 378 32316 398
rect 32272 336 32316 378
rect 32366 398 32408 436
rect 32366 378 32380 398
rect 32400 378 32408 398
rect 32366 336 32408 378
rect 32485 398 32529 436
rect 32485 378 32497 398
rect 32517 378 32529 398
rect 32485 336 32529 378
rect 32579 398 32621 436
rect 32579 378 32593 398
rect 32613 378 32621 398
rect 32579 336 32621 378
rect 32693 398 32737 436
rect 32693 378 32705 398
rect 32725 378 32737 398
rect 32693 336 32737 378
rect 32787 398 32829 436
rect 32787 378 32801 398
rect 32821 378 32829 398
rect 32787 336 32829 378
rect 32903 398 32945 436
rect 32903 378 32911 398
rect 32931 378 32945 398
rect 32903 336 32945 378
rect 32995 405 33040 436
rect 32995 398 33039 405
rect 32995 378 33007 398
rect 33027 378 33039 398
rect 32995 336 33039 378
<< ndiffc >>
rect 575 13814 593 13832
rect 11283 13808 11301 13826
rect 22248 13812 22266 13830
rect 32956 13806 32974 13824
rect 577 13715 595 13733
rect 11285 13709 11303 13727
rect 575 13558 593 13576
rect 9185 13618 9205 13638
rect 9288 13614 9308 13634
rect 9396 13614 9416 13634
rect 9499 13618 9519 13638
rect 9604 13614 9624 13634
rect 9707 13618 9727 13638
rect 9817 13614 9837 13634
rect 9920 13618 9940 13638
rect 10240 13623 10258 13641
rect 895 13491 915 13511
rect 998 13495 1018 13515
rect 1108 13491 1128 13511
rect 1211 13495 1231 13515
rect 1316 13491 1336 13511
rect 1419 13495 1439 13515
rect 1527 13495 1547 13515
rect 22250 13713 22268 13731
rect 1630 13491 1650 13511
rect 1943 13487 1963 13507
rect 577 13459 595 13477
rect 2046 13491 2066 13511
rect 2156 13487 2176 13507
rect 2259 13491 2279 13511
rect 2364 13487 2384 13507
rect 2467 13491 2487 13511
rect 2575 13491 2595 13511
rect 2678 13487 2698 13507
rect 10242 13524 10260 13542
rect 11283 13552 11301 13570
rect 19893 13612 19913 13632
rect 19996 13608 20016 13628
rect 20104 13608 20124 13628
rect 20207 13612 20227 13632
rect 20312 13608 20332 13628
rect 20415 13612 20435 13632
rect 20525 13608 20545 13628
rect 20628 13612 20648 13632
rect 20948 13617 20966 13635
rect 11603 13485 11623 13505
rect 11706 13489 11726 13509
rect 11816 13485 11836 13505
rect 11919 13489 11939 13509
rect 12024 13485 12044 13505
rect 12127 13489 12147 13509
rect 12235 13489 12255 13509
rect 32958 13707 32976 13725
rect 12338 13485 12358 13505
rect 12651 13481 12671 13501
rect 11285 13453 11303 13471
rect 12754 13485 12774 13505
rect 12864 13481 12884 13501
rect 12967 13485 12987 13505
rect 13072 13481 13092 13501
rect 13175 13485 13195 13505
rect 13283 13485 13303 13505
rect 13386 13481 13406 13501
rect 10240 13368 10258 13386
rect 20950 13518 20968 13536
rect 22248 13556 22266 13574
rect 30858 13616 30878 13636
rect 30961 13612 30981 13632
rect 31069 13612 31089 13632
rect 31172 13616 31192 13636
rect 31277 13612 31297 13632
rect 31380 13616 31400 13636
rect 31490 13612 31510 13632
rect 31593 13616 31613 13636
rect 31913 13621 31931 13639
rect 22568 13489 22588 13509
rect 22671 13493 22691 13513
rect 22781 13489 22801 13509
rect 22884 13493 22904 13513
rect 22989 13489 23009 13509
rect 23092 13493 23112 13513
rect 23200 13493 23220 13513
rect 23303 13489 23323 13509
rect 23616 13485 23636 13505
rect 22250 13457 22268 13475
rect 23719 13489 23739 13509
rect 23829 13485 23849 13505
rect 23932 13489 23952 13509
rect 24037 13485 24057 13505
rect 24140 13489 24160 13509
rect 24248 13489 24268 13509
rect 24351 13485 24371 13505
rect 20948 13362 20966 13380
rect 31915 13522 31933 13540
rect 32956 13550 32974 13568
rect 41566 13610 41586 13630
rect 41669 13606 41689 13626
rect 41777 13606 41797 13626
rect 41880 13610 41900 13630
rect 41985 13606 42005 13626
rect 42088 13610 42108 13630
rect 42198 13606 42218 13626
rect 42301 13610 42321 13630
rect 42621 13615 42639 13633
rect 33276 13483 33296 13503
rect 33379 13487 33399 13507
rect 33489 13483 33509 13503
rect 33592 13487 33612 13507
rect 33697 13483 33717 13503
rect 33800 13487 33820 13507
rect 33908 13487 33928 13507
rect 34011 13483 34031 13503
rect 34324 13479 34344 13499
rect 32958 13451 32976 13469
rect 34427 13483 34447 13503
rect 34537 13479 34557 13499
rect 34640 13483 34660 13503
rect 34745 13479 34765 13499
rect 34848 13483 34868 13503
rect 34956 13483 34976 13503
rect 35059 13479 35079 13499
rect 31913 13366 31931 13384
rect 42623 13516 42641 13534
rect 42621 13360 42639 13378
rect 10242 13269 10260 13287
rect 20950 13263 20968 13281
rect 31915 13267 31933 13285
rect 42623 13261 42641 13279
rect 575 13163 593 13181
rect 11283 13157 11301 13175
rect 22248 13161 22266 13179
rect 32956 13155 32974 13173
rect 577 13064 595 13082
rect 575 12908 593 12926
rect 11285 13058 11303 13076
rect 8137 12943 8157 12963
rect 8240 12939 8260 12959
rect 8348 12939 8368 12959
rect 8451 12943 8471 12963
rect 8556 12939 8576 12959
rect 8659 12943 8679 12963
rect 8769 12939 8789 12959
rect 10240 12973 10258 12991
rect 8872 12943 8892 12963
rect 9185 12939 9205 12959
rect 577 12809 595 12827
rect 895 12812 915 12832
rect 998 12816 1018 12836
rect 1108 12812 1128 12832
rect 1211 12816 1231 12836
rect 1316 12812 1336 12832
rect 1419 12816 1439 12836
rect 1527 12816 1547 12836
rect 9288 12935 9308 12955
rect 9396 12935 9416 12955
rect 9499 12939 9519 12959
rect 9604 12935 9624 12955
rect 9707 12939 9727 12959
rect 9817 12935 9837 12955
rect 9920 12939 9940 12959
rect 1630 12812 1650 12832
rect 3390 12807 3410 12827
rect 3493 12811 3513 12831
rect 3603 12807 3623 12827
rect 3706 12811 3726 12831
rect 3811 12807 3831 12827
rect 3914 12811 3934 12831
rect 4022 12811 4042 12831
rect 4125 12807 4145 12827
rect 10242 12874 10260 12892
rect 11283 12902 11301 12920
rect 22250 13062 22268 13080
rect 18845 12937 18865 12957
rect 18948 12933 18968 12953
rect 19056 12933 19076 12953
rect 19159 12937 19179 12957
rect 19264 12933 19284 12953
rect 19367 12937 19387 12957
rect 19477 12933 19497 12953
rect 20948 12967 20966 12985
rect 19580 12937 19600 12957
rect 19893 12933 19913 12953
rect 11285 12803 11303 12821
rect 11603 12806 11623 12826
rect 11706 12810 11726 12830
rect 11816 12806 11836 12826
rect 11919 12810 11939 12830
rect 12024 12806 12044 12826
rect 12127 12810 12147 12830
rect 12235 12810 12255 12830
rect 19996 12929 20016 12949
rect 20104 12929 20124 12949
rect 20207 12933 20227 12953
rect 20312 12929 20332 12949
rect 20415 12933 20435 12953
rect 20525 12929 20545 12949
rect 20628 12933 20648 12953
rect 12338 12806 12358 12826
rect 14098 12801 14118 12821
rect 14201 12805 14221 12825
rect 14311 12801 14331 12821
rect 14414 12805 14434 12825
rect 14519 12801 14539 12821
rect 14622 12805 14642 12825
rect 14730 12805 14750 12825
rect 14833 12801 14853 12821
rect 20950 12868 20968 12886
rect 22248 12906 22266 12924
rect 32958 13056 32976 13074
rect 10240 12717 10258 12735
rect 29810 12941 29830 12961
rect 29913 12937 29933 12957
rect 30021 12937 30041 12957
rect 30124 12941 30144 12961
rect 30229 12937 30249 12957
rect 30332 12941 30352 12961
rect 30442 12937 30462 12957
rect 31913 12971 31931 12989
rect 30545 12941 30565 12961
rect 30858 12937 30878 12957
rect 22250 12807 22268 12825
rect 22568 12810 22588 12830
rect 22671 12814 22691 12834
rect 22781 12810 22801 12830
rect 22884 12814 22904 12834
rect 22989 12810 23009 12830
rect 23092 12814 23112 12834
rect 23200 12814 23220 12834
rect 30961 12933 30981 12953
rect 31069 12933 31089 12953
rect 31172 12937 31192 12957
rect 31277 12933 31297 12953
rect 31380 12937 31400 12957
rect 31490 12933 31510 12953
rect 31593 12937 31613 12957
rect 23303 12810 23323 12830
rect 25063 12805 25083 12825
rect 25166 12809 25186 12829
rect 25276 12805 25296 12825
rect 25379 12809 25399 12829
rect 25484 12805 25504 12825
rect 25587 12809 25607 12829
rect 25695 12809 25715 12829
rect 25798 12805 25818 12825
rect 31915 12872 31933 12890
rect 32956 12900 32974 12918
rect 20948 12711 20966 12729
rect 40518 12935 40538 12955
rect 40621 12931 40641 12951
rect 40729 12931 40749 12951
rect 40832 12935 40852 12955
rect 40937 12931 40957 12951
rect 41040 12935 41060 12955
rect 41150 12931 41170 12951
rect 42621 12965 42639 12983
rect 41253 12935 41273 12955
rect 41566 12931 41586 12951
rect 32958 12801 32976 12819
rect 33276 12804 33296 12824
rect 33379 12808 33399 12828
rect 33489 12804 33509 12824
rect 33592 12808 33612 12828
rect 33697 12804 33717 12824
rect 33800 12808 33820 12828
rect 33908 12808 33928 12828
rect 41669 12927 41689 12947
rect 41777 12927 41797 12947
rect 41880 12931 41900 12951
rect 41985 12927 42005 12947
rect 42088 12931 42108 12951
rect 42198 12927 42218 12947
rect 42301 12931 42321 12951
rect 34011 12804 34031 12824
rect 35771 12799 35791 12819
rect 35874 12803 35894 12823
rect 35984 12799 36004 12819
rect 36087 12803 36107 12823
rect 36192 12799 36212 12819
rect 36295 12803 36315 12823
rect 36403 12803 36423 12823
rect 36506 12799 36526 12819
rect 42623 12866 42641 12884
rect 31913 12715 31931 12733
rect 42621 12709 42639 12727
rect 10242 12618 10260 12636
rect 20950 12612 20968 12630
rect 31915 12616 31933 12634
rect 42623 12610 42641 12628
rect 575 12367 593 12385
rect 11283 12361 11301 12379
rect 22248 12365 22266 12383
rect 32956 12359 32974 12377
rect 577 12268 595 12286
rect 11285 12262 11303 12280
rect 575 12111 593 12129
rect 6690 12176 6710 12196
rect 6793 12172 6813 12192
rect 6901 12172 6921 12192
rect 7004 12176 7024 12196
rect 7109 12172 7129 12192
rect 7212 12176 7232 12196
rect 7322 12172 7342 12192
rect 7425 12176 7445 12196
rect 9185 12171 9205 12191
rect 895 12044 915 12064
rect 998 12048 1018 12068
rect 1108 12044 1128 12064
rect 1211 12048 1231 12068
rect 1316 12044 1336 12064
rect 1419 12048 1439 12068
rect 1527 12048 1547 12068
rect 9288 12167 9308 12187
rect 9396 12167 9416 12187
rect 9499 12171 9519 12191
rect 9604 12167 9624 12187
rect 9707 12171 9727 12191
rect 9817 12167 9837 12187
rect 9920 12171 9940 12191
rect 10240 12176 10258 12194
rect 1630 12044 1650 12064
rect 1943 12040 1963 12060
rect 577 12012 595 12030
rect 2046 12044 2066 12064
rect 2156 12040 2176 12060
rect 2259 12044 2279 12064
rect 2364 12040 2384 12060
rect 2467 12044 2487 12064
rect 2575 12044 2595 12064
rect 2678 12040 2698 12060
rect 22250 12266 22268 12284
rect 10242 12077 10260 12095
rect 11283 12105 11301 12123
rect 17398 12170 17418 12190
rect 17501 12166 17521 12186
rect 17609 12166 17629 12186
rect 17712 12170 17732 12190
rect 17817 12166 17837 12186
rect 17920 12170 17940 12190
rect 18030 12166 18050 12186
rect 18133 12170 18153 12190
rect 19893 12165 19913 12185
rect 11603 12038 11623 12058
rect 11706 12042 11726 12062
rect 11816 12038 11836 12058
rect 11919 12042 11939 12062
rect 12024 12038 12044 12058
rect 12127 12042 12147 12062
rect 12235 12042 12255 12062
rect 19996 12161 20016 12181
rect 20104 12161 20124 12181
rect 20207 12165 20227 12185
rect 20312 12161 20332 12181
rect 20415 12165 20435 12185
rect 20525 12161 20545 12181
rect 20628 12165 20648 12185
rect 20948 12170 20966 12188
rect 12338 12038 12358 12058
rect 12651 12034 12671 12054
rect 11285 12006 11303 12024
rect 12754 12038 12774 12058
rect 12864 12034 12884 12054
rect 12967 12038 12987 12058
rect 13072 12034 13092 12054
rect 13175 12038 13195 12058
rect 13283 12038 13303 12058
rect 13386 12034 13406 12054
rect 32958 12260 32976 12278
rect 10240 11921 10258 11939
rect 20950 12071 20968 12089
rect 22248 12109 22266 12127
rect 28363 12174 28383 12194
rect 28466 12170 28486 12190
rect 28574 12170 28594 12190
rect 28677 12174 28697 12194
rect 28782 12170 28802 12190
rect 28885 12174 28905 12194
rect 28995 12170 29015 12190
rect 29098 12174 29118 12194
rect 30858 12169 30878 12189
rect 22568 12042 22588 12062
rect 22671 12046 22691 12066
rect 22781 12042 22801 12062
rect 22884 12046 22904 12066
rect 22989 12042 23009 12062
rect 23092 12046 23112 12066
rect 23200 12046 23220 12066
rect 30961 12165 30981 12185
rect 31069 12165 31089 12185
rect 31172 12169 31192 12189
rect 31277 12165 31297 12185
rect 31380 12169 31400 12189
rect 31490 12165 31510 12185
rect 31593 12169 31613 12189
rect 31913 12174 31931 12192
rect 23303 12042 23323 12062
rect 23616 12038 23636 12058
rect 22250 12010 22268 12028
rect 23719 12042 23739 12062
rect 23829 12038 23849 12058
rect 23932 12042 23952 12062
rect 24037 12038 24057 12058
rect 24140 12042 24160 12062
rect 24248 12042 24268 12062
rect 24351 12038 24371 12058
rect 20948 11915 20966 11933
rect 31915 12075 31933 12093
rect 32956 12103 32974 12121
rect 39071 12168 39091 12188
rect 39174 12164 39194 12184
rect 39282 12164 39302 12184
rect 39385 12168 39405 12188
rect 39490 12164 39510 12184
rect 39593 12168 39613 12188
rect 39703 12164 39723 12184
rect 39806 12168 39826 12188
rect 41566 12163 41586 12183
rect 33276 12036 33296 12056
rect 33379 12040 33399 12060
rect 33489 12036 33509 12056
rect 33592 12040 33612 12060
rect 33697 12036 33717 12056
rect 33800 12040 33820 12060
rect 33908 12040 33928 12060
rect 41669 12159 41689 12179
rect 41777 12159 41797 12179
rect 41880 12163 41900 12183
rect 41985 12159 42005 12179
rect 42088 12163 42108 12183
rect 42198 12159 42218 12179
rect 42301 12163 42321 12183
rect 42621 12168 42639 12186
rect 34011 12036 34031 12056
rect 34324 12032 34344 12052
rect 32958 12004 32976 12022
rect 34427 12036 34447 12056
rect 34537 12032 34557 12052
rect 34640 12036 34660 12056
rect 34745 12032 34765 12052
rect 34848 12036 34868 12056
rect 34956 12036 34976 12056
rect 35059 12032 35079 12052
rect 31913 11919 31931 11937
rect 42623 12069 42641 12087
rect 42621 11913 42639 11931
rect 10242 11822 10260 11840
rect 20950 11816 20968 11834
rect 31915 11820 31933 11838
rect 42623 11814 42641 11832
rect 575 11716 593 11734
rect 11283 11710 11301 11728
rect 22248 11714 22266 11732
rect 32956 11708 32974 11726
rect 577 11617 595 11635
rect 575 11461 593 11479
rect 11285 11611 11303 11629
rect 8137 11496 8157 11516
rect 8240 11492 8260 11512
rect 8348 11492 8368 11512
rect 8451 11496 8471 11516
rect 8556 11492 8576 11512
rect 8659 11496 8679 11516
rect 8769 11492 8789 11512
rect 10240 11526 10258 11544
rect 8872 11496 8892 11516
rect 9185 11492 9205 11512
rect 577 11362 595 11380
rect 895 11365 915 11385
rect 998 11369 1018 11389
rect 1108 11365 1128 11385
rect 1211 11369 1231 11389
rect 1316 11365 1336 11385
rect 1419 11369 1439 11389
rect 1527 11369 1547 11389
rect 9288 11488 9308 11508
rect 9396 11488 9416 11508
rect 9499 11492 9519 11512
rect 9604 11488 9624 11508
rect 9707 11492 9727 11512
rect 9817 11488 9837 11508
rect 9920 11492 9940 11512
rect 1630 11365 1650 11385
rect 3433 11362 3453 11382
rect 3536 11366 3556 11386
rect 3646 11362 3666 11382
rect 3749 11366 3769 11386
rect 3854 11362 3874 11382
rect 3957 11366 3977 11386
rect 4065 11366 4085 11386
rect 4168 11362 4188 11382
rect 10242 11427 10260 11445
rect 11283 11455 11301 11473
rect 22250 11615 22268 11633
rect 18845 11490 18865 11510
rect 18948 11486 18968 11506
rect 19056 11486 19076 11506
rect 19159 11490 19179 11510
rect 19264 11486 19284 11506
rect 19367 11490 19387 11510
rect 19477 11486 19497 11506
rect 20948 11520 20966 11538
rect 19580 11490 19600 11510
rect 19893 11486 19913 11506
rect 11285 11356 11303 11374
rect 11603 11359 11623 11379
rect 11706 11363 11726 11383
rect 11816 11359 11836 11379
rect 11919 11363 11939 11383
rect 12024 11359 12044 11379
rect 12127 11363 12147 11383
rect 12235 11363 12255 11383
rect 19996 11482 20016 11502
rect 20104 11482 20124 11502
rect 20207 11486 20227 11506
rect 20312 11482 20332 11502
rect 20415 11486 20435 11506
rect 20525 11482 20545 11502
rect 20628 11486 20648 11506
rect 12338 11359 12358 11379
rect 14141 11356 14161 11376
rect 14244 11360 14264 11380
rect 14354 11356 14374 11376
rect 14457 11360 14477 11380
rect 14562 11356 14582 11376
rect 14665 11360 14685 11380
rect 14773 11360 14793 11380
rect 14876 11356 14896 11376
rect 20950 11421 20968 11439
rect 22248 11459 22266 11477
rect 32958 11609 32976 11627
rect 10240 11270 10258 11288
rect 29810 11494 29830 11514
rect 29913 11490 29933 11510
rect 30021 11490 30041 11510
rect 30124 11494 30144 11514
rect 30229 11490 30249 11510
rect 30332 11494 30352 11514
rect 30442 11490 30462 11510
rect 31913 11524 31931 11542
rect 30545 11494 30565 11514
rect 30858 11490 30878 11510
rect 22250 11360 22268 11378
rect 22568 11363 22588 11383
rect 22671 11367 22691 11387
rect 22781 11363 22801 11383
rect 22884 11367 22904 11387
rect 22989 11363 23009 11383
rect 23092 11367 23112 11387
rect 23200 11367 23220 11387
rect 30961 11486 30981 11506
rect 31069 11486 31089 11506
rect 31172 11490 31192 11510
rect 31277 11486 31297 11506
rect 31380 11490 31400 11510
rect 31490 11486 31510 11506
rect 31593 11490 31613 11510
rect 23303 11363 23323 11383
rect 25106 11360 25126 11380
rect 25209 11364 25229 11384
rect 25319 11360 25339 11380
rect 25422 11364 25442 11384
rect 25527 11360 25547 11380
rect 25630 11364 25650 11384
rect 25738 11364 25758 11384
rect 25841 11360 25861 11380
rect 31915 11425 31933 11443
rect 32956 11453 32974 11471
rect 20948 11264 20966 11282
rect 40518 11488 40538 11508
rect 40621 11484 40641 11504
rect 40729 11484 40749 11504
rect 40832 11488 40852 11508
rect 40937 11484 40957 11504
rect 41040 11488 41060 11508
rect 41150 11484 41170 11504
rect 42621 11518 42639 11536
rect 41253 11488 41273 11508
rect 41566 11484 41586 11504
rect 32958 11354 32976 11372
rect 33276 11357 33296 11377
rect 33379 11361 33399 11381
rect 33489 11357 33509 11377
rect 33592 11361 33612 11381
rect 33697 11357 33717 11377
rect 33800 11361 33820 11381
rect 33908 11361 33928 11381
rect 41669 11480 41689 11500
rect 41777 11480 41797 11500
rect 41880 11484 41900 11504
rect 41985 11480 42005 11500
rect 42088 11484 42108 11504
rect 42198 11480 42218 11500
rect 42301 11484 42321 11504
rect 34011 11357 34031 11377
rect 35814 11354 35834 11374
rect 35917 11358 35937 11378
rect 36027 11354 36047 11374
rect 36130 11358 36150 11378
rect 36235 11354 36255 11374
rect 36338 11358 36358 11378
rect 36446 11358 36466 11378
rect 36549 11354 36569 11374
rect 42623 11419 42641 11437
rect 31913 11268 31931 11286
rect 42621 11262 42639 11280
rect 10242 11171 10260 11189
rect 20950 11165 20968 11183
rect 31915 11169 31933 11187
rect 42623 11163 42641 11181
rect 576 10847 594 10865
rect 11284 10841 11302 10859
rect 22249 10845 22267 10863
rect 32957 10839 32975 10857
rect 578 10748 596 10766
rect 11286 10742 11304 10760
rect 576 10591 594 10609
rect 6648 10654 6668 10674
rect 6751 10650 6771 10670
rect 6859 10650 6879 10670
rect 6962 10654 6982 10674
rect 7067 10650 7087 10670
rect 7170 10654 7190 10674
rect 7280 10650 7300 10670
rect 7383 10654 7403 10674
rect 9186 10651 9206 10671
rect 896 10524 916 10544
rect 999 10528 1019 10548
rect 1109 10524 1129 10544
rect 1212 10528 1232 10548
rect 1317 10524 1337 10544
rect 1420 10528 1440 10548
rect 1528 10528 1548 10548
rect 9289 10647 9309 10667
rect 9397 10647 9417 10667
rect 9500 10651 9520 10671
rect 9605 10647 9625 10667
rect 9708 10651 9728 10671
rect 9818 10647 9838 10667
rect 9921 10651 9941 10671
rect 10241 10656 10259 10674
rect 1631 10524 1651 10544
rect 1944 10520 1964 10540
rect 578 10492 596 10510
rect 2047 10524 2067 10544
rect 2157 10520 2177 10540
rect 2260 10524 2280 10544
rect 2365 10520 2385 10540
rect 2468 10524 2488 10544
rect 2576 10524 2596 10544
rect 2679 10520 2699 10540
rect 22251 10746 22269 10764
rect 10243 10557 10261 10575
rect 11284 10585 11302 10603
rect 17356 10648 17376 10668
rect 17459 10644 17479 10664
rect 17567 10644 17587 10664
rect 17670 10648 17690 10668
rect 17775 10644 17795 10664
rect 17878 10648 17898 10668
rect 17988 10644 18008 10664
rect 18091 10648 18111 10668
rect 19894 10645 19914 10665
rect 11604 10518 11624 10538
rect 11707 10522 11727 10542
rect 11817 10518 11837 10538
rect 11920 10522 11940 10542
rect 12025 10518 12045 10538
rect 12128 10522 12148 10542
rect 12236 10522 12256 10542
rect 19997 10641 20017 10661
rect 20105 10641 20125 10661
rect 20208 10645 20228 10665
rect 20313 10641 20333 10661
rect 20416 10645 20436 10665
rect 20526 10641 20546 10661
rect 20629 10645 20649 10665
rect 20949 10650 20967 10668
rect 12339 10518 12359 10538
rect 12652 10514 12672 10534
rect 11286 10486 11304 10504
rect 12755 10518 12775 10538
rect 12865 10514 12885 10534
rect 12968 10518 12988 10538
rect 13073 10514 13093 10534
rect 13176 10518 13196 10538
rect 13284 10518 13304 10538
rect 13387 10514 13407 10534
rect 32959 10740 32977 10758
rect 10241 10401 10259 10419
rect 20951 10551 20969 10569
rect 22249 10589 22267 10607
rect 28321 10652 28341 10672
rect 28424 10648 28444 10668
rect 28532 10648 28552 10668
rect 28635 10652 28655 10672
rect 28740 10648 28760 10668
rect 28843 10652 28863 10672
rect 28953 10648 28973 10668
rect 29056 10652 29076 10672
rect 30859 10649 30879 10669
rect 22569 10522 22589 10542
rect 22672 10526 22692 10546
rect 22782 10522 22802 10542
rect 22885 10526 22905 10546
rect 22990 10522 23010 10542
rect 23093 10526 23113 10546
rect 23201 10526 23221 10546
rect 30962 10645 30982 10665
rect 31070 10645 31090 10665
rect 31173 10649 31193 10669
rect 31278 10645 31298 10665
rect 31381 10649 31401 10669
rect 31491 10645 31511 10665
rect 31594 10649 31614 10669
rect 31914 10654 31932 10672
rect 23304 10522 23324 10542
rect 23617 10518 23637 10538
rect 22251 10490 22269 10508
rect 23720 10522 23740 10542
rect 23830 10518 23850 10538
rect 23933 10522 23953 10542
rect 24038 10518 24058 10538
rect 24141 10522 24161 10542
rect 24249 10522 24269 10542
rect 24352 10518 24372 10538
rect 20949 10395 20967 10413
rect 31916 10555 31934 10573
rect 32957 10583 32975 10601
rect 39029 10646 39049 10666
rect 39132 10642 39152 10662
rect 39240 10642 39260 10662
rect 39343 10646 39363 10666
rect 39448 10642 39468 10662
rect 39551 10646 39571 10666
rect 39661 10642 39681 10662
rect 39764 10646 39784 10666
rect 41567 10643 41587 10663
rect 33277 10516 33297 10536
rect 33380 10520 33400 10540
rect 33490 10516 33510 10536
rect 33593 10520 33613 10540
rect 33698 10516 33718 10536
rect 33801 10520 33821 10540
rect 33909 10520 33929 10540
rect 41670 10639 41690 10659
rect 41778 10639 41798 10659
rect 41881 10643 41901 10663
rect 41986 10639 42006 10659
rect 42089 10643 42109 10663
rect 42199 10639 42219 10659
rect 42302 10643 42322 10663
rect 42622 10648 42640 10666
rect 34012 10516 34032 10536
rect 34325 10512 34345 10532
rect 32959 10484 32977 10502
rect 34428 10516 34448 10536
rect 34538 10512 34558 10532
rect 34641 10516 34661 10536
rect 34746 10512 34766 10532
rect 34849 10516 34869 10536
rect 34957 10516 34977 10536
rect 35060 10512 35080 10532
rect 31914 10399 31932 10417
rect 42624 10549 42642 10567
rect 42622 10393 42640 10411
rect 10243 10302 10261 10320
rect 20951 10296 20969 10314
rect 31916 10300 31934 10318
rect 42624 10294 42642 10312
rect 576 10196 594 10214
rect 11284 10190 11302 10208
rect 22249 10194 22267 10212
rect 32957 10188 32975 10206
rect 578 10097 596 10115
rect 576 9941 594 9959
rect 11286 10091 11304 10109
rect 8138 9976 8158 9996
rect 8241 9972 8261 9992
rect 8349 9972 8369 9992
rect 8452 9976 8472 9996
rect 8557 9972 8577 9992
rect 8660 9976 8680 9996
rect 8770 9972 8790 9992
rect 10241 10006 10259 10024
rect 8873 9976 8893 9996
rect 9186 9972 9206 9992
rect 578 9842 596 9860
rect 896 9845 916 9865
rect 999 9849 1019 9869
rect 1109 9845 1129 9865
rect 1212 9849 1232 9869
rect 1317 9845 1337 9865
rect 1420 9849 1440 9869
rect 1528 9849 1548 9869
rect 9289 9968 9309 9988
rect 9397 9968 9417 9988
rect 9500 9972 9520 9992
rect 9605 9968 9625 9988
rect 9708 9972 9728 9992
rect 9818 9968 9838 9988
rect 9921 9972 9941 9992
rect 1631 9845 1651 9865
rect 3391 9840 3411 9860
rect 3494 9844 3514 9864
rect 3604 9840 3624 9860
rect 3707 9844 3727 9864
rect 3812 9840 3832 9860
rect 3915 9844 3935 9864
rect 4023 9844 4043 9864
rect 4126 9840 4146 9860
rect 10243 9907 10261 9925
rect 11284 9935 11302 9953
rect 22251 10095 22269 10113
rect 18846 9970 18866 9990
rect 18949 9966 18969 9986
rect 19057 9966 19077 9986
rect 19160 9970 19180 9990
rect 19265 9966 19285 9986
rect 19368 9970 19388 9990
rect 19478 9966 19498 9986
rect 20949 10000 20967 10018
rect 19581 9970 19601 9990
rect 19894 9966 19914 9986
rect 11286 9836 11304 9854
rect 11604 9839 11624 9859
rect 11707 9843 11727 9863
rect 11817 9839 11837 9859
rect 11920 9843 11940 9863
rect 12025 9839 12045 9859
rect 12128 9843 12148 9863
rect 12236 9843 12256 9863
rect 19997 9962 20017 9982
rect 20105 9962 20125 9982
rect 20208 9966 20228 9986
rect 20313 9962 20333 9982
rect 20416 9966 20436 9986
rect 20526 9962 20546 9982
rect 20629 9966 20649 9986
rect 12339 9839 12359 9859
rect 14099 9834 14119 9854
rect 14202 9838 14222 9858
rect 14312 9834 14332 9854
rect 14415 9838 14435 9858
rect 14520 9834 14540 9854
rect 14623 9838 14643 9858
rect 14731 9838 14751 9858
rect 14834 9834 14854 9854
rect 20951 9901 20969 9919
rect 22249 9939 22267 9957
rect 32959 10089 32977 10107
rect 10241 9750 10259 9768
rect 29811 9974 29831 9994
rect 29914 9970 29934 9990
rect 30022 9970 30042 9990
rect 30125 9974 30145 9994
rect 30230 9970 30250 9990
rect 30333 9974 30353 9994
rect 30443 9970 30463 9990
rect 31914 10004 31932 10022
rect 30546 9974 30566 9994
rect 30859 9970 30879 9990
rect 22251 9840 22269 9858
rect 22569 9843 22589 9863
rect 22672 9847 22692 9867
rect 22782 9843 22802 9863
rect 22885 9847 22905 9867
rect 22990 9843 23010 9863
rect 23093 9847 23113 9867
rect 23201 9847 23221 9867
rect 30962 9966 30982 9986
rect 31070 9966 31090 9986
rect 31173 9970 31193 9990
rect 31278 9966 31298 9986
rect 31381 9970 31401 9990
rect 31491 9966 31511 9986
rect 31594 9970 31614 9990
rect 23304 9843 23324 9863
rect 25064 9838 25084 9858
rect 25167 9842 25187 9862
rect 25277 9838 25297 9858
rect 25380 9842 25400 9862
rect 25485 9838 25505 9858
rect 25588 9842 25608 9862
rect 25696 9842 25716 9862
rect 25799 9838 25819 9858
rect 31916 9905 31934 9923
rect 32957 9933 32975 9951
rect 20949 9744 20967 9762
rect 40519 9968 40539 9988
rect 40622 9964 40642 9984
rect 40730 9964 40750 9984
rect 40833 9968 40853 9988
rect 40938 9964 40958 9984
rect 41041 9968 41061 9988
rect 41151 9964 41171 9984
rect 42622 9998 42640 10016
rect 41254 9968 41274 9988
rect 41567 9964 41587 9984
rect 32959 9834 32977 9852
rect 33277 9837 33297 9857
rect 33380 9841 33400 9861
rect 33490 9837 33510 9857
rect 33593 9841 33613 9861
rect 33698 9837 33718 9857
rect 33801 9841 33821 9861
rect 33909 9841 33929 9861
rect 41670 9960 41690 9980
rect 41778 9960 41798 9980
rect 41881 9964 41901 9984
rect 41986 9960 42006 9980
rect 42089 9964 42109 9984
rect 42199 9960 42219 9980
rect 42302 9964 42322 9984
rect 34012 9837 34032 9857
rect 35772 9832 35792 9852
rect 35875 9836 35895 9856
rect 35985 9832 36005 9852
rect 36088 9836 36108 9856
rect 36193 9832 36213 9852
rect 36296 9836 36316 9856
rect 36404 9836 36424 9856
rect 36507 9832 36527 9852
rect 42624 9899 42642 9917
rect 31914 9748 31932 9766
rect 42622 9742 42640 9760
rect 10243 9651 10261 9669
rect 20951 9645 20969 9663
rect 31916 9649 31934 9667
rect 42624 9643 42642 9661
rect 576 9400 594 9418
rect 11284 9394 11302 9412
rect 22249 9398 22267 9416
rect 32957 9392 32975 9410
rect 578 9301 596 9319
rect 11286 9295 11304 9313
rect 576 9144 594 9162
rect 6691 9209 6711 9229
rect 6794 9205 6814 9225
rect 6902 9205 6922 9225
rect 7005 9209 7025 9229
rect 7110 9205 7130 9225
rect 7213 9209 7233 9229
rect 7323 9205 7343 9225
rect 7426 9209 7446 9229
rect 9186 9204 9206 9224
rect 896 9077 916 9097
rect 999 9081 1019 9101
rect 1109 9077 1129 9097
rect 1212 9081 1232 9101
rect 1317 9077 1337 9097
rect 1420 9081 1440 9101
rect 1528 9081 1548 9101
rect 9289 9200 9309 9220
rect 9397 9200 9417 9220
rect 9500 9204 9520 9224
rect 9605 9200 9625 9220
rect 9708 9204 9728 9224
rect 9818 9200 9838 9220
rect 9921 9204 9941 9224
rect 10241 9209 10259 9227
rect 1631 9077 1651 9097
rect 1944 9073 1964 9093
rect 578 9045 596 9063
rect 2047 9077 2067 9097
rect 2157 9073 2177 9093
rect 2260 9077 2280 9097
rect 2365 9073 2385 9093
rect 2468 9077 2488 9097
rect 2576 9077 2596 9097
rect 2679 9073 2699 9093
rect 22251 9299 22269 9317
rect 10243 9110 10261 9128
rect 11284 9138 11302 9156
rect 17399 9203 17419 9223
rect 17502 9199 17522 9219
rect 17610 9199 17630 9219
rect 17713 9203 17733 9223
rect 17818 9199 17838 9219
rect 17921 9203 17941 9223
rect 18031 9199 18051 9219
rect 18134 9203 18154 9223
rect 19894 9198 19914 9218
rect 11604 9071 11624 9091
rect 11707 9075 11727 9095
rect 11817 9071 11837 9091
rect 11920 9075 11940 9095
rect 12025 9071 12045 9091
rect 12128 9075 12148 9095
rect 12236 9075 12256 9095
rect 19997 9194 20017 9214
rect 20105 9194 20125 9214
rect 20208 9198 20228 9218
rect 20313 9194 20333 9214
rect 20416 9198 20436 9218
rect 20526 9194 20546 9214
rect 20629 9198 20649 9218
rect 20949 9203 20967 9221
rect 12339 9071 12359 9091
rect 12652 9067 12672 9087
rect 11286 9039 11304 9057
rect 12755 9071 12775 9091
rect 12865 9067 12885 9087
rect 12968 9071 12988 9091
rect 13073 9067 13093 9087
rect 13176 9071 13196 9091
rect 13284 9071 13304 9091
rect 13387 9067 13407 9087
rect 32959 9293 32977 9311
rect 10241 8954 10259 8972
rect 20951 9104 20969 9122
rect 22249 9142 22267 9160
rect 28364 9207 28384 9227
rect 28467 9203 28487 9223
rect 28575 9203 28595 9223
rect 28678 9207 28698 9227
rect 28783 9203 28803 9223
rect 28886 9207 28906 9227
rect 28996 9203 29016 9223
rect 29099 9207 29119 9227
rect 30859 9202 30879 9222
rect 22569 9075 22589 9095
rect 22672 9079 22692 9099
rect 22782 9075 22802 9095
rect 22885 9079 22905 9099
rect 22990 9075 23010 9095
rect 23093 9079 23113 9099
rect 23201 9079 23221 9099
rect 30962 9198 30982 9218
rect 31070 9198 31090 9218
rect 31173 9202 31193 9222
rect 31278 9198 31298 9218
rect 31381 9202 31401 9222
rect 31491 9198 31511 9218
rect 31594 9202 31614 9222
rect 31914 9207 31932 9225
rect 23304 9075 23324 9095
rect 23617 9071 23637 9091
rect 22251 9043 22269 9061
rect 23720 9075 23740 9095
rect 23830 9071 23850 9091
rect 23933 9075 23953 9095
rect 24038 9071 24058 9091
rect 24141 9075 24161 9095
rect 24249 9075 24269 9095
rect 24352 9071 24372 9091
rect 20949 8948 20967 8966
rect 31916 9108 31934 9126
rect 32957 9136 32975 9154
rect 39072 9201 39092 9221
rect 39175 9197 39195 9217
rect 39283 9197 39303 9217
rect 39386 9201 39406 9221
rect 39491 9197 39511 9217
rect 39594 9201 39614 9221
rect 39704 9197 39724 9217
rect 39807 9201 39827 9221
rect 41567 9196 41587 9216
rect 33277 9069 33297 9089
rect 33380 9073 33400 9093
rect 33490 9069 33510 9089
rect 33593 9073 33613 9093
rect 33698 9069 33718 9089
rect 33801 9073 33821 9093
rect 33909 9073 33929 9093
rect 41670 9192 41690 9212
rect 41778 9192 41798 9212
rect 41881 9196 41901 9216
rect 41986 9192 42006 9212
rect 42089 9196 42109 9216
rect 42199 9192 42219 9212
rect 42302 9196 42322 9216
rect 42622 9201 42640 9219
rect 34012 9069 34032 9089
rect 34325 9065 34345 9085
rect 32959 9037 32977 9055
rect 34428 9069 34448 9089
rect 34538 9065 34558 9085
rect 34641 9069 34661 9089
rect 34746 9065 34766 9085
rect 34849 9069 34869 9089
rect 34957 9069 34977 9089
rect 35060 9065 35080 9085
rect 31914 8952 31932 8970
rect 42624 9102 42642 9120
rect 42622 8946 42640 8964
rect 10243 8855 10261 8873
rect 20951 8849 20969 8867
rect 31916 8853 31934 8871
rect 42624 8847 42642 8865
rect 576 8749 594 8767
rect 11284 8743 11302 8761
rect 22249 8747 22267 8765
rect 32957 8741 32975 8759
rect 578 8650 596 8668
rect 576 8494 594 8512
rect 11286 8644 11304 8662
rect 8138 8529 8158 8549
rect 8241 8525 8261 8545
rect 8349 8525 8369 8545
rect 8452 8529 8472 8549
rect 8557 8525 8577 8545
rect 8660 8529 8680 8549
rect 8770 8525 8790 8545
rect 10241 8559 10259 8577
rect 8873 8529 8893 8549
rect 9186 8525 9206 8545
rect 578 8395 596 8413
rect 896 8398 916 8418
rect 999 8402 1019 8422
rect 1109 8398 1129 8418
rect 1212 8402 1232 8422
rect 1317 8398 1337 8418
rect 1420 8402 1440 8422
rect 1528 8402 1548 8422
rect 9289 8521 9309 8541
rect 9397 8521 9417 8541
rect 9500 8525 9520 8545
rect 9605 8521 9625 8541
rect 9708 8525 9728 8545
rect 9818 8521 9838 8541
rect 9921 8525 9941 8545
rect 1631 8398 1651 8418
rect 4499 8389 4519 8409
rect 4602 8393 4622 8413
rect 4712 8389 4732 8409
rect 4815 8393 4835 8413
rect 4920 8389 4940 8409
rect 5023 8393 5043 8413
rect 5131 8393 5151 8413
rect 5234 8389 5254 8409
rect 10243 8460 10261 8478
rect 11284 8488 11302 8506
rect 22251 8648 22269 8666
rect 18846 8523 18866 8543
rect 18949 8519 18969 8539
rect 19057 8519 19077 8539
rect 19160 8523 19180 8543
rect 19265 8519 19285 8539
rect 19368 8523 19388 8543
rect 19478 8519 19498 8539
rect 20949 8553 20967 8571
rect 19581 8523 19601 8543
rect 19894 8519 19914 8539
rect 11286 8389 11304 8407
rect 11604 8392 11624 8412
rect 11707 8396 11727 8416
rect 11817 8392 11837 8412
rect 11920 8396 11940 8416
rect 12025 8392 12045 8412
rect 12128 8396 12148 8416
rect 12236 8396 12256 8416
rect 19997 8515 20017 8535
rect 20105 8515 20125 8535
rect 20208 8519 20228 8539
rect 20313 8515 20333 8535
rect 20416 8519 20436 8539
rect 20526 8515 20546 8535
rect 20629 8519 20649 8539
rect 12339 8392 12359 8412
rect 15207 8383 15227 8403
rect 15310 8387 15330 8407
rect 15420 8383 15440 8403
rect 15523 8387 15543 8407
rect 15628 8383 15648 8403
rect 15731 8387 15751 8407
rect 15839 8387 15859 8407
rect 15942 8383 15962 8403
rect 20951 8454 20969 8472
rect 22249 8492 22267 8510
rect 32959 8642 32977 8660
rect 10241 8303 10259 8321
rect 29811 8527 29831 8547
rect 29914 8523 29934 8543
rect 30022 8523 30042 8543
rect 30125 8527 30145 8547
rect 30230 8523 30250 8543
rect 30333 8527 30353 8547
rect 30443 8523 30463 8543
rect 31914 8557 31932 8575
rect 30546 8527 30566 8547
rect 30859 8523 30879 8543
rect 22251 8393 22269 8411
rect 22569 8396 22589 8416
rect 22672 8400 22692 8420
rect 22782 8396 22802 8416
rect 22885 8400 22905 8420
rect 22990 8396 23010 8416
rect 23093 8400 23113 8420
rect 23201 8400 23221 8420
rect 30962 8519 30982 8539
rect 31070 8519 31090 8539
rect 31173 8523 31193 8543
rect 31278 8519 31298 8539
rect 31381 8523 31401 8543
rect 31491 8519 31511 8539
rect 31594 8523 31614 8543
rect 23304 8396 23324 8416
rect 26172 8387 26192 8407
rect 26275 8391 26295 8411
rect 26385 8387 26405 8407
rect 26488 8391 26508 8411
rect 26593 8387 26613 8407
rect 26696 8391 26716 8411
rect 26804 8391 26824 8411
rect 26907 8387 26927 8407
rect 31916 8458 31934 8476
rect 32957 8486 32975 8504
rect 20949 8297 20967 8315
rect 40519 8521 40539 8541
rect 40622 8517 40642 8537
rect 40730 8517 40750 8537
rect 40833 8521 40853 8541
rect 40938 8517 40958 8537
rect 41041 8521 41061 8541
rect 41151 8517 41171 8537
rect 42622 8551 42640 8569
rect 41254 8521 41274 8541
rect 41567 8517 41587 8537
rect 32959 8387 32977 8405
rect 33277 8390 33297 8410
rect 33380 8394 33400 8414
rect 33490 8390 33510 8410
rect 33593 8394 33613 8414
rect 33698 8390 33718 8410
rect 33801 8394 33821 8414
rect 33909 8394 33929 8414
rect 41670 8513 41690 8533
rect 41778 8513 41798 8533
rect 41881 8517 41901 8537
rect 41986 8513 42006 8533
rect 42089 8517 42109 8537
rect 42199 8513 42219 8533
rect 42302 8517 42322 8537
rect 34012 8390 34032 8410
rect 36880 8381 36900 8401
rect 36983 8385 37003 8405
rect 37093 8381 37113 8401
rect 37196 8385 37216 8405
rect 37301 8381 37321 8401
rect 37404 8385 37424 8405
rect 37512 8385 37532 8405
rect 37615 8381 37635 8401
rect 42624 8452 42642 8470
rect 31914 8301 31932 8319
rect 42622 8295 42640 8313
rect 10243 8204 10261 8222
rect 20951 8198 20969 8216
rect 31916 8202 31934 8220
rect 42624 8196 42642 8214
rect 573 7806 591 7824
rect 11281 7800 11299 7818
rect 22246 7804 22264 7822
rect 32954 7798 32972 7816
rect 575 7707 593 7725
rect 11283 7701 11301 7719
rect 573 7550 591 7568
rect 5580 7619 5600 7639
rect 5683 7615 5703 7635
rect 5791 7615 5811 7635
rect 5894 7619 5914 7639
rect 5999 7615 6019 7635
rect 6102 7619 6122 7639
rect 6212 7615 6232 7635
rect 6315 7619 6335 7639
rect 9183 7610 9203 7630
rect 893 7483 913 7503
rect 996 7487 1016 7507
rect 1106 7483 1126 7503
rect 1209 7487 1229 7507
rect 1314 7483 1334 7503
rect 1417 7487 1437 7507
rect 1525 7487 1545 7507
rect 9286 7606 9306 7626
rect 9394 7606 9414 7626
rect 9497 7610 9517 7630
rect 9602 7606 9622 7626
rect 9705 7610 9725 7630
rect 9815 7606 9835 7626
rect 9918 7610 9938 7630
rect 10238 7615 10256 7633
rect 1628 7483 1648 7503
rect 1941 7479 1961 7499
rect 575 7451 593 7469
rect 2044 7483 2064 7503
rect 2154 7479 2174 7499
rect 2257 7483 2277 7503
rect 2362 7479 2382 7499
rect 2465 7483 2485 7503
rect 2573 7483 2593 7503
rect 2676 7479 2696 7499
rect 22248 7705 22266 7723
rect 10240 7516 10258 7534
rect 11281 7544 11299 7562
rect 16288 7613 16308 7633
rect 16391 7609 16411 7629
rect 16499 7609 16519 7629
rect 16602 7613 16622 7633
rect 16707 7609 16727 7629
rect 16810 7613 16830 7633
rect 16920 7609 16940 7629
rect 17023 7613 17043 7633
rect 19891 7604 19911 7624
rect 11601 7477 11621 7497
rect 11704 7481 11724 7501
rect 11814 7477 11834 7497
rect 11917 7481 11937 7501
rect 12022 7477 12042 7497
rect 12125 7481 12145 7501
rect 12233 7481 12253 7501
rect 19994 7600 20014 7620
rect 20102 7600 20122 7620
rect 20205 7604 20225 7624
rect 20310 7600 20330 7620
rect 20413 7604 20433 7624
rect 20523 7600 20543 7620
rect 20626 7604 20646 7624
rect 20946 7609 20964 7627
rect 12336 7477 12356 7497
rect 12649 7473 12669 7493
rect 11283 7445 11301 7463
rect 12752 7477 12772 7497
rect 12862 7473 12882 7493
rect 12965 7477 12985 7497
rect 13070 7473 13090 7493
rect 13173 7477 13193 7497
rect 13281 7477 13301 7497
rect 13384 7473 13404 7493
rect 32956 7699 32974 7717
rect 10238 7360 10256 7378
rect 20948 7510 20966 7528
rect 22246 7548 22264 7566
rect 27253 7617 27273 7637
rect 27356 7613 27376 7633
rect 27464 7613 27484 7633
rect 27567 7617 27587 7637
rect 27672 7613 27692 7633
rect 27775 7617 27795 7637
rect 27885 7613 27905 7633
rect 27988 7617 28008 7637
rect 30856 7608 30876 7628
rect 22566 7481 22586 7501
rect 22669 7485 22689 7505
rect 22779 7481 22799 7501
rect 22882 7485 22902 7505
rect 22987 7481 23007 7501
rect 23090 7485 23110 7505
rect 23198 7485 23218 7505
rect 30959 7604 30979 7624
rect 31067 7604 31087 7624
rect 31170 7608 31190 7628
rect 31275 7604 31295 7624
rect 31378 7608 31398 7628
rect 31488 7604 31508 7624
rect 31591 7608 31611 7628
rect 31911 7613 31929 7631
rect 23301 7481 23321 7501
rect 23614 7477 23634 7497
rect 22248 7449 22266 7467
rect 23717 7481 23737 7501
rect 23827 7477 23847 7497
rect 23930 7481 23950 7501
rect 24035 7477 24055 7497
rect 24138 7481 24158 7501
rect 24246 7481 24266 7501
rect 24349 7477 24369 7497
rect 20946 7354 20964 7372
rect 31913 7514 31931 7532
rect 32954 7542 32972 7560
rect 37961 7611 37981 7631
rect 38064 7607 38084 7627
rect 38172 7607 38192 7627
rect 38275 7611 38295 7631
rect 38380 7607 38400 7627
rect 38483 7611 38503 7631
rect 38593 7607 38613 7627
rect 38696 7611 38716 7631
rect 41564 7602 41584 7622
rect 33274 7475 33294 7495
rect 33377 7479 33397 7499
rect 33487 7475 33507 7495
rect 33590 7479 33610 7499
rect 33695 7475 33715 7495
rect 33798 7479 33818 7499
rect 33906 7479 33926 7499
rect 41667 7598 41687 7618
rect 41775 7598 41795 7618
rect 41878 7602 41898 7622
rect 41983 7598 42003 7618
rect 42086 7602 42106 7622
rect 42196 7598 42216 7618
rect 42299 7602 42319 7622
rect 42619 7607 42637 7625
rect 34009 7475 34029 7495
rect 34322 7471 34342 7491
rect 32956 7443 32974 7461
rect 34425 7475 34445 7495
rect 34535 7471 34555 7491
rect 34638 7475 34658 7495
rect 34743 7471 34763 7491
rect 34846 7475 34866 7495
rect 34954 7475 34974 7495
rect 35057 7471 35077 7491
rect 31911 7358 31929 7376
rect 42621 7508 42639 7526
rect 42619 7352 42637 7370
rect 10240 7261 10258 7279
rect 20948 7255 20966 7273
rect 31913 7259 31931 7277
rect 42621 7253 42639 7271
rect 573 7155 591 7173
rect 11281 7149 11299 7167
rect 22246 7153 22264 7171
rect 32954 7147 32972 7165
rect 575 7056 593 7074
rect 573 6900 591 6918
rect 11283 7050 11301 7068
rect 8135 6935 8155 6955
rect 8238 6931 8258 6951
rect 8346 6931 8366 6951
rect 8449 6935 8469 6955
rect 8554 6931 8574 6951
rect 8657 6935 8677 6955
rect 8767 6931 8787 6951
rect 10238 6965 10256 6983
rect 8870 6935 8890 6955
rect 9183 6931 9203 6951
rect 575 6801 593 6819
rect 893 6804 913 6824
rect 996 6808 1016 6828
rect 1106 6804 1126 6824
rect 1209 6808 1229 6828
rect 1314 6804 1334 6824
rect 1417 6808 1437 6828
rect 1525 6808 1545 6828
rect 9286 6927 9306 6947
rect 9394 6927 9414 6947
rect 9497 6931 9517 6951
rect 9602 6927 9622 6947
rect 9705 6931 9725 6951
rect 9815 6927 9835 6947
rect 9918 6931 9938 6951
rect 1628 6804 1648 6824
rect 3388 6799 3408 6819
rect 3491 6803 3511 6823
rect 3601 6799 3621 6819
rect 3704 6803 3724 6823
rect 3809 6799 3829 6819
rect 3912 6803 3932 6823
rect 4020 6803 4040 6823
rect 4123 6799 4143 6819
rect 10240 6866 10258 6884
rect 11281 6894 11299 6912
rect 22248 7054 22266 7072
rect 18843 6929 18863 6949
rect 18946 6925 18966 6945
rect 19054 6925 19074 6945
rect 19157 6929 19177 6949
rect 19262 6925 19282 6945
rect 19365 6929 19385 6949
rect 19475 6925 19495 6945
rect 20946 6959 20964 6977
rect 19578 6929 19598 6949
rect 19891 6925 19911 6945
rect 11283 6795 11301 6813
rect 11601 6798 11621 6818
rect 11704 6802 11724 6822
rect 11814 6798 11834 6818
rect 11917 6802 11937 6822
rect 12022 6798 12042 6818
rect 12125 6802 12145 6822
rect 12233 6802 12253 6822
rect 19994 6921 20014 6941
rect 20102 6921 20122 6941
rect 20205 6925 20225 6945
rect 20310 6921 20330 6941
rect 20413 6925 20433 6945
rect 20523 6921 20543 6941
rect 20626 6925 20646 6945
rect 12336 6798 12356 6818
rect 14096 6793 14116 6813
rect 14199 6797 14219 6817
rect 14309 6793 14329 6813
rect 14412 6797 14432 6817
rect 14517 6793 14537 6813
rect 14620 6797 14640 6817
rect 14728 6797 14748 6817
rect 14831 6793 14851 6813
rect 20948 6860 20966 6878
rect 22246 6898 22264 6916
rect 32956 7048 32974 7066
rect 10238 6709 10256 6727
rect 29808 6933 29828 6953
rect 29911 6929 29931 6949
rect 30019 6929 30039 6949
rect 30122 6933 30142 6953
rect 30227 6929 30247 6949
rect 30330 6933 30350 6953
rect 30440 6929 30460 6949
rect 31911 6963 31929 6981
rect 30543 6933 30563 6953
rect 30856 6929 30876 6949
rect 22248 6799 22266 6817
rect 22566 6802 22586 6822
rect 22669 6806 22689 6826
rect 22779 6802 22799 6822
rect 22882 6806 22902 6826
rect 22987 6802 23007 6822
rect 23090 6806 23110 6826
rect 23198 6806 23218 6826
rect 30959 6925 30979 6945
rect 31067 6925 31087 6945
rect 31170 6929 31190 6949
rect 31275 6925 31295 6945
rect 31378 6929 31398 6949
rect 31488 6925 31508 6945
rect 31591 6929 31611 6949
rect 23301 6802 23321 6822
rect 25061 6797 25081 6817
rect 25164 6801 25184 6821
rect 25274 6797 25294 6817
rect 25377 6801 25397 6821
rect 25482 6797 25502 6817
rect 25585 6801 25605 6821
rect 25693 6801 25713 6821
rect 25796 6797 25816 6817
rect 31913 6864 31931 6882
rect 32954 6892 32972 6910
rect 20946 6703 20964 6721
rect 40516 6927 40536 6947
rect 40619 6923 40639 6943
rect 40727 6923 40747 6943
rect 40830 6927 40850 6947
rect 40935 6923 40955 6943
rect 41038 6927 41058 6947
rect 41148 6923 41168 6943
rect 42619 6957 42637 6975
rect 41251 6927 41271 6947
rect 41564 6923 41584 6943
rect 32956 6793 32974 6811
rect 33274 6796 33294 6816
rect 33377 6800 33397 6820
rect 33487 6796 33507 6816
rect 33590 6800 33610 6820
rect 33695 6796 33715 6816
rect 33798 6800 33818 6820
rect 33906 6800 33926 6820
rect 41667 6919 41687 6939
rect 41775 6919 41795 6939
rect 41878 6923 41898 6943
rect 41983 6919 42003 6939
rect 42086 6923 42106 6943
rect 42196 6919 42216 6939
rect 42299 6923 42319 6943
rect 34009 6796 34029 6816
rect 35769 6791 35789 6811
rect 35872 6795 35892 6815
rect 35982 6791 36002 6811
rect 36085 6795 36105 6815
rect 36190 6791 36210 6811
rect 36293 6795 36313 6815
rect 36401 6795 36421 6815
rect 36504 6791 36524 6811
rect 42621 6858 42639 6876
rect 31911 6707 31929 6725
rect 42619 6701 42637 6719
rect 10240 6610 10258 6628
rect 20948 6604 20966 6622
rect 31913 6608 31931 6626
rect 42621 6602 42639 6620
rect 573 6359 591 6377
rect 11281 6353 11299 6371
rect 22246 6357 22264 6375
rect 32954 6351 32972 6369
rect 575 6260 593 6278
rect 11283 6254 11301 6272
rect 573 6103 591 6121
rect 6688 6168 6708 6188
rect 6791 6164 6811 6184
rect 6899 6164 6919 6184
rect 7002 6168 7022 6188
rect 7107 6164 7127 6184
rect 7210 6168 7230 6188
rect 7320 6164 7340 6184
rect 7423 6168 7443 6188
rect 9183 6163 9203 6183
rect 893 6036 913 6056
rect 996 6040 1016 6060
rect 1106 6036 1126 6056
rect 1209 6040 1229 6060
rect 1314 6036 1334 6056
rect 1417 6040 1437 6060
rect 1525 6040 1545 6060
rect 9286 6159 9306 6179
rect 9394 6159 9414 6179
rect 9497 6163 9517 6183
rect 9602 6159 9622 6179
rect 9705 6163 9725 6183
rect 9815 6159 9835 6179
rect 9918 6163 9938 6183
rect 10238 6168 10256 6186
rect 1628 6036 1648 6056
rect 1941 6032 1961 6052
rect 575 6004 593 6022
rect 2044 6036 2064 6056
rect 2154 6032 2174 6052
rect 2257 6036 2277 6056
rect 2362 6032 2382 6052
rect 2465 6036 2485 6056
rect 2573 6036 2593 6056
rect 2676 6032 2696 6052
rect 22248 6258 22266 6276
rect 10240 6069 10258 6087
rect 11281 6097 11299 6115
rect 17396 6162 17416 6182
rect 17499 6158 17519 6178
rect 17607 6158 17627 6178
rect 17710 6162 17730 6182
rect 17815 6158 17835 6178
rect 17918 6162 17938 6182
rect 18028 6158 18048 6178
rect 18131 6162 18151 6182
rect 19891 6157 19911 6177
rect 11601 6030 11621 6050
rect 11704 6034 11724 6054
rect 11814 6030 11834 6050
rect 11917 6034 11937 6054
rect 12022 6030 12042 6050
rect 12125 6034 12145 6054
rect 12233 6034 12253 6054
rect 19994 6153 20014 6173
rect 20102 6153 20122 6173
rect 20205 6157 20225 6177
rect 20310 6153 20330 6173
rect 20413 6157 20433 6177
rect 20523 6153 20543 6173
rect 20626 6157 20646 6177
rect 20946 6162 20964 6180
rect 12336 6030 12356 6050
rect 12649 6026 12669 6046
rect 11283 5998 11301 6016
rect 12752 6030 12772 6050
rect 12862 6026 12882 6046
rect 12965 6030 12985 6050
rect 13070 6026 13090 6046
rect 13173 6030 13193 6050
rect 13281 6030 13301 6050
rect 13384 6026 13404 6046
rect 32956 6252 32974 6270
rect 10238 5913 10256 5931
rect 20948 6063 20966 6081
rect 22246 6101 22264 6119
rect 28361 6166 28381 6186
rect 28464 6162 28484 6182
rect 28572 6162 28592 6182
rect 28675 6166 28695 6186
rect 28780 6162 28800 6182
rect 28883 6166 28903 6186
rect 28993 6162 29013 6182
rect 29096 6166 29116 6186
rect 30856 6161 30876 6181
rect 22566 6034 22586 6054
rect 22669 6038 22689 6058
rect 22779 6034 22799 6054
rect 22882 6038 22902 6058
rect 22987 6034 23007 6054
rect 23090 6038 23110 6058
rect 23198 6038 23218 6058
rect 30959 6157 30979 6177
rect 31067 6157 31087 6177
rect 31170 6161 31190 6181
rect 31275 6157 31295 6177
rect 31378 6161 31398 6181
rect 31488 6157 31508 6177
rect 31591 6161 31611 6181
rect 31911 6166 31929 6184
rect 23301 6034 23321 6054
rect 23614 6030 23634 6050
rect 22248 6002 22266 6020
rect 23717 6034 23737 6054
rect 23827 6030 23847 6050
rect 23930 6034 23950 6054
rect 24035 6030 24055 6050
rect 24138 6034 24158 6054
rect 24246 6034 24266 6054
rect 24349 6030 24369 6050
rect 20946 5907 20964 5925
rect 31913 6067 31931 6085
rect 32954 6095 32972 6113
rect 39069 6160 39089 6180
rect 39172 6156 39192 6176
rect 39280 6156 39300 6176
rect 39383 6160 39403 6180
rect 39488 6156 39508 6176
rect 39591 6160 39611 6180
rect 39701 6156 39721 6176
rect 39804 6160 39824 6180
rect 41564 6155 41584 6175
rect 33274 6028 33294 6048
rect 33377 6032 33397 6052
rect 33487 6028 33507 6048
rect 33590 6032 33610 6052
rect 33695 6028 33715 6048
rect 33798 6032 33818 6052
rect 33906 6032 33926 6052
rect 41667 6151 41687 6171
rect 41775 6151 41795 6171
rect 41878 6155 41898 6175
rect 41983 6151 42003 6171
rect 42086 6155 42106 6175
rect 42196 6151 42216 6171
rect 42299 6155 42319 6175
rect 42619 6160 42637 6178
rect 34009 6028 34029 6048
rect 34322 6024 34342 6044
rect 32956 5996 32974 6014
rect 34425 6028 34445 6048
rect 34535 6024 34555 6044
rect 34638 6028 34658 6048
rect 34743 6024 34763 6044
rect 34846 6028 34866 6048
rect 34954 6028 34974 6048
rect 35057 6024 35077 6044
rect 31911 5911 31929 5929
rect 42621 6061 42639 6079
rect 42619 5905 42637 5923
rect 10240 5814 10258 5832
rect 20948 5808 20966 5826
rect 31913 5812 31931 5830
rect 42621 5806 42639 5824
rect 573 5708 591 5726
rect 11281 5702 11299 5720
rect 22246 5706 22264 5724
rect 32954 5700 32972 5718
rect 575 5609 593 5627
rect 573 5453 591 5471
rect 11283 5603 11301 5621
rect 8135 5488 8155 5508
rect 8238 5484 8258 5504
rect 8346 5484 8366 5504
rect 8449 5488 8469 5508
rect 8554 5484 8574 5504
rect 8657 5488 8677 5508
rect 8767 5484 8787 5504
rect 10238 5518 10256 5536
rect 8870 5488 8890 5508
rect 9183 5484 9203 5504
rect 575 5354 593 5372
rect 893 5357 913 5377
rect 996 5361 1016 5381
rect 1106 5357 1126 5377
rect 1209 5361 1229 5381
rect 1314 5357 1334 5377
rect 1417 5361 1437 5381
rect 1525 5361 1545 5381
rect 9286 5480 9306 5500
rect 9394 5480 9414 5500
rect 9497 5484 9517 5504
rect 9602 5480 9622 5500
rect 9705 5484 9725 5504
rect 9815 5480 9835 5500
rect 9918 5484 9938 5504
rect 1628 5357 1648 5377
rect 3431 5354 3451 5374
rect 3534 5358 3554 5378
rect 3644 5354 3664 5374
rect 3747 5358 3767 5378
rect 3852 5354 3872 5374
rect 3955 5358 3975 5378
rect 4063 5358 4083 5378
rect 4166 5354 4186 5374
rect 10240 5419 10258 5437
rect 11281 5447 11299 5465
rect 22248 5607 22266 5625
rect 18843 5482 18863 5502
rect 18946 5478 18966 5498
rect 19054 5478 19074 5498
rect 19157 5482 19177 5502
rect 19262 5478 19282 5498
rect 19365 5482 19385 5502
rect 19475 5478 19495 5498
rect 20946 5512 20964 5530
rect 19578 5482 19598 5502
rect 19891 5478 19911 5498
rect 11283 5348 11301 5366
rect 11601 5351 11621 5371
rect 11704 5355 11724 5375
rect 11814 5351 11834 5371
rect 11917 5355 11937 5375
rect 12022 5351 12042 5371
rect 12125 5355 12145 5375
rect 12233 5355 12253 5375
rect 19994 5474 20014 5494
rect 20102 5474 20122 5494
rect 20205 5478 20225 5498
rect 20310 5474 20330 5494
rect 20413 5478 20433 5498
rect 20523 5474 20543 5494
rect 20626 5478 20646 5498
rect 12336 5351 12356 5371
rect 14139 5348 14159 5368
rect 14242 5352 14262 5372
rect 14352 5348 14372 5368
rect 14455 5352 14475 5372
rect 14560 5348 14580 5368
rect 14663 5352 14683 5372
rect 14771 5352 14791 5372
rect 14874 5348 14894 5368
rect 20948 5413 20966 5431
rect 22246 5451 22264 5469
rect 32956 5601 32974 5619
rect 10238 5262 10256 5280
rect 29808 5486 29828 5506
rect 29911 5482 29931 5502
rect 30019 5482 30039 5502
rect 30122 5486 30142 5506
rect 30227 5482 30247 5502
rect 30330 5486 30350 5506
rect 30440 5482 30460 5502
rect 31911 5516 31929 5534
rect 30543 5486 30563 5506
rect 30856 5482 30876 5502
rect 22248 5352 22266 5370
rect 22566 5355 22586 5375
rect 22669 5359 22689 5379
rect 22779 5355 22799 5375
rect 22882 5359 22902 5379
rect 22987 5355 23007 5375
rect 23090 5359 23110 5379
rect 23198 5359 23218 5379
rect 30959 5478 30979 5498
rect 31067 5478 31087 5498
rect 31170 5482 31190 5502
rect 31275 5478 31295 5498
rect 31378 5482 31398 5502
rect 31488 5478 31508 5498
rect 31591 5482 31611 5502
rect 23301 5355 23321 5375
rect 25104 5352 25124 5372
rect 25207 5356 25227 5376
rect 25317 5352 25337 5372
rect 25420 5356 25440 5376
rect 25525 5352 25545 5372
rect 25628 5356 25648 5376
rect 25736 5356 25756 5376
rect 25839 5352 25859 5372
rect 31913 5417 31931 5435
rect 32954 5445 32972 5463
rect 20946 5256 20964 5274
rect 40516 5480 40536 5500
rect 40619 5476 40639 5496
rect 40727 5476 40747 5496
rect 40830 5480 40850 5500
rect 40935 5476 40955 5496
rect 41038 5480 41058 5500
rect 41148 5476 41168 5496
rect 42619 5510 42637 5528
rect 41251 5480 41271 5500
rect 41564 5476 41584 5496
rect 32956 5346 32974 5364
rect 33274 5349 33294 5369
rect 33377 5353 33397 5373
rect 33487 5349 33507 5369
rect 33590 5353 33610 5373
rect 33695 5349 33715 5369
rect 33798 5353 33818 5373
rect 33906 5353 33926 5373
rect 41667 5472 41687 5492
rect 41775 5472 41795 5492
rect 41878 5476 41898 5496
rect 41983 5472 42003 5492
rect 42086 5476 42106 5496
rect 42196 5472 42216 5492
rect 42299 5476 42319 5496
rect 34009 5349 34029 5369
rect 35812 5346 35832 5366
rect 35915 5350 35935 5370
rect 36025 5346 36045 5366
rect 36128 5350 36148 5370
rect 36233 5346 36253 5366
rect 36336 5350 36356 5370
rect 36444 5350 36464 5370
rect 36547 5346 36567 5366
rect 42621 5411 42639 5429
rect 31911 5260 31929 5278
rect 42619 5254 42637 5272
rect 10240 5163 10258 5181
rect 20948 5157 20966 5175
rect 31913 5161 31931 5179
rect 42621 5155 42639 5173
rect 574 4839 592 4857
rect 11282 4833 11300 4851
rect 576 4740 594 4758
rect 22247 4837 22265 4855
rect 32955 4831 32973 4849
rect 574 4583 592 4601
rect 11284 4734 11302 4752
rect 6646 4646 6666 4666
rect 6749 4642 6769 4662
rect 6857 4642 6877 4662
rect 6960 4646 6980 4666
rect 7065 4642 7085 4662
rect 7168 4646 7188 4666
rect 7278 4642 7298 4662
rect 7381 4646 7401 4666
rect 9184 4643 9204 4663
rect 894 4516 914 4536
rect 997 4520 1017 4540
rect 1107 4516 1127 4536
rect 1210 4520 1230 4540
rect 1315 4516 1335 4536
rect 1418 4520 1438 4540
rect 1526 4520 1546 4540
rect 9287 4639 9307 4659
rect 9395 4639 9415 4659
rect 9498 4643 9518 4663
rect 9603 4639 9623 4659
rect 9706 4643 9726 4663
rect 9816 4639 9836 4659
rect 9919 4643 9939 4663
rect 10239 4648 10257 4666
rect 1629 4516 1649 4536
rect 1942 4512 1962 4532
rect 576 4484 594 4502
rect 2045 4516 2065 4536
rect 2155 4512 2175 4532
rect 2258 4516 2278 4536
rect 2363 4512 2383 4532
rect 2466 4516 2486 4536
rect 2574 4516 2594 4536
rect 2677 4512 2697 4532
rect 4844 4518 4864 4538
rect 4947 4522 4967 4542
rect 5057 4518 5077 4538
rect 5160 4522 5180 4542
rect 5265 4518 5285 4538
rect 5368 4522 5388 4542
rect 5476 4522 5496 4542
rect 5579 4518 5599 4538
rect 10241 4549 10259 4567
rect 11282 4577 11300 4595
rect 22249 4738 22267 4756
rect 17354 4640 17374 4660
rect 17457 4636 17477 4656
rect 17565 4636 17585 4656
rect 17668 4640 17688 4660
rect 17773 4636 17793 4656
rect 17876 4640 17896 4660
rect 17986 4636 18006 4656
rect 18089 4640 18109 4660
rect 19892 4637 19912 4657
rect 11602 4510 11622 4530
rect 11705 4514 11725 4534
rect 11815 4510 11835 4530
rect 11918 4514 11938 4534
rect 12023 4510 12043 4530
rect 12126 4514 12146 4534
rect 12234 4514 12254 4534
rect 19995 4633 20015 4653
rect 20103 4633 20123 4653
rect 20206 4637 20226 4657
rect 20311 4633 20331 4653
rect 20414 4637 20434 4657
rect 20524 4633 20544 4653
rect 20627 4637 20647 4657
rect 20947 4642 20965 4660
rect 12337 4510 12357 4530
rect 12650 4506 12670 4526
rect 11284 4478 11302 4496
rect 12753 4510 12773 4530
rect 12863 4506 12883 4526
rect 12966 4510 12986 4530
rect 13071 4506 13091 4526
rect 13174 4510 13194 4530
rect 13282 4510 13302 4530
rect 13385 4506 13405 4526
rect 15552 4512 15572 4532
rect 15655 4516 15675 4536
rect 15765 4512 15785 4532
rect 15868 4516 15888 4536
rect 15973 4512 15993 4532
rect 16076 4516 16096 4536
rect 16184 4516 16204 4536
rect 16287 4512 16307 4532
rect 10239 4393 10257 4411
rect 20949 4543 20967 4561
rect 22247 4581 22265 4599
rect 32957 4732 32975 4750
rect 28319 4644 28339 4664
rect 28422 4640 28442 4660
rect 28530 4640 28550 4660
rect 28633 4644 28653 4664
rect 28738 4640 28758 4660
rect 28841 4644 28861 4664
rect 28951 4640 28971 4660
rect 29054 4644 29074 4664
rect 30857 4641 30877 4661
rect 22567 4514 22587 4534
rect 22670 4518 22690 4538
rect 22780 4514 22800 4534
rect 22883 4518 22903 4538
rect 22988 4514 23008 4534
rect 23091 4518 23111 4538
rect 23199 4518 23219 4538
rect 30960 4637 30980 4657
rect 31068 4637 31088 4657
rect 31171 4641 31191 4661
rect 31276 4637 31296 4657
rect 31379 4641 31399 4661
rect 31489 4637 31509 4657
rect 31592 4641 31612 4661
rect 31912 4646 31930 4664
rect 23302 4514 23322 4534
rect 23615 4510 23635 4530
rect 22249 4482 22267 4500
rect 23718 4514 23738 4534
rect 23828 4510 23848 4530
rect 23931 4514 23951 4534
rect 24036 4510 24056 4530
rect 24139 4514 24159 4534
rect 24247 4514 24267 4534
rect 24350 4510 24370 4530
rect 26517 4516 26537 4536
rect 26620 4520 26640 4540
rect 26730 4516 26750 4536
rect 26833 4520 26853 4540
rect 26938 4516 26958 4536
rect 27041 4520 27061 4540
rect 27149 4520 27169 4540
rect 27252 4516 27272 4536
rect 20947 4387 20965 4405
rect 31914 4547 31932 4565
rect 32955 4575 32973 4593
rect 39027 4638 39047 4658
rect 39130 4634 39150 4654
rect 39238 4634 39258 4654
rect 39341 4638 39361 4658
rect 39446 4634 39466 4654
rect 39549 4638 39569 4658
rect 39659 4634 39679 4654
rect 39762 4638 39782 4658
rect 41565 4635 41585 4655
rect 33275 4508 33295 4528
rect 33378 4512 33398 4532
rect 33488 4508 33508 4528
rect 33591 4512 33611 4532
rect 33696 4508 33716 4528
rect 33799 4512 33819 4532
rect 33907 4512 33927 4532
rect 41668 4631 41688 4651
rect 41776 4631 41796 4651
rect 41879 4635 41899 4655
rect 41984 4631 42004 4651
rect 42087 4635 42107 4655
rect 42197 4631 42217 4651
rect 42300 4635 42320 4655
rect 42620 4640 42638 4658
rect 34010 4508 34030 4528
rect 34323 4504 34343 4524
rect 32957 4476 32975 4494
rect 34426 4508 34446 4528
rect 34536 4504 34556 4524
rect 34639 4508 34659 4528
rect 34744 4504 34764 4524
rect 34847 4508 34867 4528
rect 34955 4508 34975 4528
rect 35058 4504 35078 4524
rect 37225 4510 37245 4530
rect 37328 4514 37348 4534
rect 37438 4510 37458 4530
rect 37541 4514 37561 4534
rect 37646 4510 37666 4530
rect 37749 4514 37769 4534
rect 37857 4514 37877 4534
rect 37960 4510 37980 4530
rect 31912 4391 31930 4409
rect 42622 4541 42640 4559
rect 42620 4385 42638 4403
rect 10241 4294 10259 4312
rect 20949 4288 20967 4306
rect 31914 4292 31932 4310
rect 42622 4286 42640 4304
rect 574 4188 592 4206
rect 11282 4182 11300 4200
rect 22247 4186 22265 4204
rect 32955 4180 32973 4198
rect 576 4089 594 4107
rect 574 3933 592 3951
rect 11284 4083 11302 4101
rect 8136 3968 8156 3988
rect 8239 3964 8259 3984
rect 8347 3964 8367 3984
rect 8450 3968 8470 3988
rect 8555 3964 8575 3984
rect 8658 3968 8678 3988
rect 8768 3964 8788 3984
rect 10239 3998 10257 4016
rect 8871 3968 8891 3988
rect 9184 3964 9204 3984
rect 576 3834 594 3852
rect 894 3837 914 3857
rect 997 3841 1017 3861
rect 1107 3837 1127 3857
rect 1210 3841 1230 3861
rect 1315 3837 1335 3857
rect 1418 3841 1438 3861
rect 1526 3841 1546 3861
rect 9287 3960 9307 3980
rect 9395 3960 9415 3980
rect 9498 3964 9518 3984
rect 9603 3960 9623 3980
rect 9706 3964 9726 3984
rect 9816 3960 9836 3980
rect 9919 3964 9939 3984
rect 1629 3837 1649 3857
rect 3389 3832 3409 3852
rect 3492 3836 3512 3856
rect 3602 3832 3622 3852
rect 3705 3836 3725 3856
rect 3810 3832 3830 3852
rect 3913 3836 3933 3856
rect 4021 3836 4041 3856
rect 4124 3832 4144 3852
rect 10241 3899 10259 3917
rect 11282 3927 11300 3945
rect 22249 4087 22267 4105
rect 18844 3962 18864 3982
rect 18947 3958 18967 3978
rect 19055 3958 19075 3978
rect 19158 3962 19178 3982
rect 19263 3958 19283 3978
rect 19366 3962 19386 3982
rect 19476 3958 19496 3978
rect 20947 3992 20965 4010
rect 19579 3962 19599 3982
rect 19892 3958 19912 3978
rect 11284 3828 11302 3846
rect 11602 3831 11622 3851
rect 11705 3835 11725 3855
rect 11815 3831 11835 3851
rect 11918 3835 11938 3855
rect 12023 3831 12043 3851
rect 12126 3835 12146 3855
rect 12234 3835 12254 3855
rect 19995 3954 20015 3974
rect 20103 3954 20123 3974
rect 20206 3958 20226 3978
rect 20311 3954 20331 3974
rect 20414 3958 20434 3978
rect 20524 3954 20544 3974
rect 20627 3958 20647 3978
rect 12337 3831 12357 3851
rect 14097 3826 14117 3846
rect 14200 3830 14220 3850
rect 14310 3826 14330 3846
rect 14413 3830 14433 3850
rect 14518 3826 14538 3846
rect 14621 3830 14641 3850
rect 14729 3830 14749 3850
rect 14832 3826 14852 3846
rect 20949 3893 20967 3911
rect 22247 3931 22265 3949
rect 32957 4081 32975 4099
rect 10239 3742 10257 3760
rect 29809 3966 29829 3986
rect 29912 3962 29932 3982
rect 30020 3962 30040 3982
rect 30123 3966 30143 3986
rect 30228 3962 30248 3982
rect 30331 3966 30351 3986
rect 30441 3962 30461 3982
rect 31912 3996 31930 4014
rect 30544 3966 30564 3986
rect 30857 3962 30877 3982
rect 22249 3832 22267 3850
rect 22567 3835 22587 3855
rect 22670 3839 22690 3859
rect 22780 3835 22800 3855
rect 22883 3839 22903 3859
rect 22988 3835 23008 3855
rect 23091 3839 23111 3859
rect 23199 3839 23219 3859
rect 30960 3958 30980 3978
rect 31068 3958 31088 3978
rect 31171 3962 31191 3982
rect 31276 3958 31296 3978
rect 31379 3962 31399 3982
rect 31489 3958 31509 3978
rect 31592 3962 31612 3982
rect 23302 3835 23322 3855
rect 25062 3830 25082 3850
rect 25165 3834 25185 3854
rect 25275 3830 25295 3850
rect 25378 3834 25398 3854
rect 25483 3830 25503 3850
rect 25586 3834 25606 3854
rect 25694 3834 25714 3854
rect 25797 3830 25817 3850
rect 31914 3897 31932 3915
rect 32955 3925 32973 3943
rect 20947 3736 20965 3754
rect 40517 3960 40537 3980
rect 40620 3956 40640 3976
rect 40728 3956 40748 3976
rect 40831 3960 40851 3980
rect 40936 3956 40956 3976
rect 41039 3960 41059 3980
rect 41149 3956 41169 3976
rect 42620 3990 42638 4008
rect 41252 3960 41272 3980
rect 41565 3956 41585 3976
rect 32957 3826 32975 3844
rect 33275 3829 33295 3849
rect 33378 3833 33398 3853
rect 33488 3829 33508 3849
rect 33591 3833 33611 3853
rect 33696 3829 33716 3849
rect 33799 3833 33819 3853
rect 33907 3833 33927 3853
rect 41668 3952 41688 3972
rect 41776 3952 41796 3972
rect 41879 3956 41899 3976
rect 41984 3952 42004 3972
rect 42087 3956 42107 3976
rect 42197 3952 42217 3972
rect 42300 3956 42320 3976
rect 34010 3829 34030 3849
rect 35770 3824 35790 3844
rect 35873 3828 35893 3848
rect 35983 3824 36003 3844
rect 36086 3828 36106 3848
rect 36191 3824 36211 3844
rect 36294 3828 36314 3848
rect 36402 3828 36422 3848
rect 36505 3824 36525 3844
rect 42622 3891 42640 3909
rect 31912 3740 31930 3758
rect 42620 3734 42638 3752
rect 10241 3643 10259 3661
rect 20949 3637 20967 3655
rect 31914 3641 31932 3659
rect 42622 3635 42640 3653
rect 574 3392 592 3410
rect 11282 3386 11300 3404
rect 22247 3390 22265 3408
rect 32955 3384 32973 3402
rect 576 3293 594 3311
rect 11284 3287 11302 3305
rect 574 3136 592 3154
rect 6689 3201 6709 3221
rect 6792 3197 6812 3217
rect 6900 3197 6920 3217
rect 7003 3201 7023 3221
rect 7108 3197 7128 3217
rect 7211 3201 7231 3221
rect 7321 3197 7341 3217
rect 7424 3201 7444 3221
rect 9184 3196 9204 3216
rect 894 3069 914 3089
rect 997 3073 1017 3093
rect 1107 3069 1127 3089
rect 1210 3073 1230 3093
rect 1315 3069 1335 3089
rect 1418 3073 1438 3093
rect 1526 3073 1546 3093
rect 9287 3192 9307 3212
rect 9395 3192 9415 3212
rect 9498 3196 9518 3216
rect 9603 3192 9623 3212
rect 9706 3196 9726 3216
rect 9816 3192 9836 3212
rect 9919 3196 9939 3216
rect 10239 3201 10257 3219
rect 1629 3069 1649 3089
rect 1942 3065 1962 3085
rect 576 3037 594 3055
rect 2045 3069 2065 3089
rect 2155 3065 2175 3085
rect 2258 3069 2278 3089
rect 2363 3065 2383 3085
rect 2466 3069 2486 3089
rect 2574 3069 2594 3089
rect 2677 3065 2697 3085
rect 22249 3291 22267 3309
rect 10241 3102 10259 3120
rect 11282 3130 11300 3148
rect 17397 3195 17417 3215
rect 17500 3191 17520 3211
rect 17608 3191 17628 3211
rect 17711 3195 17731 3215
rect 17816 3191 17836 3211
rect 17919 3195 17939 3215
rect 18029 3191 18049 3211
rect 18132 3195 18152 3215
rect 19892 3190 19912 3210
rect 11602 3063 11622 3083
rect 11705 3067 11725 3087
rect 11815 3063 11835 3083
rect 11918 3067 11938 3087
rect 12023 3063 12043 3083
rect 12126 3067 12146 3087
rect 12234 3067 12254 3087
rect 19995 3186 20015 3206
rect 20103 3186 20123 3206
rect 20206 3190 20226 3210
rect 20311 3186 20331 3206
rect 20414 3190 20434 3210
rect 20524 3186 20544 3206
rect 20627 3190 20647 3210
rect 20947 3195 20965 3213
rect 12337 3063 12357 3083
rect 12650 3059 12670 3079
rect 11284 3031 11302 3049
rect 12753 3063 12773 3083
rect 12863 3059 12883 3079
rect 12966 3063 12986 3083
rect 13071 3059 13091 3079
rect 13174 3063 13194 3083
rect 13282 3063 13302 3083
rect 13385 3059 13405 3079
rect 32957 3285 32975 3303
rect 10239 2946 10257 2964
rect 20949 3096 20967 3114
rect 22247 3134 22265 3152
rect 28362 3199 28382 3219
rect 28465 3195 28485 3215
rect 28573 3195 28593 3215
rect 28676 3199 28696 3219
rect 28781 3195 28801 3215
rect 28884 3199 28904 3219
rect 28994 3195 29014 3215
rect 29097 3199 29117 3219
rect 30857 3194 30877 3214
rect 22567 3067 22587 3087
rect 22670 3071 22690 3091
rect 22780 3067 22800 3087
rect 22883 3071 22903 3091
rect 22988 3067 23008 3087
rect 23091 3071 23111 3091
rect 23199 3071 23219 3091
rect 30960 3190 30980 3210
rect 31068 3190 31088 3210
rect 31171 3194 31191 3214
rect 31276 3190 31296 3210
rect 31379 3194 31399 3214
rect 31489 3190 31509 3210
rect 31592 3194 31612 3214
rect 31912 3199 31930 3217
rect 23302 3067 23322 3087
rect 23615 3063 23635 3083
rect 22249 3035 22267 3053
rect 23718 3067 23738 3087
rect 23828 3063 23848 3083
rect 23931 3067 23951 3087
rect 24036 3063 24056 3083
rect 24139 3067 24159 3087
rect 24247 3067 24267 3087
rect 24350 3063 24370 3083
rect 20947 2940 20965 2958
rect 31914 3100 31932 3118
rect 32955 3128 32973 3146
rect 39070 3193 39090 3213
rect 39173 3189 39193 3209
rect 39281 3189 39301 3209
rect 39384 3193 39404 3213
rect 39489 3189 39509 3209
rect 39592 3193 39612 3213
rect 39702 3189 39722 3209
rect 39805 3193 39825 3213
rect 41565 3188 41585 3208
rect 33275 3061 33295 3081
rect 33378 3065 33398 3085
rect 33488 3061 33508 3081
rect 33591 3065 33611 3085
rect 33696 3061 33716 3081
rect 33799 3065 33819 3085
rect 33907 3065 33927 3085
rect 41668 3184 41688 3204
rect 41776 3184 41796 3204
rect 41879 3188 41899 3208
rect 41984 3184 42004 3204
rect 42087 3188 42107 3208
rect 42197 3184 42217 3204
rect 42300 3188 42320 3208
rect 42620 3193 42638 3211
rect 34010 3061 34030 3081
rect 34323 3057 34343 3077
rect 32957 3029 32975 3047
rect 34426 3061 34446 3081
rect 34536 3057 34556 3077
rect 34639 3061 34659 3081
rect 34744 3057 34764 3077
rect 34847 3061 34867 3081
rect 34955 3061 34975 3081
rect 35058 3057 35078 3077
rect 31912 2944 31930 2962
rect 42622 3094 42640 3112
rect 42620 2938 42638 2956
rect 10241 2847 10259 2865
rect 20949 2841 20967 2859
rect 31914 2845 31932 2863
rect 42622 2839 42640 2857
rect 574 2741 592 2759
rect 11282 2735 11300 2753
rect 22247 2739 22265 2757
rect 32955 2733 32973 2751
rect 576 2642 594 2660
rect 574 2486 592 2504
rect 11284 2636 11302 2654
rect 8136 2521 8156 2541
rect 8239 2517 8259 2537
rect 8347 2517 8367 2537
rect 8450 2521 8470 2541
rect 8555 2517 8575 2537
rect 8658 2521 8678 2541
rect 8768 2517 8788 2537
rect 10239 2551 10257 2569
rect 8871 2521 8891 2541
rect 9184 2517 9204 2537
rect 9287 2513 9307 2533
rect 9395 2513 9415 2533
rect 9498 2517 9518 2537
rect 9603 2513 9623 2533
rect 9706 2517 9726 2537
rect 9816 2513 9836 2533
rect 9919 2517 9939 2537
rect 576 2387 594 2405
rect 894 2390 914 2410
rect 997 2394 1017 2414
rect 1107 2390 1127 2410
rect 1210 2394 1230 2414
rect 1315 2390 1335 2410
rect 1418 2394 1438 2414
rect 1526 2394 1546 2414
rect 1629 2390 1649 2410
rect 10241 2452 10259 2470
rect 11282 2480 11300 2498
rect 22249 2640 22267 2658
rect 18844 2515 18864 2535
rect 18947 2511 18967 2531
rect 19055 2511 19075 2531
rect 19158 2515 19178 2535
rect 19263 2511 19283 2531
rect 19366 2515 19386 2535
rect 19476 2511 19496 2531
rect 20947 2545 20965 2563
rect 19579 2515 19599 2535
rect 19892 2511 19912 2531
rect 19995 2507 20015 2527
rect 20103 2507 20123 2527
rect 20206 2511 20226 2531
rect 20311 2507 20331 2527
rect 20414 2511 20434 2531
rect 20524 2507 20544 2527
rect 20627 2511 20647 2531
rect 11284 2381 11302 2399
rect 11602 2384 11622 2404
rect 11705 2388 11725 2408
rect 11815 2384 11835 2404
rect 11918 2388 11938 2408
rect 12023 2384 12043 2404
rect 12126 2388 12146 2408
rect 12234 2388 12254 2408
rect 12337 2384 12357 2404
rect 20949 2446 20967 2464
rect 22247 2484 22265 2502
rect 32957 2634 32975 2652
rect 29809 2519 29829 2539
rect 29912 2515 29932 2535
rect 30020 2515 30040 2535
rect 30123 2519 30143 2539
rect 30228 2515 30248 2535
rect 30331 2519 30351 2539
rect 30441 2515 30461 2535
rect 31912 2549 31930 2567
rect 30544 2519 30564 2539
rect 30857 2515 30877 2535
rect 10239 2295 10257 2313
rect 30960 2511 30980 2531
rect 31068 2511 31088 2531
rect 31171 2515 31191 2535
rect 31276 2511 31296 2531
rect 31379 2515 31399 2535
rect 31489 2511 31509 2531
rect 31592 2515 31612 2535
rect 22249 2385 22267 2403
rect 22567 2388 22587 2408
rect 22670 2392 22690 2412
rect 22780 2388 22800 2408
rect 22883 2392 22903 2412
rect 22988 2388 23008 2408
rect 23091 2392 23111 2412
rect 23199 2392 23219 2412
rect 23302 2388 23322 2408
rect 31914 2450 31932 2468
rect 32955 2478 32973 2496
rect 40517 2513 40537 2533
rect 40620 2509 40640 2529
rect 40728 2509 40748 2529
rect 40831 2513 40851 2533
rect 40936 2509 40956 2529
rect 41039 2513 41059 2533
rect 41149 2509 41169 2529
rect 42620 2543 42638 2561
rect 41252 2513 41272 2533
rect 41565 2509 41585 2529
rect 20947 2289 20965 2307
rect 41668 2505 41688 2525
rect 41776 2505 41796 2525
rect 41879 2509 41899 2529
rect 41984 2505 42004 2525
rect 42087 2509 42107 2529
rect 42197 2505 42217 2525
rect 42300 2509 42320 2529
rect 32957 2379 32975 2397
rect 33275 2382 33295 2402
rect 33378 2386 33398 2406
rect 33488 2382 33508 2402
rect 33591 2386 33611 2406
rect 33696 2382 33716 2402
rect 33799 2386 33819 2406
rect 33907 2386 33927 2406
rect 34010 2382 34030 2402
rect 42622 2444 42640 2462
rect 31912 2293 31930 2311
rect 42620 2287 42638 2305
rect 10241 2196 10259 2214
rect 20949 2190 20967 2208
rect 31914 2194 31932 2212
rect 42622 2188 42640 2206
rect 10605 231 10625 251
rect 10708 235 10728 255
rect 10818 231 10838 251
rect 10921 235 10941 255
rect 11026 231 11046 251
rect 11129 235 11149 255
rect 11237 235 11257 255
rect 11340 231 11360 251
rect 21242 218 21262 238
rect 21345 222 21365 242
rect 21455 218 21475 238
rect 21558 222 21578 242
rect 21663 218 21683 238
rect 21766 222 21786 242
rect 21874 222 21894 242
rect 21977 218 21997 238
rect 32278 229 32298 249
rect 32381 233 32401 253
rect 32491 229 32511 249
rect 32594 233 32614 253
rect 32699 229 32719 249
rect 32802 233 32822 253
rect 32910 233 32930 253
rect 33013 229 33033 249
<< pdiffc >>
rect 901 13640 921 13660
rect 997 13640 1017 13660
rect 1114 13640 1134 13660
rect 1210 13640 1230 13660
rect 1322 13640 1342 13660
rect 1418 13640 1438 13660
rect 1528 13640 1548 13660
rect 1624 13640 1644 13660
rect 1949 13636 1969 13656
rect 2045 13636 2065 13656
rect 2162 13636 2182 13656
rect 2258 13636 2278 13656
rect 2370 13636 2390 13656
rect 2466 13636 2486 13656
rect 2576 13636 2596 13656
rect 2672 13636 2692 13656
rect 11609 13634 11629 13654
rect 11705 13634 11725 13654
rect 11822 13634 11842 13654
rect 11918 13634 11938 13654
rect 12030 13634 12050 13654
rect 12126 13634 12146 13654
rect 12236 13634 12256 13654
rect 12332 13634 12352 13654
rect 12657 13630 12677 13650
rect 9191 13469 9211 13489
rect 9287 13469 9307 13489
rect 9397 13469 9417 13489
rect 9493 13469 9513 13489
rect 9605 13469 9625 13489
rect 9701 13469 9721 13489
rect 9818 13469 9838 13489
rect 12753 13630 12773 13650
rect 12870 13630 12890 13650
rect 12966 13630 12986 13650
rect 13078 13630 13098 13650
rect 13174 13630 13194 13650
rect 13284 13630 13304 13650
rect 13380 13630 13400 13650
rect 9914 13469 9934 13489
rect 22574 13638 22594 13658
rect 22670 13638 22690 13658
rect 22787 13638 22807 13658
rect 22883 13638 22903 13658
rect 22995 13638 23015 13658
rect 23091 13638 23111 13658
rect 23201 13638 23221 13658
rect 23297 13638 23317 13658
rect 23622 13634 23642 13654
rect 19899 13463 19919 13483
rect 19995 13463 20015 13483
rect 20105 13463 20125 13483
rect 20201 13463 20221 13483
rect 20313 13463 20333 13483
rect 20409 13463 20429 13483
rect 20526 13463 20546 13483
rect 23718 13634 23738 13654
rect 23835 13634 23855 13654
rect 23931 13634 23951 13654
rect 24043 13634 24063 13654
rect 24139 13634 24159 13654
rect 24249 13634 24269 13654
rect 24345 13634 24365 13654
rect 20622 13463 20642 13483
rect 33282 13632 33302 13652
rect 33378 13632 33398 13652
rect 33495 13632 33515 13652
rect 33591 13632 33611 13652
rect 33703 13632 33723 13652
rect 33799 13632 33819 13652
rect 33909 13632 33929 13652
rect 34005 13632 34025 13652
rect 34330 13628 34350 13648
rect 30864 13467 30884 13487
rect 30960 13467 30980 13487
rect 31070 13467 31090 13487
rect 31166 13467 31186 13487
rect 31278 13467 31298 13487
rect 31374 13467 31394 13487
rect 31491 13467 31511 13487
rect 34426 13628 34446 13648
rect 34543 13628 34563 13648
rect 34639 13628 34659 13648
rect 34751 13628 34771 13648
rect 34847 13628 34867 13648
rect 34957 13628 34977 13648
rect 35053 13628 35073 13648
rect 31587 13467 31607 13487
rect 41572 13461 41592 13481
rect 41668 13461 41688 13481
rect 41778 13461 41798 13481
rect 41874 13461 41894 13481
rect 41986 13461 42006 13481
rect 42082 13461 42102 13481
rect 42199 13461 42219 13481
rect 42295 13461 42315 13481
rect 901 12961 921 12981
rect 997 12961 1017 12981
rect 1114 12961 1134 12981
rect 1210 12961 1230 12981
rect 1322 12961 1342 12981
rect 1418 12961 1438 12981
rect 1528 12961 1548 12981
rect 1624 12961 1644 12981
rect 3396 12956 3416 12976
rect 3492 12956 3512 12976
rect 3609 12956 3629 12976
rect 3705 12956 3725 12976
rect 3817 12956 3837 12976
rect 3913 12956 3933 12976
rect 4023 12956 4043 12976
rect 4119 12956 4139 12976
rect 11609 12955 11629 12975
rect 8143 12794 8163 12814
rect 8239 12794 8259 12814
rect 8349 12794 8369 12814
rect 8445 12794 8465 12814
rect 8557 12794 8577 12814
rect 8653 12794 8673 12814
rect 8770 12794 8790 12814
rect 11705 12955 11725 12975
rect 11822 12955 11842 12975
rect 11918 12955 11938 12975
rect 12030 12955 12050 12975
rect 12126 12955 12146 12975
rect 12236 12955 12256 12975
rect 12332 12955 12352 12975
rect 14104 12950 14124 12970
rect 8866 12794 8886 12814
rect 9191 12790 9211 12810
rect 9287 12790 9307 12810
rect 9397 12790 9417 12810
rect 9493 12790 9513 12810
rect 9605 12790 9625 12810
rect 9701 12790 9721 12810
rect 9818 12790 9838 12810
rect 9914 12790 9934 12810
rect 14200 12950 14220 12970
rect 14317 12950 14337 12970
rect 14413 12950 14433 12970
rect 14525 12950 14545 12970
rect 14621 12950 14641 12970
rect 14731 12950 14751 12970
rect 14827 12950 14847 12970
rect 22574 12959 22594 12979
rect 18851 12788 18871 12808
rect 18947 12788 18967 12808
rect 19057 12788 19077 12808
rect 19153 12788 19173 12808
rect 19265 12788 19285 12808
rect 19361 12788 19381 12808
rect 19478 12788 19498 12808
rect 22670 12959 22690 12979
rect 22787 12959 22807 12979
rect 22883 12959 22903 12979
rect 22995 12959 23015 12979
rect 23091 12959 23111 12979
rect 23201 12959 23221 12979
rect 23297 12959 23317 12979
rect 25069 12954 25089 12974
rect 19574 12788 19594 12808
rect 19899 12784 19919 12804
rect 19995 12784 20015 12804
rect 20105 12784 20125 12804
rect 20201 12784 20221 12804
rect 20313 12784 20333 12804
rect 20409 12784 20429 12804
rect 20526 12784 20546 12804
rect 20622 12784 20642 12804
rect 25165 12954 25185 12974
rect 25282 12954 25302 12974
rect 25378 12954 25398 12974
rect 25490 12954 25510 12974
rect 25586 12954 25606 12974
rect 25696 12954 25716 12974
rect 25792 12954 25812 12974
rect 33282 12953 33302 12973
rect 29816 12792 29836 12812
rect 29912 12792 29932 12812
rect 30022 12792 30042 12812
rect 30118 12792 30138 12812
rect 30230 12792 30250 12812
rect 30326 12792 30346 12812
rect 30443 12792 30463 12812
rect 33378 12953 33398 12973
rect 33495 12953 33515 12973
rect 33591 12953 33611 12973
rect 33703 12953 33723 12973
rect 33799 12953 33819 12973
rect 33909 12953 33929 12973
rect 34005 12953 34025 12973
rect 35777 12948 35797 12968
rect 30539 12792 30559 12812
rect 30864 12788 30884 12808
rect 30960 12788 30980 12808
rect 31070 12788 31090 12808
rect 31166 12788 31186 12808
rect 31278 12788 31298 12808
rect 31374 12788 31394 12808
rect 31491 12788 31511 12808
rect 31587 12788 31607 12808
rect 35873 12948 35893 12968
rect 35990 12948 36010 12968
rect 36086 12948 36106 12968
rect 36198 12948 36218 12968
rect 36294 12948 36314 12968
rect 36404 12948 36424 12968
rect 36500 12948 36520 12968
rect 40524 12786 40544 12806
rect 40620 12786 40640 12806
rect 40730 12786 40750 12806
rect 40826 12786 40846 12806
rect 40938 12786 40958 12806
rect 41034 12786 41054 12806
rect 41151 12786 41171 12806
rect 41247 12786 41267 12806
rect 41572 12782 41592 12802
rect 41668 12782 41688 12802
rect 41778 12782 41798 12802
rect 41874 12782 41894 12802
rect 41986 12782 42006 12802
rect 42082 12782 42102 12802
rect 42199 12782 42219 12802
rect 42295 12782 42315 12802
rect 901 12193 921 12213
rect 997 12193 1017 12213
rect 1114 12193 1134 12213
rect 1210 12193 1230 12213
rect 1322 12193 1342 12213
rect 1418 12193 1438 12213
rect 1528 12193 1548 12213
rect 1624 12193 1644 12213
rect 1949 12189 1969 12209
rect 2045 12189 2065 12209
rect 2162 12189 2182 12209
rect 2258 12189 2278 12209
rect 2370 12189 2390 12209
rect 2466 12189 2486 12209
rect 2576 12189 2596 12209
rect 2672 12189 2692 12209
rect 6696 12027 6716 12047
rect 6792 12027 6812 12047
rect 6902 12027 6922 12047
rect 6998 12027 7018 12047
rect 7110 12027 7130 12047
rect 7206 12027 7226 12047
rect 7323 12027 7343 12047
rect 11609 12187 11629 12207
rect 11705 12187 11725 12207
rect 11822 12187 11842 12207
rect 11918 12187 11938 12207
rect 12030 12187 12050 12207
rect 12126 12187 12146 12207
rect 12236 12187 12256 12207
rect 12332 12187 12352 12207
rect 12657 12183 12677 12203
rect 7419 12027 7439 12047
rect 9191 12022 9211 12042
rect 9287 12022 9307 12042
rect 9397 12022 9417 12042
rect 9493 12022 9513 12042
rect 9605 12022 9625 12042
rect 9701 12022 9721 12042
rect 9818 12022 9838 12042
rect 12753 12183 12773 12203
rect 12870 12183 12890 12203
rect 12966 12183 12986 12203
rect 13078 12183 13098 12203
rect 13174 12183 13194 12203
rect 13284 12183 13304 12203
rect 13380 12183 13400 12203
rect 9914 12022 9934 12042
rect 17404 12021 17424 12041
rect 17500 12021 17520 12041
rect 17610 12021 17630 12041
rect 17706 12021 17726 12041
rect 17818 12021 17838 12041
rect 17914 12021 17934 12041
rect 18031 12021 18051 12041
rect 22574 12191 22594 12211
rect 22670 12191 22690 12211
rect 22787 12191 22807 12211
rect 22883 12191 22903 12211
rect 22995 12191 23015 12211
rect 23091 12191 23111 12211
rect 23201 12191 23221 12211
rect 23297 12191 23317 12211
rect 23622 12187 23642 12207
rect 18127 12021 18147 12041
rect 19899 12016 19919 12036
rect 19995 12016 20015 12036
rect 20105 12016 20125 12036
rect 20201 12016 20221 12036
rect 20313 12016 20333 12036
rect 20409 12016 20429 12036
rect 20526 12016 20546 12036
rect 23718 12187 23738 12207
rect 23835 12187 23855 12207
rect 23931 12187 23951 12207
rect 24043 12187 24063 12207
rect 24139 12187 24159 12207
rect 24249 12187 24269 12207
rect 24345 12187 24365 12207
rect 20622 12016 20642 12036
rect 28369 12025 28389 12045
rect 28465 12025 28485 12045
rect 28575 12025 28595 12045
rect 28671 12025 28691 12045
rect 28783 12025 28803 12045
rect 28879 12025 28899 12045
rect 28996 12025 29016 12045
rect 33282 12185 33302 12205
rect 33378 12185 33398 12205
rect 33495 12185 33515 12205
rect 33591 12185 33611 12205
rect 33703 12185 33723 12205
rect 33799 12185 33819 12205
rect 33909 12185 33929 12205
rect 34005 12185 34025 12205
rect 34330 12181 34350 12201
rect 29092 12025 29112 12045
rect 30864 12020 30884 12040
rect 30960 12020 30980 12040
rect 31070 12020 31090 12040
rect 31166 12020 31186 12040
rect 31278 12020 31298 12040
rect 31374 12020 31394 12040
rect 31491 12020 31511 12040
rect 34426 12181 34446 12201
rect 34543 12181 34563 12201
rect 34639 12181 34659 12201
rect 34751 12181 34771 12201
rect 34847 12181 34867 12201
rect 34957 12181 34977 12201
rect 35053 12181 35073 12201
rect 31587 12020 31607 12040
rect 39077 12019 39097 12039
rect 39173 12019 39193 12039
rect 39283 12019 39303 12039
rect 39379 12019 39399 12039
rect 39491 12019 39511 12039
rect 39587 12019 39607 12039
rect 39704 12019 39724 12039
rect 39800 12019 39820 12039
rect 41572 12014 41592 12034
rect 41668 12014 41688 12034
rect 41778 12014 41798 12034
rect 41874 12014 41894 12034
rect 41986 12014 42006 12034
rect 42082 12014 42102 12034
rect 42199 12014 42219 12034
rect 42295 12014 42315 12034
rect 901 11514 921 11534
rect 997 11514 1017 11534
rect 1114 11514 1134 11534
rect 1210 11514 1230 11534
rect 1322 11514 1342 11534
rect 1418 11514 1438 11534
rect 1528 11514 1548 11534
rect 1624 11514 1644 11534
rect 3439 11511 3459 11531
rect 3535 11511 3555 11531
rect 3652 11511 3672 11531
rect 3748 11511 3768 11531
rect 3860 11511 3880 11531
rect 3956 11511 3976 11531
rect 4066 11511 4086 11531
rect 4162 11511 4182 11531
rect 11609 11508 11629 11528
rect 8143 11347 8163 11367
rect 8239 11347 8259 11367
rect 8349 11347 8369 11367
rect 8445 11347 8465 11367
rect 8557 11347 8577 11367
rect 8653 11347 8673 11367
rect 8770 11347 8790 11367
rect 11705 11508 11725 11528
rect 11822 11508 11842 11528
rect 11918 11508 11938 11528
rect 12030 11508 12050 11528
rect 12126 11508 12146 11528
rect 12236 11508 12256 11528
rect 12332 11508 12352 11528
rect 14147 11505 14167 11525
rect 8866 11347 8886 11367
rect 9191 11343 9211 11363
rect 9287 11343 9307 11363
rect 9397 11343 9417 11363
rect 9493 11343 9513 11363
rect 9605 11343 9625 11363
rect 9701 11343 9721 11363
rect 9818 11343 9838 11363
rect 9914 11343 9934 11363
rect 14243 11505 14263 11525
rect 14360 11505 14380 11525
rect 14456 11505 14476 11525
rect 14568 11505 14588 11525
rect 14664 11505 14684 11525
rect 14774 11505 14794 11525
rect 14870 11505 14890 11525
rect 22574 11512 22594 11532
rect 18851 11341 18871 11361
rect 18947 11341 18967 11361
rect 19057 11341 19077 11361
rect 19153 11341 19173 11361
rect 19265 11341 19285 11361
rect 19361 11341 19381 11361
rect 19478 11341 19498 11361
rect 22670 11512 22690 11532
rect 22787 11512 22807 11532
rect 22883 11512 22903 11532
rect 22995 11512 23015 11532
rect 23091 11512 23111 11532
rect 23201 11512 23221 11532
rect 23297 11512 23317 11532
rect 25112 11509 25132 11529
rect 19574 11341 19594 11361
rect 19899 11337 19919 11357
rect 19995 11337 20015 11357
rect 20105 11337 20125 11357
rect 20201 11337 20221 11357
rect 20313 11337 20333 11357
rect 20409 11337 20429 11357
rect 20526 11337 20546 11357
rect 20622 11337 20642 11357
rect 25208 11509 25228 11529
rect 25325 11509 25345 11529
rect 25421 11509 25441 11529
rect 25533 11509 25553 11529
rect 25629 11509 25649 11529
rect 25739 11509 25759 11529
rect 25835 11509 25855 11529
rect 33282 11506 33302 11526
rect 29816 11345 29836 11365
rect 29912 11345 29932 11365
rect 30022 11345 30042 11365
rect 30118 11345 30138 11365
rect 30230 11345 30250 11365
rect 30326 11345 30346 11365
rect 30443 11345 30463 11365
rect 33378 11506 33398 11526
rect 33495 11506 33515 11526
rect 33591 11506 33611 11526
rect 33703 11506 33723 11526
rect 33799 11506 33819 11526
rect 33909 11506 33929 11526
rect 34005 11506 34025 11526
rect 35820 11503 35840 11523
rect 30539 11345 30559 11365
rect 30864 11341 30884 11361
rect 30960 11341 30980 11361
rect 31070 11341 31090 11361
rect 31166 11341 31186 11361
rect 31278 11341 31298 11361
rect 31374 11341 31394 11361
rect 31491 11341 31511 11361
rect 31587 11341 31607 11361
rect 35916 11503 35936 11523
rect 36033 11503 36053 11523
rect 36129 11503 36149 11523
rect 36241 11503 36261 11523
rect 36337 11503 36357 11523
rect 36447 11503 36467 11523
rect 36543 11503 36563 11523
rect 40524 11339 40544 11359
rect 40620 11339 40640 11359
rect 40730 11339 40750 11359
rect 40826 11339 40846 11359
rect 40938 11339 40958 11359
rect 41034 11339 41054 11359
rect 41151 11339 41171 11359
rect 41247 11339 41267 11359
rect 41572 11335 41592 11355
rect 41668 11335 41688 11355
rect 41778 11335 41798 11355
rect 41874 11335 41894 11355
rect 41986 11335 42006 11355
rect 42082 11335 42102 11355
rect 42199 11335 42219 11355
rect 42295 11335 42315 11355
rect 902 10673 922 10693
rect 998 10673 1018 10693
rect 1115 10673 1135 10693
rect 1211 10673 1231 10693
rect 1323 10673 1343 10693
rect 1419 10673 1439 10693
rect 1529 10673 1549 10693
rect 1625 10673 1645 10693
rect 1950 10669 1970 10689
rect 2046 10669 2066 10689
rect 2163 10669 2183 10689
rect 2259 10669 2279 10689
rect 2371 10669 2391 10689
rect 2467 10669 2487 10689
rect 2577 10669 2597 10689
rect 2673 10669 2693 10689
rect 6654 10505 6674 10525
rect 6750 10505 6770 10525
rect 6860 10505 6880 10525
rect 6956 10505 6976 10525
rect 7068 10505 7088 10525
rect 7164 10505 7184 10525
rect 7281 10505 7301 10525
rect 11610 10667 11630 10687
rect 11706 10667 11726 10687
rect 11823 10667 11843 10687
rect 11919 10667 11939 10687
rect 12031 10667 12051 10687
rect 12127 10667 12147 10687
rect 12237 10667 12257 10687
rect 12333 10667 12353 10687
rect 12658 10663 12678 10683
rect 7377 10505 7397 10525
rect 9192 10502 9212 10522
rect 9288 10502 9308 10522
rect 9398 10502 9418 10522
rect 9494 10502 9514 10522
rect 9606 10502 9626 10522
rect 9702 10502 9722 10522
rect 9819 10502 9839 10522
rect 12754 10663 12774 10683
rect 12871 10663 12891 10683
rect 12967 10663 12987 10683
rect 13079 10663 13099 10683
rect 13175 10663 13195 10683
rect 13285 10663 13305 10683
rect 13381 10663 13401 10683
rect 9915 10502 9935 10522
rect 17362 10499 17382 10519
rect 17458 10499 17478 10519
rect 17568 10499 17588 10519
rect 17664 10499 17684 10519
rect 17776 10499 17796 10519
rect 17872 10499 17892 10519
rect 17989 10499 18009 10519
rect 22575 10671 22595 10691
rect 22671 10671 22691 10691
rect 22788 10671 22808 10691
rect 22884 10671 22904 10691
rect 22996 10671 23016 10691
rect 23092 10671 23112 10691
rect 23202 10671 23222 10691
rect 23298 10671 23318 10691
rect 23623 10667 23643 10687
rect 18085 10499 18105 10519
rect 19900 10496 19920 10516
rect 19996 10496 20016 10516
rect 20106 10496 20126 10516
rect 20202 10496 20222 10516
rect 20314 10496 20334 10516
rect 20410 10496 20430 10516
rect 20527 10496 20547 10516
rect 23719 10667 23739 10687
rect 23836 10667 23856 10687
rect 23932 10667 23952 10687
rect 24044 10667 24064 10687
rect 24140 10667 24160 10687
rect 24250 10667 24270 10687
rect 24346 10667 24366 10687
rect 20623 10496 20643 10516
rect 28327 10503 28347 10523
rect 28423 10503 28443 10523
rect 28533 10503 28553 10523
rect 28629 10503 28649 10523
rect 28741 10503 28761 10523
rect 28837 10503 28857 10523
rect 28954 10503 28974 10523
rect 33283 10665 33303 10685
rect 33379 10665 33399 10685
rect 33496 10665 33516 10685
rect 33592 10665 33612 10685
rect 33704 10665 33724 10685
rect 33800 10665 33820 10685
rect 33910 10665 33930 10685
rect 34006 10665 34026 10685
rect 34331 10661 34351 10681
rect 29050 10503 29070 10523
rect 30865 10500 30885 10520
rect 30961 10500 30981 10520
rect 31071 10500 31091 10520
rect 31167 10500 31187 10520
rect 31279 10500 31299 10520
rect 31375 10500 31395 10520
rect 31492 10500 31512 10520
rect 34427 10661 34447 10681
rect 34544 10661 34564 10681
rect 34640 10661 34660 10681
rect 34752 10661 34772 10681
rect 34848 10661 34868 10681
rect 34958 10661 34978 10681
rect 35054 10661 35074 10681
rect 31588 10500 31608 10520
rect 39035 10497 39055 10517
rect 39131 10497 39151 10517
rect 39241 10497 39261 10517
rect 39337 10497 39357 10517
rect 39449 10497 39469 10517
rect 39545 10497 39565 10517
rect 39662 10497 39682 10517
rect 39758 10497 39778 10517
rect 41573 10494 41593 10514
rect 41669 10494 41689 10514
rect 41779 10494 41799 10514
rect 41875 10494 41895 10514
rect 41987 10494 42007 10514
rect 42083 10494 42103 10514
rect 42200 10494 42220 10514
rect 42296 10494 42316 10514
rect 902 9994 922 10014
rect 998 9994 1018 10014
rect 1115 9994 1135 10014
rect 1211 9994 1231 10014
rect 1323 9994 1343 10014
rect 1419 9994 1439 10014
rect 1529 9994 1549 10014
rect 1625 9994 1645 10014
rect 3397 9989 3417 10009
rect 3493 9989 3513 10009
rect 3610 9989 3630 10009
rect 3706 9989 3726 10009
rect 3818 9989 3838 10009
rect 3914 9989 3934 10009
rect 4024 9989 4044 10009
rect 4120 9989 4140 10009
rect 11610 9988 11630 10008
rect 8144 9827 8164 9847
rect 8240 9827 8260 9847
rect 8350 9827 8370 9847
rect 8446 9827 8466 9847
rect 8558 9827 8578 9847
rect 8654 9827 8674 9847
rect 8771 9827 8791 9847
rect 11706 9988 11726 10008
rect 11823 9988 11843 10008
rect 11919 9988 11939 10008
rect 12031 9988 12051 10008
rect 12127 9988 12147 10008
rect 12237 9988 12257 10008
rect 12333 9988 12353 10008
rect 14105 9983 14125 10003
rect 8867 9827 8887 9847
rect 9192 9823 9212 9843
rect 9288 9823 9308 9843
rect 9398 9823 9418 9843
rect 9494 9823 9514 9843
rect 9606 9823 9626 9843
rect 9702 9823 9722 9843
rect 9819 9823 9839 9843
rect 9915 9823 9935 9843
rect 14201 9983 14221 10003
rect 14318 9983 14338 10003
rect 14414 9983 14434 10003
rect 14526 9983 14546 10003
rect 14622 9983 14642 10003
rect 14732 9983 14752 10003
rect 14828 9983 14848 10003
rect 22575 9992 22595 10012
rect 18852 9821 18872 9841
rect 18948 9821 18968 9841
rect 19058 9821 19078 9841
rect 19154 9821 19174 9841
rect 19266 9821 19286 9841
rect 19362 9821 19382 9841
rect 19479 9821 19499 9841
rect 22671 9992 22691 10012
rect 22788 9992 22808 10012
rect 22884 9992 22904 10012
rect 22996 9992 23016 10012
rect 23092 9992 23112 10012
rect 23202 9992 23222 10012
rect 23298 9992 23318 10012
rect 25070 9987 25090 10007
rect 19575 9821 19595 9841
rect 19900 9817 19920 9837
rect 19996 9817 20016 9837
rect 20106 9817 20126 9837
rect 20202 9817 20222 9837
rect 20314 9817 20334 9837
rect 20410 9817 20430 9837
rect 20527 9817 20547 9837
rect 20623 9817 20643 9837
rect 25166 9987 25186 10007
rect 25283 9987 25303 10007
rect 25379 9987 25399 10007
rect 25491 9987 25511 10007
rect 25587 9987 25607 10007
rect 25697 9987 25717 10007
rect 25793 9987 25813 10007
rect 33283 9986 33303 10006
rect 29817 9825 29837 9845
rect 29913 9825 29933 9845
rect 30023 9825 30043 9845
rect 30119 9825 30139 9845
rect 30231 9825 30251 9845
rect 30327 9825 30347 9845
rect 30444 9825 30464 9845
rect 33379 9986 33399 10006
rect 33496 9986 33516 10006
rect 33592 9986 33612 10006
rect 33704 9986 33724 10006
rect 33800 9986 33820 10006
rect 33910 9986 33930 10006
rect 34006 9986 34026 10006
rect 35778 9981 35798 10001
rect 30540 9825 30560 9845
rect 30865 9821 30885 9841
rect 30961 9821 30981 9841
rect 31071 9821 31091 9841
rect 31167 9821 31187 9841
rect 31279 9821 31299 9841
rect 31375 9821 31395 9841
rect 31492 9821 31512 9841
rect 31588 9821 31608 9841
rect 35874 9981 35894 10001
rect 35991 9981 36011 10001
rect 36087 9981 36107 10001
rect 36199 9981 36219 10001
rect 36295 9981 36315 10001
rect 36405 9981 36425 10001
rect 36501 9981 36521 10001
rect 40525 9819 40545 9839
rect 40621 9819 40641 9839
rect 40731 9819 40751 9839
rect 40827 9819 40847 9839
rect 40939 9819 40959 9839
rect 41035 9819 41055 9839
rect 41152 9819 41172 9839
rect 41248 9819 41268 9839
rect 41573 9815 41593 9835
rect 41669 9815 41689 9835
rect 41779 9815 41799 9835
rect 41875 9815 41895 9835
rect 41987 9815 42007 9835
rect 42083 9815 42103 9835
rect 42200 9815 42220 9835
rect 42296 9815 42316 9835
rect 902 9226 922 9246
rect 998 9226 1018 9246
rect 1115 9226 1135 9246
rect 1211 9226 1231 9246
rect 1323 9226 1343 9246
rect 1419 9226 1439 9246
rect 1529 9226 1549 9246
rect 1625 9226 1645 9246
rect 1950 9222 1970 9242
rect 2046 9222 2066 9242
rect 2163 9222 2183 9242
rect 2259 9222 2279 9242
rect 2371 9222 2391 9242
rect 2467 9222 2487 9242
rect 2577 9222 2597 9242
rect 2673 9222 2693 9242
rect 6697 9060 6717 9080
rect 6793 9060 6813 9080
rect 6903 9060 6923 9080
rect 6999 9060 7019 9080
rect 7111 9060 7131 9080
rect 7207 9060 7227 9080
rect 7324 9060 7344 9080
rect 11610 9220 11630 9240
rect 11706 9220 11726 9240
rect 11823 9220 11843 9240
rect 11919 9220 11939 9240
rect 12031 9220 12051 9240
rect 12127 9220 12147 9240
rect 12237 9220 12257 9240
rect 12333 9220 12353 9240
rect 12658 9216 12678 9236
rect 7420 9060 7440 9080
rect 9192 9055 9212 9075
rect 9288 9055 9308 9075
rect 9398 9055 9418 9075
rect 9494 9055 9514 9075
rect 9606 9055 9626 9075
rect 9702 9055 9722 9075
rect 9819 9055 9839 9075
rect 12754 9216 12774 9236
rect 12871 9216 12891 9236
rect 12967 9216 12987 9236
rect 13079 9216 13099 9236
rect 13175 9216 13195 9236
rect 13285 9216 13305 9236
rect 13381 9216 13401 9236
rect 9915 9055 9935 9075
rect 17405 9054 17425 9074
rect 17501 9054 17521 9074
rect 17611 9054 17631 9074
rect 17707 9054 17727 9074
rect 17819 9054 17839 9074
rect 17915 9054 17935 9074
rect 18032 9054 18052 9074
rect 22575 9224 22595 9244
rect 22671 9224 22691 9244
rect 22788 9224 22808 9244
rect 22884 9224 22904 9244
rect 22996 9224 23016 9244
rect 23092 9224 23112 9244
rect 23202 9224 23222 9244
rect 23298 9224 23318 9244
rect 23623 9220 23643 9240
rect 18128 9054 18148 9074
rect 19900 9049 19920 9069
rect 19996 9049 20016 9069
rect 20106 9049 20126 9069
rect 20202 9049 20222 9069
rect 20314 9049 20334 9069
rect 20410 9049 20430 9069
rect 20527 9049 20547 9069
rect 23719 9220 23739 9240
rect 23836 9220 23856 9240
rect 23932 9220 23952 9240
rect 24044 9220 24064 9240
rect 24140 9220 24160 9240
rect 24250 9220 24270 9240
rect 24346 9220 24366 9240
rect 20623 9049 20643 9069
rect 28370 9058 28390 9078
rect 28466 9058 28486 9078
rect 28576 9058 28596 9078
rect 28672 9058 28692 9078
rect 28784 9058 28804 9078
rect 28880 9058 28900 9078
rect 28997 9058 29017 9078
rect 33283 9218 33303 9238
rect 33379 9218 33399 9238
rect 33496 9218 33516 9238
rect 33592 9218 33612 9238
rect 33704 9218 33724 9238
rect 33800 9218 33820 9238
rect 33910 9218 33930 9238
rect 34006 9218 34026 9238
rect 34331 9214 34351 9234
rect 29093 9058 29113 9078
rect 30865 9053 30885 9073
rect 30961 9053 30981 9073
rect 31071 9053 31091 9073
rect 31167 9053 31187 9073
rect 31279 9053 31299 9073
rect 31375 9053 31395 9073
rect 31492 9053 31512 9073
rect 34427 9214 34447 9234
rect 34544 9214 34564 9234
rect 34640 9214 34660 9234
rect 34752 9214 34772 9234
rect 34848 9214 34868 9234
rect 34958 9214 34978 9234
rect 35054 9214 35074 9234
rect 31588 9053 31608 9073
rect 39078 9052 39098 9072
rect 39174 9052 39194 9072
rect 39284 9052 39304 9072
rect 39380 9052 39400 9072
rect 39492 9052 39512 9072
rect 39588 9052 39608 9072
rect 39705 9052 39725 9072
rect 39801 9052 39821 9072
rect 41573 9047 41593 9067
rect 41669 9047 41689 9067
rect 41779 9047 41799 9067
rect 41875 9047 41895 9067
rect 41987 9047 42007 9067
rect 42083 9047 42103 9067
rect 42200 9047 42220 9067
rect 42296 9047 42316 9067
rect 902 8547 922 8567
rect 998 8547 1018 8567
rect 1115 8547 1135 8567
rect 1211 8547 1231 8567
rect 1323 8547 1343 8567
rect 1419 8547 1439 8567
rect 1529 8547 1549 8567
rect 1625 8547 1645 8567
rect 4505 8538 4525 8558
rect 4601 8538 4621 8558
rect 4718 8538 4738 8558
rect 4814 8538 4834 8558
rect 4926 8538 4946 8558
rect 5022 8538 5042 8558
rect 5132 8538 5152 8558
rect 5228 8538 5248 8558
rect 11610 8541 11630 8561
rect 8144 8380 8164 8400
rect 8240 8380 8260 8400
rect 8350 8380 8370 8400
rect 8446 8380 8466 8400
rect 8558 8380 8578 8400
rect 8654 8380 8674 8400
rect 8771 8380 8791 8400
rect 11706 8541 11726 8561
rect 11823 8541 11843 8561
rect 11919 8541 11939 8561
rect 12031 8541 12051 8561
rect 12127 8541 12147 8561
rect 12237 8541 12257 8561
rect 12333 8541 12353 8561
rect 15213 8532 15233 8552
rect 8867 8380 8887 8400
rect 9192 8376 9212 8396
rect 9288 8376 9308 8396
rect 9398 8376 9418 8396
rect 9494 8376 9514 8396
rect 9606 8376 9626 8396
rect 9702 8376 9722 8396
rect 9819 8376 9839 8396
rect 9915 8376 9935 8396
rect 15309 8532 15329 8552
rect 15426 8532 15446 8552
rect 15522 8532 15542 8552
rect 15634 8532 15654 8552
rect 15730 8532 15750 8552
rect 15840 8532 15860 8552
rect 15936 8532 15956 8552
rect 22575 8545 22595 8565
rect 18852 8374 18872 8394
rect 18948 8374 18968 8394
rect 19058 8374 19078 8394
rect 19154 8374 19174 8394
rect 19266 8374 19286 8394
rect 19362 8374 19382 8394
rect 19479 8374 19499 8394
rect 22671 8545 22691 8565
rect 22788 8545 22808 8565
rect 22884 8545 22904 8565
rect 22996 8545 23016 8565
rect 23092 8545 23112 8565
rect 23202 8545 23222 8565
rect 23298 8545 23318 8565
rect 26178 8536 26198 8556
rect 19575 8374 19595 8394
rect 19900 8370 19920 8390
rect 19996 8370 20016 8390
rect 20106 8370 20126 8390
rect 20202 8370 20222 8390
rect 20314 8370 20334 8390
rect 20410 8370 20430 8390
rect 20527 8370 20547 8390
rect 20623 8370 20643 8390
rect 26274 8536 26294 8556
rect 26391 8536 26411 8556
rect 26487 8536 26507 8556
rect 26599 8536 26619 8556
rect 26695 8536 26715 8556
rect 26805 8536 26825 8556
rect 26901 8536 26921 8556
rect 33283 8539 33303 8559
rect 29817 8378 29837 8398
rect 29913 8378 29933 8398
rect 30023 8378 30043 8398
rect 30119 8378 30139 8398
rect 30231 8378 30251 8398
rect 30327 8378 30347 8398
rect 30444 8378 30464 8398
rect 33379 8539 33399 8559
rect 33496 8539 33516 8559
rect 33592 8539 33612 8559
rect 33704 8539 33724 8559
rect 33800 8539 33820 8559
rect 33910 8539 33930 8559
rect 34006 8539 34026 8559
rect 36886 8530 36906 8550
rect 30540 8378 30560 8398
rect 30865 8374 30885 8394
rect 30961 8374 30981 8394
rect 31071 8374 31091 8394
rect 31167 8374 31187 8394
rect 31279 8374 31299 8394
rect 31375 8374 31395 8394
rect 31492 8374 31512 8394
rect 31588 8374 31608 8394
rect 36982 8530 37002 8550
rect 37099 8530 37119 8550
rect 37195 8530 37215 8550
rect 37307 8530 37327 8550
rect 37403 8530 37423 8550
rect 37513 8530 37533 8550
rect 37609 8530 37629 8550
rect 40525 8372 40545 8392
rect 40621 8372 40641 8392
rect 40731 8372 40751 8392
rect 40827 8372 40847 8392
rect 40939 8372 40959 8392
rect 41035 8372 41055 8392
rect 41152 8372 41172 8392
rect 41248 8372 41268 8392
rect 41573 8368 41593 8388
rect 41669 8368 41689 8388
rect 41779 8368 41799 8388
rect 41875 8368 41895 8388
rect 41987 8368 42007 8388
rect 42083 8368 42103 8388
rect 42200 8368 42220 8388
rect 42296 8368 42316 8388
rect 899 7632 919 7652
rect 995 7632 1015 7652
rect 1112 7632 1132 7652
rect 1208 7632 1228 7652
rect 1320 7632 1340 7652
rect 1416 7632 1436 7652
rect 1526 7632 1546 7652
rect 1622 7632 1642 7652
rect 1947 7628 1967 7648
rect 2043 7628 2063 7648
rect 2160 7628 2180 7648
rect 2256 7628 2276 7648
rect 2368 7628 2388 7648
rect 2464 7628 2484 7648
rect 2574 7628 2594 7648
rect 2670 7628 2690 7648
rect 5586 7470 5606 7490
rect 5682 7470 5702 7490
rect 5792 7470 5812 7490
rect 5888 7470 5908 7490
rect 6000 7470 6020 7490
rect 6096 7470 6116 7490
rect 6213 7470 6233 7490
rect 11607 7626 11627 7646
rect 11703 7626 11723 7646
rect 11820 7626 11840 7646
rect 11916 7626 11936 7646
rect 12028 7626 12048 7646
rect 12124 7626 12144 7646
rect 12234 7626 12254 7646
rect 12330 7626 12350 7646
rect 12655 7622 12675 7642
rect 6309 7470 6329 7490
rect 9189 7461 9209 7481
rect 9285 7461 9305 7481
rect 9395 7461 9415 7481
rect 9491 7461 9511 7481
rect 9603 7461 9623 7481
rect 9699 7461 9719 7481
rect 9816 7461 9836 7481
rect 12751 7622 12771 7642
rect 12868 7622 12888 7642
rect 12964 7622 12984 7642
rect 13076 7622 13096 7642
rect 13172 7622 13192 7642
rect 13282 7622 13302 7642
rect 13378 7622 13398 7642
rect 9912 7461 9932 7481
rect 16294 7464 16314 7484
rect 16390 7464 16410 7484
rect 16500 7464 16520 7484
rect 16596 7464 16616 7484
rect 16708 7464 16728 7484
rect 16804 7464 16824 7484
rect 16921 7464 16941 7484
rect 22572 7630 22592 7650
rect 22668 7630 22688 7650
rect 22785 7630 22805 7650
rect 22881 7630 22901 7650
rect 22993 7630 23013 7650
rect 23089 7630 23109 7650
rect 23199 7630 23219 7650
rect 23295 7630 23315 7650
rect 23620 7626 23640 7646
rect 17017 7464 17037 7484
rect 19897 7455 19917 7475
rect 19993 7455 20013 7475
rect 20103 7455 20123 7475
rect 20199 7455 20219 7475
rect 20311 7455 20331 7475
rect 20407 7455 20427 7475
rect 20524 7455 20544 7475
rect 23716 7626 23736 7646
rect 23833 7626 23853 7646
rect 23929 7626 23949 7646
rect 24041 7626 24061 7646
rect 24137 7626 24157 7646
rect 24247 7626 24267 7646
rect 24343 7626 24363 7646
rect 20620 7455 20640 7475
rect 27259 7468 27279 7488
rect 27355 7468 27375 7488
rect 27465 7468 27485 7488
rect 27561 7468 27581 7488
rect 27673 7468 27693 7488
rect 27769 7468 27789 7488
rect 27886 7468 27906 7488
rect 33280 7624 33300 7644
rect 33376 7624 33396 7644
rect 33493 7624 33513 7644
rect 33589 7624 33609 7644
rect 33701 7624 33721 7644
rect 33797 7624 33817 7644
rect 33907 7624 33927 7644
rect 34003 7624 34023 7644
rect 34328 7620 34348 7640
rect 27982 7468 28002 7488
rect 30862 7459 30882 7479
rect 30958 7459 30978 7479
rect 31068 7459 31088 7479
rect 31164 7459 31184 7479
rect 31276 7459 31296 7479
rect 31372 7459 31392 7479
rect 31489 7459 31509 7479
rect 34424 7620 34444 7640
rect 34541 7620 34561 7640
rect 34637 7620 34657 7640
rect 34749 7620 34769 7640
rect 34845 7620 34865 7640
rect 34955 7620 34975 7640
rect 35051 7620 35071 7640
rect 31585 7459 31605 7479
rect 37967 7462 37987 7482
rect 38063 7462 38083 7482
rect 38173 7462 38193 7482
rect 38269 7462 38289 7482
rect 38381 7462 38401 7482
rect 38477 7462 38497 7482
rect 38594 7462 38614 7482
rect 38690 7462 38710 7482
rect 41570 7453 41590 7473
rect 41666 7453 41686 7473
rect 41776 7453 41796 7473
rect 41872 7453 41892 7473
rect 41984 7453 42004 7473
rect 42080 7453 42100 7473
rect 42197 7453 42217 7473
rect 42293 7453 42313 7473
rect 899 6953 919 6973
rect 995 6953 1015 6973
rect 1112 6953 1132 6973
rect 1208 6953 1228 6973
rect 1320 6953 1340 6973
rect 1416 6953 1436 6973
rect 1526 6953 1546 6973
rect 1622 6953 1642 6973
rect 3394 6948 3414 6968
rect 3490 6948 3510 6968
rect 3607 6948 3627 6968
rect 3703 6948 3723 6968
rect 3815 6948 3835 6968
rect 3911 6948 3931 6968
rect 4021 6948 4041 6968
rect 4117 6948 4137 6968
rect 11607 6947 11627 6967
rect 8141 6786 8161 6806
rect 8237 6786 8257 6806
rect 8347 6786 8367 6806
rect 8443 6786 8463 6806
rect 8555 6786 8575 6806
rect 8651 6786 8671 6806
rect 8768 6786 8788 6806
rect 11703 6947 11723 6967
rect 11820 6947 11840 6967
rect 11916 6947 11936 6967
rect 12028 6947 12048 6967
rect 12124 6947 12144 6967
rect 12234 6947 12254 6967
rect 12330 6947 12350 6967
rect 14102 6942 14122 6962
rect 8864 6786 8884 6806
rect 9189 6782 9209 6802
rect 9285 6782 9305 6802
rect 9395 6782 9415 6802
rect 9491 6782 9511 6802
rect 9603 6782 9623 6802
rect 9699 6782 9719 6802
rect 9816 6782 9836 6802
rect 9912 6782 9932 6802
rect 14198 6942 14218 6962
rect 14315 6942 14335 6962
rect 14411 6942 14431 6962
rect 14523 6942 14543 6962
rect 14619 6942 14639 6962
rect 14729 6942 14749 6962
rect 14825 6942 14845 6962
rect 22572 6951 22592 6971
rect 18849 6780 18869 6800
rect 18945 6780 18965 6800
rect 19055 6780 19075 6800
rect 19151 6780 19171 6800
rect 19263 6780 19283 6800
rect 19359 6780 19379 6800
rect 19476 6780 19496 6800
rect 22668 6951 22688 6971
rect 22785 6951 22805 6971
rect 22881 6951 22901 6971
rect 22993 6951 23013 6971
rect 23089 6951 23109 6971
rect 23199 6951 23219 6971
rect 23295 6951 23315 6971
rect 25067 6946 25087 6966
rect 19572 6780 19592 6800
rect 19897 6776 19917 6796
rect 19993 6776 20013 6796
rect 20103 6776 20123 6796
rect 20199 6776 20219 6796
rect 20311 6776 20331 6796
rect 20407 6776 20427 6796
rect 20524 6776 20544 6796
rect 20620 6776 20640 6796
rect 25163 6946 25183 6966
rect 25280 6946 25300 6966
rect 25376 6946 25396 6966
rect 25488 6946 25508 6966
rect 25584 6946 25604 6966
rect 25694 6946 25714 6966
rect 25790 6946 25810 6966
rect 33280 6945 33300 6965
rect 29814 6784 29834 6804
rect 29910 6784 29930 6804
rect 30020 6784 30040 6804
rect 30116 6784 30136 6804
rect 30228 6784 30248 6804
rect 30324 6784 30344 6804
rect 30441 6784 30461 6804
rect 33376 6945 33396 6965
rect 33493 6945 33513 6965
rect 33589 6945 33609 6965
rect 33701 6945 33721 6965
rect 33797 6945 33817 6965
rect 33907 6945 33927 6965
rect 34003 6945 34023 6965
rect 35775 6940 35795 6960
rect 30537 6784 30557 6804
rect 30862 6780 30882 6800
rect 30958 6780 30978 6800
rect 31068 6780 31088 6800
rect 31164 6780 31184 6800
rect 31276 6780 31296 6800
rect 31372 6780 31392 6800
rect 31489 6780 31509 6800
rect 31585 6780 31605 6800
rect 35871 6940 35891 6960
rect 35988 6940 36008 6960
rect 36084 6940 36104 6960
rect 36196 6940 36216 6960
rect 36292 6940 36312 6960
rect 36402 6940 36422 6960
rect 36498 6940 36518 6960
rect 40522 6778 40542 6798
rect 40618 6778 40638 6798
rect 40728 6778 40748 6798
rect 40824 6778 40844 6798
rect 40936 6778 40956 6798
rect 41032 6778 41052 6798
rect 41149 6778 41169 6798
rect 41245 6778 41265 6798
rect 41570 6774 41590 6794
rect 41666 6774 41686 6794
rect 41776 6774 41796 6794
rect 41872 6774 41892 6794
rect 41984 6774 42004 6794
rect 42080 6774 42100 6794
rect 42197 6774 42217 6794
rect 42293 6774 42313 6794
rect 899 6185 919 6205
rect 995 6185 1015 6205
rect 1112 6185 1132 6205
rect 1208 6185 1228 6205
rect 1320 6185 1340 6205
rect 1416 6185 1436 6205
rect 1526 6185 1546 6205
rect 1622 6185 1642 6205
rect 1947 6181 1967 6201
rect 2043 6181 2063 6201
rect 2160 6181 2180 6201
rect 2256 6181 2276 6201
rect 2368 6181 2388 6201
rect 2464 6181 2484 6201
rect 2574 6181 2594 6201
rect 2670 6181 2690 6201
rect 6694 6019 6714 6039
rect 6790 6019 6810 6039
rect 6900 6019 6920 6039
rect 6996 6019 7016 6039
rect 7108 6019 7128 6039
rect 7204 6019 7224 6039
rect 7321 6019 7341 6039
rect 11607 6179 11627 6199
rect 11703 6179 11723 6199
rect 11820 6179 11840 6199
rect 11916 6179 11936 6199
rect 12028 6179 12048 6199
rect 12124 6179 12144 6199
rect 12234 6179 12254 6199
rect 12330 6179 12350 6199
rect 12655 6175 12675 6195
rect 7417 6019 7437 6039
rect 9189 6014 9209 6034
rect 9285 6014 9305 6034
rect 9395 6014 9415 6034
rect 9491 6014 9511 6034
rect 9603 6014 9623 6034
rect 9699 6014 9719 6034
rect 9816 6014 9836 6034
rect 12751 6175 12771 6195
rect 12868 6175 12888 6195
rect 12964 6175 12984 6195
rect 13076 6175 13096 6195
rect 13172 6175 13192 6195
rect 13282 6175 13302 6195
rect 13378 6175 13398 6195
rect 9912 6014 9932 6034
rect 17402 6013 17422 6033
rect 17498 6013 17518 6033
rect 17608 6013 17628 6033
rect 17704 6013 17724 6033
rect 17816 6013 17836 6033
rect 17912 6013 17932 6033
rect 18029 6013 18049 6033
rect 22572 6183 22592 6203
rect 22668 6183 22688 6203
rect 22785 6183 22805 6203
rect 22881 6183 22901 6203
rect 22993 6183 23013 6203
rect 23089 6183 23109 6203
rect 23199 6183 23219 6203
rect 23295 6183 23315 6203
rect 23620 6179 23640 6199
rect 18125 6013 18145 6033
rect 19897 6008 19917 6028
rect 19993 6008 20013 6028
rect 20103 6008 20123 6028
rect 20199 6008 20219 6028
rect 20311 6008 20331 6028
rect 20407 6008 20427 6028
rect 20524 6008 20544 6028
rect 23716 6179 23736 6199
rect 23833 6179 23853 6199
rect 23929 6179 23949 6199
rect 24041 6179 24061 6199
rect 24137 6179 24157 6199
rect 24247 6179 24267 6199
rect 24343 6179 24363 6199
rect 20620 6008 20640 6028
rect 28367 6017 28387 6037
rect 28463 6017 28483 6037
rect 28573 6017 28593 6037
rect 28669 6017 28689 6037
rect 28781 6017 28801 6037
rect 28877 6017 28897 6037
rect 28994 6017 29014 6037
rect 33280 6177 33300 6197
rect 33376 6177 33396 6197
rect 33493 6177 33513 6197
rect 33589 6177 33609 6197
rect 33701 6177 33721 6197
rect 33797 6177 33817 6197
rect 33907 6177 33927 6197
rect 34003 6177 34023 6197
rect 34328 6173 34348 6193
rect 29090 6017 29110 6037
rect 30862 6012 30882 6032
rect 30958 6012 30978 6032
rect 31068 6012 31088 6032
rect 31164 6012 31184 6032
rect 31276 6012 31296 6032
rect 31372 6012 31392 6032
rect 31489 6012 31509 6032
rect 34424 6173 34444 6193
rect 34541 6173 34561 6193
rect 34637 6173 34657 6193
rect 34749 6173 34769 6193
rect 34845 6173 34865 6193
rect 34955 6173 34975 6193
rect 35051 6173 35071 6193
rect 31585 6012 31605 6032
rect 39075 6011 39095 6031
rect 39171 6011 39191 6031
rect 39281 6011 39301 6031
rect 39377 6011 39397 6031
rect 39489 6011 39509 6031
rect 39585 6011 39605 6031
rect 39702 6011 39722 6031
rect 39798 6011 39818 6031
rect 41570 6006 41590 6026
rect 41666 6006 41686 6026
rect 41776 6006 41796 6026
rect 41872 6006 41892 6026
rect 41984 6006 42004 6026
rect 42080 6006 42100 6026
rect 42197 6006 42217 6026
rect 42293 6006 42313 6026
rect 899 5506 919 5526
rect 995 5506 1015 5526
rect 1112 5506 1132 5526
rect 1208 5506 1228 5526
rect 1320 5506 1340 5526
rect 1416 5506 1436 5526
rect 1526 5506 1546 5526
rect 1622 5506 1642 5526
rect 3437 5503 3457 5523
rect 3533 5503 3553 5523
rect 3650 5503 3670 5523
rect 3746 5503 3766 5523
rect 3858 5503 3878 5523
rect 3954 5503 3974 5523
rect 4064 5503 4084 5523
rect 4160 5503 4180 5523
rect 11607 5500 11627 5520
rect 8141 5339 8161 5359
rect 8237 5339 8257 5359
rect 8347 5339 8367 5359
rect 8443 5339 8463 5359
rect 8555 5339 8575 5359
rect 8651 5339 8671 5359
rect 8768 5339 8788 5359
rect 11703 5500 11723 5520
rect 11820 5500 11840 5520
rect 11916 5500 11936 5520
rect 12028 5500 12048 5520
rect 12124 5500 12144 5520
rect 12234 5500 12254 5520
rect 12330 5500 12350 5520
rect 14145 5497 14165 5517
rect 8864 5339 8884 5359
rect 9189 5335 9209 5355
rect 9285 5335 9305 5355
rect 9395 5335 9415 5355
rect 9491 5335 9511 5355
rect 9603 5335 9623 5355
rect 9699 5335 9719 5355
rect 9816 5335 9836 5355
rect 9912 5335 9932 5355
rect 14241 5497 14261 5517
rect 14358 5497 14378 5517
rect 14454 5497 14474 5517
rect 14566 5497 14586 5517
rect 14662 5497 14682 5517
rect 14772 5497 14792 5517
rect 14868 5497 14888 5517
rect 22572 5504 22592 5524
rect 18849 5333 18869 5353
rect 18945 5333 18965 5353
rect 19055 5333 19075 5353
rect 19151 5333 19171 5353
rect 19263 5333 19283 5353
rect 19359 5333 19379 5353
rect 19476 5333 19496 5353
rect 22668 5504 22688 5524
rect 22785 5504 22805 5524
rect 22881 5504 22901 5524
rect 22993 5504 23013 5524
rect 23089 5504 23109 5524
rect 23199 5504 23219 5524
rect 23295 5504 23315 5524
rect 25110 5501 25130 5521
rect 19572 5333 19592 5353
rect 19897 5329 19917 5349
rect 19993 5329 20013 5349
rect 20103 5329 20123 5349
rect 20199 5329 20219 5349
rect 20311 5329 20331 5349
rect 20407 5329 20427 5349
rect 20524 5329 20544 5349
rect 20620 5329 20640 5349
rect 25206 5501 25226 5521
rect 25323 5501 25343 5521
rect 25419 5501 25439 5521
rect 25531 5501 25551 5521
rect 25627 5501 25647 5521
rect 25737 5501 25757 5521
rect 25833 5501 25853 5521
rect 33280 5498 33300 5518
rect 29814 5337 29834 5357
rect 29910 5337 29930 5357
rect 30020 5337 30040 5357
rect 30116 5337 30136 5357
rect 30228 5337 30248 5357
rect 30324 5337 30344 5357
rect 30441 5337 30461 5357
rect 33376 5498 33396 5518
rect 33493 5498 33513 5518
rect 33589 5498 33609 5518
rect 33701 5498 33721 5518
rect 33797 5498 33817 5518
rect 33907 5498 33927 5518
rect 34003 5498 34023 5518
rect 35818 5495 35838 5515
rect 30537 5337 30557 5357
rect 30862 5333 30882 5353
rect 30958 5333 30978 5353
rect 31068 5333 31088 5353
rect 31164 5333 31184 5353
rect 31276 5333 31296 5353
rect 31372 5333 31392 5353
rect 31489 5333 31509 5353
rect 31585 5333 31605 5353
rect 35914 5495 35934 5515
rect 36031 5495 36051 5515
rect 36127 5495 36147 5515
rect 36239 5495 36259 5515
rect 36335 5495 36355 5515
rect 36445 5495 36465 5515
rect 36541 5495 36561 5515
rect 40522 5331 40542 5351
rect 40618 5331 40638 5351
rect 40728 5331 40748 5351
rect 40824 5331 40844 5351
rect 40936 5331 40956 5351
rect 41032 5331 41052 5351
rect 41149 5331 41169 5351
rect 41245 5331 41265 5351
rect 41570 5327 41590 5347
rect 41666 5327 41686 5347
rect 41776 5327 41796 5347
rect 41872 5327 41892 5347
rect 41984 5327 42004 5347
rect 42080 5327 42100 5347
rect 42197 5327 42217 5347
rect 42293 5327 42313 5347
rect 900 4665 920 4685
rect 996 4665 1016 4685
rect 1113 4665 1133 4685
rect 1209 4665 1229 4685
rect 1321 4665 1341 4685
rect 1417 4665 1437 4685
rect 1527 4665 1547 4685
rect 1623 4665 1643 4685
rect 1948 4661 1968 4681
rect 2044 4661 2064 4681
rect 2161 4661 2181 4681
rect 2257 4661 2277 4681
rect 2369 4661 2389 4681
rect 2465 4661 2485 4681
rect 2575 4661 2595 4681
rect 2671 4661 2691 4681
rect 4850 4667 4870 4687
rect 4946 4667 4966 4687
rect 5063 4667 5083 4687
rect 5159 4667 5179 4687
rect 5271 4667 5291 4687
rect 5367 4667 5387 4687
rect 5477 4667 5497 4687
rect 5573 4667 5593 4687
rect 6652 4497 6672 4517
rect 6748 4497 6768 4517
rect 6858 4497 6878 4517
rect 6954 4497 6974 4517
rect 7066 4497 7086 4517
rect 7162 4497 7182 4517
rect 7279 4497 7299 4517
rect 11608 4659 11628 4679
rect 11704 4659 11724 4679
rect 11821 4659 11841 4679
rect 11917 4659 11937 4679
rect 12029 4659 12049 4679
rect 12125 4659 12145 4679
rect 12235 4659 12255 4679
rect 12331 4659 12351 4679
rect 12656 4655 12676 4675
rect 7375 4497 7395 4517
rect 9190 4494 9210 4514
rect 9286 4494 9306 4514
rect 9396 4494 9416 4514
rect 9492 4494 9512 4514
rect 9604 4494 9624 4514
rect 9700 4494 9720 4514
rect 9817 4494 9837 4514
rect 12752 4655 12772 4675
rect 12869 4655 12889 4675
rect 12965 4655 12985 4675
rect 13077 4655 13097 4675
rect 13173 4655 13193 4675
rect 13283 4655 13303 4675
rect 13379 4655 13399 4675
rect 15558 4661 15578 4681
rect 15654 4661 15674 4681
rect 15771 4661 15791 4681
rect 15867 4661 15887 4681
rect 15979 4661 15999 4681
rect 16075 4661 16095 4681
rect 16185 4661 16205 4681
rect 16281 4661 16301 4681
rect 9913 4494 9933 4514
rect 17360 4491 17380 4511
rect 17456 4491 17476 4511
rect 17566 4491 17586 4511
rect 17662 4491 17682 4511
rect 17774 4491 17794 4511
rect 17870 4491 17890 4511
rect 17987 4491 18007 4511
rect 22573 4663 22593 4683
rect 22669 4663 22689 4683
rect 22786 4663 22806 4683
rect 22882 4663 22902 4683
rect 22994 4663 23014 4683
rect 23090 4663 23110 4683
rect 23200 4663 23220 4683
rect 23296 4663 23316 4683
rect 23621 4659 23641 4679
rect 18083 4491 18103 4511
rect 19898 4488 19918 4508
rect 19994 4488 20014 4508
rect 20104 4488 20124 4508
rect 20200 4488 20220 4508
rect 20312 4488 20332 4508
rect 20408 4488 20428 4508
rect 20525 4488 20545 4508
rect 23717 4659 23737 4679
rect 23834 4659 23854 4679
rect 23930 4659 23950 4679
rect 24042 4659 24062 4679
rect 24138 4659 24158 4679
rect 24248 4659 24268 4679
rect 24344 4659 24364 4679
rect 26523 4665 26543 4685
rect 26619 4665 26639 4685
rect 26736 4665 26756 4685
rect 26832 4665 26852 4685
rect 26944 4665 26964 4685
rect 27040 4665 27060 4685
rect 27150 4665 27170 4685
rect 27246 4665 27266 4685
rect 20621 4488 20641 4508
rect 28325 4495 28345 4515
rect 28421 4495 28441 4515
rect 28531 4495 28551 4515
rect 28627 4495 28647 4515
rect 28739 4495 28759 4515
rect 28835 4495 28855 4515
rect 28952 4495 28972 4515
rect 33281 4657 33301 4677
rect 33377 4657 33397 4677
rect 33494 4657 33514 4677
rect 33590 4657 33610 4677
rect 33702 4657 33722 4677
rect 33798 4657 33818 4677
rect 33908 4657 33928 4677
rect 34004 4657 34024 4677
rect 34329 4653 34349 4673
rect 29048 4495 29068 4515
rect 30863 4492 30883 4512
rect 30959 4492 30979 4512
rect 31069 4492 31089 4512
rect 31165 4492 31185 4512
rect 31277 4492 31297 4512
rect 31373 4492 31393 4512
rect 31490 4492 31510 4512
rect 34425 4653 34445 4673
rect 34542 4653 34562 4673
rect 34638 4653 34658 4673
rect 34750 4653 34770 4673
rect 34846 4653 34866 4673
rect 34956 4653 34976 4673
rect 35052 4653 35072 4673
rect 37231 4659 37251 4679
rect 37327 4659 37347 4679
rect 37444 4659 37464 4679
rect 37540 4659 37560 4679
rect 37652 4659 37672 4679
rect 37748 4659 37768 4679
rect 37858 4659 37878 4679
rect 37954 4659 37974 4679
rect 31586 4492 31606 4512
rect 39033 4489 39053 4509
rect 39129 4489 39149 4509
rect 39239 4489 39259 4509
rect 39335 4489 39355 4509
rect 39447 4489 39467 4509
rect 39543 4489 39563 4509
rect 39660 4489 39680 4509
rect 39756 4489 39776 4509
rect 41571 4486 41591 4506
rect 41667 4486 41687 4506
rect 41777 4486 41797 4506
rect 41873 4486 41893 4506
rect 41985 4486 42005 4506
rect 42081 4486 42101 4506
rect 42198 4486 42218 4506
rect 42294 4486 42314 4506
rect 900 3986 920 4006
rect 996 3986 1016 4006
rect 1113 3986 1133 4006
rect 1209 3986 1229 4006
rect 1321 3986 1341 4006
rect 1417 3986 1437 4006
rect 1527 3986 1547 4006
rect 1623 3986 1643 4006
rect 3395 3981 3415 4001
rect 3491 3981 3511 4001
rect 3608 3981 3628 4001
rect 3704 3981 3724 4001
rect 3816 3981 3836 4001
rect 3912 3981 3932 4001
rect 4022 3981 4042 4001
rect 4118 3981 4138 4001
rect 11608 3980 11628 4000
rect 8142 3819 8162 3839
rect 8238 3819 8258 3839
rect 8348 3819 8368 3839
rect 8444 3819 8464 3839
rect 8556 3819 8576 3839
rect 8652 3819 8672 3839
rect 8769 3819 8789 3839
rect 11704 3980 11724 4000
rect 11821 3980 11841 4000
rect 11917 3980 11937 4000
rect 12029 3980 12049 4000
rect 12125 3980 12145 4000
rect 12235 3980 12255 4000
rect 12331 3980 12351 4000
rect 14103 3975 14123 3995
rect 8865 3819 8885 3839
rect 9190 3815 9210 3835
rect 9286 3815 9306 3835
rect 9396 3815 9416 3835
rect 9492 3815 9512 3835
rect 9604 3815 9624 3835
rect 9700 3815 9720 3835
rect 9817 3815 9837 3835
rect 9913 3815 9933 3835
rect 14199 3975 14219 3995
rect 14316 3975 14336 3995
rect 14412 3975 14432 3995
rect 14524 3975 14544 3995
rect 14620 3975 14640 3995
rect 14730 3975 14750 3995
rect 14826 3975 14846 3995
rect 22573 3984 22593 4004
rect 18850 3813 18870 3833
rect 18946 3813 18966 3833
rect 19056 3813 19076 3833
rect 19152 3813 19172 3833
rect 19264 3813 19284 3833
rect 19360 3813 19380 3833
rect 19477 3813 19497 3833
rect 22669 3984 22689 4004
rect 22786 3984 22806 4004
rect 22882 3984 22902 4004
rect 22994 3984 23014 4004
rect 23090 3984 23110 4004
rect 23200 3984 23220 4004
rect 23296 3984 23316 4004
rect 25068 3979 25088 3999
rect 19573 3813 19593 3833
rect 19898 3809 19918 3829
rect 19994 3809 20014 3829
rect 20104 3809 20124 3829
rect 20200 3809 20220 3829
rect 20312 3809 20332 3829
rect 20408 3809 20428 3829
rect 20525 3809 20545 3829
rect 20621 3809 20641 3829
rect 25164 3979 25184 3999
rect 25281 3979 25301 3999
rect 25377 3979 25397 3999
rect 25489 3979 25509 3999
rect 25585 3979 25605 3999
rect 25695 3979 25715 3999
rect 25791 3979 25811 3999
rect 33281 3978 33301 3998
rect 29815 3817 29835 3837
rect 29911 3817 29931 3837
rect 30021 3817 30041 3837
rect 30117 3817 30137 3837
rect 30229 3817 30249 3837
rect 30325 3817 30345 3837
rect 30442 3817 30462 3837
rect 33377 3978 33397 3998
rect 33494 3978 33514 3998
rect 33590 3978 33610 3998
rect 33702 3978 33722 3998
rect 33798 3978 33818 3998
rect 33908 3978 33928 3998
rect 34004 3978 34024 3998
rect 35776 3973 35796 3993
rect 30538 3817 30558 3837
rect 30863 3813 30883 3833
rect 30959 3813 30979 3833
rect 31069 3813 31089 3833
rect 31165 3813 31185 3833
rect 31277 3813 31297 3833
rect 31373 3813 31393 3833
rect 31490 3813 31510 3833
rect 31586 3813 31606 3833
rect 35872 3973 35892 3993
rect 35989 3973 36009 3993
rect 36085 3973 36105 3993
rect 36197 3973 36217 3993
rect 36293 3973 36313 3993
rect 36403 3973 36423 3993
rect 36499 3973 36519 3993
rect 40523 3811 40543 3831
rect 40619 3811 40639 3831
rect 40729 3811 40749 3831
rect 40825 3811 40845 3831
rect 40937 3811 40957 3831
rect 41033 3811 41053 3831
rect 41150 3811 41170 3831
rect 41246 3811 41266 3831
rect 41571 3807 41591 3827
rect 41667 3807 41687 3827
rect 41777 3807 41797 3827
rect 41873 3807 41893 3827
rect 41985 3807 42005 3827
rect 42081 3807 42101 3827
rect 42198 3807 42218 3827
rect 42294 3807 42314 3827
rect 900 3218 920 3238
rect 996 3218 1016 3238
rect 1113 3218 1133 3238
rect 1209 3218 1229 3238
rect 1321 3218 1341 3238
rect 1417 3218 1437 3238
rect 1527 3218 1547 3238
rect 1623 3218 1643 3238
rect 1948 3214 1968 3234
rect 2044 3214 2064 3234
rect 2161 3214 2181 3234
rect 2257 3214 2277 3234
rect 2369 3214 2389 3234
rect 2465 3214 2485 3234
rect 2575 3214 2595 3234
rect 2671 3214 2691 3234
rect 6695 3052 6715 3072
rect 6791 3052 6811 3072
rect 6901 3052 6921 3072
rect 6997 3052 7017 3072
rect 7109 3052 7129 3072
rect 7205 3052 7225 3072
rect 7322 3052 7342 3072
rect 11608 3212 11628 3232
rect 11704 3212 11724 3232
rect 11821 3212 11841 3232
rect 11917 3212 11937 3232
rect 12029 3212 12049 3232
rect 12125 3212 12145 3232
rect 12235 3212 12255 3232
rect 12331 3212 12351 3232
rect 12656 3208 12676 3228
rect 7418 3052 7438 3072
rect 9190 3047 9210 3067
rect 9286 3047 9306 3067
rect 9396 3047 9416 3067
rect 9492 3047 9512 3067
rect 9604 3047 9624 3067
rect 9700 3047 9720 3067
rect 9817 3047 9837 3067
rect 12752 3208 12772 3228
rect 12869 3208 12889 3228
rect 12965 3208 12985 3228
rect 13077 3208 13097 3228
rect 13173 3208 13193 3228
rect 13283 3208 13303 3228
rect 13379 3208 13399 3228
rect 9913 3047 9933 3067
rect 17403 3046 17423 3066
rect 17499 3046 17519 3066
rect 17609 3046 17629 3066
rect 17705 3046 17725 3066
rect 17817 3046 17837 3066
rect 17913 3046 17933 3066
rect 18030 3046 18050 3066
rect 22573 3216 22593 3236
rect 22669 3216 22689 3236
rect 22786 3216 22806 3236
rect 22882 3216 22902 3236
rect 22994 3216 23014 3236
rect 23090 3216 23110 3236
rect 23200 3216 23220 3236
rect 23296 3216 23316 3236
rect 23621 3212 23641 3232
rect 18126 3046 18146 3066
rect 19898 3041 19918 3061
rect 19994 3041 20014 3061
rect 20104 3041 20124 3061
rect 20200 3041 20220 3061
rect 20312 3041 20332 3061
rect 20408 3041 20428 3061
rect 20525 3041 20545 3061
rect 23717 3212 23737 3232
rect 23834 3212 23854 3232
rect 23930 3212 23950 3232
rect 24042 3212 24062 3232
rect 24138 3212 24158 3232
rect 24248 3212 24268 3232
rect 24344 3212 24364 3232
rect 20621 3041 20641 3061
rect 28368 3050 28388 3070
rect 28464 3050 28484 3070
rect 28574 3050 28594 3070
rect 28670 3050 28690 3070
rect 28782 3050 28802 3070
rect 28878 3050 28898 3070
rect 28995 3050 29015 3070
rect 33281 3210 33301 3230
rect 33377 3210 33397 3230
rect 33494 3210 33514 3230
rect 33590 3210 33610 3230
rect 33702 3210 33722 3230
rect 33798 3210 33818 3230
rect 33908 3210 33928 3230
rect 34004 3210 34024 3230
rect 34329 3206 34349 3226
rect 29091 3050 29111 3070
rect 30863 3045 30883 3065
rect 30959 3045 30979 3065
rect 31069 3045 31089 3065
rect 31165 3045 31185 3065
rect 31277 3045 31297 3065
rect 31373 3045 31393 3065
rect 31490 3045 31510 3065
rect 34425 3206 34445 3226
rect 34542 3206 34562 3226
rect 34638 3206 34658 3226
rect 34750 3206 34770 3226
rect 34846 3206 34866 3226
rect 34956 3206 34976 3226
rect 35052 3206 35072 3226
rect 31586 3045 31606 3065
rect 39076 3044 39096 3064
rect 39172 3044 39192 3064
rect 39282 3044 39302 3064
rect 39378 3044 39398 3064
rect 39490 3044 39510 3064
rect 39586 3044 39606 3064
rect 39703 3044 39723 3064
rect 39799 3044 39819 3064
rect 41571 3039 41591 3059
rect 41667 3039 41687 3059
rect 41777 3039 41797 3059
rect 41873 3039 41893 3059
rect 41985 3039 42005 3059
rect 42081 3039 42101 3059
rect 42198 3039 42218 3059
rect 42294 3039 42314 3059
rect 900 2539 920 2559
rect 996 2539 1016 2559
rect 1113 2539 1133 2559
rect 1209 2539 1229 2559
rect 1321 2539 1341 2559
rect 1417 2539 1437 2559
rect 1527 2539 1547 2559
rect 1623 2539 1643 2559
rect 11608 2533 11628 2553
rect 8142 2372 8162 2392
rect 8238 2372 8258 2392
rect 8348 2372 8368 2392
rect 8444 2372 8464 2392
rect 8556 2372 8576 2392
rect 8652 2372 8672 2392
rect 8769 2372 8789 2392
rect 11704 2533 11724 2553
rect 11821 2533 11841 2553
rect 11917 2533 11937 2553
rect 12029 2533 12049 2553
rect 12125 2533 12145 2553
rect 12235 2533 12255 2553
rect 12331 2533 12351 2553
rect 8865 2372 8885 2392
rect 9190 2368 9210 2388
rect 9286 2368 9306 2388
rect 9396 2368 9416 2388
rect 9492 2368 9512 2388
rect 9604 2368 9624 2388
rect 9700 2368 9720 2388
rect 9817 2368 9837 2388
rect 9913 2368 9933 2388
rect 22573 2537 22593 2557
rect 18850 2366 18870 2386
rect 18946 2366 18966 2386
rect 19056 2366 19076 2386
rect 19152 2366 19172 2386
rect 19264 2366 19284 2386
rect 19360 2366 19380 2386
rect 19477 2366 19497 2386
rect 22669 2537 22689 2557
rect 22786 2537 22806 2557
rect 22882 2537 22902 2557
rect 22994 2537 23014 2557
rect 23090 2537 23110 2557
rect 23200 2537 23220 2557
rect 23296 2537 23316 2557
rect 19573 2366 19593 2386
rect 19898 2362 19918 2382
rect 19994 2362 20014 2382
rect 20104 2362 20124 2382
rect 20200 2362 20220 2382
rect 20312 2362 20332 2382
rect 20408 2362 20428 2382
rect 20525 2362 20545 2382
rect 20621 2362 20641 2382
rect 33281 2531 33301 2551
rect 29815 2370 29835 2390
rect 29911 2370 29931 2390
rect 30021 2370 30041 2390
rect 30117 2370 30137 2390
rect 30229 2370 30249 2390
rect 30325 2370 30345 2390
rect 30442 2370 30462 2390
rect 33377 2531 33397 2551
rect 33494 2531 33514 2551
rect 33590 2531 33610 2551
rect 33702 2531 33722 2551
rect 33798 2531 33818 2551
rect 33908 2531 33928 2551
rect 34004 2531 34024 2551
rect 30538 2370 30558 2390
rect 30863 2366 30883 2386
rect 30959 2366 30979 2386
rect 31069 2366 31089 2386
rect 31165 2366 31185 2386
rect 31277 2366 31297 2386
rect 31373 2366 31393 2386
rect 31490 2366 31510 2386
rect 31586 2366 31606 2386
rect 40523 2364 40543 2384
rect 40619 2364 40639 2384
rect 40729 2364 40749 2384
rect 40825 2364 40845 2384
rect 40937 2364 40957 2384
rect 41033 2364 41053 2384
rect 41150 2364 41170 2384
rect 41246 2364 41266 2384
rect 41571 2360 41591 2380
rect 41667 2360 41687 2380
rect 41777 2360 41797 2380
rect 41873 2360 41893 2380
rect 41985 2360 42005 2380
rect 42081 2360 42101 2380
rect 42198 2360 42218 2380
rect 42294 2360 42314 2380
rect 10611 380 10631 400
rect 10707 380 10727 400
rect 10824 380 10844 400
rect 10920 380 10940 400
rect 11032 380 11052 400
rect 11128 380 11148 400
rect 11238 380 11258 400
rect 11334 380 11354 400
rect 21248 367 21268 387
rect 21344 367 21364 387
rect 21461 367 21481 387
rect 21557 367 21577 387
rect 21669 367 21689 387
rect 21765 367 21785 387
rect 21875 367 21895 387
rect 21971 367 21991 387
rect 32284 378 32304 398
rect 32380 378 32400 398
rect 32497 378 32517 398
rect 32593 378 32613 398
rect 32705 378 32725 398
rect 32801 378 32821 398
rect 32911 378 32931 398
rect 33007 378 33027 398
<< psubdiff >>
rect 9755 13735 9866 13746
rect 9755 13705 9797 13735
rect 9825 13705 9866 13735
rect 20463 13729 20574 13744
rect 9755 13691 9866 13705
rect 20463 13699 20505 13729
rect 20533 13699 20574 13729
rect 31428 13733 31539 13744
rect 969 13424 1080 13438
rect 969 13394 1010 13424
rect 1038 13394 1080 13424
rect 969 13379 1080 13394
rect 2017 13420 2128 13434
rect 20463 13685 20574 13699
rect 31428 13703 31470 13733
rect 31498 13703 31539 13733
rect 42136 13727 42247 13742
rect 2017 13390 2058 13420
rect 2086 13390 2128 13420
rect 11677 13418 11788 13432
rect 2017 13375 2128 13390
rect 11677 13388 11718 13418
rect 11746 13388 11788 13418
rect 11677 13373 11788 13388
rect 12725 13414 12836 13428
rect 31428 13689 31539 13703
rect 42136 13697 42178 13727
rect 42206 13697 42247 13727
rect 12725 13384 12766 13414
rect 12794 13384 12836 13414
rect 22642 13422 22753 13436
rect 12725 13369 12836 13384
rect 22642 13392 22683 13422
rect 22711 13392 22753 13422
rect 22642 13377 22753 13392
rect 23690 13418 23801 13432
rect 42136 13683 42247 13697
rect 23690 13388 23731 13418
rect 23759 13388 23801 13418
rect 33350 13416 33461 13430
rect 23690 13373 23801 13388
rect 33350 13386 33391 13416
rect 33419 13386 33461 13416
rect 33350 13371 33461 13386
rect 34398 13412 34509 13426
rect 34398 13382 34439 13412
rect 34467 13382 34509 13412
rect 34398 13367 34509 13382
rect 8707 13060 8818 13075
rect 8707 13030 8749 13060
rect 8777 13030 8818 13060
rect 8707 13016 8818 13030
rect 9755 13056 9866 13071
rect 9755 13026 9797 13056
rect 9825 13026 9866 13056
rect 19415 13054 19526 13069
rect 9755 13012 9866 13026
rect 19415 13024 19457 13054
rect 19485 13024 19526 13054
rect 969 12745 1080 12759
rect 19415 13010 19526 13024
rect 20463 13050 20574 13065
rect 20463 13020 20505 13050
rect 20533 13020 20574 13050
rect 30380 13058 30491 13073
rect 969 12715 1010 12745
rect 1038 12715 1080 12745
rect 969 12702 1080 12715
rect 3464 12740 3575 12754
rect 20463 13006 20574 13020
rect 30380 13028 30422 13058
rect 30450 13028 30491 13058
rect 3464 12710 3505 12740
rect 3533 12710 3575 12740
rect 11677 12739 11788 12753
rect 30380 13014 30491 13028
rect 31428 13054 31539 13069
rect 31428 13024 31470 13054
rect 31498 13024 31539 13054
rect 41088 13052 41199 13067
rect 3464 12695 3575 12710
rect 11677 12709 11718 12739
rect 11746 12709 11788 12739
rect 11677 12696 11788 12709
rect 14172 12734 14283 12748
rect 31428 13010 31539 13024
rect 41088 13022 41130 13052
rect 41158 13022 41199 13052
rect 14172 12704 14213 12734
rect 14241 12704 14283 12734
rect 22642 12743 22753 12757
rect 41088 13008 41199 13022
rect 42136 13048 42247 13063
rect 42136 13018 42178 13048
rect 42206 13018 42247 13048
rect 14172 12689 14283 12704
rect 22642 12713 22683 12743
rect 22711 12713 22753 12743
rect 22642 12700 22753 12713
rect 25137 12738 25248 12752
rect 42136 13004 42247 13018
rect 25137 12708 25178 12738
rect 25206 12708 25248 12738
rect 33350 12737 33461 12751
rect 25137 12693 25248 12708
rect 33350 12707 33391 12737
rect 33419 12707 33461 12737
rect 33350 12694 33461 12707
rect 35845 12732 35956 12746
rect 35845 12702 35886 12732
rect 35914 12702 35956 12732
rect 35845 12687 35956 12702
rect 7260 12293 7371 12308
rect 7260 12263 7302 12293
rect 7330 12263 7371 12293
rect 7260 12249 7371 12263
rect 9755 12288 9866 12301
rect 9755 12258 9797 12288
rect 9825 12258 9866 12288
rect 17968 12287 18079 12302
rect 9755 12244 9866 12258
rect 17968 12257 18010 12287
rect 18038 12257 18079 12287
rect 969 11977 1080 11991
rect 17968 12243 18079 12257
rect 20463 12282 20574 12295
rect 20463 12252 20505 12282
rect 20533 12252 20574 12282
rect 28933 12291 29044 12306
rect 969 11947 1010 11977
rect 1038 11947 1080 11977
rect 969 11932 1080 11947
rect 2017 11973 2128 11987
rect 20463 12238 20574 12252
rect 28933 12261 28975 12291
rect 29003 12261 29044 12291
rect 2017 11943 2058 11973
rect 2086 11943 2128 11973
rect 11677 11971 11788 11985
rect 28933 12247 29044 12261
rect 31428 12286 31539 12299
rect 31428 12256 31470 12286
rect 31498 12256 31539 12286
rect 39641 12285 39752 12300
rect 2017 11928 2128 11943
rect 11677 11941 11718 11971
rect 11746 11941 11788 11971
rect 11677 11926 11788 11941
rect 12725 11967 12836 11981
rect 31428 12242 31539 12256
rect 39641 12255 39683 12285
rect 39711 12255 39752 12285
rect 12725 11937 12766 11967
rect 12794 11937 12836 11967
rect 22642 11975 22753 11989
rect 39641 12241 39752 12255
rect 42136 12280 42247 12293
rect 42136 12250 42178 12280
rect 42206 12250 42247 12280
rect 12725 11922 12836 11937
rect 22642 11945 22683 11975
rect 22711 11945 22753 11975
rect 22642 11930 22753 11945
rect 23690 11971 23801 11985
rect 42136 12236 42247 12250
rect 23690 11941 23731 11971
rect 23759 11941 23801 11971
rect 33350 11969 33461 11983
rect 23690 11926 23801 11941
rect 33350 11939 33391 11969
rect 33419 11939 33461 11969
rect 33350 11924 33461 11939
rect 34398 11965 34509 11979
rect 34398 11935 34439 11965
rect 34467 11935 34509 11965
rect 34398 11920 34509 11935
rect 8707 11613 8818 11628
rect 8707 11583 8749 11613
rect 8777 11583 8818 11613
rect 8707 11569 8818 11583
rect 9755 11609 9866 11624
rect 9755 11579 9797 11609
rect 9825 11579 9866 11609
rect 19415 11607 19526 11622
rect 9755 11565 9866 11579
rect 19415 11577 19457 11607
rect 19485 11577 19526 11607
rect 969 11298 1080 11312
rect 19415 11563 19526 11577
rect 20463 11603 20574 11618
rect 20463 11573 20505 11603
rect 20533 11573 20574 11603
rect 30380 11611 30491 11626
rect 969 11268 1010 11298
rect 1038 11268 1080 11298
rect 969 11253 1080 11268
rect 3507 11295 3618 11309
rect 20463 11559 20574 11573
rect 30380 11581 30422 11611
rect 30450 11581 30491 11611
rect 3507 11265 3548 11295
rect 3576 11265 3618 11295
rect 11677 11292 11788 11306
rect 30380 11567 30491 11581
rect 31428 11607 31539 11622
rect 31428 11577 31470 11607
rect 31498 11577 31539 11607
rect 41088 11605 41199 11620
rect 3507 11250 3618 11265
rect 11677 11262 11718 11292
rect 11746 11262 11788 11292
rect 11677 11247 11788 11262
rect 14215 11289 14326 11303
rect 31428 11563 31539 11577
rect 41088 11575 41130 11605
rect 41158 11575 41199 11605
rect 14215 11259 14256 11289
rect 14284 11259 14326 11289
rect 22642 11296 22753 11310
rect 41088 11561 41199 11575
rect 42136 11601 42247 11616
rect 42136 11571 42178 11601
rect 42206 11571 42247 11601
rect 14215 11244 14326 11259
rect 22642 11266 22683 11296
rect 22711 11266 22753 11296
rect 22642 11251 22753 11266
rect 25180 11293 25291 11307
rect 42136 11557 42247 11571
rect 25180 11263 25221 11293
rect 25249 11263 25291 11293
rect 33350 11290 33461 11304
rect 25180 11248 25291 11263
rect 33350 11260 33391 11290
rect 33419 11260 33461 11290
rect 33350 11245 33461 11260
rect 35888 11287 35999 11301
rect 35888 11257 35929 11287
rect 35957 11257 35999 11287
rect 35888 11242 35999 11257
rect 7218 10771 7329 10786
rect 7218 10741 7260 10771
rect 7288 10741 7329 10771
rect 7218 10727 7329 10741
rect 9756 10768 9867 10783
rect 9756 10738 9798 10768
rect 9826 10738 9867 10768
rect 17926 10765 18037 10780
rect 9756 10724 9867 10738
rect 17926 10735 17968 10765
rect 17996 10735 18037 10765
rect 970 10457 1081 10471
rect 17926 10721 18037 10735
rect 20464 10762 20575 10777
rect 20464 10732 20506 10762
rect 20534 10732 20575 10762
rect 28891 10769 29002 10784
rect 970 10427 1011 10457
rect 1039 10427 1081 10457
rect 970 10412 1081 10427
rect 2018 10453 2129 10467
rect 20464 10718 20575 10732
rect 28891 10739 28933 10769
rect 28961 10739 29002 10769
rect 2018 10423 2059 10453
rect 2087 10423 2129 10453
rect 11678 10451 11789 10465
rect 28891 10725 29002 10739
rect 31429 10766 31540 10781
rect 31429 10736 31471 10766
rect 31499 10736 31540 10766
rect 39599 10763 39710 10778
rect 2018 10408 2129 10423
rect 11678 10421 11719 10451
rect 11747 10421 11789 10451
rect 11678 10406 11789 10421
rect 12726 10447 12837 10461
rect 31429 10722 31540 10736
rect 39599 10733 39641 10763
rect 39669 10733 39710 10763
rect 12726 10417 12767 10447
rect 12795 10417 12837 10447
rect 22643 10455 22754 10469
rect 39599 10719 39710 10733
rect 42137 10760 42248 10775
rect 42137 10730 42179 10760
rect 42207 10730 42248 10760
rect 12726 10402 12837 10417
rect 22643 10425 22684 10455
rect 22712 10425 22754 10455
rect 22643 10410 22754 10425
rect 23691 10451 23802 10465
rect 42137 10716 42248 10730
rect 23691 10421 23732 10451
rect 23760 10421 23802 10451
rect 33351 10449 33462 10463
rect 23691 10406 23802 10421
rect 33351 10419 33392 10449
rect 33420 10419 33462 10449
rect 33351 10404 33462 10419
rect 34399 10445 34510 10459
rect 34399 10415 34440 10445
rect 34468 10415 34510 10445
rect 34399 10400 34510 10415
rect 8708 10093 8819 10108
rect 8708 10063 8750 10093
rect 8778 10063 8819 10093
rect 8708 10049 8819 10063
rect 9756 10089 9867 10104
rect 9756 10059 9798 10089
rect 9826 10059 9867 10089
rect 19416 10087 19527 10102
rect 9756 10045 9867 10059
rect 19416 10057 19458 10087
rect 19486 10057 19527 10087
rect 970 9778 1081 9792
rect 19416 10043 19527 10057
rect 20464 10083 20575 10098
rect 20464 10053 20506 10083
rect 20534 10053 20575 10083
rect 30381 10091 30492 10106
rect 970 9748 1011 9778
rect 1039 9748 1081 9778
rect 970 9735 1081 9748
rect 3465 9773 3576 9787
rect 20464 10039 20575 10053
rect 30381 10061 30423 10091
rect 30451 10061 30492 10091
rect 3465 9743 3506 9773
rect 3534 9743 3576 9773
rect 11678 9772 11789 9786
rect 30381 10047 30492 10061
rect 31429 10087 31540 10102
rect 31429 10057 31471 10087
rect 31499 10057 31540 10087
rect 41089 10085 41200 10100
rect 3465 9728 3576 9743
rect 11678 9742 11719 9772
rect 11747 9742 11789 9772
rect 11678 9729 11789 9742
rect 14173 9767 14284 9781
rect 31429 10043 31540 10057
rect 41089 10055 41131 10085
rect 41159 10055 41200 10085
rect 14173 9737 14214 9767
rect 14242 9737 14284 9767
rect 22643 9776 22754 9790
rect 41089 10041 41200 10055
rect 42137 10081 42248 10096
rect 42137 10051 42179 10081
rect 42207 10051 42248 10081
rect 14173 9722 14284 9737
rect 22643 9746 22684 9776
rect 22712 9746 22754 9776
rect 22643 9733 22754 9746
rect 25138 9771 25249 9785
rect 42137 10037 42248 10051
rect 25138 9741 25179 9771
rect 25207 9741 25249 9771
rect 33351 9770 33462 9784
rect 25138 9726 25249 9741
rect 33351 9740 33392 9770
rect 33420 9740 33462 9770
rect 33351 9727 33462 9740
rect 35846 9765 35957 9779
rect 35846 9735 35887 9765
rect 35915 9735 35957 9765
rect 35846 9720 35957 9735
rect 7261 9326 7372 9341
rect 7261 9296 7303 9326
rect 7331 9296 7372 9326
rect 7261 9282 7372 9296
rect 9756 9321 9867 9334
rect 9756 9291 9798 9321
rect 9826 9291 9867 9321
rect 17969 9320 18080 9335
rect 9756 9277 9867 9291
rect 17969 9290 18011 9320
rect 18039 9290 18080 9320
rect 970 9010 1081 9024
rect 17969 9276 18080 9290
rect 20464 9315 20575 9328
rect 20464 9285 20506 9315
rect 20534 9285 20575 9315
rect 28934 9324 29045 9339
rect 970 8980 1011 9010
rect 1039 8980 1081 9010
rect 970 8965 1081 8980
rect 2018 9006 2129 9020
rect 20464 9271 20575 9285
rect 28934 9294 28976 9324
rect 29004 9294 29045 9324
rect 2018 8976 2059 9006
rect 2087 8976 2129 9006
rect 11678 9004 11789 9018
rect 28934 9280 29045 9294
rect 31429 9319 31540 9332
rect 31429 9289 31471 9319
rect 31499 9289 31540 9319
rect 39642 9318 39753 9333
rect 2018 8961 2129 8976
rect 11678 8974 11719 9004
rect 11747 8974 11789 9004
rect 11678 8959 11789 8974
rect 12726 9000 12837 9014
rect 31429 9275 31540 9289
rect 39642 9288 39684 9318
rect 39712 9288 39753 9318
rect 12726 8970 12767 9000
rect 12795 8970 12837 9000
rect 22643 9008 22754 9022
rect 39642 9274 39753 9288
rect 42137 9313 42248 9326
rect 42137 9283 42179 9313
rect 42207 9283 42248 9313
rect 12726 8955 12837 8970
rect 22643 8978 22684 9008
rect 22712 8978 22754 9008
rect 22643 8963 22754 8978
rect 23691 9004 23802 9018
rect 42137 9269 42248 9283
rect 23691 8974 23732 9004
rect 23760 8974 23802 9004
rect 33351 9002 33462 9016
rect 23691 8959 23802 8974
rect 33351 8972 33392 9002
rect 33420 8972 33462 9002
rect 33351 8957 33462 8972
rect 34399 8998 34510 9012
rect 34399 8968 34440 8998
rect 34468 8968 34510 8998
rect 34399 8953 34510 8968
rect 8708 8646 8819 8661
rect 8708 8616 8750 8646
rect 8778 8616 8819 8646
rect 8708 8602 8819 8616
rect 9756 8642 9867 8657
rect 9756 8612 9798 8642
rect 9826 8612 9867 8642
rect 19416 8640 19527 8655
rect 9756 8598 9867 8612
rect 19416 8610 19458 8640
rect 19486 8610 19527 8640
rect 970 8331 1081 8345
rect 19416 8596 19527 8610
rect 20464 8636 20575 8651
rect 20464 8606 20506 8636
rect 20534 8606 20575 8636
rect 30381 8644 30492 8659
rect 20464 8592 20575 8606
rect 30381 8614 30423 8644
rect 30451 8614 30492 8644
rect 970 8301 1011 8331
rect 1039 8301 1081 8331
rect 970 8286 1081 8301
rect 4573 8322 4684 8336
rect 11678 8325 11789 8339
rect 30381 8600 30492 8614
rect 31429 8640 31540 8655
rect 31429 8610 31471 8640
rect 31499 8610 31540 8640
rect 41089 8638 41200 8653
rect 31429 8596 31540 8610
rect 41089 8608 41131 8638
rect 41159 8608 41200 8638
rect 4573 8292 4614 8322
rect 4642 8292 4684 8322
rect 4573 8277 4684 8292
rect 11678 8295 11719 8325
rect 11747 8295 11789 8325
rect 11678 8280 11789 8295
rect 15281 8316 15392 8330
rect 22643 8329 22754 8343
rect 41089 8594 41200 8608
rect 42137 8634 42248 8649
rect 42137 8604 42179 8634
rect 42207 8604 42248 8634
rect 42137 8590 42248 8604
rect 15281 8286 15322 8316
rect 15350 8286 15392 8316
rect 15281 8271 15392 8286
rect 22643 8299 22684 8329
rect 22712 8299 22754 8329
rect 22643 8284 22754 8299
rect 26246 8320 26357 8334
rect 33351 8323 33462 8337
rect 26246 8290 26287 8320
rect 26315 8290 26357 8320
rect 26246 8275 26357 8290
rect 33351 8293 33392 8323
rect 33420 8293 33462 8323
rect 33351 8278 33462 8293
rect 36954 8314 37065 8328
rect 36954 8284 36995 8314
rect 37023 8284 37065 8314
rect 36954 8269 37065 8284
rect 6150 7736 6261 7751
rect 6150 7706 6192 7736
rect 6220 7706 6261 7736
rect 6150 7692 6261 7706
rect 9753 7727 9864 7742
rect 9753 7697 9795 7727
rect 9823 7697 9864 7727
rect 16858 7730 16969 7745
rect 16858 7700 16900 7730
rect 16928 7700 16969 7730
rect 9753 7683 9864 7697
rect 16858 7686 16969 7700
rect 20461 7721 20572 7736
rect 20461 7691 20503 7721
rect 20531 7691 20572 7721
rect 27823 7734 27934 7749
rect 27823 7704 27865 7734
rect 27893 7704 27934 7734
rect 967 7416 1078 7430
rect 967 7386 1008 7416
rect 1036 7386 1078 7416
rect 967 7371 1078 7386
rect 2015 7412 2126 7426
rect 20461 7677 20572 7691
rect 27823 7690 27934 7704
rect 31426 7725 31537 7740
rect 31426 7695 31468 7725
rect 31496 7695 31537 7725
rect 38531 7728 38642 7743
rect 38531 7698 38573 7728
rect 38601 7698 38642 7728
rect 2015 7382 2056 7412
rect 2084 7382 2126 7412
rect 11675 7410 11786 7424
rect 2015 7367 2126 7382
rect 11675 7380 11716 7410
rect 11744 7380 11786 7410
rect 11675 7365 11786 7380
rect 12723 7406 12834 7420
rect 31426 7681 31537 7695
rect 38531 7684 38642 7698
rect 42134 7719 42245 7734
rect 42134 7689 42176 7719
rect 42204 7689 42245 7719
rect 12723 7376 12764 7406
rect 12792 7376 12834 7406
rect 22640 7414 22751 7428
rect 12723 7361 12834 7376
rect 22640 7384 22681 7414
rect 22709 7384 22751 7414
rect 22640 7369 22751 7384
rect 23688 7410 23799 7424
rect 42134 7675 42245 7689
rect 23688 7380 23729 7410
rect 23757 7380 23799 7410
rect 33348 7408 33459 7422
rect 23688 7365 23799 7380
rect 33348 7378 33389 7408
rect 33417 7378 33459 7408
rect 33348 7363 33459 7378
rect 34396 7404 34507 7418
rect 34396 7374 34437 7404
rect 34465 7374 34507 7404
rect 34396 7359 34507 7374
rect 8705 7052 8816 7067
rect 8705 7022 8747 7052
rect 8775 7022 8816 7052
rect 8705 7008 8816 7022
rect 9753 7048 9864 7063
rect 9753 7018 9795 7048
rect 9823 7018 9864 7048
rect 19413 7046 19524 7061
rect 9753 7004 9864 7018
rect 19413 7016 19455 7046
rect 19483 7016 19524 7046
rect 967 6737 1078 6751
rect 19413 7002 19524 7016
rect 20461 7042 20572 7057
rect 20461 7012 20503 7042
rect 20531 7012 20572 7042
rect 30378 7050 30489 7065
rect 967 6707 1008 6737
rect 1036 6707 1078 6737
rect 967 6694 1078 6707
rect 3462 6732 3573 6746
rect 20461 6998 20572 7012
rect 30378 7020 30420 7050
rect 30448 7020 30489 7050
rect 3462 6702 3503 6732
rect 3531 6702 3573 6732
rect 11675 6731 11786 6745
rect 30378 7006 30489 7020
rect 31426 7046 31537 7061
rect 31426 7016 31468 7046
rect 31496 7016 31537 7046
rect 41086 7044 41197 7059
rect 3462 6687 3573 6702
rect 11675 6701 11716 6731
rect 11744 6701 11786 6731
rect 11675 6688 11786 6701
rect 14170 6726 14281 6740
rect 31426 7002 31537 7016
rect 41086 7014 41128 7044
rect 41156 7014 41197 7044
rect 14170 6696 14211 6726
rect 14239 6696 14281 6726
rect 22640 6735 22751 6749
rect 41086 7000 41197 7014
rect 42134 7040 42245 7055
rect 42134 7010 42176 7040
rect 42204 7010 42245 7040
rect 14170 6681 14281 6696
rect 22640 6705 22681 6735
rect 22709 6705 22751 6735
rect 22640 6692 22751 6705
rect 25135 6730 25246 6744
rect 42134 6996 42245 7010
rect 25135 6700 25176 6730
rect 25204 6700 25246 6730
rect 33348 6729 33459 6743
rect 25135 6685 25246 6700
rect 33348 6699 33389 6729
rect 33417 6699 33459 6729
rect 33348 6686 33459 6699
rect 35843 6724 35954 6738
rect 35843 6694 35884 6724
rect 35912 6694 35954 6724
rect 35843 6679 35954 6694
rect 7258 6285 7369 6300
rect 7258 6255 7300 6285
rect 7328 6255 7369 6285
rect 7258 6241 7369 6255
rect 9753 6280 9864 6293
rect 9753 6250 9795 6280
rect 9823 6250 9864 6280
rect 17966 6279 18077 6294
rect 9753 6236 9864 6250
rect 17966 6249 18008 6279
rect 18036 6249 18077 6279
rect 967 5969 1078 5983
rect 17966 6235 18077 6249
rect 20461 6274 20572 6287
rect 20461 6244 20503 6274
rect 20531 6244 20572 6274
rect 28931 6283 29042 6298
rect 967 5939 1008 5969
rect 1036 5939 1078 5969
rect 967 5924 1078 5939
rect 2015 5965 2126 5979
rect 20461 6230 20572 6244
rect 28931 6253 28973 6283
rect 29001 6253 29042 6283
rect 2015 5935 2056 5965
rect 2084 5935 2126 5965
rect 11675 5963 11786 5977
rect 28931 6239 29042 6253
rect 31426 6278 31537 6291
rect 31426 6248 31468 6278
rect 31496 6248 31537 6278
rect 39639 6277 39750 6292
rect 2015 5920 2126 5935
rect 11675 5933 11716 5963
rect 11744 5933 11786 5963
rect 11675 5918 11786 5933
rect 12723 5959 12834 5973
rect 31426 6234 31537 6248
rect 39639 6247 39681 6277
rect 39709 6247 39750 6277
rect 12723 5929 12764 5959
rect 12792 5929 12834 5959
rect 22640 5967 22751 5981
rect 39639 6233 39750 6247
rect 42134 6272 42245 6285
rect 42134 6242 42176 6272
rect 42204 6242 42245 6272
rect 12723 5914 12834 5929
rect 22640 5937 22681 5967
rect 22709 5937 22751 5967
rect 22640 5922 22751 5937
rect 23688 5963 23799 5977
rect 42134 6228 42245 6242
rect 23688 5933 23729 5963
rect 23757 5933 23799 5963
rect 33348 5961 33459 5975
rect 23688 5918 23799 5933
rect 33348 5931 33389 5961
rect 33417 5931 33459 5961
rect 33348 5916 33459 5931
rect 34396 5957 34507 5971
rect 34396 5927 34437 5957
rect 34465 5927 34507 5957
rect 34396 5912 34507 5927
rect 8705 5605 8816 5620
rect 8705 5575 8747 5605
rect 8775 5575 8816 5605
rect 8705 5561 8816 5575
rect 9753 5601 9864 5616
rect 9753 5571 9795 5601
rect 9823 5571 9864 5601
rect 19413 5599 19524 5614
rect 9753 5557 9864 5571
rect 19413 5569 19455 5599
rect 19483 5569 19524 5599
rect 967 5290 1078 5304
rect 19413 5555 19524 5569
rect 20461 5595 20572 5610
rect 20461 5565 20503 5595
rect 20531 5565 20572 5595
rect 30378 5603 30489 5618
rect 967 5260 1008 5290
rect 1036 5260 1078 5290
rect 967 5245 1078 5260
rect 3505 5287 3616 5301
rect 20461 5551 20572 5565
rect 30378 5573 30420 5603
rect 30448 5573 30489 5603
rect 3505 5257 3546 5287
rect 3574 5257 3616 5287
rect 11675 5284 11786 5298
rect 30378 5559 30489 5573
rect 31426 5599 31537 5614
rect 31426 5569 31468 5599
rect 31496 5569 31537 5599
rect 41086 5597 41197 5612
rect 3505 5242 3616 5257
rect 11675 5254 11716 5284
rect 11744 5254 11786 5284
rect 11675 5239 11786 5254
rect 14213 5281 14324 5295
rect 31426 5555 31537 5569
rect 41086 5567 41128 5597
rect 41156 5567 41197 5597
rect 14213 5251 14254 5281
rect 14282 5251 14324 5281
rect 22640 5288 22751 5302
rect 41086 5553 41197 5567
rect 42134 5593 42245 5608
rect 42134 5563 42176 5593
rect 42204 5563 42245 5593
rect 14213 5236 14324 5251
rect 22640 5258 22681 5288
rect 22709 5258 22751 5288
rect 22640 5243 22751 5258
rect 25178 5285 25289 5299
rect 42134 5549 42245 5563
rect 25178 5255 25219 5285
rect 25247 5255 25289 5285
rect 33348 5282 33459 5296
rect 25178 5240 25289 5255
rect 33348 5252 33389 5282
rect 33417 5252 33459 5282
rect 33348 5237 33459 5252
rect 35886 5279 35997 5293
rect 35886 5249 35927 5279
rect 35955 5249 35997 5279
rect 35886 5234 35997 5249
rect 7216 4763 7327 4778
rect 7216 4733 7258 4763
rect 7286 4733 7327 4763
rect 7216 4719 7327 4733
rect 9754 4760 9865 4775
rect 9754 4730 9796 4760
rect 9824 4730 9865 4760
rect 17924 4757 18035 4772
rect 9754 4716 9865 4730
rect 968 4449 1079 4463
rect 968 4419 1009 4449
rect 1037 4419 1079 4449
rect 968 4404 1079 4419
rect 2016 4445 2127 4459
rect 2016 4415 2057 4445
rect 2085 4415 2127 4445
rect 2016 4400 2127 4415
rect 4918 4451 5029 4465
rect 17924 4727 17966 4757
rect 17994 4727 18035 4757
rect 4918 4421 4959 4451
rect 4987 4421 5029 4451
rect 17924 4713 18035 4727
rect 20462 4754 20573 4769
rect 20462 4724 20504 4754
rect 20532 4724 20573 4754
rect 28889 4761 29000 4776
rect 20462 4710 20573 4724
rect 11676 4443 11787 4457
rect 4918 4406 5029 4421
rect 11676 4413 11717 4443
rect 11745 4413 11787 4443
rect 11676 4398 11787 4413
rect 12724 4439 12835 4453
rect 12724 4409 12765 4439
rect 12793 4409 12835 4439
rect 12724 4394 12835 4409
rect 15626 4445 15737 4459
rect 28889 4731 28931 4761
rect 28959 4731 29000 4761
rect 15626 4415 15667 4445
rect 15695 4415 15737 4445
rect 28889 4717 29000 4731
rect 31427 4758 31538 4773
rect 31427 4728 31469 4758
rect 31497 4728 31538 4758
rect 39597 4755 39708 4770
rect 31427 4714 31538 4728
rect 22641 4447 22752 4461
rect 15626 4400 15737 4415
rect 22641 4417 22682 4447
rect 22710 4417 22752 4447
rect 22641 4402 22752 4417
rect 23689 4443 23800 4457
rect 23689 4413 23730 4443
rect 23758 4413 23800 4443
rect 23689 4398 23800 4413
rect 26591 4449 26702 4463
rect 39597 4725 39639 4755
rect 39667 4725 39708 4755
rect 26591 4419 26632 4449
rect 26660 4419 26702 4449
rect 39597 4711 39708 4725
rect 42135 4752 42246 4767
rect 42135 4722 42177 4752
rect 42205 4722 42246 4752
rect 42135 4708 42246 4722
rect 33349 4441 33460 4455
rect 26591 4404 26702 4419
rect 33349 4411 33390 4441
rect 33418 4411 33460 4441
rect 33349 4396 33460 4411
rect 34397 4437 34508 4451
rect 34397 4407 34438 4437
rect 34466 4407 34508 4437
rect 34397 4392 34508 4407
rect 37299 4443 37410 4457
rect 37299 4413 37340 4443
rect 37368 4413 37410 4443
rect 37299 4398 37410 4413
rect 8706 4085 8817 4100
rect 8706 4055 8748 4085
rect 8776 4055 8817 4085
rect 8706 4041 8817 4055
rect 9754 4081 9865 4096
rect 9754 4051 9796 4081
rect 9824 4051 9865 4081
rect 19414 4079 19525 4094
rect 9754 4037 9865 4051
rect 19414 4049 19456 4079
rect 19484 4049 19525 4079
rect 968 3770 1079 3784
rect 19414 4035 19525 4049
rect 20462 4075 20573 4090
rect 20462 4045 20504 4075
rect 20532 4045 20573 4075
rect 30379 4083 30490 4098
rect 968 3740 1009 3770
rect 1037 3740 1079 3770
rect 968 3727 1079 3740
rect 3463 3765 3574 3779
rect 20462 4031 20573 4045
rect 30379 4053 30421 4083
rect 30449 4053 30490 4083
rect 3463 3735 3504 3765
rect 3532 3735 3574 3765
rect 11676 3764 11787 3778
rect 30379 4039 30490 4053
rect 31427 4079 31538 4094
rect 31427 4049 31469 4079
rect 31497 4049 31538 4079
rect 41087 4077 41198 4092
rect 3463 3720 3574 3735
rect 11676 3734 11717 3764
rect 11745 3734 11787 3764
rect 11676 3721 11787 3734
rect 14171 3759 14282 3773
rect 31427 4035 31538 4049
rect 41087 4047 41129 4077
rect 41157 4047 41198 4077
rect 14171 3729 14212 3759
rect 14240 3729 14282 3759
rect 22641 3768 22752 3782
rect 41087 4033 41198 4047
rect 42135 4073 42246 4088
rect 42135 4043 42177 4073
rect 42205 4043 42246 4073
rect 14171 3714 14282 3729
rect 22641 3738 22682 3768
rect 22710 3738 22752 3768
rect 22641 3725 22752 3738
rect 25136 3763 25247 3777
rect 42135 4029 42246 4043
rect 25136 3733 25177 3763
rect 25205 3733 25247 3763
rect 33349 3762 33460 3776
rect 25136 3718 25247 3733
rect 33349 3732 33390 3762
rect 33418 3732 33460 3762
rect 33349 3719 33460 3732
rect 35844 3757 35955 3771
rect 35844 3727 35885 3757
rect 35913 3727 35955 3757
rect 35844 3712 35955 3727
rect 7259 3318 7370 3333
rect 7259 3288 7301 3318
rect 7329 3288 7370 3318
rect 7259 3274 7370 3288
rect 9754 3313 9865 3326
rect 9754 3283 9796 3313
rect 9824 3283 9865 3313
rect 17967 3312 18078 3327
rect 9754 3269 9865 3283
rect 17967 3282 18009 3312
rect 18037 3282 18078 3312
rect 968 3002 1079 3016
rect 17967 3268 18078 3282
rect 20462 3307 20573 3320
rect 20462 3277 20504 3307
rect 20532 3277 20573 3307
rect 28932 3316 29043 3331
rect 968 2972 1009 3002
rect 1037 2972 1079 3002
rect 968 2957 1079 2972
rect 2016 2998 2127 3012
rect 20462 3263 20573 3277
rect 28932 3286 28974 3316
rect 29002 3286 29043 3316
rect 2016 2968 2057 2998
rect 2085 2968 2127 2998
rect 11676 2996 11787 3010
rect 28932 3272 29043 3286
rect 31427 3311 31538 3324
rect 31427 3281 31469 3311
rect 31497 3281 31538 3311
rect 39640 3310 39751 3325
rect 2016 2953 2127 2968
rect 11676 2966 11717 2996
rect 11745 2966 11787 2996
rect 11676 2951 11787 2966
rect 12724 2992 12835 3006
rect 31427 3267 31538 3281
rect 39640 3280 39682 3310
rect 39710 3280 39751 3310
rect 12724 2962 12765 2992
rect 12793 2962 12835 2992
rect 22641 3000 22752 3014
rect 39640 3266 39751 3280
rect 42135 3305 42246 3318
rect 42135 3275 42177 3305
rect 42205 3275 42246 3305
rect 12724 2947 12835 2962
rect 22641 2970 22682 3000
rect 22710 2970 22752 3000
rect 22641 2955 22752 2970
rect 23689 2996 23800 3010
rect 42135 3261 42246 3275
rect 23689 2966 23730 2996
rect 23758 2966 23800 2996
rect 33349 2994 33460 3008
rect 23689 2951 23800 2966
rect 33349 2964 33390 2994
rect 33418 2964 33460 2994
rect 33349 2949 33460 2964
rect 34397 2990 34508 3004
rect 34397 2960 34438 2990
rect 34466 2960 34508 2990
rect 34397 2945 34508 2960
rect 8706 2638 8817 2653
rect 8706 2608 8748 2638
rect 8776 2608 8817 2638
rect 8706 2594 8817 2608
rect 9754 2634 9865 2649
rect 9754 2604 9796 2634
rect 9824 2604 9865 2634
rect 19414 2632 19525 2647
rect 9754 2590 9865 2604
rect 19414 2602 19456 2632
rect 19484 2602 19525 2632
rect 968 2323 1079 2337
rect 19414 2588 19525 2602
rect 20462 2628 20573 2643
rect 20462 2598 20504 2628
rect 20532 2598 20573 2628
rect 30379 2636 30490 2651
rect 20462 2584 20573 2598
rect 30379 2606 30421 2636
rect 30449 2606 30490 2636
rect 968 2293 1009 2323
rect 1037 2293 1079 2323
rect 11676 2317 11787 2331
rect 30379 2592 30490 2606
rect 31427 2632 31538 2647
rect 31427 2602 31469 2632
rect 31497 2602 31538 2632
rect 41087 2630 41198 2645
rect 31427 2588 31538 2602
rect 41087 2600 41129 2630
rect 41157 2600 41198 2630
rect 968 2278 1079 2293
rect 11676 2287 11717 2317
rect 11745 2287 11787 2317
rect 22641 2321 22752 2335
rect 41087 2586 41198 2600
rect 42135 2626 42246 2641
rect 42135 2596 42177 2626
rect 42205 2596 42246 2626
rect 42135 2582 42246 2596
rect 11676 2272 11787 2287
rect 22641 2291 22682 2321
rect 22710 2291 22752 2321
rect 33349 2315 33460 2329
rect 22641 2276 22752 2291
rect 33349 2285 33390 2315
rect 33418 2285 33460 2315
rect 33349 2270 33460 2285
rect 10679 164 10790 178
rect 10679 134 10720 164
rect 10748 134 10790 164
rect 10679 119 10790 134
rect 21316 151 21427 165
rect 21316 121 21357 151
rect 21385 121 21427 151
rect 21316 106 21427 121
rect 32352 162 32463 176
rect 32352 132 32393 162
rect 32421 132 32463 162
rect 32352 117 32463 132
<< nsubdiff >>
rect 970 13771 1080 13785
rect 970 13741 1013 13771
rect 1041 13741 1080 13771
rect 970 13726 1080 13741
rect 2018 13767 2128 13781
rect 2018 13737 2061 13767
rect 2089 13737 2128 13767
rect 11678 13765 11788 13779
rect 2018 13722 2128 13737
rect 11678 13735 11721 13765
rect 11749 13735 11788 13765
rect 11678 13720 11788 13735
rect 12726 13761 12836 13775
rect 12726 13731 12769 13761
rect 12797 13731 12836 13761
rect 22643 13769 22753 13783
rect 12726 13716 12836 13731
rect 22643 13739 22686 13769
rect 22714 13739 22753 13769
rect 22643 13724 22753 13739
rect 23691 13765 23801 13779
rect 23691 13735 23734 13765
rect 23762 13735 23801 13765
rect 33351 13763 33461 13777
rect 23691 13720 23801 13735
rect 33351 13733 33394 13763
rect 33422 13733 33461 13763
rect 33351 13718 33461 13733
rect 34399 13759 34509 13773
rect 34399 13729 34442 13759
rect 34470 13729 34509 13759
rect 34399 13714 34509 13729
rect 9755 13388 9865 13403
rect 9755 13358 9794 13388
rect 9822 13358 9865 13388
rect 9755 13344 9865 13358
rect 20463 13382 20573 13397
rect 20463 13352 20502 13382
rect 20530 13352 20573 13382
rect 20463 13338 20573 13352
rect 31428 13386 31538 13401
rect 31428 13356 31467 13386
rect 31495 13356 31538 13386
rect 31428 13342 31538 13356
rect 42136 13380 42246 13395
rect 42136 13350 42175 13380
rect 42203 13350 42246 13380
rect 42136 13336 42246 13350
rect 970 13092 1080 13106
rect 970 13062 1013 13092
rect 1041 13062 1080 13092
rect 970 13047 1080 13062
rect 3465 13087 3575 13101
rect 3465 13057 3508 13087
rect 3536 13057 3575 13087
rect 3465 13042 3575 13057
rect 11678 13086 11788 13100
rect 11678 13056 11721 13086
rect 11749 13056 11788 13086
rect 11678 13041 11788 13056
rect 14173 13081 14283 13095
rect 14173 13051 14216 13081
rect 14244 13051 14283 13081
rect 14173 13036 14283 13051
rect 22643 13090 22753 13104
rect 22643 13060 22686 13090
rect 22714 13060 22753 13090
rect 22643 13045 22753 13060
rect 25138 13085 25248 13099
rect 25138 13055 25181 13085
rect 25209 13055 25248 13085
rect 25138 13040 25248 13055
rect 33351 13084 33461 13098
rect 33351 13054 33394 13084
rect 33422 13054 33461 13084
rect 33351 13039 33461 13054
rect 35846 13079 35956 13093
rect 35846 13049 35889 13079
rect 35917 13049 35956 13079
rect 35846 13034 35956 13049
rect 8707 12713 8817 12728
rect 8707 12683 8746 12713
rect 8774 12683 8817 12713
rect 8707 12669 8817 12683
rect 9755 12709 9865 12724
rect 9755 12679 9794 12709
rect 9822 12679 9865 12709
rect 9755 12665 9865 12679
rect 19415 12707 19525 12722
rect 19415 12677 19454 12707
rect 19482 12677 19525 12707
rect 19415 12663 19525 12677
rect 20463 12703 20573 12718
rect 20463 12673 20502 12703
rect 20530 12673 20573 12703
rect 30380 12711 30490 12726
rect 20463 12659 20573 12673
rect 30380 12681 30419 12711
rect 30447 12681 30490 12711
rect 30380 12667 30490 12681
rect 31428 12707 31538 12722
rect 31428 12677 31467 12707
rect 31495 12677 31538 12707
rect 31428 12663 31538 12677
rect 41088 12705 41198 12720
rect 41088 12675 41127 12705
rect 41155 12675 41198 12705
rect 41088 12661 41198 12675
rect 42136 12701 42246 12716
rect 42136 12671 42175 12701
rect 42203 12671 42246 12701
rect 42136 12657 42246 12671
rect 970 12324 1080 12338
rect 970 12294 1013 12324
rect 1041 12294 1080 12324
rect 970 12279 1080 12294
rect 2018 12320 2128 12334
rect 2018 12290 2061 12320
rect 2089 12290 2128 12320
rect 2018 12275 2128 12290
rect 11678 12318 11788 12332
rect 11678 12288 11721 12318
rect 11749 12288 11788 12318
rect 11678 12273 11788 12288
rect 12726 12314 12836 12328
rect 12726 12284 12769 12314
rect 12797 12284 12836 12314
rect 22643 12322 22753 12336
rect 12726 12269 12836 12284
rect 22643 12292 22686 12322
rect 22714 12292 22753 12322
rect 22643 12277 22753 12292
rect 23691 12318 23801 12332
rect 23691 12288 23734 12318
rect 23762 12288 23801 12318
rect 23691 12273 23801 12288
rect 33351 12316 33461 12330
rect 33351 12286 33394 12316
rect 33422 12286 33461 12316
rect 33351 12271 33461 12286
rect 34399 12312 34509 12326
rect 34399 12282 34442 12312
rect 34470 12282 34509 12312
rect 34399 12267 34509 12282
rect 7260 11946 7370 11961
rect 7260 11916 7299 11946
rect 7327 11916 7370 11946
rect 7260 11902 7370 11916
rect 9755 11941 9865 11956
rect 9755 11911 9794 11941
rect 9822 11911 9865 11941
rect 9755 11897 9865 11911
rect 17968 11940 18078 11955
rect 17968 11910 18007 11940
rect 18035 11910 18078 11940
rect 17968 11896 18078 11910
rect 20463 11935 20573 11950
rect 20463 11905 20502 11935
rect 20530 11905 20573 11935
rect 20463 11891 20573 11905
rect 28933 11944 29043 11959
rect 28933 11914 28972 11944
rect 29000 11914 29043 11944
rect 28933 11900 29043 11914
rect 31428 11939 31538 11954
rect 31428 11909 31467 11939
rect 31495 11909 31538 11939
rect 31428 11895 31538 11909
rect 39641 11938 39751 11953
rect 39641 11908 39680 11938
rect 39708 11908 39751 11938
rect 39641 11894 39751 11908
rect 42136 11933 42246 11948
rect 42136 11903 42175 11933
rect 42203 11903 42246 11933
rect 42136 11889 42246 11903
rect 970 11645 1080 11659
rect 970 11615 1013 11645
rect 1041 11615 1080 11645
rect 970 11600 1080 11615
rect 3508 11642 3618 11656
rect 3508 11612 3551 11642
rect 3579 11612 3618 11642
rect 3508 11597 3618 11612
rect 11678 11639 11788 11653
rect 11678 11609 11721 11639
rect 11749 11609 11788 11639
rect 11678 11594 11788 11609
rect 14216 11636 14326 11650
rect 14216 11606 14259 11636
rect 14287 11606 14326 11636
rect 14216 11591 14326 11606
rect 22643 11643 22753 11657
rect 22643 11613 22686 11643
rect 22714 11613 22753 11643
rect 22643 11598 22753 11613
rect 25181 11640 25291 11654
rect 25181 11610 25224 11640
rect 25252 11610 25291 11640
rect 25181 11595 25291 11610
rect 33351 11637 33461 11651
rect 33351 11607 33394 11637
rect 33422 11607 33461 11637
rect 33351 11592 33461 11607
rect 35889 11634 35999 11648
rect 35889 11604 35932 11634
rect 35960 11604 35999 11634
rect 35889 11589 35999 11604
rect 8707 11266 8817 11281
rect 8707 11236 8746 11266
rect 8774 11236 8817 11266
rect 8707 11222 8817 11236
rect 9755 11262 9865 11277
rect 9755 11232 9794 11262
rect 9822 11232 9865 11262
rect 9755 11218 9865 11232
rect 19415 11260 19525 11275
rect 19415 11230 19454 11260
rect 19482 11230 19525 11260
rect 19415 11216 19525 11230
rect 20463 11256 20573 11271
rect 20463 11226 20502 11256
rect 20530 11226 20573 11256
rect 30380 11264 30490 11279
rect 20463 11212 20573 11226
rect 30380 11234 30419 11264
rect 30447 11234 30490 11264
rect 30380 11220 30490 11234
rect 31428 11260 31538 11275
rect 31428 11230 31467 11260
rect 31495 11230 31538 11260
rect 31428 11216 31538 11230
rect 41088 11258 41198 11273
rect 41088 11228 41127 11258
rect 41155 11228 41198 11258
rect 41088 11214 41198 11228
rect 42136 11254 42246 11269
rect 42136 11224 42175 11254
rect 42203 11224 42246 11254
rect 42136 11210 42246 11224
rect 971 10804 1081 10818
rect 971 10774 1014 10804
rect 1042 10774 1081 10804
rect 971 10759 1081 10774
rect 2019 10800 2129 10814
rect 2019 10770 2062 10800
rect 2090 10770 2129 10800
rect 2019 10755 2129 10770
rect 11679 10798 11789 10812
rect 11679 10768 11722 10798
rect 11750 10768 11789 10798
rect 11679 10753 11789 10768
rect 12727 10794 12837 10808
rect 12727 10764 12770 10794
rect 12798 10764 12837 10794
rect 22644 10802 22754 10816
rect 12727 10749 12837 10764
rect 22644 10772 22687 10802
rect 22715 10772 22754 10802
rect 22644 10757 22754 10772
rect 23692 10798 23802 10812
rect 23692 10768 23735 10798
rect 23763 10768 23802 10798
rect 23692 10753 23802 10768
rect 33352 10796 33462 10810
rect 33352 10766 33395 10796
rect 33423 10766 33462 10796
rect 33352 10751 33462 10766
rect 34400 10792 34510 10806
rect 34400 10762 34443 10792
rect 34471 10762 34510 10792
rect 34400 10747 34510 10762
rect 7218 10424 7328 10439
rect 7218 10394 7257 10424
rect 7285 10394 7328 10424
rect 7218 10380 7328 10394
rect 9756 10421 9866 10436
rect 9756 10391 9795 10421
rect 9823 10391 9866 10421
rect 9756 10377 9866 10391
rect 17926 10418 18036 10433
rect 17926 10388 17965 10418
rect 17993 10388 18036 10418
rect 17926 10374 18036 10388
rect 20464 10415 20574 10430
rect 20464 10385 20503 10415
rect 20531 10385 20574 10415
rect 20464 10371 20574 10385
rect 28891 10422 29001 10437
rect 28891 10392 28930 10422
rect 28958 10392 29001 10422
rect 28891 10378 29001 10392
rect 31429 10419 31539 10434
rect 31429 10389 31468 10419
rect 31496 10389 31539 10419
rect 31429 10375 31539 10389
rect 39599 10416 39709 10431
rect 39599 10386 39638 10416
rect 39666 10386 39709 10416
rect 39599 10372 39709 10386
rect 42137 10413 42247 10428
rect 42137 10383 42176 10413
rect 42204 10383 42247 10413
rect 42137 10369 42247 10383
rect 971 10125 1081 10139
rect 971 10095 1014 10125
rect 1042 10095 1081 10125
rect 971 10080 1081 10095
rect 3466 10120 3576 10134
rect 3466 10090 3509 10120
rect 3537 10090 3576 10120
rect 3466 10075 3576 10090
rect 11679 10119 11789 10133
rect 11679 10089 11722 10119
rect 11750 10089 11789 10119
rect 11679 10074 11789 10089
rect 14174 10114 14284 10128
rect 14174 10084 14217 10114
rect 14245 10084 14284 10114
rect 14174 10069 14284 10084
rect 22644 10123 22754 10137
rect 22644 10093 22687 10123
rect 22715 10093 22754 10123
rect 22644 10078 22754 10093
rect 25139 10118 25249 10132
rect 25139 10088 25182 10118
rect 25210 10088 25249 10118
rect 25139 10073 25249 10088
rect 33352 10117 33462 10131
rect 33352 10087 33395 10117
rect 33423 10087 33462 10117
rect 33352 10072 33462 10087
rect 35847 10112 35957 10126
rect 35847 10082 35890 10112
rect 35918 10082 35957 10112
rect 35847 10067 35957 10082
rect 8708 9746 8818 9761
rect 8708 9716 8747 9746
rect 8775 9716 8818 9746
rect 8708 9702 8818 9716
rect 9756 9742 9866 9757
rect 9756 9712 9795 9742
rect 9823 9712 9866 9742
rect 9756 9698 9866 9712
rect 19416 9740 19526 9755
rect 19416 9710 19455 9740
rect 19483 9710 19526 9740
rect 19416 9696 19526 9710
rect 20464 9736 20574 9751
rect 20464 9706 20503 9736
rect 20531 9706 20574 9736
rect 30381 9744 30491 9759
rect 20464 9692 20574 9706
rect 30381 9714 30420 9744
rect 30448 9714 30491 9744
rect 30381 9700 30491 9714
rect 31429 9740 31539 9755
rect 31429 9710 31468 9740
rect 31496 9710 31539 9740
rect 31429 9696 31539 9710
rect 41089 9738 41199 9753
rect 41089 9708 41128 9738
rect 41156 9708 41199 9738
rect 41089 9694 41199 9708
rect 42137 9734 42247 9749
rect 42137 9704 42176 9734
rect 42204 9704 42247 9734
rect 42137 9690 42247 9704
rect 971 9357 1081 9371
rect 971 9327 1014 9357
rect 1042 9327 1081 9357
rect 971 9312 1081 9327
rect 2019 9353 2129 9367
rect 2019 9323 2062 9353
rect 2090 9323 2129 9353
rect 2019 9308 2129 9323
rect 11679 9351 11789 9365
rect 11679 9321 11722 9351
rect 11750 9321 11789 9351
rect 11679 9306 11789 9321
rect 12727 9347 12837 9361
rect 12727 9317 12770 9347
rect 12798 9317 12837 9347
rect 22644 9355 22754 9369
rect 12727 9302 12837 9317
rect 22644 9325 22687 9355
rect 22715 9325 22754 9355
rect 22644 9310 22754 9325
rect 23692 9351 23802 9365
rect 23692 9321 23735 9351
rect 23763 9321 23802 9351
rect 23692 9306 23802 9321
rect 33352 9349 33462 9363
rect 33352 9319 33395 9349
rect 33423 9319 33462 9349
rect 33352 9304 33462 9319
rect 34400 9345 34510 9359
rect 34400 9315 34443 9345
rect 34471 9315 34510 9345
rect 34400 9300 34510 9315
rect 7261 8979 7371 8994
rect 7261 8949 7300 8979
rect 7328 8949 7371 8979
rect 7261 8935 7371 8949
rect 9756 8974 9866 8989
rect 9756 8944 9795 8974
rect 9823 8944 9866 8974
rect 9756 8930 9866 8944
rect 17969 8973 18079 8988
rect 17969 8943 18008 8973
rect 18036 8943 18079 8973
rect 17969 8929 18079 8943
rect 20464 8968 20574 8983
rect 20464 8938 20503 8968
rect 20531 8938 20574 8968
rect 20464 8924 20574 8938
rect 28934 8977 29044 8992
rect 28934 8947 28973 8977
rect 29001 8947 29044 8977
rect 28934 8933 29044 8947
rect 31429 8972 31539 8987
rect 31429 8942 31468 8972
rect 31496 8942 31539 8972
rect 31429 8928 31539 8942
rect 39642 8971 39752 8986
rect 39642 8941 39681 8971
rect 39709 8941 39752 8971
rect 39642 8927 39752 8941
rect 42137 8966 42247 8981
rect 42137 8936 42176 8966
rect 42204 8936 42247 8966
rect 42137 8922 42247 8936
rect 971 8678 1081 8692
rect 971 8648 1014 8678
rect 1042 8648 1081 8678
rect 971 8633 1081 8648
rect 4574 8669 4684 8683
rect 4574 8639 4617 8669
rect 4645 8639 4684 8669
rect 4574 8624 4684 8639
rect 11679 8672 11789 8686
rect 11679 8642 11722 8672
rect 11750 8642 11789 8672
rect 11679 8627 11789 8642
rect 15282 8663 15392 8677
rect 15282 8633 15325 8663
rect 15353 8633 15392 8663
rect 15282 8618 15392 8633
rect 22644 8676 22754 8690
rect 22644 8646 22687 8676
rect 22715 8646 22754 8676
rect 22644 8631 22754 8646
rect 26247 8667 26357 8681
rect 26247 8637 26290 8667
rect 26318 8637 26357 8667
rect 26247 8622 26357 8637
rect 33352 8670 33462 8684
rect 33352 8640 33395 8670
rect 33423 8640 33462 8670
rect 33352 8625 33462 8640
rect 36955 8661 37065 8675
rect 36955 8631 36998 8661
rect 37026 8631 37065 8661
rect 36955 8616 37065 8631
rect 8708 8299 8818 8314
rect 8708 8269 8747 8299
rect 8775 8269 8818 8299
rect 8708 8255 8818 8269
rect 9756 8295 9866 8310
rect 9756 8265 9795 8295
rect 9823 8265 9866 8295
rect 9756 8251 9866 8265
rect 19416 8293 19526 8308
rect 19416 8263 19455 8293
rect 19483 8263 19526 8293
rect 19416 8249 19526 8263
rect 20464 8289 20574 8304
rect 20464 8259 20503 8289
rect 20531 8259 20574 8289
rect 30381 8297 30491 8312
rect 20464 8245 20574 8259
rect 30381 8267 30420 8297
rect 30448 8267 30491 8297
rect 30381 8253 30491 8267
rect 31429 8293 31539 8308
rect 31429 8263 31468 8293
rect 31496 8263 31539 8293
rect 31429 8249 31539 8263
rect 41089 8291 41199 8306
rect 41089 8261 41128 8291
rect 41156 8261 41199 8291
rect 41089 8247 41199 8261
rect 42137 8287 42247 8302
rect 42137 8257 42176 8287
rect 42204 8257 42247 8287
rect 42137 8243 42247 8257
rect 968 7763 1078 7777
rect 968 7733 1011 7763
rect 1039 7733 1078 7763
rect 968 7718 1078 7733
rect 2016 7759 2126 7773
rect 2016 7729 2059 7759
rect 2087 7729 2126 7759
rect 2016 7714 2126 7729
rect 11676 7757 11786 7771
rect 11676 7727 11719 7757
rect 11747 7727 11786 7757
rect 11676 7712 11786 7727
rect 12724 7753 12834 7767
rect 12724 7723 12767 7753
rect 12795 7723 12834 7753
rect 22641 7761 22751 7775
rect 12724 7708 12834 7723
rect 22641 7731 22684 7761
rect 22712 7731 22751 7761
rect 22641 7716 22751 7731
rect 23689 7757 23799 7771
rect 23689 7727 23732 7757
rect 23760 7727 23799 7757
rect 23689 7712 23799 7727
rect 33349 7755 33459 7769
rect 33349 7725 33392 7755
rect 33420 7725 33459 7755
rect 33349 7710 33459 7725
rect 34397 7751 34507 7765
rect 34397 7721 34440 7751
rect 34468 7721 34507 7751
rect 34397 7706 34507 7721
rect 6150 7389 6260 7404
rect 6150 7359 6189 7389
rect 6217 7359 6260 7389
rect 6150 7345 6260 7359
rect 9753 7380 9863 7395
rect 9753 7350 9792 7380
rect 9820 7350 9863 7380
rect 9753 7336 9863 7350
rect 16858 7383 16968 7398
rect 16858 7353 16897 7383
rect 16925 7353 16968 7383
rect 16858 7339 16968 7353
rect 20461 7374 20571 7389
rect 20461 7344 20500 7374
rect 20528 7344 20571 7374
rect 20461 7330 20571 7344
rect 27823 7387 27933 7402
rect 27823 7357 27862 7387
rect 27890 7357 27933 7387
rect 27823 7343 27933 7357
rect 31426 7378 31536 7393
rect 31426 7348 31465 7378
rect 31493 7348 31536 7378
rect 31426 7334 31536 7348
rect 38531 7381 38641 7396
rect 38531 7351 38570 7381
rect 38598 7351 38641 7381
rect 38531 7337 38641 7351
rect 42134 7372 42244 7387
rect 42134 7342 42173 7372
rect 42201 7342 42244 7372
rect 42134 7328 42244 7342
rect 968 7084 1078 7098
rect 968 7054 1011 7084
rect 1039 7054 1078 7084
rect 968 7039 1078 7054
rect 3463 7079 3573 7093
rect 3463 7049 3506 7079
rect 3534 7049 3573 7079
rect 3463 7034 3573 7049
rect 11676 7078 11786 7092
rect 11676 7048 11719 7078
rect 11747 7048 11786 7078
rect 11676 7033 11786 7048
rect 14171 7073 14281 7087
rect 14171 7043 14214 7073
rect 14242 7043 14281 7073
rect 14171 7028 14281 7043
rect 22641 7082 22751 7096
rect 22641 7052 22684 7082
rect 22712 7052 22751 7082
rect 22641 7037 22751 7052
rect 25136 7077 25246 7091
rect 25136 7047 25179 7077
rect 25207 7047 25246 7077
rect 25136 7032 25246 7047
rect 33349 7076 33459 7090
rect 33349 7046 33392 7076
rect 33420 7046 33459 7076
rect 33349 7031 33459 7046
rect 35844 7071 35954 7085
rect 35844 7041 35887 7071
rect 35915 7041 35954 7071
rect 35844 7026 35954 7041
rect 8705 6705 8815 6720
rect 8705 6675 8744 6705
rect 8772 6675 8815 6705
rect 8705 6661 8815 6675
rect 9753 6701 9863 6716
rect 9753 6671 9792 6701
rect 9820 6671 9863 6701
rect 9753 6657 9863 6671
rect 19413 6699 19523 6714
rect 19413 6669 19452 6699
rect 19480 6669 19523 6699
rect 19413 6655 19523 6669
rect 20461 6695 20571 6710
rect 20461 6665 20500 6695
rect 20528 6665 20571 6695
rect 30378 6703 30488 6718
rect 20461 6651 20571 6665
rect 30378 6673 30417 6703
rect 30445 6673 30488 6703
rect 30378 6659 30488 6673
rect 31426 6699 31536 6714
rect 31426 6669 31465 6699
rect 31493 6669 31536 6699
rect 31426 6655 31536 6669
rect 41086 6697 41196 6712
rect 41086 6667 41125 6697
rect 41153 6667 41196 6697
rect 41086 6653 41196 6667
rect 42134 6693 42244 6708
rect 42134 6663 42173 6693
rect 42201 6663 42244 6693
rect 42134 6649 42244 6663
rect 968 6316 1078 6330
rect 968 6286 1011 6316
rect 1039 6286 1078 6316
rect 968 6271 1078 6286
rect 2016 6312 2126 6326
rect 2016 6282 2059 6312
rect 2087 6282 2126 6312
rect 2016 6267 2126 6282
rect 11676 6310 11786 6324
rect 11676 6280 11719 6310
rect 11747 6280 11786 6310
rect 11676 6265 11786 6280
rect 12724 6306 12834 6320
rect 12724 6276 12767 6306
rect 12795 6276 12834 6306
rect 22641 6314 22751 6328
rect 12724 6261 12834 6276
rect 22641 6284 22684 6314
rect 22712 6284 22751 6314
rect 22641 6269 22751 6284
rect 23689 6310 23799 6324
rect 23689 6280 23732 6310
rect 23760 6280 23799 6310
rect 23689 6265 23799 6280
rect 33349 6308 33459 6322
rect 33349 6278 33392 6308
rect 33420 6278 33459 6308
rect 33349 6263 33459 6278
rect 34397 6304 34507 6318
rect 34397 6274 34440 6304
rect 34468 6274 34507 6304
rect 34397 6259 34507 6274
rect 7258 5938 7368 5953
rect 7258 5908 7297 5938
rect 7325 5908 7368 5938
rect 7258 5894 7368 5908
rect 9753 5933 9863 5948
rect 9753 5903 9792 5933
rect 9820 5903 9863 5933
rect 9753 5889 9863 5903
rect 17966 5932 18076 5947
rect 17966 5902 18005 5932
rect 18033 5902 18076 5932
rect 17966 5888 18076 5902
rect 20461 5927 20571 5942
rect 20461 5897 20500 5927
rect 20528 5897 20571 5927
rect 20461 5883 20571 5897
rect 28931 5936 29041 5951
rect 28931 5906 28970 5936
rect 28998 5906 29041 5936
rect 28931 5892 29041 5906
rect 31426 5931 31536 5946
rect 31426 5901 31465 5931
rect 31493 5901 31536 5931
rect 31426 5887 31536 5901
rect 39639 5930 39749 5945
rect 39639 5900 39678 5930
rect 39706 5900 39749 5930
rect 39639 5886 39749 5900
rect 42134 5925 42244 5940
rect 42134 5895 42173 5925
rect 42201 5895 42244 5925
rect 42134 5881 42244 5895
rect 968 5637 1078 5651
rect 968 5607 1011 5637
rect 1039 5607 1078 5637
rect 968 5592 1078 5607
rect 3506 5634 3616 5648
rect 3506 5604 3549 5634
rect 3577 5604 3616 5634
rect 3506 5589 3616 5604
rect 11676 5631 11786 5645
rect 11676 5601 11719 5631
rect 11747 5601 11786 5631
rect 11676 5586 11786 5601
rect 14214 5628 14324 5642
rect 14214 5598 14257 5628
rect 14285 5598 14324 5628
rect 14214 5583 14324 5598
rect 22641 5635 22751 5649
rect 22641 5605 22684 5635
rect 22712 5605 22751 5635
rect 22641 5590 22751 5605
rect 25179 5632 25289 5646
rect 25179 5602 25222 5632
rect 25250 5602 25289 5632
rect 25179 5587 25289 5602
rect 33349 5629 33459 5643
rect 33349 5599 33392 5629
rect 33420 5599 33459 5629
rect 33349 5584 33459 5599
rect 35887 5626 35997 5640
rect 35887 5596 35930 5626
rect 35958 5596 35997 5626
rect 35887 5581 35997 5596
rect 8705 5258 8815 5273
rect 8705 5228 8744 5258
rect 8772 5228 8815 5258
rect 8705 5214 8815 5228
rect 9753 5254 9863 5269
rect 9753 5224 9792 5254
rect 9820 5224 9863 5254
rect 9753 5210 9863 5224
rect 19413 5252 19523 5267
rect 19413 5222 19452 5252
rect 19480 5222 19523 5252
rect 19413 5208 19523 5222
rect 20461 5248 20571 5263
rect 20461 5218 20500 5248
rect 20528 5218 20571 5248
rect 30378 5256 30488 5271
rect 20461 5204 20571 5218
rect 30378 5226 30417 5256
rect 30445 5226 30488 5256
rect 30378 5212 30488 5226
rect 31426 5252 31536 5267
rect 31426 5222 31465 5252
rect 31493 5222 31536 5252
rect 31426 5208 31536 5222
rect 41086 5250 41196 5265
rect 41086 5220 41125 5250
rect 41153 5220 41196 5250
rect 41086 5206 41196 5220
rect 42134 5246 42244 5261
rect 42134 5216 42173 5246
rect 42201 5216 42244 5246
rect 42134 5202 42244 5216
rect 969 4796 1079 4810
rect 969 4766 1012 4796
rect 1040 4766 1079 4796
rect 969 4751 1079 4766
rect 2017 4792 2127 4806
rect 2017 4762 2060 4792
rect 2088 4762 2127 4792
rect 2017 4747 2127 4762
rect 4919 4798 5029 4812
rect 4919 4768 4962 4798
rect 4990 4768 5029 4798
rect 4919 4753 5029 4768
rect 11677 4790 11787 4804
rect 11677 4760 11720 4790
rect 11748 4760 11787 4790
rect 11677 4745 11787 4760
rect 12725 4786 12835 4800
rect 12725 4756 12768 4786
rect 12796 4756 12835 4786
rect 12725 4741 12835 4756
rect 15627 4792 15737 4806
rect 15627 4762 15670 4792
rect 15698 4762 15737 4792
rect 22642 4794 22752 4808
rect 15627 4747 15737 4762
rect 22642 4764 22685 4794
rect 22713 4764 22752 4794
rect 22642 4749 22752 4764
rect 23690 4790 23800 4804
rect 23690 4760 23733 4790
rect 23761 4760 23800 4790
rect 23690 4745 23800 4760
rect 26592 4796 26702 4810
rect 26592 4766 26635 4796
rect 26663 4766 26702 4796
rect 26592 4751 26702 4766
rect 7216 4416 7326 4431
rect 7216 4386 7255 4416
rect 7283 4386 7326 4416
rect 7216 4372 7326 4386
rect 9754 4413 9864 4428
rect 9754 4383 9793 4413
rect 9821 4383 9864 4413
rect 9754 4369 9864 4383
rect 33350 4788 33460 4802
rect 33350 4758 33393 4788
rect 33421 4758 33460 4788
rect 33350 4743 33460 4758
rect 34398 4784 34508 4798
rect 34398 4754 34441 4784
rect 34469 4754 34508 4784
rect 34398 4739 34508 4754
rect 37300 4790 37410 4804
rect 37300 4760 37343 4790
rect 37371 4760 37410 4790
rect 37300 4745 37410 4760
rect 17924 4410 18034 4425
rect 17924 4380 17963 4410
rect 17991 4380 18034 4410
rect 17924 4366 18034 4380
rect 20462 4407 20572 4422
rect 20462 4377 20501 4407
rect 20529 4377 20572 4407
rect 20462 4363 20572 4377
rect 28889 4414 28999 4429
rect 28889 4384 28928 4414
rect 28956 4384 28999 4414
rect 28889 4370 28999 4384
rect 31427 4411 31537 4426
rect 31427 4381 31466 4411
rect 31494 4381 31537 4411
rect 31427 4367 31537 4381
rect 39597 4408 39707 4423
rect 39597 4378 39636 4408
rect 39664 4378 39707 4408
rect 39597 4364 39707 4378
rect 42135 4405 42245 4420
rect 42135 4375 42174 4405
rect 42202 4375 42245 4405
rect 42135 4361 42245 4375
rect 969 4117 1079 4131
rect 969 4087 1012 4117
rect 1040 4087 1079 4117
rect 969 4072 1079 4087
rect 3464 4112 3574 4126
rect 3464 4082 3507 4112
rect 3535 4082 3574 4112
rect 3464 4067 3574 4082
rect 11677 4111 11787 4125
rect 11677 4081 11720 4111
rect 11748 4081 11787 4111
rect 11677 4066 11787 4081
rect 14172 4106 14282 4120
rect 14172 4076 14215 4106
rect 14243 4076 14282 4106
rect 14172 4061 14282 4076
rect 22642 4115 22752 4129
rect 22642 4085 22685 4115
rect 22713 4085 22752 4115
rect 22642 4070 22752 4085
rect 25137 4110 25247 4124
rect 25137 4080 25180 4110
rect 25208 4080 25247 4110
rect 25137 4065 25247 4080
rect 33350 4109 33460 4123
rect 33350 4079 33393 4109
rect 33421 4079 33460 4109
rect 33350 4064 33460 4079
rect 35845 4104 35955 4118
rect 35845 4074 35888 4104
rect 35916 4074 35955 4104
rect 35845 4059 35955 4074
rect 8706 3738 8816 3753
rect 8706 3708 8745 3738
rect 8773 3708 8816 3738
rect 8706 3694 8816 3708
rect 9754 3734 9864 3749
rect 9754 3704 9793 3734
rect 9821 3704 9864 3734
rect 9754 3690 9864 3704
rect 19414 3732 19524 3747
rect 19414 3702 19453 3732
rect 19481 3702 19524 3732
rect 19414 3688 19524 3702
rect 20462 3728 20572 3743
rect 20462 3698 20501 3728
rect 20529 3698 20572 3728
rect 30379 3736 30489 3751
rect 20462 3684 20572 3698
rect 30379 3706 30418 3736
rect 30446 3706 30489 3736
rect 30379 3692 30489 3706
rect 31427 3732 31537 3747
rect 31427 3702 31466 3732
rect 31494 3702 31537 3732
rect 31427 3688 31537 3702
rect 41087 3730 41197 3745
rect 41087 3700 41126 3730
rect 41154 3700 41197 3730
rect 41087 3686 41197 3700
rect 42135 3726 42245 3741
rect 42135 3696 42174 3726
rect 42202 3696 42245 3726
rect 42135 3682 42245 3696
rect 969 3349 1079 3363
rect 969 3319 1012 3349
rect 1040 3319 1079 3349
rect 969 3304 1079 3319
rect 2017 3345 2127 3359
rect 2017 3315 2060 3345
rect 2088 3315 2127 3345
rect 2017 3300 2127 3315
rect 11677 3343 11787 3357
rect 11677 3313 11720 3343
rect 11748 3313 11787 3343
rect 11677 3298 11787 3313
rect 12725 3339 12835 3353
rect 12725 3309 12768 3339
rect 12796 3309 12835 3339
rect 22642 3347 22752 3361
rect 12725 3294 12835 3309
rect 22642 3317 22685 3347
rect 22713 3317 22752 3347
rect 22642 3302 22752 3317
rect 23690 3343 23800 3357
rect 23690 3313 23733 3343
rect 23761 3313 23800 3343
rect 23690 3298 23800 3313
rect 33350 3341 33460 3355
rect 33350 3311 33393 3341
rect 33421 3311 33460 3341
rect 33350 3296 33460 3311
rect 34398 3337 34508 3351
rect 34398 3307 34441 3337
rect 34469 3307 34508 3337
rect 34398 3292 34508 3307
rect 7259 2971 7369 2986
rect 7259 2941 7298 2971
rect 7326 2941 7369 2971
rect 7259 2927 7369 2941
rect 9754 2966 9864 2981
rect 9754 2936 9793 2966
rect 9821 2936 9864 2966
rect 9754 2922 9864 2936
rect 17967 2965 18077 2980
rect 17967 2935 18006 2965
rect 18034 2935 18077 2965
rect 17967 2921 18077 2935
rect 20462 2960 20572 2975
rect 20462 2930 20501 2960
rect 20529 2930 20572 2960
rect 20462 2916 20572 2930
rect 28932 2969 29042 2984
rect 28932 2939 28971 2969
rect 28999 2939 29042 2969
rect 28932 2925 29042 2939
rect 31427 2964 31537 2979
rect 31427 2934 31466 2964
rect 31494 2934 31537 2964
rect 31427 2920 31537 2934
rect 39640 2963 39750 2978
rect 39640 2933 39679 2963
rect 39707 2933 39750 2963
rect 39640 2919 39750 2933
rect 42135 2958 42245 2973
rect 42135 2928 42174 2958
rect 42202 2928 42245 2958
rect 42135 2914 42245 2928
rect 969 2670 1079 2684
rect 969 2640 1012 2670
rect 1040 2640 1079 2670
rect 969 2625 1079 2640
rect 11677 2664 11787 2678
rect 11677 2634 11720 2664
rect 11748 2634 11787 2664
rect 11677 2619 11787 2634
rect 22642 2668 22752 2682
rect 22642 2638 22685 2668
rect 22713 2638 22752 2668
rect 22642 2623 22752 2638
rect 33350 2662 33460 2676
rect 33350 2632 33393 2662
rect 33421 2632 33460 2662
rect 33350 2617 33460 2632
rect 8706 2291 8816 2306
rect 8706 2261 8745 2291
rect 8773 2261 8816 2291
rect 8706 2247 8816 2261
rect 9754 2287 9864 2302
rect 9754 2257 9793 2287
rect 9821 2257 9864 2287
rect 9754 2243 9864 2257
rect 19414 2285 19524 2300
rect 19414 2255 19453 2285
rect 19481 2255 19524 2285
rect 19414 2241 19524 2255
rect 20462 2281 20572 2296
rect 20462 2251 20501 2281
rect 20529 2251 20572 2281
rect 30379 2289 30489 2304
rect 20462 2237 20572 2251
rect 30379 2259 30418 2289
rect 30446 2259 30489 2289
rect 30379 2245 30489 2259
rect 31427 2285 31537 2300
rect 31427 2255 31466 2285
rect 31494 2255 31537 2285
rect 31427 2241 31537 2255
rect 41087 2283 41197 2298
rect 41087 2253 41126 2283
rect 41154 2253 41197 2283
rect 41087 2239 41197 2253
rect 42135 2279 42245 2294
rect 42135 2249 42174 2279
rect 42202 2249 42245 2279
rect 42135 2235 42245 2249
rect 10680 511 10790 525
rect 10680 481 10723 511
rect 10751 481 10790 511
rect 10680 466 10790 481
rect 21317 498 21427 512
rect 21317 468 21360 498
rect 21388 468 21427 498
rect 21317 453 21427 468
rect 32353 509 32463 523
rect 32353 479 32396 509
rect 32424 479 32463 509
rect 32353 464 32463 479
<< psubdiffcont >>
rect 9797 13705 9825 13735
rect 20505 13699 20533 13729
rect 1010 13394 1038 13424
rect 31470 13703 31498 13733
rect 2058 13390 2086 13420
rect 11718 13388 11746 13418
rect 42178 13697 42206 13727
rect 12766 13384 12794 13414
rect 22683 13392 22711 13422
rect 23731 13388 23759 13418
rect 33391 13386 33419 13416
rect 34439 13382 34467 13412
rect 8749 13030 8777 13060
rect 9797 13026 9825 13056
rect 19457 13024 19485 13054
rect 20505 13020 20533 13050
rect 1010 12715 1038 12745
rect 30422 13028 30450 13058
rect 3505 12710 3533 12740
rect 31470 13024 31498 13054
rect 11718 12709 11746 12739
rect 41130 13022 41158 13052
rect 14213 12704 14241 12734
rect 42178 13018 42206 13048
rect 22683 12713 22711 12743
rect 25178 12708 25206 12738
rect 33391 12707 33419 12737
rect 35886 12702 35914 12732
rect 7302 12263 7330 12293
rect 9797 12258 9825 12288
rect 18010 12257 18038 12287
rect 20505 12252 20533 12282
rect 1010 11947 1038 11977
rect 28975 12261 29003 12291
rect 2058 11943 2086 11973
rect 31470 12256 31498 12286
rect 11718 11941 11746 11971
rect 39683 12255 39711 12285
rect 12766 11937 12794 11967
rect 42178 12250 42206 12280
rect 22683 11945 22711 11975
rect 23731 11941 23759 11971
rect 33391 11939 33419 11969
rect 34439 11935 34467 11965
rect 8749 11583 8777 11613
rect 9797 11579 9825 11609
rect 19457 11577 19485 11607
rect 20505 11573 20533 11603
rect 1010 11268 1038 11298
rect 30422 11581 30450 11611
rect 3548 11265 3576 11295
rect 31470 11577 31498 11607
rect 11718 11262 11746 11292
rect 41130 11575 41158 11605
rect 14256 11259 14284 11289
rect 42178 11571 42206 11601
rect 22683 11266 22711 11296
rect 25221 11263 25249 11293
rect 33391 11260 33419 11290
rect 35929 11257 35957 11287
rect 7260 10741 7288 10771
rect 9798 10738 9826 10768
rect 17968 10735 17996 10765
rect 20506 10732 20534 10762
rect 1011 10427 1039 10457
rect 28933 10739 28961 10769
rect 2059 10423 2087 10453
rect 31471 10736 31499 10766
rect 11719 10421 11747 10451
rect 39641 10733 39669 10763
rect 12767 10417 12795 10447
rect 42179 10730 42207 10760
rect 22684 10425 22712 10455
rect 23732 10421 23760 10451
rect 33392 10419 33420 10449
rect 34440 10415 34468 10445
rect 8750 10063 8778 10093
rect 9798 10059 9826 10089
rect 19458 10057 19486 10087
rect 20506 10053 20534 10083
rect 1011 9748 1039 9778
rect 30423 10061 30451 10091
rect 3506 9743 3534 9773
rect 31471 10057 31499 10087
rect 11719 9742 11747 9772
rect 41131 10055 41159 10085
rect 14214 9737 14242 9767
rect 42179 10051 42207 10081
rect 22684 9746 22712 9776
rect 25179 9741 25207 9771
rect 33392 9740 33420 9770
rect 35887 9735 35915 9765
rect 7303 9296 7331 9326
rect 9798 9291 9826 9321
rect 18011 9290 18039 9320
rect 20506 9285 20534 9315
rect 1011 8980 1039 9010
rect 28976 9294 29004 9324
rect 2059 8976 2087 9006
rect 31471 9289 31499 9319
rect 11719 8974 11747 9004
rect 39684 9288 39712 9318
rect 12767 8970 12795 9000
rect 42179 9283 42207 9313
rect 22684 8978 22712 9008
rect 23732 8974 23760 9004
rect 33392 8972 33420 9002
rect 34440 8968 34468 8998
rect 8750 8616 8778 8646
rect 9798 8612 9826 8642
rect 19458 8610 19486 8640
rect 20506 8606 20534 8636
rect 30423 8614 30451 8644
rect 1011 8301 1039 8331
rect 31471 8610 31499 8640
rect 41131 8608 41159 8638
rect 4614 8292 4642 8322
rect 11719 8295 11747 8325
rect 42179 8604 42207 8634
rect 15322 8286 15350 8316
rect 22684 8299 22712 8329
rect 26287 8290 26315 8320
rect 33392 8293 33420 8323
rect 36995 8284 37023 8314
rect 6192 7706 6220 7736
rect 9795 7697 9823 7727
rect 16900 7700 16928 7730
rect 20503 7691 20531 7721
rect 27865 7704 27893 7734
rect 1008 7386 1036 7416
rect 31468 7695 31496 7725
rect 38573 7698 38601 7728
rect 2056 7382 2084 7412
rect 11716 7380 11744 7410
rect 42176 7689 42204 7719
rect 12764 7376 12792 7406
rect 22681 7384 22709 7414
rect 23729 7380 23757 7410
rect 33389 7378 33417 7408
rect 34437 7374 34465 7404
rect 8747 7022 8775 7052
rect 9795 7018 9823 7048
rect 19455 7016 19483 7046
rect 20503 7012 20531 7042
rect 1008 6707 1036 6737
rect 30420 7020 30448 7050
rect 3503 6702 3531 6732
rect 31468 7016 31496 7046
rect 11716 6701 11744 6731
rect 41128 7014 41156 7044
rect 14211 6696 14239 6726
rect 42176 7010 42204 7040
rect 22681 6705 22709 6735
rect 25176 6700 25204 6730
rect 33389 6699 33417 6729
rect 35884 6694 35912 6724
rect 7300 6255 7328 6285
rect 9795 6250 9823 6280
rect 18008 6249 18036 6279
rect 20503 6244 20531 6274
rect 1008 5939 1036 5969
rect 28973 6253 29001 6283
rect 2056 5935 2084 5965
rect 31468 6248 31496 6278
rect 11716 5933 11744 5963
rect 39681 6247 39709 6277
rect 12764 5929 12792 5959
rect 42176 6242 42204 6272
rect 22681 5937 22709 5967
rect 23729 5933 23757 5963
rect 33389 5931 33417 5961
rect 34437 5927 34465 5957
rect 8747 5575 8775 5605
rect 9795 5571 9823 5601
rect 19455 5569 19483 5599
rect 20503 5565 20531 5595
rect 1008 5260 1036 5290
rect 30420 5573 30448 5603
rect 3546 5257 3574 5287
rect 31468 5569 31496 5599
rect 11716 5254 11744 5284
rect 41128 5567 41156 5597
rect 14254 5251 14282 5281
rect 42176 5563 42204 5593
rect 22681 5258 22709 5288
rect 25219 5255 25247 5285
rect 33389 5252 33417 5282
rect 35927 5249 35955 5279
rect 7258 4733 7286 4763
rect 9796 4730 9824 4760
rect 1009 4419 1037 4449
rect 2057 4415 2085 4445
rect 17966 4727 17994 4757
rect 4959 4421 4987 4451
rect 20504 4724 20532 4754
rect 11717 4413 11745 4443
rect 12765 4409 12793 4439
rect 28931 4731 28959 4761
rect 15667 4415 15695 4445
rect 31469 4728 31497 4758
rect 22682 4417 22710 4447
rect 23730 4413 23758 4443
rect 39639 4725 39667 4755
rect 26632 4419 26660 4449
rect 42177 4722 42205 4752
rect 33390 4411 33418 4441
rect 34438 4407 34466 4437
rect 37340 4413 37368 4443
rect 8748 4055 8776 4085
rect 9796 4051 9824 4081
rect 19456 4049 19484 4079
rect 20504 4045 20532 4075
rect 1009 3740 1037 3770
rect 30421 4053 30449 4083
rect 3504 3735 3532 3765
rect 31469 4049 31497 4079
rect 11717 3734 11745 3764
rect 41129 4047 41157 4077
rect 14212 3729 14240 3759
rect 42177 4043 42205 4073
rect 22682 3738 22710 3768
rect 25177 3733 25205 3763
rect 33390 3732 33418 3762
rect 35885 3727 35913 3757
rect 7301 3288 7329 3318
rect 9796 3283 9824 3313
rect 18009 3282 18037 3312
rect 20504 3277 20532 3307
rect 1009 2972 1037 3002
rect 28974 3286 29002 3316
rect 2057 2968 2085 2998
rect 31469 3281 31497 3311
rect 11717 2966 11745 2996
rect 39682 3280 39710 3310
rect 12765 2962 12793 2992
rect 42177 3275 42205 3305
rect 22682 2970 22710 3000
rect 23730 2966 23758 2996
rect 33390 2964 33418 2994
rect 34438 2960 34466 2990
rect 8748 2608 8776 2638
rect 9796 2604 9824 2634
rect 19456 2602 19484 2632
rect 20504 2598 20532 2628
rect 30421 2606 30449 2636
rect 1009 2293 1037 2323
rect 31469 2602 31497 2632
rect 41129 2600 41157 2630
rect 11717 2287 11745 2317
rect 42177 2596 42205 2626
rect 22682 2291 22710 2321
rect 33390 2285 33418 2315
rect 10720 134 10748 164
rect 21357 121 21385 151
rect 32393 132 32421 162
<< nsubdiffcont >>
rect 1013 13741 1041 13771
rect 2061 13737 2089 13767
rect 11721 13735 11749 13765
rect 12769 13731 12797 13761
rect 22686 13739 22714 13769
rect 23734 13735 23762 13765
rect 33394 13733 33422 13763
rect 34442 13729 34470 13759
rect 9794 13358 9822 13388
rect 20502 13352 20530 13382
rect 31467 13356 31495 13386
rect 42175 13350 42203 13380
rect 1013 13062 1041 13092
rect 3508 13057 3536 13087
rect 11721 13056 11749 13086
rect 14216 13051 14244 13081
rect 22686 13060 22714 13090
rect 25181 13055 25209 13085
rect 33394 13054 33422 13084
rect 35889 13049 35917 13079
rect 8746 12683 8774 12713
rect 9794 12679 9822 12709
rect 19454 12677 19482 12707
rect 20502 12673 20530 12703
rect 30419 12681 30447 12711
rect 31467 12677 31495 12707
rect 41127 12675 41155 12705
rect 42175 12671 42203 12701
rect 1013 12294 1041 12324
rect 2061 12290 2089 12320
rect 11721 12288 11749 12318
rect 12769 12284 12797 12314
rect 22686 12292 22714 12322
rect 23734 12288 23762 12318
rect 33394 12286 33422 12316
rect 34442 12282 34470 12312
rect 7299 11916 7327 11946
rect 9794 11911 9822 11941
rect 18007 11910 18035 11940
rect 20502 11905 20530 11935
rect 28972 11914 29000 11944
rect 31467 11909 31495 11939
rect 39680 11908 39708 11938
rect 42175 11903 42203 11933
rect 1013 11615 1041 11645
rect 3551 11612 3579 11642
rect 11721 11609 11749 11639
rect 14259 11606 14287 11636
rect 22686 11613 22714 11643
rect 25224 11610 25252 11640
rect 33394 11607 33422 11637
rect 35932 11604 35960 11634
rect 8746 11236 8774 11266
rect 9794 11232 9822 11262
rect 19454 11230 19482 11260
rect 20502 11226 20530 11256
rect 30419 11234 30447 11264
rect 31467 11230 31495 11260
rect 41127 11228 41155 11258
rect 42175 11224 42203 11254
rect 1014 10774 1042 10804
rect 2062 10770 2090 10800
rect 11722 10768 11750 10798
rect 12770 10764 12798 10794
rect 22687 10772 22715 10802
rect 23735 10768 23763 10798
rect 33395 10766 33423 10796
rect 34443 10762 34471 10792
rect 7257 10394 7285 10424
rect 9795 10391 9823 10421
rect 17965 10388 17993 10418
rect 20503 10385 20531 10415
rect 28930 10392 28958 10422
rect 31468 10389 31496 10419
rect 39638 10386 39666 10416
rect 42176 10383 42204 10413
rect 1014 10095 1042 10125
rect 3509 10090 3537 10120
rect 11722 10089 11750 10119
rect 14217 10084 14245 10114
rect 22687 10093 22715 10123
rect 25182 10088 25210 10118
rect 33395 10087 33423 10117
rect 35890 10082 35918 10112
rect 8747 9716 8775 9746
rect 9795 9712 9823 9742
rect 19455 9710 19483 9740
rect 20503 9706 20531 9736
rect 30420 9714 30448 9744
rect 31468 9710 31496 9740
rect 41128 9708 41156 9738
rect 42176 9704 42204 9734
rect 1014 9327 1042 9357
rect 2062 9323 2090 9353
rect 11722 9321 11750 9351
rect 12770 9317 12798 9347
rect 22687 9325 22715 9355
rect 23735 9321 23763 9351
rect 33395 9319 33423 9349
rect 34443 9315 34471 9345
rect 7300 8949 7328 8979
rect 9795 8944 9823 8974
rect 18008 8943 18036 8973
rect 20503 8938 20531 8968
rect 28973 8947 29001 8977
rect 31468 8942 31496 8972
rect 39681 8941 39709 8971
rect 42176 8936 42204 8966
rect 1014 8648 1042 8678
rect 4617 8639 4645 8669
rect 11722 8642 11750 8672
rect 15325 8633 15353 8663
rect 22687 8646 22715 8676
rect 26290 8637 26318 8667
rect 33395 8640 33423 8670
rect 36998 8631 37026 8661
rect 8747 8269 8775 8299
rect 9795 8265 9823 8295
rect 19455 8263 19483 8293
rect 20503 8259 20531 8289
rect 30420 8267 30448 8297
rect 31468 8263 31496 8293
rect 41128 8261 41156 8291
rect 42176 8257 42204 8287
rect 1011 7733 1039 7763
rect 2059 7729 2087 7759
rect 11719 7727 11747 7757
rect 12767 7723 12795 7753
rect 22684 7731 22712 7761
rect 23732 7727 23760 7757
rect 33392 7725 33420 7755
rect 34440 7721 34468 7751
rect 6189 7359 6217 7389
rect 9792 7350 9820 7380
rect 16897 7353 16925 7383
rect 20500 7344 20528 7374
rect 27862 7357 27890 7387
rect 31465 7348 31493 7378
rect 38570 7351 38598 7381
rect 42173 7342 42201 7372
rect 1011 7054 1039 7084
rect 3506 7049 3534 7079
rect 11719 7048 11747 7078
rect 14214 7043 14242 7073
rect 22684 7052 22712 7082
rect 25179 7047 25207 7077
rect 33392 7046 33420 7076
rect 35887 7041 35915 7071
rect 8744 6675 8772 6705
rect 9792 6671 9820 6701
rect 19452 6669 19480 6699
rect 20500 6665 20528 6695
rect 30417 6673 30445 6703
rect 31465 6669 31493 6699
rect 41125 6667 41153 6697
rect 42173 6663 42201 6693
rect 1011 6286 1039 6316
rect 2059 6282 2087 6312
rect 11719 6280 11747 6310
rect 12767 6276 12795 6306
rect 22684 6284 22712 6314
rect 23732 6280 23760 6310
rect 33392 6278 33420 6308
rect 34440 6274 34468 6304
rect 7297 5908 7325 5938
rect 9792 5903 9820 5933
rect 18005 5902 18033 5932
rect 20500 5897 20528 5927
rect 28970 5906 28998 5936
rect 31465 5901 31493 5931
rect 39678 5900 39706 5930
rect 42173 5895 42201 5925
rect 1011 5607 1039 5637
rect 3549 5604 3577 5634
rect 11719 5601 11747 5631
rect 14257 5598 14285 5628
rect 22684 5605 22712 5635
rect 25222 5602 25250 5632
rect 33392 5599 33420 5629
rect 35930 5596 35958 5626
rect 8744 5228 8772 5258
rect 9792 5224 9820 5254
rect 19452 5222 19480 5252
rect 20500 5218 20528 5248
rect 30417 5226 30445 5256
rect 31465 5222 31493 5252
rect 41125 5220 41153 5250
rect 42173 5216 42201 5246
rect 1012 4766 1040 4796
rect 2060 4762 2088 4792
rect 4962 4768 4990 4798
rect 11720 4760 11748 4790
rect 12768 4756 12796 4786
rect 15670 4762 15698 4792
rect 22685 4764 22713 4794
rect 23733 4760 23761 4790
rect 26635 4766 26663 4796
rect 7255 4386 7283 4416
rect 9793 4383 9821 4413
rect 33393 4758 33421 4788
rect 34441 4754 34469 4784
rect 37343 4760 37371 4790
rect 17963 4380 17991 4410
rect 20501 4377 20529 4407
rect 28928 4384 28956 4414
rect 31466 4381 31494 4411
rect 39636 4378 39664 4408
rect 42174 4375 42202 4405
rect 1012 4087 1040 4117
rect 3507 4082 3535 4112
rect 11720 4081 11748 4111
rect 14215 4076 14243 4106
rect 22685 4085 22713 4115
rect 25180 4080 25208 4110
rect 33393 4079 33421 4109
rect 35888 4074 35916 4104
rect 8745 3708 8773 3738
rect 9793 3704 9821 3734
rect 19453 3702 19481 3732
rect 20501 3698 20529 3728
rect 30418 3706 30446 3736
rect 31466 3702 31494 3732
rect 41126 3700 41154 3730
rect 42174 3696 42202 3726
rect 1012 3319 1040 3349
rect 2060 3315 2088 3345
rect 11720 3313 11748 3343
rect 12768 3309 12796 3339
rect 22685 3317 22713 3347
rect 23733 3313 23761 3343
rect 33393 3311 33421 3341
rect 34441 3307 34469 3337
rect 7298 2941 7326 2971
rect 9793 2936 9821 2966
rect 18006 2935 18034 2965
rect 20501 2930 20529 2960
rect 28971 2939 28999 2969
rect 31466 2934 31494 2964
rect 39679 2933 39707 2963
rect 42174 2928 42202 2958
rect 1012 2640 1040 2670
rect 11720 2634 11748 2664
rect 22685 2638 22713 2668
rect 33393 2632 33421 2662
rect 8745 2261 8773 2291
rect 9793 2257 9821 2287
rect 19453 2255 19481 2285
rect 20501 2251 20529 2281
rect 30418 2259 30446 2289
rect 31466 2255 31494 2285
rect 41126 2253 41154 2283
rect 42174 2249 42202 2279
rect 10723 481 10751 511
rect 21360 468 21388 498
rect 32396 479 32424 509
<< poly >>
rect 933 13698 983 13711
rect 1146 13698 1196 13711
rect 1354 13698 1404 13711
rect 1562 13698 1612 13711
rect 1981 13694 2031 13707
rect 2194 13694 2244 13707
rect 2402 13694 2452 13707
rect 2610 13694 2660 13707
rect 933 13570 983 13598
rect 933 13550 946 13570
rect 966 13550 983 13570
rect 933 13521 983 13550
rect 1146 13569 1196 13598
rect 1146 13545 1157 13569
rect 1181 13545 1196 13569
rect 1146 13521 1196 13545
rect 1354 13574 1404 13598
rect 1354 13550 1366 13574
rect 1390 13550 1404 13574
rect 1354 13521 1404 13550
rect 1562 13572 1612 13598
rect 11641 13692 11691 13705
rect 11854 13692 11904 13705
rect 12062 13692 12112 13705
rect 12270 13692 12320 13705
rect 9223 13650 9273 13666
rect 9431 13650 9481 13666
rect 9639 13650 9689 13666
rect 9852 13650 9902 13666
rect 1562 13546 1580 13572
rect 1606 13546 1612 13572
rect 1562 13521 1612 13546
rect 1981 13566 2031 13594
rect 1981 13546 1994 13566
rect 2014 13546 2031 13566
rect 1981 13517 2031 13546
rect 2194 13565 2244 13594
rect 2194 13541 2205 13565
rect 2229 13541 2244 13565
rect 2194 13517 2244 13541
rect 2402 13570 2452 13594
rect 2402 13546 2414 13570
rect 2438 13546 2452 13570
rect 2402 13517 2452 13546
rect 2610 13568 2660 13594
rect 2610 13542 2628 13568
rect 2654 13542 2660 13568
rect 2610 13517 2660 13542
rect 9223 13583 9273 13608
rect 9223 13557 9229 13583
rect 9255 13557 9273 13583
rect 9223 13531 9273 13557
rect 9431 13579 9481 13608
rect 9431 13555 9445 13579
rect 9469 13555 9481 13579
rect 9431 13531 9481 13555
rect 9639 13584 9689 13608
rect 9639 13560 9654 13584
rect 9678 13560 9689 13584
rect 9639 13531 9689 13560
rect 9852 13579 9902 13608
rect 9852 13559 9869 13579
rect 9889 13559 9902 13579
rect 12689 13688 12739 13701
rect 12902 13688 12952 13701
rect 13110 13688 13160 13701
rect 13318 13688 13368 13701
rect 9852 13531 9902 13559
rect 933 13463 983 13479
rect 1146 13463 1196 13479
rect 1354 13463 1404 13479
rect 1562 13463 1612 13479
rect 1981 13459 2031 13475
rect 2194 13459 2244 13475
rect 2402 13459 2452 13475
rect 2610 13459 2660 13475
rect 11641 13564 11691 13592
rect 11641 13544 11654 13564
rect 11674 13544 11691 13564
rect 11641 13515 11691 13544
rect 11854 13563 11904 13592
rect 11854 13539 11865 13563
rect 11889 13539 11904 13563
rect 11854 13515 11904 13539
rect 12062 13568 12112 13592
rect 12062 13544 12074 13568
rect 12098 13544 12112 13568
rect 12062 13515 12112 13544
rect 12270 13566 12320 13592
rect 22606 13696 22656 13709
rect 22819 13696 22869 13709
rect 23027 13696 23077 13709
rect 23235 13696 23285 13709
rect 19931 13644 19981 13660
rect 20139 13644 20189 13660
rect 20347 13644 20397 13660
rect 20560 13644 20610 13660
rect 12270 13540 12288 13566
rect 12314 13540 12320 13566
rect 12270 13515 12320 13540
rect 12689 13560 12739 13588
rect 12689 13540 12702 13560
rect 12722 13540 12739 13560
rect 12689 13511 12739 13540
rect 12902 13559 12952 13588
rect 12902 13535 12913 13559
rect 12937 13535 12952 13559
rect 12902 13511 12952 13535
rect 13110 13564 13160 13588
rect 13110 13540 13122 13564
rect 13146 13540 13160 13564
rect 13110 13511 13160 13540
rect 13318 13562 13368 13588
rect 13318 13536 13336 13562
rect 13362 13536 13368 13562
rect 13318 13511 13368 13536
rect 19931 13577 19981 13602
rect 19931 13551 19937 13577
rect 19963 13551 19981 13577
rect 19931 13525 19981 13551
rect 20139 13573 20189 13602
rect 20139 13549 20153 13573
rect 20177 13549 20189 13573
rect 20139 13525 20189 13549
rect 20347 13578 20397 13602
rect 20347 13554 20362 13578
rect 20386 13554 20397 13578
rect 20347 13525 20397 13554
rect 20560 13573 20610 13602
rect 23654 13692 23704 13705
rect 23867 13692 23917 13705
rect 24075 13692 24125 13705
rect 24283 13692 24333 13705
rect 20560 13553 20577 13573
rect 20597 13553 20610 13573
rect 20560 13525 20610 13553
rect 11641 13457 11691 13473
rect 11854 13457 11904 13473
rect 12062 13457 12112 13473
rect 12270 13457 12320 13473
rect 12689 13453 12739 13469
rect 12902 13453 12952 13469
rect 13110 13453 13160 13469
rect 13318 13453 13368 13469
rect 9223 13418 9273 13431
rect 9431 13418 9481 13431
rect 9639 13418 9689 13431
rect 9852 13418 9902 13431
rect 22606 13568 22656 13596
rect 22606 13548 22619 13568
rect 22639 13548 22656 13568
rect 22606 13519 22656 13548
rect 22819 13567 22869 13596
rect 22819 13543 22830 13567
rect 22854 13543 22869 13567
rect 22819 13519 22869 13543
rect 23027 13572 23077 13596
rect 23027 13548 23039 13572
rect 23063 13548 23077 13572
rect 23027 13519 23077 13548
rect 23235 13570 23285 13596
rect 33314 13690 33364 13703
rect 33527 13690 33577 13703
rect 33735 13690 33785 13703
rect 33943 13690 33993 13703
rect 30896 13648 30946 13664
rect 31104 13648 31154 13664
rect 31312 13648 31362 13664
rect 31525 13648 31575 13664
rect 23235 13544 23253 13570
rect 23279 13544 23285 13570
rect 23235 13519 23285 13544
rect 23654 13564 23704 13592
rect 23654 13544 23667 13564
rect 23687 13544 23704 13564
rect 23654 13515 23704 13544
rect 23867 13563 23917 13592
rect 23867 13539 23878 13563
rect 23902 13539 23917 13563
rect 23867 13515 23917 13539
rect 24075 13568 24125 13592
rect 24075 13544 24087 13568
rect 24111 13544 24125 13568
rect 24075 13515 24125 13544
rect 24283 13566 24333 13592
rect 24283 13540 24301 13566
rect 24327 13540 24333 13566
rect 24283 13515 24333 13540
rect 30896 13581 30946 13606
rect 30896 13555 30902 13581
rect 30928 13555 30946 13581
rect 30896 13529 30946 13555
rect 31104 13577 31154 13606
rect 31104 13553 31118 13577
rect 31142 13553 31154 13577
rect 31104 13529 31154 13553
rect 31312 13582 31362 13606
rect 31312 13558 31327 13582
rect 31351 13558 31362 13582
rect 31312 13529 31362 13558
rect 31525 13577 31575 13606
rect 31525 13557 31542 13577
rect 31562 13557 31575 13577
rect 34362 13686 34412 13699
rect 34575 13686 34625 13699
rect 34783 13686 34833 13699
rect 34991 13686 35041 13699
rect 31525 13529 31575 13557
rect 22606 13461 22656 13477
rect 22819 13461 22869 13477
rect 23027 13461 23077 13477
rect 23235 13461 23285 13477
rect 23654 13457 23704 13473
rect 23867 13457 23917 13473
rect 24075 13457 24125 13473
rect 24283 13457 24333 13473
rect 19931 13412 19981 13425
rect 20139 13412 20189 13425
rect 20347 13412 20397 13425
rect 20560 13412 20610 13425
rect 33314 13562 33364 13590
rect 33314 13542 33327 13562
rect 33347 13542 33364 13562
rect 33314 13513 33364 13542
rect 33527 13561 33577 13590
rect 33527 13537 33538 13561
rect 33562 13537 33577 13561
rect 33527 13513 33577 13537
rect 33735 13566 33785 13590
rect 33735 13542 33747 13566
rect 33771 13542 33785 13566
rect 33735 13513 33785 13542
rect 33943 13564 33993 13590
rect 41604 13642 41654 13658
rect 41812 13642 41862 13658
rect 42020 13642 42070 13658
rect 42233 13642 42283 13658
rect 33943 13538 33961 13564
rect 33987 13538 33993 13564
rect 33943 13513 33993 13538
rect 34362 13558 34412 13586
rect 34362 13538 34375 13558
rect 34395 13538 34412 13558
rect 34362 13509 34412 13538
rect 34575 13557 34625 13586
rect 34575 13533 34586 13557
rect 34610 13533 34625 13557
rect 34575 13509 34625 13533
rect 34783 13562 34833 13586
rect 34783 13538 34795 13562
rect 34819 13538 34833 13562
rect 34783 13509 34833 13538
rect 34991 13560 35041 13586
rect 34991 13534 35009 13560
rect 35035 13534 35041 13560
rect 34991 13509 35041 13534
rect 41604 13575 41654 13600
rect 41604 13549 41610 13575
rect 41636 13549 41654 13575
rect 41604 13523 41654 13549
rect 41812 13571 41862 13600
rect 41812 13547 41826 13571
rect 41850 13547 41862 13571
rect 41812 13523 41862 13547
rect 42020 13576 42070 13600
rect 42020 13552 42035 13576
rect 42059 13552 42070 13576
rect 42020 13523 42070 13552
rect 42233 13571 42283 13600
rect 42233 13551 42250 13571
rect 42270 13551 42283 13571
rect 42233 13523 42283 13551
rect 33314 13455 33364 13471
rect 33527 13455 33577 13471
rect 33735 13455 33785 13471
rect 33943 13455 33993 13471
rect 34362 13451 34412 13467
rect 34575 13451 34625 13467
rect 34783 13451 34833 13467
rect 34991 13451 35041 13467
rect 30896 13416 30946 13429
rect 31104 13416 31154 13429
rect 31312 13416 31362 13429
rect 31525 13416 31575 13429
rect 41604 13410 41654 13423
rect 41812 13410 41862 13423
rect 42020 13410 42070 13423
rect 42233 13410 42283 13423
rect 933 13019 983 13032
rect 1146 13019 1196 13032
rect 1354 13019 1404 13032
rect 1562 13019 1612 13032
rect 3428 13014 3478 13027
rect 3641 13014 3691 13027
rect 3849 13014 3899 13027
rect 4057 13014 4107 13027
rect 933 12891 983 12919
rect 933 12871 946 12891
rect 966 12871 983 12891
rect 933 12842 983 12871
rect 1146 12890 1196 12919
rect 1146 12866 1157 12890
rect 1181 12866 1196 12890
rect 1146 12842 1196 12866
rect 1354 12895 1404 12919
rect 1354 12871 1366 12895
rect 1390 12871 1404 12895
rect 1354 12842 1404 12871
rect 1562 12893 1612 12919
rect 11641 13013 11691 13026
rect 11854 13013 11904 13026
rect 12062 13013 12112 13026
rect 12270 13013 12320 13026
rect 8175 12975 8225 12991
rect 8383 12975 8433 12991
rect 8591 12975 8641 12991
rect 8804 12975 8854 12991
rect 9223 12971 9273 12987
rect 9431 12971 9481 12987
rect 9639 12971 9689 12987
rect 9852 12971 9902 12987
rect 1562 12867 1580 12893
rect 1606 12867 1612 12893
rect 1562 12842 1612 12867
rect 3428 12886 3478 12914
rect 3428 12866 3441 12886
rect 3461 12866 3478 12886
rect 3428 12837 3478 12866
rect 3641 12885 3691 12914
rect 3641 12861 3652 12885
rect 3676 12861 3691 12885
rect 3641 12837 3691 12861
rect 3849 12890 3899 12914
rect 3849 12866 3861 12890
rect 3885 12866 3899 12890
rect 3849 12837 3899 12866
rect 4057 12888 4107 12914
rect 4057 12862 4075 12888
rect 4101 12862 4107 12888
rect 4057 12837 4107 12862
rect 8175 12908 8225 12933
rect 8175 12882 8181 12908
rect 8207 12882 8225 12908
rect 8175 12856 8225 12882
rect 8383 12904 8433 12933
rect 8383 12880 8397 12904
rect 8421 12880 8433 12904
rect 8383 12856 8433 12880
rect 8591 12909 8641 12933
rect 8591 12885 8606 12909
rect 8630 12885 8641 12909
rect 8591 12856 8641 12885
rect 8804 12904 8854 12933
rect 8804 12884 8821 12904
rect 8841 12884 8854 12904
rect 8804 12856 8854 12884
rect 9223 12904 9273 12929
rect 9223 12878 9229 12904
rect 9255 12878 9273 12904
rect 933 12784 983 12800
rect 1146 12784 1196 12800
rect 1354 12784 1404 12800
rect 1562 12784 1612 12800
rect 3428 12779 3478 12795
rect 3641 12779 3691 12795
rect 3849 12779 3899 12795
rect 4057 12779 4107 12795
rect 9223 12852 9273 12878
rect 9431 12900 9481 12929
rect 9431 12876 9445 12900
rect 9469 12876 9481 12900
rect 9431 12852 9481 12876
rect 9639 12905 9689 12929
rect 9639 12881 9654 12905
rect 9678 12881 9689 12905
rect 9639 12852 9689 12881
rect 9852 12900 9902 12929
rect 9852 12880 9869 12900
rect 9889 12880 9902 12900
rect 9852 12852 9902 12880
rect 14136 13008 14186 13021
rect 14349 13008 14399 13021
rect 14557 13008 14607 13021
rect 14765 13008 14815 13021
rect 11641 12885 11691 12913
rect 8175 12743 8225 12756
rect 8383 12743 8433 12756
rect 8591 12743 8641 12756
rect 8804 12743 8854 12756
rect 11641 12865 11654 12885
rect 11674 12865 11691 12885
rect 11641 12836 11691 12865
rect 11854 12884 11904 12913
rect 11854 12860 11865 12884
rect 11889 12860 11904 12884
rect 11854 12836 11904 12860
rect 12062 12889 12112 12913
rect 12062 12865 12074 12889
rect 12098 12865 12112 12889
rect 12062 12836 12112 12865
rect 12270 12887 12320 12913
rect 22606 13017 22656 13030
rect 22819 13017 22869 13030
rect 23027 13017 23077 13030
rect 23235 13017 23285 13030
rect 18883 12969 18933 12985
rect 19091 12969 19141 12985
rect 19299 12969 19349 12985
rect 19512 12969 19562 12985
rect 19931 12965 19981 12981
rect 20139 12965 20189 12981
rect 20347 12965 20397 12981
rect 20560 12965 20610 12981
rect 12270 12861 12288 12887
rect 12314 12861 12320 12887
rect 12270 12836 12320 12861
rect 14136 12880 14186 12908
rect 14136 12860 14149 12880
rect 14169 12860 14186 12880
rect 14136 12831 14186 12860
rect 14349 12879 14399 12908
rect 14349 12855 14360 12879
rect 14384 12855 14399 12879
rect 14349 12831 14399 12855
rect 14557 12884 14607 12908
rect 14557 12860 14569 12884
rect 14593 12860 14607 12884
rect 14557 12831 14607 12860
rect 14765 12882 14815 12908
rect 14765 12856 14783 12882
rect 14809 12856 14815 12882
rect 14765 12831 14815 12856
rect 18883 12902 18933 12927
rect 18883 12876 18889 12902
rect 18915 12876 18933 12902
rect 18883 12850 18933 12876
rect 19091 12898 19141 12927
rect 19091 12874 19105 12898
rect 19129 12874 19141 12898
rect 19091 12850 19141 12874
rect 19299 12903 19349 12927
rect 19299 12879 19314 12903
rect 19338 12879 19349 12903
rect 19299 12850 19349 12879
rect 19512 12898 19562 12927
rect 19512 12878 19529 12898
rect 19549 12878 19562 12898
rect 19512 12850 19562 12878
rect 19931 12898 19981 12923
rect 19931 12872 19937 12898
rect 19963 12872 19981 12898
rect 11641 12778 11691 12794
rect 11854 12778 11904 12794
rect 12062 12778 12112 12794
rect 12270 12778 12320 12794
rect 14136 12773 14186 12789
rect 14349 12773 14399 12789
rect 14557 12773 14607 12789
rect 14765 12773 14815 12789
rect 9223 12739 9273 12752
rect 9431 12739 9481 12752
rect 9639 12739 9689 12752
rect 9852 12739 9902 12752
rect 19931 12846 19981 12872
rect 20139 12894 20189 12923
rect 20139 12870 20153 12894
rect 20177 12870 20189 12894
rect 20139 12846 20189 12870
rect 20347 12899 20397 12923
rect 20347 12875 20362 12899
rect 20386 12875 20397 12899
rect 20347 12846 20397 12875
rect 20560 12894 20610 12923
rect 20560 12874 20577 12894
rect 20597 12874 20610 12894
rect 20560 12846 20610 12874
rect 25101 13012 25151 13025
rect 25314 13012 25364 13025
rect 25522 13012 25572 13025
rect 25730 13012 25780 13025
rect 22606 12889 22656 12917
rect 22606 12869 22619 12889
rect 22639 12869 22656 12889
rect 18883 12737 18933 12750
rect 19091 12737 19141 12750
rect 19299 12737 19349 12750
rect 19512 12737 19562 12750
rect 22606 12840 22656 12869
rect 22819 12888 22869 12917
rect 22819 12864 22830 12888
rect 22854 12864 22869 12888
rect 22819 12840 22869 12864
rect 23027 12893 23077 12917
rect 23027 12869 23039 12893
rect 23063 12869 23077 12893
rect 23027 12840 23077 12869
rect 23235 12891 23285 12917
rect 33314 13011 33364 13024
rect 33527 13011 33577 13024
rect 33735 13011 33785 13024
rect 33943 13011 33993 13024
rect 29848 12973 29898 12989
rect 30056 12973 30106 12989
rect 30264 12973 30314 12989
rect 30477 12973 30527 12989
rect 30896 12969 30946 12985
rect 31104 12969 31154 12985
rect 31312 12969 31362 12985
rect 31525 12969 31575 12985
rect 23235 12865 23253 12891
rect 23279 12865 23285 12891
rect 23235 12840 23285 12865
rect 25101 12884 25151 12912
rect 25101 12864 25114 12884
rect 25134 12864 25151 12884
rect 25101 12835 25151 12864
rect 25314 12883 25364 12912
rect 25314 12859 25325 12883
rect 25349 12859 25364 12883
rect 25314 12835 25364 12859
rect 25522 12888 25572 12912
rect 25522 12864 25534 12888
rect 25558 12864 25572 12888
rect 25522 12835 25572 12864
rect 25730 12886 25780 12912
rect 25730 12860 25748 12886
rect 25774 12860 25780 12886
rect 25730 12835 25780 12860
rect 29848 12906 29898 12931
rect 29848 12880 29854 12906
rect 29880 12880 29898 12906
rect 29848 12854 29898 12880
rect 30056 12902 30106 12931
rect 30056 12878 30070 12902
rect 30094 12878 30106 12902
rect 30056 12854 30106 12878
rect 30264 12907 30314 12931
rect 30264 12883 30279 12907
rect 30303 12883 30314 12907
rect 30264 12854 30314 12883
rect 30477 12902 30527 12931
rect 30477 12882 30494 12902
rect 30514 12882 30527 12902
rect 30477 12854 30527 12882
rect 30896 12902 30946 12927
rect 30896 12876 30902 12902
rect 30928 12876 30946 12902
rect 22606 12782 22656 12798
rect 22819 12782 22869 12798
rect 23027 12782 23077 12798
rect 23235 12782 23285 12798
rect 25101 12777 25151 12793
rect 25314 12777 25364 12793
rect 25522 12777 25572 12793
rect 25730 12777 25780 12793
rect 19931 12733 19981 12746
rect 20139 12733 20189 12746
rect 20347 12733 20397 12746
rect 20560 12733 20610 12746
rect 30896 12850 30946 12876
rect 31104 12898 31154 12927
rect 31104 12874 31118 12898
rect 31142 12874 31154 12898
rect 31104 12850 31154 12874
rect 31312 12903 31362 12927
rect 31312 12879 31327 12903
rect 31351 12879 31362 12903
rect 31312 12850 31362 12879
rect 31525 12898 31575 12927
rect 31525 12878 31542 12898
rect 31562 12878 31575 12898
rect 31525 12850 31575 12878
rect 35809 13006 35859 13019
rect 36022 13006 36072 13019
rect 36230 13006 36280 13019
rect 36438 13006 36488 13019
rect 33314 12883 33364 12911
rect 29848 12741 29898 12754
rect 30056 12741 30106 12754
rect 30264 12741 30314 12754
rect 30477 12741 30527 12754
rect 33314 12863 33327 12883
rect 33347 12863 33364 12883
rect 33314 12834 33364 12863
rect 33527 12882 33577 12911
rect 33527 12858 33538 12882
rect 33562 12858 33577 12882
rect 33527 12834 33577 12858
rect 33735 12887 33785 12911
rect 33735 12863 33747 12887
rect 33771 12863 33785 12887
rect 33735 12834 33785 12863
rect 33943 12885 33993 12911
rect 40556 12967 40606 12983
rect 40764 12967 40814 12983
rect 40972 12967 41022 12983
rect 41185 12967 41235 12983
rect 41604 12963 41654 12979
rect 41812 12963 41862 12979
rect 42020 12963 42070 12979
rect 42233 12963 42283 12979
rect 33943 12859 33961 12885
rect 33987 12859 33993 12885
rect 33943 12834 33993 12859
rect 35809 12878 35859 12906
rect 35809 12858 35822 12878
rect 35842 12858 35859 12878
rect 35809 12829 35859 12858
rect 36022 12877 36072 12906
rect 36022 12853 36033 12877
rect 36057 12853 36072 12877
rect 36022 12829 36072 12853
rect 36230 12882 36280 12906
rect 36230 12858 36242 12882
rect 36266 12858 36280 12882
rect 36230 12829 36280 12858
rect 36438 12880 36488 12906
rect 36438 12854 36456 12880
rect 36482 12854 36488 12880
rect 36438 12829 36488 12854
rect 40556 12900 40606 12925
rect 40556 12874 40562 12900
rect 40588 12874 40606 12900
rect 40556 12848 40606 12874
rect 40764 12896 40814 12925
rect 40764 12872 40778 12896
rect 40802 12872 40814 12896
rect 40764 12848 40814 12872
rect 40972 12901 41022 12925
rect 40972 12877 40987 12901
rect 41011 12877 41022 12901
rect 40972 12848 41022 12877
rect 41185 12896 41235 12925
rect 41185 12876 41202 12896
rect 41222 12876 41235 12896
rect 41185 12848 41235 12876
rect 41604 12896 41654 12921
rect 41604 12870 41610 12896
rect 41636 12870 41654 12896
rect 33314 12776 33364 12792
rect 33527 12776 33577 12792
rect 33735 12776 33785 12792
rect 33943 12776 33993 12792
rect 35809 12771 35859 12787
rect 36022 12771 36072 12787
rect 36230 12771 36280 12787
rect 36438 12771 36488 12787
rect 30896 12737 30946 12750
rect 31104 12737 31154 12750
rect 31312 12737 31362 12750
rect 31525 12737 31575 12750
rect 41604 12844 41654 12870
rect 41812 12892 41862 12921
rect 41812 12868 41826 12892
rect 41850 12868 41862 12892
rect 41812 12844 41862 12868
rect 42020 12897 42070 12921
rect 42020 12873 42035 12897
rect 42059 12873 42070 12897
rect 42020 12844 42070 12873
rect 42233 12892 42283 12921
rect 42233 12872 42250 12892
rect 42270 12872 42283 12892
rect 42233 12844 42283 12872
rect 40556 12735 40606 12748
rect 40764 12735 40814 12748
rect 40972 12735 41022 12748
rect 41185 12735 41235 12748
rect 41604 12731 41654 12744
rect 41812 12731 41862 12744
rect 42020 12731 42070 12744
rect 42233 12731 42283 12744
rect 933 12251 983 12264
rect 1146 12251 1196 12264
rect 1354 12251 1404 12264
rect 1562 12251 1612 12264
rect 1981 12247 2031 12260
rect 2194 12247 2244 12260
rect 2402 12247 2452 12260
rect 2610 12247 2660 12260
rect 933 12123 983 12151
rect 933 12103 946 12123
rect 966 12103 983 12123
rect 933 12074 983 12103
rect 1146 12122 1196 12151
rect 1146 12098 1157 12122
rect 1181 12098 1196 12122
rect 1146 12074 1196 12098
rect 1354 12127 1404 12151
rect 1354 12103 1366 12127
rect 1390 12103 1404 12127
rect 1354 12074 1404 12103
rect 1562 12125 1612 12151
rect 11641 12245 11691 12258
rect 11854 12245 11904 12258
rect 12062 12245 12112 12258
rect 12270 12245 12320 12258
rect 6728 12208 6778 12224
rect 6936 12208 6986 12224
rect 7144 12208 7194 12224
rect 7357 12208 7407 12224
rect 9223 12203 9273 12219
rect 9431 12203 9481 12219
rect 9639 12203 9689 12219
rect 9852 12203 9902 12219
rect 1562 12099 1580 12125
rect 1606 12099 1612 12125
rect 1562 12074 1612 12099
rect 1981 12119 2031 12147
rect 1981 12099 1994 12119
rect 2014 12099 2031 12119
rect 1981 12070 2031 12099
rect 2194 12118 2244 12147
rect 2194 12094 2205 12118
rect 2229 12094 2244 12118
rect 2194 12070 2244 12094
rect 2402 12123 2452 12147
rect 2402 12099 2414 12123
rect 2438 12099 2452 12123
rect 2402 12070 2452 12099
rect 2610 12121 2660 12147
rect 2610 12095 2628 12121
rect 2654 12095 2660 12121
rect 2610 12070 2660 12095
rect 6728 12141 6778 12166
rect 6728 12115 6734 12141
rect 6760 12115 6778 12141
rect 6728 12089 6778 12115
rect 6936 12137 6986 12166
rect 6936 12113 6950 12137
rect 6974 12113 6986 12137
rect 6936 12089 6986 12113
rect 7144 12142 7194 12166
rect 7144 12118 7159 12142
rect 7183 12118 7194 12142
rect 7144 12089 7194 12118
rect 7357 12137 7407 12166
rect 7357 12117 7374 12137
rect 7394 12117 7407 12137
rect 7357 12089 7407 12117
rect 9223 12136 9273 12161
rect 9223 12110 9229 12136
rect 9255 12110 9273 12136
rect 933 12016 983 12032
rect 1146 12016 1196 12032
rect 1354 12016 1404 12032
rect 1562 12016 1612 12032
rect 1981 12012 2031 12028
rect 2194 12012 2244 12028
rect 2402 12012 2452 12028
rect 2610 12012 2660 12028
rect 9223 12084 9273 12110
rect 9431 12132 9481 12161
rect 9431 12108 9445 12132
rect 9469 12108 9481 12132
rect 9431 12084 9481 12108
rect 9639 12137 9689 12161
rect 9639 12113 9654 12137
rect 9678 12113 9689 12137
rect 9639 12084 9689 12113
rect 9852 12132 9902 12161
rect 9852 12112 9869 12132
rect 9889 12112 9902 12132
rect 12689 12241 12739 12254
rect 12902 12241 12952 12254
rect 13110 12241 13160 12254
rect 13318 12241 13368 12254
rect 9852 12084 9902 12112
rect 6728 11976 6778 11989
rect 6936 11976 6986 11989
rect 7144 11976 7194 11989
rect 7357 11976 7407 11989
rect 11641 12117 11691 12145
rect 11641 12097 11654 12117
rect 11674 12097 11691 12117
rect 11641 12068 11691 12097
rect 11854 12116 11904 12145
rect 11854 12092 11865 12116
rect 11889 12092 11904 12116
rect 11854 12068 11904 12092
rect 12062 12121 12112 12145
rect 12062 12097 12074 12121
rect 12098 12097 12112 12121
rect 12062 12068 12112 12097
rect 12270 12119 12320 12145
rect 22606 12249 22656 12262
rect 22819 12249 22869 12262
rect 23027 12249 23077 12262
rect 23235 12249 23285 12262
rect 17436 12202 17486 12218
rect 17644 12202 17694 12218
rect 17852 12202 17902 12218
rect 18065 12202 18115 12218
rect 19931 12197 19981 12213
rect 20139 12197 20189 12213
rect 20347 12197 20397 12213
rect 20560 12197 20610 12213
rect 12270 12093 12288 12119
rect 12314 12093 12320 12119
rect 12270 12068 12320 12093
rect 12689 12113 12739 12141
rect 12689 12093 12702 12113
rect 12722 12093 12739 12113
rect 12689 12064 12739 12093
rect 12902 12112 12952 12141
rect 12902 12088 12913 12112
rect 12937 12088 12952 12112
rect 12902 12064 12952 12088
rect 13110 12117 13160 12141
rect 13110 12093 13122 12117
rect 13146 12093 13160 12117
rect 13110 12064 13160 12093
rect 13318 12115 13368 12141
rect 13318 12089 13336 12115
rect 13362 12089 13368 12115
rect 13318 12064 13368 12089
rect 17436 12135 17486 12160
rect 17436 12109 17442 12135
rect 17468 12109 17486 12135
rect 17436 12083 17486 12109
rect 17644 12131 17694 12160
rect 17644 12107 17658 12131
rect 17682 12107 17694 12131
rect 17644 12083 17694 12107
rect 17852 12136 17902 12160
rect 17852 12112 17867 12136
rect 17891 12112 17902 12136
rect 17852 12083 17902 12112
rect 18065 12131 18115 12160
rect 18065 12111 18082 12131
rect 18102 12111 18115 12131
rect 18065 12083 18115 12111
rect 19931 12130 19981 12155
rect 19931 12104 19937 12130
rect 19963 12104 19981 12130
rect 11641 12010 11691 12026
rect 11854 12010 11904 12026
rect 12062 12010 12112 12026
rect 12270 12010 12320 12026
rect 12689 12006 12739 12022
rect 12902 12006 12952 12022
rect 13110 12006 13160 12022
rect 13318 12006 13368 12022
rect 9223 11971 9273 11984
rect 9431 11971 9481 11984
rect 9639 11971 9689 11984
rect 9852 11971 9902 11984
rect 19931 12078 19981 12104
rect 20139 12126 20189 12155
rect 20139 12102 20153 12126
rect 20177 12102 20189 12126
rect 20139 12078 20189 12102
rect 20347 12131 20397 12155
rect 20347 12107 20362 12131
rect 20386 12107 20397 12131
rect 20347 12078 20397 12107
rect 20560 12126 20610 12155
rect 23654 12245 23704 12258
rect 23867 12245 23917 12258
rect 24075 12245 24125 12258
rect 24283 12245 24333 12258
rect 20560 12106 20577 12126
rect 20597 12106 20610 12126
rect 20560 12078 20610 12106
rect 17436 11970 17486 11983
rect 17644 11970 17694 11983
rect 17852 11970 17902 11983
rect 18065 11970 18115 11983
rect 22606 12121 22656 12149
rect 22606 12101 22619 12121
rect 22639 12101 22656 12121
rect 22606 12072 22656 12101
rect 22819 12120 22869 12149
rect 22819 12096 22830 12120
rect 22854 12096 22869 12120
rect 22819 12072 22869 12096
rect 23027 12125 23077 12149
rect 23027 12101 23039 12125
rect 23063 12101 23077 12125
rect 23027 12072 23077 12101
rect 23235 12123 23285 12149
rect 33314 12243 33364 12256
rect 33527 12243 33577 12256
rect 33735 12243 33785 12256
rect 33943 12243 33993 12256
rect 28401 12206 28451 12222
rect 28609 12206 28659 12222
rect 28817 12206 28867 12222
rect 29030 12206 29080 12222
rect 30896 12201 30946 12217
rect 31104 12201 31154 12217
rect 31312 12201 31362 12217
rect 31525 12201 31575 12217
rect 23235 12097 23253 12123
rect 23279 12097 23285 12123
rect 23235 12072 23285 12097
rect 23654 12117 23704 12145
rect 23654 12097 23667 12117
rect 23687 12097 23704 12117
rect 23654 12068 23704 12097
rect 23867 12116 23917 12145
rect 23867 12092 23878 12116
rect 23902 12092 23917 12116
rect 23867 12068 23917 12092
rect 24075 12121 24125 12145
rect 24075 12097 24087 12121
rect 24111 12097 24125 12121
rect 24075 12068 24125 12097
rect 24283 12119 24333 12145
rect 24283 12093 24301 12119
rect 24327 12093 24333 12119
rect 24283 12068 24333 12093
rect 28401 12139 28451 12164
rect 28401 12113 28407 12139
rect 28433 12113 28451 12139
rect 28401 12087 28451 12113
rect 28609 12135 28659 12164
rect 28609 12111 28623 12135
rect 28647 12111 28659 12135
rect 28609 12087 28659 12111
rect 28817 12140 28867 12164
rect 28817 12116 28832 12140
rect 28856 12116 28867 12140
rect 28817 12087 28867 12116
rect 29030 12135 29080 12164
rect 29030 12115 29047 12135
rect 29067 12115 29080 12135
rect 29030 12087 29080 12115
rect 30896 12134 30946 12159
rect 30896 12108 30902 12134
rect 30928 12108 30946 12134
rect 22606 12014 22656 12030
rect 22819 12014 22869 12030
rect 23027 12014 23077 12030
rect 23235 12014 23285 12030
rect 23654 12010 23704 12026
rect 23867 12010 23917 12026
rect 24075 12010 24125 12026
rect 24283 12010 24333 12026
rect 19931 11965 19981 11978
rect 20139 11965 20189 11978
rect 20347 11965 20397 11978
rect 20560 11965 20610 11978
rect 30896 12082 30946 12108
rect 31104 12130 31154 12159
rect 31104 12106 31118 12130
rect 31142 12106 31154 12130
rect 31104 12082 31154 12106
rect 31312 12135 31362 12159
rect 31312 12111 31327 12135
rect 31351 12111 31362 12135
rect 31312 12082 31362 12111
rect 31525 12130 31575 12159
rect 31525 12110 31542 12130
rect 31562 12110 31575 12130
rect 34362 12239 34412 12252
rect 34575 12239 34625 12252
rect 34783 12239 34833 12252
rect 34991 12239 35041 12252
rect 31525 12082 31575 12110
rect 28401 11974 28451 11987
rect 28609 11974 28659 11987
rect 28817 11974 28867 11987
rect 29030 11974 29080 11987
rect 33314 12115 33364 12143
rect 33314 12095 33327 12115
rect 33347 12095 33364 12115
rect 33314 12066 33364 12095
rect 33527 12114 33577 12143
rect 33527 12090 33538 12114
rect 33562 12090 33577 12114
rect 33527 12066 33577 12090
rect 33735 12119 33785 12143
rect 33735 12095 33747 12119
rect 33771 12095 33785 12119
rect 33735 12066 33785 12095
rect 33943 12117 33993 12143
rect 39109 12200 39159 12216
rect 39317 12200 39367 12216
rect 39525 12200 39575 12216
rect 39738 12200 39788 12216
rect 41604 12195 41654 12211
rect 41812 12195 41862 12211
rect 42020 12195 42070 12211
rect 42233 12195 42283 12211
rect 33943 12091 33961 12117
rect 33987 12091 33993 12117
rect 33943 12066 33993 12091
rect 34362 12111 34412 12139
rect 34362 12091 34375 12111
rect 34395 12091 34412 12111
rect 34362 12062 34412 12091
rect 34575 12110 34625 12139
rect 34575 12086 34586 12110
rect 34610 12086 34625 12110
rect 34575 12062 34625 12086
rect 34783 12115 34833 12139
rect 34783 12091 34795 12115
rect 34819 12091 34833 12115
rect 34783 12062 34833 12091
rect 34991 12113 35041 12139
rect 34991 12087 35009 12113
rect 35035 12087 35041 12113
rect 34991 12062 35041 12087
rect 39109 12133 39159 12158
rect 39109 12107 39115 12133
rect 39141 12107 39159 12133
rect 39109 12081 39159 12107
rect 39317 12129 39367 12158
rect 39317 12105 39331 12129
rect 39355 12105 39367 12129
rect 39317 12081 39367 12105
rect 39525 12134 39575 12158
rect 39525 12110 39540 12134
rect 39564 12110 39575 12134
rect 39525 12081 39575 12110
rect 39738 12129 39788 12158
rect 39738 12109 39755 12129
rect 39775 12109 39788 12129
rect 39738 12081 39788 12109
rect 41604 12128 41654 12153
rect 41604 12102 41610 12128
rect 41636 12102 41654 12128
rect 33314 12008 33364 12024
rect 33527 12008 33577 12024
rect 33735 12008 33785 12024
rect 33943 12008 33993 12024
rect 34362 12004 34412 12020
rect 34575 12004 34625 12020
rect 34783 12004 34833 12020
rect 34991 12004 35041 12020
rect 30896 11969 30946 11982
rect 31104 11969 31154 11982
rect 31312 11969 31362 11982
rect 31525 11969 31575 11982
rect 41604 12076 41654 12102
rect 41812 12124 41862 12153
rect 41812 12100 41826 12124
rect 41850 12100 41862 12124
rect 41812 12076 41862 12100
rect 42020 12129 42070 12153
rect 42020 12105 42035 12129
rect 42059 12105 42070 12129
rect 42020 12076 42070 12105
rect 42233 12124 42283 12153
rect 42233 12104 42250 12124
rect 42270 12104 42283 12124
rect 42233 12076 42283 12104
rect 39109 11968 39159 11981
rect 39317 11968 39367 11981
rect 39525 11968 39575 11981
rect 39738 11968 39788 11981
rect 41604 11963 41654 11976
rect 41812 11963 41862 11976
rect 42020 11963 42070 11976
rect 42233 11963 42283 11976
rect 933 11572 983 11585
rect 1146 11572 1196 11585
rect 1354 11572 1404 11585
rect 1562 11572 1612 11585
rect 3471 11569 3521 11582
rect 3684 11569 3734 11582
rect 3892 11569 3942 11582
rect 4100 11569 4150 11582
rect 933 11444 983 11472
rect 933 11424 946 11444
rect 966 11424 983 11444
rect 933 11395 983 11424
rect 1146 11443 1196 11472
rect 1146 11419 1157 11443
rect 1181 11419 1196 11443
rect 1146 11395 1196 11419
rect 1354 11448 1404 11472
rect 1354 11424 1366 11448
rect 1390 11424 1404 11448
rect 1354 11395 1404 11424
rect 1562 11446 1612 11472
rect 11641 11566 11691 11579
rect 11854 11566 11904 11579
rect 12062 11566 12112 11579
rect 12270 11566 12320 11579
rect 8175 11528 8225 11544
rect 8383 11528 8433 11544
rect 8591 11528 8641 11544
rect 8804 11528 8854 11544
rect 9223 11524 9273 11540
rect 9431 11524 9481 11540
rect 9639 11524 9689 11540
rect 9852 11524 9902 11540
rect 1562 11420 1580 11446
rect 1606 11420 1612 11446
rect 1562 11395 1612 11420
rect 3471 11441 3521 11469
rect 3471 11421 3484 11441
rect 3504 11421 3521 11441
rect 3471 11392 3521 11421
rect 3684 11440 3734 11469
rect 3684 11416 3695 11440
rect 3719 11416 3734 11440
rect 3684 11392 3734 11416
rect 3892 11445 3942 11469
rect 3892 11421 3904 11445
rect 3928 11421 3942 11445
rect 3892 11392 3942 11421
rect 4100 11443 4150 11469
rect 4100 11417 4118 11443
rect 4144 11417 4150 11443
rect 4100 11392 4150 11417
rect 8175 11461 8225 11486
rect 8175 11435 8181 11461
rect 8207 11435 8225 11461
rect 8175 11409 8225 11435
rect 8383 11457 8433 11486
rect 8383 11433 8397 11457
rect 8421 11433 8433 11457
rect 8383 11409 8433 11433
rect 8591 11462 8641 11486
rect 8591 11438 8606 11462
rect 8630 11438 8641 11462
rect 8591 11409 8641 11438
rect 8804 11457 8854 11486
rect 8804 11437 8821 11457
rect 8841 11437 8854 11457
rect 8804 11409 8854 11437
rect 9223 11457 9273 11482
rect 9223 11431 9229 11457
rect 9255 11431 9273 11457
rect 933 11337 983 11353
rect 1146 11337 1196 11353
rect 1354 11337 1404 11353
rect 1562 11337 1612 11353
rect 3471 11334 3521 11350
rect 3684 11334 3734 11350
rect 3892 11334 3942 11350
rect 4100 11334 4150 11350
rect 9223 11405 9273 11431
rect 9431 11453 9481 11482
rect 9431 11429 9445 11453
rect 9469 11429 9481 11453
rect 9431 11405 9481 11429
rect 9639 11458 9689 11482
rect 9639 11434 9654 11458
rect 9678 11434 9689 11458
rect 9639 11405 9689 11434
rect 9852 11453 9902 11482
rect 9852 11433 9869 11453
rect 9889 11433 9902 11453
rect 9852 11405 9902 11433
rect 14179 11563 14229 11576
rect 14392 11563 14442 11576
rect 14600 11563 14650 11576
rect 14808 11563 14858 11576
rect 11641 11438 11691 11466
rect 8175 11296 8225 11309
rect 8383 11296 8433 11309
rect 8591 11296 8641 11309
rect 8804 11296 8854 11309
rect 11641 11418 11654 11438
rect 11674 11418 11691 11438
rect 11641 11389 11691 11418
rect 11854 11437 11904 11466
rect 11854 11413 11865 11437
rect 11889 11413 11904 11437
rect 11854 11389 11904 11413
rect 12062 11442 12112 11466
rect 12062 11418 12074 11442
rect 12098 11418 12112 11442
rect 12062 11389 12112 11418
rect 12270 11440 12320 11466
rect 22606 11570 22656 11583
rect 22819 11570 22869 11583
rect 23027 11570 23077 11583
rect 23235 11570 23285 11583
rect 18883 11522 18933 11538
rect 19091 11522 19141 11538
rect 19299 11522 19349 11538
rect 19512 11522 19562 11538
rect 19931 11518 19981 11534
rect 20139 11518 20189 11534
rect 20347 11518 20397 11534
rect 20560 11518 20610 11534
rect 12270 11414 12288 11440
rect 12314 11414 12320 11440
rect 12270 11389 12320 11414
rect 14179 11435 14229 11463
rect 14179 11415 14192 11435
rect 14212 11415 14229 11435
rect 14179 11386 14229 11415
rect 14392 11434 14442 11463
rect 14392 11410 14403 11434
rect 14427 11410 14442 11434
rect 14392 11386 14442 11410
rect 14600 11439 14650 11463
rect 14600 11415 14612 11439
rect 14636 11415 14650 11439
rect 14600 11386 14650 11415
rect 14808 11437 14858 11463
rect 14808 11411 14826 11437
rect 14852 11411 14858 11437
rect 14808 11386 14858 11411
rect 18883 11455 18933 11480
rect 18883 11429 18889 11455
rect 18915 11429 18933 11455
rect 18883 11403 18933 11429
rect 19091 11451 19141 11480
rect 19091 11427 19105 11451
rect 19129 11427 19141 11451
rect 19091 11403 19141 11427
rect 19299 11456 19349 11480
rect 19299 11432 19314 11456
rect 19338 11432 19349 11456
rect 19299 11403 19349 11432
rect 19512 11451 19562 11480
rect 19512 11431 19529 11451
rect 19549 11431 19562 11451
rect 19512 11403 19562 11431
rect 19931 11451 19981 11476
rect 19931 11425 19937 11451
rect 19963 11425 19981 11451
rect 11641 11331 11691 11347
rect 11854 11331 11904 11347
rect 12062 11331 12112 11347
rect 12270 11331 12320 11347
rect 14179 11328 14229 11344
rect 14392 11328 14442 11344
rect 14600 11328 14650 11344
rect 14808 11328 14858 11344
rect 9223 11292 9273 11305
rect 9431 11292 9481 11305
rect 9639 11292 9689 11305
rect 9852 11292 9902 11305
rect 19931 11399 19981 11425
rect 20139 11447 20189 11476
rect 20139 11423 20153 11447
rect 20177 11423 20189 11447
rect 20139 11399 20189 11423
rect 20347 11452 20397 11476
rect 20347 11428 20362 11452
rect 20386 11428 20397 11452
rect 20347 11399 20397 11428
rect 20560 11447 20610 11476
rect 20560 11427 20577 11447
rect 20597 11427 20610 11447
rect 20560 11399 20610 11427
rect 25144 11567 25194 11580
rect 25357 11567 25407 11580
rect 25565 11567 25615 11580
rect 25773 11567 25823 11580
rect 22606 11442 22656 11470
rect 22606 11422 22619 11442
rect 22639 11422 22656 11442
rect 18883 11290 18933 11303
rect 19091 11290 19141 11303
rect 19299 11290 19349 11303
rect 19512 11290 19562 11303
rect 22606 11393 22656 11422
rect 22819 11441 22869 11470
rect 22819 11417 22830 11441
rect 22854 11417 22869 11441
rect 22819 11393 22869 11417
rect 23027 11446 23077 11470
rect 23027 11422 23039 11446
rect 23063 11422 23077 11446
rect 23027 11393 23077 11422
rect 23235 11444 23285 11470
rect 33314 11564 33364 11577
rect 33527 11564 33577 11577
rect 33735 11564 33785 11577
rect 33943 11564 33993 11577
rect 29848 11526 29898 11542
rect 30056 11526 30106 11542
rect 30264 11526 30314 11542
rect 30477 11526 30527 11542
rect 30896 11522 30946 11538
rect 31104 11522 31154 11538
rect 31312 11522 31362 11538
rect 31525 11522 31575 11538
rect 23235 11418 23253 11444
rect 23279 11418 23285 11444
rect 23235 11393 23285 11418
rect 25144 11439 25194 11467
rect 25144 11419 25157 11439
rect 25177 11419 25194 11439
rect 25144 11390 25194 11419
rect 25357 11438 25407 11467
rect 25357 11414 25368 11438
rect 25392 11414 25407 11438
rect 25357 11390 25407 11414
rect 25565 11443 25615 11467
rect 25565 11419 25577 11443
rect 25601 11419 25615 11443
rect 25565 11390 25615 11419
rect 25773 11441 25823 11467
rect 25773 11415 25791 11441
rect 25817 11415 25823 11441
rect 25773 11390 25823 11415
rect 29848 11459 29898 11484
rect 29848 11433 29854 11459
rect 29880 11433 29898 11459
rect 29848 11407 29898 11433
rect 30056 11455 30106 11484
rect 30056 11431 30070 11455
rect 30094 11431 30106 11455
rect 30056 11407 30106 11431
rect 30264 11460 30314 11484
rect 30264 11436 30279 11460
rect 30303 11436 30314 11460
rect 30264 11407 30314 11436
rect 30477 11455 30527 11484
rect 30477 11435 30494 11455
rect 30514 11435 30527 11455
rect 30477 11407 30527 11435
rect 30896 11455 30946 11480
rect 30896 11429 30902 11455
rect 30928 11429 30946 11455
rect 22606 11335 22656 11351
rect 22819 11335 22869 11351
rect 23027 11335 23077 11351
rect 23235 11335 23285 11351
rect 25144 11332 25194 11348
rect 25357 11332 25407 11348
rect 25565 11332 25615 11348
rect 25773 11332 25823 11348
rect 19931 11286 19981 11299
rect 20139 11286 20189 11299
rect 20347 11286 20397 11299
rect 20560 11286 20610 11299
rect 30896 11403 30946 11429
rect 31104 11451 31154 11480
rect 31104 11427 31118 11451
rect 31142 11427 31154 11451
rect 31104 11403 31154 11427
rect 31312 11456 31362 11480
rect 31312 11432 31327 11456
rect 31351 11432 31362 11456
rect 31312 11403 31362 11432
rect 31525 11451 31575 11480
rect 31525 11431 31542 11451
rect 31562 11431 31575 11451
rect 31525 11403 31575 11431
rect 35852 11561 35902 11574
rect 36065 11561 36115 11574
rect 36273 11561 36323 11574
rect 36481 11561 36531 11574
rect 33314 11436 33364 11464
rect 29848 11294 29898 11307
rect 30056 11294 30106 11307
rect 30264 11294 30314 11307
rect 30477 11294 30527 11307
rect 33314 11416 33327 11436
rect 33347 11416 33364 11436
rect 33314 11387 33364 11416
rect 33527 11435 33577 11464
rect 33527 11411 33538 11435
rect 33562 11411 33577 11435
rect 33527 11387 33577 11411
rect 33735 11440 33785 11464
rect 33735 11416 33747 11440
rect 33771 11416 33785 11440
rect 33735 11387 33785 11416
rect 33943 11438 33993 11464
rect 40556 11520 40606 11536
rect 40764 11520 40814 11536
rect 40972 11520 41022 11536
rect 41185 11520 41235 11536
rect 41604 11516 41654 11532
rect 41812 11516 41862 11532
rect 42020 11516 42070 11532
rect 42233 11516 42283 11532
rect 33943 11412 33961 11438
rect 33987 11412 33993 11438
rect 33943 11387 33993 11412
rect 35852 11433 35902 11461
rect 35852 11413 35865 11433
rect 35885 11413 35902 11433
rect 35852 11384 35902 11413
rect 36065 11432 36115 11461
rect 36065 11408 36076 11432
rect 36100 11408 36115 11432
rect 36065 11384 36115 11408
rect 36273 11437 36323 11461
rect 36273 11413 36285 11437
rect 36309 11413 36323 11437
rect 36273 11384 36323 11413
rect 36481 11435 36531 11461
rect 36481 11409 36499 11435
rect 36525 11409 36531 11435
rect 36481 11384 36531 11409
rect 40556 11453 40606 11478
rect 40556 11427 40562 11453
rect 40588 11427 40606 11453
rect 40556 11401 40606 11427
rect 40764 11449 40814 11478
rect 40764 11425 40778 11449
rect 40802 11425 40814 11449
rect 40764 11401 40814 11425
rect 40972 11454 41022 11478
rect 40972 11430 40987 11454
rect 41011 11430 41022 11454
rect 40972 11401 41022 11430
rect 41185 11449 41235 11478
rect 41185 11429 41202 11449
rect 41222 11429 41235 11449
rect 41185 11401 41235 11429
rect 41604 11449 41654 11474
rect 41604 11423 41610 11449
rect 41636 11423 41654 11449
rect 33314 11329 33364 11345
rect 33527 11329 33577 11345
rect 33735 11329 33785 11345
rect 33943 11329 33993 11345
rect 35852 11326 35902 11342
rect 36065 11326 36115 11342
rect 36273 11326 36323 11342
rect 36481 11326 36531 11342
rect 30896 11290 30946 11303
rect 31104 11290 31154 11303
rect 31312 11290 31362 11303
rect 31525 11290 31575 11303
rect 41604 11397 41654 11423
rect 41812 11445 41862 11474
rect 41812 11421 41826 11445
rect 41850 11421 41862 11445
rect 41812 11397 41862 11421
rect 42020 11450 42070 11474
rect 42020 11426 42035 11450
rect 42059 11426 42070 11450
rect 42020 11397 42070 11426
rect 42233 11445 42283 11474
rect 42233 11425 42250 11445
rect 42270 11425 42283 11445
rect 42233 11397 42283 11425
rect 40556 11288 40606 11301
rect 40764 11288 40814 11301
rect 40972 11288 41022 11301
rect 41185 11288 41235 11301
rect 41604 11284 41654 11297
rect 41812 11284 41862 11297
rect 42020 11284 42070 11297
rect 42233 11284 42283 11297
rect 934 10731 984 10744
rect 1147 10731 1197 10744
rect 1355 10731 1405 10744
rect 1563 10731 1613 10744
rect 1982 10727 2032 10740
rect 2195 10727 2245 10740
rect 2403 10727 2453 10740
rect 2611 10727 2661 10740
rect 934 10603 984 10631
rect 934 10583 947 10603
rect 967 10583 984 10603
rect 934 10554 984 10583
rect 1147 10602 1197 10631
rect 1147 10578 1158 10602
rect 1182 10578 1197 10602
rect 1147 10554 1197 10578
rect 1355 10607 1405 10631
rect 1355 10583 1367 10607
rect 1391 10583 1405 10607
rect 1355 10554 1405 10583
rect 1563 10605 1613 10631
rect 11642 10725 11692 10738
rect 11855 10725 11905 10738
rect 12063 10725 12113 10738
rect 12271 10725 12321 10738
rect 6686 10686 6736 10702
rect 6894 10686 6944 10702
rect 7102 10686 7152 10702
rect 7315 10686 7365 10702
rect 9224 10683 9274 10699
rect 9432 10683 9482 10699
rect 9640 10683 9690 10699
rect 9853 10683 9903 10699
rect 1563 10579 1581 10605
rect 1607 10579 1613 10605
rect 1563 10554 1613 10579
rect 1982 10599 2032 10627
rect 1982 10579 1995 10599
rect 2015 10579 2032 10599
rect 1982 10550 2032 10579
rect 2195 10598 2245 10627
rect 2195 10574 2206 10598
rect 2230 10574 2245 10598
rect 2195 10550 2245 10574
rect 2403 10603 2453 10627
rect 2403 10579 2415 10603
rect 2439 10579 2453 10603
rect 2403 10550 2453 10579
rect 2611 10601 2661 10627
rect 2611 10575 2629 10601
rect 2655 10575 2661 10601
rect 2611 10550 2661 10575
rect 6686 10619 6736 10644
rect 6686 10593 6692 10619
rect 6718 10593 6736 10619
rect 6686 10567 6736 10593
rect 6894 10615 6944 10644
rect 6894 10591 6908 10615
rect 6932 10591 6944 10615
rect 6894 10567 6944 10591
rect 7102 10620 7152 10644
rect 7102 10596 7117 10620
rect 7141 10596 7152 10620
rect 7102 10567 7152 10596
rect 7315 10615 7365 10644
rect 7315 10595 7332 10615
rect 7352 10595 7365 10615
rect 7315 10567 7365 10595
rect 9224 10616 9274 10641
rect 9224 10590 9230 10616
rect 9256 10590 9274 10616
rect 934 10496 984 10512
rect 1147 10496 1197 10512
rect 1355 10496 1405 10512
rect 1563 10496 1613 10512
rect 1982 10492 2032 10508
rect 2195 10492 2245 10508
rect 2403 10492 2453 10508
rect 2611 10492 2661 10508
rect 9224 10564 9274 10590
rect 9432 10612 9482 10641
rect 9432 10588 9446 10612
rect 9470 10588 9482 10612
rect 9432 10564 9482 10588
rect 9640 10617 9690 10641
rect 9640 10593 9655 10617
rect 9679 10593 9690 10617
rect 9640 10564 9690 10593
rect 9853 10612 9903 10641
rect 9853 10592 9870 10612
rect 9890 10592 9903 10612
rect 12690 10721 12740 10734
rect 12903 10721 12953 10734
rect 13111 10721 13161 10734
rect 13319 10721 13369 10734
rect 9853 10564 9903 10592
rect 6686 10454 6736 10467
rect 6894 10454 6944 10467
rect 7102 10454 7152 10467
rect 7315 10454 7365 10467
rect 11642 10597 11692 10625
rect 11642 10577 11655 10597
rect 11675 10577 11692 10597
rect 11642 10548 11692 10577
rect 11855 10596 11905 10625
rect 11855 10572 11866 10596
rect 11890 10572 11905 10596
rect 11855 10548 11905 10572
rect 12063 10601 12113 10625
rect 12063 10577 12075 10601
rect 12099 10577 12113 10601
rect 12063 10548 12113 10577
rect 12271 10599 12321 10625
rect 22607 10729 22657 10742
rect 22820 10729 22870 10742
rect 23028 10729 23078 10742
rect 23236 10729 23286 10742
rect 17394 10680 17444 10696
rect 17602 10680 17652 10696
rect 17810 10680 17860 10696
rect 18023 10680 18073 10696
rect 19932 10677 19982 10693
rect 20140 10677 20190 10693
rect 20348 10677 20398 10693
rect 20561 10677 20611 10693
rect 12271 10573 12289 10599
rect 12315 10573 12321 10599
rect 12271 10548 12321 10573
rect 12690 10593 12740 10621
rect 12690 10573 12703 10593
rect 12723 10573 12740 10593
rect 12690 10544 12740 10573
rect 12903 10592 12953 10621
rect 12903 10568 12914 10592
rect 12938 10568 12953 10592
rect 12903 10544 12953 10568
rect 13111 10597 13161 10621
rect 13111 10573 13123 10597
rect 13147 10573 13161 10597
rect 13111 10544 13161 10573
rect 13319 10595 13369 10621
rect 13319 10569 13337 10595
rect 13363 10569 13369 10595
rect 13319 10544 13369 10569
rect 17394 10613 17444 10638
rect 17394 10587 17400 10613
rect 17426 10587 17444 10613
rect 17394 10561 17444 10587
rect 17602 10609 17652 10638
rect 17602 10585 17616 10609
rect 17640 10585 17652 10609
rect 17602 10561 17652 10585
rect 17810 10614 17860 10638
rect 17810 10590 17825 10614
rect 17849 10590 17860 10614
rect 17810 10561 17860 10590
rect 18023 10609 18073 10638
rect 18023 10589 18040 10609
rect 18060 10589 18073 10609
rect 18023 10561 18073 10589
rect 19932 10610 19982 10635
rect 19932 10584 19938 10610
rect 19964 10584 19982 10610
rect 11642 10490 11692 10506
rect 11855 10490 11905 10506
rect 12063 10490 12113 10506
rect 12271 10490 12321 10506
rect 12690 10486 12740 10502
rect 12903 10486 12953 10502
rect 13111 10486 13161 10502
rect 13319 10486 13369 10502
rect 9224 10451 9274 10464
rect 9432 10451 9482 10464
rect 9640 10451 9690 10464
rect 9853 10451 9903 10464
rect 19932 10558 19982 10584
rect 20140 10606 20190 10635
rect 20140 10582 20154 10606
rect 20178 10582 20190 10606
rect 20140 10558 20190 10582
rect 20348 10611 20398 10635
rect 20348 10587 20363 10611
rect 20387 10587 20398 10611
rect 20348 10558 20398 10587
rect 20561 10606 20611 10635
rect 23655 10725 23705 10738
rect 23868 10725 23918 10738
rect 24076 10725 24126 10738
rect 24284 10725 24334 10738
rect 20561 10586 20578 10606
rect 20598 10586 20611 10606
rect 20561 10558 20611 10586
rect 17394 10448 17444 10461
rect 17602 10448 17652 10461
rect 17810 10448 17860 10461
rect 18023 10448 18073 10461
rect 22607 10601 22657 10629
rect 22607 10581 22620 10601
rect 22640 10581 22657 10601
rect 22607 10552 22657 10581
rect 22820 10600 22870 10629
rect 22820 10576 22831 10600
rect 22855 10576 22870 10600
rect 22820 10552 22870 10576
rect 23028 10605 23078 10629
rect 23028 10581 23040 10605
rect 23064 10581 23078 10605
rect 23028 10552 23078 10581
rect 23236 10603 23286 10629
rect 33315 10723 33365 10736
rect 33528 10723 33578 10736
rect 33736 10723 33786 10736
rect 33944 10723 33994 10736
rect 28359 10684 28409 10700
rect 28567 10684 28617 10700
rect 28775 10684 28825 10700
rect 28988 10684 29038 10700
rect 30897 10681 30947 10697
rect 31105 10681 31155 10697
rect 31313 10681 31363 10697
rect 31526 10681 31576 10697
rect 23236 10577 23254 10603
rect 23280 10577 23286 10603
rect 23236 10552 23286 10577
rect 23655 10597 23705 10625
rect 23655 10577 23668 10597
rect 23688 10577 23705 10597
rect 23655 10548 23705 10577
rect 23868 10596 23918 10625
rect 23868 10572 23879 10596
rect 23903 10572 23918 10596
rect 23868 10548 23918 10572
rect 24076 10601 24126 10625
rect 24076 10577 24088 10601
rect 24112 10577 24126 10601
rect 24076 10548 24126 10577
rect 24284 10599 24334 10625
rect 24284 10573 24302 10599
rect 24328 10573 24334 10599
rect 24284 10548 24334 10573
rect 28359 10617 28409 10642
rect 28359 10591 28365 10617
rect 28391 10591 28409 10617
rect 28359 10565 28409 10591
rect 28567 10613 28617 10642
rect 28567 10589 28581 10613
rect 28605 10589 28617 10613
rect 28567 10565 28617 10589
rect 28775 10618 28825 10642
rect 28775 10594 28790 10618
rect 28814 10594 28825 10618
rect 28775 10565 28825 10594
rect 28988 10613 29038 10642
rect 28988 10593 29005 10613
rect 29025 10593 29038 10613
rect 28988 10565 29038 10593
rect 30897 10614 30947 10639
rect 30897 10588 30903 10614
rect 30929 10588 30947 10614
rect 22607 10494 22657 10510
rect 22820 10494 22870 10510
rect 23028 10494 23078 10510
rect 23236 10494 23286 10510
rect 23655 10490 23705 10506
rect 23868 10490 23918 10506
rect 24076 10490 24126 10506
rect 24284 10490 24334 10506
rect 19932 10445 19982 10458
rect 20140 10445 20190 10458
rect 20348 10445 20398 10458
rect 20561 10445 20611 10458
rect 30897 10562 30947 10588
rect 31105 10610 31155 10639
rect 31105 10586 31119 10610
rect 31143 10586 31155 10610
rect 31105 10562 31155 10586
rect 31313 10615 31363 10639
rect 31313 10591 31328 10615
rect 31352 10591 31363 10615
rect 31313 10562 31363 10591
rect 31526 10610 31576 10639
rect 31526 10590 31543 10610
rect 31563 10590 31576 10610
rect 34363 10719 34413 10732
rect 34576 10719 34626 10732
rect 34784 10719 34834 10732
rect 34992 10719 35042 10732
rect 31526 10562 31576 10590
rect 28359 10452 28409 10465
rect 28567 10452 28617 10465
rect 28775 10452 28825 10465
rect 28988 10452 29038 10465
rect 33315 10595 33365 10623
rect 33315 10575 33328 10595
rect 33348 10575 33365 10595
rect 33315 10546 33365 10575
rect 33528 10594 33578 10623
rect 33528 10570 33539 10594
rect 33563 10570 33578 10594
rect 33528 10546 33578 10570
rect 33736 10599 33786 10623
rect 33736 10575 33748 10599
rect 33772 10575 33786 10599
rect 33736 10546 33786 10575
rect 33944 10597 33994 10623
rect 39067 10678 39117 10694
rect 39275 10678 39325 10694
rect 39483 10678 39533 10694
rect 39696 10678 39746 10694
rect 41605 10675 41655 10691
rect 41813 10675 41863 10691
rect 42021 10675 42071 10691
rect 42234 10675 42284 10691
rect 33944 10571 33962 10597
rect 33988 10571 33994 10597
rect 33944 10546 33994 10571
rect 34363 10591 34413 10619
rect 34363 10571 34376 10591
rect 34396 10571 34413 10591
rect 34363 10542 34413 10571
rect 34576 10590 34626 10619
rect 34576 10566 34587 10590
rect 34611 10566 34626 10590
rect 34576 10542 34626 10566
rect 34784 10595 34834 10619
rect 34784 10571 34796 10595
rect 34820 10571 34834 10595
rect 34784 10542 34834 10571
rect 34992 10593 35042 10619
rect 34992 10567 35010 10593
rect 35036 10567 35042 10593
rect 34992 10542 35042 10567
rect 39067 10611 39117 10636
rect 39067 10585 39073 10611
rect 39099 10585 39117 10611
rect 39067 10559 39117 10585
rect 39275 10607 39325 10636
rect 39275 10583 39289 10607
rect 39313 10583 39325 10607
rect 39275 10559 39325 10583
rect 39483 10612 39533 10636
rect 39483 10588 39498 10612
rect 39522 10588 39533 10612
rect 39483 10559 39533 10588
rect 39696 10607 39746 10636
rect 39696 10587 39713 10607
rect 39733 10587 39746 10607
rect 39696 10559 39746 10587
rect 41605 10608 41655 10633
rect 41605 10582 41611 10608
rect 41637 10582 41655 10608
rect 33315 10488 33365 10504
rect 33528 10488 33578 10504
rect 33736 10488 33786 10504
rect 33944 10488 33994 10504
rect 34363 10484 34413 10500
rect 34576 10484 34626 10500
rect 34784 10484 34834 10500
rect 34992 10484 35042 10500
rect 30897 10449 30947 10462
rect 31105 10449 31155 10462
rect 31313 10449 31363 10462
rect 31526 10449 31576 10462
rect 41605 10556 41655 10582
rect 41813 10604 41863 10633
rect 41813 10580 41827 10604
rect 41851 10580 41863 10604
rect 41813 10556 41863 10580
rect 42021 10609 42071 10633
rect 42021 10585 42036 10609
rect 42060 10585 42071 10609
rect 42021 10556 42071 10585
rect 42234 10604 42284 10633
rect 42234 10584 42251 10604
rect 42271 10584 42284 10604
rect 42234 10556 42284 10584
rect 39067 10446 39117 10459
rect 39275 10446 39325 10459
rect 39483 10446 39533 10459
rect 39696 10446 39746 10459
rect 41605 10443 41655 10456
rect 41813 10443 41863 10456
rect 42021 10443 42071 10456
rect 42234 10443 42284 10456
rect 934 10052 984 10065
rect 1147 10052 1197 10065
rect 1355 10052 1405 10065
rect 1563 10052 1613 10065
rect 3429 10047 3479 10060
rect 3642 10047 3692 10060
rect 3850 10047 3900 10060
rect 4058 10047 4108 10060
rect 934 9924 984 9952
rect 934 9904 947 9924
rect 967 9904 984 9924
rect 934 9875 984 9904
rect 1147 9923 1197 9952
rect 1147 9899 1158 9923
rect 1182 9899 1197 9923
rect 1147 9875 1197 9899
rect 1355 9928 1405 9952
rect 1355 9904 1367 9928
rect 1391 9904 1405 9928
rect 1355 9875 1405 9904
rect 1563 9926 1613 9952
rect 11642 10046 11692 10059
rect 11855 10046 11905 10059
rect 12063 10046 12113 10059
rect 12271 10046 12321 10059
rect 8176 10008 8226 10024
rect 8384 10008 8434 10024
rect 8592 10008 8642 10024
rect 8805 10008 8855 10024
rect 9224 10004 9274 10020
rect 9432 10004 9482 10020
rect 9640 10004 9690 10020
rect 9853 10004 9903 10020
rect 1563 9900 1581 9926
rect 1607 9900 1613 9926
rect 1563 9875 1613 9900
rect 3429 9919 3479 9947
rect 3429 9899 3442 9919
rect 3462 9899 3479 9919
rect 3429 9870 3479 9899
rect 3642 9918 3692 9947
rect 3642 9894 3653 9918
rect 3677 9894 3692 9918
rect 3642 9870 3692 9894
rect 3850 9923 3900 9947
rect 3850 9899 3862 9923
rect 3886 9899 3900 9923
rect 3850 9870 3900 9899
rect 4058 9921 4108 9947
rect 4058 9895 4076 9921
rect 4102 9895 4108 9921
rect 4058 9870 4108 9895
rect 8176 9941 8226 9966
rect 8176 9915 8182 9941
rect 8208 9915 8226 9941
rect 8176 9889 8226 9915
rect 8384 9937 8434 9966
rect 8384 9913 8398 9937
rect 8422 9913 8434 9937
rect 8384 9889 8434 9913
rect 8592 9942 8642 9966
rect 8592 9918 8607 9942
rect 8631 9918 8642 9942
rect 8592 9889 8642 9918
rect 8805 9937 8855 9966
rect 8805 9917 8822 9937
rect 8842 9917 8855 9937
rect 8805 9889 8855 9917
rect 9224 9937 9274 9962
rect 9224 9911 9230 9937
rect 9256 9911 9274 9937
rect 934 9817 984 9833
rect 1147 9817 1197 9833
rect 1355 9817 1405 9833
rect 1563 9817 1613 9833
rect 3429 9812 3479 9828
rect 3642 9812 3692 9828
rect 3850 9812 3900 9828
rect 4058 9812 4108 9828
rect 9224 9885 9274 9911
rect 9432 9933 9482 9962
rect 9432 9909 9446 9933
rect 9470 9909 9482 9933
rect 9432 9885 9482 9909
rect 9640 9938 9690 9962
rect 9640 9914 9655 9938
rect 9679 9914 9690 9938
rect 9640 9885 9690 9914
rect 9853 9933 9903 9962
rect 9853 9913 9870 9933
rect 9890 9913 9903 9933
rect 9853 9885 9903 9913
rect 14137 10041 14187 10054
rect 14350 10041 14400 10054
rect 14558 10041 14608 10054
rect 14766 10041 14816 10054
rect 11642 9918 11692 9946
rect 8176 9776 8226 9789
rect 8384 9776 8434 9789
rect 8592 9776 8642 9789
rect 8805 9776 8855 9789
rect 11642 9898 11655 9918
rect 11675 9898 11692 9918
rect 11642 9869 11692 9898
rect 11855 9917 11905 9946
rect 11855 9893 11866 9917
rect 11890 9893 11905 9917
rect 11855 9869 11905 9893
rect 12063 9922 12113 9946
rect 12063 9898 12075 9922
rect 12099 9898 12113 9922
rect 12063 9869 12113 9898
rect 12271 9920 12321 9946
rect 22607 10050 22657 10063
rect 22820 10050 22870 10063
rect 23028 10050 23078 10063
rect 23236 10050 23286 10063
rect 18884 10002 18934 10018
rect 19092 10002 19142 10018
rect 19300 10002 19350 10018
rect 19513 10002 19563 10018
rect 19932 9998 19982 10014
rect 20140 9998 20190 10014
rect 20348 9998 20398 10014
rect 20561 9998 20611 10014
rect 12271 9894 12289 9920
rect 12315 9894 12321 9920
rect 12271 9869 12321 9894
rect 14137 9913 14187 9941
rect 14137 9893 14150 9913
rect 14170 9893 14187 9913
rect 14137 9864 14187 9893
rect 14350 9912 14400 9941
rect 14350 9888 14361 9912
rect 14385 9888 14400 9912
rect 14350 9864 14400 9888
rect 14558 9917 14608 9941
rect 14558 9893 14570 9917
rect 14594 9893 14608 9917
rect 14558 9864 14608 9893
rect 14766 9915 14816 9941
rect 14766 9889 14784 9915
rect 14810 9889 14816 9915
rect 14766 9864 14816 9889
rect 18884 9935 18934 9960
rect 18884 9909 18890 9935
rect 18916 9909 18934 9935
rect 18884 9883 18934 9909
rect 19092 9931 19142 9960
rect 19092 9907 19106 9931
rect 19130 9907 19142 9931
rect 19092 9883 19142 9907
rect 19300 9936 19350 9960
rect 19300 9912 19315 9936
rect 19339 9912 19350 9936
rect 19300 9883 19350 9912
rect 19513 9931 19563 9960
rect 19513 9911 19530 9931
rect 19550 9911 19563 9931
rect 19513 9883 19563 9911
rect 19932 9931 19982 9956
rect 19932 9905 19938 9931
rect 19964 9905 19982 9931
rect 11642 9811 11692 9827
rect 11855 9811 11905 9827
rect 12063 9811 12113 9827
rect 12271 9811 12321 9827
rect 14137 9806 14187 9822
rect 14350 9806 14400 9822
rect 14558 9806 14608 9822
rect 14766 9806 14816 9822
rect 9224 9772 9274 9785
rect 9432 9772 9482 9785
rect 9640 9772 9690 9785
rect 9853 9772 9903 9785
rect 19932 9879 19982 9905
rect 20140 9927 20190 9956
rect 20140 9903 20154 9927
rect 20178 9903 20190 9927
rect 20140 9879 20190 9903
rect 20348 9932 20398 9956
rect 20348 9908 20363 9932
rect 20387 9908 20398 9932
rect 20348 9879 20398 9908
rect 20561 9927 20611 9956
rect 20561 9907 20578 9927
rect 20598 9907 20611 9927
rect 20561 9879 20611 9907
rect 25102 10045 25152 10058
rect 25315 10045 25365 10058
rect 25523 10045 25573 10058
rect 25731 10045 25781 10058
rect 22607 9922 22657 9950
rect 22607 9902 22620 9922
rect 22640 9902 22657 9922
rect 18884 9770 18934 9783
rect 19092 9770 19142 9783
rect 19300 9770 19350 9783
rect 19513 9770 19563 9783
rect 22607 9873 22657 9902
rect 22820 9921 22870 9950
rect 22820 9897 22831 9921
rect 22855 9897 22870 9921
rect 22820 9873 22870 9897
rect 23028 9926 23078 9950
rect 23028 9902 23040 9926
rect 23064 9902 23078 9926
rect 23028 9873 23078 9902
rect 23236 9924 23286 9950
rect 33315 10044 33365 10057
rect 33528 10044 33578 10057
rect 33736 10044 33786 10057
rect 33944 10044 33994 10057
rect 29849 10006 29899 10022
rect 30057 10006 30107 10022
rect 30265 10006 30315 10022
rect 30478 10006 30528 10022
rect 30897 10002 30947 10018
rect 31105 10002 31155 10018
rect 31313 10002 31363 10018
rect 31526 10002 31576 10018
rect 23236 9898 23254 9924
rect 23280 9898 23286 9924
rect 23236 9873 23286 9898
rect 25102 9917 25152 9945
rect 25102 9897 25115 9917
rect 25135 9897 25152 9917
rect 25102 9868 25152 9897
rect 25315 9916 25365 9945
rect 25315 9892 25326 9916
rect 25350 9892 25365 9916
rect 25315 9868 25365 9892
rect 25523 9921 25573 9945
rect 25523 9897 25535 9921
rect 25559 9897 25573 9921
rect 25523 9868 25573 9897
rect 25731 9919 25781 9945
rect 25731 9893 25749 9919
rect 25775 9893 25781 9919
rect 25731 9868 25781 9893
rect 29849 9939 29899 9964
rect 29849 9913 29855 9939
rect 29881 9913 29899 9939
rect 29849 9887 29899 9913
rect 30057 9935 30107 9964
rect 30057 9911 30071 9935
rect 30095 9911 30107 9935
rect 30057 9887 30107 9911
rect 30265 9940 30315 9964
rect 30265 9916 30280 9940
rect 30304 9916 30315 9940
rect 30265 9887 30315 9916
rect 30478 9935 30528 9964
rect 30478 9915 30495 9935
rect 30515 9915 30528 9935
rect 30478 9887 30528 9915
rect 30897 9935 30947 9960
rect 30897 9909 30903 9935
rect 30929 9909 30947 9935
rect 22607 9815 22657 9831
rect 22820 9815 22870 9831
rect 23028 9815 23078 9831
rect 23236 9815 23286 9831
rect 25102 9810 25152 9826
rect 25315 9810 25365 9826
rect 25523 9810 25573 9826
rect 25731 9810 25781 9826
rect 19932 9766 19982 9779
rect 20140 9766 20190 9779
rect 20348 9766 20398 9779
rect 20561 9766 20611 9779
rect 30897 9883 30947 9909
rect 31105 9931 31155 9960
rect 31105 9907 31119 9931
rect 31143 9907 31155 9931
rect 31105 9883 31155 9907
rect 31313 9936 31363 9960
rect 31313 9912 31328 9936
rect 31352 9912 31363 9936
rect 31313 9883 31363 9912
rect 31526 9931 31576 9960
rect 31526 9911 31543 9931
rect 31563 9911 31576 9931
rect 31526 9883 31576 9911
rect 35810 10039 35860 10052
rect 36023 10039 36073 10052
rect 36231 10039 36281 10052
rect 36439 10039 36489 10052
rect 33315 9916 33365 9944
rect 29849 9774 29899 9787
rect 30057 9774 30107 9787
rect 30265 9774 30315 9787
rect 30478 9774 30528 9787
rect 33315 9896 33328 9916
rect 33348 9896 33365 9916
rect 33315 9867 33365 9896
rect 33528 9915 33578 9944
rect 33528 9891 33539 9915
rect 33563 9891 33578 9915
rect 33528 9867 33578 9891
rect 33736 9920 33786 9944
rect 33736 9896 33748 9920
rect 33772 9896 33786 9920
rect 33736 9867 33786 9896
rect 33944 9918 33994 9944
rect 40557 10000 40607 10016
rect 40765 10000 40815 10016
rect 40973 10000 41023 10016
rect 41186 10000 41236 10016
rect 41605 9996 41655 10012
rect 41813 9996 41863 10012
rect 42021 9996 42071 10012
rect 42234 9996 42284 10012
rect 33944 9892 33962 9918
rect 33988 9892 33994 9918
rect 33944 9867 33994 9892
rect 35810 9911 35860 9939
rect 35810 9891 35823 9911
rect 35843 9891 35860 9911
rect 35810 9862 35860 9891
rect 36023 9910 36073 9939
rect 36023 9886 36034 9910
rect 36058 9886 36073 9910
rect 36023 9862 36073 9886
rect 36231 9915 36281 9939
rect 36231 9891 36243 9915
rect 36267 9891 36281 9915
rect 36231 9862 36281 9891
rect 36439 9913 36489 9939
rect 36439 9887 36457 9913
rect 36483 9887 36489 9913
rect 36439 9862 36489 9887
rect 40557 9933 40607 9958
rect 40557 9907 40563 9933
rect 40589 9907 40607 9933
rect 40557 9881 40607 9907
rect 40765 9929 40815 9958
rect 40765 9905 40779 9929
rect 40803 9905 40815 9929
rect 40765 9881 40815 9905
rect 40973 9934 41023 9958
rect 40973 9910 40988 9934
rect 41012 9910 41023 9934
rect 40973 9881 41023 9910
rect 41186 9929 41236 9958
rect 41186 9909 41203 9929
rect 41223 9909 41236 9929
rect 41186 9881 41236 9909
rect 41605 9929 41655 9954
rect 41605 9903 41611 9929
rect 41637 9903 41655 9929
rect 33315 9809 33365 9825
rect 33528 9809 33578 9825
rect 33736 9809 33786 9825
rect 33944 9809 33994 9825
rect 35810 9804 35860 9820
rect 36023 9804 36073 9820
rect 36231 9804 36281 9820
rect 36439 9804 36489 9820
rect 30897 9770 30947 9783
rect 31105 9770 31155 9783
rect 31313 9770 31363 9783
rect 31526 9770 31576 9783
rect 41605 9877 41655 9903
rect 41813 9925 41863 9954
rect 41813 9901 41827 9925
rect 41851 9901 41863 9925
rect 41813 9877 41863 9901
rect 42021 9930 42071 9954
rect 42021 9906 42036 9930
rect 42060 9906 42071 9930
rect 42021 9877 42071 9906
rect 42234 9925 42284 9954
rect 42234 9905 42251 9925
rect 42271 9905 42284 9925
rect 42234 9877 42284 9905
rect 40557 9768 40607 9781
rect 40765 9768 40815 9781
rect 40973 9768 41023 9781
rect 41186 9768 41236 9781
rect 41605 9764 41655 9777
rect 41813 9764 41863 9777
rect 42021 9764 42071 9777
rect 42234 9764 42284 9777
rect 934 9284 984 9297
rect 1147 9284 1197 9297
rect 1355 9284 1405 9297
rect 1563 9284 1613 9297
rect 1982 9280 2032 9293
rect 2195 9280 2245 9293
rect 2403 9280 2453 9293
rect 2611 9280 2661 9293
rect 934 9156 984 9184
rect 934 9136 947 9156
rect 967 9136 984 9156
rect 934 9107 984 9136
rect 1147 9155 1197 9184
rect 1147 9131 1158 9155
rect 1182 9131 1197 9155
rect 1147 9107 1197 9131
rect 1355 9160 1405 9184
rect 1355 9136 1367 9160
rect 1391 9136 1405 9160
rect 1355 9107 1405 9136
rect 1563 9158 1613 9184
rect 11642 9278 11692 9291
rect 11855 9278 11905 9291
rect 12063 9278 12113 9291
rect 12271 9278 12321 9291
rect 6729 9241 6779 9257
rect 6937 9241 6987 9257
rect 7145 9241 7195 9257
rect 7358 9241 7408 9257
rect 9224 9236 9274 9252
rect 9432 9236 9482 9252
rect 9640 9236 9690 9252
rect 9853 9236 9903 9252
rect 1563 9132 1581 9158
rect 1607 9132 1613 9158
rect 1563 9107 1613 9132
rect 1982 9152 2032 9180
rect 1982 9132 1995 9152
rect 2015 9132 2032 9152
rect 1982 9103 2032 9132
rect 2195 9151 2245 9180
rect 2195 9127 2206 9151
rect 2230 9127 2245 9151
rect 2195 9103 2245 9127
rect 2403 9156 2453 9180
rect 2403 9132 2415 9156
rect 2439 9132 2453 9156
rect 2403 9103 2453 9132
rect 2611 9154 2661 9180
rect 2611 9128 2629 9154
rect 2655 9128 2661 9154
rect 2611 9103 2661 9128
rect 6729 9174 6779 9199
rect 6729 9148 6735 9174
rect 6761 9148 6779 9174
rect 6729 9122 6779 9148
rect 6937 9170 6987 9199
rect 6937 9146 6951 9170
rect 6975 9146 6987 9170
rect 6937 9122 6987 9146
rect 7145 9175 7195 9199
rect 7145 9151 7160 9175
rect 7184 9151 7195 9175
rect 7145 9122 7195 9151
rect 7358 9170 7408 9199
rect 7358 9150 7375 9170
rect 7395 9150 7408 9170
rect 7358 9122 7408 9150
rect 9224 9169 9274 9194
rect 9224 9143 9230 9169
rect 9256 9143 9274 9169
rect 934 9049 984 9065
rect 1147 9049 1197 9065
rect 1355 9049 1405 9065
rect 1563 9049 1613 9065
rect 1982 9045 2032 9061
rect 2195 9045 2245 9061
rect 2403 9045 2453 9061
rect 2611 9045 2661 9061
rect 9224 9117 9274 9143
rect 9432 9165 9482 9194
rect 9432 9141 9446 9165
rect 9470 9141 9482 9165
rect 9432 9117 9482 9141
rect 9640 9170 9690 9194
rect 9640 9146 9655 9170
rect 9679 9146 9690 9170
rect 9640 9117 9690 9146
rect 9853 9165 9903 9194
rect 9853 9145 9870 9165
rect 9890 9145 9903 9165
rect 12690 9274 12740 9287
rect 12903 9274 12953 9287
rect 13111 9274 13161 9287
rect 13319 9274 13369 9287
rect 9853 9117 9903 9145
rect 6729 9009 6779 9022
rect 6937 9009 6987 9022
rect 7145 9009 7195 9022
rect 7358 9009 7408 9022
rect 11642 9150 11692 9178
rect 11642 9130 11655 9150
rect 11675 9130 11692 9150
rect 11642 9101 11692 9130
rect 11855 9149 11905 9178
rect 11855 9125 11866 9149
rect 11890 9125 11905 9149
rect 11855 9101 11905 9125
rect 12063 9154 12113 9178
rect 12063 9130 12075 9154
rect 12099 9130 12113 9154
rect 12063 9101 12113 9130
rect 12271 9152 12321 9178
rect 22607 9282 22657 9295
rect 22820 9282 22870 9295
rect 23028 9282 23078 9295
rect 23236 9282 23286 9295
rect 17437 9235 17487 9251
rect 17645 9235 17695 9251
rect 17853 9235 17903 9251
rect 18066 9235 18116 9251
rect 19932 9230 19982 9246
rect 20140 9230 20190 9246
rect 20348 9230 20398 9246
rect 20561 9230 20611 9246
rect 12271 9126 12289 9152
rect 12315 9126 12321 9152
rect 12271 9101 12321 9126
rect 12690 9146 12740 9174
rect 12690 9126 12703 9146
rect 12723 9126 12740 9146
rect 12690 9097 12740 9126
rect 12903 9145 12953 9174
rect 12903 9121 12914 9145
rect 12938 9121 12953 9145
rect 12903 9097 12953 9121
rect 13111 9150 13161 9174
rect 13111 9126 13123 9150
rect 13147 9126 13161 9150
rect 13111 9097 13161 9126
rect 13319 9148 13369 9174
rect 13319 9122 13337 9148
rect 13363 9122 13369 9148
rect 13319 9097 13369 9122
rect 17437 9168 17487 9193
rect 17437 9142 17443 9168
rect 17469 9142 17487 9168
rect 17437 9116 17487 9142
rect 17645 9164 17695 9193
rect 17645 9140 17659 9164
rect 17683 9140 17695 9164
rect 17645 9116 17695 9140
rect 17853 9169 17903 9193
rect 17853 9145 17868 9169
rect 17892 9145 17903 9169
rect 17853 9116 17903 9145
rect 18066 9164 18116 9193
rect 18066 9144 18083 9164
rect 18103 9144 18116 9164
rect 18066 9116 18116 9144
rect 19932 9163 19982 9188
rect 19932 9137 19938 9163
rect 19964 9137 19982 9163
rect 11642 9043 11692 9059
rect 11855 9043 11905 9059
rect 12063 9043 12113 9059
rect 12271 9043 12321 9059
rect 12690 9039 12740 9055
rect 12903 9039 12953 9055
rect 13111 9039 13161 9055
rect 13319 9039 13369 9055
rect 9224 9004 9274 9017
rect 9432 9004 9482 9017
rect 9640 9004 9690 9017
rect 9853 9004 9903 9017
rect 19932 9111 19982 9137
rect 20140 9159 20190 9188
rect 20140 9135 20154 9159
rect 20178 9135 20190 9159
rect 20140 9111 20190 9135
rect 20348 9164 20398 9188
rect 20348 9140 20363 9164
rect 20387 9140 20398 9164
rect 20348 9111 20398 9140
rect 20561 9159 20611 9188
rect 23655 9278 23705 9291
rect 23868 9278 23918 9291
rect 24076 9278 24126 9291
rect 24284 9278 24334 9291
rect 20561 9139 20578 9159
rect 20598 9139 20611 9159
rect 20561 9111 20611 9139
rect 17437 9003 17487 9016
rect 17645 9003 17695 9016
rect 17853 9003 17903 9016
rect 18066 9003 18116 9016
rect 22607 9154 22657 9182
rect 22607 9134 22620 9154
rect 22640 9134 22657 9154
rect 22607 9105 22657 9134
rect 22820 9153 22870 9182
rect 22820 9129 22831 9153
rect 22855 9129 22870 9153
rect 22820 9105 22870 9129
rect 23028 9158 23078 9182
rect 23028 9134 23040 9158
rect 23064 9134 23078 9158
rect 23028 9105 23078 9134
rect 23236 9156 23286 9182
rect 33315 9276 33365 9289
rect 33528 9276 33578 9289
rect 33736 9276 33786 9289
rect 33944 9276 33994 9289
rect 28402 9239 28452 9255
rect 28610 9239 28660 9255
rect 28818 9239 28868 9255
rect 29031 9239 29081 9255
rect 30897 9234 30947 9250
rect 31105 9234 31155 9250
rect 31313 9234 31363 9250
rect 31526 9234 31576 9250
rect 23236 9130 23254 9156
rect 23280 9130 23286 9156
rect 23236 9105 23286 9130
rect 23655 9150 23705 9178
rect 23655 9130 23668 9150
rect 23688 9130 23705 9150
rect 23655 9101 23705 9130
rect 23868 9149 23918 9178
rect 23868 9125 23879 9149
rect 23903 9125 23918 9149
rect 23868 9101 23918 9125
rect 24076 9154 24126 9178
rect 24076 9130 24088 9154
rect 24112 9130 24126 9154
rect 24076 9101 24126 9130
rect 24284 9152 24334 9178
rect 24284 9126 24302 9152
rect 24328 9126 24334 9152
rect 24284 9101 24334 9126
rect 28402 9172 28452 9197
rect 28402 9146 28408 9172
rect 28434 9146 28452 9172
rect 28402 9120 28452 9146
rect 28610 9168 28660 9197
rect 28610 9144 28624 9168
rect 28648 9144 28660 9168
rect 28610 9120 28660 9144
rect 28818 9173 28868 9197
rect 28818 9149 28833 9173
rect 28857 9149 28868 9173
rect 28818 9120 28868 9149
rect 29031 9168 29081 9197
rect 29031 9148 29048 9168
rect 29068 9148 29081 9168
rect 29031 9120 29081 9148
rect 30897 9167 30947 9192
rect 30897 9141 30903 9167
rect 30929 9141 30947 9167
rect 22607 9047 22657 9063
rect 22820 9047 22870 9063
rect 23028 9047 23078 9063
rect 23236 9047 23286 9063
rect 23655 9043 23705 9059
rect 23868 9043 23918 9059
rect 24076 9043 24126 9059
rect 24284 9043 24334 9059
rect 19932 8998 19982 9011
rect 20140 8998 20190 9011
rect 20348 8998 20398 9011
rect 20561 8998 20611 9011
rect 30897 9115 30947 9141
rect 31105 9163 31155 9192
rect 31105 9139 31119 9163
rect 31143 9139 31155 9163
rect 31105 9115 31155 9139
rect 31313 9168 31363 9192
rect 31313 9144 31328 9168
rect 31352 9144 31363 9168
rect 31313 9115 31363 9144
rect 31526 9163 31576 9192
rect 31526 9143 31543 9163
rect 31563 9143 31576 9163
rect 34363 9272 34413 9285
rect 34576 9272 34626 9285
rect 34784 9272 34834 9285
rect 34992 9272 35042 9285
rect 31526 9115 31576 9143
rect 28402 9007 28452 9020
rect 28610 9007 28660 9020
rect 28818 9007 28868 9020
rect 29031 9007 29081 9020
rect 33315 9148 33365 9176
rect 33315 9128 33328 9148
rect 33348 9128 33365 9148
rect 33315 9099 33365 9128
rect 33528 9147 33578 9176
rect 33528 9123 33539 9147
rect 33563 9123 33578 9147
rect 33528 9099 33578 9123
rect 33736 9152 33786 9176
rect 33736 9128 33748 9152
rect 33772 9128 33786 9152
rect 33736 9099 33786 9128
rect 33944 9150 33994 9176
rect 39110 9233 39160 9249
rect 39318 9233 39368 9249
rect 39526 9233 39576 9249
rect 39739 9233 39789 9249
rect 41605 9228 41655 9244
rect 41813 9228 41863 9244
rect 42021 9228 42071 9244
rect 42234 9228 42284 9244
rect 33944 9124 33962 9150
rect 33988 9124 33994 9150
rect 33944 9099 33994 9124
rect 34363 9144 34413 9172
rect 34363 9124 34376 9144
rect 34396 9124 34413 9144
rect 34363 9095 34413 9124
rect 34576 9143 34626 9172
rect 34576 9119 34587 9143
rect 34611 9119 34626 9143
rect 34576 9095 34626 9119
rect 34784 9148 34834 9172
rect 34784 9124 34796 9148
rect 34820 9124 34834 9148
rect 34784 9095 34834 9124
rect 34992 9146 35042 9172
rect 34992 9120 35010 9146
rect 35036 9120 35042 9146
rect 34992 9095 35042 9120
rect 39110 9166 39160 9191
rect 39110 9140 39116 9166
rect 39142 9140 39160 9166
rect 39110 9114 39160 9140
rect 39318 9162 39368 9191
rect 39318 9138 39332 9162
rect 39356 9138 39368 9162
rect 39318 9114 39368 9138
rect 39526 9167 39576 9191
rect 39526 9143 39541 9167
rect 39565 9143 39576 9167
rect 39526 9114 39576 9143
rect 39739 9162 39789 9191
rect 39739 9142 39756 9162
rect 39776 9142 39789 9162
rect 39739 9114 39789 9142
rect 41605 9161 41655 9186
rect 41605 9135 41611 9161
rect 41637 9135 41655 9161
rect 33315 9041 33365 9057
rect 33528 9041 33578 9057
rect 33736 9041 33786 9057
rect 33944 9041 33994 9057
rect 34363 9037 34413 9053
rect 34576 9037 34626 9053
rect 34784 9037 34834 9053
rect 34992 9037 35042 9053
rect 30897 9002 30947 9015
rect 31105 9002 31155 9015
rect 31313 9002 31363 9015
rect 31526 9002 31576 9015
rect 41605 9109 41655 9135
rect 41813 9157 41863 9186
rect 41813 9133 41827 9157
rect 41851 9133 41863 9157
rect 41813 9109 41863 9133
rect 42021 9162 42071 9186
rect 42021 9138 42036 9162
rect 42060 9138 42071 9162
rect 42021 9109 42071 9138
rect 42234 9157 42284 9186
rect 42234 9137 42251 9157
rect 42271 9137 42284 9157
rect 42234 9109 42284 9137
rect 39110 9001 39160 9014
rect 39318 9001 39368 9014
rect 39526 9001 39576 9014
rect 39739 9001 39789 9014
rect 41605 8996 41655 9009
rect 41813 8996 41863 9009
rect 42021 8996 42071 9009
rect 42234 8996 42284 9009
rect 934 8605 984 8618
rect 1147 8605 1197 8618
rect 1355 8605 1405 8618
rect 1563 8605 1613 8618
rect 4537 8596 4587 8609
rect 4750 8596 4800 8609
rect 4958 8596 5008 8609
rect 5166 8596 5216 8609
rect 11642 8599 11692 8612
rect 11855 8599 11905 8612
rect 12063 8599 12113 8612
rect 12271 8599 12321 8612
rect 934 8477 984 8505
rect 934 8457 947 8477
rect 967 8457 984 8477
rect 934 8428 984 8457
rect 1147 8476 1197 8505
rect 1147 8452 1158 8476
rect 1182 8452 1197 8476
rect 1147 8428 1197 8452
rect 1355 8481 1405 8505
rect 1355 8457 1367 8481
rect 1391 8457 1405 8481
rect 1355 8428 1405 8457
rect 1563 8479 1613 8505
rect 8176 8561 8226 8577
rect 8384 8561 8434 8577
rect 8592 8561 8642 8577
rect 8805 8561 8855 8577
rect 9224 8557 9274 8573
rect 9432 8557 9482 8573
rect 9640 8557 9690 8573
rect 9853 8557 9903 8573
rect 1563 8453 1581 8479
rect 1607 8453 1613 8479
rect 1563 8428 1613 8453
rect 4537 8468 4587 8496
rect 4537 8448 4550 8468
rect 4570 8448 4587 8468
rect 4537 8419 4587 8448
rect 4750 8467 4800 8496
rect 4750 8443 4761 8467
rect 4785 8443 4800 8467
rect 4750 8419 4800 8443
rect 4958 8472 5008 8496
rect 4958 8448 4970 8472
rect 4994 8448 5008 8472
rect 4958 8419 5008 8448
rect 5166 8470 5216 8496
rect 5166 8444 5184 8470
rect 5210 8444 5216 8470
rect 5166 8419 5216 8444
rect 8176 8494 8226 8519
rect 8176 8468 8182 8494
rect 8208 8468 8226 8494
rect 8176 8442 8226 8468
rect 8384 8490 8434 8519
rect 8384 8466 8398 8490
rect 8422 8466 8434 8490
rect 8384 8442 8434 8466
rect 8592 8495 8642 8519
rect 8592 8471 8607 8495
rect 8631 8471 8642 8495
rect 8592 8442 8642 8471
rect 8805 8490 8855 8519
rect 8805 8470 8822 8490
rect 8842 8470 8855 8490
rect 8805 8442 8855 8470
rect 9224 8490 9274 8515
rect 9224 8464 9230 8490
rect 9256 8464 9274 8490
rect 934 8370 984 8386
rect 1147 8370 1197 8386
rect 1355 8370 1405 8386
rect 1563 8370 1613 8386
rect 4537 8361 4587 8377
rect 4750 8361 4800 8377
rect 4958 8361 5008 8377
rect 5166 8361 5216 8377
rect 9224 8438 9274 8464
rect 9432 8486 9482 8515
rect 9432 8462 9446 8486
rect 9470 8462 9482 8486
rect 9432 8438 9482 8462
rect 9640 8491 9690 8515
rect 9640 8467 9655 8491
rect 9679 8467 9690 8491
rect 9640 8438 9690 8467
rect 9853 8486 9903 8515
rect 9853 8466 9870 8486
rect 9890 8466 9903 8486
rect 9853 8438 9903 8466
rect 15245 8590 15295 8603
rect 15458 8590 15508 8603
rect 15666 8590 15716 8603
rect 15874 8590 15924 8603
rect 22607 8603 22657 8616
rect 22820 8603 22870 8616
rect 23028 8603 23078 8616
rect 23236 8603 23286 8616
rect 11642 8471 11692 8499
rect 8176 8329 8226 8342
rect 8384 8329 8434 8342
rect 8592 8329 8642 8342
rect 8805 8329 8855 8342
rect 11642 8451 11655 8471
rect 11675 8451 11692 8471
rect 11642 8422 11692 8451
rect 11855 8470 11905 8499
rect 11855 8446 11866 8470
rect 11890 8446 11905 8470
rect 11855 8422 11905 8446
rect 12063 8475 12113 8499
rect 12063 8451 12075 8475
rect 12099 8451 12113 8475
rect 12063 8422 12113 8451
rect 12271 8473 12321 8499
rect 18884 8555 18934 8571
rect 19092 8555 19142 8571
rect 19300 8555 19350 8571
rect 19513 8555 19563 8571
rect 19932 8551 19982 8567
rect 20140 8551 20190 8567
rect 20348 8551 20398 8567
rect 20561 8551 20611 8567
rect 12271 8447 12289 8473
rect 12315 8447 12321 8473
rect 12271 8422 12321 8447
rect 15245 8462 15295 8490
rect 15245 8442 15258 8462
rect 15278 8442 15295 8462
rect 15245 8413 15295 8442
rect 15458 8461 15508 8490
rect 15458 8437 15469 8461
rect 15493 8437 15508 8461
rect 15458 8413 15508 8437
rect 15666 8466 15716 8490
rect 15666 8442 15678 8466
rect 15702 8442 15716 8466
rect 15666 8413 15716 8442
rect 15874 8464 15924 8490
rect 15874 8438 15892 8464
rect 15918 8438 15924 8464
rect 15874 8413 15924 8438
rect 18884 8488 18934 8513
rect 18884 8462 18890 8488
rect 18916 8462 18934 8488
rect 18884 8436 18934 8462
rect 19092 8484 19142 8513
rect 19092 8460 19106 8484
rect 19130 8460 19142 8484
rect 19092 8436 19142 8460
rect 19300 8489 19350 8513
rect 19300 8465 19315 8489
rect 19339 8465 19350 8489
rect 19300 8436 19350 8465
rect 19513 8484 19563 8513
rect 19513 8464 19530 8484
rect 19550 8464 19563 8484
rect 19513 8436 19563 8464
rect 19932 8484 19982 8509
rect 19932 8458 19938 8484
rect 19964 8458 19982 8484
rect 11642 8364 11692 8380
rect 11855 8364 11905 8380
rect 12063 8364 12113 8380
rect 12271 8364 12321 8380
rect 15245 8355 15295 8371
rect 15458 8355 15508 8371
rect 15666 8355 15716 8371
rect 15874 8355 15924 8371
rect 9224 8325 9274 8338
rect 9432 8325 9482 8338
rect 9640 8325 9690 8338
rect 9853 8325 9903 8338
rect 19932 8432 19982 8458
rect 20140 8480 20190 8509
rect 20140 8456 20154 8480
rect 20178 8456 20190 8480
rect 20140 8432 20190 8456
rect 20348 8485 20398 8509
rect 20348 8461 20363 8485
rect 20387 8461 20398 8485
rect 20348 8432 20398 8461
rect 20561 8480 20611 8509
rect 20561 8460 20578 8480
rect 20598 8460 20611 8480
rect 20561 8432 20611 8460
rect 26210 8594 26260 8607
rect 26423 8594 26473 8607
rect 26631 8594 26681 8607
rect 26839 8594 26889 8607
rect 33315 8597 33365 8610
rect 33528 8597 33578 8610
rect 33736 8597 33786 8610
rect 33944 8597 33994 8610
rect 22607 8475 22657 8503
rect 22607 8455 22620 8475
rect 22640 8455 22657 8475
rect 18884 8323 18934 8336
rect 19092 8323 19142 8336
rect 19300 8323 19350 8336
rect 19513 8323 19563 8336
rect 22607 8426 22657 8455
rect 22820 8474 22870 8503
rect 22820 8450 22831 8474
rect 22855 8450 22870 8474
rect 22820 8426 22870 8450
rect 23028 8479 23078 8503
rect 23028 8455 23040 8479
rect 23064 8455 23078 8479
rect 23028 8426 23078 8455
rect 23236 8477 23286 8503
rect 29849 8559 29899 8575
rect 30057 8559 30107 8575
rect 30265 8559 30315 8575
rect 30478 8559 30528 8575
rect 30897 8555 30947 8571
rect 31105 8555 31155 8571
rect 31313 8555 31363 8571
rect 31526 8555 31576 8571
rect 23236 8451 23254 8477
rect 23280 8451 23286 8477
rect 23236 8426 23286 8451
rect 26210 8466 26260 8494
rect 26210 8446 26223 8466
rect 26243 8446 26260 8466
rect 26210 8417 26260 8446
rect 26423 8465 26473 8494
rect 26423 8441 26434 8465
rect 26458 8441 26473 8465
rect 26423 8417 26473 8441
rect 26631 8470 26681 8494
rect 26631 8446 26643 8470
rect 26667 8446 26681 8470
rect 26631 8417 26681 8446
rect 26839 8468 26889 8494
rect 26839 8442 26857 8468
rect 26883 8442 26889 8468
rect 26839 8417 26889 8442
rect 29849 8492 29899 8517
rect 29849 8466 29855 8492
rect 29881 8466 29899 8492
rect 29849 8440 29899 8466
rect 30057 8488 30107 8517
rect 30057 8464 30071 8488
rect 30095 8464 30107 8488
rect 30057 8440 30107 8464
rect 30265 8493 30315 8517
rect 30265 8469 30280 8493
rect 30304 8469 30315 8493
rect 30265 8440 30315 8469
rect 30478 8488 30528 8517
rect 30478 8468 30495 8488
rect 30515 8468 30528 8488
rect 30478 8440 30528 8468
rect 30897 8488 30947 8513
rect 30897 8462 30903 8488
rect 30929 8462 30947 8488
rect 22607 8368 22657 8384
rect 22820 8368 22870 8384
rect 23028 8368 23078 8384
rect 23236 8368 23286 8384
rect 26210 8359 26260 8375
rect 26423 8359 26473 8375
rect 26631 8359 26681 8375
rect 26839 8359 26889 8375
rect 19932 8319 19982 8332
rect 20140 8319 20190 8332
rect 20348 8319 20398 8332
rect 20561 8319 20611 8332
rect 30897 8436 30947 8462
rect 31105 8484 31155 8513
rect 31105 8460 31119 8484
rect 31143 8460 31155 8484
rect 31105 8436 31155 8460
rect 31313 8489 31363 8513
rect 31313 8465 31328 8489
rect 31352 8465 31363 8489
rect 31313 8436 31363 8465
rect 31526 8484 31576 8513
rect 31526 8464 31543 8484
rect 31563 8464 31576 8484
rect 31526 8436 31576 8464
rect 36918 8588 36968 8601
rect 37131 8588 37181 8601
rect 37339 8588 37389 8601
rect 37547 8588 37597 8601
rect 33315 8469 33365 8497
rect 29849 8327 29899 8340
rect 30057 8327 30107 8340
rect 30265 8327 30315 8340
rect 30478 8327 30528 8340
rect 33315 8449 33328 8469
rect 33348 8449 33365 8469
rect 33315 8420 33365 8449
rect 33528 8468 33578 8497
rect 33528 8444 33539 8468
rect 33563 8444 33578 8468
rect 33528 8420 33578 8444
rect 33736 8473 33786 8497
rect 33736 8449 33748 8473
rect 33772 8449 33786 8473
rect 33736 8420 33786 8449
rect 33944 8471 33994 8497
rect 40557 8553 40607 8569
rect 40765 8553 40815 8569
rect 40973 8553 41023 8569
rect 41186 8553 41236 8569
rect 41605 8549 41655 8565
rect 41813 8549 41863 8565
rect 42021 8549 42071 8565
rect 42234 8549 42284 8565
rect 33944 8445 33962 8471
rect 33988 8445 33994 8471
rect 33944 8420 33994 8445
rect 36918 8460 36968 8488
rect 36918 8440 36931 8460
rect 36951 8440 36968 8460
rect 36918 8411 36968 8440
rect 37131 8459 37181 8488
rect 37131 8435 37142 8459
rect 37166 8435 37181 8459
rect 37131 8411 37181 8435
rect 37339 8464 37389 8488
rect 37339 8440 37351 8464
rect 37375 8440 37389 8464
rect 37339 8411 37389 8440
rect 37547 8462 37597 8488
rect 37547 8436 37565 8462
rect 37591 8436 37597 8462
rect 37547 8411 37597 8436
rect 40557 8486 40607 8511
rect 40557 8460 40563 8486
rect 40589 8460 40607 8486
rect 40557 8434 40607 8460
rect 40765 8482 40815 8511
rect 40765 8458 40779 8482
rect 40803 8458 40815 8482
rect 40765 8434 40815 8458
rect 40973 8487 41023 8511
rect 40973 8463 40988 8487
rect 41012 8463 41023 8487
rect 40973 8434 41023 8463
rect 41186 8482 41236 8511
rect 41186 8462 41203 8482
rect 41223 8462 41236 8482
rect 41186 8434 41236 8462
rect 41605 8482 41655 8507
rect 41605 8456 41611 8482
rect 41637 8456 41655 8482
rect 33315 8362 33365 8378
rect 33528 8362 33578 8378
rect 33736 8362 33786 8378
rect 33944 8362 33994 8378
rect 36918 8353 36968 8369
rect 37131 8353 37181 8369
rect 37339 8353 37389 8369
rect 37547 8353 37597 8369
rect 30897 8323 30947 8336
rect 31105 8323 31155 8336
rect 31313 8323 31363 8336
rect 31526 8323 31576 8336
rect 41605 8430 41655 8456
rect 41813 8478 41863 8507
rect 41813 8454 41827 8478
rect 41851 8454 41863 8478
rect 41813 8430 41863 8454
rect 42021 8483 42071 8507
rect 42021 8459 42036 8483
rect 42060 8459 42071 8483
rect 42021 8430 42071 8459
rect 42234 8478 42284 8507
rect 42234 8458 42251 8478
rect 42271 8458 42284 8478
rect 42234 8430 42284 8458
rect 40557 8321 40607 8334
rect 40765 8321 40815 8334
rect 40973 8321 41023 8334
rect 41186 8321 41236 8334
rect 41605 8317 41655 8330
rect 41813 8317 41863 8330
rect 42021 8317 42071 8330
rect 42234 8317 42284 8330
rect 931 7690 981 7703
rect 1144 7690 1194 7703
rect 1352 7690 1402 7703
rect 1560 7690 1610 7703
rect 1979 7686 2029 7699
rect 2192 7686 2242 7699
rect 2400 7686 2450 7699
rect 2608 7686 2658 7699
rect 931 7562 981 7590
rect 931 7542 944 7562
rect 964 7542 981 7562
rect 931 7513 981 7542
rect 1144 7561 1194 7590
rect 1144 7537 1155 7561
rect 1179 7537 1194 7561
rect 1144 7513 1194 7537
rect 1352 7566 1402 7590
rect 1352 7542 1364 7566
rect 1388 7542 1402 7566
rect 1352 7513 1402 7542
rect 1560 7564 1610 7590
rect 11639 7684 11689 7697
rect 11852 7684 11902 7697
rect 12060 7684 12110 7697
rect 12268 7684 12318 7697
rect 5618 7651 5668 7667
rect 5826 7651 5876 7667
rect 6034 7651 6084 7667
rect 6247 7651 6297 7667
rect 9221 7642 9271 7658
rect 9429 7642 9479 7658
rect 9637 7642 9687 7658
rect 9850 7642 9900 7658
rect 1560 7538 1578 7564
rect 1604 7538 1610 7564
rect 1560 7513 1610 7538
rect 1979 7558 2029 7586
rect 1979 7538 1992 7558
rect 2012 7538 2029 7558
rect 1979 7509 2029 7538
rect 2192 7557 2242 7586
rect 2192 7533 2203 7557
rect 2227 7533 2242 7557
rect 2192 7509 2242 7533
rect 2400 7562 2450 7586
rect 2400 7538 2412 7562
rect 2436 7538 2450 7562
rect 2400 7509 2450 7538
rect 2608 7560 2658 7586
rect 2608 7534 2626 7560
rect 2652 7534 2658 7560
rect 2608 7509 2658 7534
rect 5618 7584 5668 7609
rect 5618 7558 5624 7584
rect 5650 7558 5668 7584
rect 5618 7532 5668 7558
rect 5826 7580 5876 7609
rect 5826 7556 5840 7580
rect 5864 7556 5876 7580
rect 5826 7532 5876 7556
rect 6034 7585 6084 7609
rect 6034 7561 6049 7585
rect 6073 7561 6084 7585
rect 6034 7532 6084 7561
rect 6247 7580 6297 7609
rect 6247 7560 6264 7580
rect 6284 7560 6297 7580
rect 6247 7532 6297 7560
rect 9221 7575 9271 7600
rect 9221 7549 9227 7575
rect 9253 7549 9271 7575
rect 931 7455 981 7471
rect 1144 7455 1194 7471
rect 1352 7455 1402 7471
rect 1560 7455 1610 7471
rect 1979 7451 2029 7467
rect 2192 7451 2242 7467
rect 2400 7451 2450 7467
rect 2608 7451 2658 7467
rect 9221 7523 9271 7549
rect 9429 7571 9479 7600
rect 9429 7547 9443 7571
rect 9467 7547 9479 7571
rect 9429 7523 9479 7547
rect 9637 7576 9687 7600
rect 9637 7552 9652 7576
rect 9676 7552 9687 7576
rect 9637 7523 9687 7552
rect 9850 7571 9900 7600
rect 9850 7551 9867 7571
rect 9887 7551 9900 7571
rect 12687 7680 12737 7693
rect 12900 7680 12950 7693
rect 13108 7680 13158 7693
rect 13316 7680 13366 7693
rect 9850 7523 9900 7551
rect 5618 7419 5668 7432
rect 5826 7419 5876 7432
rect 6034 7419 6084 7432
rect 6247 7419 6297 7432
rect 11639 7556 11689 7584
rect 11639 7536 11652 7556
rect 11672 7536 11689 7556
rect 11639 7507 11689 7536
rect 11852 7555 11902 7584
rect 11852 7531 11863 7555
rect 11887 7531 11902 7555
rect 11852 7507 11902 7531
rect 12060 7560 12110 7584
rect 12060 7536 12072 7560
rect 12096 7536 12110 7560
rect 12060 7507 12110 7536
rect 12268 7558 12318 7584
rect 22604 7688 22654 7701
rect 22817 7688 22867 7701
rect 23025 7688 23075 7701
rect 23233 7688 23283 7701
rect 16326 7645 16376 7661
rect 16534 7645 16584 7661
rect 16742 7645 16792 7661
rect 16955 7645 17005 7661
rect 19929 7636 19979 7652
rect 20137 7636 20187 7652
rect 20345 7636 20395 7652
rect 20558 7636 20608 7652
rect 12268 7532 12286 7558
rect 12312 7532 12318 7558
rect 12268 7507 12318 7532
rect 12687 7552 12737 7580
rect 12687 7532 12700 7552
rect 12720 7532 12737 7552
rect 12687 7503 12737 7532
rect 12900 7551 12950 7580
rect 12900 7527 12911 7551
rect 12935 7527 12950 7551
rect 12900 7503 12950 7527
rect 13108 7556 13158 7580
rect 13108 7532 13120 7556
rect 13144 7532 13158 7556
rect 13108 7503 13158 7532
rect 13316 7554 13366 7580
rect 13316 7528 13334 7554
rect 13360 7528 13366 7554
rect 13316 7503 13366 7528
rect 16326 7578 16376 7603
rect 16326 7552 16332 7578
rect 16358 7552 16376 7578
rect 16326 7526 16376 7552
rect 16534 7574 16584 7603
rect 16534 7550 16548 7574
rect 16572 7550 16584 7574
rect 16534 7526 16584 7550
rect 16742 7579 16792 7603
rect 16742 7555 16757 7579
rect 16781 7555 16792 7579
rect 16742 7526 16792 7555
rect 16955 7574 17005 7603
rect 16955 7554 16972 7574
rect 16992 7554 17005 7574
rect 16955 7526 17005 7554
rect 19929 7569 19979 7594
rect 19929 7543 19935 7569
rect 19961 7543 19979 7569
rect 11639 7449 11689 7465
rect 11852 7449 11902 7465
rect 12060 7449 12110 7465
rect 12268 7449 12318 7465
rect 12687 7445 12737 7461
rect 12900 7445 12950 7461
rect 13108 7445 13158 7461
rect 13316 7445 13366 7461
rect 19929 7517 19979 7543
rect 20137 7565 20187 7594
rect 20137 7541 20151 7565
rect 20175 7541 20187 7565
rect 20137 7517 20187 7541
rect 20345 7570 20395 7594
rect 20345 7546 20360 7570
rect 20384 7546 20395 7570
rect 20345 7517 20395 7546
rect 20558 7565 20608 7594
rect 23652 7684 23702 7697
rect 23865 7684 23915 7697
rect 24073 7684 24123 7697
rect 24281 7684 24331 7697
rect 20558 7545 20575 7565
rect 20595 7545 20608 7565
rect 20558 7517 20608 7545
rect 9221 7410 9271 7423
rect 9429 7410 9479 7423
rect 9637 7410 9687 7423
rect 9850 7410 9900 7423
rect 16326 7413 16376 7426
rect 16534 7413 16584 7426
rect 16742 7413 16792 7426
rect 16955 7413 17005 7426
rect 22604 7560 22654 7588
rect 22604 7540 22617 7560
rect 22637 7540 22654 7560
rect 22604 7511 22654 7540
rect 22817 7559 22867 7588
rect 22817 7535 22828 7559
rect 22852 7535 22867 7559
rect 22817 7511 22867 7535
rect 23025 7564 23075 7588
rect 23025 7540 23037 7564
rect 23061 7540 23075 7564
rect 23025 7511 23075 7540
rect 23233 7562 23283 7588
rect 33312 7682 33362 7695
rect 33525 7682 33575 7695
rect 33733 7682 33783 7695
rect 33941 7682 33991 7695
rect 27291 7649 27341 7665
rect 27499 7649 27549 7665
rect 27707 7649 27757 7665
rect 27920 7649 27970 7665
rect 30894 7640 30944 7656
rect 31102 7640 31152 7656
rect 31310 7640 31360 7656
rect 31523 7640 31573 7656
rect 23233 7536 23251 7562
rect 23277 7536 23283 7562
rect 23233 7511 23283 7536
rect 23652 7556 23702 7584
rect 23652 7536 23665 7556
rect 23685 7536 23702 7556
rect 23652 7507 23702 7536
rect 23865 7555 23915 7584
rect 23865 7531 23876 7555
rect 23900 7531 23915 7555
rect 23865 7507 23915 7531
rect 24073 7560 24123 7584
rect 24073 7536 24085 7560
rect 24109 7536 24123 7560
rect 24073 7507 24123 7536
rect 24281 7558 24331 7584
rect 24281 7532 24299 7558
rect 24325 7532 24331 7558
rect 24281 7507 24331 7532
rect 27291 7582 27341 7607
rect 27291 7556 27297 7582
rect 27323 7556 27341 7582
rect 27291 7530 27341 7556
rect 27499 7578 27549 7607
rect 27499 7554 27513 7578
rect 27537 7554 27549 7578
rect 27499 7530 27549 7554
rect 27707 7583 27757 7607
rect 27707 7559 27722 7583
rect 27746 7559 27757 7583
rect 27707 7530 27757 7559
rect 27920 7578 27970 7607
rect 27920 7558 27937 7578
rect 27957 7558 27970 7578
rect 27920 7530 27970 7558
rect 30894 7573 30944 7598
rect 30894 7547 30900 7573
rect 30926 7547 30944 7573
rect 22604 7453 22654 7469
rect 22817 7453 22867 7469
rect 23025 7453 23075 7469
rect 23233 7453 23283 7469
rect 23652 7449 23702 7465
rect 23865 7449 23915 7465
rect 24073 7449 24123 7465
rect 24281 7449 24331 7465
rect 30894 7521 30944 7547
rect 31102 7569 31152 7598
rect 31102 7545 31116 7569
rect 31140 7545 31152 7569
rect 31102 7521 31152 7545
rect 31310 7574 31360 7598
rect 31310 7550 31325 7574
rect 31349 7550 31360 7574
rect 31310 7521 31360 7550
rect 31523 7569 31573 7598
rect 31523 7549 31540 7569
rect 31560 7549 31573 7569
rect 34360 7678 34410 7691
rect 34573 7678 34623 7691
rect 34781 7678 34831 7691
rect 34989 7678 35039 7691
rect 31523 7521 31573 7549
rect 19929 7404 19979 7417
rect 20137 7404 20187 7417
rect 20345 7404 20395 7417
rect 20558 7404 20608 7417
rect 27291 7417 27341 7430
rect 27499 7417 27549 7430
rect 27707 7417 27757 7430
rect 27920 7417 27970 7430
rect 33312 7554 33362 7582
rect 33312 7534 33325 7554
rect 33345 7534 33362 7554
rect 33312 7505 33362 7534
rect 33525 7553 33575 7582
rect 33525 7529 33536 7553
rect 33560 7529 33575 7553
rect 33525 7505 33575 7529
rect 33733 7558 33783 7582
rect 33733 7534 33745 7558
rect 33769 7534 33783 7558
rect 33733 7505 33783 7534
rect 33941 7556 33991 7582
rect 37999 7643 38049 7659
rect 38207 7643 38257 7659
rect 38415 7643 38465 7659
rect 38628 7643 38678 7659
rect 41602 7634 41652 7650
rect 41810 7634 41860 7650
rect 42018 7634 42068 7650
rect 42231 7634 42281 7650
rect 33941 7530 33959 7556
rect 33985 7530 33991 7556
rect 33941 7505 33991 7530
rect 34360 7550 34410 7578
rect 34360 7530 34373 7550
rect 34393 7530 34410 7550
rect 34360 7501 34410 7530
rect 34573 7549 34623 7578
rect 34573 7525 34584 7549
rect 34608 7525 34623 7549
rect 34573 7501 34623 7525
rect 34781 7554 34831 7578
rect 34781 7530 34793 7554
rect 34817 7530 34831 7554
rect 34781 7501 34831 7530
rect 34989 7552 35039 7578
rect 34989 7526 35007 7552
rect 35033 7526 35039 7552
rect 34989 7501 35039 7526
rect 37999 7576 38049 7601
rect 37999 7550 38005 7576
rect 38031 7550 38049 7576
rect 37999 7524 38049 7550
rect 38207 7572 38257 7601
rect 38207 7548 38221 7572
rect 38245 7548 38257 7572
rect 38207 7524 38257 7548
rect 38415 7577 38465 7601
rect 38415 7553 38430 7577
rect 38454 7553 38465 7577
rect 38415 7524 38465 7553
rect 38628 7572 38678 7601
rect 38628 7552 38645 7572
rect 38665 7552 38678 7572
rect 38628 7524 38678 7552
rect 41602 7567 41652 7592
rect 41602 7541 41608 7567
rect 41634 7541 41652 7567
rect 33312 7447 33362 7463
rect 33525 7447 33575 7463
rect 33733 7447 33783 7463
rect 33941 7447 33991 7463
rect 34360 7443 34410 7459
rect 34573 7443 34623 7459
rect 34781 7443 34831 7459
rect 34989 7443 35039 7459
rect 41602 7515 41652 7541
rect 41810 7563 41860 7592
rect 41810 7539 41824 7563
rect 41848 7539 41860 7563
rect 41810 7515 41860 7539
rect 42018 7568 42068 7592
rect 42018 7544 42033 7568
rect 42057 7544 42068 7568
rect 42018 7515 42068 7544
rect 42231 7563 42281 7592
rect 42231 7543 42248 7563
rect 42268 7543 42281 7563
rect 42231 7515 42281 7543
rect 30894 7408 30944 7421
rect 31102 7408 31152 7421
rect 31310 7408 31360 7421
rect 31523 7408 31573 7421
rect 37999 7411 38049 7424
rect 38207 7411 38257 7424
rect 38415 7411 38465 7424
rect 38628 7411 38678 7424
rect 41602 7402 41652 7415
rect 41810 7402 41860 7415
rect 42018 7402 42068 7415
rect 42231 7402 42281 7415
rect 931 7011 981 7024
rect 1144 7011 1194 7024
rect 1352 7011 1402 7024
rect 1560 7011 1610 7024
rect 3426 7006 3476 7019
rect 3639 7006 3689 7019
rect 3847 7006 3897 7019
rect 4055 7006 4105 7019
rect 931 6883 981 6911
rect 931 6863 944 6883
rect 964 6863 981 6883
rect 931 6834 981 6863
rect 1144 6882 1194 6911
rect 1144 6858 1155 6882
rect 1179 6858 1194 6882
rect 1144 6834 1194 6858
rect 1352 6887 1402 6911
rect 1352 6863 1364 6887
rect 1388 6863 1402 6887
rect 1352 6834 1402 6863
rect 1560 6885 1610 6911
rect 11639 7005 11689 7018
rect 11852 7005 11902 7018
rect 12060 7005 12110 7018
rect 12268 7005 12318 7018
rect 8173 6967 8223 6983
rect 8381 6967 8431 6983
rect 8589 6967 8639 6983
rect 8802 6967 8852 6983
rect 9221 6963 9271 6979
rect 9429 6963 9479 6979
rect 9637 6963 9687 6979
rect 9850 6963 9900 6979
rect 1560 6859 1578 6885
rect 1604 6859 1610 6885
rect 1560 6834 1610 6859
rect 3426 6878 3476 6906
rect 3426 6858 3439 6878
rect 3459 6858 3476 6878
rect 3426 6829 3476 6858
rect 3639 6877 3689 6906
rect 3639 6853 3650 6877
rect 3674 6853 3689 6877
rect 3639 6829 3689 6853
rect 3847 6882 3897 6906
rect 3847 6858 3859 6882
rect 3883 6858 3897 6882
rect 3847 6829 3897 6858
rect 4055 6880 4105 6906
rect 4055 6854 4073 6880
rect 4099 6854 4105 6880
rect 4055 6829 4105 6854
rect 8173 6900 8223 6925
rect 8173 6874 8179 6900
rect 8205 6874 8223 6900
rect 8173 6848 8223 6874
rect 8381 6896 8431 6925
rect 8381 6872 8395 6896
rect 8419 6872 8431 6896
rect 8381 6848 8431 6872
rect 8589 6901 8639 6925
rect 8589 6877 8604 6901
rect 8628 6877 8639 6901
rect 8589 6848 8639 6877
rect 8802 6896 8852 6925
rect 8802 6876 8819 6896
rect 8839 6876 8852 6896
rect 8802 6848 8852 6876
rect 9221 6896 9271 6921
rect 9221 6870 9227 6896
rect 9253 6870 9271 6896
rect 931 6776 981 6792
rect 1144 6776 1194 6792
rect 1352 6776 1402 6792
rect 1560 6776 1610 6792
rect 3426 6771 3476 6787
rect 3639 6771 3689 6787
rect 3847 6771 3897 6787
rect 4055 6771 4105 6787
rect 9221 6844 9271 6870
rect 9429 6892 9479 6921
rect 9429 6868 9443 6892
rect 9467 6868 9479 6892
rect 9429 6844 9479 6868
rect 9637 6897 9687 6921
rect 9637 6873 9652 6897
rect 9676 6873 9687 6897
rect 9637 6844 9687 6873
rect 9850 6892 9900 6921
rect 9850 6872 9867 6892
rect 9887 6872 9900 6892
rect 9850 6844 9900 6872
rect 14134 7000 14184 7013
rect 14347 7000 14397 7013
rect 14555 7000 14605 7013
rect 14763 7000 14813 7013
rect 11639 6877 11689 6905
rect 8173 6735 8223 6748
rect 8381 6735 8431 6748
rect 8589 6735 8639 6748
rect 8802 6735 8852 6748
rect 11639 6857 11652 6877
rect 11672 6857 11689 6877
rect 11639 6828 11689 6857
rect 11852 6876 11902 6905
rect 11852 6852 11863 6876
rect 11887 6852 11902 6876
rect 11852 6828 11902 6852
rect 12060 6881 12110 6905
rect 12060 6857 12072 6881
rect 12096 6857 12110 6881
rect 12060 6828 12110 6857
rect 12268 6879 12318 6905
rect 22604 7009 22654 7022
rect 22817 7009 22867 7022
rect 23025 7009 23075 7022
rect 23233 7009 23283 7022
rect 18881 6961 18931 6977
rect 19089 6961 19139 6977
rect 19297 6961 19347 6977
rect 19510 6961 19560 6977
rect 19929 6957 19979 6973
rect 20137 6957 20187 6973
rect 20345 6957 20395 6973
rect 20558 6957 20608 6973
rect 12268 6853 12286 6879
rect 12312 6853 12318 6879
rect 12268 6828 12318 6853
rect 14134 6872 14184 6900
rect 14134 6852 14147 6872
rect 14167 6852 14184 6872
rect 14134 6823 14184 6852
rect 14347 6871 14397 6900
rect 14347 6847 14358 6871
rect 14382 6847 14397 6871
rect 14347 6823 14397 6847
rect 14555 6876 14605 6900
rect 14555 6852 14567 6876
rect 14591 6852 14605 6876
rect 14555 6823 14605 6852
rect 14763 6874 14813 6900
rect 14763 6848 14781 6874
rect 14807 6848 14813 6874
rect 14763 6823 14813 6848
rect 18881 6894 18931 6919
rect 18881 6868 18887 6894
rect 18913 6868 18931 6894
rect 18881 6842 18931 6868
rect 19089 6890 19139 6919
rect 19089 6866 19103 6890
rect 19127 6866 19139 6890
rect 19089 6842 19139 6866
rect 19297 6895 19347 6919
rect 19297 6871 19312 6895
rect 19336 6871 19347 6895
rect 19297 6842 19347 6871
rect 19510 6890 19560 6919
rect 19510 6870 19527 6890
rect 19547 6870 19560 6890
rect 19510 6842 19560 6870
rect 19929 6890 19979 6915
rect 19929 6864 19935 6890
rect 19961 6864 19979 6890
rect 11639 6770 11689 6786
rect 11852 6770 11902 6786
rect 12060 6770 12110 6786
rect 12268 6770 12318 6786
rect 14134 6765 14184 6781
rect 14347 6765 14397 6781
rect 14555 6765 14605 6781
rect 14763 6765 14813 6781
rect 9221 6731 9271 6744
rect 9429 6731 9479 6744
rect 9637 6731 9687 6744
rect 9850 6731 9900 6744
rect 19929 6838 19979 6864
rect 20137 6886 20187 6915
rect 20137 6862 20151 6886
rect 20175 6862 20187 6886
rect 20137 6838 20187 6862
rect 20345 6891 20395 6915
rect 20345 6867 20360 6891
rect 20384 6867 20395 6891
rect 20345 6838 20395 6867
rect 20558 6886 20608 6915
rect 20558 6866 20575 6886
rect 20595 6866 20608 6886
rect 20558 6838 20608 6866
rect 25099 7004 25149 7017
rect 25312 7004 25362 7017
rect 25520 7004 25570 7017
rect 25728 7004 25778 7017
rect 22604 6881 22654 6909
rect 22604 6861 22617 6881
rect 22637 6861 22654 6881
rect 18881 6729 18931 6742
rect 19089 6729 19139 6742
rect 19297 6729 19347 6742
rect 19510 6729 19560 6742
rect 22604 6832 22654 6861
rect 22817 6880 22867 6909
rect 22817 6856 22828 6880
rect 22852 6856 22867 6880
rect 22817 6832 22867 6856
rect 23025 6885 23075 6909
rect 23025 6861 23037 6885
rect 23061 6861 23075 6885
rect 23025 6832 23075 6861
rect 23233 6883 23283 6909
rect 33312 7003 33362 7016
rect 33525 7003 33575 7016
rect 33733 7003 33783 7016
rect 33941 7003 33991 7016
rect 29846 6965 29896 6981
rect 30054 6965 30104 6981
rect 30262 6965 30312 6981
rect 30475 6965 30525 6981
rect 30894 6961 30944 6977
rect 31102 6961 31152 6977
rect 31310 6961 31360 6977
rect 31523 6961 31573 6977
rect 23233 6857 23251 6883
rect 23277 6857 23283 6883
rect 23233 6832 23283 6857
rect 25099 6876 25149 6904
rect 25099 6856 25112 6876
rect 25132 6856 25149 6876
rect 25099 6827 25149 6856
rect 25312 6875 25362 6904
rect 25312 6851 25323 6875
rect 25347 6851 25362 6875
rect 25312 6827 25362 6851
rect 25520 6880 25570 6904
rect 25520 6856 25532 6880
rect 25556 6856 25570 6880
rect 25520 6827 25570 6856
rect 25728 6878 25778 6904
rect 25728 6852 25746 6878
rect 25772 6852 25778 6878
rect 25728 6827 25778 6852
rect 29846 6898 29896 6923
rect 29846 6872 29852 6898
rect 29878 6872 29896 6898
rect 29846 6846 29896 6872
rect 30054 6894 30104 6923
rect 30054 6870 30068 6894
rect 30092 6870 30104 6894
rect 30054 6846 30104 6870
rect 30262 6899 30312 6923
rect 30262 6875 30277 6899
rect 30301 6875 30312 6899
rect 30262 6846 30312 6875
rect 30475 6894 30525 6923
rect 30475 6874 30492 6894
rect 30512 6874 30525 6894
rect 30475 6846 30525 6874
rect 30894 6894 30944 6919
rect 30894 6868 30900 6894
rect 30926 6868 30944 6894
rect 22604 6774 22654 6790
rect 22817 6774 22867 6790
rect 23025 6774 23075 6790
rect 23233 6774 23283 6790
rect 25099 6769 25149 6785
rect 25312 6769 25362 6785
rect 25520 6769 25570 6785
rect 25728 6769 25778 6785
rect 19929 6725 19979 6738
rect 20137 6725 20187 6738
rect 20345 6725 20395 6738
rect 20558 6725 20608 6738
rect 30894 6842 30944 6868
rect 31102 6890 31152 6919
rect 31102 6866 31116 6890
rect 31140 6866 31152 6890
rect 31102 6842 31152 6866
rect 31310 6895 31360 6919
rect 31310 6871 31325 6895
rect 31349 6871 31360 6895
rect 31310 6842 31360 6871
rect 31523 6890 31573 6919
rect 31523 6870 31540 6890
rect 31560 6870 31573 6890
rect 31523 6842 31573 6870
rect 35807 6998 35857 7011
rect 36020 6998 36070 7011
rect 36228 6998 36278 7011
rect 36436 6998 36486 7011
rect 33312 6875 33362 6903
rect 29846 6733 29896 6746
rect 30054 6733 30104 6746
rect 30262 6733 30312 6746
rect 30475 6733 30525 6746
rect 33312 6855 33325 6875
rect 33345 6855 33362 6875
rect 33312 6826 33362 6855
rect 33525 6874 33575 6903
rect 33525 6850 33536 6874
rect 33560 6850 33575 6874
rect 33525 6826 33575 6850
rect 33733 6879 33783 6903
rect 33733 6855 33745 6879
rect 33769 6855 33783 6879
rect 33733 6826 33783 6855
rect 33941 6877 33991 6903
rect 40554 6959 40604 6975
rect 40762 6959 40812 6975
rect 40970 6959 41020 6975
rect 41183 6959 41233 6975
rect 41602 6955 41652 6971
rect 41810 6955 41860 6971
rect 42018 6955 42068 6971
rect 42231 6955 42281 6971
rect 33941 6851 33959 6877
rect 33985 6851 33991 6877
rect 33941 6826 33991 6851
rect 35807 6870 35857 6898
rect 35807 6850 35820 6870
rect 35840 6850 35857 6870
rect 35807 6821 35857 6850
rect 36020 6869 36070 6898
rect 36020 6845 36031 6869
rect 36055 6845 36070 6869
rect 36020 6821 36070 6845
rect 36228 6874 36278 6898
rect 36228 6850 36240 6874
rect 36264 6850 36278 6874
rect 36228 6821 36278 6850
rect 36436 6872 36486 6898
rect 36436 6846 36454 6872
rect 36480 6846 36486 6872
rect 36436 6821 36486 6846
rect 40554 6892 40604 6917
rect 40554 6866 40560 6892
rect 40586 6866 40604 6892
rect 40554 6840 40604 6866
rect 40762 6888 40812 6917
rect 40762 6864 40776 6888
rect 40800 6864 40812 6888
rect 40762 6840 40812 6864
rect 40970 6893 41020 6917
rect 40970 6869 40985 6893
rect 41009 6869 41020 6893
rect 40970 6840 41020 6869
rect 41183 6888 41233 6917
rect 41183 6868 41200 6888
rect 41220 6868 41233 6888
rect 41183 6840 41233 6868
rect 41602 6888 41652 6913
rect 41602 6862 41608 6888
rect 41634 6862 41652 6888
rect 33312 6768 33362 6784
rect 33525 6768 33575 6784
rect 33733 6768 33783 6784
rect 33941 6768 33991 6784
rect 35807 6763 35857 6779
rect 36020 6763 36070 6779
rect 36228 6763 36278 6779
rect 36436 6763 36486 6779
rect 30894 6729 30944 6742
rect 31102 6729 31152 6742
rect 31310 6729 31360 6742
rect 31523 6729 31573 6742
rect 41602 6836 41652 6862
rect 41810 6884 41860 6913
rect 41810 6860 41824 6884
rect 41848 6860 41860 6884
rect 41810 6836 41860 6860
rect 42018 6889 42068 6913
rect 42018 6865 42033 6889
rect 42057 6865 42068 6889
rect 42018 6836 42068 6865
rect 42231 6884 42281 6913
rect 42231 6864 42248 6884
rect 42268 6864 42281 6884
rect 42231 6836 42281 6864
rect 40554 6727 40604 6740
rect 40762 6727 40812 6740
rect 40970 6727 41020 6740
rect 41183 6727 41233 6740
rect 41602 6723 41652 6736
rect 41810 6723 41860 6736
rect 42018 6723 42068 6736
rect 42231 6723 42281 6736
rect 931 6243 981 6256
rect 1144 6243 1194 6256
rect 1352 6243 1402 6256
rect 1560 6243 1610 6256
rect 1979 6239 2029 6252
rect 2192 6239 2242 6252
rect 2400 6239 2450 6252
rect 2608 6239 2658 6252
rect 931 6115 981 6143
rect 931 6095 944 6115
rect 964 6095 981 6115
rect 931 6066 981 6095
rect 1144 6114 1194 6143
rect 1144 6090 1155 6114
rect 1179 6090 1194 6114
rect 1144 6066 1194 6090
rect 1352 6119 1402 6143
rect 1352 6095 1364 6119
rect 1388 6095 1402 6119
rect 1352 6066 1402 6095
rect 1560 6117 1610 6143
rect 11639 6237 11689 6250
rect 11852 6237 11902 6250
rect 12060 6237 12110 6250
rect 12268 6237 12318 6250
rect 6726 6200 6776 6216
rect 6934 6200 6984 6216
rect 7142 6200 7192 6216
rect 7355 6200 7405 6216
rect 9221 6195 9271 6211
rect 9429 6195 9479 6211
rect 9637 6195 9687 6211
rect 9850 6195 9900 6211
rect 1560 6091 1578 6117
rect 1604 6091 1610 6117
rect 1560 6066 1610 6091
rect 1979 6111 2029 6139
rect 1979 6091 1992 6111
rect 2012 6091 2029 6111
rect 1979 6062 2029 6091
rect 2192 6110 2242 6139
rect 2192 6086 2203 6110
rect 2227 6086 2242 6110
rect 2192 6062 2242 6086
rect 2400 6115 2450 6139
rect 2400 6091 2412 6115
rect 2436 6091 2450 6115
rect 2400 6062 2450 6091
rect 2608 6113 2658 6139
rect 2608 6087 2626 6113
rect 2652 6087 2658 6113
rect 2608 6062 2658 6087
rect 6726 6133 6776 6158
rect 6726 6107 6732 6133
rect 6758 6107 6776 6133
rect 6726 6081 6776 6107
rect 6934 6129 6984 6158
rect 6934 6105 6948 6129
rect 6972 6105 6984 6129
rect 6934 6081 6984 6105
rect 7142 6134 7192 6158
rect 7142 6110 7157 6134
rect 7181 6110 7192 6134
rect 7142 6081 7192 6110
rect 7355 6129 7405 6158
rect 7355 6109 7372 6129
rect 7392 6109 7405 6129
rect 7355 6081 7405 6109
rect 9221 6128 9271 6153
rect 9221 6102 9227 6128
rect 9253 6102 9271 6128
rect 931 6008 981 6024
rect 1144 6008 1194 6024
rect 1352 6008 1402 6024
rect 1560 6008 1610 6024
rect 1979 6004 2029 6020
rect 2192 6004 2242 6020
rect 2400 6004 2450 6020
rect 2608 6004 2658 6020
rect 9221 6076 9271 6102
rect 9429 6124 9479 6153
rect 9429 6100 9443 6124
rect 9467 6100 9479 6124
rect 9429 6076 9479 6100
rect 9637 6129 9687 6153
rect 9637 6105 9652 6129
rect 9676 6105 9687 6129
rect 9637 6076 9687 6105
rect 9850 6124 9900 6153
rect 9850 6104 9867 6124
rect 9887 6104 9900 6124
rect 12687 6233 12737 6246
rect 12900 6233 12950 6246
rect 13108 6233 13158 6246
rect 13316 6233 13366 6246
rect 9850 6076 9900 6104
rect 6726 5968 6776 5981
rect 6934 5968 6984 5981
rect 7142 5968 7192 5981
rect 7355 5968 7405 5981
rect 11639 6109 11689 6137
rect 11639 6089 11652 6109
rect 11672 6089 11689 6109
rect 11639 6060 11689 6089
rect 11852 6108 11902 6137
rect 11852 6084 11863 6108
rect 11887 6084 11902 6108
rect 11852 6060 11902 6084
rect 12060 6113 12110 6137
rect 12060 6089 12072 6113
rect 12096 6089 12110 6113
rect 12060 6060 12110 6089
rect 12268 6111 12318 6137
rect 22604 6241 22654 6254
rect 22817 6241 22867 6254
rect 23025 6241 23075 6254
rect 23233 6241 23283 6254
rect 17434 6194 17484 6210
rect 17642 6194 17692 6210
rect 17850 6194 17900 6210
rect 18063 6194 18113 6210
rect 19929 6189 19979 6205
rect 20137 6189 20187 6205
rect 20345 6189 20395 6205
rect 20558 6189 20608 6205
rect 12268 6085 12286 6111
rect 12312 6085 12318 6111
rect 12268 6060 12318 6085
rect 12687 6105 12737 6133
rect 12687 6085 12700 6105
rect 12720 6085 12737 6105
rect 12687 6056 12737 6085
rect 12900 6104 12950 6133
rect 12900 6080 12911 6104
rect 12935 6080 12950 6104
rect 12900 6056 12950 6080
rect 13108 6109 13158 6133
rect 13108 6085 13120 6109
rect 13144 6085 13158 6109
rect 13108 6056 13158 6085
rect 13316 6107 13366 6133
rect 13316 6081 13334 6107
rect 13360 6081 13366 6107
rect 13316 6056 13366 6081
rect 17434 6127 17484 6152
rect 17434 6101 17440 6127
rect 17466 6101 17484 6127
rect 17434 6075 17484 6101
rect 17642 6123 17692 6152
rect 17642 6099 17656 6123
rect 17680 6099 17692 6123
rect 17642 6075 17692 6099
rect 17850 6128 17900 6152
rect 17850 6104 17865 6128
rect 17889 6104 17900 6128
rect 17850 6075 17900 6104
rect 18063 6123 18113 6152
rect 18063 6103 18080 6123
rect 18100 6103 18113 6123
rect 18063 6075 18113 6103
rect 19929 6122 19979 6147
rect 19929 6096 19935 6122
rect 19961 6096 19979 6122
rect 11639 6002 11689 6018
rect 11852 6002 11902 6018
rect 12060 6002 12110 6018
rect 12268 6002 12318 6018
rect 12687 5998 12737 6014
rect 12900 5998 12950 6014
rect 13108 5998 13158 6014
rect 13316 5998 13366 6014
rect 9221 5963 9271 5976
rect 9429 5963 9479 5976
rect 9637 5963 9687 5976
rect 9850 5963 9900 5976
rect 19929 6070 19979 6096
rect 20137 6118 20187 6147
rect 20137 6094 20151 6118
rect 20175 6094 20187 6118
rect 20137 6070 20187 6094
rect 20345 6123 20395 6147
rect 20345 6099 20360 6123
rect 20384 6099 20395 6123
rect 20345 6070 20395 6099
rect 20558 6118 20608 6147
rect 23652 6237 23702 6250
rect 23865 6237 23915 6250
rect 24073 6237 24123 6250
rect 24281 6237 24331 6250
rect 20558 6098 20575 6118
rect 20595 6098 20608 6118
rect 20558 6070 20608 6098
rect 17434 5962 17484 5975
rect 17642 5962 17692 5975
rect 17850 5962 17900 5975
rect 18063 5962 18113 5975
rect 22604 6113 22654 6141
rect 22604 6093 22617 6113
rect 22637 6093 22654 6113
rect 22604 6064 22654 6093
rect 22817 6112 22867 6141
rect 22817 6088 22828 6112
rect 22852 6088 22867 6112
rect 22817 6064 22867 6088
rect 23025 6117 23075 6141
rect 23025 6093 23037 6117
rect 23061 6093 23075 6117
rect 23025 6064 23075 6093
rect 23233 6115 23283 6141
rect 33312 6235 33362 6248
rect 33525 6235 33575 6248
rect 33733 6235 33783 6248
rect 33941 6235 33991 6248
rect 28399 6198 28449 6214
rect 28607 6198 28657 6214
rect 28815 6198 28865 6214
rect 29028 6198 29078 6214
rect 30894 6193 30944 6209
rect 31102 6193 31152 6209
rect 31310 6193 31360 6209
rect 31523 6193 31573 6209
rect 23233 6089 23251 6115
rect 23277 6089 23283 6115
rect 23233 6064 23283 6089
rect 23652 6109 23702 6137
rect 23652 6089 23665 6109
rect 23685 6089 23702 6109
rect 23652 6060 23702 6089
rect 23865 6108 23915 6137
rect 23865 6084 23876 6108
rect 23900 6084 23915 6108
rect 23865 6060 23915 6084
rect 24073 6113 24123 6137
rect 24073 6089 24085 6113
rect 24109 6089 24123 6113
rect 24073 6060 24123 6089
rect 24281 6111 24331 6137
rect 24281 6085 24299 6111
rect 24325 6085 24331 6111
rect 24281 6060 24331 6085
rect 28399 6131 28449 6156
rect 28399 6105 28405 6131
rect 28431 6105 28449 6131
rect 28399 6079 28449 6105
rect 28607 6127 28657 6156
rect 28607 6103 28621 6127
rect 28645 6103 28657 6127
rect 28607 6079 28657 6103
rect 28815 6132 28865 6156
rect 28815 6108 28830 6132
rect 28854 6108 28865 6132
rect 28815 6079 28865 6108
rect 29028 6127 29078 6156
rect 29028 6107 29045 6127
rect 29065 6107 29078 6127
rect 29028 6079 29078 6107
rect 30894 6126 30944 6151
rect 30894 6100 30900 6126
rect 30926 6100 30944 6126
rect 22604 6006 22654 6022
rect 22817 6006 22867 6022
rect 23025 6006 23075 6022
rect 23233 6006 23283 6022
rect 23652 6002 23702 6018
rect 23865 6002 23915 6018
rect 24073 6002 24123 6018
rect 24281 6002 24331 6018
rect 19929 5957 19979 5970
rect 20137 5957 20187 5970
rect 20345 5957 20395 5970
rect 20558 5957 20608 5970
rect 30894 6074 30944 6100
rect 31102 6122 31152 6151
rect 31102 6098 31116 6122
rect 31140 6098 31152 6122
rect 31102 6074 31152 6098
rect 31310 6127 31360 6151
rect 31310 6103 31325 6127
rect 31349 6103 31360 6127
rect 31310 6074 31360 6103
rect 31523 6122 31573 6151
rect 31523 6102 31540 6122
rect 31560 6102 31573 6122
rect 34360 6231 34410 6244
rect 34573 6231 34623 6244
rect 34781 6231 34831 6244
rect 34989 6231 35039 6244
rect 31523 6074 31573 6102
rect 28399 5966 28449 5979
rect 28607 5966 28657 5979
rect 28815 5966 28865 5979
rect 29028 5966 29078 5979
rect 33312 6107 33362 6135
rect 33312 6087 33325 6107
rect 33345 6087 33362 6107
rect 33312 6058 33362 6087
rect 33525 6106 33575 6135
rect 33525 6082 33536 6106
rect 33560 6082 33575 6106
rect 33525 6058 33575 6082
rect 33733 6111 33783 6135
rect 33733 6087 33745 6111
rect 33769 6087 33783 6111
rect 33733 6058 33783 6087
rect 33941 6109 33991 6135
rect 39107 6192 39157 6208
rect 39315 6192 39365 6208
rect 39523 6192 39573 6208
rect 39736 6192 39786 6208
rect 41602 6187 41652 6203
rect 41810 6187 41860 6203
rect 42018 6187 42068 6203
rect 42231 6187 42281 6203
rect 33941 6083 33959 6109
rect 33985 6083 33991 6109
rect 33941 6058 33991 6083
rect 34360 6103 34410 6131
rect 34360 6083 34373 6103
rect 34393 6083 34410 6103
rect 34360 6054 34410 6083
rect 34573 6102 34623 6131
rect 34573 6078 34584 6102
rect 34608 6078 34623 6102
rect 34573 6054 34623 6078
rect 34781 6107 34831 6131
rect 34781 6083 34793 6107
rect 34817 6083 34831 6107
rect 34781 6054 34831 6083
rect 34989 6105 35039 6131
rect 34989 6079 35007 6105
rect 35033 6079 35039 6105
rect 34989 6054 35039 6079
rect 39107 6125 39157 6150
rect 39107 6099 39113 6125
rect 39139 6099 39157 6125
rect 39107 6073 39157 6099
rect 39315 6121 39365 6150
rect 39315 6097 39329 6121
rect 39353 6097 39365 6121
rect 39315 6073 39365 6097
rect 39523 6126 39573 6150
rect 39523 6102 39538 6126
rect 39562 6102 39573 6126
rect 39523 6073 39573 6102
rect 39736 6121 39786 6150
rect 39736 6101 39753 6121
rect 39773 6101 39786 6121
rect 39736 6073 39786 6101
rect 41602 6120 41652 6145
rect 41602 6094 41608 6120
rect 41634 6094 41652 6120
rect 33312 6000 33362 6016
rect 33525 6000 33575 6016
rect 33733 6000 33783 6016
rect 33941 6000 33991 6016
rect 34360 5996 34410 6012
rect 34573 5996 34623 6012
rect 34781 5996 34831 6012
rect 34989 5996 35039 6012
rect 30894 5961 30944 5974
rect 31102 5961 31152 5974
rect 31310 5961 31360 5974
rect 31523 5961 31573 5974
rect 41602 6068 41652 6094
rect 41810 6116 41860 6145
rect 41810 6092 41824 6116
rect 41848 6092 41860 6116
rect 41810 6068 41860 6092
rect 42018 6121 42068 6145
rect 42018 6097 42033 6121
rect 42057 6097 42068 6121
rect 42018 6068 42068 6097
rect 42231 6116 42281 6145
rect 42231 6096 42248 6116
rect 42268 6096 42281 6116
rect 42231 6068 42281 6096
rect 39107 5960 39157 5973
rect 39315 5960 39365 5973
rect 39523 5960 39573 5973
rect 39736 5960 39786 5973
rect 41602 5955 41652 5968
rect 41810 5955 41860 5968
rect 42018 5955 42068 5968
rect 42231 5955 42281 5968
rect 931 5564 981 5577
rect 1144 5564 1194 5577
rect 1352 5564 1402 5577
rect 1560 5564 1610 5577
rect 3469 5561 3519 5574
rect 3682 5561 3732 5574
rect 3890 5561 3940 5574
rect 4098 5561 4148 5574
rect 931 5436 981 5464
rect 931 5416 944 5436
rect 964 5416 981 5436
rect 931 5387 981 5416
rect 1144 5435 1194 5464
rect 1144 5411 1155 5435
rect 1179 5411 1194 5435
rect 1144 5387 1194 5411
rect 1352 5440 1402 5464
rect 1352 5416 1364 5440
rect 1388 5416 1402 5440
rect 1352 5387 1402 5416
rect 1560 5438 1610 5464
rect 11639 5558 11689 5571
rect 11852 5558 11902 5571
rect 12060 5558 12110 5571
rect 12268 5558 12318 5571
rect 8173 5520 8223 5536
rect 8381 5520 8431 5536
rect 8589 5520 8639 5536
rect 8802 5520 8852 5536
rect 9221 5516 9271 5532
rect 9429 5516 9479 5532
rect 9637 5516 9687 5532
rect 9850 5516 9900 5532
rect 1560 5412 1578 5438
rect 1604 5412 1610 5438
rect 1560 5387 1610 5412
rect 3469 5433 3519 5461
rect 3469 5413 3482 5433
rect 3502 5413 3519 5433
rect 3469 5384 3519 5413
rect 3682 5432 3732 5461
rect 3682 5408 3693 5432
rect 3717 5408 3732 5432
rect 3682 5384 3732 5408
rect 3890 5437 3940 5461
rect 3890 5413 3902 5437
rect 3926 5413 3940 5437
rect 3890 5384 3940 5413
rect 4098 5435 4148 5461
rect 4098 5409 4116 5435
rect 4142 5409 4148 5435
rect 4098 5384 4148 5409
rect 8173 5453 8223 5478
rect 8173 5427 8179 5453
rect 8205 5427 8223 5453
rect 8173 5401 8223 5427
rect 8381 5449 8431 5478
rect 8381 5425 8395 5449
rect 8419 5425 8431 5449
rect 8381 5401 8431 5425
rect 8589 5454 8639 5478
rect 8589 5430 8604 5454
rect 8628 5430 8639 5454
rect 8589 5401 8639 5430
rect 8802 5449 8852 5478
rect 8802 5429 8819 5449
rect 8839 5429 8852 5449
rect 8802 5401 8852 5429
rect 9221 5449 9271 5474
rect 9221 5423 9227 5449
rect 9253 5423 9271 5449
rect 931 5329 981 5345
rect 1144 5329 1194 5345
rect 1352 5329 1402 5345
rect 1560 5329 1610 5345
rect 3469 5326 3519 5342
rect 3682 5326 3732 5342
rect 3890 5326 3940 5342
rect 4098 5326 4148 5342
rect 9221 5397 9271 5423
rect 9429 5445 9479 5474
rect 9429 5421 9443 5445
rect 9467 5421 9479 5445
rect 9429 5397 9479 5421
rect 9637 5450 9687 5474
rect 9637 5426 9652 5450
rect 9676 5426 9687 5450
rect 9637 5397 9687 5426
rect 9850 5445 9900 5474
rect 9850 5425 9867 5445
rect 9887 5425 9900 5445
rect 9850 5397 9900 5425
rect 14177 5555 14227 5568
rect 14390 5555 14440 5568
rect 14598 5555 14648 5568
rect 14806 5555 14856 5568
rect 11639 5430 11689 5458
rect 8173 5288 8223 5301
rect 8381 5288 8431 5301
rect 8589 5288 8639 5301
rect 8802 5288 8852 5301
rect 11639 5410 11652 5430
rect 11672 5410 11689 5430
rect 11639 5381 11689 5410
rect 11852 5429 11902 5458
rect 11852 5405 11863 5429
rect 11887 5405 11902 5429
rect 11852 5381 11902 5405
rect 12060 5434 12110 5458
rect 12060 5410 12072 5434
rect 12096 5410 12110 5434
rect 12060 5381 12110 5410
rect 12268 5432 12318 5458
rect 22604 5562 22654 5575
rect 22817 5562 22867 5575
rect 23025 5562 23075 5575
rect 23233 5562 23283 5575
rect 18881 5514 18931 5530
rect 19089 5514 19139 5530
rect 19297 5514 19347 5530
rect 19510 5514 19560 5530
rect 19929 5510 19979 5526
rect 20137 5510 20187 5526
rect 20345 5510 20395 5526
rect 20558 5510 20608 5526
rect 12268 5406 12286 5432
rect 12312 5406 12318 5432
rect 12268 5381 12318 5406
rect 14177 5427 14227 5455
rect 14177 5407 14190 5427
rect 14210 5407 14227 5427
rect 14177 5378 14227 5407
rect 14390 5426 14440 5455
rect 14390 5402 14401 5426
rect 14425 5402 14440 5426
rect 14390 5378 14440 5402
rect 14598 5431 14648 5455
rect 14598 5407 14610 5431
rect 14634 5407 14648 5431
rect 14598 5378 14648 5407
rect 14806 5429 14856 5455
rect 14806 5403 14824 5429
rect 14850 5403 14856 5429
rect 14806 5378 14856 5403
rect 18881 5447 18931 5472
rect 18881 5421 18887 5447
rect 18913 5421 18931 5447
rect 18881 5395 18931 5421
rect 19089 5443 19139 5472
rect 19089 5419 19103 5443
rect 19127 5419 19139 5443
rect 19089 5395 19139 5419
rect 19297 5448 19347 5472
rect 19297 5424 19312 5448
rect 19336 5424 19347 5448
rect 19297 5395 19347 5424
rect 19510 5443 19560 5472
rect 19510 5423 19527 5443
rect 19547 5423 19560 5443
rect 19510 5395 19560 5423
rect 19929 5443 19979 5468
rect 19929 5417 19935 5443
rect 19961 5417 19979 5443
rect 11639 5323 11689 5339
rect 11852 5323 11902 5339
rect 12060 5323 12110 5339
rect 12268 5323 12318 5339
rect 14177 5320 14227 5336
rect 14390 5320 14440 5336
rect 14598 5320 14648 5336
rect 14806 5320 14856 5336
rect 9221 5284 9271 5297
rect 9429 5284 9479 5297
rect 9637 5284 9687 5297
rect 9850 5284 9900 5297
rect 19929 5391 19979 5417
rect 20137 5439 20187 5468
rect 20137 5415 20151 5439
rect 20175 5415 20187 5439
rect 20137 5391 20187 5415
rect 20345 5444 20395 5468
rect 20345 5420 20360 5444
rect 20384 5420 20395 5444
rect 20345 5391 20395 5420
rect 20558 5439 20608 5468
rect 20558 5419 20575 5439
rect 20595 5419 20608 5439
rect 20558 5391 20608 5419
rect 25142 5559 25192 5572
rect 25355 5559 25405 5572
rect 25563 5559 25613 5572
rect 25771 5559 25821 5572
rect 22604 5434 22654 5462
rect 22604 5414 22617 5434
rect 22637 5414 22654 5434
rect 18881 5282 18931 5295
rect 19089 5282 19139 5295
rect 19297 5282 19347 5295
rect 19510 5282 19560 5295
rect 22604 5385 22654 5414
rect 22817 5433 22867 5462
rect 22817 5409 22828 5433
rect 22852 5409 22867 5433
rect 22817 5385 22867 5409
rect 23025 5438 23075 5462
rect 23025 5414 23037 5438
rect 23061 5414 23075 5438
rect 23025 5385 23075 5414
rect 23233 5436 23283 5462
rect 33312 5556 33362 5569
rect 33525 5556 33575 5569
rect 33733 5556 33783 5569
rect 33941 5556 33991 5569
rect 29846 5518 29896 5534
rect 30054 5518 30104 5534
rect 30262 5518 30312 5534
rect 30475 5518 30525 5534
rect 30894 5514 30944 5530
rect 31102 5514 31152 5530
rect 31310 5514 31360 5530
rect 31523 5514 31573 5530
rect 23233 5410 23251 5436
rect 23277 5410 23283 5436
rect 23233 5385 23283 5410
rect 25142 5431 25192 5459
rect 25142 5411 25155 5431
rect 25175 5411 25192 5431
rect 25142 5382 25192 5411
rect 25355 5430 25405 5459
rect 25355 5406 25366 5430
rect 25390 5406 25405 5430
rect 25355 5382 25405 5406
rect 25563 5435 25613 5459
rect 25563 5411 25575 5435
rect 25599 5411 25613 5435
rect 25563 5382 25613 5411
rect 25771 5433 25821 5459
rect 25771 5407 25789 5433
rect 25815 5407 25821 5433
rect 25771 5382 25821 5407
rect 29846 5451 29896 5476
rect 29846 5425 29852 5451
rect 29878 5425 29896 5451
rect 29846 5399 29896 5425
rect 30054 5447 30104 5476
rect 30054 5423 30068 5447
rect 30092 5423 30104 5447
rect 30054 5399 30104 5423
rect 30262 5452 30312 5476
rect 30262 5428 30277 5452
rect 30301 5428 30312 5452
rect 30262 5399 30312 5428
rect 30475 5447 30525 5476
rect 30475 5427 30492 5447
rect 30512 5427 30525 5447
rect 30475 5399 30525 5427
rect 30894 5447 30944 5472
rect 30894 5421 30900 5447
rect 30926 5421 30944 5447
rect 22604 5327 22654 5343
rect 22817 5327 22867 5343
rect 23025 5327 23075 5343
rect 23233 5327 23283 5343
rect 25142 5324 25192 5340
rect 25355 5324 25405 5340
rect 25563 5324 25613 5340
rect 25771 5324 25821 5340
rect 19929 5278 19979 5291
rect 20137 5278 20187 5291
rect 20345 5278 20395 5291
rect 20558 5278 20608 5291
rect 30894 5395 30944 5421
rect 31102 5443 31152 5472
rect 31102 5419 31116 5443
rect 31140 5419 31152 5443
rect 31102 5395 31152 5419
rect 31310 5448 31360 5472
rect 31310 5424 31325 5448
rect 31349 5424 31360 5448
rect 31310 5395 31360 5424
rect 31523 5443 31573 5472
rect 31523 5423 31540 5443
rect 31560 5423 31573 5443
rect 31523 5395 31573 5423
rect 35850 5553 35900 5566
rect 36063 5553 36113 5566
rect 36271 5553 36321 5566
rect 36479 5553 36529 5566
rect 33312 5428 33362 5456
rect 29846 5286 29896 5299
rect 30054 5286 30104 5299
rect 30262 5286 30312 5299
rect 30475 5286 30525 5299
rect 33312 5408 33325 5428
rect 33345 5408 33362 5428
rect 33312 5379 33362 5408
rect 33525 5427 33575 5456
rect 33525 5403 33536 5427
rect 33560 5403 33575 5427
rect 33525 5379 33575 5403
rect 33733 5432 33783 5456
rect 33733 5408 33745 5432
rect 33769 5408 33783 5432
rect 33733 5379 33783 5408
rect 33941 5430 33991 5456
rect 40554 5512 40604 5528
rect 40762 5512 40812 5528
rect 40970 5512 41020 5528
rect 41183 5512 41233 5528
rect 41602 5508 41652 5524
rect 41810 5508 41860 5524
rect 42018 5508 42068 5524
rect 42231 5508 42281 5524
rect 33941 5404 33959 5430
rect 33985 5404 33991 5430
rect 33941 5379 33991 5404
rect 35850 5425 35900 5453
rect 35850 5405 35863 5425
rect 35883 5405 35900 5425
rect 35850 5376 35900 5405
rect 36063 5424 36113 5453
rect 36063 5400 36074 5424
rect 36098 5400 36113 5424
rect 36063 5376 36113 5400
rect 36271 5429 36321 5453
rect 36271 5405 36283 5429
rect 36307 5405 36321 5429
rect 36271 5376 36321 5405
rect 36479 5427 36529 5453
rect 36479 5401 36497 5427
rect 36523 5401 36529 5427
rect 36479 5376 36529 5401
rect 40554 5445 40604 5470
rect 40554 5419 40560 5445
rect 40586 5419 40604 5445
rect 40554 5393 40604 5419
rect 40762 5441 40812 5470
rect 40762 5417 40776 5441
rect 40800 5417 40812 5441
rect 40762 5393 40812 5417
rect 40970 5446 41020 5470
rect 40970 5422 40985 5446
rect 41009 5422 41020 5446
rect 40970 5393 41020 5422
rect 41183 5441 41233 5470
rect 41183 5421 41200 5441
rect 41220 5421 41233 5441
rect 41183 5393 41233 5421
rect 41602 5441 41652 5466
rect 41602 5415 41608 5441
rect 41634 5415 41652 5441
rect 33312 5321 33362 5337
rect 33525 5321 33575 5337
rect 33733 5321 33783 5337
rect 33941 5321 33991 5337
rect 35850 5318 35900 5334
rect 36063 5318 36113 5334
rect 36271 5318 36321 5334
rect 36479 5318 36529 5334
rect 30894 5282 30944 5295
rect 31102 5282 31152 5295
rect 31310 5282 31360 5295
rect 31523 5282 31573 5295
rect 41602 5389 41652 5415
rect 41810 5437 41860 5466
rect 41810 5413 41824 5437
rect 41848 5413 41860 5437
rect 41810 5389 41860 5413
rect 42018 5442 42068 5466
rect 42018 5418 42033 5442
rect 42057 5418 42068 5442
rect 42018 5389 42068 5418
rect 42231 5437 42281 5466
rect 42231 5417 42248 5437
rect 42268 5417 42281 5437
rect 42231 5389 42281 5417
rect 40554 5280 40604 5293
rect 40762 5280 40812 5293
rect 40970 5280 41020 5293
rect 41183 5280 41233 5293
rect 41602 5276 41652 5289
rect 41810 5276 41860 5289
rect 42018 5276 42068 5289
rect 42231 5276 42281 5289
rect 932 4723 982 4736
rect 1145 4723 1195 4736
rect 1353 4723 1403 4736
rect 1561 4723 1611 4736
rect 1980 4719 2030 4732
rect 2193 4719 2243 4732
rect 2401 4719 2451 4732
rect 2609 4719 2659 4732
rect 4882 4725 4932 4738
rect 5095 4725 5145 4738
rect 5303 4725 5353 4738
rect 5511 4725 5561 4738
rect 932 4595 982 4623
rect 932 4575 945 4595
rect 965 4575 982 4595
rect 932 4546 982 4575
rect 1145 4594 1195 4623
rect 1145 4570 1156 4594
rect 1180 4570 1195 4594
rect 1145 4546 1195 4570
rect 1353 4599 1403 4623
rect 1353 4575 1365 4599
rect 1389 4575 1403 4599
rect 1353 4546 1403 4575
rect 1561 4597 1611 4623
rect 11640 4717 11690 4730
rect 11853 4717 11903 4730
rect 12061 4717 12111 4730
rect 12269 4717 12319 4730
rect 6684 4678 6734 4694
rect 6892 4678 6942 4694
rect 7100 4678 7150 4694
rect 7313 4678 7363 4694
rect 9222 4675 9272 4691
rect 9430 4675 9480 4691
rect 9638 4675 9688 4691
rect 9851 4675 9901 4691
rect 1561 4571 1579 4597
rect 1605 4571 1611 4597
rect 1561 4546 1611 4571
rect 1980 4591 2030 4619
rect 1980 4571 1993 4591
rect 2013 4571 2030 4591
rect 1980 4542 2030 4571
rect 2193 4590 2243 4619
rect 2193 4566 2204 4590
rect 2228 4566 2243 4590
rect 2193 4542 2243 4566
rect 2401 4595 2451 4619
rect 2401 4571 2413 4595
rect 2437 4571 2451 4595
rect 2401 4542 2451 4571
rect 2609 4593 2659 4619
rect 2609 4567 2627 4593
rect 2653 4567 2659 4593
rect 2609 4542 2659 4567
rect 4882 4597 4932 4625
rect 4882 4577 4895 4597
rect 4915 4577 4932 4597
rect 4882 4548 4932 4577
rect 5095 4596 5145 4625
rect 5095 4572 5106 4596
rect 5130 4572 5145 4596
rect 5095 4548 5145 4572
rect 5303 4601 5353 4625
rect 5303 4577 5315 4601
rect 5339 4577 5353 4601
rect 5303 4548 5353 4577
rect 5511 4599 5561 4625
rect 5511 4573 5529 4599
rect 5555 4573 5561 4599
rect 5511 4548 5561 4573
rect 6684 4611 6734 4636
rect 6684 4585 6690 4611
rect 6716 4585 6734 4611
rect 6684 4559 6734 4585
rect 6892 4607 6942 4636
rect 6892 4583 6906 4607
rect 6930 4583 6942 4607
rect 6892 4559 6942 4583
rect 7100 4612 7150 4636
rect 7100 4588 7115 4612
rect 7139 4588 7150 4612
rect 7100 4559 7150 4588
rect 7313 4607 7363 4636
rect 7313 4587 7330 4607
rect 7350 4587 7363 4607
rect 7313 4559 7363 4587
rect 9222 4608 9272 4633
rect 9222 4582 9228 4608
rect 9254 4582 9272 4608
rect 932 4488 982 4504
rect 1145 4488 1195 4504
rect 1353 4488 1403 4504
rect 1561 4488 1611 4504
rect 1980 4484 2030 4500
rect 2193 4484 2243 4500
rect 2401 4484 2451 4500
rect 2609 4484 2659 4500
rect 4882 4490 4932 4506
rect 5095 4490 5145 4506
rect 5303 4490 5353 4506
rect 5511 4490 5561 4506
rect 9222 4556 9272 4582
rect 9430 4604 9480 4633
rect 9430 4580 9444 4604
rect 9468 4580 9480 4604
rect 9430 4556 9480 4580
rect 9638 4609 9688 4633
rect 9638 4585 9653 4609
rect 9677 4585 9688 4609
rect 9638 4556 9688 4585
rect 9851 4604 9901 4633
rect 9851 4584 9868 4604
rect 9888 4584 9901 4604
rect 12688 4713 12738 4726
rect 12901 4713 12951 4726
rect 13109 4713 13159 4726
rect 13317 4713 13367 4726
rect 15590 4719 15640 4732
rect 15803 4719 15853 4732
rect 16011 4719 16061 4732
rect 16219 4719 16269 4732
rect 9851 4556 9901 4584
rect 6684 4446 6734 4459
rect 6892 4446 6942 4459
rect 7100 4446 7150 4459
rect 7313 4446 7363 4459
rect 11640 4589 11690 4617
rect 11640 4569 11653 4589
rect 11673 4569 11690 4589
rect 11640 4540 11690 4569
rect 11853 4588 11903 4617
rect 11853 4564 11864 4588
rect 11888 4564 11903 4588
rect 11853 4540 11903 4564
rect 12061 4593 12111 4617
rect 12061 4569 12073 4593
rect 12097 4569 12111 4593
rect 12061 4540 12111 4569
rect 12269 4591 12319 4617
rect 22605 4721 22655 4734
rect 22818 4721 22868 4734
rect 23026 4721 23076 4734
rect 23234 4721 23284 4734
rect 17392 4672 17442 4688
rect 17600 4672 17650 4688
rect 17808 4672 17858 4688
rect 18021 4672 18071 4688
rect 19930 4669 19980 4685
rect 20138 4669 20188 4685
rect 20346 4669 20396 4685
rect 20559 4669 20609 4685
rect 12269 4565 12287 4591
rect 12313 4565 12319 4591
rect 12269 4540 12319 4565
rect 12688 4585 12738 4613
rect 12688 4565 12701 4585
rect 12721 4565 12738 4585
rect 12688 4536 12738 4565
rect 12901 4584 12951 4613
rect 12901 4560 12912 4584
rect 12936 4560 12951 4584
rect 12901 4536 12951 4560
rect 13109 4589 13159 4613
rect 13109 4565 13121 4589
rect 13145 4565 13159 4589
rect 13109 4536 13159 4565
rect 13317 4587 13367 4613
rect 13317 4561 13335 4587
rect 13361 4561 13367 4587
rect 13317 4536 13367 4561
rect 15590 4591 15640 4619
rect 15590 4571 15603 4591
rect 15623 4571 15640 4591
rect 15590 4542 15640 4571
rect 15803 4590 15853 4619
rect 15803 4566 15814 4590
rect 15838 4566 15853 4590
rect 15803 4542 15853 4566
rect 16011 4595 16061 4619
rect 16011 4571 16023 4595
rect 16047 4571 16061 4595
rect 16011 4542 16061 4571
rect 16219 4593 16269 4619
rect 16219 4567 16237 4593
rect 16263 4567 16269 4593
rect 16219 4542 16269 4567
rect 17392 4605 17442 4630
rect 17392 4579 17398 4605
rect 17424 4579 17442 4605
rect 17392 4553 17442 4579
rect 17600 4601 17650 4630
rect 17600 4577 17614 4601
rect 17638 4577 17650 4601
rect 17600 4553 17650 4577
rect 17808 4606 17858 4630
rect 17808 4582 17823 4606
rect 17847 4582 17858 4606
rect 17808 4553 17858 4582
rect 18021 4601 18071 4630
rect 18021 4581 18038 4601
rect 18058 4581 18071 4601
rect 18021 4553 18071 4581
rect 19930 4602 19980 4627
rect 19930 4576 19936 4602
rect 19962 4576 19980 4602
rect 11640 4482 11690 4498
rect 11853 4482 11903 4498
rect 12061 4482 12111 4498
rect 12269 4482 12319 4498
rect 12688 4478 12738 4494
rect 12901 4478 12951 4494
rect 13109 4478 13159 4494
rect 13317 4478 13367 4494
rect 15590 4484 15640 4500
rect 15803 4484 15853 4500
rect 16011 4484 16061 4500
rect 16219 4484 16269 4500
rect 9222 4443 9272 4456
rect 9430 4443 9480 4456
rect 9638 4443 9688 4456
rect 9851 4443 9901 4456
rect 19930 4550 19980 4576
rect 20138 4598 20188 4627
rect 20138 4574 20152 4598
rect 20176 4574 20188 4598
rect 20138 4550 20188 4574
rect 20346 4603 20396 4627
rect 20346 4579 20361 4603
rect 20385 4579 20396 4603
rect 20346 4550 20396 4579
rect 20559 4598 20609 4627
rect 23653 4717 23703 4730
rect 23866 4717 23916 4730
rect 24074 4717 24124 4730
rect 24282 4717 24332 4730
rect 26555 4723 26605 4736
rect 26768 4723 26818 4736
rect 26976 4723 27026 4736
rect 27184 4723 27234 4736
rect 20559 4578 20576 4598
rect 20596 4578 20609 4598
rect 20559 4550 20609 4578
rect 17392 4440 17442 4453
rect 17600 4440 17650 4453
rect 17808 4440 17858 4453
rect 18021 4440 18071 4453
rect 22605 4593 22655 4621
rect 22605 4573 22618 4593
rect 22638 4573 22655 4593
rect 22605 4544 22655 4573
rect 22818 4592 22868 4621
rect 22818 4568 22829 4592
rect 22853 4568 22868 4592
rect 22818 4544 22868 4568
rect 23026 4597 23076 4621
rect 23026 4573 23038 4597
rect 23062 4573 23076 4597
rect 23026 4544 23076 4573
rect 23234 4595 23284 4621
rect 33313 4715 33363 4728
rect 33526 4715 33576 4728
rect 33734 4715 33784 4728
rect 33942 4715 33992 4728
rect 28357 4676 28407 4692
rect 28565 4676 28615 4692
rect 28773 4676 28823 4692
rect 28986 4676 29036 4692
rect 30895 4673 30945 4689
rect 31103 4673 31153 4689
rect 31311 4673 31361 4689
rect 31524 4673 31574 4689
rect 23234 4569 23252 4595
rect 23278 4569 23284 4595
rect 23234 4544 23284 4569
rect 23653 4589 23703 4617
rect 23653 4569 23666 4589
rect 23686 4569 23703 4589
rect 23653 4540 23703 4569
rect 23866 4588 23916 4617
rect 23866 4564 23877 4588
rect 23901 4564 23916 4588
rect 23866 4540 23916 4564
rect 24074 4593 24124 4617
rect 24074 4569 24086 4593
rect 24110 4569 24124 4593
rect 24074 4540 24124 4569
rect 24282 4591 24332 4617
rect 24282 4565 24300 4591
rect 24326 4565 24332 4591
rect 24282 4540 24332 4565
rect 26555 4595 26605 4623
rect 26555 4575 26568 4595
rect 26588 4575 26605 4595
rect 26555 4546 26605 4575
rect 26768 4594 26818 4623
rect 26768 4570 26779 4594
rect 26803 4570 26818 4594
rect 26768 4546 26818 4570
rect 26976 4599 27026 4623
rect 26976 4575 26988 4599
rect 27012 4575 27026 4599
rect 26976 4546 27026 4575
rect 27184 4597 27234 4623
rect 27184 4571 27202 4597
rect 27228 4571 27234 4597
rect 27184 4546 27234 4571
rect 28357 4609 28407 4634
rect 28357 4583 28363 4609
rect 28389 4583 28407 4609
rect 28357 4557 28407 4583
rect 28565 4605 28615 4634
rect 28565 4581 28579 4605
rect 28603 4581 28615 4605
rect 28565 4557 28615 4581
rect 28773 4610 28823 4634
rect 28773 4586 28788 4610
rect 28812 4586 28823 4610
rect 28773 4557 28823 4586
rect 28986 4605 29036 4634
rect 28986 4585 29003 4605
rect 29023 4585 29036 4605
rect 28986 4557 29036 4585
rect 30895 4606 30945 4631
rect 30895 4580 30901 4606
rect 30927 4580 30945 4606
rect 22605 4486 22655 4502
rect 22818 4486 22868 4502
rect 23026 4486 23076 4502
rect 23234 4486 23284 4502
rect 23653 4482 23703 4498
rect 23866 4482 23916 4498
rect 24074 4482 24124 4498
rect 24282 4482 24332 4498
rect 26555 4488 26605 4504
rect 26768 4488 26818 4504
rect 26976 4488 27026 4504
rect 27184 4488 27234 4504
rect 19930 4437 19980 4450
rect 20138 4437 20188 4450
rect 20346 4437 20396 4450
rect 20559 4437 20609 4450
rect 30895 4554 30945 4580
rect 31103 4602 31153 4631
rect 31103 4578 31117 4602
rect 31141 4578 31153 4602
rect 31103 4554 31153 4578
rect 31311 4607 31361 4631
rect 31311 4583 31326 4607
rect 31350 4583 31361 4607
rect 31311 4554 31361 4583
rect 31524 4602 31574 4631
rect 31524 4582 31541 4602
rect 31561 4582 31574 4602
rect 34361 4711 34411 4724
rect 34574 4711 34624 4724
rect 34782 4711 34832 4724
rect 34990 4711 35040 4724
rect 37263 4717 37313 4730
rect 37476 4717 37526 4730
rect 37684 4717 37734 4730
rect 37892 4717 37942 4730
rect 31524 4554 31574 4582
rect 28357 4444 28407 4457
rect 28565 4444 28615 4457
rect 28773 4444 28823 4457
rect 28986 4444 29036 4457
rect 33313 4587 33363 4615
rect 33313 4567 33326 4587
rect 33346 4567 33363 4587
rect 33313 4538 33363 4567
rect 33526 4586 33576 4615
rect 33526 4562 33537 4586
rect 33561 4562 33576 4586
rect 33526 4538 33576 4562
rect 33734 4591 33784 4615
rect 33734 4567 33746 4591
rect 33770 4567 33784 4591
rect 33734 4538 33784 4567
rect 33942 4589 33992 4615
rect 39065 4670 39115 4686
rect 39273 4670 39323 4686
rect 39481 4670 39531 4686
rect 39694 4670 39744 4686
rect 41603 4667 41653 4683
rect 41811 4667 41861 4683
rect 42019 4667 42069 4683
rect 42232 4667 42282 4683
rect 33942 4563 33960 4589
rect 33986 4563 33992 4589
rect 33942 4538 33992 4563
rect 34361 4583 34411 4611
rect 34361 4563 34374 4583
rect 34394 4563 34411 4583
rect 34361 4534 34411 4563
rect 34574 4582 34624 4611
rect 34574 4558 34585 4582
rect 34609 4558 34624 4582
rect 34574 4534 34624 4558
rect 34782 4587 34832 4611
rect 34782 4563 34794 4587
rect 34818 4563 34832 4587
rect 34782 4534 34832 4563
rect 34990 4585 35040 4611
rect 34990 4559 35008 4585
rect 35034 4559 35040 4585
rect 34990 4534 35040 4559
rect 37263 4589 37313 4617
rect 37263 4569 37276 4589
rect 37296 4569 37313 4589
rect 37263 4540 37313 4569
rect 37476 4588 37526 4617
rect 37476 4564 37487 4588
rect 37511 4564 37526 4588
rect 37476 4540 37526 4564
rect 37684 4593 37734 4617
rect 37684 4569 37696 4593
rect 37720 4569 37734 4593
rect 37684 4540 37734 4569
rect 37892 4591 37942 4617
rect 37892 4565 37910 4591
rect 37936 4565 37942 4591
rect 37892 4540 37942 4565
rect 39065 4603 39115 4628
rect 39065 4577 39071 4603
rect 39097 4577 39115 4603
rect 39065 4551 39115 4577
rect 39273 4599 39323 4628
rect 39273 4575 39287 4599
rect 39311 4575 39323 4599
rect 39273 4551 39323 4575
rect 39481 4604 39531 4628
rect 39481 4580 39496 4604
rect 39520 4580 39531 4604
rect 39481 4551 39531 4580
rect 39694 4599 39744 4628
rect 39694 4579 39711 4599
rect 39731 4579 39744 4599
rect 39694 4551 39744 4579
rect 41603 4600 41653 4625
rect 41603 4574 41609 4600
rect 41635 4574 41653 4600
rect 33313 4480 33363 4496
rect 33526 4480 33576 4496
rect 33734 4480 33784 4496
rect 33942 4480 33992 4496
rect 34361 4476 34411 4492
rect 34574 4476 34624 4492
rect 34782 4476 34832 4492
rect 34990 4476 35040 4492
rect 37263 4482 37313 4498
rect 37476 4482 37526 4498
rect 37684 4482 37734 4498
rect 37892 4482 37942 4498
rect 30895 4441 30945 4454
rect 31103 4441 31153 4454
rect 31311 4441 31361 4454
rect 31524 4441 31574 4454
rect 41603 4548 41653 4574
rect 41811 4596 41861 4625
rect 41811 4572 41825 4596
rect 41849 4572 41861 4596
rect 41811 4548 41861 4572
rect 42019 4601 42069 4625
rect 42019 4577 42034 4601
rect 42058 4577 42069 4601
rect 42019 4548 42069 4577
rect 42232 4596 42282 4625
rect 42232 4576 42249 4596
rect 42269 4576 42282 4596
rect 42232 4548 42282 4576
rect 39065 4438 39115 4451
rect 39273 4438 39323 4451
rect 39481 4438 39531 4451
rect 39694 4438 39744 4451
rect 41603 4435 41653 4448
rect 41811 4435 41861 4448
rect 42019 4435 42069 4448
rect 42232 4435 42282 4448
rect 932 4044 982 4057
rect 1145 4044 1195 4057
rect 1353 4044 1403 4057
rect 1561 4044 1611 4057
rect 3427 4039 3477 4052
rect 3640 4039 3690 4052
rect 3848 4039 3898 4052
rect 4056 4039 4106 4052
rect 932 3916 982 3944
rect 932 3896 945 3916
rect 965 3896 982 3916
rect 932 3867 982 3896
rect 1145 3915 1195 3944
rect 1145 3891 1156 3915
rect 1180 3891 1195 3915
rect 1145 3867 1195 3891
rect 1353 3920 1403 3944
rect 1353 3896 1365 3920
rect 1389 3896 1403 3920
rect 1353 3867 1403 3896
rect 1561 3918 1611 3944
rect 11640 4038 11690 4051
rect 11853 4038 11903 4051
rect 12061 4038 12111 4051
rect 12269 4038 12319 4051
rect 8174 4000 8224 4016
rect 8382 4000 8432 4016
rect 8590 4000 8640 4016
rect 8803 4000 8853 4016
rect 9222 3996 9272 4012
rect 9430 3996 9480 4012
rect 9638 3996 9688 4012
rect 9851 3996 9901 4012
rect 1561 3892 1579 3918
rect 1605 3892 1611 3918
rect 1561 3867 1611 3892
rect 3427 3911 3477 3939
rect 3427 3891 3440 3911
rect 3460 3891 3477 3911
rect 3427 3862 3477 3891
rect 3640 3910 3690 3939
rect 3640 3886 3651 3910
rect 3675 3886 3690 3910
rect 3640 3862 3690 3886
rect 3848 3915 3898 3939
rect 3848 3891 3860 3915
rect 3884 3891 3898 3915
rect 3848 3862 3898 3891
rect 4056 3913 4106 3939
rect 4056 3887 4074 3913
rect 4100 3887 4106 3913
rect 4056 3862 4106 3887
rect 8174 3933 8224 3958
rect 8174 3907 8180 3933
rect 8206 3907 8224 3933
rect 8174 3881 8224 3907
rect 8382 3929 8432 3958
rect 8382 3905 8396 3929
rect 8420 3905 8432 3929
rect 8382 3881 8432 3905
rect 8590 3934 8640 3958
rect 8590 3910 8605 3934
rect 8629 3910 8640 3934
rect 8590 3881 8640 3910
rect 8803 3929 8853 3958
rect 8803 3909 8820 3929
rect 8840 3909 8853 3929
rect 8803 3881 8853 3909
rect 9222 3929 9272 3954
rect 9222 3903 9228 3929
rect 9254 3903 9272 3929
rect 932 3809 982 3825
rect 1145 3809 1195 3825
rect 1353 3809 1403 3825
rect 1561 3809 1611 3825
rect 3427 3804 3477 3820
rect 3640 3804 3690 3820
rect 3848 3804 3898 3820
rect 4056 3804 4106 3820
rect 9222 3877 9272 3903
rect 9430 3925 9480 3954
rect 9430 3901 9444 3925
rect 9468 3901 9480 3925
rect 9430 3877 9480 3901
rect 9638 3930 9688 3954
rect 9638 3906 9653 3930
rect 9677 3906 9688 3930
rect 9638 3877 9688 3906
rect 9851 3925 9901 3954
rect 9851 3905 9868 3925
rect 9888 3905 9901 3925
rect 9851 3877 9901 3905
rect 14135 4033 14185 4046
rect 14348 4033 14398 4046
rect 14556 4033 14606 4046
rect 14764 4033 14814 4046
rect 11640 3910 11690 3938
rect 8174 3768 8224 3781
rect 8382 3768 8432 3781
rect 8590 3768 8640 3781
rect 8803 3768 8853 3781
rect 11640 3890 11653 3910
rect 11673 3890 11690 3910
rect 11640 3861 11690 3890
rect 11853 3909 11903 3938
rect 11853 3885 11864 3909
rect 11888 3885 11903 3909
rect 11853 3861 11903 3885
rect 12061 3914 12111 3938
rect 12061 3890 12073 3914
rect 12097 3890 12111 3914
rect 12061 3861 12111 3890
rect 12269 3912 12319 3938
rect 22605 4042 22655 4055
rect 22818 4042 22868 4055
rect 23026 4042 23076 4055
rect 23234 4042 23284 4055
rect 18882 3994 18932 4010
rect 19090 3994 19140 4010
rect 19298 3994 19348 4010
rect 19511 3994 19561 4010
rect 19930 3990 19980 4006
rect 20138 3990 20188 4006
rect 20346 3990 20396 4006
rect 20559 3990 20609 4006
rect 12269 3886 12287 3912
rect 12313 3886 12319 3912
rect 12269 3861 12319 3886
rect 14135 3905 14185 3933
rect 14135 3885 14148 3905
rect 14168 3885 14185 3905
rect 14135 3856 14185 3885
rect 14348 3904 14398 3933
rect 14348 3880 14359 3904
rect 14383 3880 14398 3904
rect 14348 3856 14398 3880
rect 14556 3909 14606 3933
rect 14556 3885 14568 3909
rect 14592 3885 14606 3909
rect 14556 3856 14606 3885
rect 14764 3907 14814 3933
rect 14764 3881 14782 3907
rect 14808 3881 14814 3907
rect 14764 3856 14814 3881
rect 18882 3927 18932 3952
rect 18882 3901 18888 3927
rect 18914 3901 18932 3927
rect 18882 3875 18932 3901
rect 19090 3923 19140 3952
rect 19090 3899 19104 3923
rect 19128 3899 19140 3923
rect 19090 3875 19140 3899
rect 19298 3928 19348 3952
rect 19298 3904 19313 3928
rect 19337 3904 19348 3928
rect 19298 3875 19348 3904
rect 19511 3923 19561 3952
rect 19511 3903 19528 3923
rect 19548 3903 19561 3923
rect 19511 3875 19561 3903
rect 19930 3923 19980 3948
rect 19930 3897 19936 3923
rect 19962 3897 19980 3923
rect 11640 3803 11690 3819
rect 11853 3803 11903 3819
rect 12061 3803 12111 3819
rect 12269 3803 12319 3819
rect 14135 3798 14185 3814
rect 14348 3798 14398 3814
rect 14556 3798 14606 3814
rect 14764 3798 14814 3814
rect 9222 3764 9272 3777
rect 9430 3764 9480 3777
rect 9638 3764 9688 3777
rect 9851 3764 9901 3777
rect 19930 3871 19980 3897
rect 20138 3919 20188 3948
rect 20138 3895 20152 3919
rect 20176 3895 20188 3919
rect 20138 3871 20188 3895
rect 20346 3924 20396 3948
rect 20346 3900 20361 3924
rect 20385 3900 20396 3924
rect 20346 3871 20396 3900
rect 20559 3919 20609 3948
rect 20559 3899 20576 3919
rect 20596 3899 20609 3919
rect 20559 3871 20609 3899
rect 25100 4037 25150 4050
rect 25313 4037 25363 4050
rect 25521 4037 25571 4050
rect 25729 4037 25779 4050
rect 22605 3914 22655 3942
rect 22605 3894 22618 3914
rect 22638 3894 22655 3914
rect 18882 3762 18932 3775
rect 19090 3762 19140 3775
rect 19298 3762 19348 3775
rect 19511 3762 19561 3775
rect 22605 3865 22655 3894
rect 22818 3913 22868 3942
rect 22818 3889 22829 3913
rect 22853 3889 22868 3913
rect 22818 3865 22868 3889
rect 23026 3918 23076 3942
rect 23026 3894 23038 3918
rect 23062 3894 23076 3918
rect 23026 3865 23076 3894
rect 23234 3916 23284 3942
rect 33313 4036 33363 4049
rect 33526 4036 33576 4049
rect 33734 4036 33784 4049
rect 33942 4036 33992 4049
rect 29847 3998 29897 4014
rect 30055 3998 30105 4014
rect 30263 3998 30313 4014
rect 30476 3998 30526 4014
rect 30895 3994 30945 4010
rect 31103 3994 31153 4010
rect 31311 3994 31361 4010
rect 31524 3994 31574 4010
rect 23234 3890 23252 3916
rect 23278 3890 23284 3916
rect 23234 3865 23284 3890
rect 25100 3909 25150 3937
rect 25100 3889 25113 3909
rect 25133 3889 25150 3909
rect 25100 3860 25150 3889
rect 25313 3908 25363 3937
rect 25313 3884 25324 3908
rect 25348 3884 25363 3908
rect 25313 3860 25363 3884
rect 25521 3913 25571 3937
rect 25521 3889 25533 3913
rect 25557 3889 25571 3913
rect 25521 3860 25571 3889
rect 25729 3911 25779 3937
rect 25729 3885 25747 3911
rect 25773 3885 25779 3911
rect 25729 3860 25779 3885
rect 29847 3931 29897 3956
rect 29847 3905 29853 3931
rect 29879 3905 29897 3931
rect 29847 3879 29897 3905
rect 30055 3927 30105 3956
rect 30055 3903 30069 3927
rect 30093 3903 30105 3927
rect 30055 3879 30105 3903
rect 30263 3932 30313 3956
rect 30263 3908 30278 3932
rect 30302 3908 30313 3932
rect 30263 3879 30313 3908
rect 30476 3927 30526 3956
rect 30476 3907 30493 3927
rect 30513 3907 30526 3927
rect 30476 3879 30526 3907
rect 30895 3927 30945 3952
rect 30895 3901 30901 3927
rect 30927 3901 30945 3927
rect 22605 3807 22655 3823
rect 22818 3807 22868 3823
rect 23026 3807 23076 3823
rect 23234 3807 23284 3823
rect 25100 3802 25150 3818
rect 25313 3802 25363 3818
rect 25521 3802 25571 3818
rect 25729 3802 25779 3818
rect 19930 3758 19980 3771
rect 20138 3758 20188 3771
rect 20346 3758 20396 3771
rect 20559 3758 20609 3771
rect 30895 3875 30945 3901
rect 31103 3923 31153 3952
rect 31103 3899 31117 3923
rect 31141 3899 31153 3923
rect 31103 3875 31153 3899
rect 31311 3928 31361 3952
rect 31311 3904 31326 3928
rect 31350 3904 31361 3928
rect 31311 3875 31361 3904
rect 31524 3923 31574 3952
rect 31524 3903 31541 3923
rect 31561 3903 31574 3923
rect 31524 3875 31574 3903
rect 35808 4031 35858 4044
rect 36021 4031 36071 4044
rect 36229 4031 36279 4044
rect 36437 4031 36487 4044
rect 33313 3908 33363 3936
rect 29847 3766 29897 3779
rect 30055 3766 30105 3779
rect 30263 3766 30313 3779
rect 30476 3766 30526 3779
rect 33313 3888 33326 3908
rect 33346 3888 33363 3908
rect 33313 3859 33363 3888
rect 33526 3907 33576 3936
rect 33526 3883 33537 3907
rect 33561 3883 33576 3907
rect 33526 3859 33576 3883
rect 33734 3912 33784 3936
rect 33734 3888 33746 3912
rect 33770 3888 33784 3912
rect 33734 3859 33784 3888
rect 33942 3910 33992 3936
rect 40555 3992 40605 4008
rect 40763 3992 40813 4008
rect 40971 3992 41021 4008
rect 41184 3992 41234 4008
rect 41603 3988 41653 4004
rect 41811 3988 41861 4004
rect 42019 3988 42069 4004
rect 42232 3988 42282 4004
rect 33942 3884 33960 3910
rect 33986 3884 33992 3910
rect 33942 3859 33992 3884
rect 35808 3903 35858 3931
rect 35808 3883 35821 3903
rect 35841 3883 35858 3903
rect 35808 3854 35858 3883
rect 36021 3902 36071 3931
rect 36021 3878 36032 3902
rect 36056 3878 36071 3902
rect 36021 3854 36071 3878
rect 36229 3907 36279 3931
rect 36229 3883 36241 3907
rect 36265 3883 36279 3907
rect 36229 3854 36279 3883
rect 36437 3905 36487 3931
rect 36437 3879 36455 3905
rect 36481 3879 36487 3905
rect 36437 3854 36487 3879
rect 40555 3925 40605 3950
rect 40555 3899 40561 3925
rect 40587 3899 40605 3925
rect 40555 3873 40605 3899
rect 40763 3921 40813 3950
rect 40763 3897 40777 3921
rect 40801 3897 40813 3921
rect 40763 3873 40813 3897
rect 40971 3926 41021 3950
rect 40971 3902 40986 3926
rect 41010 3902 41021 3926
rect 40971 3873 41021 3902
rect 41184 3921 41234 3950
rect 41184 3901 41201 3921
rect 41221 3901 41234 3921
rect 41184 3873 41234 3901
rect 41603 3921 41653 3946
rect 41603 3895 41609 3921
rect 41635 3895 41653 3921
rect 33313 3801 33363 3817
rect 33526 3801 33576 3817
rect 33734 3801 33784 3817
rect 33942 3801 33992 3817
rect 35808 3796 35858 3812
rect 36021 3796 36071 3812
rect 36229 3796 36279 3812
rect 36437 3796 36487 3812
rect 30895 3762 30945 3775
rect 31103 3762 31153 3775
rect 31311 3762 31361 3775
rect 31524 3762 31574 3775
rect 41603 3869 41653 3895
rect 41811 3917 41861 3946
rect 41811 3893 41825 3917
rect 41849 3893 41861 3917
rect 41811 3869 41861 3893
rect 42019 3922 42069 3946
rect 42019 3898 42034 3922
rect 42058 3898 42069 3922
rect 42019 3869 42069 3898
rect 42232 3917 42282 3946
rect 42232 3897 42249 3917
rect 42269 3897 42282 3917
rect 42232 3869 42282 3897
rect 40555 3760 40605 3773
rect 40763 3760 40813 3773
rect 40971 3760 41021 3773
rect 41184 3760 41234 3773
rect 41603 3756 41653 3769
rect 41811 3756 41861 3769
rect 42019 3756 42069 3769
rect 42232 3756 42282 3769
rect 932 3276 982 3289
rect 1145 3276 1195 3289
rect 1353 3276 1403 3289
rect 1561 3276 1611 3289
rect 1980 3272 2030 3285
rect 2193 3272 2243 3285
rect 2401 3272 2451 3285
rect 2609 3272 2659 3285
rect 932 3148 982 3176
rect 932 3128 945 3148
rect 965 3128 982 3148
rect 932 3099 982 3128
rect 1145 3147 1195 3176
rect 1145 3123 1156 3147
rect 1180 3123 1195 3147
rect 1145 3099 1195 3123
rect 1353 3152 1403 3176
rect 1353 3128 1365 3152
rect 1389 3128 1403 3152
rect 1353 3099 1403 3128
rect 1561 3150 1611 3176
rect 11640 3270 11690 3283
rect 11853 3270 11903 3283
rect 12061 3270 12111 3283
rect 12269 3270 12319 3283
rect 6727 3233 6777 3249
rect 6935 3233 6985 3249
rect 7143 3233 7193 3249
rect 7356 3233 7406 3249
rect 9222 3228 9272 3244
rect 9430 3228 9480 3244
rect 9638 3228 9688 3244
rect 9851 3228 9901 3244
rect 1561 3124 1579 3150
rect 1605 3124 1611 3150
rect 1561 3099 1611 3124
rect 1980 3144 2030 3172
rect 1980 3124 1993 3144
rect 2013 3124 2030 3144
rect 1980 3095 2030 3124
rect 2193 3143 2243 3172
rect 2193 3119 2204 3143
rect 2228 3119 2243 3143
rect 2193 3095 2243 3119
rect 2401 3148 2451 3172
rect 2401 3124 2413 3148
rect 2437 3124 2451 3148
rect 2401 3095 2451 3124
rect 2609 3146 2659 3172
rect 2609 3120 2627 3146
rect 2653 3120 2659 3146
rect 2609 3095 2659 3120
rect 6727 3166 6777 3191
rect 6727 3140 6733 3166
rect 6759 3140 6777 3166
rect 6727 3114 6777 3140
rect 6935 3162 6985 3191
rect 6935 3138 6949 3162
rect 6973 3138 6985 3162
rect 6935 3114 6985 3138
rect 7143 3167 7193 3191
rect 7143 3143 7158 3167
rect 7182 3143 7193 3167
rect 7143 3114 7193 3143
rect 7356 3162 7406 3191
rect 7356 3142 7373 3162
rect 7393 3142 7406 3162
rect 7356 3114 7406 3142
rect 9222 3161 9272 3186
rect 9222 3135 9228 3161
rect 9254 3135 9272 3161
rect 932 3041 982 3057
rect 1145 3041 1195 3057
rect 1353 3041 1403 3057
rect 1561 3041 1611 3057
rect 1980 3037 2030 3053
rect 2193 3037 2243 3053
rect 2401 3037 2451 3053
rect 2609 3037 2659 3053
rect 9222 3109 9272 3135
rect 9430 3157 9480 3186
rect 9430 3133 9444 3157
rect 9468 3133 9480 3157
rect 9430 3109 9480 3133
rect 9638 3162 9688 3186
rect 9638 3138 9653 3162
rect 9677 3138 9688 3162
rect 9638 3109 9688 3138
rect 9851 3157 9901 3186
rect 9851 3137 9868 3157
rect 9888 3137 9901 3157
rect 12688 3266 12738 3279
rect 12901 3266 12951 3279
rect 13109 3266 13159 3279
rect 13317 3266 13367 3279
rect 9851 3109 9901 3137
rect 6727 3001 6777 3014
rect 6935 3001 6985 3014
rect 7143 3001 7193 3014
rect 7356 3001 7406 3014
rect 11640 3142 11690 3170
rect 11640 3122 11653 3142
rect 11673 3122 11690 3142
rect 11640 3093 11690 3122
rect 11853 3141 11903 3170
rect 11853 3117 11864 3141
rect 11888 3117 11903 3141
rect 11853 3093 11903 3117
rect 12061 3146 12111 3170
rect 12061 3122 12073 3146
rect 12097 3122 12111 3146
rect 12061 3093 12111 3122
rect 12269 3144 12319 3170
rect 22605 3274 22655 3287
rect 22818 3274 22868 3287
rect 23026 3274 23076 3287
rect 23234 3274 23284 3287
rect 17435 3227 17485 3243
rect 17643 3227 17693 3243
rect 17851 3227 17901 3243
rect 18064 3227 18114 3243
rect 19930 3222 19980 3238
rect 20138 3222 20188 3238
rect 20346 3222 20396 3238
rect 20559 3222 20609 3238
rect 12269 3118 12287 3144
rect 12313 3118 12319 3144
rect 12269 3093 12319 3118
rect 12688 3138 12738 3166
rect 12688 3118 12701 3138
rect 12721 3118 12738 3138
rect 12688 3089 12738 3118
rect 12901 3137 12951 3166
rect 12901 3113 12912 3137
rect 12936 3113 12951 3137
rect 12901 3089 12951 3113
rect 13109 3142 13159 3166
rect 13109 3118 13121 3142
rect 13145 3118 13159 3142
rect 13109 3089 13159 3118
rect 13317 3140 13367 3166
rect 13317 3114 13335 3140
rect 13361 3114 13367 3140
rect 13317 3089 13367 3114
rect 17435 3160 17485 3185
rect 17435 3134 17441 3160
rect 17467 3134 17485 3160
rect 17435 3108 17485 3134
rect 17643 3156 17693 3185
rect 17643 3132 17657 3156
rect 17681 3132 17693 3156
rect 17643 3108 17693 3132
rect 17851 3161 17901 3185
rect 17851 3137 17866 3161
rect 17890 3137 17901 3161
rect 17851 3108 17901 3137
rect 18064 3156 18114 3185
rect 18064 3136 18081 3156
rect 18101 3136 18114 3156
rect 18064 3108 18114 3136
rect 19930 3155 19980 3180
rect 19930 3129 19936 3155
rect 19962 3129 19980 3155
rect 11640 3035 11690 3051
rect 11853 3035 11903 3051
rect 12061 3035 12111 3051
rect 12269 3035 12319 3051
rect 12688 3031 12738 3047
rect 12901 3031 12951 3047
rect 13109 3031 13159 3047
rect 13317 3031 13367 3047
rect 9222 2996 9272 3009
rect 9430 2996 9480 3009
rect 9638 2996 9688 3009
rect 9851 2996 9901 3009
rect 19930 3103 19980 3129
rect 20138 3151 20188 3180
rect 20138 3127 20152 3151
rect 20176 3127 20188 3151
rect 20138 3103 20188 3127
rect 20346 3156 20396 3180
rect 20346 3132 20361 3156
rect 20385 3132 20396 3156
rect 20346 3103 20396 3132
rect 20559 3151 20609 3180
rect 23653 3270 23703 3283
rect 23866 3270 23916 3283
rect 24074 3270 24124 3283
rect 24282 3270 24332 3283
rect 20559 3131 20576 3151
rect 20596 3131 20609 3151
rect 20559 3103 20609 3131
rect 17435 2995 17485 3008
rect 17643 2995 17693 3008
rect 17851 2995 17901 3008
rect 18064 2995 18114 3008
rect 22605 3146 22655 3174
rect 22605 3126 22618 3146
rect 22638 3126 22655 3146
rect 22605 3097 22655 3126
rect 22818 3145 22868 3174
rect 22818 3121 22829 3145
rect 22853 3121 22868 3145
rect 22818 3097 22868 3121
rect 23026 3150 23076 3174
rect 23026 3126 23038 3150
rect 23062 3126 23076 3150
rect 23026 3097 23076 3126
rect 23234 3148 23284 3174
rect 33313 3268 33363 3281
rect 33526 3268 33576 3281
rect 33734 3268 33784 3281
rect 33942 3268 33992 3281
rect 28400 3231 28450 3247
rect 28608 3231 28658 3247
rect 28816 3231 28866 3247
rect 29029 3231 29079 3247
rect 30895 3226 30945 3242
rect 31103 3226 31153 3242
rect 31311 3226 31361 3242
rect 31524 3226 31574 3242
rect 23234 3122 23252 3148
rect 23278 3122 23284 3148
rect 23234 3097 23284 3122
rect 23653 3142 23703 3170
rect 23653 3122 23666 3142
rect 23686 3122 23703 3142
rect 23653 3093 23703 3122
rect 23866 3141 23916 3170
rect 23866 3117 23877 3141
rect 23901 3117 23916 3141
rect 23866 3093 23916 3117
rect 24074 3146 24124 3170
rect 24074 3122 24086 3146
rect 24110 3122 24124 3146
rect 24074 3093 24124 3122
rect 24282 3144 24332 3170
rect 24282 3118 24300 3144
rect 24326 3118 24332 3144
rect 24282 3093 24332 3118
rect 28400 3164 28450 3189
rect 28400 3138 28406 3164
rect 28432 3138 28450 3164
rect 28400 3112 28450 3138
rect 28608 3160 28658 3189
rect 28608 3136 28622 3160
rect 28646 3136 28658 3160
rect 28608 3112 28658 3136
rect 28816 3165 28866 3189
rect 28816 3141 28831 3165
rect 28855 3141 28866 3165
rect 28816 3112 28866 3141
rect 29029 3160 29079 3189
rect 29029 3140 29046 3160
rect 29066 3140 29079 3160
rect 29029 3112 29079 3140
rect 30895 3159 30945 3184
rect 30895 3133 30901 3159
rect 30927 3133 30945 3159
rect 22605 3039 22655 3055
rect 22818 3039 22868 3055
rect 23026 3039 23076 3055
rect 23234 3039 23284 3055
rect 23653 3035 23703 3051
rect 23866 3035 23916 3051
rect 24074 3035 24124 3051
rect 24282 3035 24332 3051
rect 19930 2990 19980 3003
rect 20138 2990 20188 3003
rect 20346 2990 20396 3003
rect 20559 2990 20609 3003
rect 30895 3107 30945 3133
rect 31103 3155 31153 3184
rect 31103 3131 31117 3155
rect 31141 3131 31153 3155
rect 31103 3107 31153 3131
rect 31311 3160 31361 3184
rect 31311 3136 31326 3160
rect 31350 3136 31361 3160
rect 31311 3107 31361 3136
rect 31524 3155 31574 3184
rect 31524 3135 31541 3155
rect 31561 3135 31574 3155
rect 34361 3264 34411 3277
rect 34574 3264 34624 3277
rect 34782 3264 34832 3277
rect 34990 3264 35040 3277
rect 31524 3107 31574 3135
rect 28400 2999 28450 3012
rect 28608 2999 28658 3012
rect 28816 2999 28866 3012
rect 29029 2999 29079 3012
rect 33313 3140 33363 3168
rect 33313 3120 33326 3140
rect 33346 3120 33363 3140
rect 33313 3091 33363 3120
rect 33526 3139 33576 3168
rect 33526 3115 33537 3139
rect 33561 3115 33576 3139
rect 33526 3091 33576 3115
rect 33734 3144 33784 3168
rect 33734 3120 33746 3144
rect 33770 3120 33784 3144
rect 33734 3091 33784 3120
rect 33942 3142 33992 3168
rect 39108 3225 39158 3241
rect 39316 3225 39366 3241
rect 39524 3225 39574 3241
rect 39737 3225 39787 3241
rect 41603 3220 41653 3236
rect 41811 3220 41861 3236
rect 42019 3220 42069 3236
rect 42232 3220 42282 3236
rect 33942 3116 33960 3142
rect 33986 3116 33992 3142
rect 33942 3091 33992 3116
rect 34361 3136 34411 3164
rect 34361 3116 34374 3136
rect 34394 3116 34411 3136
rect 34361 3087 34411 3116
rect 34574 3135 34624 3164
rect 34574 3111 34585 3135
rect 34609 3111 34624 3135
rect 34574 3087 34624 3111
rect 34782 3140 34832 3164
rect 34782 3116 34794 3140
rect 34818 3116 34832 3140
rect 34782 3087 34832 3116
rect 34990 3138 35040 3164
rect 34990 3112 35008 3138
rect 35034 3112 35040 3138
rect 34990 3087 35040 3112
rect 39108 3158 39158 3183
rect 39108 3132 39114 3158
rect 39140 3132 39158 3158
rect 39108 3106 39158 3132
rect 39316 3154 39366 3183
rect 39316 3130 39330 3154
rect 39354 3130 39366 3154
rect 39316 3106 39366 3130
rect 39524 3159 39574 3183
rect 39524 3135 39539 3159
rect 39563 3135 39574 3159
rect 39524 3106 39574 3135
rect 39737 3154 39787 3183
rect 39737 3134 39754 3154
rect 39774 3134 39787 3154
rect 39737 3106 39787 3134
rect 41603 3153 41653 3178
rect 41603 3127 41609 3153
rect 41635 3127 41653 3153
rect 33313 3033 33363 3049
rect 33526 3033 33576 3049
rect 33734 3033 33784 3049
rect 33942 3033 33992 3049
rect 34361 3029 34411 3045
rect 34574 3029 34624 3045
rect 34782 3029 34832 3045
rect 34990 3029 35040 3045
rect 30895 2994 30945 3007
rect 31103 2994 31153 3007
rect 31311 2994 31361 3007
rect 31524 2994 31574 3007
rect 41603 3101 41653 3127
rect 41811 3149 41861 3178
rect 41811 3125 41825 3149
rect 41849 3125 41861 3149
rect 41811 3101 41861 3125
rect 42019 3154 42069 3178
rect 42019 3130 42034 3154
rect 42058 3130 42069 3154
rect 42019 3101 42069 3130
rect 42232 3149 42282 3178
rect 42232 3129 42249 3149
rect 42269 3129 42282 3149
rect 42232 3101 42282 3129
rect 39108 2993 39158 3006
rect 39316 2993 39366 3006
rect 39524 2993 39574 3006
rect 39737 2993 39787 3006
rect 41603 2988 41653 3001
rect 41811 2988 41861 3001
rect 42019 2988 42069 3001
rect 42232 2988 42282 3001
rect 932 2597 982 2610
rect 1145 2597 1195 2610
rect 1353 2597 1403 2610
rect 1561 2597 1611 2610
rect 11640 2591 11690 2604
rect 11853 2591 11903 2604
rect 12061 2591 12111 2604
rect 12269 2591 12319 2604
rect 8174 2553 8224 2569
rect 8382 2553 8432 2569
rect 8590 2553 8640 2569
rect 8803 2553 8853 2569
rect 9222 2549 9272 2565
rect 9430 2549 9480 2565
rect 9638 2549 9688 2565
rect 9851 2549 9901 2565
rect 932 2469 982 2497
rect 932 2449 945 2469
rect 965 2449 982 2469
rect 932 2420 982 2449
rect 1145 2468 1195 2497
rect 1145 2444 1156 2468
rect 1180 2444 1195 2468
rect 1145 2420 1195 2444
rect 1353 2473 1403 2497
rect 1353 2449 1365 2473
rect 1389 2449 1403 2473
rect 1353 2420 1403 2449
rect 1561 2471 1611 2497
rect 1561 2445 1579 2471
rect 1605 2445 1611 2471
rect 1561 2420 1611 2445
rect 8174 2486 8224 2511
rect 8174 2460 8180 2486
rect 8206 2460 8224 2486
rect 8174 2434 8224 2460
rect 8382 2482 8432 2511
rect 8382 2458 8396 2482
rect 8420 2458 8432 2482
rect 8382 2434 8432 2458
rect 8590 2487 8640 2511
rect 8590 2463 8605 2487
rect 8629 2463 8640 2487
rect 8590 2434 8640 2463
rect 8803 2482 8853 2511
rect 8803 2462 8820 2482
rect 8840 2462 8853 2482
rect 8803 2434 8853 2462
rect 9222 2482 9272 2507
rect 9222 2456 9228 2482
rect 9254 2456 9272 2482
rect 932 2362 982 2378
rect 1145 2362 1195 2378
rect 1353 2362 1403 2378
rect 1561 2362 1611 2378
rect 9222 2430 9272 2456
rect 9430 2478 9480 2507
rect 9430 2454 9444 2478
rect 9468 2454 9480 2478
rect 9430 2430 9480 2454
rect 9638 2483 9688 2507
rect 9638 2459 9653 2483
rect 9677 2459 9688 2483
rect 9638 2430 9688 2459
rect 9851 2478 9901 2507
rect 9851 2458 9868 2478
rect 9888 2458 9901 2478
rect 9851 2430 9901 2458
rect 22605 2595 22655 2608
rect 22818 2595 22868 2608
rect 23026 2595 23076 2608
rect 23234 2595 23284 2608
rect 18882 2547 18932 2563
rect 19090 2547 19140 2563
rect 19298 2547 19348 2563
rect 19511 2547 19561 2563
rect 19930 2543 19980 2559
rect 20138 2543 20188 2559
rect 20346 2543 20396 2559
rect 20559 2543 20609 2559
rect 11640 2463 11690 2491
rect 8174 2321 8224 2334
rect 8382 2321 8432 2334
rect 8590 2321 8640 2334
rect 8803 2321 8853 2334
rect 11640 2443 11653 2463
rect 11673 2443 11690 2463
rect 11640 2414 11690 2443
rect 11853 2462 11903 2491
rect 11853 2438 11864 2462
rect 11888 2438 11903 2462
rect 11853 2414 11903 2438
rect 12061 2467 12111 2491
rect 12061 2443 12073 2467
rect 12097 2443 12111 2467
rect 12061 2414 12111 2443
rect 12269 2465 12319 2491
rect 12269 2439 12287 2465
rect 12313 2439 12319 2465
rect 12269 2414 12319 2439
rect 18882 2480 18932 2505
rect 18882 2454 18888 2480
rect 18914 2454 18932 2480
rect 18882 2428 18932 2454
rect 19090 2476 19140 2505
rect 19090 2452 19104 2476
rect 19128 2452 19140 2476
rect 19090 2428 19140 2452
rect 19298 2481 19348 2505
rect 19298 2457 19313 2481
rect 19337 2457 19348 2481
rect 19298 2428 19348 2457
rect 19511 2476 19561 2505
rect 19511 2456 19528 2476
rect 19548 2456 19561 2476
rect 19511 2428 19561 2456
rect 19930 2476 19980 2501
rect 19930 2450 19936 2476
rect 19962 2450 19980 2476
rect 11640 2356 11690 2372
rect 11853 2356 11903 2372
rect 12061 2356 12111 2372
rect 12269 2356 12319 2372
rect 9222 2317 9272 2330
rect 9430 2317 9480 2330
rect 9638 2317 9688 2330
rect 9851 2317 9901 2330
rect 19930 2424 19980 2450
rect 20138 2472 20188 2501
rect 20138 2448 20152 2472
rect 20176 2448 20188 2472
rect 20138 2424 20188 2448
rect 20346 2477 20396 2501
rect 20346 2453 20361 2477
rect 20385 2453 20396 2477
rect 20346 2424 20396 2453
rect 20559 2472 20609 2501
rect 20559 2452 20576 2472
rect 20596 2452 20609 2472
rect 20559 2424 20609 2452
rect 33313 2589 33363 2602
rect 33526 2589 33576 2602
rect 33734 2589 33784 2602
rect 33942 2589 33992 2602
rect 29847 2551 29897 2567
rect 30055 2551 30105 2567
rect 30263 2551 30313 2567
rect 30476 2551 30526 2567
rect 30895 2547 30945 2563
rect 31103 2547 31153 2563
rect 31311 2547 31361 2563
rect 31524 2547 31574 2563
rect 22605 2467 22655 2495
rect 22605 2447 22618 2467
rect 22638 2447 22655 2467
rect 18882 2315 18932 2328
rect 19090 2315 19140 2328
rect 19298 2315 19348 2328
rect 19511 2315 19561 2328
rect 22605 2418 22655 2447
rect 22818 2466 22868 2495
rect 22818 2442 22829 2466
rect 22853 2442 22868 2466
rect 22818 2418 22868 2442
rect 23026 2471 23076 2495
rect 23026 2447 23038 2471
rect 23062 2447 23076 2471
rect 23026 2418 23076 2447
rect 23234 2469 23284 2495
rect 23234 2443 23252 2469
rect 23278 2443 23284 2469
rect 23234 2418 23284 2443
rect 29847 2484 29897 2509
rect 29847 2458 29853 2484
rect 29879 2458 29897 2484
rect 29847 2432 29897 2458
rect 30055 2480 30105 2509
rect 30055 2456 30069 2480
rect 30093 2456 30105 2480
rect 30055 2432 30105 2456
rect 30263 2485 30313 2509
rect 30263 2461 30278 2485
rect 30302 2461 30313 2485
rect 30263 2432 30313 2461
rect 30476 2480 30526 2509
rect 30476 2460 30493 2480
rect 30513 2460 30526 2480
rect 30476 2432 30526 2460
rect 30895 2480 30945 2505
rect 30895 2454 30901 2480
rect 30927 2454 30945 2480
rect 22605 2360 22655 2376
rect 22818 2360 22868 2376
rect 23026 2360 23076 2376
rect 23234 2360 23284 2376
rect 19930 2311 19980 2324
rect 20138 2311 20188 2324
rect 20346 2311 20396 2324
rect 20559 2311 20609 2324
rect 30895 2428 30945 2454
rect 31103 2476 31153 2505
rect 31103 2452 31117 2476
rect 31141 2452 31153 2476
rect 31103 2428 31153 2452
rect 31311 2481 31361 2505
rect 31311 2457 31326 2481
rect 31350 2457 31361 2481
rect 31311 2428 31361 2457
rect 31524 2476 31574 2505
rect 31524 2456 31541 2476
rect 31561 2456 31574 2476
rect 31524 2428 31574 2456
rect 40555 2545 40605 2561
rect 40763 2545 40813 2561
rect 40971 2545 41021 2561
rect 41184 2545 41234 2561
rect 41603 2541 41653 2557
rect 41811 2541 41861 2557
rect 42019 2541 42069 2557
rect 42232 2541 42282 2557
rect 33313 2461 33363 2489
rect 29847 2319 29897 2332
rect 30055 2319 30105 2332
rect 30263 2319 30313 2332
rect 30476 2319 30526 2332
rect 33313 2441 33326 2461
rect 33346 2441 33363 2461
rect 33313 2412 33363 2441
rect 33526 2460 33576 2489
rect 33526 2436 33537 2460
rect 33561 2436 33576 2460
rect 33526 2412 33576 2436
rect 33734 2465 33784 2489
rect 33734 2441 33746 2465
rect 33770 2441 33784 2465
rect 33734 2412 33784 2441
rect 33942 2463 33992 2489
rect 33942 2437 33960 2463
rect 33986 2437 33992 2463
rect 33942 2412 33992 2437
rect 40555 2478 40605 2503
rect 40555 2452 40561 2478
rect 40587 2452 40605 2478
rect 40555 2426 40605 2452
rect 40763 2474 40813 2503
rect 40763 2450 40777 2474
rect 40801 2450 40813 2474
rect 40763 2426 40813 2450
rect 40971 2479 41021 2503
rect 40971 2455 40986 2479
rect 41010 2455 41021 2479
rect 40971 2426 41021 2455
rect 41184 2474 41234 2503
rect 41184 2454 41201 2474
rect 41221 2454 41234 2474
rect 41184 2426 41234 2454
rect 41603 2474 41653 2499
rect 41603 2448 41609 2474
rect 41635 2448 41653 2474
rect 33313 2354 33363 2370
rect 33526 2354 33576 2370
rect 33734 2354 33784 2370
rect 33942 2354 33992 2370
rect 30895 2315 30945 2328
rect 31103 2315 31153 2328
rect 31311 2315 31361 2328
rect 31524 2315 31574 2328
rect 41603 2422 41653 2448
rect 41811 2470 41861 2499
rect 41811 2446 41825 2470
rect 41849 2446 41861 2470
rect 41811 2422 41861 2446
rect 42019 2475 42069 2499
rect 42019 2451 42034 2475
rect 42058 2451 42069 2475
rect 42019 2422 42069 2451
rect 42232 2470 42282 2499
rect 42232 2450 42249 2470
rect 42269 2450 42282 2470
rect 42232 2422 42282 2450
rect 40555 2313 40605 2326
rect 40763 2313 40813 2326
rect 40971 2313 41021 2326
rect 41184 2313 41234 2326
rect 41603 2309 41653 2322
rect 41811 2309 41861 2322
rect 42019 2309 42069 2322
rect 42232 2309 42282 2322
rect 10643 438 10693 451
rect 10856 438 10906 451
rect 11064 438 11114 451
rect 11272 438 11322 451
rect 21280 425 21330 438
rect 21493 425 21543 438
rect 21701 425 21751 438
rect 21909 425 21959 438
rect 32316 436 32366 449
rect 32529 436 32579 449
rect 32737 436 32787 449
rect 32945 436 32995 449
rect 10643 310 10693 338
rect 10643 290 10656 310
rect 10676 290 10693 310
rect 10643 261 10693 290
rect 10856 309 10906 338
rect 10856 285 10867 309
rect 10891 285 10906 309
rect 10856 261 10906 285
rect 11064 314 11114 338
rect 11064 290 11076 314
rect 11100 290 11114 314
rect 11064 261 11114 290
rect 11272 312 11322 338
rect 11272 286 11290 312
rect 11316 286 11322 312
rect 11272 261 11322 286
rect 21280 297 21330 325
rect 21280 277 21293 297
rect 21313 277 21330 297
rect 21280 248 21330 277
rect 21493 296 21543 325
rect 21493 272 21504 296
rect 21528 272 21543 296
rect 21493 248 21543 272
rect 21701 301 21751 325
rect 21701 277 21713 301
rect 21737 277 21751 301
rect 21701 248 21751 277
rect 21909 299 21959 325
rect 21909 273 21927 299
rect 21953 273 21959 299
rect 21909 248 21959 273
rect 32316 308 32366 336
rect 32316 288 32329 308
rect 32349 288 32366 308
rect 32316 259 32366 288
rect 32529 307 32579 336
rect 32529 283 32540 307
rect 32564 283 32579 307
rect 32529 259 32579 283
rect 32737 312 32787 336
rect 32737 288 32749 312
rect 32773 288 32787 312
rect 32737 259 32787 288
rect 32945 310 32995 336
rect 32945 284 32963 310
rect 32989 284 32995 310
rect 32945 259 32995 284
rect 10643 203 10693 219
rect 10856 203 10906 219
rect 11064 203 11114 219
rect 11272 203 11322 219
rect 21280 190 21330 206
rect 21493 190 21543 206
rect 21701 190 21751 206
rect 21909 190 21959 206
rect 32316 201 32366 217
rect 32529 201 32579 217
rect 32737 201 32787 217
rect 32945 201 32995 217
<< polycont >>
rect 946 13550 966 13570
rect 1157 13545 1181 13569
rect 1366 13550 1390 13574
rect 1580 13546 1606 13572
rect 1994 13546 2014 13566
rect 2205 13541 2229 13565
rect 2414 13546 2438 13570
rect 2628 13542 2654 13568
rect 9229 13557 9255 13583
rect 9445 13555 9469 13579
rect 9654 13560 9678 13584
rect 9869 13559 9889 13579
rect 11654 13544 11674 13564
rect 11865 13539 11889 13563
rect 12074 13544 12098 13568
rect 12288 13540 12314 13566
rect 12702 13540 12722 13560
rect 12913 13535 12937 13559
rect 13122 13540 13146 13564
rect 13336 13536 13362 13562
rect 19937 13551 19963 13577
rect 20153 13549 20177 13573
rect 20362 13554 20386 13578
rect 20577 13553 20597 13573
rect 22619 13548 22639 13568
rect 22830 13543 22854 13567
rect 23039 13548 23063 13572
rect 23253 13544 23279 13570
rect 23667 13544 23687 13564
rect 23878 13539 23902 13563
rect 24087 13544 24111 13568
rect 24301 13540 24327 13566
rect 30902 13555 30928 13581
rect 31118 13553 31142 13577
rect 31327 13558 31351 13582
rect 31542 13557 31562 13577
rect 33327 13542 33347 13562
rect 33538 13537 33562 13561
rect 33747 13542 33771 13566
rect 33961 13538 33987 13564
rect 34375 13538 34395 13558
rect 34586 13533 34610 13557
rect 34795 13538 34819 13562
rect 35009 13534 35035 13560
rect 41610 13549 41636 13575
rect 41826 13547 41850 13571
rect 42035 13552 42059 13576
rect 42250 13551 42270 13571
rect 946 12871 966 12891
rect 1157 12866 1181 12890
rect 1366 12871 1390 12895
rect 1580 12867 1606 12893
rect 3441 12866 3461 12886
rect 3652 12861 3676 12885
rect 3861 12866 3885 12890
rect 4075 12862 4101 12888
rect 8181 12882 8207 12908
rect 8397 12880 8421 12904
rect 8606 12885 8630 12909
rect 8821 12884 8841 12904
rect 9229 12878 9255 12904
rect 9445 12876 9469 12900
rect 9654 12881 9678 12905
rect 9869 12880 9889 12900
rect 11654 12865 11674 12885
rect 11865 12860 11889 12884
rect 12074 12865 12098 12889
rect 12288 12861 12314 12887
rect 14149 12860 14169 12880
rect 14360 12855 14384 12879
rect 14569 12860 14593 12884
rect 14783 12856 14809 12882
rect 18889 12876 18915 12902
rect 19105 12874 19129 12898
rect 19314 12879 19338 12903
rect 19529 12878 19549 12898
rect 19937 12872 19963 12898
rect 20153 12870 20177 12894
rect 20362 12875 20386 12899
rect 20577 12874 20597 12894
rect 22619 12869 22639 12889
rect 22830 12864 22854 12888
rect 23039 12869 23063 12893
rect 23253 12865 23279 12891
rect 25114 12864 25134 12884
rect 25325 12859 25349 12883
rect 25534 12864 25558 12888
rect 25748 12860 25774 12886
rect 29854 12880 29880 12906
rect 30070 12878 30094 12902
rect 30279 12883 30303 12907
rect 30494 12882 30514 12902
rect 30902 12876 30928 12902
rect 31118 12874 31142 12898
rect 31327 12879 31351 12903
rect 31542 12878 31562 12898
rect 33327 12863 33347 12883
rect 33538 12858 33562 12882
rect 33747 12863 33771 12887
rect 33961 12859 33987 12885
rect 35822 12858 35842 12878
rect 36033 12853 36057 12877
rect 36242 12858 36266 12882
rect 36456 12854 36482 12880
rect 40562 12874 40588 12900
rect 40778 12872 40802 12896
rect 40987 12877 41011 12901
rect 41202 12876 41222 12896
rect 41610 12870 41636 12896
rect 41826 12868 41850 12892
rect 42035 12873 42059 12897
rect 42250 12872 42270 12892
rect 946 12103 966 12123
rect 1157 12098 1181 12122
rect 1366 12103 1390 12127
rect 1580 12099 1606 12125
rect 1994 12099 2014 12119
rect 2205 12094 2229 12118
rect 2414 12099 2438 12123
rect 2628 12095 2654 12121
rect 6734 12115 6760 12141
rect 6950 12113 6974 12137
rect 7159 12118 7183 12142
rect 7374 12117 7394 12137
rect 9229 12110 9255 12136
rect 9445 12108 9469 12132
rect 9654 12113 9678 12137
rect 9869 12112 9889 12132
rect 11654 12097 11674 12117
rect 11865 12092 11889 12116
rect 12074 12097 12098 12121
rect 12288 12093 12314 12119
rect 12702 12093 12722 12113
rect 12913 12088 12937 12112
rect 13122 12093 13146 12117
rect 13336 12089 13362 12115
rect 17442 12109 17468 12135
rect 17658 12107 17682 12131
rect 17867 12112 17891 12136
rect 18082 12111 18102 12131
rect 19937 12104 19963 12130
rect 20153 12102 20177 12126
rect 20362 12107 20386 12131
rect 20577 12106 20597 12126
rect 22619 12101 22639 12121
rect 22830 12096 22854 12120
rect 23039 12101 23063 12125
rect 23253 12097 23279 12123
rect 23667 12097 23687 12117
rect 23878 12092 23902 12116
rect 24087 12097 24111 12121
rect 24301 12093 24327 12119
rect 28407 12113 28433 12139
rect 28623 12111 28647 12135
rect 28832 12116 28856 12140
rect 29047 12115 29067 12135
rect 30902 12108 30928 12134
rect 31118 12106 31142 12130
rect 31327 12111 31351 12135
rect 31542 12110 31562 12130
rect 33327 12095 33347 12115
rect 33538 12090 33562 12114
rect 33747 12095 33771 12119
rect 33961 12091 33987 12117
rect 34375 12091 34395 12111
rect 34586 12086 34610 12110
rect 34795 12091 34819 12115
rect 35009 12087 35035 12113
rect 39115 12107 39141 12133
rect 39331 12105 39355 12129
rect 39540 12110 39564 12134
rect 39755 12109 39775 12129
rect 41610 12102 41636 12128
rect 41826 12100 41850 12124
rect 42035 12105 42059 12129
rect 42250 12104 42270 12124
rect 946 11424 966 11444
rect 1157 11419 1181 11443
rect 1366 11424 1390 11448
rect 1580 11420 1606 11446
rect 3484 11421 3504 11441
rect 3695 11416 3719 11440
rect 3904 11421 3928 11445
rect 4118 11417 4144 11443
rect 8181 11435 8207 11461
rect 8397 11433 8421 11457
rect 8606 11438 8630 11462
rect 8821 11437 8841 11457
rect 9229 11431 9255 11457
rect 9445 11429 9469 11453
rect 9654 11434 9678 11458
rect 9869 11433 9889 11453
rect 11654 11418 11674 11438
rect 11865 11413 11889 11437
rect 12074 11418 12098 11442
rect 12288 11414 12314 11440
rect 14192 11415 14212 11435
rect 14403 11410 14427 11434
rect 14612 11415 14636 11439
rect 14826 11411 14852 11437
rect 18889 11429 18915 11455
rect 19105 11427 19129 11451
rect 19314 11432 19338 11456
rect 19529 11431 19549 11451
rect 19937 11425 19963 11451
rect 20153 11423 20177 11447
rect 20362 11428 20386 11452
rect 20577 11427 20597 11447
rect 22619 11422 22639 11442
rect 22830 11417 22854 11441
rect 23039 11422 23063 11446
rect 23253 11418 23279 11444
rect 25157 11419 25177 11439
rect 25368 11414 25392 11438
rect 25577 11419 25601 11443
rect 25791 11415 25817 11441
rect 29854 11433 29880 11459
rect 30070 11431 30094 11455
rect 30279 11436 30303 11460
rect 30494 11435 30514 11455
rect 30902 11429 30928 11455
rect 31118 11427 31142 11451
rect 31327 11432 31351 11456
rect 31542 11431 31562 11451
rect 33327 11416 33347 11436
rect 33538 11411 33562 11435
rect 33747 11416 33771 11440
rect 33961 11412 33987 11438
rect 35865 11413 35885 11433
rect 36076 11408 36100 11432
rect 36285 11413 36309 11437
rect 36499 11409 36525 11435
rect 40562 11427 40588 11453
rect 40778 11425 40802 11449
rect 40987 11430 41011 11454
rect 41202 11429 41222 11449
rect 41610 11423 41636 11449
rect 41826 11421 41850 11445
rect 42035 11426 42059 11450
rect 42250 11425 42270 11445
rect 947 10583 967 10603
rect 1158 10578 1182 10602
rect 1367 10583 1391 10607
rect 1581 10579 1607 10605
rect 1995 10579 2015 10599
rect 2206 10574 2230 10598
rect 2415 10579 2439 10603
rect 2629 10575 2655 10601
rect 6692 10593 6718 10619
rect 6908 10591 6932 10615
rect 7117 10596 7141 10620
rect 7332 10595 7352 10615
rect 9230 10590 9256 10616
rect 9446 10588 9470 10612
rect 9655 10593 9679 10617
rect 9870 10592 9890 10612
rect 11655 10577 11675 10597
rect 11866 10572 11890 10596
rect 12075 10577 12099 10601
rect 12289 10573 12315 10599
rect 12703 10573 12723 10593
rect 12914 10568 12938 10592
rect 13123 10573 13147 10597
rect 13337 10569 13363 10595
rect 17400 10587 17426 10613
rect 17616 10585 17640 10609
rect 17825 10590 17849 10614
rect 18040 10589 18060 10609
rect 19938 10584 19964 10610
rect 20154 10582 20178 10606
rect 20363 10587 20387 10611
rect 20578 10586 20598 10606
rect 22620 10581 22640 10601
rect 22831 10576 22855 10600
rect 23040 10581 23064 10605
rect 23254 10577 23280 10603
rect 23668 10577 23688 10597
rect 23879 10572 23903 10596
rect 24088 10577 24112 10601
rect 24302 10573 24328 10599
rect 28365 10591 28391 10617
rect 28581 10589 28605 10613
rect 28790 10594 28814 10618
rect 29005 10593 29025 10613
rect 30903 10588 30929 10614
rect 31119 10586 31143 10610
rect 31328 10591 31352 10615
rect 31543 10590 31563 10610
rect 33328 10575 33348 10595
rect 33539 10570 33563 10594
rect 33748 10575 33772 10599
rect 33962 10571 33988 10597
rect 34376 10571 34396 10591
rect 34587 10566 34611 10590
rect 34796 10571 34820 10595
rect 35010 10567 35036 10593
rect 39073 10585 39099 10611
rect 39289 10583 39313 10607
rect 39498 10588 39522 10612
rect 39713 10587 39733 10607
rect 41611 10582 41637 10608
rect 41827 10580 41851 10604
rect 42036 10585 42060 10609
rect 42251 10584 42271 10604
rect 947 9904 967 9924
rect 1158 9899 1182 9923
rect 1367 9904 1391 9928
rect 1581 9900 1607 9926
rect 3442 9899 3462 9919
rect 3653 9894 3677 9918
rect 3862 9899 3886 9923
rect 4076 9895 4102 9921
rect 8182 9915 8208 9941
rect 8398 9913 8422 9937
rect 8607 9918 8631 9942
rect 8822 9917 8842 9937
rect 9230 9911 9256 9937
rect 9446 9909 9470 9933
rect 9655 9914 9679 9938
rect 9870 9913 9890 9933
rect 11655 9898 11675 9918
rect 11866 9893 11890 9917
rect 12075 9898 12099 9922
rect 12289 9894 12315 9920
rect 14150 9893 14170 9913
rect 14361 9888 14385 9912
rect 14570 9893 14594 9917
rect 14784 9889 14810 9915
rect 18890 9909 18916 9935
rect 19106 9907 19130 9931
rect 19315 9912 19339 9936
rect 19530 9911 19550 9931
rect 19938 9905 19964 9931
rect 20154 9903 20178 9927
rect 20363 9908 20387 9932
rect 20578 9907 20598 9927
rect 22620 9902 22640 9922
rect 22831 9897 22855 9921
rect 23040 9902 23064 9926
rect 23254 9898 23280 9924
rect 25115 9897 25135 9917
rect 25326 9892 25350 9916
rect 25535 9897 25559 9921
rect 25749 9893 25775 9919
rect 29855 9913 29881 9939
rect 30071 9911 30095 9935
rect 30280 9916 30304 9940
rect 30495 9915 30515 9935
rect 30903 9909 30929 9935
rect 31119 9907 31143 9931
rect 31328 9912 31352 9936
rect 31543 9911 31563 9931
rect 33328 9896 33348 9916
rect 33539 9891 33563 9915
rect 33748 9896 33772 9920
rect 33962 9892 33988 9918
rect 35823 9891 35843 9911
rect 36034 9886 36058 9910
rect 36243 9891 36267 9915
rect 36457 9887 36483 9913
rect 40563 9907 40589 9933
rect 40779 9905 40803 9929
rect 40988 9910 41012 9934
rect 41203 9909 41223 9929
rect 41611 9903 41637 9929
rect 41827 9901 41851 9925
rect 42036 9906 42060 9930
rect 42251 9905 42271 9925
rect 947 9136 967 9156
rect 1158 9131 1182 9155
rect 1367 9136 1391 9160
rect 1581 9132 1607 9158
rect 1995 9132 2015 9152
rect 2206 9127 2230 9151
rect 2415 9132 2439 9156
rect 2629 9128 2655 9154
rect 6735 9148 6761 9174
rect 6951 9146 6975 9170
rect 7160 9151 7184 9175
rect 7375 9150 7395 9170
rect 9230 9143 9256 9169
rect 9446 9141 9470 9165
rect 9655 9146 9679 9170
rect 9870 9145 9890 9165
rect 11655 9130 11675 9150
rect 11866 9125 11890 9149
rect 12075 9130 12099 9154
rect 12289 9126 12315 9152
rect 12703 9126 12723 9146
rect 12914 9121 12938 9145
rect 13123 9126 13147 9150
rect 13337 9122 13363 9148
rect 17443 9142 17469 9168
rect 17659 9140 17683 9164
rect 17868 9145 17892 9169
rect 18083 9144 18103 9164
rect 19938 9137 19964 9163
rect 20154 9135 20178 9159
rect 20363 9140 20387 9164
rect 20578 9139 20598 9159
rect 22620 9134 22640 9154
rect 22831 9129 22855 9153
rect 23040 9134 23064 9158
rect 23254 9130 23280 9156
rect 23668 9130 23688 9150
rect 23879 9125 23903 9149
rect 24088 9130 24112 9154
rect 24302 9126 24328 9152
rect 28408 9146 28434 9172
rect 28624 9144 28648 9168
rect 28833 9149 28857 9173
rect 29048 9148 29068 9168
rect 30903 9141 30929 9167
rect 31119 9139 31143 9163
rect 31328 9144 31352 9168
rect 31543 9143 31563 9163
rect 33328 9128 33348 9148
rect 33539 9123 33563 9147
rect 33748 9128 33772 9152
rect 33962 9124 33988 9150
rect 34376 9124 34396 9144
rect 34587 9119 34611 9143
rect 34796 9124 34820 9148
rect 35010 9120 35036 9146
rect 39116 9140 39142 9166
rect 39332 9138 39356 9162
rect 39541 9143 39565 9167
rect 39756 9142 39776 9162
rect 41611 9135 41637 9161
rect 41827 9133 41851 9157
rect 42036 9138 42060 9162
rect 42251 9137 42271 9157
rect 947 8457 967 8477
rect 1158 8452 1182 8476
rect 1367 8457 1391 8481
rect 1581 8453 1607 8479
rect 4550 8448 4570 8468
rect 4761 8443 4785 8467
rect 4970 8448 4994 8472
rect 5184 8444 5210 8470
rect 8182 8468 8208 8494
rect 8398 8466 8422 8490
rect 8607 8471 8631 8495
rect 8822 8470 8842 8490
rect 9230 8464 9256 8490
rect 9446 8462 9470 8486
rect 9655 8467 9679 8491
rect 9870 8466 9890 8486
rect 11655 8451 11675 8471
rect 11866 8446 11890 8470
rect 12075 8451 12099 8475
rect 12289 8447 12315 8473
rect 15258 8442 15278 8462
rect 15469 8437 15493 8461
rect 15678 8442 15702 8466
rect 15892 8438 15918 8464
rect 18890 8462 18916 8488
rect 19106 8460 19130 8484
rect 19315 8465 19339 8489
rect 19530 8464 19550 8484
rect 19938 8458 19964 8484
rect 20154 8456 20178 8480
rect 20363 8461 20387 8485
rect 20578 8460 20598 8480
rect 22620 8455 22640 8475
rect 22831 8450 22855 8474
rect 23040 8455 23064 8479
rect 23254 8451 23280 8477
rect 26223 8446 26243 8466
rect 26434 8441 26458 8465
rect 26643 8446 26667 8470
rect 26857 8442 26883 8468
rect 29855 8466 29881 8492
rect 30071 8464 30095 8488
rect 30280 8469 30304 8493
rect 30495 8468 30515 8488
rect 30903 8462 30929 8488
rect 31119 8460 31143 8484
rect 31328 8465 31352 8489
rect 31543 8464 31563 8484
rect 33328 8449 33348 8469
rect 33539 8444 33563 8468
rect 33748 8449 33772 8473
rect 33962 8445 33988 8471
rect 36931 8440 36951 8460
rect 37142 8435 37166 8459
rect 37351 8440 37375 8464
rect 37565 8436 37591 8462
rect 40563 8460 40589 8486
rect 40779 8458 40803 8482
rect 40988 8463 41012 8487
rect 41203 8462 41223 8482
rect 41611 8456 41637 8482
rect 41827 8454 41851 8478
rect 42036 8459 42060 8483
rect 42251 8458 42271 8478
rect 944 7542 964 7562
rect 1155 7537 1179 7561
rect 1364 7542 1388 7566
rect 1578 7538 1604 7564
rect 1992 7538 2012 7558
rect 2203 7533 2227 7557
rect 2412 7538 2436 7562
rect 2626 7534 2652 7560
rect 5624 7558 5650 7584
rect 5840 7556 5864 7580
rect 6049 7561 6073 7585
rect 6264 7560 6284 7580
rect 9227 7549 9253 7575
rect 9443 7547 9467 7571
rect 9652 7552 9676 7576
rect 9867 7551 9887 7571
rect 11652 7536 11672 7556
rect 11863 7531 11887 7555
rect 12072 7536 12096 7560
rect 12286 7532 12312 7558
rect 12700 7532 12720 7552
rect 12911 7527 12935 7551
rect 13120 7532 13144 7556
rect 13334 7528 13360 7554
rect 16332 7552 16358 7578
rect 16548 7550 16572 7574
rect 16757 7555 16781 7579
rect 16972 7554 16992 7574
rect 19935 7543 19961 7569
rect 20151 7541 20175 7565
rect 20360 7546 20384 7570
rect 20575 7545 20595 7565
rect 22617 7540 22637 7560
rect 22828 7535 22852 7559
rect 23037 7540 23061 7564
rect 23251 7536 23277 7562
rect 23665 7536 23685 7556
rect 23876 7531 23900 7555
rect 24085 7536 24109 7560
rect 24299 7532 24325 7558
rect 27297 7556 27323 7582
rect 27513 7554 27537 7578
rect 27722 7559 27746 7583
rect 27937 7558 27957 7578
rect 30900 7547 30926 7573
rect 31116 7545 31140 7569
rect 31325 7550 31349 7574
rect 31540 7549 31560 7569
rect 33325 7534 33345 7554
rect 33536 7529 33560 7553
rect 33745 7534 33769 7558
rect 33959 7530 33985 7556
rect 34373 7530 34393 7550
rect 34584 7525 34608 7549
rect 34793 7530 34817 7554
rect 35007 7526 35033 7552
rect 38005 7550 38031 7576
rect 38221 7548 38245 7572
rect 38430 7553 38454 7577
rect 38645 7552 38665 7572
rect 41608 7541 41634 7567
rect 41824 7539 41848 7563
rect 42033 7544 42057 7568
rect 42248 7543 42268 7563
rect 944 6863 964 6883
rect 1155 6858 1179 6882
rect 1364 6863 1388 6887
rect 1578 6859 1604 6885
rect 3439 6858 3459 6878
rect 3650 6853 3674 6877
rect 3859 6858 3883 6882
rect 4073 6854 4099 6880
rect 8179 6874 8205 6900
rect 8395 6872 8419 6896
rect 8604 6877 8628 6901
rect 8819 6876 8839 6896
rect 9227 6870 9253 6896
rect 9443 6868 9467 6892
rect 9652 6873 9676 6897
rect 9867 6872 9887 6892
rect 11652 6857 11672 6877
rect 11863 6852 11887 6876
rect 12072 6857 12096 6881
rect 12286 6853 12312 6879
rect 14147 6852 14167 6872
rect 14358 6847 14382 6871
rect 14567 6852 14591 6876
rect 14781 6848 14807 6874
rect 18887 6868 18913 6894
rect 19103 6866 19127 6890
rect 19312 6871 19336 6895
rect 19527 6870 19547 6890
rect 19935 6864 19961 6890
rect 20151 6862 20175 6886
rect 20360 6867 20384 6891
rect 20575 6866 20595 6886
rect 22617 6861 22637 6881
rect 22828 6856 22852 6880
rect 23037 6861 23061 6885
rect 23251 6857 23277 6883
rect 25112 6856 25132 6876
rect 25323 6851 25347 6875
rect 25532 6856 25556 6880
rect 25746 6852 25772 6878
rect 29852 6872 29878 6898
rect 30068 6870 30092 6894
rect 30277 6875 30301 6899
rect 30492 6874 30512 6894
rect 30900 6868 30926 6894
rect 31116 6866 31140 6890
rect 31325 6871 31349 6895
rect 31540 6870 31560 6890
rect 33325 6855 33345 6875
rect 33536 6850 33560 6874
rect 33745 6855 33769 6879
rect 33959 6851 33985 6877
rect 35820 6850 35840 6870
rect 36031 6845 36055 6869
rect 36240 6850 36264 6874
rect 36454 6846 36480 6872
rect 40560 6866 40586 6892
rect 40776 6864 40800 6888
rect 40985 6869 41009 6893
rect 41200 6868 41220 6888
rect 41608 6862 41634 6888
rect 41824 6860 41848 6884
rect 42033 6865 42057 6889
rect 42248 6864 42268 6884
rect 944 6095 964 6115
rect 1155 6090 1179 6114
rect 1364 6095 1388 6119
rect 1578 6091 1604 6117
rect 1992 6091 2012 6111
rect 2203 6086 2227 6110
rect 2412 6091 2436 6115
rect 2626 6087 2652 6113
rect 6732 6107 6758 6133
rect 6948 6105 6972 6129
rect 7157 6110 7181 6134
rect 7372 6109 7392 6129
rect 9227 6102 9253 6128
rect 9443 6100 9467 6124
rect 9652 6105 9676 6129
rect 9867 6104 9887 6124
rect 11652 6089 11672 6109
rect 11863 6084 11887 6108
rect 12072 6089 12096 6113
rect 12286 6085 12312 6111
rect 12700 6085 12720 6105
rect 12911 6080 12935 6104
rect 13120 6085 13144 6109
rect 13334 6081 13360 6107
rect 17440 6101 17466 6127
rect 17656 6099 17680 6123
rect 17865 6104 17889 6128
rect 18080 6103 18100 6123
rect 19935 6096 19961 6122
rect 20151 6094 20175 6118
rect 20360 6099 20384 6123
rect 20575 6098 20595 6118
rect 22617 6093 22637 6113
rect 22828 6088 22852 6112
rect 23037 6093 23061 6117
rect 23251 6089 23277 6115
rect 23665 6089 23685 6109
rect 23876 6084 23900 6108
rect 24085 6089 24109 6113
rect 24299 6085 24325 6111
rect 28405 6105 28431 6131
rect 28621 6103 28645 6127
rect 28830 6108 28854 6132
rect 29045 6107 29065 6127
rect 30900 6100 30926 6126
rect 31116 6098 31140 6122
rect 31325 6103 31349 6127
rect 31540 6102 31560 6122
rect 33325 6087 33345 6107
rect 33536 6082 33560 6106
rect 33745 6087 33769 6111
rect 33959 6083 33985 6109
rect 34373 6083 34393 6103
rect 34584 6078 34608 6102
rect 34793 6083 34817 6107
rect 35007 6079 35033 6105
rect 39113 6099 39139 6125
rect 39329 6097 39353 6121
rect 39538 6102 39562 6126
rect 39753 6101 39773 6121
rect 41608 6094 41634 6120
rect 41824 6092 41848 6116
rect 42033 6097 42057 6121
rect 42248 6096 42268 6116
rect 944 5416 964 5436
rect 1155 5411 1179 5435
rect 1364 5416 1388 5440
rect 1578 5412 1604 5438
rect 3482 5413 3502 5433
rect 3693 5408 3717 5432
rect 3902 5413 3926 5437
rect 4116 5409 4142 5435
rect 8179 5427 8205 5453
rect 8395 5425 8419 5449
rect 8604 5430 8628 5454
rect 8819 5429 8839 5449
rect 9227 5423 9253 5449
rect 9443 5421 9467 5445
rect 9652 5426 9676 5450
rect 9867 5425 9887 5445
rect 11652 5410 11672 5430
rect 11863 5405 11887 5429
rect 12072 5410 12096 5434
rect 12286 5406 12312 5432
rect 14190 5407 14210 5427
rect 14401 5402 14425 5426
rect 14610 5407 14634 5431
rect 14824 5403 14850 5429
rect 18887 5421 18913 5447
rect 19103 5419 19127 5443
rect 19312 5424 19336 5448
rect 19527 5423 19547 5443
rect 19935 5417 19961 5443
rect 20151 5415 20175 5439
rect 20360 5420 20384 5444
rect 20575 5419 20595 5439
rect 22617 5414 22637 5434
rect 22828 5409 22852 5433
rect 23037 5414 23061 5438
rect 23251 5410 23277 5436
rect 25155 5411 25175 5431
rect 25366 5406 25390 5430
rect 25575 5411 25599 5435
rect 25789 5407 25815 5433
rect 29852 5425 29878 5451
rect 30068 5423 30092 5447
rect 30277 5428 30301 5452
rect 30492 5427 30512 5447
rect 30900 5421 30926 5447
rect 31116 5419 31140 5443
rect 31325 5424 31349 5448
rect 31540 5423 31560 5443
rect 33325 5408 33345 5428
rect 33536 5403 33560 5427
rect 33745 5408 33769 5432
rect 33959 5404 33985 5430
rect 35863 5405 35883 5425
rect 36074 5400 36098 5424
rect 36283 5405 36307 5429
rect 36497 5401 36523 5427
rect 40560 5419 40586 5445
rect 40776 5417 40800 5441
rect 40985 5422 41009 5446
rect 41200 5421 41220 5441
rect 41608 5415 41634 5441
rect 41824 5413 41848 5437
rect 42033 5418 42057 5442
rect 42248 5417 42268 5437
rect 945 4575 965 4595
rect 1156 4570 1180 4594
rect 1365 4575 1389 4599
rect 1579 4571 1605 4597
rect 1993 4571 2013 4591
rect 2204 4566 2228 4590
rect 2413 4571 2437 4595
rect 2627 4567 2653 4593
rect 4895 4577 4915 4597
rect 5106 4572 5130 4596
rect 5315 4577 5339 4601
rect 5529 4573 5555 4599
rect 6690 4585 6716 4611
rect 6906 4583 6930 4607
rect 7115 4588 7139 4612
rect 7330 4587 7350 4607
rect 9228 4582 9254 4608
rect 9444 4580 9468 4604
rect 9653 4585 9677 4609
rect 9868 4584 9888 4604
rect 11653 4569 11673 4589
rect 11864 4564 11888 4588
rect 12073 4569 12097 4593
rect 12287 4565 12313 4591
rect 12701 4565 12721 4585
rect 12912 4560 12936 4584
rect 13121 4565 13145 4589
rect 13335 4561 13361 4587
rect 15603 4571 15623 4591
rect 15814 4566 15838 4590
rect 16023 4571 16047 4595
rect 16237 4567 16263 4593
rect 17398 4579 17424 4605
rect 17614 4577 17638 4601
rect 17823 4582 17847 4606
rect 18038 4581 18058 4601
rect 19936 4576 19962 4602
rect 20152 4574 20176 4598
rect 20361 4579 20385 4603
rect 20576 4578 20596 4598
rect 22618 4573 22638 4593
rect 22829 4568 22853 4592
rect 23038 4573 23062 4597
rect 23252 4569 23278 4595
rect 23666 4569 23686 4589
rect 23877 4564 23901 4588
rect 24086 4569 24110 4593
rect 24300 4565 24326 4591
rect 26568 4575 26588 4595
rect 26779 4570 26803 4594
rect 26988 4575 27012 4599
rect 27202 4571 27228 4597
rect 28363 4583 28389 4609
rect 28579 4581 28603 4605
rect 28788 4586 28812 4610
rect 29003 4585 29023 4605
rect 30901 4580 30927 4606
rect 31117 4578 31141 4602
rect 31326 4583 31350 4607
rect 31541 4582 31561 4602
rect 33326 4567 33346 4587
rect 33537 4562 33561 4586
rect 33746 4567 33770 4591
rect 33960 4563 33986 4589
rect 34374 4563 34394 4583
rect 34585 4558 34609 4582
rect 34794 4563 34818 4587
rect 35008 4559 35034 4585
rect 37276 4569 37296 4589
rect 37487 4564 37511 4588
rect 37696 4569 37720 4593
rect 37910 4565 37936 4591
rect 39071 4577 39097 4603
rect 39287 4575 39311 4599
rect 39496 4580 39520 4604
rect 39711 4579 39731 4599
rect 41609 4574 41635 4600
rect 41825 4572 41849 4596
rect 42034 4577 42058 4601
rect 42249 4576 42269 4596
rect 945 3896 965 3916
rect 1156 3891 1180 3915
rect 1365 3896 1389 3920
rect 1579 3892 1605 3918
rect 3440 3891 3460 3911
rect 3651 3886 3675 3910
rect 3860 3891 3884 3915
rect 4074 3887 4100 3913
rect 8180 3907 8206 3933
rect 8396 3905 8420 3929
rect 8605 3910 8629 3934
rect 8820 3909 8840 3929
rect 9228 3903 9254 3929
rect 9444 3901 9468 3925
rect 9653 3906 9677 3930
rect 9868 3905 9888 3925
rect 11653 3890 11673 3910
rect 11864 3885 11888 3909
rect 12073 3890 12097 3914
rect 12287 3886 12313 3912
rect 14148 3885 14168 3905
rect 14359 3880 14383 3904
rect 14568 3885 14592 3909
rect 14782 3881 14808 3907
rect 18888 3901 18914 3927
rect 19104 3899 19128 3923
rect 19313 3904 19337 3928
rect 19528 3903 19548 3923
rect 19936 3897 19962 3923
rect 20152 3895 20176 3919
rect 20361 3900 20385 3924
rect 20576 3899 20596 3919
rect 22618 3894 22638 3914
rect 22829 3889 22853 3913
rect 23038 3894 23062 3918
rect 23252 3890 23278 3916
rect 25113 3889 25133 3909
rect 25324 3884 25348 3908
rect 25533 3889 25557 3913
rect 25747 3885 25773 3911
rect 29853 3905 29879 3931
rect 30069 3903 30093 3927
rect 30278 3908 30302 3932
rect 30493 3907 30513 3927
rect 30901 3901 30927 3927
rect 31117 3899 31141 3923
rect 31326 3904 31350 3928
rect 31541 3903 31561 3923
rect 33326 3888 33346 3908
rect 33537 3883 33561 3907
rect 33746 3888 33770 3912
rect 33960 3884 33986 3910
rect 35821 3883 35841 3903
rect 36032 3878 36056 3902
rect 36241 3883 36265 3907
rect 36455 3879 36481 3905
rect 40561 3899 40587 3925
rect 40777 3897 40801 3921
rect 40986 3902 41010 3926
rect 41201 3901 41221 3921
rect 41609 3895 41635 3921
rect 41825 3893 41849 3917
rect 42034 3898 42058 3922
rect 42249 3897 42269 3917
rect 945 3128 965 3148
rect 1156 3123 1180 3147
rect 1365 3128 1389 3152
rect 1579 3124 1605 3150
rect 1993 3124 2013 3144
rect 2204 3119 2228 3143
rect 2413 3124 2437 3148
rect 2627 3120 2653 3146
rect 6733 3140 6759 3166
rect 6949 3138 6973 3162
rect 7158 3143 7182 3167
rect 7373 3142 7393 3162
rect 9228 3135 9254 3161
rect 9444 3133 9468 3157
rect 9653 3138 9677 3162
rect 9868 3137 9888 3157
rect 11653 3122 11673 3142
rect 11864 3117 11888 3141
rect 12073 3122 12097 3146
rect 12287 3118 12313 3144
rect 12701 3118 12721 3138
rect 12912 3113 12936 3137
rect 13121 3118 13145 3142
rect 13335 3114 13361 3140
rect 17441 3134 17467 3160
rect 17657 3132 17681 3156
rect 17866 3137 17890 3161
rect 18081 3136 18101 3156
rect 19936 3129 19962 3155
rect 20152 3127 20176 3151
rect 20361 3132 20385 3156
rect 20576 3131 20596 3151
rect 22618 3126 22638 3146
rect 22829 3121 22853 3145
rect 23038 3126 23062 3150
rect 23252 3122 23278 3148
rect 23666 3122 23686 3142
rect 23877 3117 23901 3141
rect 24086 3122 24110 3146
rect 24300 3118 24326 3144
rect 28406 3138 28432 3164
rect 28622 3136 28646 3160
rect 28831 3141 28855 3165
rect 29046 3140 29066 3160
rect 30901 3133 30927 3159
rect 31117 3131 31141 3155
rect 31326 3136 31350 3160
rect 31541 3135 31561 3155
rect 33326 3120 33346 3140
rect 33537 3115 33561 3139
rect 33746 3120 33770 3144
rect 33960 3116 33986 3142
rect 34374 3116 34394 3136
rect 34585 3111 34609 3135
rect 34794 3116 34818 3140
rect 35008 3112 35034 3138
rect 39114 3132 39140 3158
rect 39330 3130 39354 3154
rect 39539 3135 39563 3159
rect 39754 3134 39774 3154
rect 41609 3127 41635 3153
rect 41825 3125 41849 3149
rect 42034 3130 42058 3154
rect 42249 3129 42269 3149
rect 945 2449 965 2469
rect 1156 2444 1180 2468
rect 1365 2449 1389 2473
rect 1579 2445 1605 2471
rect 8180 2460 8206 2486
rect 8396 2458 8420 2482
rect 8605 2463 8629 2487
rect 8820 2462 8840 2482
rect 9228 2456 9254 2482
rect 9444 2454 9468 2478
rect 9653 2459 9677 2483
rect 9868 2458 9888 2478
rect 11653 2443 11673 2463
rect 11864 2438 11888 2462
rect 12073 2443 12097 2467
rect 12287 2439 12313 2465
rect 18888 2454 18914 2480
rect 19104 2452 19128 2476
rect 19313 2457 19337 2481
rect 19528 2456 19548 2476
rect 19936 2450 19962 2476
rect 20152 2448 20176 2472
rect 20361 2453 20385 2477
rect 20576 2452 20596 2472
rect 22618 2447 22638 2467
rect 22829 2442 22853 2466
rect 23038 2447 23062 2471
rect 23252 2443 23278 2469
rect 29853 2458 29879 2484
rect 30069 2456 30093 2480
rect 30278 2461 30302 2485
rect 30493 2460 30513 2480
rect 30901 2454 30927 2480
rect 31117 2452 31141 2476
rect 31326 2457 31350 2481
rect 31541 2456 31561 2476
rect 33326 2441 33346 2461
rect 33537 2436 33561 2460
rect 33746 2441 33770 2465
rect 33960 2437 33986 2463
rect 40561 2452 40587 2478
rect 40777 2450 40801 2474
rect 40986 2455 41010 2479
rect 41201 2454 41221 2474
rect 41609 2448 41635 2474
rect 41825 2446 41849 2470
rect 42034 2451 42058 2475
rect 42249 2450 42269 2470
rect 10656 290 10676 310
rect 10867 285 10891 309
rect 11076 290 11100 314
rect 11290 286 11316 312
rect 21293 277 21313 297
rect 21504 272 21528 296
rect 21713 277 21737 301
rect 21927 273 21953 299
rect 32329 288 32349 308
rect 32540 283 32564 307
rect 32749 288 32773 312
rect 32963 284 32989 310
<< ndiffres >>
rect 554 13832 611 13851
rect 554 13829 575 13832
rect 460 13814 575 13829
rect 593 13814 611 13832
rect 11262 13826 11319 13845
rect 22227 13830 22284 13849
rect 22227 13827 22248 13830
rect 11262 13823 11283 13826
rect 460 13791 611 13814
rect 11168 13808 11283 13823
rect 11301 13808 11319 13826
rect 460 13755 502 13791
rect 11168 13785 11319 13808
rect 22133 13812 22248 13827
rect 22266 13812 22284 13830
rect 32935 13824 32992 13843
rect 32935 13821 32956 13824
rect 22133 13789 22284 13812
rect 32841 13806 32956 13821
rect 32974 13806 32992 13824
rect 459 13754 559 13755
rect 459 13733 615 13754
rect 459 13715 577 13733
rect 595 13715 615 13733
rect 11168 13749 11210 13785
rect 11167 13748 11267 13749
rect 459 13711 615 13715
rect 554 13695 615 13711
rect 11167 13727 11323 13748
rect 11167 13709 11285 13727
rect 11303 13709 11323 13727
rect 22133 13753 22175 13789
rect 32841 13783 32992 13806
rect 22132 13752 22232 13753
rect 11167 13705 11323 13709
rect 554 13576 611 13595
rect 554 13573 575 13576
rect 460 13558 575 13573
rect 593 13558 611 13576
rect 460 13535 611 13558
rect 460 13499 502 13535
rect 11262 13689 11323 13705
rect 10220 13645 10281 13661
rect 10220 13641 10376 13645
rect 10220 13623 10240 13641
rect 10258 13623 10376 13641
rect 459 13498 559 13499
rect 459 13477 615 13498
rect 10220 13602 10376 13623
rect 10276 13601 10376 13602
rect 10333 13565 10375 13601
rect 22132 13731 22288 13752
rect 22132 13713 22250 13731
rect 22268 13713 22288 13731
rect 32841 13747 32883 13783
rect 32840 13746 32940 13747
rect 22132 13709 22288 13713
rect 11262 13570 11319 13589
rect 11262 13567 11283 13570
rect 10224 13542 10375 13565
rect 459 13459 577 13477
rect 595 13459 615 13477
rect 459 13455 615 13459
rect 554 13439 615 13455
rect 10224 13524 10242 13542
rect 10260 13527 10375 13542
rect 11168 13552 11283 13567
rect 11301 13552 11319 13570
rect 11168 13529 11319 13552
rect 10260 13524 10281 13527
rect 10224 13505 10281 13524
rect 11168 13493 11210 13529
rect 22227 13693 22288 13709
rect 20928 13639 20989 13655
rect 20928 13635 21084 13639
rect 20928 13617 20948 13635
rect 20966 13617 21084 13635
rect 11167 13492 11267 13493
rect 11167 13471 11323 13492
rect 20928 13596 21084 13617
rect 32840 13725 32996 13746
rect 32840 13707 32958 13725
rect 32976 13707 32996 13725
rect 32840 13703 32996 13707
rect 20984 13595 21084 13596
rect 21041 13559 21083 13595
rect 22227 13574 22284 13593
rect 22227 13571 22248 13574
rect 20932 13536 21083 13559
rect 11167 13453 11285 13471
rect 11303 13453 11323 13471
rect 11167 13449 11323 13453
rect 11262 13433 11323 13449
rect 10220 13390 10281 13406
rect 10220 13386 10376 13390
rect 10220 13368 10240 13386
rect 10258 13368 10376 13386
rect 20932 13518 20950 13536
rect 20968 13521 21083 13536
rect 22133 13556 22248 13571
rect 22266 13556 22284 13574
rect 22133 13533 22284 13556
rect 20968 13518 20989 13521
rect 20932 13499 20989 13518
rect 22133 13497 22175 13533
rect 32935 13687 32996 13703
rect 31893 13643 31954 13659
rect 31893 13639 32049 13643
rect 31893 13621 31913 13639
rect 31931 13621 32049 13639
rect 22132 13496 22232 13497
rect 22132 13475 22288 13496
rect 31893 13600 32049 13621
rect 31949 13599 32049 13600
rect 32006 13563 32048 13599
rect 32935 13568 32992 13587
rect 32935 13565 32956 13568
rect 31897 13540 32048 13563
rect 22132 13457 22250 13475
rect 22268 13457 22288 13475
rect 22132 13453 22288 13457
rect 22227 13437 22288 13453
rect 10220 13347 10376 13368
rect 10276 13346 10376 13347
rect 10333 13310 10375 13346
rect 20928 13384 20989 13400
rect 20928 13380 21084 13384
rect 20928 13362 20948 13380
rect 20966 13362 21084 13380
rect 31897 13522 31915 13540
rect 31933 13525 32048 13540
rect 32841 13550 32956 13565
rect 32974 13550 32992 13568
rect 32841 13527 32992 13550
rect 31933 13522 31954 13525
rect 31897 13503 31954 13522
rect 32841 13491 32883 13527
rect 42601 13637 42662 13653
rect 42601 13633 42757 13637
rect 42601 13615 42621 13633
rect 42639 13615 42757 13633
rect 32840 13490 32940 13491
rect 32840 13469 32996 13490
rect 42601 13594 42757 13615
rect 42657 13593 42757 13594
rect 42714 13557 42756 13593
rect 42605 13534 42756 13557
rect 32840 13451 32958 13469
rect 32976 13451 32996 13469
rect 32840 13447 32996 13451
rect 32935 13431 32996 13447
rect 20928 13341 21084 13362
rect 31893 13388 31954 13404
rect 31893 13384 32049 13388
rect 31893 13366 31913 13384
rect 31931 13366 32049 13384
rect 42605 13516 42623 13534
rect 42641 13519 42756 13534
rect 42641 13516 42662 13519
rect 42605 13497 42662 13516
rect 31893 13345 32049 13366
rect 31949 13344 32049 13345
rect 20984 13340 21084 13341
rect 10224 13287 10375 13310
rect 21041 13304 21083 13340
rect 32006 13308 32048 13344
rect 42601 13382 42662 13398
rect 42601 13378 42757 13382
rect 42601 13360 42621 13378
rect 42639 13360 42757 13378
rect 42601 13339 42757 13360
rect 42657 13338 42757 13339
rect 10224 13269 10242 13287
rect 10260 13272 10375 13287
rect 20932 13281 21083 13304
rect 10260 13269 10281 13272
rect 10224 13250 10281 13269
rect 20932 13263 20950 13281
rect 20968 13266 21083 13281
rect 31897 13285 32048 13308
rect 42714 13302 42756 13338
rect 31897 13267 31915 13285
rect 31933 13270 32048 13285
rect 42605 13279 42756 13302
rect 31933 13267 31954 13270
rect 20968 13263 20989 13266
rect 20932 13244 20989 13263
rect 31897 13248 31954 13267
rect 42605 13261 42623 13279
rect 42641 13264 42756 13279
rect 42641 13261 42662 13264
rect 42605 13242 42662 13261
rect 554 13181 611 13200
rect 554 13178 575 13181
rect 460 13163 575 13178
rect 593 13163 611 13181
rect 11262 13175 11319 13194
rect 22227 13179 22284 13198
rect 22227 13176 22248 13179
rect 11262 13172 11283 13175
rect 460 13140 611 13163
rect 11168 13157 11283 13172
rect 11301 13157 11319 13175
rect 460 13104 502 13140
rect 11168 13134 11319 13157
rect 22133 13161 22248 13176
rect 22266 13161 22284 13179
rect 32935 13173 32992 13192
rect 32935 13170 32956 13173
rect 22133 13138 22284 13161
rect 32841 13155 32956 13170
rect 32974 13155 32992 13173
rect 459 13103 559 13104
rect 459 13082 615 13103
rect 459 13064 577 13082
rect 595 13064 615 13082
rect 459 13060 615 13064
rect 554 13044 615 13060
rect 11168 13098 11210 13134
rect 22133 13102 22175 13138
rect 32841 13132 32992 13155
rect 22132 13101 22232 13102
rect 11167 13097 11267 13098
rect 11167 13076 11323 13097
rect 554 12926 611 12945
rect 554 12923 575 12926
rect 460 12908 575 12923
rect 593 12908 611 12926
rect 11167 13058 11285 13076
rect 11303 13058 11323 13076
rect 11167 13054 11323 13058
rect 11262 13038 11323 13054
rect 22132 13080 22288 13101
rect 460 12885 611 12908
rect 460 12849 502 12885
rect 459 12848 559 12849
rect 459 12827 615 12848
rect 10220 12995 10281 13011
rect 10220 12991 10376 12995
rect 10220 12973 10240 12991
rect 10258 12973 10376 12991
rect 459 12809 577 12827
rect 595 12809 615 12827
rect 459 12805 615 12809
rect 554 12789 615 12805
rect 10220 12952 10376 12973
rect 10276 12951 10376 12952
rect 10333 12915 10375 12951
rect 11262 12920 11319 12939
rect 11262 12917 11283 12920
rect 10224 12892 10375 12915
rect 10224 12874 10242 12892
rect 10260 12877 10375 12892
rect 11168 12902 11283 12917
rect 11301 12902 11319 12920
rect 22132 13062 22250 13080
rect 22268 13062 22288 13080
rect 22132 13058 22288 13062
rect 22227 13042 22288 13058
rect 32841 13096 32883 13132
rect 32840 13095 32940 13096
rect 32840 13074 32996 13095
rect 11168 12879 11319 12902
rect 10260 12874 10281 12877
rect 10224 12855 10281 12874
rect 11168 12843 11210 12879
rect 11167 12842 11267 12843
rect 11167 12821 11323 12842
rect 20928 12989 20989 13005
rect 20928 12985 21084 12989
rect 20928 12967 20948 12985
rect 20966 12967 21084 12985
rect 11167 12803 11285 12821
rect 11303 12803 11323 12821
rect 11167 12799 11323 12803
rect 11262 12783 11323 12799
rect 20928 12946 21084 12967
rect 20984 12945 21084 12946
rect 10220 12739 10281 12755
rect 21041 12909 21083 12945
rect 22227 12924 22284 12943
rect 22227 12921 22248 12924
rect 20932 12886 21083 12909
rect 20932 12868 20950 12886
rect 20968 12871 21083 12886
rect 22133 12906 22248 12921
rect 22266 12906 22284 12924
rect 32840 13056 32958 13074
rect 32976 13056 32996 13074
rect 32840 13052 32996 13056
rect 32935 13036 32996 13052
rect 22133 12883 22284 12906
rect 20968 12868 20989 12871
rect 20932 12849 20989 12868
rect 22133 12847 22175 12883
rect 22132 12846 22232 12847
rect 10220 12735 10376 12739
rect 10220 12717 10240 12735
rect 10258 12717 10376 12735
rect 10220 12696 10376 12717
rect 22132 12825 22288 12846
rect 31893 12993 31954 13009
rect 31893 12989 32049 12993
rect 31893 12971 31913 12989
rect 31931 12971 32049 12989
rect 22132 12807 22250 12825
rect 22268 12807 22288 12825
rect 22132 12803 22288 12807
rect 22227 12787 22288 12803
rect 31893 12950 32049 12971
rect 31949 12949 32049 12950
rect 20928 12733 20989 12749
rect 32006 12913 32048 12949
rect 32935 12918 32992 12937
rect 32935 12915 32956 12918
rect 31897 12890 32048 12913
rect 31897 12872 31915 12890
rect 31933 12875 32048 12890
rect 32841 12900 32956 12915
rect 32974 12900 32992 12918
rect 32841 12877 32992 12900
rect 31933 12872 31954 12875
rect 31897 12853 31954 12872
rect 20928 12729 21084 12733
rect 10276 12695 10376 12696
rect 10333 12659 10375 12695
rect 20928 12711 20948 12729
rect 20966 12711 21084 12729
rect 20928 12690 21084 12711
rect 32841 12841 32883 12877
rect 32840 12840 32940 12841
rect 32840 12819 32996 12840
rect 42601 12987 42662 13003
rect 42601 12983 42757 12987
rect 42601 12965 42621 12983
rect 42639 12965 42757 12983
rect 32840 12801 32958 12819
rect 32976 12801 32996 12819
rect 32840 12797 32996 12801
rect 32935 12781 32996 12797
rect 42601 12944 42757 12965
rect 42657 12943 42757 12944
rect 31893 12737 31954 12753
rect 42714 12907 42756 12943
rect 42605 12884 42756 12907
rect 42605 12866 42623 12884
rect 42641 12869 42756 12884
rect 42641 12866 42662 12869
rect 42605 12847 42662 12866
rect 31893 12733 32049 12737
rect 20984 12689 21084 12690
rect 10224 12636 10375 12659
rect 21041 12653 21083 12689
rect 31893 12715 31913 12733
rect 31931 12715 32049 12733
rect 31893 12694 32049 12715
rect 42601 12731 42662 12747
rect 42601 12727 42757 12731
rect 31949 12693 32049 12694
rect 32006 12657 32048 12693
rect 42601 12709 42621 12727
rect 42639 12709 42757 12727
rect 42601 12688 42757 12709
rect 42657 12687 42757 12688
rect 10224 12618 10242 12636
rect 10260 12621 10375 12636
rect 20932 12630 21083 12653
rect 10260 12618 10281 12621
rect 10224 12599 10281 12618
rect 20932 12612 20950 12630
rect 20968 12615 21083 12630
rect 31897 12634 32048 12657
rect 42714 12651 42756 12687
rect 31897 12616 31915 12634
rect 31933 12619 32048 12634
rect 42605 12628 42756 12651
rect 31933 12616 31954 12619
rect 20968 12612 20989 12615
rect 20932 12593 20989 12612
rect 31897 12597 31954 12616
rect 42605 12610 42623 12628
rect 42641 12613 42756 12628
rect 42641 12610 42662 12613
rect 42605 12591 42662 12610
rect 554 12385 611 12404
rect 554 12382 575 12385
rect 460 12367 575 12382
rect 593 12367 611 12385
rect 11262 12379 11319 12398
rect 22227 12383 22284 12402
rect 22227 12380 22248 12383
rect 11262 12376 11283 12379
rect 460 12344 611 12367
rect 11168 12361 11283 12376
rect 11301 12361 11319 12379
rect 460 12308 502 12344
rect 11168 12338 11319 12361
rect 22133 12365 22248 12380
rect 22266 12365 22284 12383
rect 32935 12377 32992 12396
rect 32935 12374 32956 12377
rect 22133 12342 22284 12365
rect 32841 12359 32956 12374
rect 32974 12359 32992 12377
rect 459 12307 559 12308
rect 459 12286 615 12307
rect 459 12268 577 12286
rect 595 12268 615 12286
rect 11168 12302 11210 12338
rect 11167 12301 11267 12302
rect 459 12264 615 12268
rect 554 12248 615 12264
rect 11167 12280 11323 12301
rect 11167 12262 11285 12280
rect 11303 12262 11323 12280
rect 22133 12306 22175 12342
rect 32841 12336 32992 12359
rect 22132 12305 22232 12306
rect 11167 12258 11323 12262
rect 554 12129 611 12148
rect 554 12126 575 12129
rect 460 12111 575 12126
rect 593 12111 611 12129
rect 460 12088 611 12111
rect 460 12052 502 12088
rect 11262 12242 11323 12258
rect 459 12051 559 12052
rect 459 12030 615 12051
rect 10220 12198 10281 12214
rect 10220 12194 10376 12198
rect 10220 12176 10240 12194
rect 10258 12176 10376 12194
rect 459 12012 577 12030
rect 595 12012 615 12030
rect 459 12008 615 12012
rect 554 11992 615 12008
rect 10220 12155 10376 12176
rect 10276 12154 10376 12155
rect 10333 12118 10375 12154
rect 22132 12284 22288 12305
rect 22132 12266 22250 12284
rect 22268 12266 22288 12284
rect 32841 12300 32883 12336
rect 32840 12299 32940 12300
rect 22132 12262 22288 12266
rect 11262 12123 11319 12142
rect 11262 12120 11283 12123
rect 10224 12095 10375 12118
rect 10224 12077 10242 12095
rect 10260 12080 10375 12095
rect 11168 12105 11283 12120
rect 11301 12105 11319 12123
rect 11168 12082 11319 12105
rect 10260 12077 10281 12080
rect 10224 12058 10281 12077
rect 11168 12046 11210 12082
rect 22227 12246 22288 12262
rect 11167 12045 11267 12046
rect 11167 12024 11323 12045
rect 20928 12192 20989 12208
rect 20928 12188 21084 12192
rect 20928 12170 20948 12188
rect 20966 12170 21084 12188
rect 11167 12006 11285 12024
rect 11303 12006 11323 12024
rect 11167 12002 11323 12006
rect 11262 11986 11323 12002
rect 20928 12149 21084 12170
rect 32840 12278 32996 12299
rect 32840 12260 32958 12278
rect 32976 12260 32996 12278
rect 32840 12256 32996 12260
rect 20984 12148 21084 12149
rect 21041 12112 21083 12148
rect 22227 12127 22284 12146
rect 22227 12124 22248 12127
rect 20932 12089 21083 12112
rect 10220 11943 10281 11959
rect 10220 11939 10376 11943
rect 10220 11921 10240 11939
rect 10258 11921 10376 11939
rect 20932 12071 20950 12089
rect 20968 12074 21083 12089
rect 22133 12109 22248 12124
rect 22266 12109 22284 12127
rect 22133 12086 22284 12109
rect 20968 12071 20989 12074
rect 20932 12052 20989 12071
rect 22133 12050 22175 12086
rect 32935 12240 32996 12256
rect 22132 12049 22232 12050
rect 22132 12028 22288 12049
rect 31893 12196 31954 12212
rect 31893 12192 32049 12196
rect 31893 12174 31913 12192
rect 31931 12174 32049 12192
rect 22132 12010 22250 12028
rect 22268 12010 22288 12028
rect 22132 12006 22288 12010
rect 22227 11990 22288 12006
rect 31893 12153 32049 12174
rect 31949 12152 32049 12153
rect 32006 12116 32048 12152
rect 32935 12121 32992 12140
rect 32935 12118 32956 12121
rect 31897 12093 32048 12116
rect 10220 11900 10376 11921
rect 10276 11899 10376 11900
rect 10333 11863 10375 11899
rect 20928 11937 20989 11953
rect 20928 11933 21084 11937
rect 20928 11915 20948 11933
rect 20966 11915 21084 11933
rect 31897 12075 31915 12093
rect 31933 12078 32048 12093
rect 32841 12103 32956 12118
rect 32974 12103 32992 12121
rect 32841 12080 32992 12103
rect 31933 12075 31954 12078
rect 31897 12056 31954 12075
rect 32841 12044 32883 12080
rect 32840 12043 32940 12044
rect 32840 12022 32996 12043
rect 42601 12190 42662 12206
rect 42601 12186 42757 12190
rect 42601 12168 42621 12186
rect 42639 12168 42757 12186
rect 32840 12004 32958 12022
rect 32976 12004 32996 12022
rect 32840 12000 32996 12004
rect 32935 11984 32996 12000
rect 42601 12147 42757 12168
rect 42657 12146 42757 12147
rect 42714 12110 42756 12146
rect 42605 12087 42756 12110
rect 20928 11894 21084 11915
rect 31893 11941 31954 11957
rect 31893 11937 32049 11941
rect 31893 11919 31913 11937
rect 31931 11919 32049 11937
rect 42605 12069 42623 12087
rect 42641 12072 42756 12087
rect 42641 12069 42662 12072
rect 42605 12050 42662 12069
rect 31893 11898 32049 11919
rect 31949 11897 32049 11898
rect 20984 11893 21084 11894
rect 10224 11840 10375 11863
rect 21041 11857 21083 11893
rect 32006 11861 32048 11897
rect 42601 11935 42662 11951
rect 42601 11931 42757 11935
rect 42601 11913 42621 11931
rect 42639 11913 42757 11931
rect 42601 11892 42757 11913
rect 42657 11891 42757 11892
rect 10224 11822 10242 11840
rect 10260 11825 10375 11840
rect 20932 11834 21083 11857
rect 10260 11822 10281 11825
rect 10224 11803 10281 11822
rect 20932 11816 20950 11834
rect 20968 11819 21083 11834
rect 31897 11838 32048 11861
rect 42714 11855 42756 11891
rect 31897 11820 31915 11838
rect 31933 11823 32048 11838
rect 42605 11832 42756 11855
rect 31933 11820 31954 11823
rect 20968 11816 20989 11819
rect 20932 11797 20989 11816
rect 31897 11801 31954 11820
rect 42605 11814 42623 11832
rect 42641 11817 42756 11832
rect 42641 11814 42662 11817
rect 42605 11795 42662 11814
rect 554 11734 611 11753
rect 554 11731 575 11734
rect 460 11716 575 11731
rect 593 11716 611 11734
rect 11262 11728 11319 11747
rect 22227 11732 22284 11751
rect 22227 11729 22248 11732
rect 11262 11725 11283 11728
rect 460 11693 611 11716
rect 11168 11710 11283 11725
rect 11301 11710 11319 11728
rect 460 11657 502 11693
rect 11168 11687 11319 11710
rect 22133 11714 22248 11729
rect 22266 11714 22284 11732
rect 32935 11726 32992 11745
rect 32935 11723 32956 11726
rect 22133 11691 22284 11714
rect 32841 11708 32956 11723
rect 32974 11708 32992 11726
rect 459 11656 559 11657
rect 459 11635 615 11656
rect 459 11617 577 11635
rect 595 11617 615 11635
rect 459 11613 615 11617
rect 554 11597 615 11613
rect 11168 11651 11210 11687
rect 22133 11655 22175 11691
rect 32841 11685 32992 11708
rect 22132 11654 22232 11655
rect 11167 11650 11267 11651
rect 11167 11629 11323 11650
rect 554 11479 611 11498
rect 554 11476 575 11479
rect 460 11461 575 11476
rect 593 11461 611 11479
rect 11167 11611 11285 11629
rect 11303 11611 11323 11629
rect 11167 11607 11323 11611
rect 11262 11591 11323 11607
rect 22132 11633 22288 11654
rect 460 11438 611 11461
rect 460 11402 502 11438
rect 459 11401 559 11402
rect 459 11380 615 11401
rect 10220 11548 10281 11564
rect 10220 11544 10376 11548
rect 10220 11526 10240 11544
rect 10258 11526 10376 11544
rect 459 11362 577 11380
rect 595 11362 615 11380
rect 459 11358 615 11362
rect 554 11342 615 11358
rect 10220 11505 10376 11526
rect 10276 11504 10376 11505
rect 10333 11468 10375 11504
rect 11262 11473 11319 11492
rect 11262 11470 11283 11473
rect 10224 11445 10375 11468
rect 10224 11427 10242 11445
rect 10260 11430 10375 11445
rect 11168 11455 11283 11470
rect 11301 11455 11319 11473
rect 22132 11615 22250 11633
rect 22268 11615 22288 11633
rect 22132 11611 22288 11615
rect 22227 11595 22288 11611
rect 32841 11649 32883 11685
rect 32840 11648 32940 11649
rect 32840 11627 32996 11648
rect 11168 11432 11319 11455
rect 10260 11427 10281 11430
rect 10224 11408 10281 11427
rect 11168 11396 11210 11432
rect 11167 11395 11267 11396
rect 11167 11374 11323 11395
rect 20928 11542 20989 11558
rect 20928 11538 21084 11542
rect 20928 11520 20948 11538
rect 20966 11520 21084 11538
rect 11167 11356 11285 11374
rect 11303 11356 11323 11374
rect 11167 11352 11323 11356
rect 11262 11336 11323 11352
rect 20928 11499 21084 11520
rect 20984 11498 21084 11499
rect 10220 11292 10281 11308
rect 21041 11462 21083 11498
rect 22227 11477 22284 11496
rect 22227 11474 22248 11477
rect 20932 11439 21083 11462
rect 20932 11421 20950 11439
rect 20968 11424 21083 11439
rect 22133 11459 22248 11474
rect 22266 11459 22284 11477
rect 32840 11609 32958 11627
rect 32976 11609 32996 11627
rect 32840 11605 32996 11609
rect 32935 11589 32996 11605
rect 22133 11436 22284 11459
rect 20968 11421 20989 11424
rect 20932 11402 20989 11421
rect 22133 11400 22175 11436
rect 22132 11399 22232 11400
rect 10220 11288 10376 11292
rect 10220 11270 10240 11288
rect 10258 11270 10376 11288
rect 10220 11249 10376 11270
rect 10276 11248 10376 11249
rect 10333 11212 10375 11248
rect 22132 11378 22288 11399
rect 31893 11546 31954 11562
rect 31893 11542 32049 11546
rect 31893 11524 31913 11542
rect 31931 11524 32049 11542
rect 22132 11360 22250 11378
rect 22268 11360 22288 11378
rect 22132 11356 22288 11360
rect 22227 11340 22288 11356
rect 31893 11503 32049 11524
rect 31949 11502 32049 11503
rect 20928 11286 20989 11302
rect 32006 11466 32048 11502
rect 32935 11471 32992 11490
rect 32935 11468 32956 11471
rect 31897 11443 32048 11466
rect 31897 11425 31915 11443
rect 31933 11428 32048 11443
rect 32841 11453 32956 11468
rect 32974 11453 32992 11471
rect 32841 11430 32992 11453
rect 31933 11425 31954 11428
rect 31897 11406 31954 11425
rect 20928 11282 21084 11286
rect 20928 11264 20948 11282
rect 20966 11264 21084 11282
rect 20928 11243 21084 11264
rect 32841 11394 32883 11430
rect 32840 11393 32940 11394
rect 32840 11372 32996 11393
rect 42601 11540 42662 11556
rect 42601 11536 42757 11540
rect 42601 11518 42621 11536
rect 42639 11518 42757 11536
rect 32840 11354 32958 11372
rect 32976 11354 32996 11372
rect 32840 11350 32996 11354
rect 32935 11334 32996 11350
rect 42601 11497 42757 11518
rect 42657 11496 42757 11497
rect 31893 11290 31954 11306
rect 42714 11460 42756 11496
rect 42605 11437 42756 11460
rect 42605 11419 42623 11437
rect 42641 11422 42756 11437
rect 42641 11419 42662 11422
rect 42605 11400 42662 11419
rect 31893 11286 32049 11290
rect 20984 11242 21084 11243
rect 10224 11189 10375 11212
rect 21041 11206 21083 11242
rect 31893 11268 31913 11286
rect 31931 11268 32049 11286
rect 31893 11247 32049 11268
rect 31949 11246 32049 11247
rect 32006 11210 32048 11246
rect 42601 11284 42662 11300
rect 42601 11280 42757 11284
rect 42601 11262 42621 11280
rect 42639 11262 42757 11280
rect 42601 11241 42757 11262
rect 42657 11240 42757 11241
rect 10224 11171 10242 11189
rect 10260 11174 10375 11189
rect 20932 11183 21083 11206
rect 10260 11171 10281 11174
rect 10224 11152 10281 11171
rect 20932 11165 20950 11183
rect 20968 11168 21083 11183
rect 31897 11187 32048 11210
rect 42714 11204 42756 11240
rect 31897 11169 31915 11187
rect 31933 11172 32048 11187
rect 42605 11181 42756 11204
rect 31933 11169 31954 11172
rect 20968 11165 20989 11168
rect 20932 11146 20989 11165
rect 31897 11150 31954 11169
rect 42605 11163 42623 11181
rect 42641 11166 42756 11181
rect 42641 11163 42662 11166
rect 42605 11144 42662 11163
rect 555 10865 612 10884
rect 555 10862 576 10865
rect 461 10847 576 10862
rect 594 10847 612 10865
rect 11263 10859 11320 10878
rect 22228 10863 22285 10882
rect 22228 10860 22249 10863
rect 11263 10856 11284 10859
rect 461 10824 612 10847
rect 11169 10841 11284 10856
rect 11302 10841 11320 10859
rect 461 10788 503 10824
rect 11169 10818 11320 10841
rect 22134 10845 22249 10860
rect 22267 10845 22285 10863
rect 32936 10857 32993 10876
rect 32936 10854 32957 10857
rect 22134 10822 22285 10845
rect 32842 10839 32957 10854
rect 32975 10839 32993 10857
rect 460 10787 560 10788
rect 460 10766 616 10787
rect 460 10748 578 10766
rect 596 10748 616 10766
rect 460 10744 616 10748
rect 555 10728 616 10744
rect 11169 10782 11211 10818
rect 11168 10781 11268 10782
rect 11168 10760 11324 10781
rect 11168 10742 11286 10760
rect 11304 10742 11324 10760
rect 22134 10786 22176 10822
rect 32842 10816 32993 10839
rect 22133 10785 22233 10786
rect 11168 10738 11324 10742
rect 555 10609 612 10628
rect 555 10606 576 10609
rect 461 10591 576 10606
rect 594 10591 612 10609
rect 461 10568 612 10591
rect 461 10532 503 10568
rect 11263 10722 11324 10738
rect 460 10531 560 10532
rect 460 10510 616 10531
rect 10221 10678 10282 10694
rect 10221 10674 10377 10678
rect 10221 10656 10241 10674
rect 10259 10656 10377 10674
rect 460 10492 578 10510
rect 596 10492 616 10510
rect 460 10488 616 10492
rect 555 10472 616 10488
rect 10221 10635 10377 10656
rect 10277 10634 10377 10635
rect 10334 10598 10376 10634
rect 22133 10764 22289 10785
rect 22133 10746 22251 10764
rect 22269 10746 22289 10764
rect 22133 10742 22289 10746
rect 11263 10603 11320 10622
rect 11263 10600 11284 10603
rect 10225 10575 10376 10598
rect 10225 10557 10243 10575
rect 10261 10560 10376 10575
rect 11169 10585 11284 10600
rect 11302 10585 11320 10603
rect 11169 10562 11320 10585
rect 10261 10557 10282 10560
rect 10225 10538 10282 10557
rect 11169 10526 11211 10562
rect 22228 10726 22289 10742
rect 11168 10525 11268 10526
rect 11168 10504 11324 10525
rect 20929 10672 20990 10688
rect 20929 10668 21085 10672
rect 20929 10650 20949 10668
rect 20967 10650 21085 10668
rect 11168 10486 11286 10504
rect 11304 10486 11324 10504
rect 11168 10482 11324 10486
rect 11263 10466 11324 10482
rect 20929 10629 21085 10650
rect 32842 10780 32884 10816
rect 32841 10779 32941 10780
rect 32841 10758 32997 10779
rect 32841 10740 32959 10758
rect 32977 10740 32997 10758
rect 32841 10736 32997 10740
rect 20985 10628 21085 10629
rect 21042 10592 21084 10628
rect 22228 10607 22285 10626
rect 22228 10604 22249 10607
rect 20933 10569 21084 10592
rect 10221 10423 10282 10439
rect 10221 10419 10377 10423
rect 10221 10401 10241 10419
rect 10259 10401 10377 10419
rect 20933 10551 20951 10569
rect 20969 10554 21084 10569
rect 22134 10589 22249 10604
rect 22267 10589 22285 10607
rect 22134 10566 22285 10589
rect 20969 10551 20990 10554
rect 20933 10532 20990 10551
rect 22134 10530 22176 10566
rect 32936 10720 32997 10736
rect 22133 10529 22233 10530
rect 22133 10508 22289 10529
rect 31894 10676 31955 10692
rect 31894 10672 32050 10676
rect 31894 10654 31914 10672
rect 31932 10654 32050 10672
rect 22133 10490 22251 10508
rect 22269 10490 22289 10508
rect 22133 10486 22289 10490
rect 22228 10470 22289 10486
rect 31894 10633 32050 10654
rect 31950 10632 32050 10633
rect 32007 10596 32049 10632
rect 32936 10601 32993 10620
rect 32936 10598 32957 10601
rect 31898 10573 32049 10596
rect 10221 10380 10377 10401
rect 10277 10379 10377 10380
rect 10334 10343 10376 10379
rect 20929 10417 20990 10433
rect 20929 10413 21085 10417
rect 20929 10395 20949 10413
rect 20967 10395 21085 10413
rect 31898 10555 31916 10573
rect 31934 10558 32049 10573
rect 32842 10583 32957 10598
rect 32975 10583 32993 10601
rect 32842 10560 32993 10583
rect 31934 10555 31955 10558
rect 31898 10536 31955 10555
rect 32842 10524 32884 10560
rect 32841 10523 32941 10524
rect 32841 10502 32997 10523
rect 42602 10670 42663 10686
rect 42602 10666 42758 10670
rect 42602 10648 42622 10666
rect 42640 10648 42758 10666
rect 32841 10484 32959 10502
rect 32977 10484 32997 10502
rect 32841 10480 32997 10484
rect 32936 10464 32997 10480
rect 42602 10627 42758 10648
rect 42658 10626 42758 10627
rect 42715 10590 42757 10626
rect 42606 10567 42757 10590
rect 20929 10374 21085 10395
rect 31894 10421 31955 10437
rect 31894 10417 32050 10421
rect 31894 10399 31914 10417
rect 31932 10399 32050 10417
rect 42606 10549 42624 10567
rect 42642 10552 42757 10567
rect 42642 10549 42663 10552
rect 42606 10530 42663 10549
rect 31894 10378 32050 10399
rect 31950 10377 32050 10378
rect 20985 10373 21085 10374
rect 10225 10320 10376 10343
rect 21042 10337 21084 10373
rect 32007 10341 32049 10377
rect 42602 10415 42663 10431
rect 42602 10411 42758 10415
rect 42602 10393 42622 10411
rect 42640 10393 42758 10411
rect 42602 10372 42758 10393
rect 42658 10371 42758 10372
rect 10225 10302 10243 10320
rect 10261 10305 10376 10320
rect 20933 10314 21084 10337
rect 10261 10302 10282 10305
rect 10225 10283 10282 10302
rect 20933 10296 20951 10314
rect 20969 10299 21084 10314
rect 31898 10318 32049 10341
rect 42715 10335 42757 10371
rect 31898 10300 31916 10318
rect 31934 10303 32049 10318
rect 42606 10312 42757 10335
rect 31934 10300 31955 10303
rect 20969 10296 20990 10299
rect 20933 10277 20990 10296
rect 31898 10281 31955 10300
rect 42606 10294 42624 10312
rect 42642 10297 42757 10312
rect 42642 10294 42663 10297
rect 42606 10275 42663 10294
rect 555 10214 612 10233
rect 555 10211 576 10214
rect 461 10196 576 10211
rect 594 10196 612 10214
rect 11263 10208 11320 10227
rect 22228 10212 22285 10231
rect 22228 10209 22249 10212
rect 11263 10205 11284 10208
rect 461 10173 612 10196
rect 11169 10190 11284 10205
rect 11302 10190 11320 10208
rect 461 10137 503 10173
rect 11169 10167 11320 10190
rect 22134 10194 22249 10209
rect 22267 10194 22285 10212
rect 32936 10206 32993 10225
rect 32936 10203 32957 10206
rect 22134 10171 22285 10194
rect 32842 10188 32957 10203
rect 32975 10188 32993 10206
rect 460 10136 560 10137
rect 460 10115 616 10136
rect 460 10097 578 10115
rect 596 10097 616 10115
rect 460 10093 616 10097
rect 555 10077 616 10093
rect 11169 10131 11211 10167
rect 22134 10135 22176 10171
rect 32842 10165 32993 10188
rect 22133 10134 22233 10135
rect 11168 10130 11268 10131
rect 11168 10109 11324 10130
rect 555 9959 612 9978
rect 555 9956 576 9959
rect 461 9941 576 9956
rect 594 9941 612 9959
rect 11168 10091 11286 10109
rect 11304 10091 11324 10109
rect 11168 10087 11324 10091
rect 11263 10071 11324 10087
rect 22133 10113 22289 10134
rect 461 9918 612 9941
rect 461 9882 503 9918
rect 460 9881 560 9882
rect 460 9860 616 9881
rect 10221 10028 10282 10044
rect 10221 10024 10377 10028
rect 10221 10006 10241 10024
rect 10259 10006 10377 10024
rect 460 9842 578 9860
rect 596 9842 616 9860
rect 460 9838 616 9842
rect 555 9822 616 9838
rect 10221 9985 10377 10006
rect 10277 9984 10377 9985
rect 10334 9948 10376 9984
rect 11263 9953 11320 9972
rect 11263 9950 11284 9953
rect 10225 9925 10376 9948
rect 10225 9907 10243 9925
rect 10261 9910 10376 9925
rect 11169 9935 11284 9950
rect 11302 9935 11320 9953
rect 22133 10095 22251 10113
rect 22269 10095 22289 10113
rect 22133 10091 22289 10095
rect 22228 10075 22289 10091
rect 32842 10129 32884 10165
rect 32841 10128 32941 10129
rect 32841 10107 32997 10128
rect 11169 9912 11320 9935
rect 10261 9907 10282 9910
rect 10225 9888 10282 9907
rect 11169 9876 11211 9912
rect 11168 9875 11268 9876
rect 11168 9854 11324 9875
rect 20929 10022 20990 10038
rect 20929 10018 21085 10022
rect 20929 10000 20949 10018
rect 20967 10000 21085 10018
rect 11168 9836 11286 9854
rect 11304 9836 11324 9854
rect 11168 9832 11324 9836
rect 11263 9816 11324 9832
rect 20929 9979 21085 10000
rect 20985 9978 21085 9979
rect 10221 9772 10282 9788
rect 21042 9942 21084 9978
rect 22228 9957 22285 9976
rect 22228 9954 22249 9957
rect 20933 9919 21084 9942
rect 20933 9901 20951 9919
rect 20969 9904 21084 9919
rect 22134 9939 22249 9954
rect 22267 9939 22285 9957
rect 32841 10089 32959 10107
rect 32977 10089 32997 10107
rect 32841 10085 32997 10089
rect 32936 10069 32997 10085
rect 22134 9916 22285 9939
rect 20969 9901 20990 9904
rect 20933 9882 20990 9901
rect 22134 9880 22176 9916
rect 22133 9879 22233 9880
rect 10221 9768 10377 9772
rect 10221 9750 10241 9768
rect 10259 9750 10377 9768
rect 10221 9729 10377 9750
rect 22133 9858 22289 9879
rect 31894 10026 31955 10042
rect 31894 10022 32050 10026
rect 31894 10004 31914 10022
rect 31932 10004 32050 10022
rect 22133 9840 22251 9858
rect 22269 9840 22289 9858
rect 22133 9836 22289 9840
rect 22228 9820 22289 9836
rect 31894 9983 32050 10004
rect 31950 9982 32050 9983
rect 20929 9766 20990 9782
rect 32007 9946 32049 9982
rect 32936 9951 32993 9970
rect 32936 9948 32957 9951
rect 31898 9923 32049 9946
rect 31898 9905 31916 9923
rect 31934 9908 32049 9923
rect 32842 9933 32957 9948
rect 32975 9933 32993 9951
rect 32842 9910 32993 9933
rect 31934 9905 31955 9908
rect 31898 9886 31955 9905
rect 20929 9762 21085 9766
rect 10277 9728 10377 9729
rect 10334 9692 10376 9728
rect 20929 9744 20949 9762
rect 20967 9744 21085 9762
rect 20929 9723 21085 9744
rect 32842 9874 32884 9910
rect 32841 9873 32941 9874
rect 32841 9852 32997 9873
rect 42602 10020 42663 10036
rect 42602 10016 42758 10020
rect 42602 9998 42622 10016
rect 42640 9998 42758 10016
rect 32841 9834 32959 9852
rect 32977 9834 32997 9852
rect 32841 9830 32997 9834
rect 32936 9814 32997 9830
rect 42602 9977 42758 9998
rect 42658 9976 42758 9977
rect 31894 9770 31955 9786
rect 42715 9940 42757 9976
rect 42606 9917 42757 9940
rect 42606 9899 42624 9917
rect 42642 9902 42757 9917
rect 42642 9899 42663 9902
rect 42606 9880 42663 9899
rect 31894 9766 32050 9770
rect 20985 9722 21085 9723
rect 10225 9669 10376 9692
rect 21042 9686 21084 9722
rect 31894 9748 31914 9766
rect 31932 9748 32050 9766
rect 31894 9727 32050 9748
rect 42602 9764 42663 9780
rect 42602 9760 42758 9764
rect 31950 9726 32050 9727
rect 32007 9690 32049 9726
rect 42602 9742 42622 9760
rect 42640 9742 42758 9760
rect 42602 9721 42758 9742
rect 42658 9720 42758 9721
rect 10225 9651 10243 9669
rect 10261 9654 10376 9669
rect 20933 9663 21084 9686
rect 10261 9651 10282 9654
rect 10225 9632 10282 9651
rect 20933 9645 20951 9663
rect 20969 9648 21084 9663
rect 31898 9667 32049 9690
rect 42715 9684 42757 9720
rect 31898 9649 31916 9667
rect 31934 9652 32049 9667
rect 42606 9661 42757 9684
rect 31934 9649 31955 9652
rect 20969 9645 20990 9648
rect 20933 9626 20990 9645
rect 31898 9630 31955 9649
rect 42606 9643 42624 9661
rect 42642 9646 42757 9661
rect 42642 9643 42663 9646
rect 42606 9624 42663 9643
rect 555 9418 612 9437
rect 555 9415 576 9418
rect 461 9400 576 9415
rect 594 9400 612 9418
rect 11263 9412 11320 9431
rect 22228 9416 22285 9435
rect 22228 9413 22249 9416
rect 11263 9409 11284 9412
rect 461 9377 612 9400
rect 11169 9394 11284 9409
rect 11302 9394 11320 9412
rect 461 9341 503 9377
rect 11169 9371 11320 9394
rect 22134 9398 22249 9413
rect 22267 9398 22285 9416
rect 32936 9410 32993 9429
rect 32936 9407 32957 9410
rect 22134 9375 22285 9398
rect 32842 9392 32957 9407
rect 32975 9392 32993 9410
rect 460 9340 560 9341
rect 460 9319 616 9340
rect 460 9301 578 9319
rect 596 9301 616 9319
rect 11169 9335 11211 9371
rect 11168 9334 11268 9335
rect 460 9297 616 9301
rect 555 9281 616 9297
rect 11168 9313 11324 9334
rect 11168 9295 11286 9313
rect 11304 9295 11324 9313
rect 22134 9339 22176 9375
rect 32842 9369 32993 9392
rect 22133 9338 22233 9339
rect 11168 9291 11324 9295
rect 555 9162 612 9181
rect 555 9159 576 9162
rect 461 9144 576 9159
rect 594 9144 612 9162
rect 461 9121 612 9144
rect 461 9085 503 9121
rect 11263 9275 11324 9291
rect 460 9084 560 9085
rect 460 9063 616 9084
rect 10221 9231 10282 9247
rect 10221 9227 10377 9231
rect 10221 9209 10241 9227
rect 10259 9209 10377 9227
rect 460 9045 578 9063
rect 596 9045 616 9063
rect 460 9041 616 9045
rect 555 9025 616 9041
rect 10221 9188 10377 9209
rect 10277 9187 10377 9188
rect 10334 9151 10376 9187
rect 22133 9317 22289 9338
rect 22133 9299 22251 9317
rect 22269 9299 22289 9317
rect 32842 9333 32884 9369
rect 32841 9332 32941 9333
rect 22133 9295 22289 9299
rect 11263 9156 11320 9175
rect 11263 9153 11284 9156
rect 10225 9128 10376 9151
rect 10225 9110 10243 9128
rect 10261 9113 10376 9128
rect 11169 9138 11284 9153
rect 11302 9138 11320 9156
rect 11169 9115 11320 9138
rect 10261 9110 10282 9113
rect 10225 9091 10282 9110
rect 11169 9079 11211 9115
rect 22228 9279 22289 9295
rect 11168 9078 11268 9079
rect 11168 9057 11324 9078
rect 20929 9225 20990 9241
rect 20929 9221 21085 9225
rect 20929 9203 20949 9221
rect 20967 9203 21085 9221
rect 11168 9039 11286 9057
rect 11304 9039 11324 9057
rect 11168 9035 11324 9039
rect 11263 9019 11324 9035
rect 20929 9182 21085 9203
rect 32841 9311 32997 9332
rect 32841 9293 32959 9311
rect 32977 9293 32997 9311
rect 32841 9289 32997 9293
rect 20985 9181 21085 9182
rect 21042 9145 21084 9181
rect 22228 9160 22285 9179
rect 22228 9157 22249 9160
rect 20933 9122 21084 9145
rect 10221 8976 10282 8992
rect 10221 8972 10377 8976
rect 10221 8954 10241 8972
rect 10259 8954 10377 8972
rect 20933 9104 20951 9122
rect 20969 9107 21084 9122
rect 22134 9142 22249 9157
rect 22267 9142 22285 9160
rect 22134 9119 22285 9142
rect 20969 9104 20990 9107
rect 20933 9085 20990 9104
rect 22134 9083 22176 9119
rect 32936 9273 32997 9289
rect 22133 9082 22233 9083
rect 22133 9061 22289 9082
rect 31894 9229 31955 9245
rect 31894 9225 32050 9229
rect 31894 9207 31914 9225
rect 31932 9207 32050 9225
rect 22133 9043 22251 9061
rect 22269 9043 22289 9061
rect 22133 9039 22289 9043
rect 22228 9023 22289 9039
rect 31894 9186 32050 9207
rect 31950 9185 32050 9186
rect 32007 9149 32049 9185
rect 32936 9154 32993 9173
rect 32936 9151 32957 9154
rect 31898 9126 32049 9149
rect 10221 8933 10377 8954
rect 10277 8932 10377 8933
rect 10334 8896 10376 8932
rect 20929 8970 20990 8986
rect 20929 8966 21085 8970
rect 20929 8948 20949 8966
rect 20967 8948 21085 8966
rect 31898 9108 31916 9126
rect 31934 9111 32049 9126
rect 32842 9136 32957 9151
rect 32975 9136 32993 9154
rect 32842 9113 32993 9136
rect 31934 9108 31955 9111
rect 31898 9089 31955 9108
rect 32842 9077 32884 9113
rect 32841 9076 32941 9077
rect 32841 9055 32997 9076
rect 42602 9223 42663 9239
rect 42602 9219 42758 9223
rect 42602 9201 42622 9219
rect 42640 9201 42758 9219
rect 32841 9037 32959 9055
rect 32977 9037 32997 9055
rect 32841 9033 32997 9037
rect 32936 9017 32997 9033
rect 42602 9180 42758 9201
rect 42658 9179 42758 9180
rect 42715 9143 42757 9179
rect 42606 9120 42757 9143
rect 20929 8927 21085 8948
rect 31894 8974 31955 8990
rect 31894 8970 32050 8974
rect 31894 8952 31914 8970
rect 31932 8952 32050 8970
rect 42606 9102 42624 9120
rect 42642 9105 42757 9120
rect 42642 9102 42663 9105
rect 42606 9083 42663 9102
rect 31894 8931 32050 8952
rect 31950 8930 32050 8931
rect 20985 8926 21085 8927
rect 10225 8873 10376 8896
rect 21042 8890 21084 8926
rect 32007 8894 32049 8930
rect 42602 8968 42663 8984
rect 42602 8964 42758 8968
rect 42602 8946 42622 8964
rect 42640 8946 42758 8964
rect 42602 8925 42758 8946
rect 42658 8924 42758 8925
rect 10225 8855 10243 8873
rect 10261 8858 10376 8873
rect 20933 8867 21084 8890
rect 10261 8855 10282 8858
rect 10225 8836 10282 8855
rect 20933 8849 20951 8867
rect 20969 8852 21084 8867
rect 31898 8871 32049 8894
rect 42715 8888 42757 8924
rect 31898 8853 31916 8871
rect 31934 8856 32049 8871
rect 42606 8865 42757 8888
rect 31934 8853 31955 8856
rect 20969 8849 20990 8852
rect 20933 8830 20990 8849
rect 31898 8834 31955 8853
rect 42606 8847 42624 8865
rect 42642 8850 42757 8865
rect 42642 8847 42663 8850
rect 42606 8828 42663 8847
rect 555 8767 612 8786
rect 555 8764 576 8767
rect 461 8749 576 8764
rect 594 8749 612 8767
rect 11263 8761 11320 8780
rect 22228 8765 22285 8784
rect 22228 8762 22249 8765
rect 11263 8758 11284 8761
rect 461 8726 612 8749
rect 11169 8743 11284 8758
rect 11302 8743 11320 8761
rect 461 8690 503 8726
rect 11169 8720 11320 8743
rect 22134 8747 22249 8762
rect 22267 8747 22285 8765
rect 32936 8759 32993 8778
rect 32936 8756 32957 8759
rect 22134 8724 22285 8747
rect 32842 8741 32957 8756
rect 32975 8741 32993 8759
rect 460 8689 560 8690
rect 460 8668 616 8689
rect 460 8650 578 8668
rect 596 8650 616 8668
rect 460 8646 616 8650
rect 555 8630 616 8646
rect 11169 8684 11211 8720
rect 22134 8688 22176 8724
rect 32842 8718 32993 8741
rect 22133 8687 22233 8688
rect 11168 8683 11268 8684
rect 11168 8662 11324 8683
rect 555 8512 612 8531
rect 555 8509 576 8512
rect 461 8494 576 8509
rect 594 8494 612 8512
rect 11168 8644 11286 8662
rect 11304 8644 11324 8662
rect 11168 8640 11324 8644
rect 11263 8624 11324 8640
rect 22133 8666 22289 8687
rect 461 8471 612 8494
rect 461 8435 503 8471
rect 460 8434 560 8435
rect 460 8413 616 8434
rect 10221 8581 10282 8597
rect 10221 8577 10377 8581
rect 10221 8559 10241 8577
rect 10259 8559 10377 8577
rect 460 8395 578 8413
rect 596 8395 616 8413
rect 460 8391 616 8395
rect 555 8375 616 8391
rect 10221 8538 10377 8559
rect 10277 8537 10377 8538
rect 10334 8501 10376 8537
rect 11263 8506 11320 8525
rect 11263 8503 11284 8506
rect 10225 8478 10376 8501
rect 10225 8460 10243 8478
rect 10261 8463 10376 8478
rect 11169 8488 11284 8503
rect 11302 8488 11320 8506
rect 22133 8648 22251 8666
rect 22269 8648 22289 8666
rect 22133 8644 22289 8648
rect 22228 8628 22289 8644
rect 32842 8682 32884 8718
rect 32841 8681 32941 8682
rect 32841 8660 32997 8681
rect 11169 8465 11320 8488
rect 10261 8460 10282 8463
rect 10225 8441 10282 8460
rect 11169 8429 11211 8465
rect 11168 8428 11268 8429
rect 11168 8407 11324 8428
rect 20929 8575 20990 8591
rect 20929 8571 21085 8575
rect 20929 8553 20949 8571
rect 20967 8553 21085 8571
rect 11168 8389 11286 8407
rect 11304 8389 11324 8407
rect 11168 8385 11324 8389
rect 11263 8369 11324 8385
rect 20929 8532 21085 8553
rect 20985 8531 21085 8532
rect 10221 8325 10282 8341
rect 21042 8495 21084 8531
rect 22228 8510 22285 8529
rect 22228 8507 22249 8510
rect 20933 8472 21084 8495
rect 20933 8454 20951 8472
rect 20969 8457 21084 8472
rect 22134 8492 22249 8507
rect 22267 8492 22285 8510
rect 32841 8642 32959 8660
rect 32977 8642 32997 8660
rect 32841 8638 32997 8642
rect 32936 8622 32997 8638
rect 22134 8469 22285 8492
rect 20969 8454 20990 8457
rect 20933 8435 20990 8454
rect 22134 8433 22176 8469
rect 22133 8432 22233 8433
rect 10221 8321 10377 8325
rect 10221 8303 10241 8321
rect 10259 8303 10377 8321
rect 10221 8282 10377 8303
rect 10277 8281 10377 8282
rect 10334 8245 10376 8281
rect 22133 8411 22289 8432
rect 31894 8579 31955 8595
rect 31894 8575 32050 8579
rect 31894 8557 31914 8575
rect 31932 8557 32050 8575
rect 22133 8393 22251 8411
rect 22269 8393 22289 8411
rect 22133 8389 22289 8393
rect 22228 8373 22289 8389
rect 31894 8536 32050 8557
rect 31950 8535 32050 8536
rect 20929 8319 20990 8335
rect 32007 8499 32049 8535
rect 32936 8504 32993 8523
rect 32936 8501 32957 8504
rect 31898 8476 32049 8499
rect 31898 8458 31916 8476
rect 31934 8461 32049 8476
rect 32842 8486 32957 8501
rect 32975 8486 32993 8504
rect 32842 8463 32993 8486
rect 31934 8458 31955 8461
rect 31898 8439 31955 8458
rect 20929 8315 21085 8319
rect 20929 8297 20949 8315
rect 20967 8297 21085 8315
rect 20929 8276 21085 8297
rect 32842 8427 32884 8463
rect 32841 8426 32941 8427
rect 32841 8405 32997 8426
rect 42602 8573 42663 8589
rect 42602 8569 42758 8573
rect 42602 8551 42622 8569
rect 42640 8551 42758 8569
rect 32841 8387 32959 8405
rect 32977 8387 32997 8405
rect 32841 8383 32997 8387
rect 32936 8367 32997 8383
rect 42602 8530 42758 8551
rect 42658 8529 42758 8530
rect 31894 8323 31955 8339
rect 42715 8493 42757 8529
rect 42606 8470 42757 8493
rect 42606 8452 42624 8470
rect 42642 8455 42757 8470
rect 42642 8452 42663 8455
rect 42606 8433 42663 8452
rect 31894 8319 32050 8323
rect 20985 8275 21085 8276
rect 10225 8222 10376 8245
rect 21042 8239 21084 8275
rect 31894 8301 31914 8319
rect 31932 8301 32050 8319
rect 31894 8280 32050 8301
rect 31950 8279 32050 8280
rect 32007 8243 32049 8279
rect 42602 8317 42663 8333
rect 42602 8313 42758 8317
rect 42602 8295 42622 8313
rect 42640 8295 42758 8313
rect 42602 8274 42758 8295
rect 42658 8273 42758 8274
rect 10225 8204 10243 8222
rect 10261 8207 10376 8222
rect 20933 8216 21084 8239
rect 10261 8204 10282 8207
rect 10225 8185 10282 8204
rect 20933 8198 20951 8216
rect 20969 8201 21084 8216
rect 31898 8220 32049 8243
rect 42715 8237 42757 8273
rect 31898 8202 31916 8220
rect 31934 8205 32049 8220
rect 42606 8214 42757 8237
rect 31934 8202 31955 8205
rect 20969 8198 20990 8201
rect 20933 8179 20990 8198
rect 31898 8183 31955 8202
rect 42606 8196 42624 8214
rect 42642 8199 42757 8214
rect 42642 8196 42663 8199
rect 42606 8177 42663 8196
rect 552 7824 609 7843
rect 552 7821 573 7824
rect 458 7806 573 7821
rect 591 7806 609 7824
rect 11260 7818 11317 7837
rect 22225 7822 22282 7841
rect 22225 7819 22246 7822
rect 11260 7815 11281 7818
rect 458 7783 609 7806
rect 11166 7800 11281 7815
rect 11299 7800 11317 7818
rect 458 7747 500 7783
rect 11166 7777 11317 7800
rect 22131 7804 22246 7819
rect 22264 7804 22282 7822
rect 32933 7816 32990 7835
rect 32933 7813 32954 7816
rect 22131 7781 22282 7804
rect 32839 7798 32954 7813
rect 32972 7798 32990 7816
rect 457 7746 557 7747
rect 457 7725 613 7746
rect 457 7707 575 7725
rect 593 7707 613 7725
rect 457 7703 613 7707
rect 552 7687 613 7703
rect 11166 7741 11208 7777
rect 11165 7740 11265 7741
rect 11165 7719 11321 7740
rect 11165 7701 11283 7719
rect 11301 7701 11321 7719
rect 22131 7745 22173 7781
rect 32839 7775 32990 7798
rect 22130 7744 22230 7745
rect 11165 7697 11321 7701
rect 552 7568 609 7587
rect 552 7565 573 7568
rect 458 7550 573 7565
rect 591 7550 609 7568
rect 458 7527 609 7550
rect 458 7491 500 7527
rect 11260 7681 11321 7697
rect 457 7490 557 7491
rect 457 7469 613 7490
rect 10218 7637 10279 7653
rect 10218 7633 10374 7637
rect 10218 7615 10238 7633
rect 10256 7615 10374 7633
rect 457 7451 575 7469
rect 593 7451 613 7469
rect 457 7447 613 7451
rect 552 7431 613 7447
rect 10218 7594 10374 7615
rect 10274 7593 10374 7594
rect 10331 7557 10373 7593
rect 22130 7723 22286 7744
rect 22130 7705 22248 7723
rect 22266 7705 22286 7723
rect 22130 7701 22286 7705
rect 11260 7562 11317 7581
rect 11260 7559 11281 7562
rect 10222 7534 10373 7557
rect 10222 7516 10240 7534
rect 10258 7519 10373 7534
rect 11166 7544 11281 7559
rect 11299 7544 11317 7562
rect 11166 7521 11317 7544
rect 10258 7516 10279 7519
rect 10222 7497 10279 7516
rect 11166 7485 11208 7521
rect 22225 7685 22286 7701
rect 11165 7484 11265 7485
rect 11165 7463 11321 7484
rect 20926 7631 20987 7647
rect 20926 7627 21082 7631
rect 20926 7609 20946 7627
rect 20964 7609 21082 7627
rect 11165 7445 11283 7463
rect 11301 7445 11321 7463
rect 11165 7441 11321 7445
rect 11260 7425 11321 7441
rect 20926 7588 21082 7609
rect 32839 7739 32881 7775
rect 32838 7738 32938 7739
rect 32838 7717 32994 7738
rect 32838 7699 32956 7717
rect 32974 7699 32994 7717
rect 32838 7695 32994 7699
rect 20982 7587 21082 7588
rect 21039 7551 21081 7587
rect 22225 7566 22282 7585
rect 22225 7563 22246 7566
rect 20930 7528 21081 7551
rect 10218 7382 10279 7398
rect 10218 7378 10374 7382
rect 10218 7360 10238 7378
rect 10256 7360 10374 7378
rect 20930 7510 20948 7528
rect 20966 7513 21081 7528
rect 22131 7548 22246 7563
rect 22264 7548 22282 7566
rect 22131 7525 22282 7548
rect 20966 7510 20987 7513
rect 20930 7491 20987 7510
rect 22131 7489 22173 7525
rect 32933 7679 32994 7695
rect 22130 7488 22230 7489
rect 22130 7467 22286 7488
rect 31891 7635 31952 7651
rect 31891 7631 32047 7635
rect 31891 7613 31911 7631
rect 31929 7613 32047 7631
rect 22130 7449 22248 7467
rect 22266 7449 22286 7467
rect 22130 7445 22286 7449
rect 22225 7429 22286 7445
rect 31891 7592 32047 7613
rect 31947 7591 32047 7592
rect 32004 7555 32046 7591
rect 32933 7560 32990 7579
rect 32933 7557 32954 7560
rect 31895 7532 32046 7555
rect 10218 7339 10374 7360
rect 10274 7338 10374 7339
rect 10331 7302 10373 7338
rect 20926 7376 20987 7392
rect 20926 7372 21082 7376
rect 20926 7354 20946 7372
rect 20964 7354 21082 7372
rect 31895 7514 31913 7532
rect 31931 7517 32046 7532
rect 32839 7542 32954 7557
rect 32972 7542 32990 7560
rect 32839 7519 32990 7542
rect 31931 7514 31952 7517
rect 31895 7495 31952 7514
rect 32839 7483 32881 7519
rect 32838 7482 32938 7483
rect 32838 7461 32994 7482
rect 42599 7629 42660 7645
rect 42599 7625 42755 7629
rect 42599 7607 42619 7625
rect 42637 7607 42755 7625
rect 32838 7443 32956 7461
rect 32974 7443 32994 7461
rect 32838 7439 32994 7443
rect 32933 7423 32994 7439
rect 42599 7586 42755 7607
rect 42655 7585 42755 7586
rect 42712 7549 42754 7585
rect 42603 7526 42754 7549
rect 20926 7333 21082 7354
rect 31891 7380 31952 7396
rect 31891 7376 32047 7380
rect 31891 7358 31911 7376
rect 31929 7358 32047 7376
rect 42603 7508 42621 7526
rect 42639 7511 42754 7526
rect 42639 7508 42660 7511
rect 42603 7489 42660 7508
rect 31891 7337 32047 7358
rect 31947 7336 32047 7337
rect 20982 7332 21082 7333
rect 10222 7279 10373 7302
rect 21039 7296 21081 7332
rect 32004 7300 32046 7336
rect 42599 7374 42660 7390
rect 42599 7370 42755 7374
rect 42599 7352 42619 7370
rect 42637 7352 42755 7370
rect 42599 7331 42755 7352
rect 42655 7330 42755 7331
rect 10222 7261 10240 7279
rect 10258 7264 10373 7279
rect 20930 7273 21081 7296
rect 10258 7261 10279 7264
rect 10222 7242 10279 7261
rect 20930 7255 20948 7273
rect 20966 7258 21081 7273
rect 31895 7277 32046 7300
rect 42712 7294 42754 7330
rect 31895 7259 31913 7277
rect 31931 7262 32046 7277
rect 42603 7271 42754 7294
rect 31931 7259 31952 7262
rect 20966 7255 20987 7258
rect 20930 7236 20987 7255
rect 31895 7240 31952 7259
rect 42603 7253 42621 7271
rect 42639 7256 42754 7271
rect 42639 7253 42660 7256
rect 42603 7234 42660 7253
rect 552 7173 609 7192
rect 552 7170 573 7173
rect 458 7155 573 7170
rect 591 7155 609 7173
rect 11260 7167 11317 7186
rect 22225 7171 22282 7190
rect 22225 7168 22246 7171
rect 11260 7164 11281 7167
rect 458 7132 609 7155
rect 11166 7149 11281 7164
rect 11299 7149 11317 7167
rect 458 7096 500 7132
rect 11166 7126 11317 7149
rect 22131 7153 22246 7168
rect 22264 7153 22282 7171
rect 32933 7165 32990 7184
rect 32933 7162 32954 7165
rect 22131 7130 22282 7153
rect 32839 7147 32954 7162
rect 32972 7147 32990 7165
rect 457 7095 557 7096
rect 457 7074 613 7095
rect 457 7056 575 7074
rect 593 7056 613 7074
rect 457 7052 613 7056
rect 552 7036 613 7052
rect 11166 7090 11208 7126
rect 22131 7094 22173 7130
rect 32839 7124 32990 7147
rect 22130 7093 22230 7094
rect 11165 7089 11265 7090
rect 11165 7068 11321 7089
rect 552 6918 609 6937
rect 552 6915 573 6918
rect 458 6900 573 6915
rect 591 6900 609 6918
rect 11165 7050 11283 7068
rect 11301 7050 11321 7068
rect 11165 7046 11321 7050
rect 11260 7030 11321 7046
rect 22130 7072 22286 7093
rect 458 6877 609 6900
rect 458 6841 500 6877
rect 457 6840 557 6841
rect 457 6819 613 6840
rect 10218 6987 10279 7003
rect 10218 6983 10374 6987
rect 10218 6965 10238 6983
rect 10256 6965 10374 6983
rect 457 6801 575 6819
rect 593 6801 613 6819
rect 457 6797 613 6801
rect 552 6781 613 6797
rect 10218 6944 10374 6965
rect 10274 6943 10374 6944
rect 10331 6907 10373 6943
rect 11260 6912 11317 6931
rect 11260 6909 11281 6912
rect 10222 6884 10373 6907
rect 10222 6866 10240 6884
rect 10258 6869 10373 6884
rect 11166 6894 11281 6909
rect 11299 6894 11317 6912
rect 22130 7054 22248 7072
rect 22266 7054 22286 7072
rect 22130 7050 22286 7054
rect 22225 7034 22286 7050
rect 32839 7088 32881 7124
rect 32838 7087 32938 7088
rect 32838 7066 32994 7087
rect 11166 6871 11317 6894
rect 10258 6866 10279 6869
rect 10222 6847 10279 6866
rect 11166 6835 11208 6871
rect 11165 6834 11265 6835
rect 11165 6813 11321 6834
rect 20926 6981 20987 6997
rect 20926 6977 21082 6981
rect 20926 6959 20946 6977
rect 20964 6959 21082 6977
rect 11165 6795 11283 6813
rect 11301 6795 11321 6813
rect 11165 6791 11321 6795
rect 11260 6775 11321 6791
rect 20926 6938 21082 6959
rect 20982 6937 21082 6938
rect 10218 6731 10279 6747
rect 21039 6901 21081 6937
rect 22225 6916 22282 6935
rect 22225 6913 22246 6916
rect 20930 6878 21081 6901
rect 20930 6860 20948 6878
rect 20966 6863 21081 6878
rect 22131 6898 22246 6913
rect 22264 6898 22282 6916
rect 32838 7048 32956 7066
rect 32974 7048 32994 7066
rect 32838 7044 32994 7048
rect 32933 7028 32994 7044
rect 22131 6875 22282 6898
rect 20966 6860 20987 6863
rect 20930 6841 20987 6860
rect 22131 6839 22173 6875
rect 22130 6838 22230 6839
rect 10218 6727 10374 6731
rect 10218 6709 10238 6727
rect 10256 6709 10374 6727
rect 10218 6688 10374 6709
rect 22130 6817 22286 6838
rect 31891 6985 31952 7001
rect 31891 6981 32047 6985
rect 31891 6963 31911 6981
rect 31929 6963 32047 6981
rect 22130 6799 22248 6817
rect 22266 6799 22286 6817
rect 22130 6795 22286 6799
rect 22225 6779 22286 6795
rect 31891 6942 32047 6963
rect 31947 6941 32047 6942
rect 20926 6725 20987 6741
rect 32004 6905 32046 6941
rect 32933 6910 32990 6929
rect 32933 6907 32954 6910
rect 31895 6882 32046 6905
rect 31895 6864 31913 6882
rect 31931 6867 32046 6882
rect 32839 6892 32954 6907
rect 32972 6892 32990 6910
rect 32839 6869 32990 6892
rect 31931 6864 31952 6867
rect 31895 6845 31952 6864
rect 20926 6721 21082 6725
rect 10274 6687 10374 6688
rect 10331 6651 10373 6687
rect 20926 6703 20946 6721
rect 20964 6703 21082 6721
rect 20926 6682 21082 6703
rect 32839 6833 32881 6869
rect 32838 6832 32938 6833
rect 32838 6811 32994 6832
rect 42599 6979 42660 6995
rect 42599 6975 42755 6979
rect 42599 6957 42619 6975
rect 42637 6957 42755 6975
rect 32838 6793 32956 6811
rect 32974 6793 32994 6811
rect 32838 6789 32994 6793
rect 32933 6773 32994 6789
rect 42599 6936 42755 6957
rect 42655 6935 42755 6936
rect 31891 6729 31952 6745
rect 42712 6899 42754 6935
rect 42603 6876 42754 6899
rect 42603 6858 42621 6876
rect 42639 6861 42754 6876
rect 42639 6858 42660 6861
rect 42603 6839 42660 6858
rect 31891 6725 32047 6729
rect 20982 6681 21082 6682
rect 10222 6628 10373 6651
rect 21039 6645 21081 6681
rect 31891 6707 31911 6725
rect 31929 6707 32047 6725
rect 31891 6686 32047 6707
rect 42599 6723 42660 6739
rect 42599 6719 42755 6723
rect 31947 6685 32047 6686
rect 32004 6649 32046 6685
rect 42599 6701 42619 6719
rect 42637 6701 42755 6719
rect 42599 6680 42755 6701
rect 42655 6679 42755 6680
rect 10222 6610 10240 6628
rect 10258 6613 10373 6628
rect 20930 6622 21081 6645
rect 10258 6610 10279 6613
rect 10222 6591 10279 6610
rect 20930 6604 20948 6622
rect 20966 6607 21081 6622
rect 31895 6626 32046 6649
rect 42712 6643 42754 6679
rect 31895 6608 31913 6626
rect 31931 6611 32046 6626
rect 42603 6620 42754 6643
rect 31931 6608 31952 6611
rect 20966 6604 20987 6607
rect 20930 6585 20987 6604
rect 31895 6589 31952 6608
rect 42603 6602 42621 6620
rect 42639 6605 42754 6620
rect 42639 6602 42660 6605
rect 42603 6583 42660 6602
rect 552 6377 609 6396
rect 552 6374 573 6377
rect 458 6359 573 6374
rect 591 6359 609 6377
rect 11260 6371 11317 6390
rect 22225 6375 22282 6394
rect 22225 6372 22246 6375
rect 11260 6368 11281 6371
rect 458 6336 609 6359
rect 11166 6353 11281 6368
rect 11299 6353 11317 6371
rect 458 6300 500 6336
rect 11166 6330 11317 6353
rect 22131 6357 22246 6372
rect 22264 6357 22282 6375
rect 32933 6369 32990 6388
rect 32933 6366 32954 6369
rect 22131 6334 22282 6357
rect 32839 6351 32954 6366
rect 32972 6351 32990 6369
rect 457 6299 557 6300
rect 457 6278 613 6299
rect 457 6260 575 6278
rect 593 6260 613 6278
rect 11166 6294 11208 6330
rect 11165 6293 11265 6294
rect 457 6256 613 6260
rect 552 6240 613 6256
rect 11165 6272 11321 6293
rect 11165 6254 11283 6272
rect 11301 6254 11321 6272
rect 22131 6298 22173 6334
rect 32839 6328 32990 6351
rect 22130 6297 22230 6298
rect 11165 6250 11321 6254
rect 552 6121 609 6140
rect 552 6118 573 6121
rect 458 6103 573 6118
rect 591 6103 609 6121
rect 458 6080 609 6103
rect 458 6044 500 6080
rect 11260 6234 11321 6250
rect 457 6043 557 6044
rect 457 6022 613 6043
rect 10218 6190 10279 6206
rect 10218 6186 10374 6190
rect 10218 6168 10238 6186
rect 10256 6168 10374 6186
rect 457 6004 575 6022
rect 593 6004 613 6022
rect 457 6000 613 6004
rect 552 5984 613 6000
rect 10218 6147 10374 6168
rect 10274 6146 10374 6147
rect 10331 6110 10373 6146
rect 22130 6276 22286 6297
rect 22130 6258 22248 6276
rect 22266 6258 22286 6276
rect 32839 6292 32881 6328
rect 32838 6291 32938 6292
rect 22130 6254 22286 6258
rect 11260 6115 11317 6134
rect 11260 6112 11281 6115
rect 10222 6087 10373 6110
rect 10222 6069 10240 6087
rect 10258 6072 10373 6087
rect 11166 6097 11281 6112
rect 11299 6097 11317 6115
rect 11166 6074 11317 6097
rect 10258 6069 10279 6072
rect 10222 6050 10279 6069
rect 11166 6038 11208 6074
rect 22225 6238 22286 6254
rect 11165 6037 11265 6038
rect 11165 6016 11321 6037
rect 20926 6184 20987 6200
rect 20926 6180 21082 6184
rect 20926 6162 20946 6180
rect 20964 6162 21082 6180
rect 11165 5998 11283 6016
rect 11301 5998 11321 6016
rect 11165 5994 11321 5998
rect 11260 5978 11321 5994
rect 20926 6141 21082 6162
rect 32838 6270 32994 6291
rect 32838 6252 32956 6270
rect 32974 6252 32994 6270
rect 32838 6248 32994 6252
rect 20982 6140 21082 6141
rect 21039 6104 21081 6140
rect 22225 6119 22282 6138
rect 22225 6116 22246 6119
rect 20930 6081 21081 6104
rect 10218 5935 10279 5951
rect 10218 5931 10374 5935
rect 10218 5913 10238 5931
rect 10256 5913 10374 5931
rect 20930 6063 20948 6081
rect 20966 6066 21081 6081
rect 22131 6101 22246 6116
rect 22264 6101 22282 6119
rect 22131 6078 22282 6101
rect 20966 6063 20987 6066
rect 20930 6044 20987 6063
rect 22131 6042 22173 6078
rect 32933 6232 32994 6248
rect 22130 6041 22230 6042
rect 22130 6020 22286 6041
rect 31891 6188 31952 6204
rect 31891 6184 32047 6188
rect 31891 6166 31911 6184
rect 31929 6166 32047 6184
rect 22130 6002 22248 6020
rect 22266 6002 22286 6020
rect 22130 5998 22286 6002
rect 22225 5982 22286 5998
rect 31891 6145 32047 6166
rect 31947 6144 32047 6145
rect 32004 6108 32046 6144
rect 32933 6113 32990 6132
rect 32933 6110 32954 6113
rect 31895 6085 32046 6108
rect 10218 5892 10374 5913
rect 10274 5891 10374 5892
rect 10331 5855 10373 5891
rect 20926 5929 20987 5945
rect 20926 5925 21082 5929
rect 20926 5907 20946 5925
rect 20964 5907 21082 5925
rect 31895 6067 31913 6085
rect 31931 6070 32046 6085
rect 32839 6095 32954 6110
rect 32972 6095 32990 6113
rect 32839 6072 32990 6095
rect 31931 6067 31952 6070
rect 31895 6048 31952 6067
rect 32839 6036 32881 6072
rect 32838 6035 32938 6036
rect 32838 6014 32994 6035
rect 42599 6182 42660 6198
rect 42599 6178 42755 6182
rect 42599 6160 42619 6178
rect 42637 6160 42755 6178
rect 32838 5996 32956 6014
rect 32974 5996 32994 6014
rect 32838 5992 32994 5996
rect 32933 5976 32994 5992
rect 42599 6139 42755 6160
rect 42655 6138 42755 6139
rect 42712 6102 42754 6138
rect 42603 6079 42754 6102
rect 20926 5886 21082 5907
rect 31891 5933 31952 5949
rect 31891 5929 32047 5933
rect 31891 5911 31911 5929
rect 31929 5911 32047 5929
rect 42603 6061 42621 6079
rect 42639 6064 42754 6079
rect 42639 6061 42660 6064
rect 42603 6042 42660 6061
rect 31891 5890 32047 5911
rect 31947 5889 32047 5890
rect 20982 5885 21082 5886
rect 10222 5832 10373 5855
rect 21039 5849 21081 5885
rect 32004 5853 32046 5889
rect 42599 5927 42660 5943
rect 42599 5923 42755 5927
rect 42599 5905 42619 5923
rect 42637 5905 42755 5923
rect 42599 5884 42755 5905
rect 42655 5883 42755 5884
rect 10222 5814 10240 5832
rect 10258 5817 10373 5832
rect 20930 5826 21081 5849
rect 10258 5814 10279 5817
rect 10222 5795 10279 5814
rect 20930 5808 20948 5826
rect 20966 5811 21081 5826
rect 31895 5830 32046 5853
rect 42712 5847 42754 5883
rect 31895 5812 31913 5830
rect 31931 5815 32046 5830
rect 42603 5824 42754 5847
rect 31931 5812 31952 5815
rect 20966 5808 20987 5811
rect 20930 5789 20987 5808
rect 31895 5793 31952 5812
rect 42603 5806 42621 5824
rect 42639 5809 42754 5824
rect 42639 5806 42660 5809
rect 42603 5787 42660 5806
rect 552 5726 609 5745
rect 552 5723 573 5726
rect 458 5708 573 5723
rect 591 5708 609 5726
rect 11260 5720 11317 5739
rect 22225 5724 22282 5743
rect 22225 5721 22246 5724
rect 11260 5717 11281 5720
rect 458 5685 609 5708
rect 11166 5702 11281 5717
rect 11299 5702 11317 5720
rect 458 5649 500 5685
rect 11166 5679 11317 5702
rect 22131 5706 22246 5721
rect 22264 5706 22282 5724
rect 32933 5718 32990 5737
rect 32933 5715 32954 5718
rect 22131 5683 22282 5706
rect 32839 5700 32954 5715
rect 32972 5700 32990 5718
rect 457 5648 557 5649
rect 457 5627 613 5648
rect 457 5609 575 5627
rect 593 5609 613 5627
rect 457 5605 613 5609
rect 552 5589 613 5605
rect 11166 5643 11208 5679
rect 22131 5647 22173 5683
rect 32839 5677 32990 5700
rect 22130 5646 22230 5647
rect 11165 5642 11265 5643
rect 11165 5621 11321 5642
rect 552 5471 609 5490
rect 552 5468 573 5471
rect 458 5453 573 5468
rect 591 5453 609 5471
rect 11165 5603 11283 5621
rect 11301 5603 11321 5621
rect 11165 5599 11321 5603
rect 11260 5583 11321 5599
rect 22130 5625 22286 5646
rect 458 5430 609 5453
rect 458 5394 500 5430
rect 457 5393 557 5394
rect 457 5372 613 5393
rect 10218 5540 10279 5556
rect 10218 5536 10374 5540
rect 10218 5518 10238 5536
rect 10256 5518 10374 5536
rect 457 5354 575 5372
rect 593 5354 613 5372
rect 457 5350 613 5354
rect 552 5334 613 5350
rect 10218 5497 10374 5518
rect 10274 5496 10374 5497
rect 10331 5460 10373 5496
rect 11260 5465 11317 5484
rect 11260 5462 11281 5465
rect 10222 5437 10373 5460
rect 10222 5419 10240 5437
rect 10258 5422 10373 5437
rect 11166 5447 11281 5462
rect 11299 5447 11317 5465
rect 22130 5607 22248 5625
rect 22266 5607 22286 5625
rect 22130 5603 22286 5607
rect 22225 5587 22286 5603
rect 32839 5641 32881 5677
rect 32838 5640 32938 5641
rect 32838 5619 32994 5640
rect 11166 5424 11317 5447
rect 10258 5419 10279 5422
rect 10222 5400 10279 5419
rect 11166 5388 11208 5424
rect 11165 5387 11265 5388
rect 11165 5366 11321 5387
rect 20926 5534 20987 5550
rect 20926 5530 21082 5534
rect 20926 5512 20946 5530
rect 20964 5512 21082 5530
rect 11165 5348 11283 5366
rect 11301 5348 11321 5366
rect 11165 5344 11321 5348
rect 11260 5328 11321 5344
rect 20926 5491 21082 5512
rect 20982 5490 21082 5491
rect 10218 5284 10279 5300
rect 21039 5454 21081 5490
rect 22225 5469 22282 5488
rect 22225 5466 22246 5469
rect 20930 5431 21081 5454
rect 20930 5413 20948 5431
rect 20966 5416 21081 5431
rect 22131 5451 22246 5466
rect 22264 5451 22282 5469
rect 32838 5601 32956 5619
rect 32974 5601 32994 5619
rect 32838 5597 32994 5601
rect 32933 5581 32994 5597
rect 22131 5428 22282 5451
rect 20966 5413 20987 5416
rect 20930 5394 20987 5413
rect 22131 5392 22173 5428
rect 22130 5391 22230 5392
rect 10218 5280 10374 5284
rect 10218 5262 10238 5280
rect 10256 5262 10374 5280
rect 10218 5241 10374 5262
rect 10274 5240 10374 5241
rect 10331 5204 10373 5240
rect 22130 5370 22286 5391
rect 31891 5538 31952 5554
rect 31891 5534 32047 5538
rect 31891 5516 31911 5534
rect 31929 5516 32047 5534
rect 22130 5352 22248 5370
rect 22266 5352 22286 5370
rect 22130 5348 22286 5352
rect 22225 5332 22286 5348
rect 31891 5495 32047 5516
rect 31947 5494 32047 5495
rect 20926 5278 20987 5294
rect 32004 5458 32046 5494
rect 32933 5463 32990 5482
rect 32933 5460 32954 5463
rect 31895 5435 32046 5458
rect 31895 5417 31913 5435
rect 31931 5420 32046 5435
rect 32839 5445 32954 5460
rect 32972 5445 32990 5463
rect 32839 5422 32990 5445
rect 31931 5417 31952 5420
rect 31895 5398 31952 5417
rect 20926 5274 21082 5278
rect 20926 5256 20946 5274
rect 20964 5256 21082 5274
rect 20926 5235 21082 5256
rect 32839 5386 32881 5422
rect 32838 5385 32938 5386
rect 32838 5364 32994 5385
rect 42599 5532 42660 5548
rect 42599 5528 42755 5532
rect 42599 5510 42619 5528
rect 42637 5510 42755 5528
rect 32838 5346 32956 5364
rect 32974 5346 32994 5364
rect 32838 5342 32994 5346
rect 32933 5326 32994 5342
rect 42599 5489 42755 5510
rect 42655 5488 42755 5489
rect 31891 5282 31952 5298
rect 42712 5452 42754 5488
rect 42603 5429 42754 5452
rect 42603 5411 42621 5429
rect 42639 5414 42754 5429
rect 42639 5411 42660 5414
rect 42603 5392 42660 5411
rect 31891 5278 32047 5282
rect 20982 5234 21082 5235
rect 10222 5181 10373 5204
rect 21039 5198 21081 5234
rect 31891 5260 31911 5278
rect 31929 5260 32047 5278
rect 31891 5239 32047 5260
rect 31947 5238 32047 5239
rect 32004 5202 32046 5238
rect 42599 5276 42660 5292
rect 42599 5272 42755 5276
rect 42599 5254 42619 5272
rect 42637 5254 42755 5272
rect 42599 5233 42755 5254
rect 42655 5232 42755 5233
rect 10222 5163 10240 5181
rect 10258 5166 10373 5181
rect 20930 5175 21081 5198
rect 10258 5163 10279 5166
rect 10222 5144 10279 5163
rect 20930 5157 20948 5175
rect 20966 5160 21081 5175
rect 31895 5179 32046 5202
rect 42712 5196 42754 5232
rect 31895 5161 31913 5179
rect 31931 5164 32046 5179
rect 42603 5173 42754 5196
rect 31931 5161 31952 5164
rect 20966 5157 20987 5160
rect 20930 5138 20987 5157
rect 31895 5142 31952 5161
rect 42603 5155 42621 5173
rect 42639 5158 42754 5173
rect 42639 5155 42660 5158
rect 42603 5136 42660 5155
rect 553 4857 610 4876
rect 553 4854 574 4857
rect 459 4839 574 4854
rect 592 4839 610 4857
rect 11261 4851 11318 4870
rect 22226 4855 22283 4874
rect 22226 4852 22247 4855
rect 11261 4848 11282 4851
rect 459 4816 610 4839
rect 11167 4833 11282 4848
rect 11300 4833 11318 4851
rect 459 4780 501 4816
rect 458 4779 558 4780
rect 458 4758 614 4779
rect 458 4740 576 4758
rect 594 4740 614 4758
rect 11167 4810 11318 4833
rect 22132 4837 22247 4852
rect 22265 4837 22283 4855
rect 32934 4849 32991 4868
rect 32934 4846 32955 4849
rect 22132 4814 22283 4837
rect 32840 4831 32955 4846
rect 32973 4831 32991 4849
rect 458 4736 614 4740
rect 553 4720 614 4736
rect 553 4601 610 4620
rect 553 4598 574 4601
rect 459 4583 574 4598
rect 592 4583 610 4601
rect 459 4560 610 4583
rect 459 4524 501 4560
rect 11167 4774 11209 4810
rect 11166 4773 11266 4774
rect 11166 4752 11322 4773
rect 11166 4734 11284 4752
rect 11302 4734 11322 4752
rect 22132 4778 22174 4814
rect 22131 4777 22231 4778
rect 11166 4730 11322 4734
rect 11261 4714 11322 4730
rect 458 4523 558 4524
rect 458 4502 614 4523
rect 10219 4670 10280 4686
rect 10219 4666 10375 4670
rect 10219 4648 10239 4666
rect 10257 4648 10375 4666
rect 458 4484 576 4502
rect 594 4484 614 4502
rect 458 4480 614 4484
rect 553 4464 614 4480
rect 10219 4627 10375 4648
rect 10275 4626 10375 4627
rect 10332 4590 10374 4626
rect 11261 4595 11318 4614
rect 11261 4592 11282 4595
rect 10223 4567 10374 4590
rect 10223 4549 10241 4567
rect 10259 4552 10374 4567
rect 11167 4577 11282 4592
rect 11300 4577 11318 4595
rect 11167 4554 11318 4577
rect 10259 4549 10280 4552
rect 10223 4530 10280 4549
rect 11167 4518 11209 4554
rect 22131 4756 22287 4777
rect 22131 4738 22249 4756
rect 22267 4738 22287 4756
rect 32840 4808 32991 4831
rect 22131 4734 22287 4738
rect 22226 4718 22287 4734
rect 11166 4517 11266 4518
rect 11166 4496 11322 4517
rect 20927 4664 20988 4680
rect 20927 4660 21083 4664
rect 20927 4642 20947 4660
rect 20965 4642 21083 4660
rect 11166 4478 11284 4496
rect 11302 4478 11322 4496
rect 11166 4474 11322 4478
rect 11261 4458 11322 4474
rect 10219 4415 10280 4431
rect 10219 4411 10375 4415
rect 10219 4393 10239 4411
rect 10257 4393 10375 4411
rect 20927 4621 21083 4642
rect 20983 4620 21083 4621
rect 21040 4584 21082 4620
rect 22226 4599 22283 4618
rect 22226 4596 22247 4599
rect 20931 4561 21082 4584
rect 20931 4543 20949 4561
rect 20967 4546 21082 4561
rect 22132 4581 22247 4596
rect 22265 4581 22283 4599
rect 22132 4558 22283 4581
rect 20967 4543 20988 4546
rect 20931 4524 20988 4543
rect 22132 4522 22174 4558
rect 32840 4772 32882 4808
rect 32839 4771 32939 4772
rect 32839 4750 32995 4771
rect 32839 4732 32957 4750
rect 32975 4732 32995 4750
rect 32839 4728 32995 4732
rect 32934 4712 32995 4728
rect 22131 4521 22231 4522
rect 22131 4500 22287 4521
rect 31892 4668 31953 4684
rect 31892 4664 32048 4668
rect 31892 4646 31912 4664
rect 31930 4646 32048 4664
rect 22131 4482 22249 4500
rect 22267 4482 22287 4500
rect 22131 4478 22287 4482
rect 22226 4462 22287 4478
rect 10219 4372 10375 4393
rect 10275 4371 10375 4372
rect 10332 4335 10374 4371
rect 20927 4409 20988 4425
rect 20927 4405 21083 4409
rect 20927 4387 20947 4405
rect 20965 4387 21083 4405
rect 31892 4625 32048 4646
rect 31948 4624 32048 4625
rect 32005 4588 32047 4624
rect 32934 4593 32991 4612
rect 32934 4590 32955 4593
rect 31896 4565 32047 4588
rect 31896 4547 31914 4565
rect 31932 4550 32047 4565
rect 32840 4575 32955 4590
rect 32973 4575 32991 4593
rect 32840 4552 32991 4575
rect 31932 4547 31953 4550
rect 31896 4528 31953 4547
rect 32840 4516 32882 4552
rect 32839 4515 32939 4516
rect 32839 4494 32995 4515
rect 42600 4662 42661 4678
rect 42600 4658 42756 4662
rect 42600 4640 42620 4658
rect 42638 4640 42756 4658
rect 32839 4476 32957 4494
rect 32975 4476 32995 4494
rect 32839 4472 32995 4476
rect 32934 4456 32995 4472
rect 20927 4366 21083 4387
rect 31892 4413 31953 4429
rect 31892 4409 32048 4413
rect 31892 4391 31912 4409
rect 31930 4391 32048 4409
rect 42600 4619 42756 4640
rect 42656 4618 42756 4619
rect 42713 4582 42755 4618
rect 42604 4559 42755 4582
rect 42604 4541 42622 4559
rect 42640 4544 42755 4559
rect 42640 4541 42661 4544
rect 42604 4522 42661 4541
rect 31892 4370 32048 4391
rect 31948 4369 32048 4370
rect 20983 4365 21083 4366
rect 10223 4312 10374 4335
rect 21040 4329 21082 4365
rect 32005 4333 32047 4369
rect 42600 4407 42661 4423
rect 42600 4403 42756 4407
rect 42600 4385 42620 4403
rect 42638 4385 42756 4403
rect 42600 4364 42756 4385
rect 42656 4363 42756 4364
rect 10223 4294 10241 4312
rect 10259 4297 10374 4312
rect 20931 4306 21082 4329
rect 10259 4294 10280 4297
rect 10223 4275 10280 4294
rect 20931 4288 20949 4306
rect 20967 4291 21082 4306
rect 31896 4310 32047 4333
rect 42713 4327 42755 4363
rect 31896 4292 31914 4310
rect 31932 4295 32047 4310
rect 42604 4304 42755 4327
rect 31932 4292 31953 4295
rect 20967 4288 20988 4291
rect 20931 4269 20988 4288
rect 31896 4273 31953 4292
rect 42604 4286 42622 4304
rect 42640 4289 42755 4304
rect 42640 4286 42661 4289
rect 42604 4267 42661 4286
rect 553 4206 610 4225
rect 553 4203 574 4206
rect 459 4188 574 4203
rect 592 4188 610 4206
rect 11261 4200 11318 4219
rect 22226 4204 22283 4223
rect 22226 4201 22247 4204
rect 11261 4197 11282 4200
rect 459 4165 610 4188
rect 11167 4182 11282 4197
rect 11300 4182 11318 4200
rect 459 4129 501 4165
rect 11167 4159 11318 4182
rect 22132 4186 22247 4201
rect 22265 4186 22283 4204
rect 32934 4198 32991 4217
rect 32934 4195 32955 4198
rect 22132 4163 22283 4186
rect 32840 4180 32955 4195
rect 32973 4180 32991 4198
rect 458 4128 558 4129
rect 458 4107 614 4128
rect 458 4089 576 4107
rect 594 4089 614 4107
rect 458 4085 614 4089
rect 553 4069 614 4085
rect 11167 4123 11209 4159
rect 22132 4127 22174 4163
rect 32840 4157 32991 4180
rect 22131 4126 22231 4127
rect 11166 4122 11266 4123
rect 11166 4101 11322 4122
rect 553 3951 610 3970
rect 553 3948 574 3951
rect 459 3933 574 3948
rect 592 3933 610 3951
rect 11166 4083 11284 4101
rect 11302 4083 11322 4101
rect 11166 4079 11322 4083
rect 11261 4063 11322 4079
rect 22131 4105 22287 4126
rect 459 3910 610 3933
rect 459 3874 501 3910
rect 458 3873 558 3874
rect 458 3852 614 3873
rect 10219 4020 10280 4036
rect 10219 4016 10375 4020
rect 10219 3998 10239 4016
rect 10257 3998 10375 4016
rect 458 3834 576 3852
rect 594 3834 614 3852
rect 458 3830 614 3834
rect 553 3814 614 3830
rect 10219 3977 10375 3998
rect 10275 3976 10375 3977
rect 10332 3940 10374 3976
rect 11261 3945 11318 3964
rect 11261 3942 11282 3945
rect 10223 3917 10374 3940
rect 10223 3899 10241 3917
rect 10259 3902 10374 3917
rect 11167 3927 11282 3942
rect 11300 3927 11318 3945
rect 22131 4087 22249 4105
rect 22267 4087 22287 4105
rect 22131 4083 22287 4087
rect 22226 4067 22287 4083
rect 32840 4121 32882 4157
rect 32839 4120 32939 4121
rect 32839 4099 32995 4120
rect 11167 3904 11318 3927
rect 10259 3899 10280 3902
rect 10223 3880 10280 3899
rect 11167 3868 11209 3904
rect 11166 3867 11266 3868
rect 11166 3846 11322 3867
rect 20927 4014 20988 4030
rect 20927 4010 21083 4014
rect 20927 3992 20947 4010
rect 20965 3992 21083 4010
rect 11166 3828 11284 3846
rect 11302 3828 11322 3846
rect 11166 3824 11322 3828
rect 11261 3808 11322 3824
rect 20927 3971 21083 3992
rect 20983 3970 21083 3971
rect 10219 3764 10280 3780
rect 21040 3934 21082 3970
rect 22226 3949 22283 3968
rect 22226 3946 22247 3949
rect 20931 3911 21082 3934
rect 20931 3893 20949 3911
rect 20967 3896 21082 3911
rect 22132 3931 22247 3946
rect 22265 3931 22283 3949
rect 32839 4081 32957 4099
rect 32975 4081 32995 4099
rect 32839 4077 32995 4081
rect 32934 4061 32995 4077
rect 22132 3908 22283 3931
rect 20967 3893 20988 3896
rect 20931 3874 20988 3893
rect 22132 3872 22174 3908
rect 22131 3871 22231 3872
rect 10219 3760 10375 3764
rect 10219 3742 10239 3760
rect 10257 3742 10375 3760
rect 10219 3721 10375 3742
rect 22131 3850 22287 3871
rect 31892 4018 31953 4034
rect 31892 4014 32048 4018
rect 31892 3996 31912 4014
rect 31930 3996 32048 4014
rect 22131 3832 22249 3850
rect 22267 3832 22287 3850
rect 22131 3828 22287 3832
rect 22226 3812 22287 3828
rect 31892 3975 32048 3996
rect 31948 3974 32048 3975
rect 20927 3758 20988 3774
rect 32005 3938 32047 3974
rect 32934 3943 32991 3962
rect 32934 3940 32955 3943
rect 31896 3915 32047 3938
rect 31896 3897 31914 3915
rect 31932 3900 32047 3915
rect 32840 3925 32955 3940
rect 32973 3925 32991 3943
rect 32840 3902 32991 3925
rect 31932 3897 31953 3900
rect 31896 3878 31953 3897
rect 20927 3754 21083 3758
rect 10275 3720 10375 3721
rect 10332 3684 10374 3720
rect 20927 3736 20947 3754
rect 20965 3736 21083 3754
rect 20927 3715 21083 3736
rect 32840 3866 32882 3902
rect 32839 3865 32939 3866
rect 32839 3844 32995 3865
rect 42600 4012 42661 4028
rect 42600 4008 42756 4012
rect 42600 3990 42620 4008
rect 42638 3990 42756 4008
rect 32839 3826 32957 3844
rect 32975 3826 32995 3844
rect 32839 3822 32995 3826
rect 32934 3806 32995 3822
rect 42600 3969 42756 3990
rect 42656 3968 42756 3969
rect 31892 3762 31953 3778
rect 42713 3932 42755 3968
rect 42604 3909 42755 3932
rect 42604 3891 42622 3909
rect 42640 3894 42755 3909
rect 42640 3891 42661 3894
rect 42604 3872 42661 3891
rect 31892 3758 32048 3762
rect 20983 3714 21083 3715
rect 10223 3661 10374 3684
rect 21040 3678 21082 3714
rect 31892 3740 31912 3758
rect 31930 3740 32048 3758
rect 31892 3719 32048 3740
rect 42600 3756 42661 3772
rect 42600 3752 42756 3756
rect 31948 3718 32048 3719
rect 32005 3682 32047 3718
rect 42600 3734 42620 3752
rect 42638 3734 42756 3752
rect 42600 3713 42756 3734
rect 42656 3712 42756 3713
rect 10223 3643 10241 3661
rect 10259 3646 10374 3661
rect 20931 3655 21082 3678
rect 10259 3643 10280 3646
rect 10223 3624 10280 3643
rect 20931 3637 20949 3655
rect 20967 3640 21082 3655
rect 31896 3659 32047 3682
rect 42713 3676 42755 3712
rect 31896 3641 31914 3659
rect 31932 3644 32047 3659
rect 42604 3653 42755 3676
rect 31932 3641 31953 3644
rect 20967 3637 20988 3640
rect 20931 3618 20988 3637
rect 31896 3622 31953 3641
rect 42604 3635 42622 3653
rect 42640 3638 42755 3653
rect 42640 3635 42661 3638
rect 42604 3616 42661 3635
rect 553 3410 610 3429
rect 553 3407 574 3410
rect 459 3392 574 3407
rect 592 3392 610 3410
rect 11261 3404 11318 3423
rect 22226 3408 22283 3427
rect 22226 3405 22247 3408
rect 11261 3401 11282 3404
rect 459 3369 610 3392
rect 11167 3386 11282 3401
rect 11300 3386 11318 3404
rect 459 3333 501 3369
rect 11167 3363 11318 3386
rect 22132 3390 22247 3405
rect 22265 3390 22283 3408
rect 32934 3402 32991 3421
rect 32934 3399 32955 3402
rect 22132 3367 22283 3390
rect 32840 3384 32955 3399
rect 32973 3384 32991 3402
rect 458 3332 558 3333
rect 458 3311 614 3332
rect 458 3293 576 3311
rect 594 3293 614 3311
rect 11167 3327 11209 3363
rect 11166 3326 11266 3327
rect 458 3289 614 3293
rect 553 3273 614 3289
rect 11166 3305 11322 3326
rect 11166 3287 11284 3305
rect 11302 3287 11322 3305
rect 22132 3331 22174 3367
rect 32840 3361 32991 3384
rect 22131 3330 22231 3331
rect 11166 3283 11322 3287
rect 553 3154 610 3173
rect 553 3151 574 3154
rect 459 3136 574 3151
rect 592 3136 610 3154
rect 459 3113 610 3136
rect 459 3077 501 3113
rect 11261 3267 11322 3283
rect 458 3076 558 3077
rect 458 3055 614 3076
rect 10219 3223 10280 3239
rect 10219 3219 10375 3223
rect 10219 3201 10239 3219
rect 10257 3201 10375 3219
rect 458 3037 576 3055
rect 594 3037 614 3055
rect 458 3033 614 3037
rect 553 3017 614 3033
rect 10219 3180 10375 3201
rect 10275 3179 10375 3180
rect 10332 3143 10374 3179
rect 22131 3309 22287 3330
rect 22131 3291 22249 3309
rect 22267 3291 22287 3309
rect 32840 3325 32882 3361
rect 32839 3324 32939 3325
rect 22131 3287 22287 3291
rect 11261 3148 11318 3167
rect 11261 3145 11282 3148
rect 10223 3120 10374 3143
rect 10223 3102 10241 3120
rect 10259 3105 10374 3120
rect 11167 3130 11282 3145
rect 11300 3130 11318 3148
rect 11167 3107 11318 3130
rect 10259 3102 10280 3105
rect 10223 3083 10280 3102
rect 11167 3071 11209 3107
rect 22226 3271 22287 3287
rect 11166 3070 11266 3071
rect 11166 3049 11322 3070
rect 20927 3217 20988 3233
rect 20927 3213 21083 3217
rect 20927 3195 20947 3213
rect 20965 3195 21083 3213
rect 11166 3031 11284 3049
rect 11302 3031 11322 3049
rect 11166 3027 11322 3031
rect 11261 3011 11322 3027
rect 20927 3174 21083 3195
rect 32839 3303 32995 3324
rect 32839 3285 32957 3303
rect 32975 3285 32995 3303
rect 32839 3281 32995 3285
rect 20983 3173 21083 3174
rect 21040 3137 21082 3173
rect 22226 3152 22283 3171
rect 22226 3149 22247 3152
rect 20931 3114 21082 3137
rect 10219 2968 10280 2984
rect 10219 2964 10375 2968
rect 10219 2946 10239 2964
rect 10257 2946 10375 2964
rect 20931 3096 20949 3114
rect 20967 3099 21082 3114
rect 22132 3134 22247 3149
rect 22265 3134 22283 3152
rect 22132 3111 22283 3134
rect 20967 3096 20988 3099
rect 20931 3077 20988 3096
rect 22132 3075 22174 3111
rect 32934 3265 32995 3281
rect 22131 3074 22231 3075
rect 22131 3053 22287 3074
rect 31892 3221 31953 3237
rect 31892 3217 32048 3221
rect 31892 3199 31912 3217
rect 31930 3199 32048 3217
rect 22131 3035 22249 3053
rect 22267 3035 22287 3053
rect 22131 3031 22287 3035
rect 22226 3015 22287 3031
rect 31892 3178 32048 3199
rect 31948 3177 32048 3178
rect 32005 3141 32047 3177
rect 32934 3146 32991 3165
rect 32934 3143 32955 3146
rect 31896 3118 32047 3141
rect 10219 2925 10375 2946
rect 10275 2924 10375 2925
rect 10332 2888 10374 2924
rect 20927 2962 20988 2978
rect 20927 2958 21083 2962
rect 20927 2940 20947 2958
rect 20965 2940 21083 2958
rect 31896 3100 31914 3118
rect 31932 3103 32047 3118
rect 32840 3128 32955 3143
rect 32973 3128 32991 3146
rect 32840 3105 32991 3128
rect 31932 3100 31953 3103
rect 31896 3081 31953 3100
rect 32840 3069 32882 3105
rect 32839 3068 32939 3069
rect 32839 3047 32995 3068
rect 42600 3215 42661 3231
rect 42600 3211 42756 3215
rect 42600 3193 42620 3211
rect 42638 3193 42756 3211
rect 32839 3029 32957 3047
rect 32975 3029 32995 3047
rect 32839 3025 32995 3029
rect 32934 3009 32995 3025
rect 42600 3172 42756 3193
rect 42656 3171 42756 3172
rect 42713 3135 42755 3171
rect 42604 3112 42755 3135
rect 20927 2919 21083 2940
rect 31892 2966 31953 2982
rect 31892 2962 32048 2966
rect 31892 2944 31912 2962
rect 31930 2944 32048 2962
rect 42604 3094 42622 3112
rect 42640 3097 42755 3112
rect 42640 3094 42661 3097
rect 42604 3075 42661 3094
rect 31892 2923 32048 2944
rect 31948 2922 32048 2923
rect 20983 2918 21083 2919
rect 10223 2865 10374 2888
rect 21040 2882 21082 2918
rect 32005 2886 32047 2922
rect 42600 2960 42661 2976
rect 42600 2956 42756 2960
rect 42600 2938 42620 2956
rect 42638 2938 42756 2956
rect 42600 2917 42756 2938
rect 42656 2916 42756 2917
rect 10223 2847 10241 2865
rect 10259 2850 10374 2865
rect 20931 2859 21082 2882
rect 10259 2847 10280 2850
rect 10223 2828 10280 2847
rect 20931 2841 20949 2859
rect 20967 2844 21082 2859
rect 31896 2863 32047 2886
rect 42713 2880 42755 2916
rect 31896 2845 31914 2863
rect 31932 2848 32047 2863
rect 42604 2857 42755 2880
rect 31932 2845 31953 2848
rect 20967 2841 20988 2844
rect 20931 2822 20988 2841
rect 31896 2826 31953 2845
rect 42604 2839 42622 2857
rect 42640 2842 42755 2857
rect 42640 2839 42661 2842
rect 42604 2820 42661 2839
rect 553 2759 610 2778
rect 553 2756 574 2759
rect 459 2741 574 2756
rect 592 2741 610 2759
rect 11261 2753 11318 2772
rect 22226 2757 22283 2776
rect 22226 2754 22247 2757
rect 11261 2750 11282 2753
rect 459 2718 610 2741
rect 11167 2735 11282 2750
rect 11300 2735 11318 2753
rect 459 2682 501 2718
rect 11167 2712 11318 2735
rect 22132 2739 22247 2754
rect 22265 2739 22283 2757
rect 32934 2751 32991 2770
rect 32934 2748 32955 2751
rect 22132 2716 22283 2739
rect 32840 2733 32955 2748
rect 32973 2733 32991 2751
rect 458 2681 558 2682
rect 458 2660 614 2681
rect 458 2642 576 2660
rect 594 2642 614 2660
rect 458 2638 614 2642
rect 553 2622 614 2638
rect 11167 2676 11209 2712
rect 22132 2680 22174 2716
rect 32840 2710 32991 2733
rect 22131 2679 22231 2680
rect 11166 2675 11266 2676
rect 11166 2654 11322 2675
rect 553 2504 610 2523
rect 553 2501 574 2504
rect 459 2486 574 2501
rect 592 2486 610 2504
rect 11166 2636 11284 2654
rect 11302 2636 11322 2654
rect 11166 2632 11322 2636
rect 11261 2616 11322 2632
rect 22131 2658 22287 2679
rect 10219 2573 10280 2589
rect 10219 2569 10375 2573
rect 10219 2551 10239 2569
rect 10257 2551 10375 2569
rect 459 2463 610 2486
rect 459 2427 501 2463
rect 458 2426 558 2427
rect 458 2405 614 2426
rect 10219 2530 10375 2551
rect 10275 2529 10375 2530
rect 458 2387 576 2405
rect 594 2387 614 2405
rect 458 2383 614 2387
rect 553 2367 614 2383
rect 10332 2493 10374 2529
rect 11261 2498 11318 2517
rect 11261 2495 11282 2498
rect 10223 2470 10374 2493
rect 10223 2452 10241 2470
rect 10259 2455 10374 2470
rect 11167 2480 11282 2495
rect 11300 2480 11318 2498
rect 22131 2640 22249 2658
rect 22267 2640 22287 2658
rect 22131 2636 22287 2640
rect 22226 2620 22287 2636
rect 32840 2674 32882 2710
rect 32839 2673 32939 2674
rect 32839 2652 32995 2673
rect 20927 2567 20988 2583
rect 20927 2563 21083 2567
rect 20927 2545 20947 2563
rect 20965 2545 21083 2563
rect 11167 2457 11318 2480
rect 10259 2452 10280 2455
rect 10223 2433 10280 2452
rect 11167 2421 11209 2457
rect 11166 2420 11266 2421
rect 11166 2399 11322 2420
rect 20927 2524 21083 2545
rect 20983 2523 21083 2524
rect 11166 2381 11284 2399
rect 11302 2381 11322 2399
rect 11166 2377 11322 2381
rect 11261 2361 11322 2377
rect 10219 2317 10280 2333
rect 21040 2487 21082 2523
rect 22226 2502 22283 2521
rect 22226 2499 22247 2502
rect 20931 2464 21082 2487
rect 20931 2446 20949 2464
rect 20967 2449 21082 2464
rect 22132 2484 22247 2499
rect 22265 2484 22283 2502
rect 32839 2634 32957 2652
rect 32975 2634 32995 2652
rect 32839 2630 32995 2634
rect 32934 2614 32995 2630
rect 31892 2571 31953 2587
rect 31892 2567 32048 2571
rect 31892 2549 31912 2567
rect 31930 2549 32048 2567
rect 22132 2461 22283 2484
rect 20967 2446 20988 2449
rect 20931 2427 20988 2446
rect 22132 2425 22174 2461
rect 22131 2424 22231 2425
rect 10219 2313 10375 2317
rect 10219 2295 10239 2313
rect 10257 2295 10375 2313
rect 10219 2274 10375 2295
rect 10275 2273 10375 2274
rect 22131 2403 22287 2424
rect 31892 2528 32048 2549
rect 31948 2527 32048 2528
rect 22131 2385 22249 2403
rect 22267 2385 22287 2403
rect 22131 2381 22287 2385
rect 22226 2365 22287 2381
rect 20927 2311 20988 2327
rect 32005 2491 32047 2527
rect 32934 2496 32991 2515
rect 32934 2493 32955 2496
rect 31896 2468 32047 2491
rect 31896 2450 31914 2468
rect 31932 2453 32047 2468
rect 32840 2478 32955 2493
rect 32973 2478 32991 2496
rect 42600 2565 42661 2581
rect 42600 2561 42756 2565
rect 42600 2543 42620 2561
rect 42638 2543 42756 2561
rect 32840 2455 32991 2478
rect 31932 2450 31953 2453
rect 31896 2431 31953 2450
rect 20927 2307 21083 2311
rect 10332 2237 10374 2273
rect 20927 2289 20947 2307
rect 20965 2289 21083 2307
rect 20927 2268 21083 2289
rect 32840 2419 32882 2455
rect 32839 2418 32939 2419
rect 32839 2397 32995 2418
rect 42600 2522 42756 2543
rect 42656 2521 42756 2522
rect 32839 2379 32957 2397
rect 32975 2379 32995 2397
rect 32839 2375 32995 2379
rect 32934 2359 32995 2375
rect 31892 2315 31953 2331
rect 42713 2485 42755 2521
rect 42604 2462 42755 2485
rect 42604 2444 42622 2462
rect 42640 2447 42755 2462
rect 42640 2444 42661 2447
rect 42604 2425 42661 2444
rect 31892 2311 32048 2315
rect 20983 2267 21083 2268
rect 10223 2214 10374 2237
rect 21040 2231 21082 2267
rect 31892 2293 31912 2311
rect 31930 2293 32048 2311
rect 31892 2272 32048 2293
rect 31948 2271 32048 2272
rect 42600 2309 42661 2325
rect 42600 2305 42756 2309
rect 32005 2235 32047 2271
rect 42600 2287 42620 2305
rect 42638 2287 42756 2305
rect 42600 2266 42756 2287
rect 42656 2265 42756 2266
rect 10223 2196 10241 2214
rect 10259 2199 10374 2214
rect 20931 2208 21082 2231
rect 10259 2196 10280 2199
rect 10223 2177 10280 2196
rect 20931 2190 20949 2208
rect 20967 2193 21082 2208
rect 31896 2212 32047 2235
rect 42713 2229 42755 2265
rect 31896 2194 31914 2212
rect 31932 2197 32047 2212
rect 42604 2206 42755 2229
rect 31932 2194 31953 2197
rect 20967 2190 20988 2193
rect 20931 2171 20988 2190
rect 31896 2175 31953 2194
rect 42604 2188 42622 2206
rect 42640 2191 42755 2206
rect 42640 2188 42661 2191
rect 42604 2169 42661 2188
<< locali >>
rect 2930 14456 2995 14467
rect 2930 14408 2943 14456
rect 2980 14408 2995 14456
rect 2930 14395 2995 14408
rect 553 13832 612 14215
rect 11261 13966 11320 13971
rect 3143 13915 3854 13917
rect 2516 13914 3854 13915
rect 1466 13913 1538 13914
rect 1465 13905 1564 13913
rect 1465 13902 1517 13905
rect 1465 13867 1473 13902
rect 1498 13867 1517 13902
rect 1542 13894 1564 13905
rect 2515 13906 3854 13914
rect 2515 13903 2567 13906
rect 1542 13893 2409 13894
rect 1542 13867 2410 13893
rect 1465 13857 2410 13867
rect 1465 13855 1564 13857
rect 553 13814 575 13832
rect 593 13814 612 13832
rect 553 13792 612 13814
rect 820 13828 1352 13833
rect 820 13808 1706 13828
rect 1726 13808 1729 13828
rect 2365 13824 2410 13857
rect 2515 13868 2523 13903
rect 2548 13868 2567 13903
rect 2592 13868 3854 13906
rect 2515 13859 3854 13868
rect 2515 13856 2604 13859
rect 3143 13857 3854 13859
rect 820 13804 1729 13808
rect 820 13757 863 13804
rect 1313 13803 1729 13804
rect 2361 13804 2754 13824
rect 2774 13804 2777 13824
rect 1313 13802 1654 13803
rect 970 13771 1080 13785
rect 970 13768 1013 13771
rect 970 13763 974 13768
rect 808 13756 863 13757
rect 552 13733 863 13756
rect 552 13715 577 13733
rect 595 13721 863 13733
rect 892 13741 974 13763
rect 1003 13741 1013 13768
rect 1041 13744 1048 13771
rect 1077 13763 1080 13771
rect 1077 13744 1142 13763
rect 1041 13741 1142 13744
rect 892 13739 1142 13741
rect 595 13715 617 13721
rect 552 13576 617 13715
rect 892 13660 929 13739
rect 970 13726 1080 13739
rect 1044 13670 1075 13671
rect 892 13640 901 13660
rect 921 13640 929 13660
rect 552 13558 575 13576
rect 593 13558 617 13576
rect 552 13541 617 13558
rect 772 13622 840 13635
rect 892 13630 929 13640
rect 988 13660 1075 13670
rect 988 13640 997 13660
rect 1017 13640 1075 13660
rect 988 13631 1075 13640
rect 988 13630 1025 13631
rect 772 13580 779 13622
rect 828 13580 840 13622
rect 772 13577 840 13580
rect 1044 13578 1075 13631
rect 1105 13660 1142 13739
rect 1257 13670 1288 13671
rect 1105 13640 1114 13660
rect 1134 13640 1142 13660
rect 1105 13630 1142 13640
rect 1201 13663 1288 13670
rect 1201 13660 1262 13663
rect 1201 13640 1210 13660
rect 1230 13643 1262 13660
rect 1283 13643 1288 13663
rect 1230 13640 1288 13643
rect 1201 13633 1288 13640
rect 1313 13660 1350 13802
rect 1616 13801 1653 13802
rect 2361 13799 2777 13804
rect 2361 13798 2702 13799
rect 2018 13767 2128 13781
rect 2018 13764 2061 13767
rect 2018 13759 2022 13764
rect 1940 13737 2022 13759
rect 2051 13737 2061 13764
rect 2089 13740 2096 13767
rect 2125 13759 2128 13767
rect 2125 13740 2190 13759
rect 2089 13737 2190 13740
rect 1940 13735 2190 13737
rect 1465 13670 1501 13671
rect 1313 13640 1322 13660
rect 1342 13640 1350 13660
rect 1201 13631 1257 13633
rect 1201 13630 1238 13631
rect 1313 13630 1350 13640
rect 1409 13660 1557 13670
rect 1657 13667 1753 13669
rect 1409 13640 1418 13660
rect 1438 13640 1528 13660
rect 1548 13640 1557 13660
rect 1409 13634 1557 13640
rect 1409 13631 1473 13634
rect 1409 13630 1446 13631
rect 1465 13604 1473 13631
rect 1494 13631 1557 13634
rect 1615 13660 1753 13667
rect 1615 13640 1624 13660
rect 1644 13640 1753 13660
rect 1615 13631 1753 13640
rect 1940 13656 1977 13735
rect 2018 13722 2128 13735
rect 2092 13666 2123 13667
rect 1940 13636 1949 13656
rect 1969 13636 1977 13656
rect 1494 13604 1501 13631
rect 1520 13630 1557 13631
rect 1616 13630 1653 13631
rect 1465 13579 1501 13604
rect 936 13577 977 13578
rect 772 13570 977 13577
rect 772 13559 946 13570
rect 772 13526 780 13559
rect 773 13517 780 13526
rect 829 13550 946 13559
rect 966 13550 977 13570
rect 829 13542 977 13550
rect 1044 13574 1403 13578
rect 1044 13569 1366 13574
rect 1044 13545 1157 13569
rect 1181 13550 1366 13569
rect 1390 13550 1403 13574
rect 1181 13545 1403 13550
rect 1044 13542 1403 13545
rect 1465 13542 1500 13579
rect 1568 13576 1668 13579
rect 1568 13572 1635 13576
rect 1568 13546 1580 13572
rect 1606 13550 1635 13572
rect 1661 13550 1668 13576
rect 1606 13546 1668 13550
rect 1568 13542 1668 13546
rect 829 13526 840 13542
rect 829 13517 837 13526
rect 1044 13521 1075 13542
rect 1465 13521 1501 13542
rect 887 13520 924 13521
rect 552 13477 617 13496
rect 552 13459 577 13477
rect 595 13459 617 13477
rect 552 13258 617 13459
rect 773 13333 837 13517
rect 886 13511 924 13520
rect 886 13491 895 13511
rect 915 13491 924 13511
rect 886 13483 924 13491
rect 990 13515 1075 13521
rect 1100 13520 1137 13521
rect 990 13495 998 13515
rect 1018 13495 1075 13515
rect 990 13487 1075 13495
rect 1099 13511 1137 13520
rect 1099 13491 1108 13511
rect 1128 13491 1137 13511
rect 990 13486 1026 13487
rect 1099 13483 1137 13491
rect 1203 13515 1288 13521
rect 1308 13520 1345 13521
rect 1203 13495 1211 13515
rect 1231 13514 1288 13515
rect 1231 13495 1260 13514
rect 1203 13494 1260 13495
rect 1281 13494 1288 13514
rect 1203 13487 1288 13494
rect 1307 13511 1345 13520
rect 1307 13491 1316 13511
rect 1336 13491 1345 13511
rect 1203 13486 1239 13487
rect 1307 13483 1345 13491
rect 1411 13515 1555 13521
rect 1411 13495 1419 13515
rect 1439 13495 1527 13515
rect 1547 13495 1555 13515
rect 1411 13487 1555 13495
rect 1411 13486 1447 13487
rect 1519 13486 1555 13487
rect 1621 13520 1658 13521
rect 1621 13519 1659 13520
rect 1621 13511 1685 13519
rect 1621 13491 1630 13511
rect 1650 13497 1685 13511
rect 1705 13497 1708 13517
rect 1650 13492 1708 13497
rect 1650 13491 1685 13492
rect 887 13454 924 13483
rect 888 13452 924 13454
rect 1100 13452 1137 13483
rect 888 13430 1137 13452
rect 969 13424 1080 13430
rect 969 13416 1010 13424
rect 969 13396 977 13416
rect 996 13396 1010 13416
rect 969 13394 1010 13396
rect 1038 13416 1080 13424
rect 1038 13396 1054 13416
rect 1073 13396 1080 13416
rect 1038 13394 1080 13396
rect 969 13379 1080 13394
rect 773 13323 841 13333
rect 773 13290 790 13323
rect 830 13290 841 13323
rect 773 13278 841 13290
rect 773 13276 837 13278
rect 1308 13259 1345 13483
rect 1621 13479 1685 13491
rect 1725 13261 1752 13631
rect 1940 13626 1977 13636
rect 2036 13656 2123 13666
rect 2036 13636 2045 13656
rect 2065 13636 2123 13656
rect 2036 13627 2123 13636
rect 2036 13626 2073 13627
rect 1816 13613 1886 13618
rect 1811 13607 1886 13613
rect 1811 13574 1819 13607
rect 1872 13574 1886 13607
rect 2092 13574 2123 13627
rect 2153 13656 2190 13735
rect 2305 13666 2336 13667
rect 2153 13636 2162 13656
rect 2182 13636 2190 13656
rect 2153 13626 2190 13636
rect 2249 13659 2336 13666
rect 2249 13656 2310 13659
rect 2249 13636 2258 13656
rect 2278 13639 2310 13656
rect 2331 13639 2336 13659
rect 2278 13636 2336 13639
rect 2249 13629 2336 13636
rect 2361 13656 2398 13798
rect 2664 13797 2701 13798
rect 2513 13666 2549 13667
rect 2361 13636 2370 13656
rect 2390 13636 2398 13656
rect 2249 13627 2305 13629
rect 2249 13626 2286 13627
rect 2361 13626 2398 13636
rect 2457 13656 2605 13666
rect 2705 13663 2801 13665
rect 2457 13636 2466 13656
rect 2486 13636 2576 13656
rect 2596 13636 2605 13656
rect 2457 13630 2605 13636
rect 2457 13627 2521 13630
rect 2457 13626 2494 13627
rect 2513 13600 2521 13627
rect 2542 13627 2605 13630
rect 2663 13656 2801 13663
rect 2663 13636 2672 13656
rect 2692 13636 2801 13656
rect 2663 13627 2801 13636
rect 2542 13600 2549 13627
rect 2568 13626 2605 13627
rect 2664 13626 2701 13627
rect 2513 13575 2549 13600
rect 1811 13573 1894 13574
rect 1984 13573 2025 13574
rect 1811 13566 2025 13573
rect 1811 13549 1994 13566
rect 1811 13516 1824 13549
rect 1877 13546 1994 13549
rect 2014 13546 2025 13566
rect 1877 13538 2025 13546
rect 2092 13570 2451 13574
rect 2092 13565 2414 13570
rect 2092 13541 2205 13565
rect 2229 13546 2414 13565
rect 2438 13546 2451 13570
rect 2229 13541 2451 13546
rect 2092 13538 2451 13541
rect 2513 13538 2548 13575
rect 2616 13572 2716 13575
rect 2616 13568 2683 13572
rect 2616 13542 2628 13568
rect 2654 13546 2683 13568
rect 2709 13546 2716 13572
rect 2654 13542 2716 13546
rect 2616 13538 2716 13542
rect 1877 13516 1894 13538
rect 2092 13517 2123 13538
rect 2513 13517 2549 13538
rect 1935 13516 1972 13517
rect 1811 13502 1894 13516
rect 1584 13259 1752 13261
rect 1308 13258 1752 13259
rect 552 13228 1752 13258
rect 1822 13292 1894 13502
rect 1934 13507 1972 13516
rect 1934 13487 1943 13507
rect 1963 13487 1972 13507
rect 1934 13479 1972 13487
rect 2038 13511 2123 13517
rect 2148 13516 2185 13517
rect 2038 13491 2046 13511
rect 2066 13491 2123 13511
rect 2038 13483 2123 13491
rect 2147 13507 2185 13516
rect 2147 13487 2156 13507
rect 2176 13487 2185 13507
rect 2038 13482 2074 13483
rect 2147 13479 2185 13487
rect 2251 13511 2336 13517
rect 2356 13516 2393 13517
rect 2251 13491 2259 13511
rect 2279 13510 2336 13511
rect 2279 13491 2308 13510
rect 2251 13490 2308 13491
rect 2329 13490 2336 13510
rect 2251 13483 2336 13490
rect 2355 13507 2393 13516
rect 2355 13487 2364 13507
rect 2384 13487 2393 13507
rect 2251 13482 2287 13483
rect 2355 13479 2393 13487
rect 2459 13511 2603 13517
rect 2459 13491 2467 13511
rect 2487 13491 2575 13511
rect 2595 13491 2603 13511
rect 2459 13483 2603 13491
rect 2459 13482 2495 13483
rect 2567 13482 2603 13483
rect 2669 13516 2706 13517
rect 2669 13515 2707 13516
rect 2669 13507 2733 13515
rect 2669 13487 2678 13507
rect 2698 13493 2733 13507
rect 2753 13493 2756 13513
rect 2698 13488 2756 13493
rect 2698 13487 2733 13488
rect 1935 13450 1972 13479
rect 1936 13448 1972 13450
rect 2148 13448 2185 13479
rect 1936 13426 2185 13448
rect 2017 13420 2128 13426
rect 2017 13412 2058 13420
rect 2017 13392 2025 13412
rect 2044 13392 2058 13412
rect 2017 13390 2058 13392
rect 2086 13412 2128 13420
rect 2086 13392 2102 13412
rect 2121 13392 2128 13412
rect 2086 13390 2128 13392
rect 2017 13375 2128 13390
rect 1822 13253 1841 13292
rect 1886 13253 1894 13292
rect 1822 13236 1894 13253
rect 2356 13280 2393 13479
rect 2669 13475 2733 13487
rect 2356 13274 2397 13280
rect 2773 13276 2800 13627
rect 3095 13614 3190 13640
rect 2931 13592 2995 13611
rect 2931 13553 2944 13592
rect 2978 13553 2995 13592
rect 2931 13534 2995 13553
rect 2632 13274 2800 13276
rect 2356 13248 2800 13274
rect 552 13181 617 13228
rect 552 13163 575 13181
rect 593 13163 617 13181
rect 1465 13208 1500 13210
rect 1465 13206 1569 13208
rect 2358 13206 2397 13248
rect 2632 13247 2800 13248
rect 1465 13199 2399 13206
rect 1465 13198 1516 13199
rect 1465 13178 1468 13198
rect 1493 13179 1516 13198
rect 1548 13179 2399 13199
rect 1493 13178 2399 13179
rect 1465 13171 2399 13178
rect 1738 13170 2399 13171
rect 552 13142 617 13163
rect 829 13153 869 13156
rect 829 13149 1732 13153
rect 829 13129 1706 13149
rect 1726 13129 1732 13149
rect 829 13126 1732 13129
rect 553 13082 618 13102
rect 553 13064 577 13082
rect 595 13064 618 13082
rect 553 13037 618 13064
rect 829 13037 869 13126
rect 1313 13124 1729 13126
rect 1313 13123 1654 13124
rect 970 13092 1080 13106
rect 970 13089 1013 13092
rect 970 13084 974 13089
rect 552 13002 869 13037
rect 892 13062 974 13084
rect 1003 13062 1013 13089
rect 1041 13065 1048 13092
rect 1077 13084 1080 13092
rect 1077 13065 1142 13084
rect 1041 13062 1142 13065
rect 892 13060 1142 13062
rect 553 12926 618 13002
rect 892 12981 929 13060
rect 970 13047 1080 13060
rect 1044 12991 1075 12992
rect 892 12961 901 12981
rect 921 12961 929 12981
rect 892 12951 929 12961
rect 988 12981 1075 12991
rect 988 12961 997 12981
rect 1017 12961 1075 12981
rect 988 12952 1075 12961
rect 988 12951 1025 12952
rect 553 12908 575 12926
rect 593 12908 618 12926
rect 553 12887 618 12908
rect 766 12906 831 12915
rect 766 12869 776 12906
rect 816 12898 831 12906
rect 1044 12899 1075 12952
rect 1105 12981 1142 13060
rect 1257 12991 1288 12992
rect 1105 12961 1114 12981
rect 1134 12961 1142 12981
rect 1105 12951 1142 12961
rect 1201 12984 1288 12991
rect 1201 12981 1262 12984
rect 1201 12961 1210 12981
rect 1230 12964 1262 12981
rect 1283 12964 1288 12984
rect 1230 12961 1288 12964
rect 1201 12954 1288 12961
rect 1313 12981 1350 13123
rect 1616 13122 1653 13123
rect 2933 13063 2995 13534
rect 3095 13573 3121 13614
rect 3157 13573 3190 13614
rect 3095 13277 3190 13573
rect 3095 13233 3110 13277
rect 3170 13233 3190 13277
rect 3095 13213 3190 13233
rect 3807 13144 3850 13857
rect 4883 13747 5776 13787
rect 4883 13680 4916 13747
rect 5002 13680 5784 13747
rect 8949 13683 9019 13936
rect 9488 13933 9529 13935
rect 9760 13933 9864 13935
rect 10200 13933 11323 13966
rect 32934 13964 32993 13969
rect 9081 13898 11323 13933
rect 13851 13909 14562 13911
rect 12174 13907 12246 13908
rect 13732 13907 14562 13909
rect 9081 13884 9109 13898
rect 9083 13753 9109 13884
rect 9488 13896 11323 13898
rect 9488 13895 9631 13896
rect 9889 13895 11323 13896
rect 4883 13612 5784 13680
rect 4892 13611 4998 13612
rect 5667 13518 5784 13612
rect 8941 13632 9021 13683
rect 8941 13606 8957 13632
rect 8997 13606 9021 13632
rect 8941 13587 9021 13606
rect 8941 13561 8960 13587
rect 9000 13561 9021 13587
rect 8941 13534 9021 13561
rect 3807 13124 4201 13144
rect 4221 13124 4224 13144
rect 3808 13119 4224 13124
rect 3808 13118 4149 13119
rect 3465 13087 3575 13101
rect 3465 13084 3508 13087
rect 3465 13079 3469 13084
rect 2928 13011 3003 13063
rect 3387 13057 3469 13079
rect 3498 13057 3508 13084
rect 3536 13060 3543 13087
rect 3572 13079 3575 13087
rect 3572 13060 3637 13079
rect 3536 13057 3637 13060
rect 3387 13055 3637 13057
rect 3297 13011 3343 13012
rect 1465 12991 1501 12992
rect 1313 12961 1322 12981
rect 1342 12961 1350 12981
rect 1201 12952 1257 12954
rect 1201 12951 1238 12952
rect 1313 12951 1350 12961
rect 1409 12981 1557 12991
rect 1657 12988 1753 12990
rect 1409 12961 1418 12981
rect 1438 12961 1528 12981
rect 1548 12961 1557 12981
rect 1409 12955 1557 12961
rect 1409 12952 1473 12955
rect 1409 12951 1446 12952
rect 1465 12925 1473 12952
rect 1494 12952 1557 12955
rect 1615 12981 1753 12988
rect 1615 12961 1624 12981
rect 1644 12961 1753 12981
rect 1615 12952 1753 12961
rect 2928 12976 3343 13011
rect 1494 12925 1501 12952
rect 1520 12951 1557 12952
rect 1616 12951 1653 12952
rect 1465 12900 1501 12925
rect 936 12898 977 12899
rect 816 12891 977 12898
rect 816 12871 946 12891
rect 966 12871 977 12891
rect 816 12869 977 12871
rect 766 12863 977 12869
rect 1044 12895 1403 12899
rect 1044 12890 1366 12895
rect 1044 12866 1157 12890
rect 1181 12871 1366 12890
rect 1390 12871 1403 12895
rect 1181 12866 1403 12871
rect 1044 12863 1403 12866
rect 1465 12863 1500 12900
rect 1568 12897 1668 12900
rect 1568 12893 1635 12897
rect 1568 12867 1580 12893
rect 1606 12871 1635 12893
rect 1661 12871 1668 12897
rect 1606 12867 1668 12871
rect 1568 12863 1668 12867
rect 766 12850 833 12863
rect 558 12827 614 12847
rect 558 12809 577 12827
rect 595 12809 614 12827
rect 558 12696 614 12809
rect 766 12829 780 12850
rect 816 12829 833 12850
rect 1044 12842 1075 12863
rect 1465 12842 1501 12863
rect 887 12841 924 12842
rect 766 12822 833 12829
rect 886 12832 924 12841
rect 558 12558 613 12696
rect 766 12670 831 12822
rect 886 12812 895 12832
rect 915 12812 924 12832
rect 886 12804 924 12812
rect 990 12836 1075 12842
rect 1100 12841 1137 12842
rect 990 12816 998 12836
rect 1018 12816 1075 12836
rect 990 12808 1075 12816
rect 1099 12832 1137 12841
rect 1099 12812 1108 12832
rect 1128 12812 1137 12832
rect 990 12807 1026 12808
rect 1099 12804 1137 12812
rect 1203 12836 1288 12842
rect 1308 12841 1345 12842
rect 1203 12816 1211 12836
rect 1231 12835 1288 12836
rect 1231 12816 1260 12835
rect 1203 12815 1260 12816
rect 1281 12815 1288 12835
rect 1203 12808 1288 12815
rect 1307 12832 1345 12841
rect 1307 12812 1316 12832
rect 1336 12812 1345 12832
rect 1203 12807 1239 12808
rect 1307 12804 1345 12812
rect 1411 12836 1555 12842
rect 1411 12816 1419 12836
rect 1439 12816 1527 12836
rect 1547 12816 1555 12836
rect 1411 12808 1555 12816
rect 1411 12807 1447 12808
rect 1519 12807 1555 12808
rect 1621 12841 1658 12842
rect 1621 12840 1659 12841
rect 1621 12832 1685 12840
rect 1621 12812 1630 12832
rect 1650 12818 1685 12832
rect 1705 12818 1708 12838
rect 1650 12813 1708 12818
rect 1650 12812 1685 12813
rect 887 12775 924 12804
rect 888 12773 924 12775
rect 1100 12773 1137 12804
rect 888 12751 1137 12773
rect 969 12745 1080 12751
rect 969 12737 1010 12745
rect 969 12717 977 12737
rect 996 12717 1010 12737
rect 969 12715 1010 12717
rect 1038 12737 1080 12745
rect 1038 12717 1054 12737
rect 1073 12717 1080 12737
rect 1038 12715 1080 12717
rect 969 12702 1080 12715
rect 1308 12705 1345 12804
rect 1621 12800 1685 12812
rect 759 12660 880 12670
rect 759 12658 828 12660
rect 759 12617 772 12658
rect 809 12619 828 12658
rect 865 12619 880 12660
rect 809 12617 880 12619
rect 759 12599 880 12617
rect 551 12555 615 12558
rect 971 12555 1075 12561
rect 1306 12555 1347 12705
rect 1725 12697 1752 12952
rect 1814 12942 1894 12953
rect 1814 12916 1831 12942
rect 1871 12916 1894 12942
rect 1814 12889 1894 12916
rect 1814 12863 1835 12889
rect 1875 12863 1894 12889
rect 1814 12844 1894 12863
rect 1814 12818 1838 12844
rect 1878 12818 1894 12844
rect 1814 12767 1894 12818
rect 551 12552 1347 12555
rect 1726 12566 1752 12697
rect 1726 12552 1754 12566
rect 551 12517 1754 12552
rect 1816 12559 1886 12767
rect 2928 12692 3003 12976
rect 3297 12893 3343 12976
rect 3387 12976 3424 13055
rect 3465 13042 3575 13055
rect 3539 12986 3570 12987
rect 3387 12956 3396 12976
rect 3416 12956 3424 12976
rect 3387 12946 3424 12956
rect 3483 12976 3570 12986
rect 3483 12956 3492 12976
rect 3512 12956 3570 12976
rect 3483 12947 3570 12956
rect 3483 12946 3520 12947
rect 3539 12894 3570 12947
rect 3600 12976 3637 13055
rect 3752 12986 3783 12987
rect 3600 12956 3609 12976
rect 3629 12956 3637 12976
rect 3600 12946 3637 12956
rect 3696 12979 3783 12986
rect 3696 12976 3757 12979
rect 3696 12956 3705 12976
rect 3725 12959 3757 12976
rect 3778 12959 3783 12979
rect 3725 12956 3783 12959
rect 3696 12949 3783 12956
rect 3808 12976 3845 13118
rect 4111 13117 4148 13118
rect 3960 12986 3996 12987
rect 3808 12956 3817 12976
rect 3837 12956 3845 12976
rect 3696 12947 3752 12949
rect 3696 12946 3733 12947
rect 3808 12946 3845 12956
rect 3904 12976 4052 12986
rect 4152 12983 4248 12985
rect 3904 12956 3913 12976
rect 3933 12956 4023 12976
rect 4043 12956 4052 12976
rect 3904 12950 4052 12956
rect 3904 12947 3968 12950
rect 3904 12946 3941 12947
rect 3960 12920 3968 12947
rect 3989 12947 4052 12950
rect 4110 12976 4248 12983
rect 4110 12956 4119 12976
rect 4139 12956 4248 12976
rect 4110 12947 4248 12956
rect 3989 12920 3996 12947
rect 4015 12946 4052 12947
rect 4111 12946 4148 12947
rect 3960 12895 3996 12920
rect 3431 12893 3472 12894
rect 3297 12886 3472 12893
rect 3095 12860 3181 12879
rect 3095 12819 3110 12860
rect 3164 12819 3181 12860
rect 3297 12866 3441 12886
rect 3461 12866 3472 12886
rect 3297 12858 3472 12866
rect 3539 12890 3898 12894
rect 3539 12885 3861 12890
rect 3539 12861 3652 12885
rect 3676 12866 3861 12885
rect 3885 12866 3898 12890
rect 3676 12861 3898 12866
rect 3539 12858 3898 12861
rect 3960 12858 3995 12895
rect 4063 12892 4163 12895
rect 4063 12888 4130 12892
rect 4063 12862 4075 12888
rect 4101 12866 4130 12888
rect 4156 12866 4163 12892
rect 4101 12862 4163 12866
rect 4063 12858 4163 12862
rect 3297 12854 3343 12858
rect 3539 12837 3570 12858
rect 3960 12837 3996 12858
rect 3382 12836 3419 12837
rect 3095 12783 3181 12819
rect 3381 12827 3419 12836
rect 3381 12807 3390 12827
rect 3410 12807 3419 12827
rect 3381 12799 3419 12807
rect 3485 12831 3570 12837
rect 3595 12836 3632 12837
rect 3485 12811 3493 12831
rect 3513 12811 3570 12831
rect 3485 12803 3570 12811
rect 3594 12827 3632 12836
rect 3594 12807 3603 12827
rect 3623 12807 3632 12827
rect 3485 12802 3521 12803
rect 3594 12799 3632 12807
rect 3698 12831 3783 12837
rect 3803 12836 3840 12837
rect 3698 12811 3706 12831
rect 3726 12830 3783 12831
rect 3726 12811 3755 12830
rect 3698 12810 3755 12811
rect 3776 12810 3783 12830
rect 3698 12803 3783 12810
rect 3802 12827 3840 12836
rect 3802 12807 3811 12827
rect 3831 12807 3840 12827
rect 3698 12802 3734 12803
rect 3802 12799 3840 12807
rect 3906 12831 4050 12837
rect 3906 12811 3914 12831
rect 3934 12811 4022 12831
rect 4042 12811 4050 12831
rect 3906 12803 4050 12811
rect 3906 12802 3942 12803
rect 551 12456 615 12517
rect 971 12515 1075 12517
rect 1306 12515 1347 12517
rect 1816 12514 1837 12559
rect 1817 12493 1837 12514
rect 1867 12514 1886 12559
rect 2923 12650 3003 12692
rect 1867 12493 1884 12514
rect 1817 12474 1884 12493
rect 1466 12466 1538 12467
rect 1465 12458 1564 12466
rect 553 12385 612 12456
rect 1465 12455 1517 12458
rect 1465 12420 1473 12455
rect 1498 12420 1517 12455
rect 1542 12447 1564 12458
rect 1542 12446 2409 12447
rect 1542 12420 2410 12446
rect 1465 12410 2410 12420
rect 1465 12408 1564 12410
rect 553 12367 575 12385
rect 593 12367 612 12385
rect 553 12345 612 12367
rect 820 12381 1352 12386
rect 820 12361 1706 12381
rect 1726 12361 1729 12381
rect 2365 12377 2410 12410
rect 820 12357 1729 12361
rect 820 12310 863 12357
rect 1313 12356 1729 12357
rect 2361 12357 2754 12377
rect 2774 12357 2777 12377
rect 1313 12355 1654 12356
rect 970 12324 1080 12338
rect 970 12321 1013 12324
rect 970 12316 974 12321
rect 808 12309 863 12310
rect 552 12286 863 12309
rect 552 12268 577 12286
rect 595 12274 863 12286
rect 892 12294 974 12316
rect 1003 12294 1013 12321
rect 1041 12297 1048 12324
rect 1077 12316 1080 12324
rect 1077 12297 1142 12316
rect 1041 12294 1142 12297
rect 892 12292 1142 12294
rect 595 12268 617 12274
rect 552 12129 617 12268
rect 892 12213 929 12292
rect 970 12279 1080 12292
rect 1044 12223 1075 12224
rect 892 12193 901 12213
rect 921 12193 929 12213
rect 552 12111 575 12129
rect 593 12111 617 12129
rect 552 12094 617 12111
rect 772 12175 840 12188
rect 892 12183 929 12193
rect 988 12213 1075 12223
rect 988 12193 997 12213
rect 1017 12193 1075 12213
rect 988 12184 1075 12193
rect 988 12183 1025 12184
rect 772 12133 779 12175
rect 828 12133 840 12175
rect 772 12130 840 12133
rect 1044 12131 1075 12184
rect 1105 12213 1142 12292
rect 1257 12223 1288 12224
rect 1105 12193 1114 12213
rect 1134 12193 1142 12213
rect 1105 12183 1142 12193
rect 1201 12216 1288 12223
rect 1201 12213 1262 12216
rect 1201 12193 1210 12213
rect 1230 12196 1262 12213
rect 1283 12196 1288 12216
rect 1230 12193 1288 12196
rect 1201 12186 1288 12193
rect 1313 12213 1350 12355
rect 1616 12354 1653 12355
rect 2361 12352 2777 12357
rect 2361 12351 2702 12352
rect 2018 12320 2128 12334
rect 2018 12317 2061 12320
rect 2018 12312 2022 12317
rect 1940 12290 2022 12312
rect 2051 12290 2061 12317
rect 2089 12293 2096 12320
rect 2125 12312 2128 12320
rect 2125 12293 2190 12312
rect 2089 12290 2190 12293
rect 1940 12288 2190 12290
rect 1465 12223 1501 12224
rect 1313 12193 1322 12213
rect 1342 12193 1350 12213
rect 1201 12184 1257 12186
rect 1201 12183 1238 12184
rect 1313 12183 1350 12193
rect 1409 12213 1557 12223
rect 1657 12220 1753 12222
rect 1409 12193 1418 12213
rect 1438 12193 1528 12213
rect 1548 12193 1557 12213
rect 1409 12187 1557 12193
rect 1409 12184 1473 12187
rect 1409 12183 1446 12184
rect 1465 12157 1473 12184
rect 1494 12184 1557 12187
rect 1615 12213 1753 12220
rect 1615 12193 1624 12213
rect 1644 12193 1753 12213
rect 1615 12184 1753 12193
rect 1940 12209 1977 12288
rect 2018 12275 2128 12288
rect 2092 12219 2123 12220
rect 1940 12189 1949 12209
rect 1969 12189 1977 12209
rect 1494 12157 1501 12184
rect 1520 12183 1557 12184
rect 1616 12183 1653 12184
rect 1465 12132 1501 12157
rect 936 12130 977 12131
rect 772 12123 977 12130
rect 772 12112 946 12123
rect 772 12079 780 12112
rect 773 12070 780 12079
rect 829 12103 946 12112
rect 966 12103 977 12123
rect 829 12095 977 12103
rect 1044 12127 1403 12131
rect 1044 12122 1366 12127
rect 1044 12098 1157 12122
rect 1181 12103 1366 12122
rect 1390 12103 1403 12127
rect 1181 12098 1403 12103
rect 1044 12095 1403 12098
rect 1465 12095 1500 12132
rect 1568 12129 1668 12132
rect 1568 12125 1635 12129
rect 1568 12099 1580 12125
rect 1606 12103 1635 12125
rect 1661 12103 1668 12129
rect 1606 12099 1668 12103
rect 1568 12095 1668 12099
rect 829 12079 840 12095
rect 829 12070 837 12079
rect 1044 12074 1075 12095
rect 1465 12074 1501 12095
rect 887 12073 924 12074
rect 552 12030 617 12049
rect 552 12012 577 12030
rect 595 12012 617 12030
rect 552 11811 617 12012
rect 773 11886 837 12070
rect 886 12064 924 12073
rect 886 12044 895 12064
rect 915 12044 924 12064
rect 886 12036 924 12044
rect 990 12068 1075 12074
rect 1100 12073 1137 12074
rect 990 12048 998 12068
rect 1018 12048 1075 12068
rect 990 12040 1075 12048
rect 1099 12064 1137 12073
rect 1099 12044 1108 12064
rect 1128 12044 1137 12064
rect 990 12039 1026 12040
rect 1099 12036 1137 12044
rect 1203 12068 1288 12074
rect 1308 12073 1345 12074
rect 1203 12048 1211 12068
rect 1231 12067 1288 12068
rect 1231 12048 1260 12067
rect 1203 12047 1260 12048
rect 1281 12047 1288 12067
rect 1203 12040 1288 12047
rect 1307 12064 1345 12073
rect 1307 12044 1316 12064
rect 1336 12044 1345 12064
rect 1203 12039 1239 12040
rect 1307 12036 1345 12044
rect 1411 12068 1555 12074
rect 1411 12048 1419 12068
rect 1439 12048 1527 12068
rect 1547 12048 1555 12068
rect 1411 12040 1555 12048
rect 1411 12039 1447 12040
rect 1519 12039 1555 12040
rect 1621 12073 1658 12074
rect 1621 12072 1659 12073
rect 1621 12064 1685 12072
rect 1621 12044 1630 12064
rect 1650 12050 1685 12064
rect 1705 12050 1708 12070
rect 1650 12045 1708 12050
rect 1650 12044 1685 12045
rect 887 12007 924 12036
rect 888 12005 924 12007
rect 1100 12005 1137 12036
rect 888 11983 1137 12005
rect 969 11977 1080 11983
rect 969 11969 1010 11977
rect 969 11949 977 11969
rect 996 11949 1010 11969
rect 969 11947 1010 11949
rect 1038 11969 1080 11977
rect 1038 11949 1054 11969
rect 1073 11949 1080 11969
rect 1038 11947 1080 11949
rect 969 11932 1080 11947
rect 773 11876 841 11886
rect 773 11843 790 11876
rect 830 11843 841 11876
rect 773 11831 841 11843
rect 773 11829 837 11831
rect 1308 11812 1345 12036
rect 1621 12032 1685 12044
rect 1725 11814 1752 12184
rect 1940 12179 1977 12189
rect 2036 12209 2123 12219
rect 2036 12189 2045 12209
rect 2065 12189 2123 12209
rect 2036 12180 2123 12189
rect 2036 12179 2073 12180
rect 1816 12166 1886 12171
rect 1811 12160 1886 12166
rect 1811 12127 1819 12160
rect 1872 12127 1886 12160
rect 2092 12127 2123 12180
rect 2153 12209 2190 12288
rect 2305 12219 2336 12220
rect 2153 12189 2162 12209
rect 2182 12189 2190 12209
rect 2153 12179 2190 12189
rect 2249 12212 2336 12219
rect 2249 12209 2310 12212
rect 2249 12189 2258 12209
rect 2278 12192 2310 12209
rect 2331 12192 2336 12212
rect 2278 12189 2336 12192
rect 2249 12182 2336 12189
rect 2361 12209 2398 12351
rect 2664 12350 2701 12351
rect 2513 12219 2549 12220
rect 2361 12189 2370 12209
rect 2390 12189 2398 12209
rect 2249 12180 2305 12182
rect 2249 12179 2286 12180
rect 2361 12179 2398 12189
rect 2457 12209 2605 12219
rect 2705 12216 2801 12218
rect 2457 12189 2466 12209
rect 2486 12189 2576 12209
rect 2596 12189 2605 12209
rect 2457 12183 2605 12189
rect 2457 12180 2521 12183
rect 2457 12179 2494 12180
rect 2513 12153 2521 12180
rect 2542 12180 2605 12183
rect 2663 12209 2801 12216
rect 2663 12189 2672 12209
rect 2692 12189 2801 12209
rect 2663 12180 2801 12189
rect 2542 12153 2549 12180
rect 2568 12179 2605 12180
rect 2664 12179 2701 12180
rect 2513 12128 2549 12153
rect 1811 12126 1894 12127
rect 1984 12126 2025 12127
rect 1811 12119 2025 12126
rect 1811 12102 1994 12119
rect 1811 12069 1824 12102
rect 1877 12099 1994 12102
rect 2014 12099 2025 12119
rect 1877 12091 2025 12099
rect 2092 12123 2451 12127
rect 2092 12118 2414 12123
rect 2092 12094 2205 12118
rect 2229 12099 2414 12118
rect 2438 12099 2451 12123
rect 2229 12094 2451 12099
rect 2092 12091 2451 12094
rect 2513 12091 2548 12128
rect 2616 12125 2716 12128
rect 2616 12121 2683 12125
rect 2616 12095 2628 12121
rect 2654 12099 2683 12121
rect 2709 12099 2716 12125
rect 2654 12095 2716 12099
rect 2616 12091 2716 12095
rect 1877 12069 1894 12091
rect 2092 12070 2123 12091
rect 2513 12070 2549 12091
rect 1935 12069 1972 12070
rect 1811 12055 1894 12069
rect 1584 11812 1752 11814
rect 1308 11811 1752 11812
rect 552 11781 1752 11811
rect 1822 11845 1894 12055
rect 1934 12060 1972 12069
rect 1934 12040 1943 12060
rect 1963 12040 1972 12060
rect 1934 12032 1972 12040
rect 2038 12064 2123 12070
rect 2148 12069 2185 12070
rect 2038 12044 2046 12064
rect 2066 12044 2123 12064
rect 2038 12036 2123 12044
rect 2147 12060 2185 12069
rect 2147 12040 2156 12060
rect 2176 12040 2185 12060
rect 2038 12035 2074 12036
rect 2147 12032 2185 12040
rect 2251 12064 2336 12070
rect 2356 12069 2393 12070
rect 2251 12044 2259 12064
rect 2279 12063 2336 12064
rect 2279 12044 2308 12063
rect 2251 12043 2308 12044
rect 2329 12043 2336 12063
rect 2251 12036 2336 12043
rect 2355 12060 2393 12069
rect 2355 12040 2364 12060
rect 2384 12040 2393 12060
rect 2251 12035 2287 12036
rect 2355 12032 2393 12040
rect 2459 12064 2603 12070
rect 2459 12044 2467 12064
rect 2487 12044 2575 12064
rect 2595 12044 2603 12064
rect 2459 12036 2603 12044
rect 2459 12035 2495 12036
rect 2567 12035 2603 12036
rect 2669 12069 2706 12070
rect 2669 12068 2707 12069
rect 2669 12060 2733 12068
rect 2669 12040 2678 12060
rect 2698 12046 2733 12060
rect 2753 12046 2756 12066
rect 2698 12041 2756 12046
rect 2698 12040 2733 12041
rect 1935 12003 1972 12032
rect 1936 12001 1972 12003
rect 2148 12001 2185 12032
rect 1936 11979 2185 12001
rect 2017 11973 2128 11979
rect 2017 11965 2058 11973
rect 2017 11945 2025 11965
rect 2044 11945 2058 11965
rect 2017 11943 2058 11945
rect 2086 11965 2128 11973
rect 2086 11945 2102 11965
rect 2121 11945 2128 11965
rect 2086 11943 2128 11945
rect 2017 11928 2128 11943
rect 1822 11806 1841 11845
rect 1886 11806 1894 11845
rect 1822 11789 1894 11806
rect 2356 11833 2393 12032
rect 2669 12028 2733 12040
rect 2356 11827 2397 11833
rect 2773 11829 2800 12180
rect 2923 12050 3002 12650
rect 3099 12198 3178 12783
rect 3382 12770 3419 12799
rect 3383 12768 3419 12770
rect 3595 12768 3632 12799
rect 3383 12746 3632 12768
rect 3464 12740 3575 12746
rect 3464 12732 3505 12740
rect 3464 12712 3472 12732
rect 3491 12712 3505 12732
rect 3464 12710 3505 12712
rect 3533 12732 3575 12740
rect 3533 12712 3549 12732
rect 3568 12712 3575 12732
rect 3533 12710 3575 12712
rect 3464 12695 3575 12710
rect 3803 12684 3840 12799
rect 3796 12572 3843 12684
rect 3964 12644 3994 12803
rect 4014 12802 4050 12803
rect 4116 12836 4153 12837
rect 4116 12835 4154 12836
rect 4116 12827 4180 12835
rect 4116 12807 4125 12827
rect 4145 12813 4180 12827
rect 4200 12813 4203 12833
rect 4145 12808 4203 12813
rect 4145 12807 4180 12808
rect 4116 12795 4180 12807
rect 3964 12640 4050 12644
rect 3964 12622 3979 12640
rect 4031 12622 4050 12640
rect 3964 12613 4050 12622
rect 4220 12574 4247 12947
rect 4079 12572 4247 12574
rect 3796 12546 4247 12572
rect 3796 12468 3843 12546
rect 4079 12545 4247 12546
rect 3741 12467 3843 12468
rect 3740 12459 3843 12467
rect 3740 12456 3792 12459
rect 3740 12421 3748 12456
rect 3773 12421 3792 12456
rect 3817 12421 3843 12459
rect 3740 12415 3843 12421
rect 4003 12460 4039 12464
rect 4003 12437 4011 12460
rect 4035 12437 4039 12460
rect 4003 12416 4039 12437
rect 3740 12411 3839 12415
rect 4003 12393 4011 12416
rect 4035 12393 4039 12416
rect 2632 11827 2800 11829
rect 2356 11801 2800 11827
rect 552 11734 617 11781
rect 552 11716 575 11734
rect 593 11716 617 11734
rect 1465 11761 1500 11763
rect 1465 11759 1569 11761
rect 2358 11759 2397 11801
rect 2632 11800 2800 11801
rect 1465 11752 2399 11759
rect 1465 11751 1516 11752
rect 1465 11731 1468 11751
rect 1493 11732 1516 11751
rect 1548 11732 2399 11752
rect 1493 11731 2399 11732
rect 1465 11724 2399 11731
rect 1738 11723 2399 11724
rect 552 11695 617 11716
rect 829 11706 869 11709
rect 829 11702 1732 11706
rect 829 11682 1706 11702
rect 1726 11682 1732 11702
rect 829 11679 1732 11682
rect 553 11635 618 11655
rect 553 11617 577 11635
rect 595 11617 618 11635
rect 553 11590 618 11617
rect 829 11590 869 11679
rect 1313 11677 1729 11679
rect 1313 11676 1654 11677
rect 970 11645 1080 11659
rect 970 11642 1013 11645
rect 970 11637 974 11642
rect 552 11555 869 11590
rect 892 11615 974 11637
rect 1003 11615 1013 11642
rect 1041 11618 1048 11645
rect 1077 11637 1080 11645
rect 1077 11618 1142 11637
rect 1041 11615 1142 11618
rect 892 11613 1142 11615
rect 553 11479 618 11555
rect 892 11534 929 11613
rect 970 11600 1080 11613
rect 1044 11544 1075 11545
rect 892 11514 901 11534
rect 921 11514 929 11534
rect 892 11504 929 11514
rect 988 11534 1075 11544
rect 988 11514 997 11534
rect 1017 11514 1075 11534
rect 988 11505 1075 11514
rect 988 11504 1025 11505
rect 553 11461 575 11479
rect 593 11461 618 11479
rect 553 11440 618 11461
rect 766 11459 831 11468
rect 766 11422 776 11459
rect 816 11451 831 11459
rect 1044 11452 1075 11505
rect 1105 11534 1142 11613
rect 1257 11544 1288 11545
rect 1105 11514 1114 11534
rect 1134 11514 1142 11534
rect 1105 11504 1142 11514
rect 1201 11537 1288 11544
rect 1201 11534 1262 11537
rect 1201 11514 1210 11534
rect 1230 11517 1262 11534
rect 1283 11517 1288 11537
rect 1230 11514 1288 11517
rect 1201 11507 1288 11514
rect 1313 11534 1350 11676
rect 1616 11675 1653 11676
rect 1465 11544 1501 11545
rect 1313 11514 1322 11534
rect 1342 11514 1350 11534
rect 1201 11505 1257 11507
rect 1201 11504 1238 11505
rect 1313 11504 1350 11514
rect 1409 11534 1557 11544
rect 1657 11541 1753 11543
rect 1409 11514 1418 11534
rect 1438 11514 1528 11534
rect 1548 11514 1557 11534
rect 1409 11508 1557 11514
rect 1409 11505 1473 11508
rect 1409 11504 1446 11505
rect 1465 11478 1473 11505
rect 1494 11505 1557 11508
rect 1615 11534 1753 11541
rect 1615 11514 1624 11534
rect 1644 11514 1753 11534
rect 1615 11505 1753 11514
rect 1494 11478 1501 11505
rect 1520 11504 1557 11505
rect 1616 11504 1653 11505
rect 1465 11453 1501 11478
rect 936 11451 977 11452
rect 816 11444 977 11451
rect 816 11424 946 11444
rect 966 11424 977 11444
rect 816 11422 977 11424
rect 766 11416 977 11422
rect 1044 11448 1403 11452
rect 1044 11443 1366 11448
rect 1044 11419 1157 11443
rect 1181 11424 1366 11443
rect 1390 11424 1403 11448
rect 1181 11419 1403 11424
rect 1044 11416 1403 11419
rect 1465 11416 1500 11453
rect 1568 11450 1668 11453
rect 1568 11446 1635 11450
rect 1568 11420 1580 11446
rect 1606 11424 1635 11446
rect 1661 11424 1668 11450
rect 1606 11420 1668 11424
rect 1568 11416 1668 11420
rect 766 11403 833 11416
rect 558 11380 614 11400
rect 558 11362 577 11380
rect 595 11362 614 11380
rect 558 11249 614 11362
rect 766 11382 780 11403
rect 816 11382 833 11403
rect 1044 11395 1075 11416
rect 1465 11395 1501 11416
rect 887 11394 924 11395
rect 766 11375 833 11382
rect 886 11385 924 11394
rect 558 11120 613 11249
rect 766 11223 831 11375
rect 886 11365 895 11385
rect 915 11365 924 11385
rect 886 11357 924 11365
rect 990 11389 1075 11395
rect 1100 11394 1137 11395
rect 990 11369 998 11389
rect 1018 11369 1075 11389
rect 990 11361 1075 11369
rect 1099 11385 1137 11394
rect 1099 11365 1108 11385
rect 1128 11365 1137 11385
rect 990 11360 1026 11361
rect 1099 11357 1137 11365
rect 1203 11389 1288 11395
rect 1308 11394 1345 11395
rect 1203 11369 1211 11389
rect 1231 11388 1288 11389
rect 1231 11369 1260 11388
rect 1203 11368 1260 11369
rect 1281 11368 1288 11388
rect 1203 11361 1288 11368
rect 1307 11385 1345 11394
rect 1307 11365 1316 11385
rect 1336 11365 1345 11385
rect 1203 11360 1239 11361
rect 1307 11357 1345 11365
rect 1411 11389 1555 11395
rect 1411 11369 1419 11389
rect 1439 11369 1527 11389
rect 1547 11369 1555 11389
rect 1411 11361 1555 11369
rect 1411 11360 1447 11361
rect 1519 11360 1555 11361
rect 1621 11394 1658 11395
rect 1621 11393 1659 11394
rect 1621 11385 1685 11393
rect 1621 11365 1630 11385
rect 1650 11371 1685 11385
rect 1705 11371 1708 11391
rect 1650 11366 1708 11371
rect 1650 11365 1685 11366
rect 887 11328 924 11357
rect 888 11326 924 11328
rect 1100 11326 1137 11357
rect 888 11304 1137 11326
rect 969 11298 1080 11304
rect 969 11290 1010 11298
rect 969 11270 977 11290
rect 996 11270 1010 11290
rect 969 11268 1010 11270
rect 1038 11290 1080 11298
rect 1038 11270 1054 11290
rect 1073 11270 1080 11290
rect 1038 11268 1080 11270
rect 969 11253 1080 11268
rect 1308 11258 1345 11357
rect 1621 11353 1685 11365
rect 971 11244 1075 11253
rect 759 11213 880 11223
rect 759 11211 828 11213
rect 759 11170 772 11211
rect 809 11172 828 11211
rect 865 11172 880 11213
rect 809 11170 880 11172
rect 759 11152 880 11170
rect 552 11108 613 11120
rect 1306 11108 1347 11258
rect 1725 11250 1752 11505
rect 1814 11495 1894 11506
rect 1814 11469 1831 11495
rect 1871 11469 1894 11495
rect 1814 11442 1894 11469
rect 1814 11416 1835 11442
rect 1875 11416 1894 11442
rect 1814 11397 1894 11416
rect 1814 11371 1838 11397
rect 1878 11371 1894 11397
rect 1814 11320 1894 11371
rect 552 11105 1347 11108
rect 1726 11119 1752 11250
rect 1816 11164 1886 11320
rect 1815 11148 1891 11164
rect 1726 11105 1754 11119
rect 552 11070 1754 11105
rect 1815 11111 1830 11148
rect 1874 11111 1891 11148
rect 1815 11091 1891 11111
rect 2929 11141 2999 12050
rect 3098 11485 3179 12198
rect 4003 12084 4039 12393
rect 3927 12055 4040 12084
rect 3927 11699 3958 12055
rect 3997 11800 4988 11825
rect 3997 11795 4057 11800
rect 3997 11774 4016 11795
rect 4036 11779 4057 11795
rect 4077 11779 4988 11800
rect 4036 11774 4988 11779
rect 3997 11766 4988 11774
rect 4002 11743 4108 11766
rect 4002 11740 4107 11743
rect 3851 11679 4244 11699
rect 4264 11679 4267 11699
rect 3851 11674 4267 11679
rect 3851 11673 4192 11674
rect 3508 11642 3618 11656
rect 3508 11639 3551 11642
rect 3508 11634 3512 11639
rect 3430 11612 3512 11634
rect 3541 11612 3551 11639
rect 3579 11615 3586 11642
rect 3615 11634 3618 11642
rect 3615 11615 3680 11634
rect 3579 11612 3680 11615
rect 3430 11610 3680 11612
rect 3430 11531 3467 11610
rect 3508 11597 3618 11610
rect 3582 11541 3613 11542
rect 3430 11511 3439 11531
rect 3459 11511 3467 11531
rect 3430 11501 3467 11511
rect 3526 11531 3613 11541
rect 3526 11511 3535 11531
rect 3555 11511 3613 11531
rect 3526 11502 3613 11511
rect 3526 11501 3563 11502
rect 3096 11449 3188 11485
rect 3582 11449 3613 11502
rect 3643 11531 3680 11610
rect 3795 11541 3826 11542
rect 3643 11511 3652 11531
rect 3672 11511 3680 11531
rect 3643 11501 3680 11511
rect 3739 11534 3826 11541
rect 3739 11531 3800 11534
rect 3739 11511 3748 11531
rect 3768 11514 3800 11531
rect 3821 11514 3826 11534
rect 3768 11511 3826 11514
rect 3739 11504 3826 11511
rect 3851 11531 3888 11673
rect 4154 11672 4191 11673
rect 4003 11541 4039 11542
rect 3851 11511 3860 11531
rect 3880 11511 3888 11531
rect 3739 11502 3795 11504
rect 3739 11501 3776 11502
rect 3851 11501 3888 11511
rect 3947 11531 4095 11541
rect 4195 11538 4291 11540
rect 3947 11511 3956 11531
rect 3976 11511 4066 11531
rect 4086 11511 4095 11531
rect 3947 11505 4095 11511
rect 3947 11502 4011 11505
rect 3947 11501 3984 11502
rect 4003 11475 4011 11502
rect 4032 11502 4095 11505
rect 4153 11531 4291 11538
rect 4153 11511 4162 11531
rect 4182 11511 4291 11531
rect 4153 11502 4291 11511
rect 4032 11475 4039 11502
rect 4058 11501 4095 11502
rect 4154 11501 4191 11502
rect 4003 11450 4039 11475
rect 3096 11448 3432 11449
rect 3474 11448 3515 11449
rect 3096 11441 3515 11448
rect 3096 11421 3484 11441
rect 3504 11421 3515 11441
rect 3096 11413 3515 11421
rect 3582 11445 3941 11449
rect 3582 11440 3904 11445
rect 3582 11416 3695 11440
rect 3719 11421 3904 11440
rect 3928 11421 3941 11445
rect 3719 11416 3941 11421
rect 3582 11413 3941 11416
rect 4003 11413 4038 11450
rect 4106 11447 4206 11450
rect 4106 11443 4173 11447
rect 4106 11417 4118 11443
rect 4144 11421 4173 11443
rect 4199 11421 4206 11447
rect 4144 11417 4206 11421
rect 4106 11413 4206 11417
rect 3096 11409 3432 11413
rect 2929 11091 3001 11141
rect 552 10995 613 11070
rect 971 11068 1075 11070
rect 1306 11068 1347 11070
rect 1815 11025 1825 11091
rect 1879 11025 1891 11091
rect 1815 11001 1891 11025
rect 554 10865 613 10995
rect 1467 10946 1539 10947
rect 1466 10938 1565 10946
rect 1466 10935 1518 10938
rect 1466 10900 1474 10935
rect 1499 10900 1518 10935
rect 1543 10927 1565 10938
rect 1543 10926 2410 10927
rect 1543 10900 2411 10926
rect 1466 10890 2411 10900
rect 1466 10888 1565 10890
rect 554 10847 576 10865
rect 594 10847 613 10865
rect 554 10825 613 10847
rect 821 10861 1353 10866
rect 821 10841 1707 10861
rect 1727 10841 1730 10861
rect 2366 10857 2411 10890
rect 821 10837 1730 10841
rect 821 10790 864 10837
rect 1314 10836 1730 10837
rect 2362 10837 2755 10857
rect 2775 10837 2778 10857
rect 1314 10835 1655 10836
rect 971 10804 1081 10818
rect 971 10801 1014 10804
rect 971 10796 975 10801
rect 809 10789 864 10790
rect 553 10766 864 10789
rect 553 10748 578 10766
rect 596 10754 864 10766
rect 893 10774 975 10796
rect 1004 10774 1014 10801
rect 1042 10777 1049 10804
rect 1078 10796 1081 10804
rect 1078 10777 1143 10796
rect 1042 10774 1143 10777
rect 893 10772 1143 10774
rect 596 10748 618 10754
rect 553 10609 618 10748
rect 893 10693 930 10772
rect 971 10759 1081 10772
rect 1045 10703 1076 10704
rect 893 10673 902 10693
rect 922 10673 930 10693
rect 553 10591 576 10609
rect 594 10591 618 10609
rect 553 10574 618 10591
rect 773 10655 841 10668
rect 893 10663 930 10673
rect 989 10693 1076 10703
rect 989 10673 998 10693
rect 1018 10673 1076 10693
rect 989 10664 1076 10673
rect 989 10663 1026 10664
rect 773 10613 780 10655
rect 829 10613 841 10655
rect 773 10610 841 10613
rect 1045 10611 1076 10664
rect 1106 10693 1143 10772
rect 1258 10703 1289 10704
rect 1106 10673 1115 10693
rect 1135 10673 1143 10693
rect 1106 10663 1143 10673
rect 1202 10696 1289 10703
rect 1202 10693 1263 10696
rect 1202 10673 1211 10693
rect 1231 10676 1263 10693
rect 1284 10676 1289 10696
rect 1231 10673 1289 10676
rect 1202 10666 1289 10673
rect 1314 10693 1351 10835
rect 1617 10834 1654 10835
rect 2362 10832 2778 10837
rect 2362 10831 2703 10832
rect 2019 10800 2129 10814
rect 2019 10797 2062 10800
rect 2019 10792 2023 10797
rect 1941 10770 2023 10792
rect 2052 10770 2062 10797
rect 2090 10773 2097 10800
rect 2126 10792 2129 10800
rect 2126 10773 2191 10792
rect 2090 10770 2191 10773
rect 1941 10768 2191 10770
rect 1466 10703 1502 10704
rect 1314 10673 1323 10693
rect 1343 10673 1351 10693
rect 1202 10664 1258 10666
rect 1202 10663 1239 10664
rect 1314 10663 1351 10673
rect 1410 10693 1558 10703
rect 1658 10700 1754 10702
rect 1410 10673 1419 10693
rect 1439 10673 1529 10693
rect 1549 10673 1558 10693
rect 1410 10667 1558 10673
rect 1410 10664 1474 10667
rect 1410 10663 1447 10664
rect 1466 10637 1474 10664
rect 1495 10664 1558 10667
rect 1616 10693 1754 10700
rect 1616 10673 1625 10693
rect 1645 10673 1754 10693
rect 1616 10664 1754 10673
rect 1941 10689 1978 10768
rect 2019 10755 2129 10768
rect 2093 10699 2124 10700
rect 1941 10669 1950 10689
rect 1970 10669 1978 10689
rect 1495 10637 1502 10664
rect 1521 10663 1558 10664
rect 1617 10663 1654 10664
rect 1466 10612 1502 10637
rect 937 10610 978 10611
rect 773 10603 978 10610
rect 773 10592 947 10603
rect 773 10559 781 10592
rect 774 10550 781 10559
rect 830 10583 947 10592
rect 967 10583 978 10603
rect 830 10575 978 10583
rect 1045 10607 1404 10611
rect 1045 10602 1367 10607
rect 1045 10578 1158 10602
rect 1182 10583 1367 10602
rect 1391 10583 1404 10607
rect 1182 10578 1404 10583
rect 1045 10575 1404 10578
rect 1466 10575 1501 10612
rect 1569 10609 1669 10612
rect 1569 10605 1636 10609
rect 1569 10579 1581 10605
rect 1607 10583 1636 10605
rect 1662 10583 1669 10609
rect 1607 10579 1669 10583
rect 1569 10575 1669 10579
rect 830 10559 841 10575
rect 830 10550 838 10559
rect 1045 10554 1076 10575
rect 1466 10554 1502 10575
rect 888 10553 925 10554
rect 553 10510 618 10529
rect 553 10492 578 10510
rect 596 10492 618 10510
rect 553 10291 618 10492
rect 774 10366 838 10550
rect 887 10544 925 10553
rect 887 10524 896 10544
rect 916 10524 925 10544
rect 887 10516 925 10524
rect 991 10548 1076 10554
rect 1101 10553 1138 10554
rect 991 10528 999 10548
rect 1019 10528 1076 10548
rect 991 10520 1076 10528
rect 1100 10544 1138 10553
rect 1100 10524 1109 10544
rect 1129 10524 1138 10544
rect 991 10519 1027 10520
rect 1100 10516 1138 10524
rect 1204 10548 1289 10554
rect 1309 10553 1346 10554
rect 1204 10528 1212 10548
rect 1232 10547 1289 10548
rect 1232 10528 1261 10547
rect 1204 10527 1261 10528
rect 1282 10527 1289 10547
rect 1204 10520 1289 10527
rect 1308 10544 1346 10553
rect 1308 10524 1317 10544
rect 1337 10524 1346 10544
rect 1204 10519 1240 10520
rect 1308 10516 1346 10524
rect 1412 10548 1556 10554
rect 1412 10528 1420 10548
rect 1440 10528 1528 10548
rect 1548 10528 1556 10548
rect 1412 10520 1556 10528
rect 1412 10519 1448 10520
rect 1520 10519 1556 10520
rect 1622 10553 1659 10554
rect 1622 10552 1660 10553
rect 1622 10544 1686 10552
rect 1622 10524 1631 10544
rect 1651 10530 1686 10544
rect 1706 10530 1709 10550
rect 1651 10525 1709 10530
rect 1651 10524 1686 10525
rect 888 10487 925 10516
rect 889 10485 925 10487
rect 1101 10485 1138 10516
rect 889 10463 1138 10485
rect 970 10457 1081 10463
rect 970 10449 1011 10457
rect 970 10429 978 10449
rect 997 10429 1011 10449
rect 970 10427 1011 10429
rect 1039 10449 1081 10457
rect 1039 10429 1055 10449
rect 1074 10429 1081 10449
rect 1039 10427 1081 10429
rect 970 10412 1081 10427
rect 774 10356 842 10366
rect 774 10323 791 10356
rect 831 10323 842 10356
rect 774 10311 842 10323
rect 774 10309 838 10311
rect 1309 10292 1346 10516
rect 1622 10512 1686 10524
rect 1726 10294 1753 10664
rect 1941 10659 1978 10669
rect 2037 10689 2124 10699
rect 2037 10669 2046 10689
rect 2066 10669 2124 10689
rect 2037 10660 2124 10669
rect 2037 10659 2074 10660
rect 1817 10646 1887 10651
rect 1812 10640 1887 10646
rect 1812 10607 1820 10640
rect 1873 10607 1887 10640
rect 2093 10607 2124 10660
rect 2154 10689 2191 10768
rect 2306 10699 2337 10700
rect 2154 10669 2163 10689
rect 2183 10669 2191 10689
rect 2154 10659 2191 10669
rect 2250 10692 2337 10699
rect 2250 10689 2311 10692
rect 2250 10669 2259 10689
rect 2279 10672 2311 10689
rect 2332 10672 2337 10692
rect 2279 10669 2337 10672
rect 2250 10662 2337 10669
rect 2362 10689 2399 10831
rect 2665 10830 2702 10831
rect 2514 10699 2550 10700
rect 2362 10669 2371 10689
rect 2391 10669 2399 10689
rect 2250 10660 2306 10662
rect 2250 10659 2287 10660
rect 2362 10659 2399 10669
rect 2458 10689 2606 10699
rect 2706 10696 2802 10698
rect 2458 10669 2467 10689
rect 2487 10669 2577 10689
rect 2597 10669 2606 10689
rect 2458 10663 2606 10669
rect 2458 10660 2522 10663
rect 2458 10659 2495 10660
rect 2514 10633 2522 10660
rect 2543 10660 2606 10663
rect 2664 10689 2802 10696
rect 2664 10669 2673 10689
rect 2693 10669 2802 10689
rect 2664 10660 2802 10669
rect 2543 10633 2550 10660
rect 2569 10659 2606 10660
rect 2665 10659 2702 10660
rect 2514 10608 2550 10633
rect 1812 10606 1895 10607
rect 1985 10606 2026 10607
rect 1812 10599 2026 10606
rect 1812 10582 1995 10599
rect 1812 10549 1825 10582
rect 1878 10579 1995 10582
rect 2015 10579 2026 10599
rect 1878 10571 2026 10579
rect 2093 10603 2452 10607
rect 2093 10598 2415 10603
rect 2093 10574 2206 10598
rect 2230 10579 2415 10598
rect 2439 10579 2452 10603
rect 2230 10574 2452 10579
rect 2093 10571 2452 10574
rect 2514 10571 2549 10608
rect 2617 10605 2717 10608
rect 2617 10601 2684 10605
rect 2617 10575 2629 10601
rect 2655 10579 2684 10601
rect 2710 10579 2717 10605
rect 2655 10575 2717 10579
rect 2617 10571 2717 10575
rect 1878 10549 1895 10571
rect 2093 10550 2124 10571
rect 2514 10550 2550 10571
rect 1936 10549 1973 10550
rect 1812 10535 1895 10549
rect 1585 10292 1753 10294
rect 1309 10291 1753 10292
rect 553 10261 1753 10291
rect 1823 10325 1895 10535
rect 1935 10540 1973 10549
rect 1935 10520 1944 10540
rect 1964 10520 1973 10540
rect 1935 10512 1973 10520
rect 2039 10544 2124 10550
rect 2149 10549 2186 10550
rect 2039 10524 2047 10544
rect 2067 10524 2124 10544
rect 2039 10516 2124 10524
rect 2148 10540 2186 10549
rect 2148 10520 2157 10540
rect 2177 10520 2186 10540
rect 2039 10515 2075 10516
rect 2148 10512 2186 10520
rect 2252 10544 2337 10550
rect 2357 10549 2394 10550
rect 2252 10524 2260 10544
rect 2280 10543 2337 10544
rect 2280 10524 2309 10543
rect 2252 10523 2309 10524
rect 2330 10523 2337 10543
rect 2252 10516 2337 10523
rect 2356 10540 2394 10549
rect 2356 10520 2365 10540
rect 2385 10520 2394 10540
rect 2252 10515 2288 10516
rect 2356 10512 2394 10520
rect 2460 10544 2604 10550
rect 2460 10524 2468 10544
rect 2488 10524 2576 10544
rect 2596 10524 2604 10544
rect 2460 10516 2604 10524
rect 2460 10515 2496 10516
rect 2568 10515 2604 10516
rect 2670 10549 2707 10550
rect 2670 10548 2708 10549
rect 2670 10540 2734 10548
rect 2670 10520 2679 10540
rect 2699 10526 2734 10540
rect 2754 10526 2757 10546
rect 2699 10521 2757 10526
rect 2699 10520 2734 10521
rect 1936 10483 1973 10512
rect 1937 10481 1973 10483
rect 2149 10481 2186 10512
rect 1937 10459 2186 10481
rect 2018 10453 2129 10459
rect 2018 10445 2059 10453
rect 2018 10425 2026 10445
rect 2045 10425 2059 10445
rect 2018 10423 2059 10425
rect 2087 10445 2129 10453
rect 2087 10425 2103 10445
rect 2122 10425 2129 10445
rect 2087 10423 2129 10425
rect 2018 10408 2129 10423
rect 1823 10286 1842 10325
rect 1887 10286 1895 10325
rect 1823 10269 1895 10286
rect 2357 10313 2394 10512
rect 2670 10508 2734 10520
rect 2357 10307 2398 10313
rect 2774 10309 2801 10660
rect 2930 10612 3001 11091
rect 2930 10528 2999 10612
rect 2633 10307 2801 10309
rect 2357 10281 2801 10307
rect 553 10214 618 10261
rect 553 10196 576 10214
rect 594 10196 618 10214
rect 1466 10241 1501 10243
rect 1466 10239 1570 10241
rect 2359 10239 2398 10281
rect 2633 10280 2801 10281
rect 1466 10232 2400 10239
rect 1466 10231 1517 10232
rect 1466 10211 1469 10231
rect 1494 10212 1517 10231
rect 1549 10212 2400 10232
rect 1494 10211 2400 10212
rect 1466 10204 2400 10211
rect 1739 10203 2400 10204
rect 553 10175 618 10196
rect 830 10186 870 10189
rect 830 10182 1733 10186
rect 830 10162 1707 10182
rect 1727 10162 1733 10182
rect 830 10159 1733 10162
rect 554 10115 619 10135
rect 554 10097 578 10115
rect 596 10097 619 10115
rect 554 10070 619 10097
rect 830 10070 870 10159
rect 1314 10157 1730 10159
rect 1314 10156 1655 10157
rect 971 10125 1081 10139
rect 971 10122 1014 10125
rect 971 10117 975 10122
rect 553 10035 870 10070
rect 893 10095 975 10117
rect 1004 10095 1014 10122
rect 1042 10098 1049 10125
rect 1078 10117 1081 10125
rect 1078 10098 1143 10117
rect 1042 10095 1143 10098
rect 893 10093 1143 10095
rect 554 9959 619 10035
rect 893 10014 930 10093
rect 971 10080 1081 10093
rect 1045 10024 1076 10025
rect 893 9994 902 10014
rect 922 9994 930 10014
rect 893 9984 930 9994
rect 989 10014 1076 10024
rect 989 9994 998 10014
rect 1018 9994 1076 10014
rect 989 9985 1076 9994
rect 989 9984 1026 9985
rect 554 9941 576 9959
rect 594 9941 619 9959
rect 554 9920 619 9941
rect 767 9939 832 9948
rect 767 9902 777 9939
rect 817 9931 832 9939
rect 1045 9932 1076 9985
rect 1106 10014 1143 10093
rect 1258 10024 1289 10025
rect 1106 9994 1115 10014
rect 1135 9994 1143 10014
rect 1106 9984 1143 9994
rect 1202 10017 1289 10024
rect 1202 10014 1263 10017
rect 1202 9994 1211 10014
rect 1231 9997 1263 10014
rect 1284 9997 1289 10017
rect 1231 9994 1289 9997
rect 1202 9987 1289 9994
rect 1314 10014 1351 10156
rect 1617 10155 1654 10156
rect 1466 10024 1502 10025
rect 1314 9994 1323 10014
rect 1343 9994 1351 10014
rect 1202 9985 1258 9987
rect 1202 9984 1239 9985
rect 1314 9984 1351 9994
rect 1410 10014 1558 10024
rect 1658 10021 1754 10023
rect 1410 9994 1419 10014
rect 1439 9994 1529 10014
rect 1549 9994 1558 10014
rect 1410 9988 1558 9994
rect 1410 9985 1474 9988
rect 1410 9984 1447 9985
rect 1466 9958 1474 9985
rect 1495 9985 1558 9988
rect 1616 10014 1754 10021
rect 1616 9994 1625 10014
rect 1645 9994 1754 10014
rect 2934 10012 2996 10528
rect 1616 9985 1754 9994
rect 1495 9958 1502 9985
rect 1521 9984 1558 9985
rect 1617 9984 1654 9985
rect 1466 9933 1502 9958
rect 937 9931 978 9932
rect 817 9924 978 9931
rect 817 9904 947 9924
rect 967 9904 978 9924
rect 817 9902 978 9904
rect 767 9896 978 9902
rect 1045 9928 1404 9932
rect 1045 9923 1367 9928
rect 1045 9899 1158 9923
rect 1182 9904 1367 9923
rect 1391 9904 1404 9928
rect 1182 9899 1404 9904
rect 1045 9896 1404 9899
rect 1466 9896 1501 9933
rect 1569 9930 1669 9933
rect 1569 9926 1636 9930
rect 1569 9900 1581 9926
rect 1607 9904 1636 9926
rect 1662 9904 1669 9930
rect 1607 9900 1669 9904
rect 1569 9896 1669 9900
rect 767 9883 834 9896
rect 559 9860 615 9880
rect 559 9842 578 9860
rect 596 9842 615 9860
rect 559 9729 615 9842
rect 767 9862 781 9883
rect 817 9862 834 9883
rect 1045 9875 1076 9896
rect 1466 9875 1502 9896
rect 888 9874 925 9875
rect 767 9855 834 9862
rect 887 9865 925 9874
rect 559 9591 614 9729
rect 767 9703 832 9855
rect 887 9845 896 9865
rect 916 9845 925 9865
rect 887 9837 925 9845
rect 991 9869 1076 9875
rect 1101 9874 1138 9875
rect 991 9849 999 9869
rect 1019 9849 1076 9869
rect 991 9841 1076 9849
rect 1100 9865 1138 9874
rect 1100 9845 1109 9865
rect 1129 9845 1138 9865
rect 991 9840 1027 9841
rect 1100 9837 1138 9845
rect 1204 9869 1289 9875
rect 1309 9874 1346 9875
rect 1204 9849 1212 9869
rect 1232 9868 1289 9869
rect 1232 9849 1261 9868
rect 1204 9848 1261 9849
rect 1282 9848 1289 9868
rect 1204 9841 1289 9848
rect 1308 9865 1346 9874
rect 1308 9845 1317 9865
rect 1337 9845 1346 9865
rect 1204 9840 1240 9841
rect 1308 9837 1346 9845
rect 1412 9869 1556 9875
rect 1412 9849 1420 9869
rect 1440 9849 1528 9869
rect 1548 9849 1556 9869
rect 1412 9841 1556 9849
rect 1412 9840 1448 9841
rect 1520 9840 1556 9841
rect 1622 9874 1659 9875
rect 1622 9873 1660 9874
rect 1622 9865 1686 9873
rect 1622 9845 1631 9865
rect 1651 9851 1686 9865
rect 1706 9851 1709 9871
rect 1651 9846 1709 9851
rect 1651 9845 1686 9846
rect 888 9808 925 9837
rect 889 9806 925 9808
rect 1101 9806 1138 9837
rect 889 9784 1138 9806
rect 970 9778 1081 9784
rect 970 9770 1011 9778
rect 970 9750 978 9770
rect 997 9750 1011 9770
rect 970 9748 1011 9750
rect 1039 9770 1081 9778
rect 1039 9750 1055 9770
rect 1074 9750 1081 9770
rect 1039 9748 1081 9750
rect 970 9735 1081 9748
rect 1309 9738 1346 9837
rect 1622 9833 1686 9845
rect 760 9693 881 9703
rect 760 9691 829 9693
rect 760 9650 773 9691
rect 810 9652 829 9691
rect 866 9652 881 9693
rect 810 9650 881 9652
rect 760 9632 881 9650
rect 552 9588 616 9591
rect 972 9588 1076 9594
rect 1307 9588 1348 9738
rect 1726 9730 1753 9985
rect 1815 9975 1895 9986
rect 1815 9949 1832 9975
rect 1872 9949 1895 9975
rect 1815 9922 1895 9949
rect 1815 9896 1836 9922
rect 1876 9896 1895 9922
rect 1815 9877 1895 9896
rect 1815 9851 1839 9877
rect 1879 9851 1895 9877
rect 1815 9800 1895 9851
rect 2918 9977 2996 10012
rect 2918 9915 3000 9977
rect 2918 9892 2946 9915
rect 2972 9892 3000 9915
rect 2918 9872 3000 9892
rect 552 9585 1348 9588
rect 1727 9599 1753 9730
rect 1727 9585 1755 9599
rect 552 9550 1755 9585
rect 1817 9592 1887 9800
rect 552 9489 616 9550
rect 972 9548 1076 9550
rect 1307 9548 1348 9550
rect 1817 9547 1838 9592
rect 1818 9526 1838 9547
rect 1868 9547 1887 9592
rect 1868 9526 1885 9547
rect 1818 9507 1885 9526
rect 1467 9499 1539 9500
rect 1466 9491 1565 9499
rect 554 9418 613 9489
rect 1466 9488 1518 9491
rect 1466 9453 1474 9488
rect 1499 9453 1518 9488
rect 1543 9480 1565 9491
rect 1543 9479 2410 9480
rect 1543 9453 2411 9479
rect 1466 9443 2411 9453
rect 1466 9441 1565 9443
rect 554 9400 576 9418
rect 594 9400 613 9418
rect 554 9378 613 9400
rect 821 9414 1353 9419
rect 821 9394 1707 9414
rect 1727 9394 1730 9414
rect 2366 9410 2411 9443
rect 821 9390 1730 9394
rect 821 9343 864 9390
rect 1314 9389 1730 9390
rect 2362 9390 2755 9410
rect 2775 9390 2778 9410
rect 1314 9388 1655 9389
rect 971 9357 1081 9371
rect 971 9354 1014 9357
rect 971 9349 975 9354
rect 809 9342 864 9343
rect 553 9319 864 9342
rect 553 9301 578 9319
rect 596 9307 864 9319
rect 893 9327 975 9349
rect 1004 9327 1014 9354
rect 1042 9330 1049 9357
rect 1078 9349 1081 9357
rect 1078 9330 1143 9349
rect 1042 9327 1143 9330
rect 893 9325 1143 9327
rect 596 9301 618 9307
rect 553 9162 618 9301
rect 893 9246 930 9325
rect 971 9312 1081 9325
rect 1045 9256 1076 9257
rect 893 9226 902 9246
rect 922 9226 930 9246
rect 553 9144 576 9162
rect 594 9144 618 9162
rect 553 9127 618 9144
rect 773 9208 841 9221
rect 893 9216 930 9226
rect 989 9246 1076 9256
rect 989 9226 998 9246
rect 1018 9226 1076 9246
rect 989 9217 1076 9226
rect 989 9216 1026 9217
rect 773 9166 780 9208
rect 829 9166 841 9208
rect 773 9163 841 9166
rect 1045 9164 1076 9217
rect 1106 9246 1143 9325
rect 1258 9256 1289 9257
rect 1106 9226 1115 9246
rect 1135 9226 1143 9246
rect 1106 9216 1143 9226
rect 1202 9249 1289 9256
rect 1202 9246 1263 9249
rect 1202 9226 1211 9246
rect 1231 9229 1263 9246
rect 1284 9229 1289 9249
rect 1231 9226 1289 9229
rect 1202 9219 1289 9226
rect 1314 9246 1351 9388
rect 1617 9387 1654 9388
rect 2362 9385 2778 9390
rect 2362 9384 2703 9385
rect 2019 9353 2129 9367
rect 2019 9350 2062 9353
rect 2019 9345 2023 9350
rect 1941 9323 2023 9345
rect 2052 9323 2062 9350
rect 2090 9326 2097 9353
rect 2126 9345 2129 9353
rect 2126 9326 2191 9345
rect 2090 9323 2191 9326
rect 1941 9321 2191 9323
rect 1466 9256 1502 9257
rect 1314 9226 1323 9246
rect 1343 9226 1351 9246
rect 1202 9217 1258 9219
rect 1202 9216 1239 9217
rect 1314 9216 1351 9226
rect 1410 9246 1558 9256
rect 1658 9253 1754 9255
rect 1410 9226 1419 9246
rect 1439 9226 1529 9246
rect 1549 9226 1558 9246
rect 1410 9220 1558 9226
rect 1410 9217 1474 9220
rect 1410 9216 1447 9217
rect 1466 9190 1474 9217
rect 1495 9217 1558 9220
rect 1616 9246 1754 9253
rect 1616 9226 1625 9246
rect 1645 9226 1754 9246
rect 1616 9217 1754 9226
rect 1941 9242 1978 9321
rect 2019 9308 2129 9321
rect 2093 9252 2124 9253
rect 1941 9222 1950 9242
rect 1970 9222 1978 9242
rect 1495 9190 1502 9217
rect 1521 9216 1558 9217
rect 1617 9216 1654 9217
rect 1466 9165 1502 9190
rect 937 9163 978 9164
rect 773 9156 978 9163
rect 773 9145 947 9156
rect 773 9112 781 9145
rect 774 9103 781 9112
rect 830 9136 947 9145
rect 967 9136 978 9156
rect 830 9128 978 9136
rect 1045 9160 1404 9164
rect 1045 9155 1367 9160
rect 1045 9131 1158 9155
rect 1182 9136 1367 9155
rect 1391 9136 1404 9160
rect 1182 9131 1404 9136
rect 1045 9128 1404 9131
rect 1466 9128 1501 9165
rect 1569 9162 1669 9165
rect 1569 9158 1636 9162
rect 1569 9132 1581 9158
rect 1607 9136 1636 9158
rect 1662 9136 1669 9162
rect 1607 9132 1669 9136
rect 1569 9128 1669 9132
rect 830 9112 841 9128
rect 830 9103 838 9112
rect 1045 9107 1076 9128
rect 1466 9107 1502 9128
rect 888 9106 925 9107
rect 553 9063 618 9082
rect 553 9045 578 9063
rect 596 9045 618 9063
rect 553 8844 618 9045
rect 774 8919 838 9103
rect 887 9097 925 9106
rect 887 9077 896 9097
rect 916 9077 925 9097
rect 887 9069 925 9077
rect 991 9101 1076 9107
rect 1101 9106 1138 9107
rect 991 9081 999 9101
rect 1019 9081 1076 9101
rect 991 9073 1076 9081
rect 1100 9097 1138 9106
rect 1100 9077 1109 9097
rect 1129 9077 1138 9097
rect 991 9072 1027 9073
rect 1100 9069 1138 9077
rect 1204 9101 1289 9107
rect 1309 9106 1346 9107
rect 1204 9081 1212 9101
rect 1232 9100 1289 9101
rect 1232 9081 1261 9100
rect 1204 9080 1261 9081
rect 1282 9080 1289 9100
rect 1204 9073 1289 9080
rect 1308 9097 1346 9106
rect 1308 9077 1317 9097
rect 1337 9077 1346 9097
rect 1204 9072 1240 9073
rect 1308 9069 1346 9077
rect 1412 9101 1556 9107
rect 1412 9081 1420 9101
rect 1440 9081 1528 9101
rect 1548 9081 1556 9101
rect 1412 9073 1556 9081
rect 1412 9072 1448 9073
rect 1520 9072 1556 9073
rect 1622 9106 1659 9107
rect 1622 9105 1660 9106
rect 1622 9097 1686 9105
rect 1622 9077 1631 9097
rect 1651 9083 1686 9097
rect 1706 9083 1709 9103
rect 1651 9078 1709 9083
rect 1651 9077 1686 9078
rect 888 9040 925 9069
rect 889 9038 925 9040
rect 1101 9038 1138 9069
rect 889 9016 1138 9038
rect 970 9010 1081 9016
rect 970 9002 1011 9010
rect 970 8982 978 9002
rect 997 8982 1011 9002
rect 970 8980 1011 8982
rect 1039 9002 1081 9010
rect 1039 8982 1055 9002
rect 1074 8982 1081 9002
rect 1039 8980 1081 8982
rect 970 8965 1081 8980
rect 774 8909 842 8919
rect 774 8876 791 8909
rect 831 8876 842 8909
rect 774 8864 842 8876
rect 774 8862 838 8864
rect 1309 8845 1346 9069
rect 1622 9065 1686 9077
rect 1726 8847 1753 9217
rect 1941 9212 1978 9222
rect 2037 9242 2124 9252
rect 2037 9222 2046 9242
rect 2066 9222 2124 9242
rect 2037 9213 2124 9222
rect 2037 9212 2074 9213
rect 1817 9199 1887 9204
rect 1812 9193 1887 9199
rect 1812 9160 1820 9193
rect 1873 9160 1887 9193
rect 2093 9160 2124 9213
rect 2154 9242 2191 9321
rect 2306 9252 2337 9253
rect 2154 9222 2163 9242
rect 2183 9222 2191 9242
rect 2154 9212 2191 9222
rect 2250 9245 2337 9252
rect 2250 9242 2311 9245
rect 2250 9222 2259 9242
rect 2279 9225 2311 9242
rect 2332 9225 2337 9245
rect 2279 9222 2337 9225
rect 2250 9215 2337 9222
rect 2362 9242 2399 9384
rect 2665 9383 2702 9384
rect 2514 9252 2550 9253
rect 2362 9222 2371 9242
rect 2391 9222 2399 9242
rect 2250 9213 2306 9215
rect 2250 9212 2287 9213
rect 2362 9212 2399 9222
rect 2458 9242 2606 9252
rect 2706 9249 2802 9251
rect 2458 9222 2467 9242
rect 2487 9222 2577 9242
rect 2597 9222 2606 9242
rect 2458 9216 2606 9222
rect 2458 9213 2522 9216
rect 2458 9212 2495 9213
rect 2514 9186 2522 9213
rect 2543 9213 2606 9216
rect 2664 9242 2802 9249
rect 2664 9222 2673 9242
rect 2693 9222 2802 9242
rect 2664 9213 2802 9222
rect 2543 9186 2550 9213
rect 2569 9212 2606 9213
rect 2665 9212 2702 9213
rect 2514 9161 2550 9186
rect 1812 9159 1895 9160
rect 1985 9159 2026 9160
rect 1812 9152 2026 9159
rect 1812 9135 1995 9152
rect 1812 9102 1825 9135
rect 1878 9132 1995 9135
rect 2015 9132 2026 9152
rect 1878 9124 2026 9132
rect 2093 9156 2452 9160
rect 2093 9151 2415 9156
rect 2093 9127 2206 9151
rect 2230 9132 2415 9151
rect 2439 9132 2452 9156
rect 2230 9127 2452 9132
rect 2093 9124 2452 9127
rect 2514 9124 2549 9161
rect 2617 9158 2717 9161
rect 2617 9154 2684 9158
rect 2617 9128 2629 9154
rect 2655 9132 2684 9154
rect 2710 9132 2717 9158
rect 2655 9128 2717 9132
rect 2617 9124 2717 9128
rect 1878 9102 1895 9124
rect 2093 9103 2124 9124
rect 2514 9103 2550 9124
rect 1936 9102 1973 9103
rect 1812 9088 1895 9102
rect 1585 8845 1753 8847
rect 1309 8844 1753 8845
rect 553 8814 1753 8844
rect 1823 8878 1895 9088
rect 1935 9093 1973 9102
rect 1935 9073 1944 9093
rect 1964 9073 1973 9093
rect 1935 9065 1973 9073
rect 2039 9097 2124 9103
rect 2149 9102 2186 9103
rect 2039 9077 2047 9097
rect 2067 9077 2124 9097
rect 2039 9069 2124 9077
rect 2148 9093 2186 9102
rect 2148 9073 2157 9093
rect 2177 9073 2186 9093
rect 2039 9068 2075 9069
rect 2148 9065 2186 9073
rect 2252 9097 2337 9103
rect 2357 9102 2394 9103
rect 2252 9077 2260 9097
rect 2280 9096 2337 9097
rect 2280 9077 2309 9096
rect 2252 9076 2309 9077
rect 2330 9076 2337 9096
rect 2252 9069 2337 9076
rect 2356 9093 2394 9102
rect 2356 9073 2365 9093
rect 2385 9073 2394 9093
rect 2252 9068 2288 9069
rect 2356 9065 2394 9073
rect 2460 9097 2604 9103
rect 2460 9077 2468 9097
rect 2488 9077 2576 9097
rect 2596 9077 2604 9097
rect 2460 9069 2604 9077
rect 2460 9068 2496 9069
rect 2568 9068 2604 9069
rect 2670 9102 2707 9103
rect 2670 9101 2708 9102
rect 2670 9093 2734 9101
rect 2670 9073 2679 9093
rect 2699 9079 2734 9093
rect 2754 9079 2757 9099
rect 2699 9074 2757 9079
rect 2699 9073 2734 9074
rect 1936 9036 1973 9065
rect 1937 9034 1973 9036
rect 2149 9034 2186 9065
rect 1937 9012 2186 9034
rect 2018 9006 2129 9012
rect 2018 8998 2059 9006
rect 2018 8978 2026 8998
rect 2045 8978 2059 8998
rect 2018 8976 2059 8978
rect 2087 8998 2129 9006
rect 2087 8978 2103 8998
rect 2122 8978 2129 8998
rect 2087 8976 2129 8978
rect 2018 8961 2129 8976
rect 1823 8839 1842 8878
rect 1887 8839 1895 8878
rect 1823 8822 1895 8839
rect 2357 8866 2394 9065
rect 2670 9061 2734 9073
rect 2357 8860 2398 8866
rect 2774 8862 2801 9213
rect 2633 8860 2801 8862
rect 2357 8834 2801 8860
rect 553 8767 618 8814
rect 553 8749 576 8767
rect 594 8749 618 8767
rect 1466 8794 1501 8796
rect 1466 8792 1570 8794
rect 2359 8792 2398 8834
rect 2633 8833 2801 8834
rect 1466 8785 2400 8792
rect 1466 8784 1517 8785
rect 1466 8764 1469 8784
rect 1494 8765 1517 8784
rect 1549 8765 2400 8785
rect 1494 8764 2400 8765
rect 1466 8757 2400 8764
rect 1739 8756 2400 8757
rect 553 8728 618 8749
rect 830 8739 870 8742
rect 830 8735 1733 8739
rect 830 8715 1707 8735
rect 1727 8715 1733 8735
rect 830 8712 1733 8715
rect 554 8668 619 8688
rect 554 8650 578 8668
rect 596 8650 619 8668
rect 554 8623 619 8650
rect 830 8623 870 8712
rect 1314 8710 1730 8712
rect 1314 8709 1655 8710
rect 971 8678 1081 8692
rect 971 8675 1014 8678
rect 971 8670 975 8675
rect 553 8588 870 8623
rect 893 8648 975 8670
rect 1004 8648 1014 8675
rect 1042 8651 1049 8678
rect 1078 8670 1081 8678
rect 1078 8651 1143 8670
rect 1042 8648 1143 8651
rect 893 8646 1143 8648
rect 554 8512 619 8588
rect 893 8567 930 8646
rect 971 8633 1081 8646
rect 1045 8577 1076 8578
rect 893 8547 902 8567
rect 922 8547 930 8567
rect 893 8537 930 8547
rect 989 8567 1076 8577
rect 989 8547 998 8567
rect 1018 8547 1076 8567
rect 989 8538 1076 8547
rect 989 8537 1026 8538
rect 554 8494 576 8512
rect 594 8494 619 8512
rect 554 8473 619 8494
rect 767 8492 832 8501
rect 767 8455 777 8492
rect 817 8484 832 8492
rect 1045 8485 1076 8538
rect 1106 8567 1143 8646
rect 1258 8577 1289 8578
rect 1106 8547 1115 8567
rect 1135 8547 1143 8567
rect 1106 8537 1143 8547
rect 1202 8570 1289 8577
rect 1202 8567 1263 8570
rect 1202 8547 1211 8567
rect 1231 8550 1263 8567
rect 1284 8550 1289 8570
rect 1231 8547 1289 8550
rect 1202 8540 1289 8547
rect 1314 8567 1351 8709
rect 1617 8708 1654 8709
rect 1466 8577 1502 8578
rect 1314 8547 1323 8567
rect 1343 8547 1351 8567
rect 1202 8538 1258 8540
rect 1202 8537 1239 8538
rect 1314 8537 1351 8547
rect 1410 8567 1558 8577
rect 1658 8574 1754 8576
rect 1410 8547 1419 8567
rect 1439 8547 1529 8567
rect 1549 8547 1558 8567
rect 1410 8541 1558 8547
rect 1410 8538 1474 8541
rect 1410 8537 1447 8538
rect 1466 8511 1474 8538
rect 1495 8538 1558 8541
rect 1616 8567 1754 8574
rect 1616 8547 1625 8567
rect 1645 8547 1754 8567
rect 1616 8538 1754 8547
rect 1495 8511 1502 8538
rect 1521 8537 1558 8538
rect 1617 8537 1654 8538
rect 1466 8486 1502 8511
rect 937 8484 978 8485
rect 817 8477 978 8484
rect 817 8457 947 8477
rect 967 8457 978 8477
rect 817 8455 978 8457
rect 767 8449 978 8455
rect 1045 8481 1404 8485
rect 1045 8476 1367 8481
rect 1045 8452 1158 8476
rect 1182 8457 1367 8476
rect 1391 8457 1404 8481
rect 1182 8452 1404 8457
rect 1045 8449 1404 8452
rect 1466 8449 1501 8486
rect 1569 8483 1669 8486
rect 1569 8479 1636 8483
rect 1569 8453 1581 8479
rect 1607 8457 1636 8479
rect 1662 8457 1669 8483
rect 1607 8453 1669 8457
rect 1569 8449 1669 8453
rect 767 8436 834 8449
rect 559 8413 615 8433
rect 559 8395 578 8413
rect 596 8395 615 8413
rect 559 8282 615 8395
rect 767 8415 781 8436
rect 817 8415 834 8436
rect 1045 8428 1076 8449
rect 1466 8428 1502 8449
rect 888 8427 925 8428
rect 767 8408 834 8415
rect 887 8418 925 8427
rect 559 8175 614 8282
rect 767 8256 832 8408
rect 887 8398 896 8418
rect 916 8398 925 8418
rect 887 8390 925 8398
rect 991 8422 1076 8428
rect 1101 8427 1138 8428
rect 991 8402 999 8422
rect 1019 8402 1076 8422
rect 991 8394 1076 8402
rect 1100 8418 1138 8427
rect 1100 8398 1109 8418
rect 1129 8398 1138 8418
rect 991 8393 1027 8394
rect 1100 8390 1138 8398
rect 1204 8422 1289 8428
rect 1309 8427 1346 8428
rect 1204 8402 1212 8422
rect 1232 8421 1289 8422
rect 1232 8402 1261 8421
rect 1204 8401 1261 8402
rect 1282 8401 1289 8421
rect 1204 8394 1289 8401
rect 1308 8418 1346 8427
rect 1308 8398 1317 8418
rect 1337 8398 1346 8418
rect 1204 8393 1240 8394
rect 1308 8390 1346 8398
rect 1412 8422 1556 8428
rect 1412 8402 1420 8422
rect 1440 8402 1528 8422
rect 1548 8402 1556 8422
rect 1412 8394 1556 8402
rect 1412 8393 1448 8394
rect 1520 8393 1556 8394
rect 1622 8427 1659 8428
rect 1622 8426 1660 8427
rect 1622 8418 1686 8426
rect 1622 8398 1631 8418
rect 1651 8404 1686 8418
rect 1706 8404 1709 8424
rect 1651 8399 1709 8404
rect 1651 8398 1686 8399
rect 888 8361 925 8390
rect 889 8359 925 8361
rect 1101 8359 1138 8390
rect 889 8337 1138 8359
rect 970 8331 1081 8337
rect 970 8323 1011 8331
rect 970 8303 978 8323
rect 997 8303 1011 8323
rect 970 8301 1011 8303
rect 1039 8323 1081 8331
rect 1039 8303 1055 8323
rect 1074 8303 1081 8323
rect 1039 8301 1081 8303
rect 970 8286 1081 8301
rect 1309 8291 1346 8390
rect 1622 8386 1686 8398
rect 972 8283 1076 8286
rect 760 8246 881 8256
rect 760 8244 829 8246
rect 760 8203 773 8244
rect 810 8205 829 8244
rect 866 8205 881 8246
rect 810 8203 881 8205
rect 760 8185 881 8203
rect 552 8141 617 8175
rect 972 8141 1076 8143
rect 1307 8141 1348 8291
rect 1726 8283 1753 8538
rect 1815 8528 1895 8539
rect 1815 8502 1832 8528
rect 1872 8502 1895 8528
rect 1815 8475 1895 8502
rect 1815 8449 1836 8475
rect 1876 8449 1895 8475
rect 1815 8430 1895 8449
rect 1815 8404 1839 8430
rect 1879 8404 1895 8430
rect 1815 8353 1895 8404
rect 552 8138 1348 8141
rect 1727 8152 1753 8283
rect 1817 8153 1887 8353
rect 1727 8138 1755 8152
rect 552 8103 1755 8138
rect 1816 8131 1888 8153
rect 552 7946 617 8103
rect 972 8101 1076 8103
rect 1307 8101 1348 8103
rect 1816 8083 1830 8131
rect 1876 8083 1888 8131
rect 1816 8066 1888 8083
rect 2918 8033 2990 9872
rect 3096 8105 3188 11409
rect 3582 11392 3613 11413
rect 4003 11392 4039 11413
rect 3425 11391 3462 11392
rect 3424 11382 3462 11391
rect 3424 11362 3433 11382
rect 3453 11362 3462 11382
rect 3424 11354 3462 11362
rect 3528 11386 3613 11392
rect 3638 11391 3675 11392
rect 3528 11366 3536 11386
rect 3556 11366 3613 11386
rect 3528 11358 3613 11366
rect 3637 11382 3675 11391
rect 3637 11362 3646 11382
rect 3666 11362 3675 11382
rect 3528 11357 3564 11358
rect 3637 11354 3675 11362
rect 3741 11386 3826 11392
rect 3846 11391 3883 11392
rect 3741 11366 3749 11386
rect 3769 11385 3826 11386
rect 3769 11366 3798 11385
rect 3741 11365 3798 11366
rect 3819 11365 3826 11385
rect 3741 11358 3826 11365
rect 3845 11382 3883 11391
rect 3845 11362 3854 11382
rect 3874 11362 3883 11382
rect 3741 11357 3777 11358
rect 3845 11354 3883 11362
rect 3949 11386 4093 11392
rect 3949 11366 3957 11386
rect 3977 11366 4065 11386
rect 4085 11366 4093 11386
rect 3949 11358 4093 11366
rect 3949 11357 3985 11358
rect 4057 11357 4093 11358
rect 4159 11391 4196 11392
rect 4159 11390 4197 11391
rect 4159 11382 4223 11390
rect 4159 11362 4168 11382
rect 4188 11368 4223 11382
rect 4243 11368 4246 11388
rect 4188 11363 4246 11368
rect 4188 11362 4223 11363
rect 3425 11325 3462 11354
rect 3426 11323 3462 11325
rect 3638 11323 3675 11354
rect 3426 11301 3675 11323
rect 3507 11295 3618 11301
rect 3507 11287 3548 11295
rect 3507 11267 3515 11287
rect 3534 11267 3548 11287
rect 3507 11265 3548 11267
rect 3576 11287 3618 11295
rect 3576 11267 3592 11287
rect 3611 11267 3618 11287
rect 3576 11265 3618 11267
rect 3507 11250 3618 11265
rect 3846 11233 3883 11354
rect 4159 11350 4223 11362
rect 3964 11233 3993 11237
rect 4263 11235 4290 11502
rect 4122 11233 4290 11235
rect 3846 11207 4290 11233
rect 3805 10939 3850 10948
rect 3805 10901 3815 10939
rect 3840 10901 3850 10939
rect 3805 10890 3850 10901
rect 3808 10882 3850 10890
rect 3808 10177 3851 10882
rect 3964 10268 3993 11207
rect 4122 11206 4290 11207
rect 3962 10247 3999 10268
rect 3962 10210 3973 10247
rect 3990 10210 3999 10247
rect 3962 10200 3999 10210
rect 3808 10157 4202 10177
rect 4222 10157 4225 10177
rect 3809 10152 4225 10157
rect 3809 10151 4150 10152
rect 3466 10120 3576 10134
rect 3466 10117 3509 10120
rect 3466 10112 3470 10117
rect 3388 10090 3470 10112
rect 3499 10090 3509 10117
rect 3537 10093 3544 10120
rect 3573 10112 3576 10120
rect 3573 10093 3638 10112
rect 3537 10090 3638 10093
rect 3388 10088 3638 10090
rect 3388 10009 3425 10088
rect 3466 10075 3576 10088
rect 3540 10019 3571 10020
rect 3388 9989 3397 10009
rect 3417 9989 3425 10009
rect 3388 9979 3425 9989
rect 3484 10009 3571 10019
rect 3484 9989 3493 10009
rect 3513 9989 3571 10009
rect 3484 9980 3571 9989
rect 3484 9979 3521 9980
rect 3540 9927 3571 9980
rect 3601 10009 3638 10088
rect 3753 10019 3784 10020
rect 3601 9989 3610 10009
rect 3630 9989 3638 10009
rect 3601 9979 3638 9989
rect 3697 10012 3784 10019
rect 3697 10009 3758 10012
rect 3697 9989 3706 10009
rect 3726 9992 3758 10009
rect 3779 9992 3784 10012
rect 3726 9989 3784 9992
rect 3697 9982 3784 9989
rect 3809 10009 3846 10151
rect 4112 10150 4149 10151
rect 3961 10019 3997 10020
rect 3809 9989 3818 10009
rect 3838 9989 3846 10009
rect 3697 9980 3753 9982
rect 3697 9979 3734 9980
rect 3809 9979 3846 9989
rect 3905 10009 4053 10019
rect 4153 10016 4249 10018
rect 3905 9989 3914 10009
rect 3934 9989 4024 10009
rect 4044 9989 4053 10009
rect 3905 9983 4053 9989
rect 3905 9980 3969 9983
rect 3905 9979 3942 9980
rect 3961 9953 3969 9980
rect 3990 9980 4053 9983
rect 4111 10009 4249 10016
rect 4111 9989 4120 10009
rect 4140 9989 4249 10009
rect 4111 9980 4249 9989
rect 3990 9953 3997 9980
rect 4016 9979 4053 9980
rect 4112 9979 4149 9980
rect 3961 9928 3997 9953
rect 3432 9926 3473 9927
rect 3352 9921 3473 9926
rect 3303 9919 3473 9921
rect 3303 9908 3442 9919
rect 3303 9885 3326 9908
rect 3352 9899 3442 9908
rect 3462 9899 3473 9919
rect 3352 9891 3473 9899
rect 3540 9923 3899 9927
rect 3540 9918 3862 9923
rect 3540 9894 3653 9918
rect 3677 9899 3862 9918
rect 3886 9899 3899 9923
rect 3677 9894 3899 9899
rect 3540 9891 3899 9894
rect 3961 9891 3996 9928
rect 4064 9925 4164 9928
rect 4064 9921 4131 9925
rect 4064 9895 4076 9921
rect 4102 9899 4131 9921
rect 4157 9899 4164 9925
rect 4102 9895 4164 9899
rect 4064 9891 4164 9895
rect 3352 9885 3360 9891
rect 3303 9877 3360 9885
rect 3540 9870 3571 9891
rect 3961 9870 3997 9891
rect 3383 9869 3420 9870
rect 3382 9860 3420 9869
rect 3382 9840 3391 9860
rect 3411 9840 3420 9860
rect 3382 9832 3420 9840
rect 3486 9864 3571 9870
rect 3596 9869 3633 9870
rect 3486 9844 3494 9864
rect 3514 9844 3571 9864
rect 3486 9836 3571 9844
rect 3595 9860 3633 9869
rect 3595 9840 3604 9860
rect 3624 9840 3633 9860
rect 3486 9835 3522 9836
rect 3595 9832 3633 9840
rect 3699 9864 3784 9870
rect 3804 9869 3841 9870
rect 3699 9844 3707 9864
rect 3727 9863 3784 9864
rect 3727 9844 3756 9863
rect 3699 9843 3756 9844
rect 3777 9843 3784 9863
rect 3699 9836 3784 9843
rect 3803 9860 3841 9869
rect 3803 9840 3812 9860
rect 3832 9840 3841 9860
rect 3699 9835 3735 9836
rect 3803 9832 3841 9840
rect 3907 9864 4051 9870
rect 3907 9844 3915 9864
rect 3935 9844 4023 9864
rect 4043 9844 4051 9864
rect 3907 9836 4051 9844
rect 3907 9835 3943 9836
rect 4015 9835 4051 9836
rect 4117 9869 4154 9870
rect 4117 9868 4155 9869
rect 4117 9860 4181 9868
rect 4117 9840 4126 9860
rect 4146 9846 4181 9860
rect 4201 9846 4204 9866
rect 4146 9841 4204 9846
rect 4146 9840 4181 9841
rect 3383 9803 3420 9832
rect 3384 9801 3420 9803
rect 3596 9801 3633 9832
rect 3384 9779 3633 9801
rect 3465 9773 3576 9779
rect 3465 9765 3506 9773
rect 3465 9745 3473 9765
rect 3492 9745 3506 9765
rect 3465 9743 3506 9745
rect 3534 9765 3576 9773
rect 3534 9745 3550 9765
rect 3569 9745 3576 9765
rect 3534 9743 3576 9745
rect 3465 9728 3576 9743
rect 3804 9717 3841 9832
rect 4117 9828 4181 9840
rect 3797 9711 3844 9717
rect 4221 9713 4248 9980
rect 4080 9711 4248 9713
rect 3797 9685 4248 9711
rect 3797 9550 3844 9685
rect 4080 9684 4248 9685
rect 3795 9501 3854 9550
rect 3795 9473 3813 9501
rect 3841 9473 3854 9501
rect 3795 9463 3854 9473
rect 4910 8726 4988 11766
rect 4910 8706 5310 8726
rect 5330 8706 5333 8726
rect 4910 8704 5333 8706
rect 4917 8701 5333 8704
rect 4917 8700 5258 8701
rect 4574 8669 4684 8683
rect 4574 8666 4617 8669
rect 4574 8661 4578 8666
rect 4496 8639 4578 8661
rect 4607 8639 4617 8666
rect 4645 8642 4652 8669
rect 4681 8661 4684 8669
rect 4681 8642 4746 8661
rect 4645 8639 4746 8642
rect 4496 8637 4746 8639
rect 4496 8558 4533 8637
rect 4574 8624 4684 8637
rect 4648 8568 4679 8569
rect 4496 8538 4505 8558
rect 4525 8538 4533 8558
rect 4496 8528 4533 8538
rect 4592 8558 4679 8568
rect 4592 8538 4601 8558
rect 4621 8538 4679 8558
rect 4592 8529 4679 8538
rect 4592 8528 4629 8529
rect 4366 8475 4477 8478
rect 4648 8476 4679 8529
rect 4709 8558 4746 8637
rect 4861 8568 4892 8569
rect 4709 8538 4718 8558
rect 4738 8538 4746 8558
rect 4709 8528 4746 8538
rect 4805 8561 4892 8568
rect 4805 8558 4866 8561
rect 4805 8538 4814 8558
rect 4834 8541 4866 8558
rect 4887 8541 4892 8561
rect 4834 8538 4892 8541
rect 4805 8531 4892 8538
rect 4917 8558 4954 8700
rect 5220 8699 5257 8700
rect 5069 8568 5105 8569
rect 4917 8538 4926 8558
rect 4946 8538 4954 8558
rect 4805 8529 4861 8531
rect 4805 8528 4842 8529
rect 4917 8528 4954 8538
rect 5013 8558 5161 8568
rect 5261 8565 5357 8567
rect 5013 8538 5022 8558
rect 5042 8538 5132 8558
rect 5152 8538 5161 8558
rect 5013 8532 5161 8538
rect 5013 8529 5077 8532
rect 5013 8528 5050 8529
rect 5069 8502 5077 8529
rect 5098 8529 5161 8532
rect 5219 8558 5357 8565
rect 5219 8538 5228 8558
rect 5248 8538 5357 8558
rect 5219 8529 5357 8538
rect 5098 8502 5105 8529
rect 5124 8528 5161 8529
rect 5220 8528 5257 8529
rect 5069 8477 5105 8502
rect 4540 8475 4581 8476
rect 4366 8468 4581 8475
rect 4366 8467 4431 8468
rect 4366 8443 4374 8467
rect 4398 8444 4431 8467
rect 4455 8448 4550 8468
rect 4570 8448 4581 8468
rect 4455 8444 4581 8448
rect 4398 8443 4581 8444
rect 4366 8440 4581 8443
rect 4648 8472 5007 8476
rect 4648 8467 4970 8472
rect 4648 8443 4761 8467
rect 4785 8448 4970 8467
rect 4994 8448 5007 8472
rect 4785 8443 5007 8448
rect 4648 8440 5007 8443
rect 5069 8440 5104 8477
rect 5172 8474 5272 8477
rect 5172 8470 5239 8474
rect 5172 8444 5184 8470
rect 5210 8448 5239 8470
rect 5265 8448 5272 8474
rect 5210 8444 5272 8448
rect 5172 8440 5272 8444
rect 4366 8436 4477 8440
rect 4648 8419 4679 8440
rect 5069 8419 5105 8440
rect 4491 8418 4528 8419
rect 4490 8409 4528 8418
rect 4490 8389 4499 8409
rect 4519 8389 4528 8409
rect 4490 8381 4528 8389
rect 4594 8413 4679 8419
rect 4704 8418 4741 8419
rect 4594 8393 4602 8413
rect 4622 8393 4679 8413
rect 4594 8385 4679 8393
rect 4703 8409 4741 8418
rect 4703 8389 4712 8409
rect 4732 8389 4741 8409
rect 4594 8384 4630 8385
rect 4703 8381 4741 8389
rect 4807 8413 4892 8419
rect 4912 8418 4949 8419
rect 4807 8393 4815 8413
rect 4835 8412 4892 8413
rect 4835 8393 4864 8412
rect 4807 8392 4864 8393
rect 4885 8392 4892 8412
rect 4807 8385 4892 8392
rect 4911 8409 4949 8418
rect 4911 8389 4920 8409
rect 4940 8389 4949 8409
rect 4807 8384 4843 8385
rect 4911 8381 4949 8389
rect 5015 8413 5159 8419
rect 5015 8393 5023 8413
rect 5043 8412 5131 8413
rect 5043 8393 5077 8412
rect 5015 8390 5077 8393
rect 5101 8393 5131 8412
rect 5151 8393 5159 8413
rect 5101 8390 5159 8393
rect 5015 8385 5159 8390
rect 5015 8384 5051 8385
rect 5123 8384 5159 8385
rect 5225 8418 5262 8419
rect 5225 8417 5263 8418
rect 5225 8409 5289 8417
rect 5225 8389 5234 8409
rect 5254 8395 5289 8409
rect 5309 8395 5312 8415
rect 5254 8390 5312 8395
rect 5254 8389 5289 8390
rect 4491 8352 4528 8381
rect 4492 8350 4528 8352
rect 4704 8350 4741 8381
rect 4492 8328 4741 8350
rect 4573 8322 4684 8328
rect 4573 8314 4614 8322
rect 4573 8294 4581 8314
rect 4600 8294 4614 8314
rect 4573 8292 4614 8294
rect 4642 8314 4684 8322
rect 4642 8294 4658 8314
rect 4677 8294 4684 8314
rect 4642 8292 4684 8294
rect 4573 8277 4684 8292
rect 4912 8266 4949 8381
rect 5225 8377 5289 8389
rect 4908 8260 4963 8266
rect 5329 8262 5356 8529
rect 5188 8260 5356 8262
rect 4908 8235 5356 8260
rect 5669 8320 5775 13518
rect 8941 13508 8964 13534
rect 9004 13508 9021 13534
rect 8941 13497 9021 13508
rect 9083 13498 9110 13753
rect 9488 13745 9529 13895
rect 10200 13864 11323 13895
rect 12173 13899 12272 13907
rect 12173 13896 12225 13899
rect 9955 13833 10076 13851
rect 9955 13831 10026 13833
rect 9955 13790 9970 13831
rect 10007 13792 10026 13831
rect 10063 13792 10076 13833
rect 10007 13790 10076 13792
rect 9955 13780 10076 13790
rect 9150 13638 9214 13650
rect 9490 13646 9527 13745
rect 9755 13735 9866 13746
rect 9755 13733 9797 13735
rect 9755 13713 9762 13733
rect 9781 13713 9797 13733
rect 9755 13705 9797 13713
rect 9825 13733 9866 13735
rect 9825 13713 9839 13733
rect 9858 13713 9866 13733
rect 9825 13705 9866 13713
rect 9755 13699 9866 13705
rect 9698 13677 9947 13699
rect 9698 13646 9735 13677
rect 9911 13675 9947 13677
rect 9911 13646 9948 13675
rect 9150 13637 9185 13638
rect 9127 13632 9185 13637
rect 9127 13612 9130 13632
rect 9150 13618 9185 13632
rect 9205 13618 9214 13638
rect 9150 13610 9214 13618
rect 9176 13609 9214 13610
rect 9177 13608 9214 13609
rect 9280 13642 9316 13643
rect 9388 13642 9424 13643
rect 9280 13634 9424 13642
rect 9280 13614 9288 13634
rect 9308 13614 9396 13634
rect 9416 13614 9424 13634
rect 9280 13608 9424 13614
rect 9490 13638 9528 13646
rect 9596 13642 9632 13643
rect 9490 13618 9499 13638
rect 9519 13618 9528 13638
rect 9490 13609 9528 13618
rect 9547 13635 9632 13642
rect 9547 13615 9554 13635
rect 9575 13634 9632 13635
rect 9575 13615 9604 13634
rect 9547 13614 9604 13615
rect 9624 13614 9632 13634
rect 9490 13608 9527 13609
rect 9547 13608 9632 13614
rect 9698 13638 9736 13646
rect 9809 13642 9845 13643
rect 9698 13618 9707 13638
rect 9727 13618 9736 13638
rect 9698 13609 9736 13618
rect 9760 13634 9845 13642
rect 9760 13614 9817 13634
rect 9837 13614 9845 13634
rect 9698 13608 9735 13609
rect 9760 13608 9845 13614
rect 9911 13638 9949 13646
rect 9911 13618 9920 13638
rect 9940 13618 9949 13638
rect 10004 13628 10069 13780
rect 10222 13754 10277 13864
rect 11261 13826 11320 13864
rect 12173 13861 12181 13896
rect 12206 13861 12225 13896
rect 12250 13888 12272 13899
rect 13223 13900 14562 13907
rect 13223 13897 13275 13900
rect 12250 13887 13117 13888
rect 12250 13861 13118 13887
rect 12173 13851 13118 13861
rect 12173 13849 12272 13851
rect 11261 13808 11283 13826
rect 11301 13808 11320 13826
rect 11261 13786 11320 13808
rect 11528 13822 12060 13827
rect 11528 13802 12414 13822
rect 12434 13802 12437 13822
rect 13073 13818 13118 13851
rect 13223 13862 13231 13897
rect 13256 13862 13275 13897
rect 13300 13862 14562 13900
rect 13223 13853 14562 13862
rect 13223 13850 13312 13853
rect 13851 13851 14562 13853
rect 11528 13798 12437 13802
rect 9911 13609 9949 13618
rect 10002 13621 10069 13628
rect 9911 13608 9948 13609
rect 9334 13587 9370 13608
rect 9760 13587 9791 13608
rect 10002 13600 10019 13621
rect 10055 13600 10069 13621
rect 10221 13641 10277 13754
rect 11528 13751 11571 13798
rect 12021 13797 12437 13798
rect 13069 13798 13462 13818
rect 13482 13798 13485 13818
rect 12021 13796 12362 13797
rect 11678 13765 11788 13779
rect 11678 13762 11721 13765
rect 11678 13757 11682 13762
rect 11516 13750 11571 13751
rect 10221 13623 10240 13641
rect 10258 13623 10277 13641
rect 10221 13603 10277 13623
rect 11260 13727 11571 13750
rect 11260 13709 11285 13727
rect 11303 13715 11571 13727
rect 11600 13735 11682 13757
rect 11711 13735 11721 13762
rect 11749 13738 11756 13765
rect 11785 13757 11788 13765
rect 11785 13738 11850 13757
rect 11749 13735 11850 13738
rect 11600 13733 11850 13735
rect 11303 13709 11325 13715
rect 10002 13587 10069 13600
rect 9167 13583 9267 13587
rect 9167 13579 9229 13583
rect 9167 13553 9174 13579
rect 9200 13557 9229 13579
rect 9255 13557 9267 13583
rect 9200 13553 9267 13557
rect 9167 13550 9267 13553
rect 9335 13550 9370 13587
rect 9432 13584 9791 13587
rect 9432 13579 9654 13584
rect 9432 13555 9445 13579
rect 9469 13560 9654 13579
rect 9678 13560 9791 13584
rect 9469 13555 9791 13560
rect 9432 13551 9791 13555
rect 9858 13581 10069 13587
rect 9858 13579 10019 13581
rect 9858 13559 9869 13579
rect 9889 13559 10019 13579
rect 9858 13552 10019 13559
rect 9858 13551 9899 13552
rect 9334 13525 9370 13550
rect 9182 13498 9219 13499
rect 9278 13498 9315 13499
rect 9334 13498 9341 13525
rect 9082 13489 9220 13498
rect 9082 13469 9191 13489
rect 9211 13469 9220 13489
rect 9082 13462 9220 13469
rect 9278 13495 9341 13498
rect 9362 13498 9370 13525
rect 9389 13498 9426 13499
rect 9362 13495 9426 13498
rect 9278 13489 9426 13495
rect 9278 13469 9287 13489
rect 9307 13469 9397 13489
rect 9417 13469 9426 13489
rect 9082 13460 9178 13462
rect 9278 13459 9426 13469
rect 9485 13489 9522 13499
rect 9597 13498 9634 13499
rect 9578 13496 9634 13498
rect 9485 13469 9493 13489
rect 9513 13469 9522 13489
rect 9334 13458 9370 13459
rect 9182 13327 9219 13328
rect 9485 13327 9522 13469
rect 9547 13489 9634 13496
rect 9547 13486 9605 13489
rect 9547 13466 9552 13486
rect 9573 13469 9605 13486
rect 9625 13469 9634 13489
rect 9573 13466 9634 13469
rect 9547 13459 9634 13466
rect 9693 13489 9730 13499
rect 9693 13469 9701 13489
rect 9721 13469 9730 13489
rect 9547 13458 9578 13459
rect 9693 13390 9730 13469
rect 9760 13498 9791 13551
rect 10004 13544 10019 13552
rect 10059 13544 10069 13581
rect 11260 13570 11325 13709
rect 11600 13654 11637 13733
rect 11678 13720 11788 13733
rect 11752 13664 11783 13665
rect 11600 13634 11609 13654
rect 11629 13634 11637 13654
rect 10004 13535 10069 13544
rect 10217 13542 10282 13563
rect 10217 13524 10242 13542
rect 10260 13524 10282 13542
rect 11260 13552 11283 13570
rect 11301 13552 11325 13570
rect 11260 13535 11325 13552
rect 11480 13616 11548 13629
rect 11600 13624 11637 13634
rect 11696 13654 11783 13664
rect 11696 13634 11705 13654
rect 11725 13634 11783 13654
rect 11696 13625 11783 13634
rect 11696 13624 11733 13625
rect 11480 13574 11487 13616
rect 11536 13574 11548 13616
rect 11480 13571 11548 13574
rect 11752 13572 11783 13625
rect 11813 13654 11850 13733
rect 11965 13664 11996 13665
rect 11813 13634 11822 13654
rect 11842 13634 11850 13654
rect 11813 13624 11850 13634
rect 11909 13657 11996 13664
rect 11909 13654 11970 13657
rect 11909 13634 11918 13654
rect 11938 13637 11970 13654
rect 11991 13637 11996 13657
rect 11938 13634 11996 13637
rect 11909 13627 11996 13634
rect 12021 13654 12058 13796
rect 12324 13795 12361 13796
rect 13069 13793 13485 13798
rect 13069 13792 13410 13793
rect 12726 13761 12836 13775
rect 12726 13758 12769 13761
rect 12726 13753 12730 13758
rect 12648 13731 12730 13753
rect 12759 13731 12769 13758
rect 12797 13734 12804 13761
rect 12833 13753 12836 13761
rect 12833 13734 12898 13753
rect 12797 13731 12898 13734
rect 12648 13729 12898 13731
rect 12173 13664 12209 13665
rect 12021 13634 12030 13654
rect 12050 13634 12058 13654
rect 11909 13625 11965 13627
rect 11909 13624 11946 13625
rect 12021 13624 12058 13634
rect 12117 13654 12265 13664
rect 12365 13661 12461 13663
rect 12117 13634 12126 13654
rect 12146 13634 12236 13654
rect 12256 13634 12265 13654
rect 12117 13628 12265 13634
rect 12117 13625 12181 13628
rect 12117 13624 12154 13625
rect 12173 13598 12181 13625
rect 12202 13625 12265 13628
rect 12323 13654 12461 13661
rect 12323 13634 12332 13654
rect 12352 13634 12461 13654
rect 12323 13625 12461 13634
rect 12648 13650 12685 13729
rect 12726 13716 12836 13729
rect 12800 13660 12831 13661
rect 12648 13630 12657 13650
rect 12677 13630 12685 13650
rect 12202 13598 12209 13625
rect 12228 13624 12265 13625
rect 12324 13624 12361 13625
rect 12173 13573 12209 13598
rect 11644 13571 11685 13572
rect 11480 13564 11685 13571
rect 11480 13553 11654 13564
rect 9810 13498 9847 13499
rect 9760 13489 9847 13498
rect 9760 13469 9818 13489
rect 9838 13469 9847 13489
rect 9760 13459 9847 13469
rect 9906 13489 9943 13499
rect 9906 13469 9914 13489
rect 9934 13469 9943 13489
rect 9760 13458 9791 13459
rect 9755 13390 9865 13403
rect 9906 13390 9943 13469
rect 10217 13448 10282 13524
rect 11480 13520 11488 13553
rect 11481 13511 11488 13520
rect 11537 13544 11654 13553
rect 11674 13544 11685 13564
rect 11537 13536 11685 13544
rect 11752 13568 12111 13572
rect 11752 13563 12074 13568
rect 11752 13539 11865 13563
rect 11889 13544 12074 13563
rect 12098 13544 12111 13568
rect 11889 13539 12111 13544
rect 11752 13536 12111 13539
rect 12173 13536 12208 13573
rect 12276 13570 12376 13573
rect 12276 13566 12343 13570
rect 12276 13540 12288 13566
rect 12314 13544 12343 13566
rect 12369 13544 12376 13570
rect 12314 13540 12376 13544
rect 12276 13536 12376 13540
rect 11537 13520 11548 13536
rect 11537 13511 11545 13520
rect 11752 13515 11783 13536
rect 12173 13515 12209 13536
rect 11595 13514 11632 13515
rect 11260 13471 11325 13490
rect 11260 13453 11285 13471
rect 11303 13453 11325 13471
rect 9693 13388 9943 13390
rect 9693 13385 9794 13388
rect 9693 13366 9758 13385
rect 9755 13358 9758 13366
rect 9787 13358 9794 13385
rect 9822 13361 9832 13388
rect 9861 13366 9943 13388
rect 9966 13413 10283 13448
rect 9861 13361 9865 13366
rect 9822 13358 9865 13361
rect 9755 13344 9865 13358
rect 9181 13326 9522 13327
rect 9106 13324 9522 13326
rect 9966 13324 10006 13413
rect 10217 13386 10282 13413
rect 10217 13368 10240 13386
rect 10258 13368 10282 13386
rect 10217 13348 10282 13368
rect 9103 13321 10006 13324
rect 9103 13301 9109 13321
rect 9129 13301 10006 13321
rect 9103 13297 10006 13301
rect 9966 13294 10006 13297
rect 10218 13287 10283 13308
rect 8436 13279 9097 13280
rect 8436 13272 9370 13279
rect 8436 13271 9342 13272
rect 8436 13251 9287 13271
rect 9319 13252 9342 13271
rect 9367 13252 9370 13272
rect 9319 13251 9370 13252
rect 8436 13244 9370 13251
rect 8035 13202 8203 13203
rect 8438 13202 8477 13244
rect 9266 13242 9370 13244
rect 9335 13240 9370 13242
rect 10218 13269 10242 13287
rect 10260 13269 10283 13287
rect 10218 13222 10283 13269
rect 8035 13176 8479 13202
rect 8035 13174 8203 13176
rect 8035 12823 8062 13174
rect 8438 13170 8479 13176
rect 8102 12963 8166 12975
rect 8442 12971 8479 13170
rect 8941 13197 9013 13214
rect 8941 13158 8949 13197
rect 8994 13158 9013 13197
rect 8707 13060 8818 13075
rect 8707 13058 8749 13060
rect 8707 13038 8714 13058
rect 8733 13038 8749 13058
rect 8707 13030 8749 13038
rect 8777 13058 8818 13060
rect 8777 13038 8791 13058
rect 8810 13038 8818 13058
rect 8777 13030 8818 13038
rect 8707 13024 8818 13030
rect 8650 13002 8899 13024
rect 8650 12971 8687 13002
rect 8863 13000 8899 13002
rect 8863 12971 8900 13000
rect 8102 12962 8137 12963
rect 8079 12957 8137 12962
rect 8079 12937 8082 12957
rect 8102 12943 8137 12957
rect 8157 12943 8166 12963
rect 8102 12935 8166 12943
rect 8128 12934 8166 12935
rect 8129 12933 8166 12934
rect 8232 12967 8268 12968
rect 8340 12967 8376 12968
rect 8232 12959 8376 12967
rect 8232 12939 8240 12959
rect 8260 12939 8348 12959
rect 8368 12939 8376 12959
rect 8232 12933 8376 12939
rect 8442 12963 8480 12971
rect 8548 12967 8584 12968
rect 8442 12943 8451 12963
rect 8471 12943 8480 12963
rect 8442 12934 8480 12943
rect 8499 12960 8584 12967
rect 8499 12940 8506 12960
rect 8527 12959 8584 12960
rect 8527 12940 8556 12959
rect 8499 12939 8556 12940
rect 8576 12939 8584 12959
rect 8442 12933 8479 12934
rect 8499 12933 8584 12939
rect 8650 12963 8688 12971
rect 8761 12967 8797 12968
rect 8650 12943 8659 12963
rect 8679 12943 8688 12963
rect 8650 12934 8688 12943
rect 8712 12959 8797 12967
rect 8712 12939 8769 12959
rect 8789 12939 8797 12959
rect 8650 12933 8687 12934
rect 8712 12933 8797 12939
rect 8863 12963 8901 12971
rect 8863 12943 8872 12963
rect 8892 12943 8901 12963
rect 8863 12934 8901 12943
rect 8941 12948 9013 13158
rect 9083 13192 10283 13222
rect 9083 13191 9527 13192
rect 9083 13189 9251 13191
rect 8941 12934 9024 12948
rect 8863 12933 8900 12934
rect 8286 12912 8322 12933
rect 8712 12912 8743 12933
rect 8941 12912 8958 12934
rect 8119 12908 8219 12912
rect 8119 12904 8181 12908
rect 8119 12878 8126 12904
rect 8152 12882 8181 12904
rect 8207 12882 8219 12908
rect 8152 12878 8219 12882
rect 8119 12875 8219 12878
rect 8287 12875 8322 12912
rect 8384 12909 8743 12912
rect 8384 12904 8606 12909
rect 8384 12880 8397 12904
rect 8421 12885 8606 12904
rect 8630 12885 8743 12909
rect 8421 12880 8743 12885
rect 8384 12876 8743 12880
rect 8810 12904 8958 12912
rect 8810 12884 8821 12904
rect 8841 12901 8958 12904
rect 9011 12901 9024 12934
rect 8841 12884 9024 12901
rect 8810 12877 9024 12884
rect 8810 12876 8851 12877
rect 8941 12876 9024 12877
rect 8286 12850 8322 12875
rect 8134 12823 8171 12824
rect 8230 12823 8267 12824
rect 8286 12823 8293 12850
rect 8034 12814 8172 12823
rect 8034 12794 8143 12814
rect 8163 12794 8172 12814
rect 8034 12787 8172 12794
rect 8230 12820 8293 12823
rect 8314 12823 8322 12850
rect 8341 12823 8378 12824
rect 8314 12820 8378 12823
rect 8230 12814 8378 12820
rect 8230 12794 8239 12814
rect 8259 12794 8349 12814
rect 8369 12794 8378 12814
rect 8034 12785 8130 12787
rect 8230 12784 8378 12794
rect 8437 12814 8474 12824
rect 8549 12823 8586 12824
rect 8530 12821 8586 12823
rect 8437 12794 8445 12814
rect 8465 12794 8474 12814
rect 8286 12783 8322 12784
rect 8134 12652 8171 12653
rect 8437 12652 8474 12794
rect 8499 12814 8586 12821
rect 8499 12811 8557 12814
rect 8499 12791 8504 12811
rect 8525 12794 8557 12811
rect 8577 12794 8586 12814
rect 8525 12791 8586 12794
rect 8499 12784 8586 12791
rect 8645 12814 8682 12824
rect 8645 12794 8653 12814
rect 8673 12794 8682 12814
rect 8499 12783 8530 12784
rect 8645 12715 8682 12794
rect 8712 12823 8743 12876
rect 8949 12843 8963 12876
rect 9016 12843 9024 12876
rect 8949 12837 9024 12843
rect 8949 12832 9019 12837
rect 8762 12823 8799 12824
rect 8712 12814 8799 12823
rect 8712 12794 8770 12814
rect 8790 12794 8799 12814
rect 8712 12784 8799 12794
rect 8858 12814 8895 12824
rect 9083 12819 9110 13189
rect 9150 12959 9214 12971
rect 9490 12967 9527 13191
rect 9998 13172 10062 13174
rect 9994 13160 10062 13172
rect 9994 13127 10005 13160
rect 10045 13127 10062 13160
rect 9994 13117 10062 13127
rect 9755 13056 9866 13071
rect 9755 13054 9797 13056
rect 9755 13034 9762 13054
rect 9781 13034 9797 13054
rect 9755 13026 9797 13034
rect 9825 13054 9866 13056
rect 9825 13034 9839 13054
rect 9858 13034 9866 13054
rect 9825 13026 9866 13034
rect 9755 13020 9866 13026
rect 9698 12998 9947 13020
rect 9698 12967 9735 12998
rect 9911 12996 9947 12998
rect 9911 12967 9948 12996
rect 9150 12958 9185 12959
rect 9127 12953 9185 12958
rect 9127 12933 9130 12953
rect 9150 12939 9185 12953
rect 9205 12939 9214 12959
rect 9150 12931 9214 12939
rect 9176 12930 9214 12931
rect 9177 12929 9214 12930
rect 9280 12963 9316 12964
rect 9388 12963 9424 12964
rect 9280 12955 9424 12963
rect 9280 12935 9288 12955
rect 9308 12935 9396 12955
rect 9416 12935 9424 12955
rect 9280 12929 9424 12935
rect 9490 12959 9528 12967
rect 9596 12963 9632 12964
rect 9490 12939 9499 12959
rect 9519 12939 9528 12959
rect 9490 12930 9528 12939
rect 9547 12956 9632 12963
rect 9547 12936 9554 12956
rect 9575 12955 9632 12956
rect 9575 12936 9604 12955
rect 9547 12935 9604 12936
rect 9624 12935 9632 12955
rect 9490 12929 9527 12930
rect 9547 12929 9632 12935
rect 9698 12959 9736 12967
rect 9809 12963 9845 12964
rect 9698 12939 9707 12959
rect 9727 12939 9736 12959
rect 9698 12930 9736 12939
rect 9760 12955 9845 12963
rect 9760 12935 9817 12955
rect 9837 12935 9845 12955
rect 9698 12929 9735 12930
rect 9760 12929 9845 12935
rect 9911 12959 9949 12967
rect 9911 12939 9920 12959
rect 9940 12939 9949 12959
rect 9911 12930 9949 12939
rect 9998 12933 10062 13117
rect 10218 12991 10283 13192
rect 11260 13252 11325 13453
rect 11481 13327 11545 13511
rect 11594 13505 11632 13514
rect 11594 13485 11603 13505
rect 11623 13485 11632 13505
rect 11594 13477 11632 13485
rect 11698 13509 11783 13515
rect 11808 13514 11845 13515
rect 11698 13489 11706 13509
rect 11726 13489 11783 13509
rect 11698 13481 11783 13489
rect 11807 13505 11845 13514
rect 11807 13485 11816 13505
rect 11836 13485 11845 13505
rect 11698 13480 11734 13481
rect 11807 13477 11845 13485
rect 11911 13509 11996 13515
rect 12016 13514 12053 13515
rect 11911 13489 11919 13509
rect 11939 13508 11996 13509
rect 11939 13489 11968 13508
rect 11911 13488 11968 13489
rect 11989 13488 11996 13508
rect 11911 13481 11996 13488
rect 12015 13505 12053 13514
rect 12015 13485 12024 13505
rect 12044 13485 12053 13505
rect 11911 13480 11947 13481
rect 12015 13477 12053 13485
rect 12119 13509 12263 13515
rect 12119 13489 12127 13509
rect 12147 13489 12235 13509
rect 12255 13489 12263 13509
rect 12119 13481 12263 13489
rect 12119 13480 12155 13481
rect 12227 13480 12263 13481
rect 12329 13514 12366 13515
rect 12329 13513 12367 13514
rect 12329 13505 12393 13513
rect 12329 13485 12338 13505
rect 12358 13491 12393 13505
rect 12413 13491 12416 13511
rect 12358 13486 12416 13491
rect 12358 13485 12393 13486
rect 11595 13448 11632 13477
rect 11596 13446 11632 13448
rect 11808 13446 11845 13477
rect 11596 13424 11845 13446
rect 11677 13418 11788 13424
rect 11677 13410 11718 13418
rect 11677 13390 11685 13410
rect 11704 13390 11718 13410
rect 11677 13388 11718 13390
rect 11746 13410 11788 13418
rect 11746 13390 11762 13410
rect 11781 13390 11788 13410
rect 11746 13388 11788 13390
rect 11677 13373 11788 13388
rect 11481 13317 11549 13327
rect 11481 13284 11498 13317
rect 11538 13284 11549 13317
rect 11481 13272 11549 13284
rect 11481 13270 11545 13272
rect 12016 13253 12053 13477
rect 12329 13473 12393 13485
rect 12433 13255 12460 13625
rect 12648 13620 12685 13630
rect 12744 13650 12831 13660
rect 12744 13630 12753 13650
rect 12773 13630 12831 13650
rect 12744 13621 12831 13630
rect 12744 13620 12781 13621
rect 12524 13607 12594 13612
rect 12519 13601 12594 13607
rect 12519 13568 12527 13601
rect 12580 13568 12594 13601
rect 12800 13568 12831 13621
rect 12861 13650 12898 13729
rect 13013 13660 13044 13661
rect 12861 13630 12870 13650
rect 12890 13630 12898 13650
rect 12861 13620 12898 13630
rect 12957 13653 13044 13660
rect 12957 13650 13018 13653
rect 12957 13630 12966 13650
rect 12986 13633 13018 13650
rect 13039 13633 13044 13653
rect 12986 13630 13044 13633
rect 12957 13623 13044 13630
rect 13069 13650 13106 13792
rect 13372 13791 13409 13792
rect 13221 13660 13257 13661
rect 13069 13630 13078 13650
rect 13098 13630 13106 13650
rect 12957 13621 13013 13623
rect 12957 13620 12994 13621
rect 13069 13620 13106 13630
rect 13165 13650 13313 13660
rect 13413 13657 13509 13659
rect 13165 13630 13174 13650
rect 13194 13630 13284 13650
rect 13304 13630 13313 13650
rect 13165 13624 13313 13630
rect 13165 13621 13229 13624
rect 13165 13620 13202 13621
rect 13221 13594 13229 13621
rect 13250 13621 13313 13624
rect 13371 13650 13509 13657
rect 13371 13630 13380 13650
rect 13400 13630 13509 13650
rect 13371 13621 13509 13630
rect 13250 13594 13257 13621
rect 13276 13620 13313 13621
rect 13372 13620 13409 13621
rect 13221 13569 13257 13594
rect 12519 13567 12602 13568
rect 12692 13567 12733 13568
rect 12519 13560 12733 13567
rect 12519 13543 12702 13560
rect 12519 13510 12532 13543
rect 12585 13540 12702 13543
rect 12722 13540 12733 13560
rect 12585 13532 12733 13540
rect 12800 13564 13159 13568
rect 12800 13559 13122 13564
rect 12800 13535 12913 13559
rect 12937 13540 13122 13559
rect 13146 13540 13159 13564
rect 12937 13535 13159 13540
rect 12800 13532 13159 13535
rect 13221 13532 13256 13569
rect 13324 13566 13424 13569
rect 13324 13562 13391 13566
rect 13324 13536 13336 13562
rect 13362 13540 13391 13562
rect 13417 13540 13424 13566
rect 13362 13536 13424 13540
rect 13324 13532 13424 13536
rect 12585 13510 12602 13532
rect 12800 13511 12831 13532
rect 13221 13511 13257 13532
rect 12643 13510 12680 13511
rect 12519 13496 12602 13510
rect 12292 13253 12460 13255
rect 12016 13252 12460 13253
rect 11260 13222 12460 13252
rect 12530 13286 12602 13496
rect 12642 13501 12680 13510
rect 12642 13481 12651 13501
rect 12671 13481 12680 13501
rect 12642 13473 12680 13481
rect 12746 13505 12831 13511
rect 12856 13510 12893 13511
rect 12746 13485 12754 13505
rect 12774 13485 12831 13505
rect 12746 13477 12831 13485
rect 12855 13501 12893 13510
rect 12855 13481 12864 13501
rect 12884 13481 12893 13501
rect 12746 13476 12782 13477
rect 12855 13473 12893 13481
rect 12959 13505 13044 13511
rect 13064 13510 13101 13511
rect 12959 13485 12967 13505
rect 12987 13504 13044 13505
rect 12987 13485 13016 13504
rect 12959 13484 13016 13485
rect 13037 13484 13044 13504
rect 12959 13477 13044 13484
rect 13063 13501 13101 13510
rect 13063 13481 13072 13501
rect 13092 13481 13101 13501
rect 12959 13476 12995 13477
rect 13063 13473 13101 13481
rect 13167 13505 13311 13511
rect 13167 13485 13175 13505
rect 13195 13485 13283 13505
rect 13303 13485 13311 13505
rect 13167 13477 13311 13485
rect 13167 13476 13203 13477
rect 13275 13476 13311 13477
rect 13377 13510 13414 13511
rect 13377 13509 13415 13510
rect 13377 13501 13441 13509
rect 13377 13481 13386 13501
rect 13406 13487 13441 13501
rect 13461 13487 13464 13507
rect 13406 13482 13464 13487
rect 13406 13481 13441 13482
rect 12643 13444 12680 13473
rect 12644 13442 12680 13444
rect 12856 13442 12893 13473
rect 12644 13420 12893 13442
rect 12725 13414 12836 13420
rect 12725 13406 12766 13414
rect 12725 13386 12733 13406
rect 12752 13386 12766 13406
rect 12725 13384 12766 13386
rect 12794 13406 12836 13414
rect 12794 13386 12810 13406
rect 12829 13386 12836 13406
rect 12794 13384 12836 13386
rect 12725 13369 12836 13384
rect 12530 13247 12549 13286
rect 12594 13247 12602 13286
rect 12530 13230 12602 13247
rect 13064 13274 13101 13473
rect 13377 13469 13441 13481
rect 13064 13268 13105 13274
rect 13481 13270 13508 13621
rect 13803 13608 13898 13634
rect 13639 13586 13703 13605
rect 13639 13547 13652 13586
rect 13686 13547 13703 13586
rect 13639 13528 13703 13547
rect 13340 13268 13508 13270
rect 13064 13242 13508 13268
rect 11260 13175 11325 13222
rect 11260 13157 11283 13175
rect 11301 13157 11325 13175
rect 12173 13202 12208 13204
rect 12173 13200 12277 13202
rect 13066 13200 13105 13242
rect 13340 13241 13508 13242
rect 12173 13193 13107 13200
rect 12173 13192 12224 13193
rect 12173 13172 12176 13192
rect 12201 13173 12224 13192
rect 12256 13173 13107 13193
rect 12201 13172 13107 13173
rect 12173 13165 13107 13172
rect 12446 13164 13107 13165
rect 11260 13136 11325 13157
rect 11537 13147 11577 13150
rect 11537 13143 12440 13147
rect 11537 13123 12414 13143
rect 12434 13123 12440 13143
rect 11537 13120 12440 13123
rect 11261 13076 11326 13096
rect 11261 13058 11285 13076
rect 11303 13058 11326 13076
rect 11261 13031 11326 13058
rect 11537 13031 11577 13120
rect 12021 13118 12437 13120
rect 12021 13117 12362 13118
rect 11678 13086 11788 13100
rect 11678 13083 11721 13086
rect 11678 13078 11682 13083
rect 11260 12996 11577 13031
rect 11600 13056 11682 13078
rect 11711 13056 11721 13083
rect 11749 13059 11756 13086
rect 11785 13078 11788 13086
rect 11785 13059 11850 13078
rect 11749 13056 11850 13059
rect 11600 13054 11850 13056
rect 10218 12973 10240 12991
rect 10258 12973 10283 12991
rect 10218 12954 10283 12973
rect 9911 12929 9948 12930
rect 9334 12908 9370 12929
rect 9760 12908 9791 12929
rect 9998 12924 10006 12933
rect 9995 12908 10006 12924
rect 9167 12904 9267 12908
rect 9167 12900 9229 12904
rect 9167 12874 9174 12900
rect 9200 12878 9229 12900
rect 9255 12878 9267 12904
rect 9200 12874 9267 12878
rect 9167 12871 9267 12874
rect 9335 12871 9370 12908
rect 9432 12905 9791 12908
rect 9432 12900 9654 12905
rect 9432 12876 9445 12900
rect 9469 12881 9654 12900
rect 9678 12881 9791 12905
rect 9469 12876 9791 12881
rect 9432 12872 9791 12876
rect 9858 12900 10006 12908
rect 9858 12880 9869 12900
rect 9889 12891 10006 12900
rect 10055 12924 10062 12933
rect 10055 12891 10063 12924
rect 11261 12920 11326 12996
rect 11600 12975 11637 13054
rect 11678 13041 11788 13054
rect 11752 12985 11783 12986
rect 11600 12955 11609 12975
rect 11629 12955 11637 12975
rect 11600 12945 11637 12955
rect 11696 12975 11783 12985
rect 11696 12955 11705 12975
rect 11725 12955 11783 12975
rect 11696 12946 11783 12955
rect 11696 12945 11733 12946
rect 9889 12880 10063 12891
rect 9858 12873 10063 12880
rect 9858 12872 9899 12873
rect 9334 12846 9370 12871
rect 9182 12819 9219 12820
rect 9278 12819 9315 12820
rect 9334 12819 9341 12846
rect 8858 12794 8866 12814
rect 8886 12794 8895 12814
rect 8712 12783 8743 12784
rect 8707 12715 8817 12728
rect 8858 12715 8895 12794
rect 9082 12810 9220 12819
rect 9082 12790 9191 12810
rect 9211 12790 9220 12810
rect 9082 12783 9220 12790
rect 9278 12816 9341 12819
rect 9362 12819 9370 12846
rect 9389 12819 9426 12820
rect 9362 12816 9426 12819
rect 9278 12810 9426 12816
rect 9278 12790 9287 12810
rect 9307 12790 9397 12810
rect 9417 12790 9426 12810
rect 9082 12781 9178 12783
rect 9278 12780 9426 12790
rect 9485 12810 9522 12820
rect 9597 12819 9634 12820
rect 9578 12817 9634 12819
rect 9485 12790 9493 12810
rect 9513 12790 9522 12810
rect 9334 12779 9370 12780
rect 8645 12713 8895 12715
rect 8645 12710 8746 12713
rect 8645 12691 8710 12710
rect 8707 12683 8710 12691
rect 8739 12683 8746 12710
rect 8774 12686 8784 12713
rect 8813 12691 8895 12713
rect 8813 12686 8817 12691
rect 8774 12683 8817 12686
rect 8707 12669 8817 12683
rect 8133 12651 8474 12652
rect 8058 12646 8474 12651
rect 9182 12648 9219 12649
rect 9485 12648 9522 12790
rect 9547 12810 9634 12817
rect 9547 12807 9605 12810
rect 9547 12787 9552 12807
rect 9573 12790 9605 12807
rect 9625 12790 9634 12810
rect 9573 12787 9634 12790
rect 9547 12780 9634 12787
rect 9693 12810 9730 12820
rect 9693 12790 9701 12810
rect 9721 12790 9730 12810
rect 9547 12779 9578 12780
rect 9693 12711 9730 12790
rect 9760 12819 9791 12872
rect 9995 12870 10063 12873
rect 9995 12828 10007 12870
rect 10056 12828 10063 12870
rect 9810 12819 9847 12820
rect 9760 12810 9847 12819
rect 9760 12790 9818 12810
rect 9838 12790 9847 12810
rect 9760 12780 9847 12790
rect 9906 12810 9943 12820
rect 9995 12815 10063 12828
rect 10218 12892 10283 12909
rect 10218 12874 10242 12892
rect 10260 12874 10283 12892
rect 11261 12902 11283 12920
rect 11301 12902 11326 12920
rect 11261 12881 11326 12902
rect 11474 12900 11539 12909
rect 9906 12790 9914 12810
rect 9934 12790 9943 12810
rect 9760 12779 9791 12780
rect 9755 12711 9865 12724
rect 9906 12711 9943 12790
rect 10218 12735 10283 12874
rect 11474 12863 11484 12900
rect 11524 12892 11539 12900
rect 11752 12893 11783 12946
rect 11813 12975 11850 13054
rect 11965 12985 11996 12986
rect 11813 12955 11822 12975
rect 11842 12955 11850 12975
rect 11813 12945 11850 12955
rect 11909 12978 11996 12985
rect 11909 12975 11970 12978
rect 11909 12955 11918 12975
rect 11938 12958 11970 12975
rect 11991 12958 11996 12978
rect 11938 12955 11996 12958
rect 11909 12948 11996 12955
rect 12021 12975 12058 13117
rect 12324 13116 12361 13117
rect 13641 13057 13703 13528
rect 13803 13567 13829 13608
rect 13865 13567 13898 13608
rect 13803 13271 13898 13567
rect 13803 13227 13818 13271
rect 13878 13227 13898 13271
rect 13803 13207 13898 13227
rect 14515 13138 14558 13851
rect 15098 13793 15244 13804
rect 15098 13777 16480 13793
rect 15098 13772 16507 13777
rect 15098 13766 15190 13772
rect 15098 13669 15130 13766
rect 15168 13675 15190 13766
rect 15228 13675 16507 13772
rect 19657 13677 19727 13930
rect 20196 13927 20237 13929
rect 20468 13927 20572 13929
rect 22226 13927 22285 13934
rect 19789 13892 22285 13927
rect 24816 13913 25527 13915
rect 24189 13912 25527 13913
rect 23139 13911 23211 13912
rect 19789 13878 19817 13892
rect 19791 13747 19817 13878
rect 20196 13889 22285 13892
rect 15168 13669 16507 13675
rect 15098 13642 16507 13669
rect 16377 13567 16507 13642
rect 19649 13626 19729 13677
rect 19649 13600 19665 13626
rect 19705 13600 19729 13626
rect 19649 13581 19729 13600
rect 14515 13118 14909 13138
rect 14929 13118 14932 13138
rect 14516 13113 14932 13118
rect 14516 13112 14857 13113
rect 14173 13081 14283 13095
rect 14173 13078 14216 13081
rect 14173 13073 14177 13078
rect 13636 13005 13711 13057
rect 14095 13051 14177 13073
rect 14206 13051 14216 13078
rect 14244 13054 14251 13081
rect 14280 13073 14283 13081
rect 14280 13054 14345 13073
rect 14244 13051 14345 13054
rect 14095 13049 14345 13051
rect 14005 13005 14051 13006
rect 12173 12985 12209 12986
rect 12021 12955 12030 12975
rect 12050 12955 12058 12975
rect 11909 12946 11965 12948
rect 11909 12945 11946 12946
rect 12021 12945 12058 12955
rect 12117 12975 12265 12985
rect 12365 12982 12461 12984
rect 12117 12955 12126 12975
rect 12146 12955 12236 12975
rect 12256 12955 12265 12975
rect 12117 12949 12265 12955
rect 12117 12946 12181 12949
rect 12117 12945 12154 12946
rect 12173 12919 12181 12946
rect 12202 12946 12265 12949
rect 12323 12975 12461 12982
rect 12323 12955 12332 12975
rect 12352 12955 12461 12975
rect 12323 12946 12461 12955
rect 13636 12970 14051 13005
rect 12202 12919 12209 12946
rect 12228 12945 12265 12946
rect 12324 12945 12361 12946
rect 12173 12894 12209 12919
rect 11644 12892 11685 12893
rect 11524 12885 11685 12892
rect 11524 12865 11654 12885
rect 11674 12865 11685 12885
rect 11524 12863 11685 12865
rect 11474 12857 11685 12863
rect 11752 12889 12111 12893
rect 11752 12884 12074 12889
rect 11752 12860 11865 12884
rect 11889 12865 12074 12884
rect 12098 12865 12111 12889
rect 11889 12860 12111 12865
rect 11752 12857 12111 12860
rect 12173 12857 12208 12894
rect 12276 12891 12376 12894
rect 12276 12887 12343 12891
rect 12276 12861 12288 12887
rect 12314 12865 12343 12887
rect 12369 12865 12376 12891
rect 12314 12861 12376 12865
rect 12276 12857 12376 12861
rect 11474 12844 11541 12857
rect 10218 12729 10240 12735
rect 9693 12709 9943 12711
rect 9693 12706 9794 12709
rect 9693 12687 9758 12706
rect 9755 12679 9758 12687
rect 9787 12679 9794 12706
rect 9822 12682 9832 12709
rect 9861 12687 9943 12709
rect 9972 12717 10240 12729
rect 10258 12717 10283 12735
rect 9972 12694 10283 12717
rect 11266 12821 11322 12841
rect 11266 12803 11285 12821
rect 11303 12803 11322 12821
rect 9972 12693 10027 12694
rect 9861 12682 9865 12687
rect 9822 12679 9865 12682
rect 9755 12665 9865 12679
rect 9181 12647 9522 12648
rect 8058 12626 8061 12646
rect 8081 12626 8474 12646
rect 9106 12646 9522 12647
rect 9972 12646 10015 12693
rect 11266 12690 11322 12803
rect 11474 12823 11488 12844
rect 11524 12823 11541 12844
rect 11752 12836 11783 12857
rect 12173 12836 12209 12857
rect 11595 12835 11632 12836
rect 11474 12816 11541 12823
rect 11594 12826 11632 12835
rect 9106 12642 10015 12646
rect 8425 12593 8470 12626
rect 9106 12622 9109 12642
rect 9129 12622 10015 12642
rect 9483 12617 10015 12622
rect 10223 12636 10282 12658
rect 10223 12618 10242 12636
rect 10260 12618 10282 12636
rect 9271 12593 9370 12595
rect 8425 12583 9370 12593
rect 6982 12563 7041 12573
rect 6982 12535 6995 12563
rect 7023 12535 7041 12563
rect 8425 12557 9293 12583
rect 8426 12556 9293 12557
rect 9271 12545 9293 12556
rect 9318 12548 9337 12583
rect 9362 12548 9370 12583
rect 9318 12545 9370 12548
rect 10223 12547 10282 12618
rect 11266 12552 11321 12690
rect 11474 12664 11539 12816
rect 11594 12806 11603 12826
rect 11623 12806 11632 12826
rect 11594 12798 11632 12806
rect 11698 12830 11783 12836
rect 11808 12835 11845 12836
rect 11698 12810 11706 12830
rect 11726 12810 11783 12830
rect 11698 12802 11783 12810
rect 11807 12826 11845 12835
rect 11807 12806 11816 12826
rect 11836 12806 11845 12826
rect 11698 12801 11734 12802
rect 11807 12798 11845 12806
rect 11911 12830 11996 12836
rect 12016 12835 12053 12836
rect 11911 12810 11919 12830
rect 11939 12829 11996 12830
rect 11939 12810 11968 12829
rect 11911 12809 11968 12810
rect 11989 12809 11996 12829
rect 11911 12802 11996 12809
rect 12015 12826 12053 12835
rect 12015 12806 12024 12826
rect 12044 12806 12053 12826
rect 11911 12801 11947 12802
rect 12015 12798 12053 12806
rect 12119 12830 12263 12836
rect 12119 12810 12127 12830
rect 12147 12810 12235 12830
rect 12255 12810 12263 12830
rect 12119 12802 12263 12810
rect 12119 12801 12155 12802
rect 12227 12801 12263 12802
rect 12329 12835 12366 12836
rect 12329 12834 12367 12835
rect 12329 12826 12393 12834
rect 12329 12806 12338 12826
rect 12358 12812 12393 12826
rect 12413 12812 12416 12832
rect 12358 12807 12416 12812
rect 12358 12806 12393 12807
rect 11595 12769 11632 12798
rect 11596 12767 11632 12769
rect 11808 12767 11845 12798
rect 11596 12745 11845 12767
rect 11677 12739 11788 12745
rect 11677 12731 11718 12739
rect 11677 12711 11685 12731
rect 11704 12711 11718 12731
rect 11677 12709 11718 12711
rect 11746 12731 11788 12739
rect 11746 12711 11762 12731
rect 11781 12711 11788 12731
rect 11746 12709 11788 12711
rect 11677 12696 11788 12709
rect 12016 12699 12053 12798
rect 12329 12794 12393 12806
rect 11467 12654 11588 12664
rect 11467 12652 11536 12654
rect 11467 12611 11480 12652
rect 11517 12613 11536 12652
rect 11573 12613 11588 12654
rect 11517 12611 11588 12613
rect 11467 12593 11588 12611
rect 11259 12549 11323 12552
rect 11679 12549 11783 12555
rect 12014 12549 12055 12699
rect 12433 12691 12460 12946
rect 12522 12936 12602 12947
rect 12522 12910 12539 12936
rect 12579 12910 12602 12936
rect 12522 12883 12602 12910
rect 12522 12857 12543 12883
rect 12583 12857 12602 12883
rect 12522 12838 12602 12857
rect 12522 12812 12546 12838
rect 12586 12812 12602 12838
rect 12522 12761 12602 12812
rect 9271 12537 9370 12545
rect 9297 12536 9369 12537
rect 6982 12486 7041 12535
rect 8951 12510 9018 12529
rect 8951 12489 8968 12510
rect 6588 12351 6756 12352
rect 6992 12351 7039 12486
rect 6588 12325 7039 12351
rect 6588 12323 6756 12325
rect 6588 12056 6615 12323
rect 6992 12319 7039 12325
rect 8949 12444 8968 12489
rect 8998 12489 9018 12510
rect 8998 12444 9019 12489
rect 9488 12486 9529 12488
rect 9760 12486 9864 12488
rect 10220 12486 10284 12547
rect 6655 12196 6719 12208
rect 6995 12204 7032 12319
rect 7260 12293 7371 12308
rect 7260 12291 7302 12293
rect 7260 12271 7267 12291
rect 7286 12271 7302 12291
rect 7260 12263 7302 12271
rect 7330 12291 7371 12293
rect 7330 12271 7344 12291
rect 7363 12271 7371 12291
rect 7330 12263 7371 12271
rect 7260 12257 7371 12263
rect 7203 12235 7452 12257
rect 8949 12236 9019 12444
rect 9081 12451 10284 12486
rect 9081 12437 9109 12451
rect 9083 12306 9109 12437
rect 9488 12448 10284 12451
rect 11259 12546 12055 12549
rect 12434 12560 12460 12691
rect 12434 12546 12462 12560
rect 11259 12511 12462 12546
rect 12524 12553 12594 12761
rect 13636 12686 13711 12970
rect 14005 12887 14051 12970
rect 14095 12970 14132 13049
rect 14173 13036 14283 13049
rect 14247 12980 14278 12981
rect 14095 12950 14104 12970
rect 14124 12950 14132 12970
rect 14095 12940 14132 12950
rect 14191 12970 14278 12980
rect 14191 12950 14200 12970
rect 14220 12950 14278 12970
rect 14191 12941 14278 12950
rect 14191 12940 14228 12941
rect 14247 12888 14278 12941
rect 14308 12970 14345 13049
rect 14460 12980 14491 12981
rect 14308 12950 14317 12970
rect 14337 12950 14345 12970
rect 14308 12940 14345 12950
rect 14404 12973 14491 12980
rect 14404 12970 14465 12973
rect 14404 12950 14413 12970
rect 14433 12953 14465 12970
rect 14486 12953 14491 12973
rect 14433 12950 14491 12953
rect 14404 12943 14491 12950
rect 14516 12970 14553 13112
rect 14819 13111 14856 13112
rect 14668 12980 14704 12981
rect 14516 12950 14525 12970
rect 14545 12950 14553 12970
rect 14404 12941 14460 12943
rect 14404 12940 14441 12941
rect 14516 12940 14553 12950
rect 14612 12970 14760 12980
rect 14860 12977 14956 12979
rect 14612 12950 14621 12970
rect 14641 12950 14731 12970
rect 14751 12950 14760 12970
rect 14612 12944 14760 12950
rect 14612 12941 14676 12944
rect 14612 12940 14649 12941
rect 14668 12914 14676 12941
rect 14697 12941 14760 12944
rect 14818 12970 14956 12977
rect 14818 12950 14827 12970
rect 14847 12950 14956 12970
rect 14818 12941 14956 12950
rect 14697 12914 14704 12941
rect 14723 12940 14760 12941
rect 14819 12940 14856 12941
rect 14668 12889 14704 12914
rect 14139 12887 14180 12888
rect 14005 12880 14180 12887
rect 13803 12854 13889 12873
rect 13803 12813 13818 12854
rect 13872 12813 13889 12854
rect 14005 12860 14149 12880
rect 14169 12860 14180 12880
rect 14005 12852 14180 12860
rect 14247 12884 14606 12888
rect 14247 12879 14569 12884
rect 14247 12855 14360 12879
rect 14384 12860 14569 12879
rect 14593 12860 14606 12884
rect 14384 12855 14606 12860
rect 14247 12852 14606 12855
rect 14668 12852 14703 12889
rect 14771 12886 14871 12889
rect 14771 12882 14838 12886
rect 14771 12856 14783 12882
rect 14809 12860 14838 12882
rect 14864 12860 14871 12886
rect 14809 12856 14871 12860
rect 14771 12852 14871 12856
rect 14005 12848 14051 12852
rect 14247 12831 14278 12852
rect 14668 12831 14704 12852
rect 14090 12830 14127 12831
rect 13803 12777 13889 12813
rect 14089 12821 14127 12830
rect 14089 12801 14098 12821
rect 14118 12801 14127 12821
rect 14089 12793 14127 12801
rect 14193 12825 14278 12831
rect 14303 12830 14340 12831
rect 14193 12805 14201 12825
rect 14221 12805 14278 12825
rect 14193 12797 14278 12805
rect 14302 12821 14340 12830
rect 14302 12801 14311 12821
rect 14331 12801 14340 12821
rect 14193 12796 14229 12797
rect 14302 12793 14340 12801
rect 14406 12825 14491 12831
rect 14511 12830 14548 12831
rect 14406 12805 14414 12825
rect 14434 12824 14491 12825
rect 14434 12805 14463 12824
rect 14406 12804 14463 12805
rect 14484 12804 14491 12824
rect 14406 12797 14491 12804
rect 14510 12821 14548 12830
rect 14510 12801 14519 12821
rect 14539 12801 14548 12821
rect 14406 12796 14442 12797
rect 14510 12793 14548 12801
rect 14614 12825 14758 12831
rect 14614 12805 14622 12825
rect 14642 12805 14730 12825
rect 14750 12805 14758 12825
rect 14614 12797 14758 12805
rect 14614 12796 14650 12797
rect 11259 12450 11323 12511
rect 11679 12509 11783 12511
rect 12014 12509 12055 12511
rect 12524 12508 12545 12553
rect 12525 12487 12545 12508
rect 12575 12508 12594 12553
rect 13631 12644 13711 12686
rect 12575 12487 12592 12508
rect 12525 12468 12592 12487
rect 12174 12460 12246 12461
rect 12173 12452 12272 12460
rect 7203 12204 7240 12235
rect 7416 12233 7452 12235
rect 7416 12204 7453 12233
rect 6655 12195 6690 12196
rect 6632 12190 6690 12195
rect 6632 12170 6635 12190
rect 6655 12176 6690 12190
rect 6710 12176 6719 12196
rect 6655 12168 6719 12176
rect 6681 12167 6719 12168
rect 6682 12166 6719 12167
rect 6785 12200 6821 12201
rect 6893 12200 6929 12201
rect 6785 12192 6929 12200
rect 6785 12172 6793 12192
rect 6813 12172 6901 12192
rect 6921 12172 6929 12192
rect 6785 12166 6929 12172
rect 6995 12196 7033 12204
rect 7101 12200 7137 12201
rect 6995 12176 7004 12196
rect 7024 12176 7033 12196
rect 6995 12167 7033 12176
rect 7052 12193 7137 12200
rect 7052 12173 7059 12193
rect 7080 12192 7137 12193
rect 7080 12173 7109 12192
rect 7052 12172 7109 12173
rect 7129 12172 7137 12192
rect 6995 12166 7032 12167
rect 7052 12166 7137 12172
rect 7203 12196 7241 12204
rect 7314 12200 7350 12201
rect 7203 12176 7212 12196
rect 7232 12176 7241 12196
rect 7203 12167 7241 12176
rect 7265 12192 7350 12200
rect 7265 12172 7322 12192
rect 7342 12172 7350 12192
rect 7203 12166 7240 12167
rect 7265 12166 7350 12172
rect 7416 12196 7454 12204
rect 7416 12176 7425 12196
rect 7445 12176 7454 12196
rect 7416 12167 7454 12176
rect 8941 12185 9021 12236
rect 7416 12166 7453 12167
rect 6839 12145 6875 12166
rect 7265 12145 7296 12166
rect 7476 12151 7533 12159
rect 7476 12145 7484 12151
rect 6672 12141 6772 12145
rect 6672 12137 6734 12141
rect 6672 12111 6679 12137
rect 6705 12115 6734 12137
rect 6760 12115 6772 12141
rect 6705 12111 6772 12115
rect 6672 12108 6772 12111
rect 6840 12108 6875 12145
rect 6937 12142 7296 12145
rect 6937 12137 7159 12142
rect 6937 12113 6950 12137
rect 6974 12118 7159 12137
rect 7183 12118 7296 12142
rect 6974 12113 7296 12118
rect 6937 12109 7296 12113
rect 7363 12137 7484 12145
rect 7363 12117 7374 12137
rect 7394 12128 7484 12137
rect 7510 12128 7533 12151
rect 7394 12117 7533 12128
rect 7363 12115 7533 12117
rect 7836 12144 7908 12164
rect 7836 12121 7864 12144
rect 7890 12121 7908 12144
rect 7363 12110 7484 12115
rect 7363 12109 7404 12110
rect 6839 12083 6875 12108
rect 6687 12056 6724 12057
rect 6783 12056 6820 12057
rect 6839 12056 6846 12083
rect 6587 12047 6725 12056
rect 6587 12027 6696 12047
rect 6716 12027 6725 12047
rect 6587 12020 6725 12027
rect 6783 12053 6846 12056
rect 6867 12056 6875 12083
rect 6894 12056 6931 12057
rect 6867 12053 6931 12056
rect 6783 12047 6931 12053
rect 6783 12027 6792 12047
rect 6812 12027 6902 12047
rect 6922 12027 6931 12047
rect 6587 12018 6683 12020
rect 6783 12017 6931 12027
rect 6990 12047 7027 12057
rect 7102 12056 7139 12057
rect 7083 12054 7139 12056
rect 6990 12027 6998 12047
rect 7018 12027 7027 12047
rect 6839 12016 6875 12017
rect 6687 11885 6724 11886
rect 6990 11885 7027 12027
rect 7052 12047 7139 12054
rect 7052 12044 7110 12047
rect 7052 12024 7057 12044
rect 7078 12027 7110 12044
rect 7130 12027 7139 12047
rect 7078 12024 7139 12027
rect 7052 12017 7139 12024
rect 7198 12047 7235 12057
rect 7198 12027 7206 12047
rect 7226 12027 7235 12047
rect 7052 12016 7083 12017
rect 7198 11948 7235 12027
rect 7265 12056 7296 12109
rect 7836 12059 7908 12121
rect 8941 12159 8957 12185
rect 8997 12159 9021 12185
rect 8941 12140 9021 12159
rect 8941 12114 8960 12140
rect 9000 12114 9021 12140
rect 8941 12087 9021 12114
rect 8941 12061 8964 12087
rect 9004 12061 9021 12087
rect 7315 12056 7352 12057
rect 7265 12047 7352 12056
rect 7265 12027 7323 12047
rect 7343 12027 7352 12047
rect 7265 12017 7352 12027
rect 7411 12047 7448 12057
rect 7411 12027 7419 12047
rect 7439 12027 7448 12047
rect 7265 12016 7296 12017
rect 7260 11948 7370 11961
rect 7411 11948 7448 12027
rect 7198 11946 7448 11948
rect 7198 11943 7299 11946
rect 7198 11924 7263 11943
rect 7260 11916 7263 11924
rect 7292 11916 7299 11943
rect 7327 11919 7337 11946
rect 7366 11924 7448 11946
rect 7366 11919 7370 11924
rect 7327 11916 7370 11919
rect 7260 11902 7370 11916
rect 6686 11884 7027 11885
rect 6611 11879 7027 11884
rect 6611 11859 6614 11879
rect 6634 11859 7028 11879
rect 6837 11826 6874 11836
rect 6837 11789 6846 11826
rect 6863 11789 6874 11826
rect 6837 11768 6874 11789
rect 6546 10829 6714 10830
rect 6843 10829 6872 11768
rect 6985 11154 7028 11859
rect 7840 11508 7902 12059
rect 8941 12050 9021 12061
rect 9083 12051 9110 12306
rect 9488 12298 9529 12448
rect 9760 12442 9864 12448
rect 10220 12445 10284 12448
rect 9955 12386 10076 12404
rect 9955 12384 10026 12386
rect 9955 12343 9970 12384
rect 10007 12345 10026 12384
rect 10063 12345 10076 12386
rect 10007 12343 10076 12345
rect 9955 12333 10076 12343
rect 9150 12191 9214 12203
rect 9490 12199 9527 12298
rect 9755 12288 9866 12301
rect 9755 12286 9797 12288
rect 9755 12266 9762 12286
rect 9781 12266 9797 12286
rect 9755 12258 9797 12266
rect 9825 12286 9866 12288
rect 9825 12266 9839 12286
rect 9858 12266 9866 12286
rect 9825 12258 9866 12266
rect 9755 12252 9866 12258
rect 9698 12230 9947 12252
rect 9698 12199 9735 12230
rect 9911 12228 9947 12230
rect 9911 12199 9948 12228
rect 9150 12190 9185 12191
rect 9127 12185 9185 12190
rect 9127 12165 9130 12185
rect 9150 12171 9185 12185
rect 9205 12171 9214 12191
rect 9150 12163 9214 12171
rect 9176 12162 9214 12163
rect 9177 12161 9214 12162
rect 9280 12195 9316 12196
rect 9388 12195 9424 12196
rect 9280 12187 9424 12195
rect 9280 12167 9288 12187
rect 9308 12167 9396 12187
rect 9416 12167 9424 12187
rect 9280 12161 9424 12167
rect 9490 12191 9528 12199
rect 9596 12195 9632 12196
rect 9490 12171 9499 12191
rect 9519 12171 9528 12191
rect 9490 12162 9528 12171
rect 9547 12188 9632 12195
rect 9547 12168 9554 12188
rect 9575 12187 9632 12188
rect 9575 12168 9604 12187
rect 9547 12167 9604 12168
rect 9624 12167 9632 12187
rect 9490 12161 9527 12162
rect 9547 12161 9632 12167
rect 9698 12191 9736 12199
rect 9809 12195 9845 12196
rect 9698 12171 9707 12191
rect 9727 12171 9736 12191
rect 9698 12162 9736 12171
rect 9760 12187 9845 12195
rect 9760 12167 9817 12187
rect 9837 12167 9845 12187
rect 9698 12161 9735 12162
rect 9760 12161 9845 12167
rect 9911 12191 9949 12199
rect 9911 12171 9920 12191
rect 9940 12171 9949 12191
rect 10004 12181 10069 12333
rect 10222 12307 10277 12445
rect 11261 12379 11320 12450
rect 12173 12449 12225 12452
rect 12173 12414 12181 12449
rect 12206 12414 12225 12449
rect 12250 12441 12272 12452
rect 12250 12440 13117 12441
rect 12250 12414 13118 12440
rect 12173 12404 13118 12414
rect 12173 12402 12272 12404
rect 11261 12361 11283 12379
rect 11301 12361 11320 12379
rect 11261 12339 11320 12361
rect 11528 12375 12060 12380
rect 11528 12355 12414 12375
rect 12434 12355 12437 12375
rect 13073 12371 13118 12404
rect 11528 12351 12437 12355
rect 9911 12162 9949 12171
rect 10002 12174 10069 12181
rect 9911 12161 9948 12162
rect 9334 12140 9370 12161
rect 9760 12140 9791 12161
rect 10002 12153 10019 12174
rect 10055 12153 10069 12174
rect 10221 12194 10277 12307
rect 11528 12304 11571 12351
rect 12021 12350 12437 12351
rect 13069 12351 13462 12371
rect 13482 12351 13485 12371
rect 12021 12349 12362 12350
rect 11678 12318 11788 12332
rect 11678 12315 11721 12318
rect 11678 12310 11682 12315
rect 11516 12303 11571 12304
rect 10221 12176 10240 12194
rect 10258 12176 10277 12194
rect 10221 12156 10277 12176
rect 11260 12280 11571 12303
rect 11260 12262 11285 12280
rect 11303 12268 11571 12280
rect 11600 12288 11682 12310
rect 11711 12288 11721 12315
rect 11749 12291 11756 12318
rect 11785 12310 11788 12318
rect 11785 12291 11850 12310
rect 11749 12288 11850 12291
rect 11600 12286 11850 12288
rect 11303 12262 11325 12268
rect 10002 12140 10069 12153
rect 9167 12136 9267 12140
rect 9167 12132 9229 12136
rect 9167 12106 9174 12132
rect 9200 12110 9229 12132
rect 9255 12110 9267 12136
rect 9200 12106 9267 12110
rect 9167 12103 9267 12106
rect 9335 12103 9370 12140
rect 9432 12137 9791 12140
rect 9432 12132 9654 12137
rect 9432 12108 9445 12132
rect 9469 12113 9654 12132
rect 9678 12113 9791 12137
rect 9469 12108 9791 12113
rect 9432 12104 9791 12108
rect 9858 12134 10069 12140
rect 9858 12132 10019 12134
rect 9858 12112 9869 12132
rect 9889 12112 10019 12132
rect 9858 12105 10019 12112
rect 9858 12104 9899 12105
rect 9334 12078 9370 12103
rect 9182 12051 9219 12052
rect 9278 12051 9315 12052
rect 9334 12051 9341 12078
rect 9082 12042 9220 12051
rect 9082 12022 9191 12042
rect 9211 12022 9220 12042
rect 9082 12015 9220 12022
rect 9278 12048 9341 12051
rect 9362 12051 9370 12078
rect 9389 12051 9426 12052
rect 9362 12048 9426 12051
rect 9278 12042 9426 12048
rect 9278 12022 9287 12042
rect 9307 12022 9397 12042
rect 9417 12022 9426 12042
rect 9082 12013 9178 12015
rect 9278 12012 9426 12022
rect 9485 12042 9522 12052
rect 9597 12051 9634 12052
rect 9578 12049 9634 12051
rect 9485 12022 9493 12042
rect 9513 12022 9522 12042
rect 9334 12011 9370 12012
rect 9182 11880 9219 11881
rect 9485 11880 9522 12022
rect 9547 12042 9634 12049
rect 9547 12039 9605 12042
rect 9547 12019 9552 12039
rect 9573 12022 9605 12039
rect 9625 12022 9634 12042
rect 9573 12019 9634 12022
rect 9547 12012 9634 12019
rect 9693 12042 9730 12052
rect 9693 12022 9701 12042
rect 9721 12022 9730 12042
rect 9547 12011 9578 12012
rect 9693 11943 9730 12022
rect 9760 12051 9791 12104
rect 10004 12097 10019 12105
rect 10059 12097 10069 12134
rect 11260 12123 11325 12262
rect 11600 12207 11637 12286
rect 11678 12273 11788 12286
rect 11752 12217 11783 12218
rect 11600 12187 11609 12207
rect 11629 12187 11637 12207
rect 10004 12088 10069 12097
rect 10217 12095 10282 12116
rect 10217 12077 10242 12095
rect 10260 12077 10282 12095
rect 11260 12105 11283 12123
rect 11301 12105 11325 12123
rect 11260 12088 11325 12105
rect 11480 12169 11548 12182
rect 11600 12177 11637 12187
rect 11696 12207 11783 12217
rect 11696 12187 11705 12207
rect 11725 12187 11783 12207
rect 11696 12178 11783 12187
rect 11696 12177 11733 12178
rect 11480 12127 11487 12169
rect 11536 12127 11548 12169
rect 11480 12124 11548 12127
rect 11752 12125 11783 12178
rect 11813 12207 11850 12286
rect 11965 12217 11996 12218
rect 11813 12187 11822 12207
rect 11842 12187 11850 12207
rect 11813 12177 11850 12187
rect 11909 12210 11996 12217
rect 11909 12207 11970 12210
rect 11909 12187 11918 12207
rect 11938 12190 11970 12207
rect 11991 12190 11996 12210
rect 11938 12187 11996 12190
rect 11909 12180 11996 12187
rect 12021 12207 12058 12349
rect 12324 12348 12361 12349
rect 13069 12346 13485 12351
rect 13069 12345 13410 12346
rect 12726 12314 12836 12328
rect 12726 12311 12769 12314
rect 12726 12306 12730 12311
rect 12648 12284 12730 12306
rect 12759 12284 12769 12311
rect 12797 12287 12804 12314
rect 12833 12306 12836 12314
rect 12833 12287 12898 12306
rect 12797 12284 12898 12287
rect 12648 12282 12898 12284
rect 12173 12217 12209 12218
rect 12021 12187 12030 12207
rect 12050 12187 12058 12207
rect 11909 12178 11965 12180
rect 11909 12177 11946 12178
rect 12021 12177 12058 12187
rect 12117 12207 12265 12217
rect 12365 12214 12461 12216
rect 12117 12187 12126 12207
rect 12146 12187 12236 12207
rect 12256 12187 12265 12207
rect 12117 12181 12265 12187
rect 12117 12178 12181 12181
rect 12117 12177 12154 12178
rect 12173 12151 12181 12178
rect 12202 12178 12265 12181
rect 12323 12207 12461 12214
rect 12323 12187 12332 12207
rect 12352 12187 12461 12207
rect 12323 12178 12461 12187
rect 12648 12203 12685 12282
rect 12726 12269 12836 12282
rect 12800 12213 12831 12214
rect 12648 12183 12657 12203
rect 12677 12183 12685 12203
rect 12202 12151 12209 12178
rect 12228 12177 12265 12178
rect 12324 12177 12361 12178
rect 12173 12126 12209 12151
rect 11644 12124 11685 12125
rect 11480 12117 11685 12124
rect 11480 12106 11654 12117
rect 9810 12051 9847 12052
rect 9760 12042 9847 12051
rect 9760 12022 9818 12042
rect 9838 12022 9847 12042
rect 9760 12012 9847 12022
rect 9906 12042 9943 12052
rect 9906 12022 9914 12042
rect 9934 12022 9943 12042
rect 9760 12011 9791 12012
rect 9755 11943 9865 11956
rect 9906 11943 9943 12022
rect 10217 12001 10282 12077
rect 11480 12073 11488 12106
rect 11481 12064 11488 12073
rect 11537 12097 11654 12106
rect 11674 12097 11685 12117
rect 11537 12089 11685 12097
rect 11752 12121 12111 12125
rect 11752 12116 12074 12121
rect 11752 12092 11865 12116
rect 11889 12097 12074 12116
rect 12098 12097 12111 12121
rect 11889 12092 12111 12097
rect 11752 12089 12111 12092
rect 12173 12089 12208 12126
rect 12276 12123 12376 12126
rect 12276 12119 12343 12123
rect 12276 12093 12288 12119
rect 12314 12097 12343 12119
rect 12369 12097 12376 12123
rect 12314 12093 12376 12097
rect 12276 12089 12376 12093
rect 11537 12073 11548 12089
rect 11537 12064 11545 12073
rect 11752 12068 11783 12089
rect 12173 12068 12209 12089
rect 11595 12067 11632 12068
rect 11260 12024 11325 12043
rect 11260 12006 11285 12024
rect 11303 12006 11325 12024
rect 9693 11941 9943 11943
rect 9693 11938 9794 11941
rect 9693 11919 9758 11938
rect 9755 11911 9758 11919
rect 9787 11911 9794 11938
rect 9822 11914 9832 11941
rect 9861 11919 9943 11941
rect 9966 11966 10283 12001
rect 9861 11914 9865 11919
rect 9822 11911 9865 11914
rect 9755 11897 9865 11911
rect 9181 11879 9522 11880
rect 9106 11877 9522 11879
rect 9966 11877 10006 11966
rect 10217 11939 10282 11966
rect 10217 11921 10240 11939
rect 10258 11921 10282 11939
rect 10217 11901 10282 11921
rect 9103 11874 10006 11877
rect 9103 11854 9109 11874
rect 9129 11854 10006 11874
rect 9103 11850 10006 11854
rect 9966 11847 10006 11850
rect 10218 11840 10283 11861
rect 8436 11832 9097 11833
rect 8436 11825 9370 11832
rect 8436 11824 9342 11825
rect 8436 11804 9287 11824
rect 9319 11805 9342 11824
rect 9367 11805 9370 11825
rect 9319 11804 9370 11805
rect 8436 11797 9370 11804
rect 8035 11755 8203 11756
rect 8438 11755 8477 11797
rect 9266 11795 9370 11797
rect 9335 11793 9370 11795
rect 10218 11822 10242 11840
rect 10260 11822 10283 11840
rect 10218 11775 10283 11822
rect 8035 11729 8479 11755
rect 8035 11727 8203 11729
rect 7837 11424 7906 11508
rect 6986 11146 7028 11154
rect 6986 11135 7031 11146
rect 6986 11097 6996 11135
rect 7021 11097 7031 11135
rect 6986 11088 7031 11097
rect 7835 10945 7906 11424
rect 8035 11376 8062 11727
rect 8438 11723 8479 11729
rect 8102 11516 8166 11528
rect 8442 11524 8479 11723
rect 8941 11750 9013 11767
rect 8941 11711 8949 11750
rect 8994 11711 9013 11750
rect 8707 11613 8818 11628
rect 8707 11611 8749 11613
rect 8707 11591 8714 11611
rect 8733 11591 8749 11611
rect 8707 11583 8749 11591
rect 8777 11611 8818 11613
rect 8777 11591 8791 11611
rect 8810 11591 8818 11611
rect 8777 11583 8818 11591
rect 8707 11577 8818 11583
rect 8650 11555 8899 11577
rect 8650 11524 8687 11555
rect 8863 11553 8899 11555
rect 8863 11524 8900 11553
rect 8102 11515 8137 11516
rect 8079 11510 8137 11515
rect 8079 11490 8082 11510
rect 8102 11496 8137 11510
rect 8157 11496 8166 11516
rect 8102 11488 8166 11496
rect 8128 11487 8166 11488
rect 8129 11486 8166 11487
rect 8232 11520 8268 11521
rect 8340 11520 8376 11521
rect 8232 11512 8376 11520
rect 8232 11492 8240 11512
rect 8260 11492 8348 11512
rect 8368 11492 8376 11512
rect 8232 11486 8376 11492
rect 8442 11516 8480 11524
rect 8548 11520 8584 11521
rect 8442 11496 8451 11516
rect 8471 11496 8480 11516
rect 8442 11487 8480 11496
rect 8499 11513 8584 11520
rect 8499 11493 8506 11513
rect 8527 11512 8584 11513
rect 8527 11493 8556 11512
rect 8499 11492 8556 11493
rect 8576 11492 8584 11512
rect 8442 11486 8479 11487
rect 8499 11486 8584 11492
rect 8650 11516 8688 11524
rect 8761 11520 8797 11521
rect 8650 11496 8659 11516
rect 8679 11496 8688 11516
rect 8650 11487 8688 11496
rect 8712 11512 8797 11520
rect 8712 11492 8769 11512
rect 8789 11492 8797 11512
rect 8650 11486 8687 11487
rect 8712 11486 8797 11492
rect 8863 11516 8901 11524
rect 8863 11496 8872 11516
rect 8892 11496 8901 11516
rect 8863 11487 8901 11496
rect 8941 11501 9013 11711
rect 9083 11745 10283 11775
rect 9083 11744 9527 11745
rect 9083 11742 9251 11744
rect 8941 11487 9024 11501
rect 8863 11486 8900 11487
rect 8286 11465 8322 11486
rect 8712 11465 8743 11486
rect 8941 11465 8958 11487
rect 8119 11461 8219 11465
rect 8119 11457 8181 11461
rect 8119 11431 8126 11457
rect 8152 11435 8181 11457
rect 8207 11435 8219 11461
rect 8152 11431 8219 11435
rect 8119 11428 8219 11431
rect 8287 11428 8322 11465
rect 8384 11462 8743 11465
rect 8384 11457 8606 11462
rect 8384 11433 8397 11457
rect 8421 11438 8606 11457
rect 8630 11438 8743 11462
rect 8421 11433 8743 11438
rect 8384 11429 8743 11433
rect 8810 11457 8958 11465
rect 8810 11437 8821 11457
rect 8841 11454 8958 11457
rect 9011 11454 9024 11487
rect 8841 11437 9024 11454
rect 8810 11430 9024 11437
rect 8810 11429 8851 11430
rect 8941 11429 9024 11430
rect 8286 11403 8322 11428
rect 8134 11376 8171 11377
rect 8230 11376 8267 11377
rect 8286 11376 8293 11403
rect 8034 11367 8172 11376
rect 8034 11347 8143 11367
rect 8163 11347 8172 11367
rect 8034 11340 8172 11347
rect 8230 11373 8293 11376
rect 8314 11376 8322 11403
rect 8341 11376 8378 11377
rect 8314 11373 8378 11376
rect 8230 11367 8378 11373
rect 8230 11347 8239 11367
rect 8259 11347 8349 11367
rect 8369 11347 8378 11367
rect 8034 11338 8130 11340
rect 8230 11337 8378 11347
rect 8437 11367 8474 11377
rect 8549 11376 8586 11377
rect 8530 11374 8586 11376
rect 8437 11347 8445 11367
rect 8465 11347 8474 11367
rect 8286 11336 8322 11337
rect 8134 11205 8171 11206
rect 8437 11205 8474 11347
rect 8499 11367 8586 11374
rect 8499 11364 8557 11367
rect 8499 11344 8504 11364
rect 8525 11347 8557 11364
rect 8577 11347 8586 11367
rect 8525 11344 8586 11347
rect 8499 11337 8586 11344
rect 8645 11367 8682 11377
rect 8645 11347 8653 11367
rect 8673 11347 8682 11367
rect 8499 11336 8530 11337
rect 8645 11268 8682 11347
rect 8712 11376 8743 11429
rect 8949 11396 8963 11429
rect 9016 11396 9024 11429
rect 8949 11390 9024 11396
rect 8949 11385 9019 11390
rect 8762 11376 8799 11377
rect 8712 11367 8799 11376
rect 8712 11347 8770 11367
rect 8790 11347 8799 11367
rect 8712 11337 8799 11347
rect 8858 11367 8895 11377
rect 9083 11372 9110 11742
rect 9150 11512 9214 11524
rect 9490 11520 9527 11744
rect 9998 11725 10062 11727
rect 9994 11713 10062 11725
rect 9994 11680 10005 11713
rect 10045 11680 10062 11713
rect 9994 11670 10062 11680
rect 9755 11609 9866 11624
rect 9755 11607 9797 11609
rect 9755 11587 9762 11607
rect 9781 11587 9797 11607
rect 9755 11579 9797 11587
rect 9825 11607 9866 11609
rect 9825 11587 9839 11607
rect 9858 11587 9866 11607
rect 9825 11579 9866 11587
rect 9755 11573 9866 11579
rect 9698 11551 9947 11573
rect 9698 11520 9735 11551
rect 9911 11549 9947 11551
rect 9911 11520 9948 11549
rect 9150 11511 9185 11512
rect 9127 11506 9185 11511
rect 9127 11486 9130 11506
rect 9150 11492 9185 11506
rect 9205 11492 9214 11512
rect 9150 11484 9214 11492
rect 9176 11483 9214 11484
rect 9177 11482 9214 11483
rect 9280 11516 9316 11517
rect 9388 11516 9424 11517
rect 9280 11508 9424 11516
rect 9280 11488 9288 11508
rect 9308 11488 9396 11508
rect 9416 11488 9424 11508
rect 9280 11482 9424 11488
rect 9490 11512 9528 11520
rect 9596 11516 9632 11517
rect 9490 11492 9499 11512
rect 9519 11492 9528 11512
rect 9490 11483 9528 11492
rect 9547 11509 9632 11516
rect 9547 11489 9554 11509
rect 9575 11508 9632 11509
rect 9575 11489 9604 11508
rect 9547 11488 9604 11489
rect 9624 11488 9632 11508
rect 9490 11482 9527 11483
rect 9547 11482 9632 11488
rect 9698 11512 9736 11520
rect 9809 11516 9845 11517
rect 9698 11492 9707 11512
rect 9727 11492 9736 11512
rect 9698 11483 9736 11492
rect 9760 11508 9845 11516
rect 9760 11488 9817 11508
rect 9837 11488 9845 11508
rect 9698 11482 9735 11483
rect 9760 11482 9845 11488
rect 9911 11512 9949 11520
rect 9911 11492 9920 11512
rect 9940 11492 9949 11512
rect 9911 11483 9949 11492
rect 9998 11486 10062 11670
rect 10218 11544 10283 11745
rect 11260 11805 11325 12006
rect 11481 11880 11545 12064
rect 11594 12058 11632 12067
rect 11594 12038 11603 12058
rect 11623 12038 11632 12058
rect 11594 12030 11632 12038
rect 11698 12062 11783 12068
rect 11808 12067 11845 12068
rect 11698 12042 11706 12062
rect 11726 12042 11783 12062
rect 11698 12034 11783 12042
rect 11807 12058 11845 12067
rect 11807 12038 11816 12058
rect 11836 12038 11845 12058
rect 11698 12033 11734 12034
rect 11807 12030 11845 12038
rect 11911 12062 11996 12068
rect 12016 12067 12053 12068
rect 11911 12042 11919 12062
rect 11939 12061 11996 12062
rect 11939 12042 11968 12061
rect 11911 12041 11968 12042
rect 11989 12041 11996 12061
rect 11911 12034 11996 12041
rect 12015 12058 12053 12067
rect 12015 12038 12024 12058
rect 12044 12038 12053 12058
rect 11911 12033 11947 12034
rect 12015 12030 12053 12038
rect 12119 12062 12263 12068
rect 12119 12042 12127 12062
rect 12147 12042 12235 12062
rect 12255 12042 12263 12062
rect 12119 12034 12263 12042
rect 12119 12033 12155 12034
rect 12227 12033 12263 12034
rect 12329 12067 12366 12068
rect 12329 12066 12367 12067
rect 12329 12058 12393 12066
rect 12329 12038 12338 12058
rect 12358 12044 12393 12058
rect 12413 12044 12416 12064
rect 12358 12039 12416 12044
rect 12358 12038 12393 12039
rect 11595 12001 11632 12030
rect 11596 11999 11632 12001
rect 11808 11999 11845 12030
rect 11596 11977 11845 11999
rect 11677 11971 11788 11977
rect 11677 11963 11718 11971
rect 11677 11943 11685 11963
rect 11704 11943 11718 11963
rect 11677 11941 11718 11943
rect 11746 11963 11788 11971
rect 11746 11943 11762 11963
rect 11781 11943 11788 11963
rect 11746 11941 11788 11943
rect 11677 11926 11788 11941
rect 11481 11870 11549 11880
rect 11481 11837 11498 11870
rect 11538 11837 11549 11870
rect 11481 11825 11549 11837
rect 11481 11823 11545 11825
rect 12016 11806 12053 12030
rect 12329 12026 12393 12038
rect 12433 11808 12460 12178
rect 12648 12173 12685 12183
rect 12744 12203 12831 12213
rect 12744 12183 12753 12203
rect 12773 12183 12831 12203
rect 12744 12174 12831 12183
rect 12744 12173 12781 12174
rect 12524 12160 12594 12165
rect 12519 12154 12594 12160
rect 12519 12121 12527 12154
rect 12580 12121 12594 12154
rect 12800 12121 12831 12174
rect 12861 12203 12898 12282
rect 13013 12213 13044 12214
rect 12861 12183 12870 12203
rect 12890 12183 12898 12203
rect 12861 12173 12898 12183
rect 12957 12206 13044 12213
rect 12957 12203 13018 12206
rect 12957 12183 12966 12203
rect 12986 12186 13018 12203
rect 13039 12186 13044 12206
rect 12986 12183 13044 12186
rect 12957 12176 13044 12183
rect 13069 12203 13106 12345
rect 13372 12344 13409 12345
rect 13221 12213 13257 12214
rect 13069 12183 13078 12203
rect 13098 12183 13106 12203
rect 12957 12174 13013 12176
rect 12957 12173 12994 12174
rect 13069 12173 13106 12183
rect 13165 12203 13313 12213
rect 13413 12210 13509 12212
rect 13165 12183 13174 12203
rect 13194 12183 13284 12203
rect 13304 12183 13313 12203
rect 13165 12177 13313 12183
rect 13165 12174 13229 12177
rect 13165 12173 13202 12174
rect 13221 12147 13229 12174
rect 13250 12174 13313 12177
rect 13371 12203 13509 12210
rect 13371 12183 13380 12203
rect 13400 12183 13509 12203
rect 13371 12174 13509 12183
rect 13250 12147 13257 12174
rect 13276 12173 13313 12174
rect 13372 12173 13409 12174
rect 13221 12122 13257 12147
rect 12519 12120 12602 12121
rect 12692 12120 12733 12121
rect 12519 12113 12733 12120
rect 12519 12096 12702 12113
rect 12519 12063 12532 12096
rect 12585 12093 12702 12096
rect 12722 12093 12733 12113
rect 12585 12085 12733 12093
rect 12800 12117 13159 12121
rect 12800 12112 13122 12117
rect 12800 12088 12913 12112
rect 12937 12093 13122 12112
rect 13146 12093 13159 12117
rect 12937 12088 13159 12093
rect 12800 12085 13159 12088
rect 13221 12085 13256 12122
rect 13324 12119 13424 12122
rect 13324 12115 13391 12119
rect 13324 12089 13336 12115
rect 13362 12093 13391 12115
rect 13417 12093 13424 12119
rect 13362 12089 13424 12093
rect 13324 12085 13424 12089
rect 12585 12063 12602 12085
rect 12800 12064 12831 12085
rect 13221 12064 13257 12085
rect 12643 12063 12680 12064
rect 12519 12049 12602 12063
rect 12292 11806 12460 11808
rect 12016 11805 12460 11806
rect 11260 11775 12460 11805
rect 12530 11839 12602 12049
rect 12642 12054 12680 12063
rect 12642 12034 12651 12054
rect 12671 12034 12680 12054
rect 12642 12026 12680 12034
rect 12746 12058 12831 12064
rect 12856 12063 12893 12064
rect 12746 12038 12754 12058
rect 12774 12038 12831 12058
rect 12746 12030 12831 12038
rect 12855 12054 12893 12063
rect 12855 12034 12864 12054
rect 12884 12034 12893 12054
rect 12746 12029 12782 12030
rect 12855 12026 12893 12034
rect 12959 12058 13044 12064
rect 13064 12063 13101 12064
rect 12959 12038 12967 12058
rect 12987 12057 13044 12058
rect 12987 12038 13016 12057
rect 12959 12037 13016 12038
rect 13037 12037 13044 12057
rect 12959 12030 13044 12037
rect 13063 12054 13101 12063
rect 13063 12034 13072 12054
rect 13092 12034 13101 12054
rect 12959 12029 12995 12030
rect 13063 12026 13101 12034
rect 13167 12058 13311 12064
rect 13167 12038 13175 12058
rect 13195 12038 13283 12058
rect 13303 12038 13311 12058
rect 13167 12030 13311 12038
rect 13167 12029 13203 12030
rect 13275 12029 13311 12030
rect 13377 12063 13414 12064
rect 13377 12062 13415 12063
rect 13377 12054 13441 12062
rect 13377 12034 13386 12054
rect 13406 12040 13441 12054
rect 13461 12040 13464 12060
rect 13406 12035 13464 12040
rect 13406 12034 13441 12035
rect 12643 11997 12680 12026
rect 12644 11995 12680 11997
rect 12856 11995 12893 12026
rect 12644 11973 12893 11995
rect 12725 11967 12836 11973
rect 12725 11959 12766 11967
rect 12725 11939 12733 11959
rect 12752 11939 12766 11959
rect 12725 11937 12766 11939
rect 12794 11959 12836 11967
rect 12794 11939 12810 11959
rect 12829 11939 12836 11959
rect 12794 11937 12836 11939
rect 12725 11922 12836 11937
rect 12530 11800 12549 11839
rect 12594 11800 12602 11839
rect 12530 11783 12602 11800
rect 13064 11827 13101 12026
rect 13377 12022 13441 12034
rect 13064 11821 13105 11827
rect 13481 11823 13508 12174
rect 13631 12044 13710 12644
rect 13807 12192 13886 12777
rect 14090 12764 14127 12793
rect 14091 12762 14127 12764
rect 14303 12762 14340 12793
rect 14091 12740 14340 12762
rect 14172 12734 14283 12740
rect 14172 12726 14213 12734
rect 14172 12706 14180 12726
rect 14199 12706 14213 12726
rect 14172 12704 14213 12706
rect 14241 12726 14283 12734
rect 14241 12706 14257 12726
rect 14276 12706 14283 12726
rect 14241 12704 14283 12706
rect 14172 12689 14283 12704
rect 14511 12678 14548 12793
rect 14504 12566 14551 12678
rect 14672 12638 14702 12797
rect 14722 12796 14758 12797
rect 14824 12830 14861 12831
rect 14824 12829 14862 12830
rect 14824 12821 14888 12829
rect 14824 12801 14833 12821
rect 14853 12807 14888 12821
rect 14908 12807 14911 12827
rect 14853 12802 14911 12807
rect 14853 12801 14888 12802
rect 14824 12789 14888 12801
rect 14672 12634 14758 12638
rect 14672 12616 14687 12634
rect 14739 12616 14758 12634
rect 14672 12607 14758 12616
rect 14928 12568 14955 12941
rect 14787 12566 14955 12568
rect 14504 12540 14955 12566
rect 14504 12462 14551 12540
rect 14787 12539 14955 12540
rect 14449 12461 14551 12462
rect 14448 12453 14551 12461
rect 14448 12450 14500 12453
rect 14448 12415 14456 12450
rect 14481 12415 14500 12450
rect 14525 12415 14551 12453
rect 14448 12409 14551 12415
rect 14711 12454 14747 12458
rect 14711 12431 14719 12454
rect 14743 12431 14747 12454
rect 14711 12410 14747 12431
rect 14448 12405 14547 12409
rect 14711 12387 14719 12410
rect 14743 12387 14747 12410
rect 13340 11821 13508 11823
rect 13064 11795 13508 11821
rect 11260 11728 11325 11775
rect 11260 11710 11283 11728
rect 11301 11710 11325 11728
rect 12173 11755 12208 11757
rect 12173 11753 12277 11755
rect 13066 11753 13105 11795
rect 13340 11794 13508 11795
rect 12173 11746 13107 11753
rect 12173 11745 12224 11746
rect 12173 11725 12176 11745
rect 12201 11726 12224 11745
rect 12256 11726 13107 11746
rect 12201 11725 13107 11726
rect 12173 11718 13107 11725
rect 12446 11717 13107 11718
rect 11260 11689 11325 11710
rect 11537 11700 11577 11703
rect 11537 11696 12440 11700
rect 11537 11676 12414 11696
rect 12434 11676 12440 11696
rect 11537 11673 12440 11676
rect 11261 11629 11326 11649
rect 11261 11611 11285 11629
rect 11303 11611 11326 11629
rect 11261 11584 11326 11611
rect 11537 11584 11577 11673
rect 12021 11671 12437 11673
rect 12021 11670 12362 11671
rect 11678 11639 11788 11653
rect 11678 11636 11721 11639
rect 11678 11631 11682 11636
rect 11260 11549 11577 11584
rect 11600 11609 11682 11631
rect 11711 11609 11721 11636
rect 11749 11612 11756 11639
rect 11785 11631 11788 11639
rect 11785 11612 11850 11631
rect 11749 11609 11850 11612
rect 11600 11607 11850 11609
rect 10218 11526 10240 11544
rect 10258 11526 10283 11544
rect 10218 11507 10283 11526
rect 9911 11482 9948 11483
rect 9334 11461 9370 11482
rect 9760 11461 9791 11482
rect 9998 11477 10006 11486
rect 9995 11461 10006 11477
rect 9167 11457 9267 11461
rect 9167 11453 9229 11457
rect 9167 11427 9174 11453
rect 9200 11431 9229 11453
rect 9255 11431 9267 11457
rect 9200 11427 9267 11431
rect 9167 11424 9267 11427
rect 9335 11424 9370 11461
rect 9432 11458 9791 11461
rect 9432 11453 9654 11458
rect 9432 11429 9445 11453
rect 9469 11434 9654 11453
rect 9678 11434 9791 11458
rect 9469 11429 9791 11434
rect 9432 11425 9791 11429
rect 9858 11453 10006 11461
rect 9858 11433 9869 11453
rect 9889 11444 10006 11453
rect 10055 11477 10062 11486
rect 10055 11444 10063 11477
rect 11261 11473 11326 11549
rect 11600 11528 11637 11607
rect 11678 11594 11788 11607
rect 11752 11538 11783 11539
rect 11600 11508 11609 11528
rect 11629 11508 11637 11528
rect 11600 11498 11637 11508
rect 11696 11528 11783 11538
rect 11696 11508 11705 11528
rect 11725 11508 11783 11528
rect 11696 11499 11783 11508
rect 11696 11498 11733 11499
rect 9889 11433 10063 11444
rect 9858 11426 10063 11433
rect 9858 11425 9899 11426
rect 9334 11399 9370 11424
rect 9182 11372 9219 11373
rect 9278 11372 9315 11373
rect 9334 11372 9341 11399
rect 8858 11347 8866 11367
rect 8886 11347 8895 11367
rect 8712 11336 8743 11337
rect 8707 11268 8817 11281
rect 8858 11268 8895 11347
rect 9082 11363 9220 11372
rect 9082 11343 9191 11363
rect 9211 11343 9220 11363
rect 9082 11336 9220 11343
rect 9278 11369 9341 11372
rect 9362 11372 9370 11399
rect 9389 11372 9426 11373
rect 9362 11369 9426 11372
rect 9278 11363 9426 11369
rect 9278 11343 9287 11363
rect 9307 11343 9397 11363
rect 9417 11343 9426 11363
rect 9082 11334 9178 11336
rect 9278 11333 9426 11343
rect 9485 11363 9522 11373
rect 9597 11372 9634 11373
rect 9578 11370 9634 11372
rect 9485 11343 9493 11363
rect 9513 11343 9522 11363
rect 9334 11332 9370 11333
rect 8645 11266 8895 11268
rect 8645 11263 8746 11266
rect 8645 11244 8710 11263
rect 8707 11236 8710 11244
rect 8739 11236 8746 11263
rect 8774 11239 8784 11266
rect 8813 11244 8895 11266
rect 8813 11239 8817 11244
rect 8774 11236 8817 11239
rect 8707 11222 8817 11236
rect 8133 11204 8474 11205
rect 8058 11199 8474 11204
rect 9182 11201 9219 11202
rect 9485 11201 9522 11343
rect 9547 11363 9634 11370
rect 9547 11360 9605 11363
rect 9547 11340 9552 11360
rect 9573 11343 9605 11360
rect 9625 11343 9634 11363
rect 9573 11340 9634 11343
rect 9547 11333 9634 11340
rect 9693 11363 9730 11373
rect 9693 11343 9701 11363
rect 9721 11343 9730 11363
rect 9547 11332 9578 11333
rect 9693 11264 9730 11343
rect 9760 11372 9791 11425
rect 9995 11423 10063 11426
rect 9995 11381 10007 11423
rect 10056 11381 10063 11423
rect 9810 11372 9847 11373
rect 9760 11363 9847 11372
rect 9760 11343 9818 11363
rect 9838 11343 9847 11363
rect 9760 11333 9847 11343
rect 9906 11363 9943 11373
rect 9995 11368 10063 11381
rect 10218 11445 10283 11462
rect 10218 11427 10242 11445
rect 10260 11427 10283 11445
rect 11261 11455 11283 11473
rect 11301 11455 11326 11473
rect 11261 11434 11326 11455
rect 11474 11453 11539 11462
rect 9906 11343 9914 11363
rect 9934 11343 9943 11363
rect 9760 11332 9791 11333
rect 9755 11264 9865 11277
rect 9906 11264 9943 11343
rect 10218 11288 10283 11427
rect 11474 11416 11484 11453
rect 11524 11445 11539 11453
rect 11752 11446 11783 11499
rect 11813 11528 11850 11607
rect 11965 11538 11996 11539
rect 11813 11508 11822 11528
rect 11842 11508 11850 11528
rect 11813 11498 11850 11508
rect 11909 11531 11996 11538
rect 11909 11528 11970 11531
rect 11909 11508 11918 11528
rect 11938 11511 11970 11528
rect 11991 11511 11996 11531
rect 11938 11508 11996 11511
rect 11909 11501 11996 11508
rect 12021 11528 12058 11670
rect 12324 11669 12361 11670
rect 12173 11538 12209 11539
rect 12021 11508 12030 11528
rect 12050 11508 12058 11528
rect 11909 11499 11965 11501
rect 11909 11498 11946 11499
rect 12021 11498 12058 11508
rect 12117 11528 12265 11538
rect 12365 11535 12461 11537
rect 12117 11508 12126 11528
rect 12146 11508 12236 11528
rect 12256 11508 12265 11528
rect 12117 11502 12265 11508
rect 12117 11499 12181 11502
rect 12117 11498 12154 11499
rect 12173 11472 12181 11499
rect 12202 11499 12265 11502
rect 12323 11528 12461 11535
rect 12323 11508 12332 11528
rect 12352 11508 12461 11528
rect 12323 11499 12461 11508
rect 12202 11472 12209 11499
rect 12228 11498 12265 11499
rect 12324 11498 12361 11499
rect 12173 11447 12209 11472
rect 11644 11445 11685 11446
rect 11524 11438 11685 11445
rect 11524 11418 11654 11438
rect 11674 11418 11685 11438
rect 11524 11416 11685 11418
rect 11474 11410 11685 11416
rect 11752 11442 12111 11446
rect 11752 11437 12074 11442
rect 11752 11413 11865 11437
rect 11889 11418 12074 11437
rect 12098 11418 12111 11442
rect 11889 11413 12111 11418
rect 11752 11410 12111 11413
rect 12173 11410 12208 11447
rect 12276 11444 12376 11447
rect 12276 11440 12343 11444
rect 12276 11414 12288 11440
rect 12314 11418 12343 11440
rect 12369 11418 12376 11444
rect 12314 11414 12376 11418
rect 12276 11410 12376 11414
rect 11474 11397 11541 11410
rect 10218 11282 10240 11288
rect 9693 11262 9943 11264
rect 9693 11259 9794 11262
rect 9693 11240 9758 11259
rect 9755 11232 9758 11240
rect 9787 11232 9794 11259
rect 9822 11235 9832 11262
rect 9861 11240 9943 11262
rect 9972 11270 10240 11282
rect 10258 11270 10283 11288
rect 9972 11247 10283 11270
rect 11266 11374 11322 11394
rect 11266 11356 11285 11374
rect 11303 11356 11322 11374
rect 9972 11246 10027 11247
rect 9861 11235 9865 11240
rect 9822 11232 9865 11235
rect 9755 11218 9865 11232
rect 9181 11200 9522 11201
rect 8058 11179 8061 11199
rect 8081 11179 8474 11199
rect 9106 11199 9522 11200
rect 9972 11199 10015 11246
rect 11266 11243 11322 11356
rect 11474 11376 11488 11397
rect 11524 11376 11541 11397
rect 11752 11389 11783 11410
rect 12173 11389 12209 11410
rect 11595 11388 11632 11389
rect 11474 11369 11541 11376
rect 11594 11379 11632 11388
rect 9106 11195 10015 11199
rect 8425 11146 8470 11179
rect 9106 11175 9109 11195
rect 9129 11175 10015 11195
rect 9483 11170 10015 11175
rect 10223 11189 10282 11211
rect 10223 11171 10242 11189
rect 10260 11171 10282 11189
rect 9271 11146 9370 11148
rect 8425 11136 9370 11146
rect 8425 11110 9293 11136
rect 8426 11109 9293 11110
rect 9271 11098 9293 11109
rect 9318 11101 9337 11136
rect 9362 11101 9370 11136
rect 9318 11098 9370 11101
rect 9271 11090 9370 11098
rect 9297 11089 9369 11090
rect 10223 11041 10282 11171
rect 11266 11114 11321 11243
rect 11474 11217 11539 11369
rect 11594 11359 11603 11379
rect 11623 11359 11632 11379
rect 11594 11351 11632 11359
rect 11698 11383 11783 11389
rect 11808 11388 11845 11389
rect 11698 11363 11706 11383
rect 11726 11363 11783 11383
rect 11698 11355 11783 11363
rect 11807 11379 11845 11388
rect 11807 11359 11816 11379
rect 11836 11359 11845 11379
rect 11698 11354 11734 11355
rect 11807 11351 11845 11359
rect 11911 11383 11996 11389
rect 12016 11388 12053 11389
rect 11911 11363 11919 11383
rect 11939 11382 11996 11383
rect 11939 11363 11968 11382
rect 11911 11362 11968 11363
rect 11989 11362 11996 11382
rect 11911 11355 11996 11362
rect 12015 11379 12053 11388
rect 12015 11359 12024 11379
rect 12044 11359 12053 11379
rect 11911 11354 11947 11355
rect 12015 11351 12053 11359
rect 12119 11383 12263 11389
rect 12119 11363 12127 11383
rect 12147 11363 12235 11383
rect 12255 11363 12263 11383
rect 12119 11355 12263 11363
rect 12119 11354 12155 11355
rect 12227 11354 12263 11355
rect 12329 11388 12366 11389
rect 12329 11387 12367 11388
rect 12329 11379 12393 11387
rect 12329 11359 12338 11379
rect 12358 11365 12393 11379
rect 12413 11365 12416 11385
rect 12358 11360 12416 11365
rect 12358 11359 12393 11360
rect 11595 11322 11632 11351
rect 11596 11320 11632 11322
rect 11808 11320 11845 11351
rect 11596 11298 11845 11320
rect 11677 11292 11788 11298
rect 11677 11284 11718 11292
rect 11677 11264 11685 11284
rect 11704 11264 11718 11284
rect 11677 11262 11718 11264
rect 11746 11284 11788 11292
rect 11746 11264 11762 11284
rect 11781 11264 11788 11284
rect 11746 11262 11788 11264
rect 11677 11247 11788 11262
rect 12016 11252 12053 11351
rect 12329 11347 12393 11359
rect 11679 11238 11783 11247
rect 11467 11207 11588 11217
rect 11467 11205 11536 11207
rect 11467 11164 11480 11205
rect 11517 11166 11536 11205
rect 11573 11166 11588 11207
rect 11517 11164 11588 11166
rect 11467 11146 11588 11164
rect 11260 11102 11321 11114
rect 12014 11102 12055 11252
rect 12433 11244 12460 11499
rect 12522 11489 12602 11500
rect 12522 11463 12539 11489
rect 12579 11463 12602 11489
rect 12522 11436 12602 11463
rect 12522 11410 12543 11436
rect 12583 11410 12602 11436
rect 12522 11391 12602 11410
rect 12522 11365 12546 11391
rect 12586 11365 12602 11391
rect 12522 11314 12602 11365
rect 11260 11099 12055 11102
rect 12434 11113 12460 11244
rect 12524 11158 12594 11314
rect 12523 11142 12599 11158
rect 12434 11099 12462 11113
rect 11260 11064 12462 11099
rect 12523 11105 12538 11142
rect 12582 11105 12599 11142
rect 12523 11085 12599 11105
rect 13637 11135 13707 12044
rect 13806 11479 13887 12192
rect 14711 12078 14747 12387
rect 14635 12049 14748 12078
rect 14635 11693 14666 12049
rect 14705 11794 15696 11819
rect 14705 11789 14765 11794
rect 14705 11768 14724 11789
rect 14744 11773 14765 11789
rect 14785 11773 15696 11794
rect 14744 11768 15696 11773
rect 14705 11760 15696 11768
rect 14710 11737 14816 11760
rect 14710 11734 14815 11737
rect 14559 11673 14952 11693
rect 14972 11673 14975 11693
rect 14559 11668 14975 11673
rect 14559 11667 14900 11668
rect 14216 11636 14326 11650
rect 14216 11633 14259 11636
rect 14216 11628 14220 11633
rect 14138 11606 14220 11628
rect 14249 11606 14259 11633
rect 14287 11609 14294 11636
rect 14323 11628 14326 11636
rect 14323 11609 14388 11628
rect 14287 11606 14388 11609
rect 14138 11604 14388 11606
rect 14138 11525 14175 11604
rect 14216 11591 14326 11604
rect 14290 11535 14321 11536
rect 14138 11505 14147 11525
rect 14167 11505 14175 11525
rect 14138 11495 14175 11505
rect 14234 11525 14321 11535
rect 14234 11505 14243 11525
rect 14263 11505 14321 11525
rect 14234 11496 14321 11505
rect 14234 11495 14271 11496
rect 13804 11443 13896 11479
rect 14290 11443 14321 11496
rect 14351 11525 14388 11604
rect 14503 11535 14534 11536
rect 14351 11505 14360 11525
rect 14380 11505 14388 11525
rect 14351 11495 14388 11505
rect 14447 11528 14534 11535
rect 14447 11525 14508 11528
rect 14447 11505 14456 11525
rect 14476 11508 14508 11525
rect 14529 11508 14534 11528
rect 14476 11505 14534 11508
rect 14447 11498 14534 11505
rect 14559 11525 14596 11667
rect 14862 11666 14899 11667
rect 14711 11535 14747 11536
rect 14559 11505 14568 11525
rect 14588 11505 14596 11525
rect 14447 11496 14503 11498
rect 14447 11495 14484 11496
rect 14559 11495 14596 11505
rect 14655 11525 14803 11535
rect 14903 11532 14999 11534
rect 14655 11505 14664 11525
rect 14684 11505 14774 11525
rect 14794 11505 14803 11525
rect 14655 11499 14803 11505
rect 14655 11496 14719 11499
rect 14655 11495 14692 11496
rect 14711 11469 14719 11496
rect 14740 11496 14803 11499
rect 14861 11525 14999 11532
rect 14861 11505 14870 11525
rect 14890 11505 14999 11525
rect 14861 11496 14999 11505
rect 14740 11469 14747 11496
rect 14766 11495 14803 11496
rect 14862 11495 14899 11496
rect 14711 11444 14747 11469
rect 13804 11442 14140 11443
rect 14182 11442 14223 11443
rect 13804 11435 14223 11442
rect 13804 11415 14192 11435
rect 14212 11415 14223 11435
rect 13804 11407 14223 11415
rect 14290 11439 14649 11443
rect 14290 11434 14612 11439
rect 14290 11410 14403 11434
rect 14427 11415 14612 11434
rect 14636 11415 14649 11439
rect 14427 11410 14649 11415
rect 14290 11407 14649 11410
rect 14711 11407 14746 11444
rect 14814 11441 14914 11444
rect 14814 11437 14881 11441
rect 14814 11411 14826 11437
rect 14852 11415 14881 11437
rect 14907 11415 14914 11441
rect 14852 11411 14914 11415
rect 14814 11407 14914 11411
rect 13804 11403 14140 11407
rect 13637 11085 13709 11135
rect 8945 11011 9021 11035
rect 8945 10945 8957 11011
rect 9011 10945 9021 11011
rect 9489 10966 9530 10968
rect 9761 10966 9865 10968
rect 10223 10966 10284 11041
rect 11260 10989 11321 11064
rect 11679 11062 11783 11064
rect 12014 11062 12055 11064
rect 12523 11019 12533 11085
rect 12587 11019 12599 11085
rect 12523 10995 12599 11019
rect 7835 10895 7907 10945
rect 6546 10803 6990 10829
rect 6546 10801 6714 10803
rect 6546 10534 6573 10801
rect 6843 10799 6872 10803
rect 6613 10674 6677 10686
rect 6953 10682 6990 10803
rect 7218 10771 7329 10786
rect 7218 10769 7260 10771
rect 7218 10749 7225 10769
rect 7244 10749 7260 10769
rect 7218 10741 7260 10749
rect 7288 10769 7329 10771
rect 7288 10749 7302 10769
rect 7321 10749 7329 10769
rect 7288 10741 7329 10749
rect 7218 10735 7329 10741
rect 7161 10713 7410 10735
rect 7161 10682 7198 10713
rect 7374 10711 7410 10713
rect 7374 10682 7411 10711
rect 6613 10673 6648 10674
rect 6590 10668 6648 10673
rect 6590 10648 6593 10668
rect 6613 10654 6648 10668
rect 6668 10654 6677 10674
rect 6613 10646 6677 10654
rect 6639 10645 6677 10646
rect 6640 10644 6677 10645
rect 6743 10678 6779 10679
rect 6851 10678 6887 10679
rect 6743 10670 6887 10678
rect 6743 10650 6751 10670
rect 6771 10650 6859 10670
rect 6879 10650 6887 10670
rect 6743 10644 6887 10650
rect 6953 10674 6991 10682
rect 7059 10678 7095 10679
rect 6953 10654 6962 10674
rect 6982 10654 6991 10674
rect 6953 10645 6991 10654
rect 7010 10671 7095 10678
rect 7010 10651 7017 10671
rect 7038 10670 7095 10671
rect 7038 10651 7067 10670
rect 7010 10650 7067 10651
rect 7087 10650 7095 10670
rect 6953 10644 6990 10645
rect 7010 10644 7095 10650
rect 7161 10674 7199 10682
rect 7272 10678 7308 10679
rect 7161 10654 7170 10674
rect 7190 10654 7199 10674
rect 7161 10645 7199 10654
rect 7223 10670 7308 10678
rect 7223 10650 7280 10670
rect 7300 10650 7308 10670
rect 7161 10644 7198 10645
rect 7223 10644 7308 10650
rect 7374 10674 7412 10682
rect 7374 10654 7383 10674
rect 7403 10654 7412 10674
rect 7374 10645 7412 10654
rect 7374 10644 7411 10645
rect 6797 10623 6833 10644
rect 7223 10623 7254 10644
rect 7404 10623 7738 10627
rect 6630 10619 6730 10623
rect 6630 10615 6692 10619
rect 6630 10589 6637 10615
rect 6663 10593 6692 10615
rect 6718 10593 6730 10619
rect 6663 10589 6730 10593
rect 6630 10586 6730 10589
rect 6798 10586 6833 10623
rect 6895 10620 7254 10623
rect 6895 10615 7117 10620
rect 6895 10591 6908 10615
rect 6932 10596 7117 10615
rect 7141 10596 7254 10620
rect 6932 10591 7254 10596
rect 6895 10587 7254 10591
rect 7321 10615 7738 10623
rect 7321 10595 7332 10615
rect 7352 10595 7738 10615
rect 7321 10588 7738 10595
rect 7321 10587 7362 10588
rect 7404 10587 7738 10588
rect 6797 10561 6833 10586
rect 6645 10534 6682 10535
rect 6741 10534 6778 10535
rect 6797 10534 6804 10561
rect 6545 10525 6683 10534
rect 6545 10505 6654 10525
rect 6674 10505 6683 10525
rect 6545 10498 6683 10505
rect 6741 10531 6804 10534
rect 6825 10534 6833 10561
rect 6852 10534 6889 10535
rect 6825 10531 6889 10534
rect 6741 10525 6889 10531
rect 6741 10505 6750 10525
rect 6770 10505 6860 10525
rect 6880 10505 6889 10525
rect 6545 10496 6641 10498
rect 6741 10495 6889 10505
rect 6948 10525 6985 10535
rect 7060 10534 7097 10535
rect 7041 10532 7097 10534
rect 6948 10505 6956 10525
rect 6976 10505 6985 10525
rect 6797 10494 6833 10495
rect 6645 10363 6682 10364
rect 6948 10363 6985 10505
rect 7010 10525 7097 10532
rect 7010 10522 7068 10525
rect 7010 10502 7015 10522
rect 7036 10505 7068 10522
rect 7088 10505 7097 10525
rect 7036 10502 7097 10505
rect 7010 10495 7097 10502
rect 7156 10525 7193 10535
rect 7156 10505 7164 10525
rect 7184 10505 7193 10525
rect 7010 10494 7041 10495
rect 7156 10426 7193 10505
rect 7223 10534 7254 10587
rect 7273 10534 7310 10535
rect 7223 10525 7310 10534
rect 7223 10505 7281 10525
rect 7301 10505 7310 10525
rect 7223 10495 7310 10505
rect 7369 10525 7406 10535
rect 7369 10505 7377 10525
rect 7397 10505 7406 10525
rect 7223 10494 7254 10495
rect 7218 10426 7328 10439
rect 7369 10426 7406 10505
rect 7156 10424 7406 10426
rect 7156 10421 7257 10424
rect 7156 10402 7221 10421
rect 7218 10394 7221 10402
rect 7250 10394 7257 10421
rect 7285 10397 7295 10424
rect 7324 10402 7406 10424
rect 7324 10397 7328 10402
rect 7285 10394 7328 10397
rect 7218 10380 7328 10394
rect 6644 10362 6985 10363
rect 6569 10357 6985 10362
rect 6569 10337 6572 10357
rect 6592 10337 6985 10357
rect 6878 9972 6909 10337
rect 6796 9943 6909 9972
rect 6797 9643 6833 9943
rect 7657 9838 7738 10587
rect 7837 9986 7907 10895
rect 8945 10925 9021 10945
rect 8945 10888 8962 10925
rect 9006 10888 9021 10925
rect 9082 10931 10284 10966
rect 9082 10917 9110 10931
rect 8945 10872 9021 10888
rect 8950 10716 9020 10872
rect 9084 10786 9110 10917
rect 9489 10928 10284 10931
rect 8942 10665 9022 10716
rect 8942 10639 8958 10665
rect 8998 10639 9022 10665
rect 8942 10620 9022 10639
rect 8942 10594 8961 10620
rect 9001 10594 9022 10620
rect 8942 10567 9022 10594
rect 8942 10541 8965 10567
rect 9005 10541 9022 10567
rect 8942 10530 9022 10541
rect 9084 10531 9111 10786
rect 9489 10778 9530 10928
rect 10223 10916 10284 10928
rect 9956 10866 10077 10884
rect 9956 10864 10027 10866
rect 9956 10823 9971 10864
rect 10008 10825 10027 10864
rect 10064 10825 10077 10866
rect 10008 10823 10077 10825
rect 9956 10813 10077 10823
rect 9761 10783 9865 10792
rect 9151 10671 9215 10683
rect 9491 10679 9528 10778
rect 9756 10768 9867 10783
rect 9756 10766 9798 10768
rect 9756 10746 9763 10766
rect 9782 10746 9798 10766
rect 9756 10738 9798 10746
rect 9826 10766 9867 10768
rect 9826 10746 9840 10766
rect 9859 10746 9867 10766
rect 9826 10738 9867 10746
rect 9756 10732 9867 10738
rect 9699 10710 9948 10732
rect 9699 10679 9736 10710
rect 9912 10708 9948 10710
rect 9912 10679 9949 10708
rect 9151 10670 9186 10671
rect 9128 10665 9186 10670
rect 9128 10645 9131 10665
rect 9151 10651 9186 10665
rect 9206 10651 9215 10671
rect 9151 10643 9215 10651
rect 9177 10642 9215 10643
rect 9178 10641 9215 10642
rect 9281 10675 9317 10676
rect 9389 10675 9425 10676
rect 9281 10667 9425 10675
rect 9281 10647 9289 10667
rect 9309 10647 9397 10667
rect 9417 10647 9425 10667
rect 9281 10641 9425 10647
rect 9491 10671 9529 10679
rect 9597 10675 9633 10676
rect 9491 10651 9500 10671
rect 9520 10651 9529 10671
rect 9491 10642 9529 10651
rect 9548 10668 9633 10675
rect 9548 10648 9555 10668
rect 9576 10667 9633 10668
rect 9576 10648 9605 10667
rect 9548 10647 9605 10648
rect 9625 10647 9633 10667
rect 9491 10641 9528 10642
rect 9548 10641 9633 10647
rect 9699 10671 9737 10679
rect 9810 10675 9846 10676
rect 9699 10651 9708 10671
rect 9728 10651 9737 10671
rect 9699 10642 9737 10651
rect 9761 10667 9846 10675
rect 9761 10647 9818 10667
rect 9838 10647 9846 10667
rect 9699 10641 9736 10642
rect 9761 10641 9846 10647
rect 9912 10671 9950 10679
rect 9912 10651 9921 10671
rect 9941 10651 9950 10671
rect 10005 10661 10070 10813
rect 10223 10787 10278 10916
rect 11262 10859 11321 10989
rect 12175 10940 12247 10941
rect 12174 10932 12273 10940
rect 12174 10929 12226 10932
rect 12174 10894 12182 10929
rect 12207 10894 12226 10929
rect 12251 10921 12273 10932
rect 12251 10920 13118 10921
rect 12251 10894 13119 10920
rect 12174 10884 13119 10894
rect 12174 10882 12273 10884
rect 11262 10841 11284 10859
rect 11302 10841 11321 10859
rect 11262 10819 11321 10841
rect 11529 10855 12061 10860
rect 11529 10835 12415 10855
rect 12435 10835 12438 10855
rect 13074 10851 13119 10884
rect 11529 10831 12438 10835
rect 9912 10642 9950 10651
rect 10003 10654 10070 10661
rect 9912 10641 9949 10642
rect 9335 10620 9371 10641
rect 9761 10620 9792 10641
rect 10003 10633 10020 10654
rect 10056 10633 10070 10654
rect 10222 10674 10278 10787
rect 11529 10784 11572 10831
rect 12022 10830 12438 10831
rect 13070 10831 13463 10851
rect 13483 10831 13486 10851
rect 12022 10829 12363 10830
rect 11679 10798 11789 10812
rect 11679 10795 11722 10798
rect 11679 10790 11683 10795
rect 11517 10783 11572 10784
rect 10222 10656 10241 10674
rect 10259 10656 10278 10674
rect 10222 10636 10278 10656
rect 11261 10760 11572 10783
rect 11261 10742 11286 10760
rect 11304 10748 11572 10760
rect 11601 10768 11683 10790
rect 11712 10768 11722 10795
rect 11750 10771 11757 10798
rect 11786 10790 11789 10798
rect 11786 10771 11851 10790
rect 11750 10768 11851 10771
rect 11601 10766 11851 10768
rect 11304 10742 11326 10748
rect 10003 10620 10070 10633
rect 9168 10616 9268 10620
rect 9168 10612 9230 10616
rect 9168 10586 9175 10612
rect 9201 10590 9230 10612
rect 9256 10590 9268 10616
rect 9201 10586 9268 10590
rect 9168 10583 9268 10586
rect 9336 10583 9371 10620
rect 9433 10617 9792 10620
rect 9433 10612 9655 10617
rect 9433 10588 9446 10612
rect 9470 10593 9655 10612
rect 9679 10593 9792 10617
rect 9470 10588 9792 10593
rect 9433 10584 9792 10588
rect 9859 10614 10070 10620
rect 9859 10612 10020 10614
rect 9859 10592 9870 10612
rect 9890 10592 10020 10612
rect 9859 10585 10020 10592
rect 9859 10584 9900 10585
rect 9335 10558 9371 10583
rect 9183 10531 9220 10532
rect 9279 10531 9316 10532
rect 9335 10531 9342 10558
rect 9083 10522 9221 10531
rect 9083 10502 9192 10522
rect 9212 10502 9221 10522
rect 9083 10495 9221 10502
rect 9279 10528 9342 10531
rect 9363 10531 9371 10558
rect 9390 10531 9427 10532
rect 9363 10528 9427 10531
rect 9279 10522 9427 10528
rect 9279 10502 9288 10522
rect 9308 10502 9398 10522
rect 9418 10502 9427 10522
rect 9083 10493 9179 10495
rect 9279 10492 9427 10502
rect 9486 10522 9523 10532
rect 9598 10531 9635 10532
rect 9579 10529 9635 10531
rect 9486 10502 9494 10522
rect 9514 10502 9523 10522
rect 9335 10491 9371 10492
rect 9183 10360 9220 10361
rect 9486 10360 9523 10502
rect 9548 10522 9635 10529
rect 9548 10519 9606 10522
rect 9548 10499 9553 10519
rect 9574 10502 9606 10519
rect 9626 10502 9635 10522
rect 9574 10499 9635 10502
rect 9548 10492 9635 10499
rect 9694 10522 9731 10532
rect 9694 10502 9702 10522
rect 9722 10502 9731 10522
rect 9548 10491 9579 10492
rect 9694 10423 9731 10502
rect 9761 10531 9792 10584
rect 10005 10577 10020 10585
rect 10060 10577 10070 10614
rect 11261 10603 11326 10742
rect 11601 10687 11638 10766
rect 11679 10753 11789 10766
rect 11753 10697 11784 10698
rect 11601 10667 11610 10687
rect 11630 10667 11638 10687
rect 10005 10568 10070 10577
rect 10218 10575 10283 10596
rect 10218 10557 10243 10575
rect 10261 10557 10283 10575
rect 11261 10585 11284 10603
rect 11302 10585 11326 10603
rect 11261 10568 11326 10585
rect 11481 10649 11549 10662
rect 11601 10657 11638 10667
rect 11697 10687 11784 10697
rect 11697 10667 11706 10687
rect 11726 10667 11784 10687
rect 11697 10658 11784 10667
rect 11697 10657 11734 10658
rect 11481 10607 11488 10649
rect 11537 10607 11549 10649
rect 11481 10604 11549 10607
rect 11753 10605 11784 10658
rect 11814 10687 11851 10766
rect 11966 10697 11997 10698
rect 11814 10667 11823 10687
rect 11843 10667 11851 10687
rect 11814 10657 11851 10667
rect 11910 10690 11997 10697
rect 11910 10687 11971 10690
rect 11910 10667 11919 10687
rect 11939 10670 11971 10687
rect 11992 10670 11997 10690
rect 11939 10667 11997 10670
rect 11910 10660 11997 10667
rect 12022 10687 12059 10829
rect 12325 10828 12362 10829
rect 13070 10826 13486 10831
rect 13070 10825 13411 10826
rect 12727 10794 12837 10808
rect 12727 10791 12770 10794
rect 12727 10786 12731 10791
rect 12649 10764 12731 10786
rect 12760 10764 12770 10791
rect 12798 10767 12805 10794
rect 12834 10786 12837 10794
rect 12834 10767 12899 10786
rect 12798 10764 12899 10767
rect 12649 10762 12899 10764
rect 12174 10697 12210 10698
rect 12022 10667 12031 10687
rect 12051 10667 12059 10687
rect 11910 10658 11966 10660
rect 11910 10657 11947 10658
rect 12022 10657 12059 10667
rect 12118 10687 12266 10697
rect 12366 10694 12462 10696
rect 12118 10667 12127 10687
rect 12147 10667 12237 10687
rect 12257 10667 12266 10687
rect 12118 10661 12266 10667
rect 12118 10658 12182 10661
rect 12118 10657 12155 10658
rect 12174 10631 12182 10658
rect 12203 10658 12266 10661
rect 12324 10687 12462 10694
rect 12324 10667 12333 10687
rect 12353 10667 12462 10687
rect 12324 10658 12462 10667
rect 12649 10683 12686 10762
rect 12727 10749 12837 10762
rect 12801 10693 12832 10694
rect 12649 10663 12658 10683
rect 12678 10663 12686 10683
rect 12203 10631 12210 10658
rect 12229 10657 12266 10658
rect 12325 10657 12362 10658
rect 12174 10606 12210 10631
rect 11645 10604 11686 10605
rect 11481 10597 11686 10604
rect 11481 10586 11655 10597
rect 9811 10531 9848 10532
rect 9761 10522 9848 10531
rect 9761 10502 9819 10522
rect 9839 10502 9848 10522
rect 9761 10492 9848 10502
rect 9907 10522 9944 10532
rect 9907 10502 9915 10522
rect 9935 10502 9944 10522
rect 9761 10491 9792 10492
rect 9756 10423 9866 10436
rect 9907 10423 9944 10502
rect 10218 10481 10283 10557
rect 11481 10553 11489 10586
rect 11482 10544 11489 10553
rect 11538 10577 11655 10586
rect 11675 10577 11686 10597
rect 11538 10569 11686 10577
rect 11753 10601 12112 10605
rect 11753 10596 12075 10601
rect 11753 10572 11866 10596
rect 11890 10577 12075 10596
rect 12099 10577 12112 10601
rect 11890 10572 12112 10577
rect 11753 10569 12112 10572
rect 12174 10569 12209 10606
rect 12277 10603 12377 10606
rect 12277 10599 12344 10603
rect 12277 10573 12289 10599
rect 12315 10577 12344 10599
rect 12370 10577 12377 10603
rect 12315 10573 12377 10577
rect 12277 10569 12377 10573
rect 11538 10553 11549 10569
rect 11538 10544 11546 10553
rect 11753 10548 11784 10569
rect 12174 10548 12210 10569
rect 11596 10547 11633 10548
rect 11261 10504 11326 10523
rect 11261 10486 11286 10504
rect 11304 10486 11326 10504
rect 9694 10421 9944 10423
rect 9694 10418 9795 10421
rect 9694 10399 9759 10418
rect 9756 10391 9759 10399
rect 9788 10391 9795 10418
rect 9823 10394 9833 10421
rect 9862 10399 9944 10421
rect 9967 10446 10284 10481
rect 9862 10394 9866 10399
rect 9823 10391 9866 10394
rect 9756 10377 9866 10391
rect 9182 10359 9523 10360
rect 9107 10357 9523 10359
rect 9967 10357 10007 10446
rect 10218 10419 10283 10446
rect 10218 10401 10241 10419
rect 10259 10401 10283 10419
rect 10218 10381 10283 10401
rect 9104 10354 10007 10357
rect 9104 10334 9110 10354
rect 9130 10334 10007 10354
rect 9104 10330 10007 10334
rect 9967 10327 10007 10330
rect 10219 10320 10284 10341
rect 8437 10312 9098 10313
rect 8437 10305 9371 10312
rect 8437 10304 9343 10305
rect 8437 10284 9288 10304
rect 9320 10285 9343 10304
rect 9368 10285 9371 10305
rect 9320 10284 9371 10285
rect 8437 10277 9371 10284
rect 8036 10235 8204 10236
rect 8439 10235 8478 10277
rect 9267 10275 9371 10277
rect 9336 10273 9371 10275
rect 10219 10302 10243 10320
rect 10261 10302 10284 10320
rect 10219 10255 10284 10302
rect 8036 10209 8480 10235
rect 8036 10207 8204 10209
rect 6797 9620 6801 9643
rect 6825 9620 6833 9643
rect 6997 9621 7096 9625
rect 6797 9599 6833 9620
rect 6797 9576 6801 9599
rect 6825 9576 6833 9599
rect 6797 9572 6833 9576
rect 6993 9615 7096 9621
rect 6993 9577 7019 9615
rect 7044 9580 7063 9615
rect 7088 9580 7096 9615
rect 7044 9577 7096 9580
rect 6993 9569 7096 9577
rect 6993 9568 7095 9569
rect 6589 9490 6757 9491
rect 6993 9490 7040 9568
rect 6589 9464 7040 9490
rect 6589 9462 6757 9464
rect 6589 9089 6616 9462
rect 6786 9414 6872 9423
rect 6786 9396 6805 9414
rect 6857 9396 6872 9414
rect 6786 9392 6872 9396
rect 6656 9229 6720 9241
rect 6656 9228 6691 9229
rect 6633 9223 6691 9228
rect 6633 9203 6636 9223
rect 6656 9209 6691 9223
rect 6711 9209 6720 9229
rect 6656 9201 6720 9209
rect 6682 9200 6720 9201
rect 6683 9199 6720 9200
rect 6786 9233 6822 9234
rect 6842 9233 6872 9392
rect 6993 9352 7040 9464
rect 6996 9237 7033 9352
rect 7261 9326 7372 9341
rect 7261 9324 7303 9326
rect 7261 9304 7268 9324
rect 7287 9304 7303 9324
rect 7261 9296 7303 9304
rect 7331 9324 7372 9326
rect 7331 9304 7345 9324
rect 7364 9304 7372 9324
rect 7331 9296 7372 9304
rect 7261 9290 7372 9296
rect 7204 9268 7453 9290
rect 7204 9237 7241 9268
rect 7417 9266 7453 9268
rect 7417 9237 7454 9266
rect 7658 9253 7737 9838
rect 7834 9386 7913 9986
rect 8036 9856 8063 10207
rect 8439 10203 8480 10209
rect 8103 9996 8167 10008
rect 8443 10004 8480 10203
rect 8942 10230 9014 10247
rect 8942 10191 8950 10230
rect 8995 10191 9014 10230
rect 8708 10093 8819 10108
rect 8708 10091 8750 10093
rect 8708 10071 8715 10091
rect 8734 10071 8750 10091
rect 8708 10063 8750 10071
rect 8778 10091 8819 10093
rect 8778 10071 8792 10091
rect 8811 10071 8819 10091
rect 8778 10063 8819 10071
rect 8708 10057 8819 10063
rect 8651 10035 8900 10057
rect 8651 10004 8688 10035
rect 8864 10033 8900 10035
rect 8864 10004 8901 10033
rect 8103 9995 8138 9996
rect 8080 9990 8138 9995
rect 8080 9970 8083 9990
rect 8103 9976 8138 9990
rect 8158 9976 8167 9996
rect 8103 9968 8167 9976
rect 8129 9967 8167 9968
rect 8130 9966 8167 9967
rect 8233 10000 8269 10001
rect 8341 10000 8377 10001
rect 8233 9992 8377 10000
rect 8233 9972 8241 9992
rect 8261 9972 8349 9992
rect 8369 9972 8377 9992
rect 8233 9966 8377 9972
rect 8443 9996 8481 10004
rect 8549 10000 8585 10001
rect 8443 9976 8452 9996
rect 8472 9976 8481 9996
rect 8443 9967 8481 9976
rect 8500 9993 8585 10000
rect 8500 9973 8507 9993
rect 8528 9992 8585 9993
rect 8528 9973 8557 9992
rect 8500 9972 8557 9973
rect 8577 9972 8585 9992
rect 8443 9966 8480 9967
rect 8500 9966 8585 9972
rect 8651 9996 8689 10004
rect 8762 10000 8798 10001
rect 8651 9976 8660 9996
rect 8680 9976 8689 9996
rect 8651 9967 8689 9976
rect 8713 9992 8798 10000
rect 8713 9972 8770 9992
rect 8790 9972 8798 9992
rect 8651 9966 8688 9967
rect 8713 9966 8798 9972
rect 8864 9996 8902 10004
rect 8864 9976 8873 9996
rect 8893 9976 8902 9996
rect 8864 9967 8902 9976
rect 8942 9981 9014 10191
rect 9084 10225 10284 10255
rect 9084 10224 9528 10225
rect 9084 10222 9252 10224
rect 8942 9967 9025 9981
rect 8864 9966 8901 9967
rect 8287 9945 8323 9966
rect 8713 9945 8744 9966
rect 8942 9945 8959 9967
rect 8120 9941 8220 9945
rect 8120 9937 8182 9941
rect 8120 9911 8127 9937
rect 8153 9915 8182 9937
rect 8208 9915 8220 9941
rect 8153 9911 8220 9915
rect 8120 9908 8220 9911
rect 8288 9908 8323 9945
rect 8385 9942 8744 9945
rect 8385 9937 8607 9942
rect 8385 9913 8398 9937
rect 8422 9918 8607 9937
rect 8631 9918 8744 9942
rect 8422 9913 8744 9918
rect 8385 9909 8744 9913
rect 8811 9937 8959 9945
rect 8811 9917 8822 9937
rect 8842 9934 8959 9937
rect 9012 9934 9025 9967
rect 8842 9917 9025 9934
rect 8811 9910 9025 9917
rect 8811 9909 8852 9910
rect 8942 9909 9025 9910
rect 8287 9883 8323 9908
rect 8135 9856 8172 9857
rect 8231 9856 8268 9857
rect 8287 9856 8294 9883
rect 8035 9847 8173 9856
rect 8035 9827 8144 9847
rect 8164 9827 8173 9847
rect 8035 9820 8173 9827
rect 8231 9853 8294 9856
rect 8315 9856 8323 9883
rect 8342 9856 8379 9857
rect 8315 9853 8379 9856
rect 8231 9847 8379 9853
rect 8231 9827 8240 9847
rect 8260 9827 8350 9847
rect 8370 9827 8379 9847
rect 8035 9818 8131 9820
rect 8231 9817 8379 9827
rect 8438 9847 8475 9857
rect 8550 9856 8587 9857
rect 8531 9854 8587 9856
rect 8438 9827 8446 9847
rect 8466 9827 8475 9847
rect 8287 9816 8323 9817
rect 8135 9685 8172 9686
rect 8438 9685 8475 9827
rect 8500 9847 8587 9854
rect 8500 9844 8558 9847
rect 8500 9824 8505 9844
rect 8526 9827 8558 9844
rect 8578 9827 8587 9847
rect 8526 9824 8587 9827
rect 8500 9817 8587 9824
rect 8646 9847 8683 9857
rect 8646 9827 8654 9847
rect 8674 9827 8683 9847
rect 8500 9816 8531 9817
rect 8646 9748 8683 9827
rect 8713 9856 8744 9909
rect 8950 9876 8964 9909
rect 9017 9876 9025 9909
rect 8950 9870 9025 9876
rect 8950 9865 9020 9870
rect 8763 9856 8800 9857
rect 8713 9847 8800 9856
rect 8713 9827 8771 9847
rect 8791 9827 8800 9847
rect 8713 9817 8800 9827
rect 8859 9847 8896 9857
rect 9084 9852 9111 10222
rect 9151 9992 9215 10004
rect 9491 10000 9528 10224
rect 9999 10205 10063 10207
rect 9995 10193 10063 10205
rect 9995 10160 10006 10193
rect 10046 10160 10063 10193
rect 9995 10150 10063 10160
rect 9756 10089 9867 10104
rect 9756 10087 9798 10089
rect 9756 10067 9763 10087
rect 9782 10067 9798 10087
rect 9756 10059 9798 10067
rect 9826 10087 9867 10089
rect 9826 10067 9840 10087
rect 9859 10067 9867 10087
rect 9826 10059 9867 10067
rect 9756 10053 9867 10059
rect 9699 10031 9948 10053
rect 9699 10000 9736 10031
rect 9912 10029 9948 10031
rect 9912 10000 9949 10029
rect 9151 9991 9186 9992
rect 9128 9986 9186 9991
rect 9128 9966 9131 9986
rect 9151 9972 9186 9986
rect 9206 9972 9215 9992
rect 9151 9964 9215 9972
rect 9177 9963 9215 9964
rect 9178 9962 9215 9963
rect 9281 9996 9317 9997
rect 9389 9996 9425 9997
rect 9281 9988 9425 9996
rect 9281 9968 9289 9988
rect 9309 9968 9397 9988
rect 9417 9968 9425 9988
rect 9281 9962 9425 9968
rect 9491 9992 9529 10000
rect 9597 9996 9633 9997
rect 9491 9972 9500 9992
rect 9520 9972 9529 9992
rect 9491 9963 9529 9972
rect 9548 9989 9633 9996
rect 9548 9969 9555 9989
rect 9576 9988 9633 9989
rect 9576 9969 9605 9988
rect 9548 9968 9605 9969
rect 9625 9968 9633 9988
rect 9491 9962 9528 9963
rect 9548 9962 9633 9968
rect 9699 9992 9737 10000
rect 9810 9996 9846 9997
rect 9699 9972 9708 9992
rect 9728 9972 9737 9992
rect 9699 9963 9737 9972
rect 9761 9988 9846 9996
rect 9761 9968 9818 9988
rect 9838 9968 9846 9988
rect 9699 9962 9736 9963
rect 9761 9962 9846 9968
rect 9912 9992 9950 10000
rect 9912 9972 9921 9992
rect 9941 9972 9950 9992
rect 9912 9963 9950 9972
rect 9999 9966 10063 10150
rect 10219 10024 10284 10225
rect 11261 10285 11326 10486
rect 11482 10360 11546 10544
rect 11595 10538 11633 10547
rect 11595 10518 11604 10538
rect 11624 10518 11633 10538
rect 11595 10510 11633 10518
rect 11699 10542 11784 10548
rect 11809 10547 11846 10548
rect 11699 10522 11707 10542
rect 11727 10522 11784 10542
rect 11699 10514 11784 10522
rect 11808 10538 11846 10547
rect 11808 10518 11817 10538
rect 11837 10518 11846 10538
rect 11699 10513 11735 10514
rect 11808 10510 11846 10518
rect 11912 10542 11997 10548
rect 12017 10547 12054 10548
rect 11912 10522 11920 10542
rect 11940 10541 11997 10542
rect 11940 10522 11969 10541
rect 11912 10521 11969 10522
rect 11990 10521 11997 10541
rect 11912 10514 11997 10521
rect 12016 10538 12054 10547
rect 12016 10518 12025 10538
rect 12045 10518 12054 10538
rect 11912 10513 11948 10514
rect 12016 10510 12054 10518
rect 12120 10542 12264 10548
rect 12120 10522 12128 10542
rect 12148 10522 12236 10542
rect 12256 10522 12264 10542
rect 12120 10514 12264 10522
rect 12120 10513 12156 10514
rect 12228 10513 12264 10514
rect 12330 10547 12367 10548
rect 12330 10546 12368 10547
rect 12330 10538 12394 10546
rect 12330 10518 12339 10538
rect 12359 10524 12394 10538
rect 12414 10524 12417 10544
rect 12359 10519 12417 10524
rect 12359 10518 12394 10519
rect 11596 10481 11633 10510
rect 11597 10479 11633 10481
rect 11809 10479 11846 10510
rect 11597 10457 11846 10479
rect 11678 10451 11789 10457
rect 11678 10443 11719 10451
rect 11678 10423 11686 10443
rect 11705 10423 11719 10443
rect 11678 10421 11719 10423
rect 11747 10443 11789 10451
rect 11747 10423 11763 10443
rect 11782 10423 11789 10443
rect 11747 10421 11789 10423
rect 11678 10406 11789 10421
rect 11482 10350 11550 10360
rect 11482 10317 11499 10350
rect 11539 10317 11550 10350
rect 11482 10305 11550 10317
rect 11482 10303 11546 10305
rect 12017 10286 12054 10510
rect 12330 10506 12394 10518
rect 12434 10288 12461 10658
rect 12649 10653 12686 10663
rect 12745 10683 12832 10693
rect 12745 10663 12754 10683
rect 12774 10663 12832 10683
rect 12745 10654 12832 10663
rect 12745 10653 12782 10654
rect 12525 10640 12595 10645
rect 12520 10634 12595 10640
rect 12520 10601 12528 10634
rect 12581 10601 12595 10634
rect 12801 10601 12832 10654
rect 12862 10683 12899 10762
rect 13014 10693 13045 10694
rect 12862 10663 12871 10683
rect 12891 10663 12899 10683
rect 12862 10653 12899 10663
rect 12958 10686 13045 10693
rect 12958 10683 13019 10686
rect 12958 10663 12967 10683
rect 12987 10666 13019 10683
rect 13040 10666 13045 10686
rect 12987 10663 13045 10666
rect 12958 10656 13045 10663
rect 13070 10683 13107 10825
rect 13373 10824 13410 10825
rect 13222 10693 13258 10694
rect 13070 10663 13079 10683
rect 13099 10663 13107 10683
rect 12958 10654 13014 10656
rect 12958 10653 12995 10654
rect 13070 10653 13107 10663
rect 13166 10683 13314 10693
rect 13414 10690 13510 10692
rect 13166 10663 13175 10683
rect 13195 10663 13285 10683
rect 13305 10663 13314 10683
rect 13166 10657 13314 10663
rect 13166 10654 13230 10657
rect 13166 10653 13203 10654
rect 13222 10627 13230 10654
rect 13251 10654 13314 10657
rect 13372 10683 13510 10690
rect 13372 10663 13381 10683
rect 13401 10663 13510 10683
rect 13372 10654 13510 10663
rect 13251 10627 13258 10654
rect 13277 10653 13314 10654
rect 13373 10653 13410 10654
rect 13222 10602 13258 10627
rect 12520 10600 12603 10601
rect 12693 10600 12734 10601
rect 12520 10593 12734 10600
rect 12520 10576 12703 10593
rect 12520 10543 12533 10576
rect 12586 10573 12703 10576
rect 12723 10573 12734 10593
rect 12586 10565 12734 10573
rect 12801 10597 13160 10601
rect 12801 10592 13123 10597
rect 12801 10568 12914 10592
rect 12938 10573 13123 10592
rect 13147 10573 13160 10597
rect 12938 10568 13160 10573
rect 12801 10565 13160 10568
rect 13222 10565 13257 10602
rect 13325 10599 13425 10602
rect 13325 10595 13392 10599
rect 13325 10569 13337 10595
rect 13363 10573 13392 10595
rect 13418 10573 13425 10599
rect 13363 10569 13425 10573
rect 13325 10565 13425 10569
rect 12586 10543 12603 10565
rect 12801 10544 12832 10565
rect 13222 10544 13258 10565
rect 12644 10543 12681 10544
rect 12520 10529 12603 10543
rect 12293 10286 12461 10288
rect 12017 10285 12461 10286
rect 11261 10255 12461 10285
rect 12531 10319 12603 10529
rect 12643 10534 12681 10543
rect 12643 10514 12652 10534
rect 12672 10514 12681 10534
rect 12643 10506 12681 10514
rect 12747 10538 12832 10544
rect 12857 10543 12894 10544
rect 12747 10518 12755 10538
rect 12775 10518 12832 10538
rect 12747 10510 12832 10518
rect 12856 10534 12894 10543
rect 12856 10514 12865 10534
rect 12885 10514 12894 10534
rect 12747 10509 12783 10510
rect 12856 10506 12894 10514
rect 12960 10538 13045 10544
rect 13065 10543 13102 10544
rect 12960 10518 12968 10538
rect 12988 10537 13045 10538
rect 12988 10518 13017 10537
rect 12960 10517 13017 10518
rect 13038 10517 13045 10537
rect 12960 10510 13045 10517
rect 13064 10534 13102 10543
rect 13064 10514 13073 10534
rect 13093 10514 13102 10534
rect 12960 10509 12996 10510
rect 13064 10506 13102 10514
rect 13168 10538 13312 10544
rect 13168 10518 13176 10538
rect 13196 10518 13284 10538
rect 13304 10518 13312 10538
rect 13168 10510 13312 10518
rect 13168 10509 13204 10510
rect 13276 10509 13312 10510
rect 13378 10543 13415 10544
rect 13378 10542 13416 10543
rect 13378 10534 13442 10542
rect 13378 10514 13387 10534
rect 13407 10520 13442 10534
rect 13462 10520 13465 10540
rect 13407 10515 13465 10520
rect 13407 10514 13442 10515
rect 12644 10477 12681 10506
rect 12645 10475 12681 10477
rect 12857 10475 12894 10506
rect 12645 10453 12894 10475
rect 12726 10447 12837 10453
rect 12726 10439 12767 10447
rect 12726 10419 12734 10439
rect 12753 10419 12767 10439
rect 12726 10417 12767 10419
rect 12795 10439 12837 10447
rect 12795 10419 12811 10439
rect 12830 10419 12837 10439
rect 12795 10417 12837 10419
rect 12726 10402 12837 10417
rect 12531 10280 12550 10319
rect 12595 10280 12603 10319
rect 12531 10263 12603 10280
rect 13065 10307 13102 10506
rect 13378 10502 13442 10514
rect 13065 10301 13106 10307
rect 13482 10303 13509 10654
rect 13638 10606 13709 11085
rect 13638 10522 13707 10606
rect 13341 10301 13509 10303
rect 13065 10275 13509 10301
rect 11261 10208 11326 10255
rect 11261 10190 11284 10208
rect 11302 10190 11326 10208
rect 12174 10235 12209 10237
rect 12174 10233 12278 10235
rect 13067 10233 13106 10275
rect 13341 10274 13509 10275
rect 12174 10226 13108 10233
rect 12174 10225 12225 10226
rect 12174 10205 12177 10225
rect 12202 10206 12225 10225
rect 12257 10206 13108 10226
rect 12202 10205 13108 10206
rect 12174 10198 13108 10205
rect 12447 10197 13108 10198
rect 11261 10169 11326 10190
rect 11538 10180 11578 10183
rect 11538 10176 12441 10180
rect 11538 10156 12415 10176
rect 12435 10156 12441 10176
rect 11538 10153 12441 10156
rect 11262 10109 11327 10129
rect 11262 10091 11286 10109
rect 11304 10091 11327 10109
rect 11262 10064 11327 10091
rect 11538 10064 11578 10153
rect 12022 10151 12438 10153
rect 12022 10150 12363 10151
rect 11679 10119 11789 10133
rect 11679 10116 11722 10119
rect 11679 10111 11683 10116
rect 11261 10029 11578 10064
rect 11601 10089 11683 10111
rect 11712 10089 11722 10116
rect 11750 10092 11757 10119
rect 11786 10111 11789 10119
rect 11786 10092 11851 10111
rect 11750 10089 11851 10092
rect 11601 10087 11851 10089
rect 10219 10006 10241 10024
rect 10259 10006 10284 10024
rect 10219 9987 10284 10006
rect 9912 9962 9949 9963
rect 9335 9941 9371 9962
rect 9761 9941 9792 9962
rect 9999 9957 10007 9966
rect 9996 9941 10007 9957
rect 9168 9937 9268 9941
rect 9168 9933 9230 9937
rect 9168 9907 9175 9933
rect 9201 9911 9230 9933
rect 9256 9911 9268 9937
rect 9201 9907 9268 9911
rect 9168 9904 9268 9907
rect 9336 9904 9371 9941
rect 9433 9938 9792 9941
rect 9433 9933 9655 9938
rect 9433 9909 9446 9933
rect 9470 9914 9655 9933
rect 9679 9914 9792 9938
rect 9470 9909 9792 9914
rect 9433 9905 9792 9909
rect 9859 9933 10007 9941
rect 9859 9913 9870 9933
rect 9890 9924 10007 9933
rect 10056 9957 10063 9966
rect 10056 9924 10064 9957
rect 11262 9953 11327 10029
rect 11601 10008 11638 10087
rect 11679 10074 11789 10087
rect 11753 10018 11784 10019
rect 11601 9988 11610 10008
rect 11630 9988 11638 10008
rect 11601 9978 11638 9988
rect 11697 10008 11784 10018
rect 11697 9988 11706 10008
rect 11726 9988 11784 10008
rect 11697 9979 11784 9988
rect 11697 9978 11734 9979
rect 9890 9913 10064 9924
rect 9859 9906 10064 9913
rect 9859 9905 9900 9906
rect 9335 9879 9371 9904
rect 9183 9852 9220 9853
rect 9279 9852 9316 9853
rect 9335 9852 9342 9879
rect 8859 9827 8867 9847
rect 8887 9827 8896 9847
rect 8713 9816 8744 9817
rect 8708 9748 8818 9761
rect 8859 9748 8896 9827
rect 9083 9843 9221 9852
rect 9083 9823 9192 9843
rect 9212 9823 9221 9843
rect 9083 9816 9221 9823
rect 9279 9849 9342 9852
rect 9363 9852 9371 9879
rect 9390 9852 9427 9853
rect 9363 9849 9427 9852
rect 9279 9843 9427 9849
rect 9279 9823 9288 9843
rect 9308 9823 9398 9843
rect 9418 9823 9427 9843
rect 9083 9814 9179 9816
rect 9279 9813 9427 9823
rect 9486 9843 9523 9853
rect 9598 9852 9635 9853
rect 9579 9850 9635 9852
rect 9486 9823 9494 9843
rect 9514 9823 9523 9843
rect 9335 9812 9371 9813
rect 8646 9746 8896 9748
rect 8646 9743 8747 9746
rect 8646 9724 8711 9743
rect 8708 9716 8711 9724
rect 8740 9716 8747 9743
rect 8775 9719 8785 9746
rect 8814 9724 8896 9746
rect 8814 9719 8818 9724
rect 8775 9716 8818 9719
rect 8708 9702 8818 9716
rect 8134 9684 8475 9685
rect 8059 9679 8475 9684
rect 9183 9681 9220 9682
rect 9486 9681 9523 9823
rect 9548 9843 9635 9850
rect 9548 9840 9606 9843
rect 9548 9820 9553 9840
rect 9574 9823 9606 9840
rect 9626 9823 9635 9843
rect 9574 9820 9635 9823
rect 9548 9813 9635 9820
rect 9694 9843 9731 9853
rect 9694 9823 9702 9843
rect 9722 9823 9731 9843
rect 9548 9812 9579 9813
rect 9694 9744 9731 9823
rect 9761 9852 9792 9905
rect 9996 9903 10064 9906
rect 9996 9861 10008 9903
rect 10057 9861 10064 9903
rect 9811 9852 9848 9853
rect 9761 9843 9848 9852
rect 9761 9823 9819 9843
rect 9839 9823 9848 9843
rect 9761 9813 9848 9823
rect 9907 9843 9944 9853
rect 9996 9848 10064 9861
rect 10219 9925 10284 9942
rect 10219 9907 10243 9925
rect 10261 9907 10284 9925
rect 11262 9935 11284 9953
rect 11302 9935 11327 9953
rect 11262 9914 11327 9935
rect 11475 9933 11540 9942
rect 9907 9823 9915 9843
rect 9935 9823 9944 9843
rect 9761 9812 9792 9813
rect 9756 9744 9866 9757
rect 9907 9744 9944 9823
rect 10219 9768 10284 9907
rect 11475 9896 11485 9933
rect 11525 9925 11540 9933
rect 11753 9926 11784 9979
rect 11814 10008 11851 10087
rect 11966 10018 11997 10019
rect 11814 9988 11823 10008
rect 11843 9988 11851 10008
rect 11814 9978 11851 9988
rect 11910 10011 11997 10018
rect 11910 10008 11971 10011
rect 11910 9988 11919 10008
rect 11939 9991 11971 10008
rect 11992 9991 11997 10011
rect 11939 9988 11997 9991
rect 11910 9981 11997 9988
rect 12022 10008 12059 10150
rect 12325 10149 12362 10150
rect 12174 10018 12210 10019
rect 12022 9988 12031 10008
rect 12051 9988 12059 10008
rect 11910 9979 11966 9981
rect 11910 9978 11947 9979
rect 12022 9978 12059 9988
rect 12118 10008 12266 10018
rect 12366 10015 12462 10017
rect 12118 9988 12127 10008
rect 12147 9988 12237 10008
rect 12257 9988 12266 10008
rect 12118 9982 12266 9988
rect 12118 9979 12182 9982
rect 12118 9978 12155 9979
rect 12174 9952 12182 9979
rect 12203 9979 12266 9982
rect 12324 10008 12462 10015
rect 12324 9988 12333 10008
rect 12353 9988 12462 10008
rect 13642 10006 13704 10522
rect 12324 9979 12462 9988
rect 12203 9952 12210 9979
rect 12229 9978 12266 9979
rect 12325 9978 12362 9979
rect 12174 9927 12210 9952
rect 11645 9925 11686 9926
rect 11525 9918 11686 9925
rect 11525 9898 11655 9918
rect 11675 9898 11686 9918
rect 11525 9896 11686 9898
rect 11475 9890 11686 9896
rect 11753 9922 12112 9926
rect 11753 9917 12075 9922
rect 11753 9893 11866 9917
rect 11890 9898 12075 9917
rect 12099 9898 12112 9922
rect 11890 9893 12112 9898
rect 11753 9890 12112 9893
rect 12174 9890 12209 9927
rect 12277 9924 12377 9927
rect 12277 9920 12344 9924
rect 12277 9894 12289 9920
rect 12315 9898 12344 9920
rect 12370 9898 12377 9924
rect 12315 9894 12377 9898
rect 12277 9890 12377 9894
rect 11475 9877 11542 9890
rect 10219 9762 10241 9768
rect 9694 9742 9944 9744
rect 9694 9739 9795 9742
rect 9694 9720 9759 9739
rect 9756 9712 9759 9720
rect 9788 9712 9795 9739
rect 9823 9715 9833 9742
rect 9862 9720 9944 9742
rect 9973 9750 10241 9762
rect 10259 9750 10284 9768
rect 9973 9727 10284 9750
rect 11267 9854 11323 9874
rect 11267 9836 11286 9854
rect 11304 9836 11323 9854
rect 9973 9726 10028 9727
rect 9862 9715 9866 9720
rect 9823 9712 9866 9715
rect 9756 9698 9866 9712
rect 9182 9680 9523 9681
rect 8059 9659 8062 9679
rect 8082 9659 8475 9679
rect 9107 9679 9523 9680
rect 9973 9679 10016 9726
rect 11267 9723 11323 9836
rect 11475 9856 11489 9877
rect 11525 9856 11542 9877
rect 11753 9869 11784 9890
rect 12174 9869 12210 9890
rect 11596 9868 11633 9869
rect 11475 9849 11542 9856
rect 11595 9859 11633 9868
rect 9107 9675 10016 9679
rect 8426 9626 8471 9659
rect 9107 9655 9110 9675
rect 9130 9655 10016 9675
rect 9484 9650 10016 9655
rect 10224 9669 10283 9691
rect 10224 9651 10243 9669
rect 10261 9651 10283 9669
rect 9272 9626 9371 9628
rect 8426 9616 9371 9626
rect 8426 9590 9294 9616
rect 8427 9589 9294 9590
rect 9272 9578 9294 9589
rect 9319 9581 9338 9616
rect 9363 9581 9371 9616
rect 9319 9578 9371 9581
rect 10224 9580 10283 9651
rect 11267 9585 11322 9723
rect 11475 9697 11540 9849
rect 11595 9839 11604 9859
rect 11624 9839 11633 9859
rect 11595 9831 11633 9839
rect 11699 9863 11784 9869
rect 11809 9868 11846 9869
rect 11699 9843 11707 9863
rect 11727 9843 11784 9863
rect 11699 9835 11784 9843
rect 11808 9859 11846 9868
rect 11808 9839 11817 9859
rect 11837 9839 11846 9859
rect 11699 9834 11735 9835
rect 11808 9831 11846 9839
rect 11912 9863 11997 9869
rect 12017 9868 12054 9869
rect 11912 9843 11920 9863
rect 11940 9862 11997 9863
rect 11940 9843 11969 9862
rect 11912 9842 11969 9843
rect 11990 9842 11997 9862
rect 11912 9835 11997 9842
rect 12016 9859 12054 9868
rect 12016 9839 12025 9859
rect 12045 9839 12054 9859
rect 11912 9834 11948 9835
rect 12016 9831 12054 9839
rect 12120 9863 12264 9869
rect 12120 9843 12128 9863
rect 12148 9843 12236 9863
rect 12256 9843 12264 9863
rect 12120 9835 12264 9843
rect 12120 9834 12156 9835
rect 12228 9834 12264 9835
rect 12330 9868 12367 9869
rect 12330 9867 12368 9868
rect 12330 9859 12394 9867
rect 12330 9839 12339 9859
rect 12359 9845 12394 9859
rect 12414 9845 12417 9865
rect 12359 9840 12417 9845
rect 12359 9839 12394 9840
rect 11596 9802 11633 9831
rect 11597 9800 11633 9802
rect 11809 9800 11846 9831
rect 11597 9778 11846 9800
rect 11678 9772 11789 9778
rect 11678 9764 11719 9772
rect 11678 9744 11686 9764
rect 11705 9744 11719 9764
rect 11678 9742 11719 9744
rect 11747 9764 11789 9772
rect 11747 9744 11763 9764
rect 11782 9744 11789 9764
rect 11747 9742 11789 9744
rect 11678 9729 11789 9742
rect 12017 9732 12054 9831
rect 12330 9827 12394 9839
rect 11468 9687 11589 9697
rect 11468 9685 11537 9687
rect 11468 9644 11481 9685
rect 11518 9646 11537 9685
rect 11574 9646 11589 9687
rect 11518 9644 11589 9646
rect 11468 9626 11589 9644
rect 11260 9582 11324 9585
rect 11680 9582 11784 9588
rect 12015 9582 12056 9732
rect 12434 9724 12461 9979
rect 12523 9969 12603 9980
rect 12523 9943 12540 9969
rect 12580 9943 12603 9969
rect 12523 9916 12603 9943
rect 12523 9890 12544 9916
rect 12584 9890 12603 9916
rect 12523 9871 12603 9890
rect 12523 9845 12547 9871
rect 12587 9845 12603 9871
rect 12523 9794 12603 9845
rect 13626 9971 13704 10006
rect 13626 9909 13708 9971
rect 13626 9886 13654 9909
rect 13680 9886 13708 9909
rect 13626 9866 13708 9886
rect 9272 9570 9371 9578
rect 9298 9569 9370 9570
rect 8952 9543 9019 9562
rect 8952 9522 8969 9543
rect 7833 9344 7913 9386
rect 8950 9477 8969 9522
rect 8999 9522 9019 9543
rect 8999 9477 9020 9522
rect 9489 9519 9530 9521
rect 9761 9519 9865 9521
rect 10221 9519 10285 9580
rect 6894 9233 6930 9234
rect 6786 9225 6930 9233
rect 6786 9205 6794 9225
rect 6814 9205 6902 9225
rect 6922 9205 6930 9225
rect 6786 9199 6930 9205
rect 6996 9229 7034 9237
rect 7102 9233 7138 9234
rect 6996 9209 7005 9229
rect 7025 9209 7034 9229
rect 6996 9200 7034 9209
rect 7053 9226 7138 9233
rect 7053 9206 7060 9226
rect 7081 9225 7138 9226
rect 7081 9206 7110 9225
rect 7053 9205 7110 9206
rect 7130 9205 7138 9225
rect 6996 9199 7033 9200
rect 7053 9199 7138 9205
rect 7204 9229 7242 9237
rect 7315 9233 7351 9234
rect 7204 9209 7213 9229
rect 7233 9209 7242 9229
rect 7204 9200 7242 9209
rect 7266 9225 7351 9233
rect 7266 9205 7323 9225
rect 7343 9205 7351 9225
rect 7204 9199 7241 9200
rect 7266 9199 7351 9205
rect 7417 9229 7455 9237
rect 7417 9209 7426 9229
rect 7446 9209 7455 9229
rect 7417 9200 7455 9209
rect 7655 9217 7741 9253
rect 7417 9199 7454 9200
rect 6840 9178 6876 9199
rect 7266 9178 7297 9199
rect 7493 9178 7539 9182
rect 6673 9174 6773 9178
rect 6673 9170 6735 9174
rect 6673 9144 6680 9170
rect 6706 9148 6735 9170
rect 6761 9148 6773 9174
rect 6706 9144 6773 9148
rect 6673 9141 6773 9144
rect 6841 9141 6876 9178
rect 6938 9175 7297 9178
rect 6938 9170 7160 9175
rect 6938 9146 6951 9170
rect 6975 9151 7160 9170
rect 7184 9151 7297 9175
rect 6975 9146 7297 9151
rect 6938 9142 7297 9146
rect 7364 9170 7539 9178
rect 7364 9150 7375 9170
rect 7395 9150 7539 9170
rect 7655 9176 7672 9217
rect 7726 9176 7741 9217
rect 7655 9157 7741 9176
rect 7364 9143 7539 9150
rect 7364 9142 7405 9143
rect 6840 9116 6876 9141
rect 6688 9089 6725 9090
rect 6784 9089 6821 9090
rect 6840 9089 6847 9116
rect 6588 9080 6726 9089
rect 6588 9060 6697 9080
rect 6717 9060 6726 9080
rect 6588 9053 6726 9060
rect 6784 9086 6847 9089
rect 6868 9089 6876 9116
rect 6895 9089 6932 9090
rect 6868 9086 6932 9089
rect 6784 9080 6932 9086
rect 6784 9060 6793 9080
rect 6813 9060 6903 9080
rect 6923 9060 6932 9080
rect 6588 9051 6684 9053
rect 6784 9050 6932 9060
rect 6991 9080 7028 9090
rect 7103 9089 7140 9090
rect 7084 9087 7140 9089
rect 6991 9060 6999 9080
rect 7019 9060 7028 9080
rect 6840 9049 6876 9050
rect 6688 8918 6725 8919
rect 6991 8918 7028 9060
rect 7053 9080 7140 9087
rect 7053 9077 7111 9080
rect 7053 9057 7058 9077
rect 7079 9060 7111 9077
rect 7131 9060 7140 9080
rect 7079 9057 7140 9060
rect 7053 9050 7140 9057
rect 7199 9080 7236 9090
rect 7199 9060 7207 9080
rect 7227 9060 7236 9080
rect 7053 9049 7084 9050
rect 7199 8981 7236 9060
rect 7266 9089 7297 9142
rect 7316 9089 7353 9090
rect 7266 9080 7353 9089
rect 7266 9060 7324 9080
rect 7344 9060 7353 9080
rect 7266 9050 7353 9060
rect 7412 9080 7449 9090
rect 7412 9060 7420 9080
rect 7440 9060 7449 9080
rect 7266 9049 7297 9050
rect 7261 8981 7371 8994
rect 7412 8981 7449 9060
rect 7493 9060 7539 9143
rect 7833 9060 7908 9344
rect 8950 9269 9020 9477
rect 9082 9484 10285 9519
rect 9082 9470 9110 9484
rect 9084 9339 9110 9470
rect 9489 9481 10285 9484
rect 11260 9579 12056 9582
rect 12435 9593 12461 9724
rect 12435 9579 12463 9593
rect 11260 9544 12463 9579
rect 12525 9586 12595 9794
rect 11260 9483 11324 9544
rect 11680 9542 11784 9544
rect 12015 9542 12056 9544
rect 12525 9541 12546 9586
rect 12526 9520 12546 9541
rect 12576 9541 12595 9586
rect 12576 9520 12593 9541
rect 12526 9501 12593 9520
rect 12175 9493 12247 9494
rect 12174 9485 12273 9493
rect 8942 9218 9022 9269
rect 8942 9192 8958 9218
rect 8998 9192 9022 9218
rect 8942 9173 9022 9192
rect 8942 9147 8961 9173
rect 9001 9147 9022 9173
rect 8942 9120 9022 9147
rect 8942 9094 8965 9120
rect 9005 9094 9022 9120
rect 8942 9083 9022 9094
rect 9084 9084 9111 9339
rect 9489 9331 9530 9481
rect 9761 9475 9865 9481
rect 10221 9478 10285 9481
rect 9956 9419 10077 9437
rect 9956 9417 10027 9419
rect 9956 9376 9971 9417
rect 10008 9378 10027 9417
rect 10064 9378 10077 9419
rect 10008 9376 10077 9378
rect 9956 9366 10077 9376
rect 9151 9224 9215 9236
rect 9491 9232 9528 9331
rect 9756 9321 9867 9334
rect 9756 9319 9798 9321
rect 9756 9299 9763 9319
rect 9782 9299 9798 9319
rect 9756 9291 9798 9299
rect 9826 9319 9867 9321
rect 9826 9299 9840 9319
rect 9859 9299 9867 9319
rect 9826 9291 9867 9299
rect 9756 9285 9867 9291
rect 9699 9263 9948 9285
rect 9699 9232 9736 9263
rect 9912 9261 9948 9263
rect 9912 9232 9949 9261
rect 9151 9223 9186 9224
rect 9128 9218 9186 9223
rect 9128 9198 9131 9218
rect 9151 9204 9186 9218
rect 9206 9204 9215 9224
rect 9151 9196 9215 9204
rect 9177 9195 9215 9196
rect 9178 9194 9215 9195
rect 9281 9228 9317 9229
rect 9389 9228 9425 9229
rect 9281 9220 9425 9228
rect 9281 9200 9289 9220
rect 9309 9200 9397 9220
rect 9417 9200 9425 9220
rect 9281 9194 9425 9200
rect 9491 9224 9529 9232
rect 9597 9228 9633 9229
rect 9491 9204 9500 9224
rect 9520 9204 9529 9224
rect 9491 9195 9529 9204
rect 9548 9221 9633 9228
rect 9548 9201 9555 9221
rect 9576 9220 9633 9221
rect 9576 9201 9605 9220
rect 9548 9200 9605 9201
rect 9625 9200 9633 9220
rect 9491 9194 9528 9195
rect 9548 9194 9633 9200
rect 9699 9224 9737 9232
rect 9810 9228 9846 9229
rect 9699 9204 9708 9224
rect 9728 9204 9737 9224
rect 9699 9195 9737 9204
rect 9761 9220 9846 9228
rect 9761 9200 9818 9220
rect 9838 9200 9846 9220
rect 9699 9194 9736 9195
rect 9761 9194 9846 9200
rect 9912 9224 9950 9232
rect 9912 9204 9921 9224
rect 9941 9204 9950 9224
rect 10005 9214 10070 9366
rect 10223 9340 10278 9478
rect 11262 9412 11321 9483
rect 12174 9482 12226 9485
rect 12174 9447 12182 9482
rect 12207 9447 12226 9482
rect 12251 9474 12273 9485
rect 12251 9473 13118 9474
rect 12251 9447 13119 9473
rect 12174 9437 13119 9447
rect 12174 9435 12273 9437
rect 11262 9394 11284 9412
rect 11302 9394 11321 9412
rect 11262 9372 11321 9394
rect 11529 9408 12061 9413
rect 11529 9388 12415 9408
rect 12435 9388 12438 9408
rect 13074 9404 13119 9437
rect 11529 9384 12438 9388
rect 9912 9195 9950 9204
rect 10003 9207 10070 9214
rect 9912 9194 9949 9195
rect 9335 9173 9371 9194
rect 9761 9173 9792 9194
rect 10003 9186 10020 9207
rect 10056 9186 10070 9207
rect 10222 9227 10278 9340
rect 11529 9337 11572 9384
rect 12022 9383 12438 9384
rect 13070 9384 13463 9404
rect 13483 9384 13486 9404
rect 12022 9382 12363 9383
rect 11679 9351 11789 9365
rect 11679 9348 11722 9351
rect 11679 9343 11683 9348
rect 11517 9336 11572 9337
rect 10222 9209 10241 9227
rect 10259 9209 10278 9227
rect 10222 9189 10278 9209
rect 11261 9313 11572 9336
rect 11261 9295 11286 9313
rect 11304 9301 11572 9313
rect 11601 9321 11683 9343
rect 11712 9321 11722 9348
rect 11750 9324 11757 9351
rect 11786 9343 11789 9351
rect 11786 9324 11851 9343
rect 11750 9321 11851 9324
rect 11601 9319 11851 9321
rect 11304 9295 11326 9301
rect 10003 9173 10070 9186
rect 9168 9169 9268 9173
rect 9168 9165 9230 9169
rect 9168 9139 9175 9165
rect 9201 9143 9230 9165
rect 9256 9143 9268 9169
rect 9201 9139 9268 9143
rect 9168 9136 9268 9139
rect 9336 9136 9371 9173
rect 9433 9170 9792 9173
rect 9433 9165 9655 9170
rect 9433 9141 9446 9165
rect 9470 9146 9655 9165
rect 9679 9146 9792 9170
rect 9470 9141 9792 9146
rect 9433 9137 9792 9141
rect 9859 9167 10070 9173
rect 9859 9165 10020 9167
rect 9859 9145 9870 9165
rect 9890 9145 10020 9165
rect 9859 9138 10020 9145
rect 9859 9137 9900 9138
rect 9335 9111 9371 9136
rect 9183 9084 9220 9085
rect 9279 9084 9316 9085
rect 9335 9084 9342 9111
rect 7493 9025 7908 9060
rect 9083 9075 9221 9084
rect 9083 9055 9192 9075
rect 9212 9055 9221 9075
rect 9083 9048 9221 9055
rect 9279 9081 9342 9084
rect 9363 9084 9371 9111
rect 9390 9084 9427 9085
rect 9363 9081 9427 9084
rect 9279 9075 9427 9081
rect 9279 9055 9288 9075
rect 9308 9055 9398 9075
rect 9418 9055 9427 9075
rect 9083 9046 9179 9048
rect 9279 9045 9427 9055
rect 9486 9075 9523 9085
rect 9598 9084 9635 9085
rect 9579 9082 9635 9084
rect 9486 9055 9494 9075
rect 9514 9055 9523 9075
rect 9335 9044 9371 9045
rect 7493 9024 7539 9025
rect 7199 8979 7449 8981
rect 7199 8976 7300 8979
rect 7199 8957 7264 8976
rect 7261 8949 7264 8957
rect 7293 8949 7300 8976
rect 7328 8952 7338 8979
rect 7367 8957 7449 8979
rect 7833 8973 7908 9025
rect 7367 8952 7371 8957
rect 7328 8949 7371 8952
rect 7261 8935 7371 8949
rect 6687 8917 7028 8918
rect 6612 8912 7028 8917
rect 6612 8892 6615 8912
rect 6635 8892 7029 8912
rect 5669 8245 6475 8320
rect 4908 8201 4917 8235
rect 4946 8234 5356 8235
rect 4946 8201 4963 8234
rect 5188 8233 5356 8234
rect 4908 8175 4963 8201
rect 4908 8141 4916 8175
rect 4945 8141 4963 8175
rect 4908 8129 4963 8141
rect 3104 8084 3188 8105
rect 3104 8056 3132 8084
rect 3176 8056 3188 8084
rect 2918 8005 2992 8033
rect 2918 7957 2941 8005
rect 2978 7957 2992 8005
rect 3104 8027 3188 8056
rect 3104 7999 3129 8027
rect 3173 7999 3188 8027
rect 3104 7974 3188 7999
rect 5244 7988 5332 7992
rect 2918 7948 2992 7957
rect 551 7898 617 7946
rect 2928 7944 2992 7948
rect 5244 7971 5508 7988
rect 5244 7917 5424 7971
rect 5487 7917 5508 7971
rect 3141 7907 3852 7909
rect 2514 7906 3852 7907
rect 1464 7905 1536 7906
rect 551 7824 610 7898
rect 1463 7897 1562 7905
rect 1463 7894 1515 7897
rect 1463 7859 1471 7894
rect 1496 7859 1515 7894
rect 1540 7886 1562 7897
rect 2513 7898 3852 7906
rect 2513 7895 2565 7898
rect 1540 7885 2407 7886
rect 1540 7859 2408 7885
rect 1463 7849 2408 7859
rect 1463 7847 1562 7849
rect 551 7806 573 7824
rect 591 7806 610 7824
rect 551 7784 610 7806
rect 818 7820 1350 7825
rect 818 7800 1704 7820
rect 1724 7800 1727 7820
rect 2363 7816 2408 7849
rect 2513 7860 2521 7895
rect 2546 7860 2565 7895
rect 2590 7860 3852 7898
rect 2513 7851 3852 7860
rect 2513 7848 2602 7851
rect 3141 7849 3852 7851
rect 5244 7900 5508 7917
rect 818 7796 1727 7800
rect 818 7749 861 7796
rect 1311 7795 1727 7796
rect 2359 7796 2752 7816
rect 2772 7796 2775 7816
rect 1311 7794 1652 7795
rect 968 7763 1078 7777
rect 968 7760 1011 7763
rect 968 7755 972 7760
rect 806 7748 861 7749
rect 550 7725 861 7748
rect 550 7707 575 7725
rect 593 7713 861 7725
rect 890 7733 972 7755
rect 1001 7733 1011 7760
rect 1039 7736 1046 7763
rect 1075 7755 1078 7763
rect 1075 7736 1140 7755
rect 1039 7733 1140 7736
rect 890 7731 1140 7733
rect 593 7707 615 7713
rect 550 7568 615 7707
rect 890 7652 927 7731
rect 968 7718 1078 7731
rect 1042 7662 1073 7663
rect 890 7632 899 7652
rect 919 7632 927 7652
rect 550 7550 573 7568
rect 591 7550 615 7568
rect 550 7533 615 7550
rect 770 7614 838 7627
rect 890 7622 927 7632
rect 986 7652 1073 7662
rect 986 7632 995 7652
rect 1015 7632 1073 7652
rect 986 7623 1073 7632
rect 986 7622 1023 7623
rect 770 7572 777 7614
rect 826 7572 838 7614
rect 770 7569 838 7572
rect 1042 7570 1073 7623
rect 1103 7652 1140 7731
rect 1255 7662 1286 7663
rect 1103 7632 1112 7652
rect 1132 7632 1140 7652
rect 1103 7622 1140 7632
rect 1199 7655 1286 7662
rect 1199 7652 1260 7655
rect 1199 7632 1208 7652
rect 1228 7635 1260 7652
rect 1281 7635 1286 7655
rect 1228 7632 1286 7635
rect 1199 7625 1286 7632
rect 1311 7652 1348 7794
rect 1614 7793 1651 7794
rect 2359 7791 2775 7796
rect 2359 7790 2700 7791
rect 2016 7759 2126 7773
rect 2016 7756 2059 7759
rect 2016 7751 2020 7756
rect 1938 7729 2020 7751
rect 2049 7729 2059 7756
rect 2087 7732 2094 7759
rect 2123 7751 2126 7759
rect 2123 7732 2188 7751
rect 2087 7729 2188 7732
rect 1938 7727 2188 7729
rect 1463 7662 1499 7663
rect 1311 7632 1320 7652
rect 1340 7632 1348 7652
rect 1199 7623 1255 7625
rect 1199 7622 1236 7623
rect 1311 7622 1348 7632
rect 1407 7652 1555 7662
rect 1655 7659 1751 7661
rect 1407 7632 1416 7652
rect 1436 7632 1526 7652
rect 1546 7632 1555 7652
rect 1407 7626 1555 7632
rect 1407 7623 1471 7626
rect 1407 7622 1444 7623
rect 1463 7596 1471 7623
rect 1492 7623 1555 7626
rect 1613 7652 1751 7659
rect 1613 7632 1622 7652
rect 1642 7632 1751 7652
rect 1613 7623 1751 7632
rect 1938 7648 1975 7727
rect 2016 7714 2126 7727
rect 2090 7658 2121 7659
rect 1938 7628 1947 7648
rect 1967 7628 1975 7648
rect 1492 7596 1499 7623
rect 1518 7622 1555 7623
rect 1614 7622 1651 7623
rect 1463 7571 1499 7596
rect 934 7569 975 7570
rect 770 7562 975 7569
rect 770 7551 944 7562
rect 770 7518 778 7551
rect 771 7509 778 7518
rect 827 7542 944 7551
rect 964 7542 975 7562
rect 827 7534 975 7542
rect 1042 7566 1401 7570
rect 1042 7561 1364 7566
rect 1042 7537 1155 7561
rect 1179 7542 1364 7561
rect 1388 7542 1401 7566
rect 1179 7537 1401 7542
rect 1042 7534 1401 7537
rect 1463 7534 1498 7571
rect 1566 7568 1666 7571
rect 1566 7564 1633 7568
rect 1566 7538 1578 7564
rect 1604 7542 1633 7564
rect 1659 7542 1666 7568
rect 1604 7538 1666 7542
rect 1566 7534 1666 7538
rect 827 7518 838 7534
rect 827 7509 835 7518
rect 1042 7513 1073 7534
rect 1463 7513 1499 7534
rect 885 7512 922 7513
rect 550 7469 615 7488
rect 550 7451 575 7469
rect 593 7451 615 7469
rect 550 7250 615 7451
rect 771 7325 835 7509
rect 884 7503 922 7512
rect 884 7483 893 7503
rect 913 7483 922 7503
rect 884 7475 922 7483
rect 988 7507 1073 7513
rect 1098 7512 1135 7513
rect 988 7487 996 7507
rect 1016 7487 1073 7507
rect 988 7479 1073 7487
rect 1097 7503 1135 7512
rect 1097 7483 1106 7503
rect 1126 7483 1135 7503
rect 988 7478 1024 7479
rect 1097 7475 1135 7483
rect 1201 7507 1286 7513
rect 1306 7512 1343 7513
rect 1201 7487 1209 7507
rect 1229 7506 1286 7507
rect 1229 7487 1258 7506
rect 1201 7486 1258 7487
rect 1279 7486 1286 7506
rect 1201 7479 1286 7486
rect 1305 7503 1343 7512
rect 1305 7483 1314 7503
rect 1334 7483 1343 7503
rect 1201 7478 1237 7479
rect 1305 7475 1343 7483
rect 1409 7507 1553 7513
rect 1409 7487 1417 7507
rect 1437 7487 1525 7507
rect 1545 7487 1553 7507
rect 1409 7479 1553 7487
rect 1409 7478 1445 7479
rect 1517 7478 1553 7479
rect 1619 7512 1656 7513
rect 1619 7511 1657 7512
rect 1619 7503 1683 7511
rect 1619 7483 1628 7503
rect 1648 7489 1683 7503
rect 1703 7489 1706 7509
rect 1648 7484 1706 7489
rect 1648 7483 1683 7484
rect 885 7446 922 7475
rect 886 7444 922 7446
rect 1098 7444 1135 7475
rect 886 7422 1135 7444
rect 967 7416 1078 7422
rect 967 7408 1008 7416
rect 967 7388 975 7408
rect 994 7388 1008 7408
rect 967 7386 1008 7388
rect 1036 7408 1078 7416
rect 1036 7388 1052 7408
rect 1071 7388 1078 7408
rect 1036 7386 1078 7388
rect 967 7371 1078 7386
rect 771 7315 839 7325
rect 771 7282 788 7315
rect 828 7282 839 7315
rect 771 7270 839 7282
rect 771 7268 835 7270
rect 1306 7251 1343 7475
rect 1619 7471 1683 7483
rect 1723 7253 1750 7623
rect 1938 7618 1975 7628
rect 2034 7648 2121 7658
rect 2034 7628 2043 7648
rect 2063 7628 2121 7648
rect 2034 7619 2121 7628
rect 2034 7618 2071 7619
rect 1814 7605 1884 7610
rect 1809 7599 1884 7605
rect 1809 7566 1817 7599
rect 1870 7566 1884 7599
rect 2090 7566 2121 7619
rect 2151 7648 2188 7727
rect 2303 7658 2334 7659
rect 2151 7628 2160 7648
rect 2180 7628 2188 7648
rect 2151 7618 2188 7628
rect 2247 7651 2334 7658
rect 2247 7648 2308 7651
rect 2247 7628 2256 7648
rect 2276 7631 2308 7648
rect 2329 7631 2334 7651
rect 2276 7628 2334 7631
rect 2247 7621 2334 7628
rect 2359 7648 2396 7790
rect 2662 7789 2699 7790
rect 2511 7658 2547 7659
rect 2359 7628 2368 7648
rect 2388 7628 2396 7648
rect 2247 7619 2303 7621
rect 2247 7618 2284 7619
rect 2359 7618 2396 7628
rect 2455 7648 2603 7658
rect 2703 7655 2799 7657
rect 2455 7628 2464 7648
rect 2484 7628 2574 7648
rect 2594 7628 2603 7648
rect 2455 7622 2603 7628
rect 2455 7619 2519 7622
rect 2455 7618 2492 7619
rect 2511 7592 2519 7619
rect 2540 7619 2603 7622
rect 2661 7648 2799 7655
rect 2661 7628 2670 7648
rect 2690 7628 2799 7648
rect 2661 7619 2799 7628
rect 2540 7592 2547 7619
rect 2566 7618 2603 7619
rect 2662 7618 2699 7619
rect 2511 7567 2547 7592
rect 1809 7565 1892 7566
rect 1982 7565 2023 7566
rect 1809 7558 2023 7565
rect 1809 7541 1992 7558
rect 1809 7508 1822 7541
rect 1875 7538 1992 7541
rect 2012 7538 2023 7558
rect 1875 7530 2023 7538
rect 2090 7562 2449 7566
rect 2090 7557 2412 7562
rect 2090 7533 2203 7557
rect 2227 7538 2412 7557
rect 2436 7538 2449 7562
rect 2227 7533 2449 7538
rect 2090 7530 2449 7533
rect 2511 7530 2546 7567
rect 2614 7564 2714 7567
rect 2614 7560 2681 7564
rect 2614 7534 2626 7560
rect 2652 7538 2681 7560
rect 2707 7538 2714 7564
rect 2652 7534 2714 7538
rect 2614 7530 2714 7534
rect 1875 7508 1892 7530
rect 2090 7509 2121 7530
rect 2511 7509 2547 7530
rect 1933 7508 1970 7509
rect 1809 7494 1892 7508
rect 1582 7251 1750 7253
rect 1306 7250 1750 7251
rect 550 7220 1750 7250
rect 1820 7284 1892 7494
rect 1932 7499 1970 7508
rect 1932 7479 1941 7499
rect 1961 7479 1970 7499
rect 1932 7471 1970 7479
rect 2036 7503 2121 7509
rect 2146 7508 2183 7509
rect 2036 7483 2044 7503
rect 2064 7483 2121 7503
rect 2036 7475 2121 7483
rect 2145 7499 2183 7508
rect 2145 7479 2154 7499
rect 2174 7479 2183 7499
rect 2036 7474 2072 7475
rect 2145 7471 2183 7479
rect 2249 7503 2334 7509
rect 2354 7508 2391 7509
rect 2249 7483 2257 7503
rect 2277 7502 2334 7503
rect 2277 7483 2306 7502
rect 2249 7482 2306 7483
rect 2327 7482 2334 7502
rect 2249 7475 2334 7482
rect 2353 7499 2391 7508
rect 2353 7479 2362 7499
rect 2382 7479 2391 7499
rect 2249 7474 2285 7475
rect 2353 7471 2391 7479
rect 2457 7503 2601 7509
rect 2457 7483 2465 7503
rect 2485 7483 2573 7503
rect 2593 7483 2601 7503
rect 2457 7475 2601 7483
rect 2457 7474 2493 7475
rect 2565 7474 2601 7475
rect 2667 7508 2704 7509
rect 2667 7507 2705 7508
rect 2667 7499 2731 7507
rect 2667 7479 2676 7499
rect 2696 7485 2731 7499
rect 2751 7485 2754 7505
rect 2696 7480 2754 7485
rect 2696 7479 2731 7480
rect 1933 7442 1970 7471
rect 1934 7440 1970 7442
rect 2146 7440 2183 7471
rect 1934 7418 2183 7440
rect 2015 7412 2126 7418
rect 2015 7404 2056 7412
rect 2015 7384 2023 7404
rect 2042 7384 2056 7404
rect 2015 7382 2056 7384
rect 2084 7404 2126 7412
rect 2084 7384 2100 7404
rect 2119 7384 2126 7404
rect 2084 7382 2126 7384
rect 2015 7367 2126 7382
rect 1820 7245 1839 7284
rect 1884 7245 1892 7284
rect 1820 7228 1892 7245
rect 2354 7272 2391 7471
rect 2667 7467 2731 7479
rect 2354 7266 2395 7272
rect 2771 7268 2798 7619
rect 3093 7606 3188 7632
rect 2929 7584 2993 7603
rect 2929 7545 2942 7584
rect 2976 7545 2993 7584
rect 2929 7526 2993 7545
rect 2630 7266 2798 7268
rect 2354 7240 2798 7266
rect 550 7173 615 7220
rect 550 7155 573 7173
rect 591 7155 615 7173
rect 1463 7200 1498 7202
rect 1463 7198 1567 7200
rect 2356 7198 2395 7240
rect 2630 7239 2798 7240
rect 1463 7191 2397 7198
rect 1463 7190 1514 7191
rect 1463 7170 1466 7190
rect 1491 7171 1514 7190
rect 1546 7171 2397 7191
rect 1491 7170 2397 7171
rect 1463 7163 2397 7170
rect 1736 7162 2397 7163
rect 550 7134 615 7155
rect 827 7145 867 7148
rect 827 7141 1730 7145
rect 827 7121 1704 7141
rect 1724 7121 1730 7141
rect 827 7118 1730 7121
rect 551 7074 616 7094
rect 551 7056 575 7074
rect 593 7056 616 7074
rect 551 7029 616 7056
rect 827 7029 867 7118
rect 1311 7116 1727 7118
rect 1311 7115 1652 7116
rect 968 7084 1078 7098
rect 968 7081 1011 7084
rect 968 7076 972 7081
rect 550 6994 867 7029
rect 890 7054 972 7076
rect 1001 7054 1011 7081
rect 1039 7057 1046 7084
rect 1075 7076 1078 7084
rect 1075 7057 1140 7076
rect 1039 7054 1140 7057
rect 890 7052 1140 7054
rect 551 6918 616 6994
rect 890 6973 927 7052
rect 968 7039 1078 7052
rect 1042 6983 1073 6984
rect 890 6953 899 6973
rect 919 6953 927 6973
rect 890 6943 927 6953
rect 986 6973 1073 6983
rect 986 6953 995 6973
rect 1015 6953 1073 6973
rect 986 6944 1073 6953
rect 986 6943 1023 6944
rect 551 6900 573 6918
rect 591 6900 616 6918
rect 551 6879 616 6900
rect 764 6898 829 6907
rect 764 6861 774 6898
rect 814 6890 829 6898
rect 1042 6891 1073 6944
rect 1103 6973 1140 7052
rect 1255 6983 1286 6984
rect 1103 6953 1112 6973
rect 1132 6953 1140 6973
rect 1103 6943 1140 6953
rect 1199 6976 1286 6983
rect 1199 6973 1260 6976
rect 1199 6953 1208 6973
rect 1228 6956 1260 6973
rect 1281 6956 1286 6976
rect 1228 6953 1286 6956
rect 1199 6946 1286 6953
rect 1311 6973 1348 7115
rect 1614 7114 1651 7115
rect 2931 7055 2993 7526
rect 3093 7565 3119 7606
rect 3155 7565 3188 7606
rect 3093 7269 3188 7565
rect 3093 7225 3108 7269
rect 3168 7225 3188 7269
rect 3093 7205 3188 7225
rect 3805 7136 3848 7849
rect 3805 7116 4199 7136
rect 4219 7116 4222 7136
rect 3806 7111 4222 7116
rect 3806 7110 4147 7111
rect 3463 7079 3573 7093
rect 3463 7076 3506 7079
rect 3463 7071 3467 7076
rect 2926 7003 3001 7055
rect 3385 7049 3467 7071
rect 3496 7049 3506 7076
rect 3534 7052 3541 7079
rect 3570 7071 3573 7079
rect 3570 7052 3635 7071
rect 3534 7049 3635 7052
rect 3385 7047 3635 7049
rect 3295 7003 3341 7004
rect 1463 6983 1499 6984
rect 1311 6953 1320 6973
rect 1340 6953 1348 6973
rect 1199 6944 1255 6946
rect 1199 6943 1236 6944
rect 1311 6943 1348 6953
rect 1407 6973 1555 6983
rect 1655 6980 1751 6982
rect 1407 6953 1416 6973
rect 1436 6953 1526 6973
rect 1546 6953 1555 6973
rect 1407 6947 1555 6953
rect 1407 6944 1471 6947
rect 1407 6943 1444 6944
rect 1463 6917 1471 6944
rect 1492 6944 1555 6947
rect 1613 6973 1751 6980
rect 1613 6953 1622 6973
rect 1642 6953 1751 6973
rect 1613 6944 1751 6953
rect 2926 6968 3341 7003
rect 1492 6917 1499 6944
rect 1518 6943 1555 6944
rect 1614 6943 1651 6944
rect 1463 6892 1499 6917
rect 934 6890 975 6891
rect 814 6883 975 6890
rect 814 6863 944 6883
rect 964 6863 975 6883
rect 814 6861 975 6863
rect 764 6855 975 6861
rect 1042 6887 1401 6891
rect 1042 6882 1364 6887
rect 1042 6858 1155 6882
rect 1179 6863 1364 6882
rect 1388 6863 1401 6887
rect 1179 6858 1401 6863
rect 1042 6855 1401 6858
rect 1463 6855 1498 6892
rect 1566 6889 1666 6892
rect 1566 6885 1633 6889
rect 1566 6859 1578 6885
rect 1604 6863 1633 6885
rect 1659 6863 1666 6889
rect 1604 6859 1666 6863
rect 1566 6855 1666 6859
rect 764 6842 831 6855
rect 556 6819 612 6839
rect 556 6801 575 6819
rect 593 6801 612 6819
rect 556 6688 612 6801
rect 764 6821 778 6842
rect 814 6821 831 6842
rect 1042 6834 1073 6855
rect 1463 6834 1499 6855
rect 885 6833 922 6834
rect 764 6814 831 6821
rect 884 6824 922 6833
rect 556 6550 611 6688
rect 764 6662 829 6814
rect 884 6804 893 6824
rect 913 6804 922 6824
rect 884 6796 922 6804
rect 988 6828 1073 6834
rect 1098 6833 1135 6834
rect 988 6808 996 6828
rect 1016 6808 1073 6828
rect 988 6800 1073 6808
rect 1097 6824 1135 6833
rect 1097 6804 1106 6824
rect 1126 6804 1135 6824
rect 988 6799 1024 6800
rect 1097 6796 1135 6804
rect 1201 6828 1286 6834
rect 1306 6833 1343 6834
rect 1201 6808 1209 6828
rect 1229 6827 1286 6828
rect 1229 6808 1258 6827
rect 1201 6807 1258 6808
rect 1279 6807 1286 6827
rect 1201 6800 1286 6807
rect 1305 6824 1343 6833
rect 1305 6804 1314 6824
rect 1334 6804 1343 6824
rect 1201 6799 1237 6800
rect 1305 6796 1343 6804
rect 1409 6828 1553 6834
rect 1409 6808 1417 6828
rect 1437 6808 1525 6828
rect 1545 6808 1553 6828
rect 1409 6800 1553 6808
rect 1409 6799 1445 6800
rect 1517 6799 1553 6800
rect 1619 6833 1656 6834
rect 1619 6832 1657 6833
rect 1619 6824 1683 6832
rect 1619 6804 1628 6824
rect 1648 6810 1683 6824
rect 1703 6810 1706 6830
rect 1648 6805 1706 6810
rect 1648 6804 1683 6805
rect 885 6767 922 6796
rect 886 6765 922 6767
rect 1098 6765 1135 6796
rect 886 6743 1135 6765
rect 967 6737 1078 6743
rect 967 6729 1008 6737
rect 967 6709 975 6729
rect 994 6709 1008 6729
rect 967 6707 1008 6709
rect 1036 6729 1078 6737
rect 1036 6709 1052 6729
rect 1071 6709 1078 6729
rect 1036 6707 1078 6709
rect 967 6694 1078 6707
rect 1306 6697 1343 6796
rect 1619 6792 1683 6804
rect 757 6652 878 6662
rect 757 6650 826 6652
rect 757 6609 770 6650
rect 807 6611 826 6650
rect 863 6611 878 6652
rect 807 6609 878 6611
rect 757 6591 878 6609
rect 549 6547 613 6550
rect 969 6547 1073 6553
rect 1304 6547 1345 6697
rect 1723 6689 1750 6944
rect 1812 6934 1892 6945
rect 1812 6908 1829 6934
rect 1869 6908 1892 6934
rect 1812 6881 1892 6908
rect 1812 6855 1833 6881
rect 1873 6855 1892 6881
rect 1812 6836 1892 6855
rect 1812 6810 1836 6836
rect 1876 6810 1892 6836
rect 1812 6759 1892 6810
rect 549 6544 1345 6547
rect 1724 6558 1750 6689
rect 1724 6544 1752 6558
rect 549 6509 1752 6544
rect 1814 6551 1884 6759
rect 2926 6684 3001 6968
rect 3295 6885 3341 6968
rect 3385 6968 3422 7047
rect 3463 7034 3573 7047
rect 3537 6978 3568 6979
rect 3385 6948 3394 6968
rect 3414 6948 3422 6968
rect 3385 6938 3422 6948
rect 3481 6968 3568 6978
rect 3481 6948 3490 6968
rect 3510 6948 3568 6968
rect 3481 6939 3568 6948
rect 3481 6938 3518 6939
rect 3537 6886 3568 6939
rect 3598 6968 3635 7047
rect 3750 6978 3781 6979
rect 3598 6948 3607 6968
rect 3627 6948 3635 6968
rect 3598 6938 3635 6948
rect 3694 6971 3781 6978
rect 3694 6968 3755 6971
rect 3694 6948 3703 6968
rect 3723 6951 3755 6968
rect 3776 6951 3781 6971
rect 3723 6948 3781 6951
rect 3694 6941 3781 6948
rect 3806 6968 3843 7110
rect 4109 7109 4146 7110
rect 3958 6978 3994 6979
rect 3806 6948 3815 6968
rect 3835 6948 3843 6968
rect 3694 6939 3750 6941
rect 3694 6938 3731 6939
rect 3806 6938 3843 6948
rect 3902 6968 4050 6978
rect 4150 6975 4246 6977
rect 3902 6948 3911 6968
rect 3931 6948 4021 6968
rect 4041 6948 4050 6968
rect 3902 6942 4050 6948
rect 3902 6939 3966 6942
rect 3902 6938 3939 6939
rect 3958 6912 3966 6939
rect 3987 6939 4050 6942
rect 4108 6968 4246 6975
rect 4108 6948 4117 6968
rect 4137 6948 4246 6968
rect 4108 6939 4246 6948
rect 3987 6912 3994 6939
rect 4013 6938 4050 6939
rect 4109 6938 4146 6939
rect 3958 6887 3994 6912
rect 3429 6885 3470 6886
rect 3295 6878 3470 6885
rect 3093 6852 3179 6871
rect 3093 6811 3108 6852
rect 3162 6811 3179 6852
rect 3295 6858 3439 6878
rect 3459 6858 3470 6878
rect 3295 6850 3470 6858
rect 3537 6882 3896 6886
rect 3537 6877 3859 6882
rect 3537 6853 3650 6877
rect 3674 6858 3859 6877
rect 3883 6858 3896 6882
rect 3674 6853 3896 6858
rect 3537 6850 3896 6853
rect 3958 6850 3993 6887
rect 4061 6884 4161 6887
rect 4061 6880 4128 6884
rect 4061 6854 4073 6880
rect 4099 6858 4128 6880
rect 4154 6858 4161 6884
rect 4099 6854 4161 6858
rect 4061 6850 4161 6854
rect 3295 6846 3341 6850
rect 3537 6829 3568 6850
rect 3958 6829 3994 6850
rect 3380 6828 3417 6829
rect 3093 6775 3179 6811
rect 3379 6819 3417 6828
rect 3379 6799 3388 6819
rect 3408 6799 3417 6819
rect 3379 6791 3417 6799
rect 3483 6823 3568 6829
rect 3593 6828 3630 6829
rect 3483 6803 3491 6823
rect 3511 6803 3568 6823
rect 3483 6795 3568 6803
rect 3592 6819 3630 6828
rect 3592 6799 3601 6819
rect 3621 6799 3630 6819
rect 3483 6794 3519 6795
rect 3592 6791 3630 6799
rect 3696 6823 3781 6829
rect 3801 6828 3838 6829
rect 3696 6803 3704 6823
rect 3724 6822 3781 6823
rect 3724 6803 3753 6822
rect 3696 6802 3753 6803
rect 3774 6802 3781 6822
rect 3696 6795 3781 6802
rect 3800 6819 3838 6828
rect 3800 6799 3809 6819
rect 3829 6799 3838 6819
rect 3696 6794 3732 6795
rect 3800 6791 3838 6799
rect 3904 6823 4048 6829
rect 3904 6803 3912 6823
rect 3932 6803 4020 6823
rect 4040 6803 4048 6823
rect 3904 6795 4048 6803
rect 3904 6794 3940 6795
rect 549 6448 613 6509
rect 969 6507 1073 6509
rect 1304 6507 1345 6509
rect 1814 6506 1835 6551
rect 1815 6485 1835 6506
rect 1865 6506 1884 6551
rect 2921 6642 3001 6684
rect 1865 6485 1882 6506
rect 1815 6466 1882 6485
rect 1464 6458 1536 6459
rect 1463 6450 1562 6458
rect 551 6377 610 6448
rect 1463 6447 1515 6450
rect 1463 6412 1471 6447
rect 1496 6412 1515 6447
rect 1540 6439 1562 6450
rect 1540 6438 2407 6439
rect 1540 6412 2408 6438
rect 1463 6402 2408 6412
rect 1463 6400 1562 6402
rect 551 6359 573 6377
rect 591 6359 610 6377
rect 551 6337 610 6359
rect 818 6373 1350 6378
rect 818 6353 1704 6373
rect 1724 6353 1727 6373
rect 2363 6369 2408 6402
rect 818 6349 1727 6353
rect 818 6302 861 6349
rect 1311 6348 1727 6349
rect 2359 6349 2752 6369
rect 2772 6349 2775 6369
rect 1311 6347 1652 6348
rect 968 6316 1078 6330
rect 968 6313 1011 6316
rect 968 6308 972 6313
rect 806 6301 861 6302
rect 550 6278 861 6301
rect 550 6260 575 6278
rect 593 6266 861 6278
rect 890 6286 972 6308
rect 1001 6286 1011 6313
rect 1039 6289 1046 6316
rect 1075 6308 1078 6316
rect 1075 6289 1140 6308
rect 1039 6286 1140 6289
rect 890 6284 1140 6286
rect 593 6260 615 6266
rect 550 6121 615 6260
rect 890 6205 927 6284
rect 968 6271 1078 6284
rect 1042 6215 1073 6216
rect 890 6185 899 6205
rect 919 6185 927 6205
rect 550 6103 573 6121
rect 591 6103 615 6121
rect 550 6086 615 6103
rect 770 6167 838 6180
rect 890 6175 927 6185
rect 986 6205 1073 6215
rect 986 6185 995 6205
rect 1015 6185 1073 6205
rect 986 6176 1073 6185
rect 986 6175 1023 6176
rect 770 6125 777 6167
rect 826 6125 838 6167
rect 770 6122 838 6125
rect 1042 6123 1073 6176
rect 1103 6205 1140 6284
rect 1255 6215 1286 6216
rect 1103 6185 1112 6205
rect 1132 6185 1140 6205
rect 1103 6175 1140 6185
rect 1199 6208 1286 6215
rect 1199 6205 1260 6208
rect 1199 6185 1208 6205
rect 1228 6188 1260 6205
rect 1281 6188 1286 6208
rect 1228 6185 1286 6188
rect 1199 6178 1286 6185
rect 1311 6205 1348 6347
rect 1614 6346 1651 6347
rect 2359 6344 2775 6349
rect 2359 6343 2700 6344
rect 2016 6312 2126 6326
rect 2016 6309 2059 6312
rect 2016 6304 2020 6309
rect 1938 6282 2020 6304
rect 2049 6282 2059 6309
rect 2087 6285 2094 6312
rect 2123 6304 2126 6312
rect 2123 6285 2188 6304
rect 2087 6282 2188 6285
rect 1938 6280 2188 6282
rect 1463 6215 1499 6216
rect 1311 6185 1320 6205
rect 1340 6185 1348 6205
rect 1199 6176 1255 6178
rect 1199 6175 1236 6176
rect 1311 6175 1348 6185
rect 1407 6205 1555 6215
rect 1655 6212 1751 6214
rect 1407 6185 1416 6205
rect 1436 6185 1526 6205
rect 1546 6185 1555 6205
rect 1407 6179 1555 6185
rect 1407 6176 1471 6179
rect 1407 6175 1444 6176
rect 1463 6149 1471 6176
rect 1492 6176 1555 6179
rect 1613 6205 1751 6212
rect 1613 6185 1622 6205
rect 1642 6185 1751 6205
rect 1613 6176 1751 6185
rect 1938 6201 1975 6280
rect 2016 6267 2126 6280
rect 2090 6211 2121 6212
rect 1938 6181 1947 6201
rect 1967 6181 1975 6201
rect 1492 6149 1499 6176
rect 1518 6175 1555 6176
rect 1614 6175 1651 6176
rect 1463 6124 1499 6149
rect 934 6122 975 6123
rect 770 6115 975 6122
rect 770 6104 944 6115
rect 770 6071 778 6104
rect 771 6062 778 6071
rect 827 6095 944 6104
rect 964 6095 975 6115
rect 827 6087 975 6095
rect 1042 6119 1401 6123
rect 1042 6114 1364 6119
rect 1042 6090 1155 6114
rect 1179 6095 1364 6114
rect 1388 6095 1401 6119
rect 1179 6090 1401 6095
rect 1042 6087 1401 6090
rect 1463 6087 1498 6124
rect 1566 6121 1666 6124
rect 1566 6117 1633 6121
rect 1566 6091 1578 6117
rect 1604 6095 1633 6117
rect 1659 6095 1666 6121
rect 1604 6091 1666 6095
rect 1566 6087 1666 6091
rect 827 6071 838 6087
rect 827 6062 835 6071
rect 1042 6066 1073 6087
rect 1463 6066 1499 6087
rect 885 6065 922 6066
rect 550 6022 615 6041
rect 550 6004 575 6022
rect 593 6004 615 6022
rect 550 5803 615 6004
rect 771 5878 835 6062
rect 884 6056 922 6065
rect 884 6036 893 6056
rect 913 6036 922 6056
rect 884 6028 922 6036
rect 988 6060 1073 6066
rect 1098 6065 1135 6066
rect 988 6040 996 6060
rect 1016 6040 1073 6060
rect 988 6032 1073 6040
rect 1097 6056 1135 6065
rect 1097 6036 1106 6056
rect 1126 6036 1135 6056
rect 988 6031 1024 6032
rect 1097 6028 1135 6036
rect 1201 6060 1286 6066
rect 1306 6065 1343 6066
rect 1201 6040 1209 6060
rect 1229 6059 1286 6060
rect 1229 6040 1258 6059
rect 1201 6039 1258 6040
rect 1279 6039 1286 6059
rect 1201 6032 1286 6039
rect 1305 6056 1343 6065
rect 1305 6036 1314 6056
rect 1334 6036 1343 6056
rect 1201 6031 1237 6032
rect 1305 6028 1343 6036
rect 1409 6060 1553 6066
rect 1409 6040 1417 6060
rect 1437 6040 1525 6060
rect 1545 6040 1553 6060
rect 1409 6032 1553 6040
rect 1409 6031 1445 6032
rect 1517 6031 1553 6032
rect 1619 6065 1656 6066
rect 1619 6064 1657 6065
rect 1619 6056 1683 6064
rect 1619 6036 1628 6056
rect 1648 6042 1683 6056
rect 1703 6042 1706 6062
rect 1648 6037 1706 6042
rect 1648 6036 1683 6037
rect 885 5999 922 6028
rect 886 5997 922 5999
rect 1098 5997 1135 6028
rect 886 5975 1135 5997
rect 967 5969 1078 5975
rect 967 5961 1008 5969
rect 967 5941 975 5961
rect 994 5941 1008 5961
rect 967 5939 1008 5941
rect 1036 5961 1078 5969
rect 1036 5941 1052 5961
rect 1071 5941 1078 5961
rect 1036 5939 1078 5941
rect 967 5924 1078 5939
rect 771 5868 839 5878
rect 771 5835 788 5868
rect 828 5835 839 5868
rect 771 5823 839 5835
rect 771 5821 835 5823
rect 1306 5804 1343 6028
rect 1619 6024 1683 6036
rect 1723 5806 1750 6176
rect 1938 6171 1975 6181
rect 2034 6201 2121 6211
rect 2034 6181 2043 6201
rect 2063 6181 2121 6201
rect 2034 6172 2121 6181
rect 2034 6171 2071 6172
rect 1814 6158 1884 6163
rect 1809 6152 1884 6158
rect 1809 6119 1817 6152
rect 1870 6119 1884 6152
rect 2090 6119 2121 6172
rect 2151 6201 2188 6280
rect 2303 6211 2334 6212
rect 2151 6181 2160 6201
rect 2180 6181 2188 6201
rect 2151 6171 2188 6181
rect 2247 6204 2334 6211
rect 2247 6201 2308 6204
rect 2247 6181 2256 6201
rect 2276 6184 2308 6201
rect 2329 6184 2334 6204
rect 2276 6181 2334 6184
rect 2247 6174 2334 6181
rect 2359 6201 2396 6343
rect 2662 6342 2699 6343
rect 2511 6211 2547 6212
rect 2359 6181 2368 6201
rect 2388 6181 2396 6201
rect 2247 6172 2303 6174
rect 2247 6171 2284 6172
rect 2359 6171 2396 6181
rect 2455 6201 2603 6211
rect 2703 6208 2799 6210
rect 2455 6181 2464 6201
rect 2484 6181 2574 6201
rect 2594 6181 2603 6201
rect 2455 6175 2603 6181
rect 2455 6172 2519 6175
rect 2455 6171 2492 6172
rect 2511 6145 2519 6172
rect 2540 6172 2603 6175
rect 2661 6201 2799 6208
rect 2661 6181 2670 6201
rect 2690 6181 2799 6201
rect 2661 6172 2799 6181
rect 2540 6145 2547 6172
rect 2566 6171 2603 6172
rect 2662 6171 2699 6172
rect 2511 6120 2547 6145
rect 1809 6118 1892 6119
rect 1982 6118 2023 6119
rect 1809 6111 2023 6118
rect 1809 6094 1992 6111
rect 1809 6061 1822 6094
rect 1875 6091 1992 6094
rect 2012 6091 2023 6111
rect 1875 6083 2023 6091
rect 2090 6115 2449 6119
rect 2090 6110 2412 6115
rect 2090 6086 2203 6110
rect 2227 6091 2412 6110
rect 2436 6091 2449 6115
rect 2227 6086 2449 6091
rect 2090 6083 2449 6086
rect 2511 6083 2546 6120
rect 2614 6117 2714 6120
rect 2614 6113 2681 6117
rect 2614 6087 2626 6113
rect 2652 6091 2681 6113
rect 2707 6091 2714 6117
rect 2652 6087 2714 6091
rect 2614 6083 2714 6087
rect 1875 6061 1892 6083
rect 2090 6062 2121 6083
rect 2511 6062 2547 6083
rect 1933 6061 1970 6062
rect 1809 6047 1892 6061
rect 1582 5804 1750 5806
rect 1306 5803 1750 5804
rect 550 5773 1750 5803
rect 1820 5837 1892 6047
rect 1932 6052 1970 6061
rect 1932 6032 1941 6052
rect 1961 6032 1970 6052
rect 1932 6024 1970 6032
rect 2036 6056 2121 6062
rect 2146 6061 2183 6062
rect 2036 6036 2044 6056
rect 2064 6036 2121 6056
rect 2036 6028 2121 6036
rect 2145 6052 2183 6061
rect 2145 6032 2154 6052
rect 2174 6032 2183 6052
rect 2036 6027 2072 6028
rect 2145 6024 2183 6032
rect 2249 6056 2334 6062
rect 2354 6061 2391 6062
rect 2249 6036 2257 6056
rect 2277 6055 2334 6056
rect 2277 6036 2306 6055
rect 2249 6035 2306 6036
rect 2327 6035 2334 6055
rect 2249 6028 2334 6035
rect 2353 6052 2391 6061
rect 2353 6032 2362 6052
rect 2382 6032 2391 6052
rect 2249 6027 2285 6028
rect 2353 6024 2391 6032
rect 2457 6056 2601 6062
rect 2457 6036 2465 6056
rect 2485 6036 2573 6056
rect 2593 6036 2601 6056
rect 2457 6028 2601 6036
rect 2457 6027 2493 6028
rect 2565 6027 2601 6028
rect 2667 6061 2704 6062
rect 2667 6060 2705 6061
rect 2667 6052 2731 6060
rect 2667 6032 2676 6052
rect 2696 6038 2731 6052
rect 2751 6038 2754 6058
rect 2696 6033 2754 6038
rect 2696 6032 2731 6033
rect 1933 5995 1970 6024
rect 1934 5993 1970 5995
rect 2146 5993 2183 6024
rect 1934 5971 2183 5993
rect 2015 5965 2126 5971
rect 2015 5957 2056 5965
rect 2015 5937 2023 5957
rect 2042 5937 2056 5957
rect 2015 5935 2056 5937
rect 2084 5957 2126 5965
rect 2084 5937 2100 5957
rect 2119 5937 2126 5957
rect 2084 5935 2126 5937
rect 2015 5920 2126 5935
rect 1820 5798 1839 5837
rect 1884 5798 1892 5837
rect 1820 5781 1892 5798
rect 2354 5825 2391 6024
rect 2667 6020 2731 6032
rect 2354 5819 2395 5825
rect 2771 5821 2798 6172
rect 2921 6042 3000 6642
rect 3097 6190 3176 6775
rect 3380 6762 3417 6791
rect 3381 6760 3417 6762
rect 3593 6760 3630 6791
rect 3381 6738 3630 6760
rect 3462 6732 3573 6738
rect 3462 6724 3503 6732
rect 3462 6704 3470 6724
rect 3489 6704 3503 6724
rect 3462 6702 3503 6704
rect 3531 6724 3573 6732
rect 3531 6704 3547 6724
rect 3566 6704 3573 6724
rect 3531 6702 3573 6704
rect 3462 6687 3573 6702
rect 3801 6676 3838 6791
rect 3794 6564 3841 6676
rect 3962 6636 3992 6795
rect 4012 6794 4048 6795
rect 4114 6828 4151 6829
rect 4114 6827 4152 6828
rect 4114 6819 4178 6827
rect 4114 6799 4123 6819
rect 4143 6805 4178 6819
rect 4198 6805 4201 6825
rect 4143 6800 4201 6805
rect 4143 6799 4178 6800
rect 4114 6787 4178 6799
rect 3962 6632 4048 6636
rect 3962 6614 3977 6632
rect 4029 6614 4048 6632
rect 3962 6605 4048 6614
rect 4218 6566 4245 6939
rect 4077 6564 4245 6566
rect 3794 6538 4245 6564
rect 3794 6460 3841 6538
rect 4077 6537 4245 6538
rect 3739 6459 3841 6460
rect 3738 6451 3841 6459
rect 3738 6448 3790 6451
rect 3738 6413 3746 6448
rect 3771 6413 3790 6448
rect 3815 6413 3841 6451
rect 3738 6407 3841 6413
rect 4001 6452 4037 6456
rect 4001 6429 4009 6452
rect 4033 6429 4037 6452
rect 4001 6408 4037 6429
rect 3738 6403 3837 6407
rect 4001 6385 4009 6408
rect 4033 6385 4037 6408
rect 2630 5819 2798 5821
rect 2354 5793 2798 5819
rect 550 5726 615 5773
rect 550 5708 573 5726
rect 591 5708 615 5726
rect 1463 5753 1498 5755
rect 1463 5751 1567 5753
rect 2356 5751 2395 5793
rect 2630 5792 2798 5793
rect 1463 5744 2397 5751
rect 1463 5743 1514 5744
rect 1463 5723 1466 5743
rect 1491 5724 1514 5743
rect 1546 5724 2397 5744
rect 1491 5723 2397 5724
rect 1463 5716 2397 5723
rect 1736 5715 2397 5716
rect 550 5687 615 5708
rect 827 5698 867 5701
rect 827 5694 1730 5698
rect 827 5674 1704 5694
rect 1724 5674 1730 5694
rect 827 5671 1730 5674
rect 551 5627 616 5647
rect 551 5609 575 5627
rect 593 5609 616 5627
rect 551 5582 616 5609
rect 827 5582 867 5671
rect 1311 5669 1727 5671
rect 1311 5668 1652 5669
rect 968 5637 1078 5651
rect 968 5634 1011 5637
rect 968 5629 972 5634
rect 550 5547 867 5582
rect 890 5607 972 5629
rect 1001 5607 1011 5634
rect 1039 5610 1046 5637
rect 1075 5629 1078 5637
rect 1075 5610 1140 5629
rect 1039 5607 1140 5610
rect 890 5605 1140 5607
rect 551 5471 616 5547
rect 890 5526 927 5605
rect 968 5592 1078 5605
rect 1042 5536 1073 5537
rect 890 5506 899 5526
rect 919 5506 927 5526
rect 890 5496 927 5506
rect 986 5526 1073 5536
rect 986 5506 995 5526
rect 1015 5506 1073 5526
rect 986 5497 1073 5506
rect 986 5496 1023 5497
rect 551 5453 573 5471
rect 591 5453 616 5471
rect 551 5432 616 5453
rect 764 5451 829 5460
rect 764 5414 774 5451
rect 814 5443 829 5451
rect 1042 5444 1073 5497
rect 1103 5526 1140 5605
rect 1255 5536 1286 5537
rect 1103 5506 1112 5526
rect 1132 5506 1140 5526
rect 1103 5496 1140 5506
rect 1199 5529 1286 5536
rect 1199 5526 1260 5529
rect 1199 5506 1208 5526
rect 1228 5509 1260 5526
rect 1281 5509 1286 5529
rect 1228 5506 1286 5509
rect 1199 5499 1286 5506
rect 1311 5526 1348 5668
rect 1614 5667 1651 5668
rect 1463 5536 1499 5537
rect 1311 5506 1320 5526
rect 1340 5506 1348 5526
rect 1199 5497 1255 5499
rect 1199 5496 1236 5497
rect 1311 5496 1348 5506
rect 1407 5526 1555 5536
rect 1655 5533 1751 5535
rect 1407 5506 1416 5526
rect 1436 5506 1526 5526
rect 1546 5506 1555 5526
rect 1407 5500 1555 5506
rect 1407 5497 1471 5500
rect 1407 5496 1444 5497
rect 1463 5470 1471 5497
rect 1492 5497 1555 5500
rect 1613 5526 1751 5533
rect 1613 5506 1622 5526
rect 1642 5506 1751 5526
rect 1613 5497 1751 5506
rect 1492 5470 1499 5497
rect 1518 5496 1555 5497
rect 1614 5496 1651 5497
rect 1463 5445 1499 5470
rect 934 5443 975 5444
rect 814 5436 975 5443
rect 814 5416 944 5436
rect 964 5416 975 5436
rect 814 5414 975 5416
rect 764 5408 975 5414
rect 1042 5440 1401 5444
rect 1042 5435 1364 5440
rect 1042 5411 1155 5435
rect 1179 5416 1364 5435
rect 1388 5416 1401 5440
rect 1179 5411 1401 5416
rect 1042 5408 1401 5411
rect 1463 5408 1498 5445
rect 1566 5442 1666 5445
rect 1566 5438 1633 5442
rect 1566 5412 1578 5438
rect 1604 5416 1633 5438
rect 1659 5416 1666 5442
rect 1604 5412 1666 5416
rect 1566 5408 1666 5412
rect 764 5395 831 5408
rect 556 5372 612 5392
rect 556 5354 575 5372
rect 593 5354 612 5372
rect 556 5241 612 5354
rect 764 5374 778 5395
rect 814 5374 831 5395
rect 1042 5387 1073 5408
rect 1463 5387 1499 5408
rect 885 5386 922 5387
rect 764 5367 831 5374
rect 884 5377 922 5386
rect 556 5112 611 5241
rect 764 5215 829 5367
rect 884 5357 893 5377
rect 913 5357 922 5377
rect 884 5349 922 5357
rect 988 5381 1073 5387
rect 1098 5386 1135 5387
rect 988 5361 996 5381
rect 1016 5361 1073 5381
rect 988 5353 1073 5361
rect 1097 5377 1135 5386
rect 1097 5357 1106 5377
rect 1126 5357 1135 5377
rect 988 5352 1024 5353
rect 1097 5349 1135 5357
rect 1201 5381 1286 5387
rect 1306 5386 1343 5387
rect 1201 5361 1209 5381
rect 1229 5380 1286 5381
rect 1229 5361 1258 5380
rect 1201 5360 1258 5361
rect 1279 5360 1286 5380
rect 1201 5353 1286 5360
rect 1305 5377 1343 5386
rect 1305 5357 1314 5377
rect 1334 5357 1343 5377
rect 1201 5352 1237 5353
rect 1305 5349 1343 5357
rect 1409 5381 1553 5387
rect 1409 5361 1417 5381
rect 1437 5361 1525 5381
rect 1545 5361 1553 5381
rect 1409 5353 1553 5361
rect 1409 5352 1445 5353
rect 1517 5352 1553 5353
rect 1619 5386 1656 5387
rect 1619 5385 1657 5386
rect 1619 5377 1683 5385
rect 1619 5357 1628 5377
rect 1648 5363 1683 5377
rect 1703 5363 1706 5383
rect 1648 5358 1706 5363
rect 1648 5357 1683 5358
rect 885 5320 922 5349
rect 886 5318 922 5320
rect 1098 5318 1135 5349
rect 886 5296 1135 5318
rect 967 5290 1078 5296
rect 967 5282 1008 5290
rect 967 5262 975 5282
rect 994 5262 1008 5282
rect 967 5260 1008 5262
rect 1036 5282 1078 5290
rect 1036 5262 1052 5282
rect 1071 5262 1078 5282
rect 1036 5260 1078 5262
rect 967 5245 1078 5260
rect 1306 5250 1343 5349
rect 1619 5345 1683 5357
rect 969 5236 1073 5245
rect 757 5205 878 5215
rect 757 5203 826 5205
rect 757 5162 770 5203
rect 807 5164 826 5203
rect 863 5164 878 5205
rect 807 5162 878 5164
rect 757 5144 878 5162
rect 550 5100 611 5112
rect 1304 5100 1345 5250
rect 1723 5242 1750 5497
rect 1812 5487 1892 5498
rect 1812 5461 1829 5487
rect 1869 5461 1892 5487
rect 1812 5434 1892 5461
rect 1812 5408 1833 5434
rect 1873 5408 1892 5434
rect 1812 5389 1892 5408
rect 1812 5363 1836 5389
rect 1876 5363 1892 5389
rect 1812 5312 1892 5363
rect 550 5097 1345 5100
rect 1724 5111 1750 5242
rect 1814 5156 1884 5312
rect 1813 5140 1889 5156
rect 1724 5097 1752 5111
rect 550 5062 1752 5097
rect 1813 5103 1828 5140
rect 1872 5103 1889 5140
rect 1813 5083 1889 5103
rect 2927 5133 2997 6042
rect 3096 5521 3177 6190
rect 4001 6085 4037 6385
rect 3925 6056 4038 6085
rect 3925 5691 3956 6056
rect 3849 5671 4242 5691
rect 4262 5671 4265 5691
rect 3849 5666 4265 5671
rect 3849 5665 4190 5666
rect 3506 5634 3616 5648
rect 3506 5631 3549 5634
rect 3506 5626 3510 5631
rect 3428 5604 3510 5626
rect 3539 5604 3549 5631
rect 3577 5607 3584 5634
rect 3613 5626 3616 5634
rect 3613 5607 3678 5626
rect 3577 5604 3678 5607
rect 3428 5602 3678 5604
rect 3428 5523 3465 5602
rect 3506 5589 3616 5602
rect 3580 5533 3611 5534
rect 3090 5441 3189 5521
rect 3428 5503 3437 5523
rect 3457 5503 3465 5523
rect 3428 5493 3465 5503
rect 3524 5523 3611 5533
rect 3524 5503 3533 5523
rect 3553 5503 3611 5523
rect 3524 5494 3611 5503
rect 3524 5493 3561 5494
rect 3580 5441 3611 5494
rect 3641 5523 3678 5602
rect 3793 5533 3824 5534
rect 3641 5503 3650 5523
rect 3670 5503 3678 5523
rect 3641 5493 3678 5503
rect 3737 5526 3824 5533
rect 3737 5523 3798 5526
rect 3737 5503 3746 5523
rect 3766 5506 3798 5523
rect 3819 5506 3824 5526
rect 3766 5503 3824 5506
rect 3737 5496 3824 5503
rect 3849 5523 3886 5665
rect 4152 5664 4189 5665
rect 4001 5533 4037 5534
rect 3849 5503 3858 5523
rect 3878 5503 3886 5523
rect 3737 5494 3793 5496
rect 3737 5493 3774 5494
rect 3849 5493 3886 5503
rect 3945 5523 4093 5533
rect 4193 5530 4289 5532
rect 3945 5503 3954 5523
rect 3974 5503 4064 5523
rect 4084 5503 4093 5523
rect 3945 5497 4093 5503
rect 3945 5494 4009 5497
rect 3945 5493 3982 5494
rect 4001 5467 4009 5494
rect 4030 5494 4093 5497
rect 4151 5523 4289 5530
rect 4151 5503 4160 5523
rect 4180 5503 4289 5523
rect 4151 5494 4289 5503
rect 4030 5467 4037 5494
rect 4056 5493 4093 5494
rect 4152 5493 4189 5494
rect 4001 5442 4037 5467
rect 3090 5440 3430 5441
rect 3472 5440 3513 5441
rect 3090 5433 3513 5440
rect 3090 5413 3482 5433
rect 3502 5413 3513 5433
rect 3090 5405 3513 5413
rect 3580 5437 3939 5441
rect 3580 5432 3902 5437
rect 3580 5408 3693 5432
rect 3717 5413 3902 5432
rect 3926 5413 3939 5437
rect 3717 5408 3939 5413
rect 3580 5405 3939 5408
rect 4001 5405 4036 5442
rect 4104 5439 4204 5442
rect 4104 5435 4171 5439
rect 4104 5409 4116 5435
rect 4142 5413 4171 5435
rect 4197 5413 4204 5439
rect 4142 5409 4204 5413
rect 4104 5405 4204 5409
rect 3090 5401 3430 5405
rect 2927 5083 2999 5133
rect 550 4987 611 5062
rect 969 5060 1073 5062
rect 1304 5060 1345 5062
rect 1813 5017 1823 5083
rect 1877 5017 1889 5083
rect 1813 4993 1889 5017
rect 552 4857 611 4987
rect 1465 4938 1537 4939
rect 1464 4930 1563 4938
rect 1464 4927 1516 4930
rect 1464 4892 1472 4927
rect 1497 4892 1516 4927
rect 1541 4919 1563 4930
rect 1541 4918 2408 4919
rect 1541 4892 2409 4918
rect 1464 4882 2409 4892
rect 1464 4880 1563 4882
rect 552 4839 574 4857
rect 592 4839 611 4857
rect 552 4817 611 4839
rect 819 4853 1351 4858
rect 819 4833 1705 4853
rect 1725 4833 1728 4853
rect 2364 4849 2409 4882
rect 819 4829 1728 4833
rect 819 4782 862 4829
rect 1312 4828 1728 4829
rect 2360 4829 2753 4849
rect 2773 4829 2776 4849
rect 1312 4827 1653 4828
rect 969 4796 1079 4810
rect 969 4793 1012 4796
rect 969 4788 973 4793
rect 807 4781 862 4782
rect 551 4758 862 4781
rect 551 4740 576 4758
rect 594 4746 862 4758
rect 891 4766 973 4788
rect 1002 4766 1012 4793
rect 1040 4769 1047 4796
rect 1076 4788 1079 4796
rect 1076 4769 1141 4788
rect 1040 4766 1141 4769
rect 891 4764 1141 4766
rect 594 4740 616 4746
rect 551 4601 616 4740
rect 891 4685 928 4764
rect 969 4751 1079 4764
rect 1043 4695 1074 4696
rect 891 4665 900 4685
rect 920 4665 928 4685
rect 551 4583 574 4601
rect 592 4583 616 4601
rect 551 4566 616 4583
rect 771 4647 839 4660
rect 891 4655 928 4665
rect 987 4685 1074 4695
rect 987 4665 996 4685
rect 1016 4665 1074 4685
rect 987 4656 1074 4665
rect 987 4655 1024 4656
rect 771 4605 778 4647
rect 827 4605 839 4647
rect 771 4602 839 4605
rect 1043 4603 1074 4656
rect 1104 4685 1141 4764
rect 1256 4695 1287 4696
rect 1104 4665 1113 4685
rect 1133 4665 1141 4685
rect 1104 4655 1141 4665
rect 1200 4688 1287 4695
rect 1200 4685 1261 4688
rect 1200 4665 1209 4685
rect 1229 4668 1261 4685
rect 1282 4668 1287 4688
rect 1229 4665 1287 4668
rect 1200 4658 1287 4665
rect 1312 4685 1349 4827
rect 1615 4826 1652 4827
rect 2360 4824 2776 4829
rect 2360 4823 2701 4824
rect 2017 4792 2127 4806
rect 2017 4789 2060 4792
rect 2017 4784 2021 4789
rect 1939 4762 2021 4784
rect 2050 4762 2060 4789
rect 2088 4765 2095 4792
rect 2124 4784 2127 4792
rect 2124 4765 2189 4784
rect 2088 4762 2189 4765
rect 1939 4760 2189 4762
rect 1464 4695 1500 4696
rect 1312 4665 1321 4685
rect 1341 4665 1349 4685
rect 1200 4656 1256 4658
rect 1200 4655 1237 4656
rect 1312 4655 1349 4665
rect 1408 4685 1556 4695
rect 1656 4692 1752 4694
rect 1408 4665 1417 4685
rect 1437 4665 1527 4685
rect 1547 4665 1556 4685
rect 1408 4659 1556 4665
rect 1408 4656 1472 4659
rect 1408 4655 1445 4656
rect 1464 4629 1472 4656
rect 1493 4656 1556 4659
rect 1614 4685 1752 4692
rect 1614 4665 1623 4685
rect 1643 4665 1752 4685
rect 1614 4656 1752 4665
rect 1939 4681 1976 4760
rect 2017 4747 2127 4760
rect 2091 4691 2122 4692
rect 1939 4661 1948 4681
rect 1968 4661 1976 4681
rect 1493 4629 1500 4656
rect 1519 4655 1556 4656
rect 1615 4655 1652 4656
rect 1464 4604 1500 4629
rect 935 4602 976 4603
rect 771 4595 976 4602
rect 771 4584 945 4595
rect 771 4551 779 4584
rect 772 4542 779 4551
rect 828 4575 945 4584
rect 965 4575 976 4595
rect 828 4567 976 4575
rect 1043 4599 1402 4603
rect 1043 4594 1365 4599
rect 1043 4570 1156 4594
rect 1180 4575 1365 4594
rect 1389 4575 1402 4599
rect 1180 4570 1402 4575
rect 1043 4567 1402 4570
rect 1464 4567 1499 4604
rect 1567 4601 1667 4604
rect 1567 4597 1634 4601
rect 1567 4571 1579 4597
rect 1605 4575 1634 4597
rect 1660 4575 1667 4601
rect 1605 4571 1667 4575
rect 1567 4567 1667 4571
rect 828 4551 839 4567
rect 828 4542 836 4551
rect 1043 4546 1074 4567
rect 1464 4546 1500 4567
rect 886 4545 923 4546
rect 551 4502 616 4521
rect 551 4484 576 4502
rect 594 4484 616 4502
rect 551 4283 616 4484
rect 772 4358 836 4542
rect 885 4536 923 4545
rect 885 4516 894 4536
rect 914 4516 923 4536
rect 885 4508 923 4516
rect 989 4540 1074 4546
rect 1099 4545 1136 4546
rect 989 4520 997 4540
rect 1017 4520 1074 4540
rect 989 4512 1074 4520
rect 1098 4536 1136 4545
rect 1098 4516 1107 4536
rect 1127 4516 1136 4536
rect 989 4511 1025 4512
rect 1098 4508 1136 4516
rect 1202 4540 1287 4546
rect 1307 4545 1344 4546
rect 1202 4520 1210 4540
rect 1230 4539 1287 4540
rect 1230 4520 1259 4539
rect 1202 4519 1259 4520
rect 1280 4519 1287 4539
rect 1202 4512 1287 4519
rect 1306 4536 1344 4545
rect 1306 4516 1315 4536
rect 1335 4516 1344 4536
rect 1202 4511 1238 4512
rect 1306 4508 1344 4516
rect 1410 4540 1554 4546
rect 1410 4520 1418 4540
rect 1438 4520 1526 4540
rect 1546 4520 1554 4540
rect 1410 4512 1554 4520
rect 1410 4511 1446 4512
rect 1518 4511 1554 4512
rect 1620 4545 1657 4546
rect 1620 4544 1658 4545
rect 1620 4536 1684 4544
rect 1620 4516 1629 4536
rect 1649 4522 1684 4536
rect 1704 4522 1707 4542
rect 1649 4517 1707 4522
rect 1649 4516 1684 4517
rect 886 4479 923 4508
rect 887 4477 923 4479
rect 1099 4477 1136 4508
rect 887 4455 1136 4477
rect 968 4449 1079 4455
rect 968 4441 1009 4449
rect 968 4421 976 4441
rect 995 4421 1009 4441
rect 968 4419 1009 4421
rect 1037 4441 1079 4449
rect 1037 4421 1053 4441
rect 1072 4421 1079 4441
rect 1037 4419 1079 4421
rect 968 4404 1079 4419
rect 772 4348 840 4358
rect 772 4315 789 4348
rect 829 4315 840 4348
rect 772 4303 840 4315
rect 772 4301 836 4303
rect 1307 4284 1344 4508
rect 1620 4504 1684 4516
rect 1724 4286 1751 4656
rect 1939 4651 1976 4661
rect 2035 4681 2122 4691
rect 2035 4661 2044 4681
rect 2064 4661 2122 4681
rect 2035 4652 2122 4661
rect 2035 4651 2072 4652
rect 1815 4638 1885 4643
rect 1810 4632 1885 4638
rect 1810 4599 1818 4632
rect 1871 4599 1885 4632
rect 2091 4599 2122 4652
rect 2152 4681 2189 4760
rect 2304 4691 2335 4692
rect 2152 4661 2161 4681
rect 2181 4661 2189 4681
rect 2152 4651 2189 4661
rect 2248 4684 2335 4691
rect 2248 4681 2309 4684
rect 2248 4661 2257 4681
rect 2277 4664 2309 4681
rect 2330 4664 2335 4684
rect 2277 4661 2335 4664
rect 2248 4654 2335 4661
rect 2360 4681 2397 4823
rect 2663 4822 2700 4823
rect 2512 4691 2548 4692
rect 2360 4661 2369 4681
rect 2389 4661 2397 4681
rect 2248 4652 2304 4654
rect 2248 4651 2285 4652
rect 2360 4651 2397 4661
rect 2456 4681 2604 4691
rect 2704 4688 2800 4690
rect 2456 4661 2465 4681
rect 2485 4661 2575 4681
rect 2595 4661 2604 4681
rect 2456 4655 2604 4661
rect 2456 4652 2520 4655
rect 2456 4651 2493 4652
rect 2512 4625 2520 4652
rect 2541 4652 2604 4655
rect 2662 4681 2800 4688
rect 2662 4661 2671 4681
rect 2691 4661 2800 4681
rect 2662 4652 2800 4661
rect 2541 4625 2548 4652
rect 2567 4651 2604 4652
rect 2663 4651 2700 4652
rect 2512 4600 2548 4625
rect 1810 4598 1893 4599
rect 1983 4598 2024 4599
rect 1810 4591 2024 4598
rect 1810 4574 1993 4591
rect 1810 4541 1823 4574
rect 1876 4571 1993 4574
rect 2013 4571 2024 4591
rect 1876 4563 2024 4571
rect 2091 4595 2450 4599
rect 2091 4590 2413 4595
rect 2091 4566 2204 4590
rect 2228 4571 2413 4590
rect 2437 4571 2450 4595
rect 2228 4566 2450 4571
rect 2091 4563 2450 4566
rect 2512 4563 2547 4600
rect 2615 4597 2715 4600
rect 2615 4593 2682 4597
rect 2615 4567 2627 4593
rect 2653 4571 2682 4593
rect 2708 4571 2715 4597
rect 2653 4567 2715 4571
rect 2615 4563 2715 4567
rect 1876 4541 1893 4563
rect 2091 4542 2122 4563
rect 2512 4542 2548 4563
rect 1934 4541 1971 4542
rect 1810 4527 1893 4541
rect 1583 4284 1751 4286
rect 1307 4283 1751 4284
rect 551 4253 1751 4283
rect 1821 4317 1893 4527
rect 1933 4532 1971 4541
rect 1933 4512 1942 4532
rect 1962 4512 1971 4532
rect 1933 4504 1971 4512
rect 2037 4536 2122 4542
rect 2147 4541 2184 4542
rect 2037 4516 2045 4536
rect 2065 4516 2122 4536
rect 2037 4508 2122 4516
rect 2146 4532 2184 4541
rect 2146 4512 2155 4532
rect 2175 4512 2184 4532
rect 2037 4507 2073 4508
rect 2146 4504 2184 4512
rect 2250 4536 2335 4542
rect 2355 4541 2392 4542
rect 2250 4516 2258 4536
rect 2278 4535 2335 4536
rect 2278 4516 2307 4535
rect 2250 4515 2307 4516
rect 2328 4515 2335 4535
rect 2250 4508 2335 4515
rect 2354 4532 2392 4541
rect 2354 4512 2363 4532
rect 2383 4512 2392 4532
rect 2250 4507 2286 4508
rect 2354 4504 2392 4512
rect 2458 4536 2602 4542
rect 2458 4516 2466 4536
rect 2486 4516 2574 4536
rect 2594 4516 2602 4536
rect 2458 4508 2602 4516
rect 2458 4507 2494 4508
rect 2566 4507 2602 4508
rect 2668 4541 2705 4542
rect 2668 4540 2706 4541
rect 2668 4532 2732 4540
rect 2668 4512 2677 4532
rect 2697 4518 2732 4532
rect 2752 4518 2755 4538
rect 2697 4513 2755 4518
rect 2697 4512 2732 4513
rect 1934 4475 1971 4504
rect 1935 4473 1971 4475
rect 2147 4473 2184 4504
rect 1935 4451 2184 4473
rect 2016 4445 2127 4451
rect 2016 4437 2057 4445
rect 2016 4417 2024 4437
rect 2043 4417 2057 4437
rect 2016 4415 2057 4417
rect 2085 4437 2127 4445
rect 2085 4417 2101 4437
rect 2120 4417 2127 4437
rect 2085 4415 2127 4417
rect 2016 4400 2127 4415
rect 1821 4278 1840 4317
rect 1885 4278 1893 4317
rect 1821 4261 1893 4278
rect 2355 4305 2392 4504
rect 2668 4500 2732 4512
rect 2355 4299 2396 4305
rect 2772 4301 2799 4652
rect 2928 4604 2999 5083
rect 2928 4520 2997 4604
rect 2631 4299 2799 4301
rect 2355 4273 2799 4299
rect 551 4206 616 4253
rect 551 4188 574 4206
rect 592 4188 616 4206
rect 1464 4233 1499 4235
rect 1464 4231 1568 4233
rect 2357 4231 2396 4273
rect 2631 4272 2799 4273
rect 1464 4224 2398 4231
rect 1464 4223 1515 4224
rect 1464 4203 1467 4223
rect 1492 4204 1515 4223
rect 1547 4204 2398 4224
rect 1492 4203 2398 4204
rect 1464 4196 2398 4203
rect 1737 4195 2398 4196
rect 551 4167 616 4188
rect 828 4178 868 4181
rect 828 4174 1731 4178
rect 828 4154 1705 4174
rect 1725 4154 1731 4174
rect 828 4151 1731 4154
rect 552 4107 617 4127
rect 552 4089 576 4107
rect 594 4089 617 4107
rect 552 4062 617 4089
rect 828 4062 868 4151
rect 1312 4149 1728 4151
rect 1312 4148 1653 4149
rect 969 4117 1079 4131
rect 969 4114 1012 4117
rect 969 4109 973 4114
rect 551 4027 868 4062
rect 891 4087 973 4109
rect 1002 4087 1012 4114
rect 1040 4090 1047 4117
rect 1076 4109 1079 4117
rect 1076 4090 1141 4109
rect 1040 4087 1141 4090
rect 891 4085 1141 4087
rect 552 3951 617 4027
rect 891 4006 928 4085
rect 969 4072 1079 4085
rect 1043 4016 1074 4017
rect 891 3986 900 4006
rect 920 3986 928 4006
rect 891 3976 928 3986
rect 987 4006 1074 4016
rect 987 3986 996 4006
rect 1016 3986 1074 4006
rect 987 3977 1074 3986
rect 987 3976 1024 3977
rect 552 3933 574 3951
rect 592 3933 617 3951
rect 552 3912 617 3933
rect 765 3931 830 3940
rect 765 3894 775 3931
rect 815 3923 830 3931
rect 1043 3924 1074 3977
rect 1104 4006 1141 4085
rect 1256 4016 1287 4017
rect 1104 3986 1113 4006
rect 1133 3986 1141 4006
rect 1104 3976 1141 3986
rect 1200 4009 1287 4016
rect 1200 4006 1261 4009
rect 1200 3986 1209 4006
rect 1229 3989 1261 4006
rect 1282 3989 1287 4009
rect 1229 3986 1287 3989
rect 1200 3979 1287 3986
rect 1312 4006 1349 4148
rect 1615 4147 1652 4148
rect 1464 4016 1500 4017
rect 1312 3986 1321 4006
rect 1341 3986 1349 4006
rect 1200 3977 1256 3979
rect 1200 3976 1237 3977
rect 1312 3976 1349 3986
rect 1408 4006 1556 4016
rect 1656 4013 1752 4015
rect 1408 3986 1417 4006
rect 1437 3986 1527 4006
rect 1547 3986 1556 4006
rect 1408 3980 1556 3986
rect 1408 3977 1472 3980
rect 1408 3976 1445 3977
rect 1464 3950 1472 3977
rect 1493 3977 1556 3980
rect 1614 4006 1752 4013
rect 2932 4008 2994 4520
rect 1614 3986 1623 4006
rect 1643 3986 1752 4006
rect 1614 3977 1752 3986
rect 1493 3950 1500 3977
rect 1519 3976 1556 3977
rect 1615 3976 1652 3977
rect 1464 3925 1500 3950
rect 935 3923 976 3924
rect 815 3916 976 3923
rect 815 3896 945 3916
rect 965 3896 976 3916
rect 815 3894 976 3896
rect 765 3888 976 3894
rect 1043 3920 1402 3924
rect 1043 3915 1365 3920
rect 1043 3891 1156 3915
rect 1180 3896 1365 3915
rect 1389 3896 1402 3920
rect 1180 3891 1402 3896
rect 1043 3888 1402 3891
rect 1464 3888 1499 3925
rect 1567 3922 1667 3925
rect 1567 3918 1634 3922
rect 1567 3892 1579 3918
rect 1605 3896 1634 3918
rect 1660 3896 1667 3922
rect 1605 3892 1667 3896
rect 1567 3888 1667 3892
rect 765 3875 832 3888
rect 557 3852 613 3872
rect 557 3834 576 3852
rect 594 3834 613 3852
rect 557 3721 613 3834
rect 765 3854 779 3875
rect 815 3854 832 3875
rect 1043 3867 1074 3888
rect 1464 3867 1500 3888
rect 886 3866 923 3867
rect 765 3847 832 3854
rect 885 3857 923 3866
rect 557 3583 612 3721
rect 765 3695 830 3847
rect 885 3837 894 3857
rect 914 3837 923 3857
rect 885 3829 923 3837
rect 989 3861 1074 3867
rect 1099 3866 1136 3867
rect 989 3841 997 3861
rect 1017 3841 1074 3861
rect 989 3833 1074 3841
rect 1098 3857 1136 3866
rect 1098 3837 1107 3857
rect 1127 3837 1136 3857
rect 989 3832 1025 3833
rect 1098 3829 1136 3837
rect 1202 3861 1287 3867
rect 1307 3866 1344 3867
rect 1202 3841 1210 3861
rect 1230 3860 1287 3861
rect 1230 3841 1259 3860
rect 1202 3840 1259 3841
rect 1280 3840 1287 3860
rect 1202 3833 1287 3840
rect 1306 3857 1344 3866
rect 1306 3837 1315 3857
rect 1335 3837 1344 3857
rect 1202 3832 1238 3833
rect 1306 3829 1344 3837
rect 1410 3861 1554 3867
rect 1410 3841 1418 3861
rect 1438 3841 1526 3861
rect 1546 3841 1554 3861
rect 1410 3833 1554 3841
rect 1410 3832 1446 3833
rect 1518 3832 1554 3833
rect 1620 3866 1657 3867
rect 1620 3865 1658 3866
rect 1620 3857 1684 3865
rect 1620 3837 1629 3857
rect 1649 3843 1684 3857
rect 1704 3843 1707 3863
rect 1649 3838 1707 3843
rect 1649 3837 1684 3838
rect 886 3800 923 3829
rect 887 3798 923 3800
rect 1099 3798 1136 3829
rect 887 3776 1136 3798
rect 968 3770 1079 3776
rect 968 3762 1009 3770
rect 968 3742 976 3762
rect 995 3742 1009 3762
rect 968 3740 1009 3742
rect 1037 3762 1079 3770
rect 1037 3742 1053 3762
rect 1072 3742 1079 3762
rect 1037 3740 1079 3742
rect 968 3727 1079 3740
rect 1307 3730 1344 3829
rect 1620 3825 1684 3837
rect 758 3685 879 3695
rect 758 3683 827 3685
rect 758 3642 771 3683
rect 808 3644 827 3683
rect 864 3644 879 3685
rect 808 3642 879 3644
rect 758 3624 879 3642
rect 550 3580 614 3583
rect 970 3580 1074 3586
rect 1305 3580 1346 3730
rect 1724 3722 1751 3977
rect 1813 3967 1893 3978
rect 1813 3941 1830 3967
rect 1870 3941 1893 3967
rect 1813 3914 1893 3941
rect 2936 3969 2994 4008
rect 2936 3934 2998 3969
rect 1813 3888 1834 3914
rect 1874 3888 1893 3914
rect 1813 3869 1893 3888
rect 1813 3843 1837 3869
rect 1877 3843 1893 3869
rect 1813 3792 1893 3843
rect 2885 3907 2998 3934
rect 2885 3905 2944 3907
rect 2885 3874 2899 3905
rect 2924 3884 2944 3905
rect 2970 3884 2998 3907
rect 2924 3874 2998 3884
rect 2885 3864 2998 3874
rect 550 3577 1346 3580
rect 1725 3591 1751 3722
rect 1725 3577 1753 3591
rect 550 3542 1753 3577
rect 1815 3584 1885 3792
rect 550 3481 614 3542
rect 970 3540 1074 3542
rect 1305 3540 1346 3542
rect 1815 3539 1836 3584
rect 1816 3518 1836 3539
rect 1866 3539 1885 3584
rect 1866 3518 1883 3539
rect 1816 3499 1883 3518
rect 1465 3491 1537 3492
rect 1464 3483 1563 3491
rect 552 3410 611 3481
rect 1464 3480 1516 3483
rect 1464 3445 1472 3480
rect 1497 3445 1516 3480
rect 1541 3472 1563 3483
rect 1541 3471 2408 3472
rect 1541 3445 2409 3471
rect 1464 3435 2409 3445
rect 1464 3433 1563 3435
rect 552 3392 574 3410
rect 592 3392 611 3410
rect 552 3370 611 3392
rect 819 3406 1351 3411
rect 819 3386 1705 3406
rect 1725 3386 1728 3406
rect 2364 3402 2409 3435
rect 819 3382 1728 3386
rect 819 3335 862 3382
rect 1312 3381 1728 3382
rect 2360 3382 2753 3402
rect 2773 3382 2776 3402
rect 1312 3380 1653 3381
rect 969 3349 1079 3363
rect 969 3346 1012 3349
rect 969 3341 973 3346
rect 807 3334 862 3335
rect 551 3311 862 3334
rect 551 3293 576 3311
rect 594 3299 862 3311
rect 891 3319 973 3341
rect 1002 3319 1012 3346
rect 1040 3322 1047 3349
rect 1076 3341 1079 3349
rect 1076 3322 1141 3341
rect 1040 3319 1141 3322
rect 891 3317 1141 3319
rect 594 3293 616 3299
rect 551 3154 616 3293
rect 891 3238 928 3317
rect 969 3304 1079 3317
rect 1043 3248 1074 3249
rect 891 3218 900 3238
rect 920 3218 928 3238
rect 551 3136 574 3154
rect 592 3136 616 3154
rect 551 3119 616 3136
rect 771 3200 839 3213
rect 891 3208 928 3218
rect 987 3238 1074 3248
rect 987 3218 996 3238
rect 1016 3218 1074 3238
rect 987 3209 1074 3218
rect 987 3208 1024 3209
rect 771 3158 778 3200
rect 827 3158 839 3200
rect 771 3155 839 3158
rect 1043 3156 1074 3209
rect 1104 3238 1141 3317
rect 1256 3248 1287 3249
rect 1104 3218 1113 3238
rect 1133 3218 1141 3238
rect 1104 3208 1141 3218
rect 1200 3241 1287 3248
rect 1200 3238 1261 3241
rect 1200 3218 1209 3238
rect 1229 3221 1261 3238
rect 1282 3221 1287 3241
rect 1229 3218 1287 3221
rect 1200 3211 1287 3218
rect 1312 3238 1349 3380
rect 1615 3379 1652 3380
rect 2360 3377 2776 3382
rect 2360 3376 2701 3377
rect 2017 3345 2127 3359
rect 2017 3342 2060 3345
rect 2017 3337 2021 3342
rect 1939 3315 2021 3337
rect 2050 3315 2060 3342
rect 2088 3318 2095 3345
rect 2124 3337 2127 3345
rect 2124 3318 2189 3337
rect 2088 3315 2189 3318
rect 1939 3313 2189 3315
rect 1464 3248 1500 3249
rect 1312 3218 1321 3238
rect 1341 3218 1349 3238
rect 1200 3209 1256 3211
rect 1200 3208 1237 3209
rect 1312 3208 1349 3218
rect 1408 3238 1556 3248
rect 1656 3245 1752 3247
rect 1408 3218 1417 3238
rect 1437 3218 1527 3238
rect 1547 3218 1556 3238
rect 1408 3212 1556 3218
rect 1408 3209 1472 3212
rect 1408 3208 1445 3209
rect 1464 3182 1472 3209
rect 1493 3209 1556 3212
rect 1614 3238 1752 3245
rect 1614 3218 1623 3238
rect 1643 3218 1752 3238
rect 1614 3209 1752 3218
rect 1939 3234 1976 3313
rect 2017 3300 2127 3313
rect 2091 3244 2122 3245
rect 1939 3214 1948 3234
rect 1968 3214 1976 3234
rect 1493 3182 1500 3209
rect 1519 3208 1556 3209
rect 1615 3208 1652 3209
rect 1464 3157 1500 3182
rect 935 3155 976 3156
rect 771 3148 976 3155
rect 771 3137 945 3148
rect 771 3104 779 3137
rect 772 3095 779 3104
rect 828 3128 945 3137
rect 965 3128 976 3148
rect 828 3120 976 3128
rect 1043 3152 1402 3156
rect 1043 3147 1365 3152
rect 1043 3123 1156 3147
rect 1180 3128 1365 3147
rect 1389 3128 1402 3152
rect 1180 3123 1402 3128
rect 1043 3120 1402 3123
rect 1464 3120 1499 3157
rect 1567 3154 1667 3157
rect 1567 3150 1634 3154
rect 1567 3124 1579 3150
rect 1605 3128 1634 3150
rect 1660 3128 1667 3154
rect 1605 3124 1667 3128
rect 1567 3120 1667 3124
rect 828 3104 839 3120
rect 828 3095 836 3104
rect 1043 3099 1074 3120
rect 1464 3099 1500 3120
rect 886 3098 923 3099
rect 551 3055 616 3074
rect 551 3037 576 3055
rect 594 3037 616 3055
rect 551 2836 616 3037
rect 772 2911 836 3095
rect 885 3089 923 3098
rect 885 3069 894 3089
rect 914 3069 923 3089
rect 885 3061 923 3069
rect 989 3093 1074 3099
rect 1099 3098 1136 3099
rect 989 3073 997 3093
rect 1017 3073 1074 3093
rect 989 3065 1074 3073
rect 1098 3089 1136 3098
rect 1098 3069 1107 3089
rect 1127 3069 1136 3089
rect 989 3064 1025 3065
rect 1098 3061 1136 3069
rect 1202 3093 1287 3099
rect 1307 3098 1344 3099
rect 1202 3073 1210 3093
rect 1230 3092 1287 3093
rect 1230 3073 1259 3092
rect 1202 3072 1259 3073
rect 1280 3072 1287 3092
rect 1202 3065 1287 3072
rect 1306 3089 1344 3098
rect 1306 3069 1315 3089
rect 1335 3069 1344 3089
rect 1202 3064 1238 3065
rect 1306 3061 1344 3069
rect 1410 3093 1554 3099
rect 1410 3073 1418 3093
rect 1438 3073 1526 3093
rect 1546 3073 1554 3093
rect 1410 3065 1554 3073
rect 1410 3064 1446 3065
rect 1518 3064 1554 3065
rect 1620 3098 1657 3099
rect 1620 3097 1658 3098
rect 1620 3089 1684 3097
rect 1620 3069 1629 3089
rect 1649 3075 1684 3089
rect 1704 3075 1707 3095
rect 1649 3070 1707 3075
rect 1649 3069 1684 3070
rect 886 3032 923 3061
rect 887 3030 923 3032
rect 1099 3030 1136 3061
rect 887 3008 1136 3030
rect 968 3002 1079 3008
rect 968 2994 1009 3002
rect 968 2974 976 2994
rect 995 2974 1009 2994
rect 968 2972 1009 2974
rect 1037 2994 1079 3002
rect 1037 2974 1053 2994
rect 1072 2974 1079 2994
rect 1037 2972 1079 2974
rect 968 2957 1079 2972
rect 772 2901 840 2911
rect 772 2868 789 2901
rect 829 2868 840 2901
rect 772 2856 840 2868
rect 772 2854 836 2856
rect 1307 2837 1344 3061
rect 1620 3057 1684 3069
rect 1724 2839 1751 3209
rect 1939 3204 1976 3214
rect 2035 3234 2122 3244
rect 2035 3214 2044 3234
rect 2064 3214 2122 3234
rect 2035 3205 2122 3214
rect 2035 3204 2072 3205
rect 1815 3191 1885 3196
rect 1810 3185 1885 3191
rect 1810 3152 1818 3185
rect 1871 3152 1885 3185
rect 2091 3152 2122 3205
rect 2152 3234 2189 3313
rect 2304 3244 2335 3245
rect 2152 3214 2161 3234
rect 2181 3214 2189 3234
rect 2152 3204 2189 3214
rect 2248 3237 2335 3244
rect 2248 3234 2309 3237
rect 2248 3214 2257 3234
rect 2277 3217 2309 3234
rect 2330 3217 2335 3237
rect 2277 3214 2335 3217
rect 2248 3207 2335 3214
rect 2360 3234 2397 3376
rect 2663 3375 2700 3376
rect 2512 3244 2548 3245
rect 2360 3214 2369 3234
rect 2389 3214 2397 3234
rect 2248 3205 2304 3207
rect 2248 3204 2285 3205
rect 2360 3204 2397 3214
rect 2456 3234 2604 3244
rect 2704 3241 2800 3243
rect 2456 3214 2465 3234
rect 2485 3214 2575 3234
rect 2595 3214 2604 3234
rect 2456 3208 2604 3214
rect 2456 3205 2520 3208
rect 2456 3204 2493 3205
rect 2512 3178 2520 3205
rect 2541 3205 2604 3208
rect 2662 3234 2800 3241
rect 2662 3214 2671 3234
rect 2691 3214 2800 3234
rect 2662 3205 2800 3214
rect 2541 3178 2548 3205
rect 2567 3204 2604 3205
rect 2663 3204 2700 3205
rect 2512 3153 2548 3178
rect 1810 3151 1893 3152
rect 1983 3151 2024 3152
rect 1810 3144 2024 3151
rect 1810 3127 1993 3144
rect 1810 3094 1823 3127
rect 1876 3124 1993 3127
rect 2013 3124 2024 3144
rect 1876 3116 2024 3124
rect 2091 3148 2450 3152
rect 2091 3143 2413 3148
rect 2091 3119 2204 3143
rect 2228 3124 2413 3143
rect 2437 3124 2450 3148
rect 2228 3119 2450 3124
rect 2091 3116 2450 3119
rect 2512 3116 2547 3153
rect 2615 3150 2715 3153
rect 2615 3146 2682 3150
rect 2615 3120 2627 3146
rect 2653 3124 2682 3146
rect 2708 3124 2715 3150
rect 2653 3120 2715 3124
rect 2615 3116 2715 3120
rect 1876 3094 1893 3116
rect 2091 3095 2122 3116
rect 2512 3095 2548 3116
rect 1934 3094 1971 3095
rect 1810 3080 1893 3094
rect 1583 2837 1751 2839
rect 1307 2836 1751 2837
rect 551 2806 1751 2836
rect 1821 2870 1893 3080
rect 1933 3085 1971 3094
rect 1933 3065 1942 3085
rect 1962 3065 1971 3085
rect 1933 3057 1971 3065
rect 2037 3089 2122 3095
rect 2147 3094 2184 3095
rect 2037 3069 2045 3089
rect 2065 3069 2122 3089
rect 2037 3061 2122 3069
rect 2146 3085 2184 3094
rect 2146 3065 2155 3085
rect 2175 3065 2184 3085
rect 2037 3060 2073 3061
rect 2146 3057 2184 3065
rect 2250 3089 2335 3095
rect 2355 3094 2392 3095
rect 2250 3069 2258 3089
rect 2278 3088 2335 3089
rect 2278 3069 2307 3088
rect 2250 3068 2307 3069
rect 2328 3068 2335 3088
rect 2250 3061 2335 3068
rect 2354 3085 2392 3094
rect 2354 3065 2363 3085
rect 2383 3065 2392 3085
rect 2250 3060 2286 3061
rect 2354 3057 2392 3065
rect 2458 3089 2602 3095
rect 2458 3069 2466 3089
rect 2486 3069 2574 3089
rect 2594 3069 2602 3089
rect 2458 3061 2602 3069
rect 2458 3060 2494 3061
rect 2566 3060 2602 3061
rect 2668 3094 2705 3095
rect 2668 3093 2706 3094
rect 2668 3085 2732 3093
rect 2668 3065 2677 3085
rect 2697 3071 2732 3085
rect 2752 3071 2755 3091
rect 2697 3066 2755 3071
rect 2697 3065 2732 3066
rect 1934 3028 1971 3057
rect 1935 3026 1971 3028
rect 2147 3026 2184 3057
rect 1935 3004 2184 3026
rect 2016 2998 2127 3004
rect 2016 2990 2057 2998
rect 2016 2970 2024 2990
rect 2043 2970 2057 2990
rect 2016 2968 2057 2970
rect 2085 2990 2127 2998
rect 2085 2970 2101 2990
rect 2120 2970 2127 2990
rect 2085 2968 2127 2970
rect 2016 2953 2127 2968
rect 1821 2831 1840 2870
rect 1885 2831 1893 2870
rect 1821 2814 1893 2831
rect 2355 2858 2392 3057
rect 2668 3053 2732 3065
rect 2355 2852 2396 2858
rect 2772 2854 2799 3205
rect 2631 2852 2799 2854
rect 2355 2826 2799 2852
rect 551 2759 616 2806
rect 551 2741 574 2759
rect 592 2741 616 2759
rect 1464 2786 1499 2788
rect 1464 2784 1568 2786
rect 2357 2784 2396 2826
rect 2631 2825 2799 2826
rect 1464 2777 2398 2784
rect 1464 2776 1515 2777
rect 1464 2756 1467 2776
rect 1492 2757 1515 2776
rect 1547 2757 2398 2777
rect 1492 2756 2398 2757
rect 1464 2749 2398 2756
rect 1737 2748 2398 2749
rect 551 2720 616 2741
rect 828 2731 868 2734
rect 828 2727 1731 2731
rect 828 2707 1705 2727
rect 1725 2707 1731 2727
rect 828 2704 1731 2707
rect 552 2660 617 2680
rect 552 2642 576 2660
rect 594 2642 617 2660
rect 552 2615 617 2642
rect 828 2615 868 2704
rect 1312 2702 1728 2704
rect 1312 2701 1653 2702
rect 969 2670 1079 2684
rect 969 2667 1012 2670
rect 969 2662 973 2667
rect 551 2580 868 2615
rect 891 2640 973 2662
rect 1002 2640 1012 2667
rect 1040 2643 1047 2670
rect 1076 2662 1079 2670
rect 1076 2643 1141 2662
rect 1040 2640 1141 2643
rect 891 2638 1141 2640
rect 552 2504 617 2580
rect 891 2559 928 2638
rect 969 2625 1079 2638
rect 1043 2569 1074 2570
rect 891 2539 900 2559
rect 920 2539 928 2559
rect 891 2529 928 2539
rect 987 2559 1074 2569
rect 987 2539 996 2559
rect 1016 2539 1074 2559
rect 987 2530 1074 2539
rect 987 2529 1024 2530
rect 552 2486 574 2504
rect 592 2486 617 2504
rect 552 2465 617 2486
rect 765 2484 830 2493
rect 765 2447 775 2484
rect 815 2476 830 2484
rect 1043 2477 1074 2530
rect 1104 2559 1141 2638
rect 1256 2569 1287 2570
rect 1104 2539 1113 2559
rect 1133 2539 1141 2559
rect 1104 2529 1141 2539
rect 1200 2562 1287 2569
rect 1200 2559 1261 2562
rect 1200 2539 1209 2559
rect 1229 2542 1261 2559
rect 1282 2542 1287 2562
rect 1229 2539 1287 2542
rect 1200 2532 1287 2539
rect 1312 2559 1349 2701
rect 1615 2700 1652 2701
rect 1464 2569 1500 2570
rect 1312 2539 1321 2559
rect 1341 2539 1349 2559
rect 1200 2530 1256 2532
rect 1200 2529 1237 2530
rect 1312 2529 1349 2539
rect 1408 2559 1556 2569
rect 1656 2566 1752 2568
rect 1408 2539 1417 2559
rect 1437 2539 1527 2559
rect 1547 2539 1556 2559
rect 1408 2533 1556 2539
rect 1408 2530 1472 2533
rect 1408 2529 1445 2530
rect 1464 2503 1472 2530
rect 1493 2530 1556 2533
rect 1614 2559 1752 2566
rect 1614 2539 1623 2559
rect 1643 2539 1752 2559
rect 1614 2530 1752 2539
rect 1493 2503 1500 2530
rect 1519 2529 1556 2530
rect 1615 2529 1652 2530
rect 1464 2478 1500 2503
rect 935 2476 976 2477
rect 815 2469 976 2476
rect 815 2449 945 2469
rect 965 2449 976 2469
rect 815 2447 976 2449
rect 765 2441 976 2447
rect 1043 2473 1402 2477
rect 1043 2468 1365 2473
rect 1043 2444 1156 2468
rect 1180 2449 1365 2468
rect 1389 2449 1402 2473
rect 1180 2444 1402 2449
rect 1043 2441 1402 2444
rect 1464 2441 1499 2478
rect 1567 2475 1667 2478
rect 1567 2471 1634 2475
rect 1567 2445 1579 2471
rect 1605 2449 1634 2471
rect 1660 2449 1667 2475
rect 1605 2445 1667 2449
rect 1567 2441 1667 2445
rect 765 2428 832 2441
rect 557 2405 613 2425
rect 557 2387 576 2405
rect 594 2387 613 2405
rect 557 2352 613 2387
rect 519 2274 613 2352
rect 765 2407 779 2428
rect 815 2407 832 2428
rect 1043 2420 1074 2441
rect 1464 2420 1500 2441
rect 886 2419 923 2420
rect 765 2400 832 2407
rect 885 2410 923 2419
rect 519 2133 612 2274
rect 765 2248 830 2400
rect 885 2390 894 2410
rect 914 2390 923 2410
rect 885 2382 923 2390
rect 989 2414 1074 2420
rect 1099 2419 1136 2420
rect 989 2394 997 2414
rect 1017 2394 1074 2414
rect 989 2386 1074 2394
rect 1098 2410 1136 2419
rect 1098 2390 1107 2410
rect 1127 2390 1136 2410
rect 989 2385 1025 2386
rect 1098 2382 1136 2390
rect 1202 2414 1287 2420
rect 1307 2419 1344 2420
rect 1202 2394 1210 2414
rect 1230 2413 1287 2414
rect 1230 2394 1259 2413
rect 1202 2393 1259 2394
rect 1280 2393 1287 2413
rect 1202 2386 1287 2393
rect 1306 2410 1344 2419
rect 1306 2390 1315 2410
rect 1335 2390 1344 2410
rect 1202 2385 1238 2386
rect 1306 2382 1344 2390
rect 1410 2414 1554 2420
rect 1410 2394 1418 2414
rect 1438 2394 1526 2414
rect 1546 2394 1554 2414
rect 1410 2386 1554 2394
rect 1410 2385 1446 2386
rect 1518 2385 1554 2386
rect 1620 2419 1657 2420
rect 1620 2418 1658 2419
rect 1620 2410 1684 2418
rect 1620 2390 1629 2410
rect 1649 2396 1684 2410
rect 1704 2396 1707 2416
rect 1649 2391 1707 2396
rect 1649 2390 1684 2391
rect 886 2353 923 2382
rect 887 2351 923 2353
rect 1099 2351 1136 2382
rect 887 2329 1136 2351
rect 968 2323 1079 2329
rect 968 2315 1009 2323
rect 968 2295 976 2315
rect 995 2295 1009 2315
rect 968 2293 1009 2295
rect 1037 2315 1079 2323
rect 1037 2295 1053 2315
rect 1072 2295 1079 2315
rect 1037 2293 1079 2295
rect 968 2278 1079 2293
rect 1307 2283 1344 2382
rect 1620 2378 1684 2390
rect 1724 2339 1751 2530
rect 970 2269 1074 2278
rect 758 2238 879 2248
rect 758 2236 827 2238
rect 758 2195 771 2236
rect 808 2197 827 2236
rect 864 2197 879 2238
rect 808 2195 879 2197
rect 758 2177 879 2195
rect 970 2133 1074 2142
rect 1305 2133 1346 2283
rect 519 2131 1346 2133
rect 527 2130 1346 2131
rect 1725 2249 1750 2339
rect 2885 2307 2984 3864
rect 3090 2500 3189 5401
rect 3580 5384 3611 5405
rect 4001 5384 4037 5405
rect 3423 5383 3460 5384
rect 3422 5374 3460 5383
rect 3422 5354 3431 5374
rect 3451 5354 3460 5374
rect 3422 5346 3460 5354
rect 3526 5378 3611 5384
rect 3636 5383 3673 5384
rect 3526 5358 3534 5378
rect 3554 5358 3611 5378
rect 3526 5350 3611 5358
rect 3635 5374 3673 5383
rect 3635 5354 3644 5374
rect 3664 5354 3673 5374
rect 3526 5349 3562 5350
rect 3635 5346 3673 5354
rect 3739 5378 3824 5384
rect 3844 5383 3881 5384
rect 3739 5358 3747 5378
rect 3767 5377 3824 5378
rect 3767 5358 3796 5377
rect 3739 5357 3796 5358
rect 3817 5357 3824 5377
rect 3739 5350 3824 5357
rect 3843 5374 3881 5383
rect 3843 5354 3852 5374
rect 3872 5354 3881 5374
rect 3739 5349 3775 5350
rect 3843 5346 3881 5354
rect 3947 5378 4091 5384
rect 3947 5358 3955 5378
rect 3975 5358 4063 5378
rect 4083 5358 4091 5378
rect 3947 5350 4091 5358
rect 3947 5349 3983 5350
rect 4055 5349 4091 5350
rect 4157 5383 4194 5384
rect 4157 5382 4195 5383
rect 4157 5374 4221 5382
rect 4157 5354 4166 5374
rect 4186 5360 4221 5374
rect 4241 5360 4244 5380
rect 4186 5355 4244 5360
rect 4186 5354 4221 5355
rect 3423 5317 3460 5346
rect 3424 5315 3460 5317
rect 3636 5315 3673 5346
rect 3424 5293 3673 5315
rect 3505 5287 3616 5293
rect 3505 5279 3546 5287
rect 3505 5259 3513 5279
rect 3532 5259 3546 5279
rect 3505 5257 3546 5259
rect 3574 5279 3616 5287
rect 3574 5259 3590 5279
rect 3609 5259 3616 5279
rect 3574 5257 3616 5259
rect 3505 5242 3616 5257
rect 3844 5225 3881 5346
rect 4157 5342 4221 5354
rect 3962 5225 3991 5229
rect 4261 5227 4288 5494
rect 4120 5225 4288 5227
rect 3844 5199 4288 5225
rect 3803 4931 3848 4940
rect 3803 4893 3813 4931
rect 3838 4893 3848 4931
rect 3803 4882 3848 4893
rect 3806 4874 3848 4882
rect 3806 4169 3849 4874
rect 3962 4260 3991 5199
rect 4120 5198 4288 5199
rect 4692 5049 4776 5053
rect 5244 5049 5332 7900
rect 5871 7887 5926 7899
rect 5871 7853 5889 7887
rect 5918 7853 5926 7887
rect 5871 7827 5926 7853
rect 5478 7794 5646 7795
rect 5871 7794 5888 7827
rect 5478 7793 5888 7794
rect 5917 7793 5926 7827
rect 5478 7768 5926 7793
rect 5478 7766 5646 7768
rect 5478 7499 5505 7766
rect 5871 7762 5926 7768
rect 5545 7639 5609 7651
rect 5885 7647 5922 7762
rect 6150 7736 6261 7751
rect 6150 7734 6192 7736
rect 6150 7714 6157 7734
rect 6176 7714 6192 7734
rect 6150 7706 6192 7714
rect 6220 7734 6261 7736
rect 6220 7714 6234 7734
rect 6253 7714 6261 7734
rect 6220 7706 6261 7714
rect 6150 7700 6261 7706
rect 6093 7678 6342 7700
rect 6093 7647 6130 7678
rect 6306 7676 6342 7678
rect 6306 7647 6343 7676
rect 5545 7638 5580 7639
rect 5522 7633 5580 7638
rect 5522 7613 5525 7633
rect 5545 7619 5580 7633
rect 5600 7619 5609 7639
rect 5545 7611 5609 7619
rect 5571 7610 5609 7611
rect 5572 7609 5609 7610
rect 5675 7643 5711 7644
rect 5783 7643 5819 7644
rect 5675 7635 5819 7643
rect 5675 7615 5683 7635
rect 5703 7615 5791 7635
rect 5811 7615 5819 7635
rect 5675 7609 5819 7615
rect 5885 7639 5923 7647
rect 5991 7643 6027 7644
rect 5885 7619 5894 7639
rect 5914 7619 5923 7639
rect 5885 7610 5923 7619
rect 5942 7636 6027 7643
rect 5942 7616 5949 7636
rect 5970 7635 6027 7636
rect 5970 7616 5999 7635
rect 5942 7615 5999 7616
rect 6019 7615 6027 7635
rect 5885 7609 5922 7610
rect 5942 7609 6027 7615
rect 6093 7639 6131 7647
rect 6204 7643 6240 7644
rect 6093 7619 6102 7639
rect 6122 7619 6131 7639
rect 6093 7610 6131 7619
rect 6155 7635 6240 7643
rect 6155 7615 6212 7635
rect 6232 7615 6240 7635
rect 6093 7609 6130 7610
rect 6155 7609 6240 7615
rect 6306 7639 6344 7647
rect 6306 7619 6315 7639
rect 6335 7619 6344 7639
rect 6306 7610 6344 7619
rect 6306 7609 6343 7610
rect 5729 7588 5765 7609
rect 6155 7588 6186 7609
rect 6400 7592 6471 8245
rect 6986 8179 7029 8892
rect 7646 8803 7741 8823
rect 7646 8759 7666 8803
rect 7726 8759 7741 8803
rect 7646 8463 7741 8759
rect 7646 8422 7679 8463
rect 7715 8422 7741 8463
rect 7841 8502 7903 8973
rect 9183 8913 9220 8914
rect 9486 8913 9523 9055
rect 9548 9075 9635 9082
rect 9548 9072 9606 9075
rect 9548 9052 9553 9072
rect 9574 9055 9606 9072
rect 9626 9055 9635 9075
rect 9574 9052 9635 9055
rect 9548 9045 9635 9052
rect 9694 9075 9731 9085
rect 9694 9055 9702 9075
rect 9722 9055 9731 9075
rect 9548 9044 9579 9045
rect 9694 8976 9731 9055
rect 9761 9084 9792 9137
rect 10005 9130 10020 9138
rect 10060 9130 10070 9167
rect 11261 9156 11326 9295
rect 11601 9240 11638 9319
rect 11679 9306 11789 9319
rect 11753 9250 11784 9251
rect 11601 9220 11610 9240
rect 11630 9220 11638 9240
rect 10005 9121 10070 9130
rect 10218 9128 10283 9149
rect 10218 9110 10243 9128
rect 10261 9110 10283 9128
rect 11261 9138 11284 9156
rect 11302 9138 11326 9156
rect 11261 9121 11326 9138
rect 11481 9202 11549 9215
rect 11601 9210 11638 9220
rect 11697 9240 11784 9250
rect 11697 9220 11706 9240
rect 11726 9220 11784 9240
rect 11697 9211 11784 9220
rect 11697 9210 11734 9211
rect 11481 9160 11488 9202
rect 11537 9160 11549 9202
rect 11481 9157 11549 9160
rect 11753 9158 11784 9211
rect 11814 9240 11851 9319
rect 11966 9250 11997 9251
rect 11814 9220 11823 9240
rect 11843 9220 11851 9240
rect 11814 9210 11851 9220
rect 11910 9243 11997 9250
rect 11910 9240 11971 9243
rect 11910 9220 11919 9240
rect 11939 9223 11971 9240
rect 11992 9223 11997 9243
rect 11939 9220 11997 9223
rect 11910 9213 11997 9220
rect 12022 9240 12059 9382
rect 12325 9381 12362 9382
rect 13070 9379 13486 9384
rect 13070 9378 13411 9379
rect 12727 9347 12837 9361
rect 12727 9344 12770 9347
rect 12727 9339 12731 9344
rect 12649 9317 12731 9339
rect 12760 9317 12770 9344
rect 12798 9320 12805 9347
rect 12834 9339 12837 9347
rect 12834 9320 12899 9339
rect 12798 9317 12899 9320
rect 12649 9315 12899 9317
rect 12174 9250 12210 9251
rect 12022 9220 12031 9240
rect 12051 9220 12059 9240
rect 11910 9211 11966 9213
rect 11910 9210 11947 9211
rect 12022 9210 12059 9220
rect 12118 9240 12266 9250
rect 12366 9247 12462 9249
rect 12118 9220 12127 9240
rect 12147 9220 12237 9240
rect 12257 9220 12266 9240
rect 12118 9214 12266 9220
rect 12118 9211 12182 9214
rect 12118 9210 12155 9211
rect 12174 9184 12182 9211
rect 12203 9211 12266 9214
rect 12324 9240 12462 9247
rect 12324 9220 12333 9240
rect 12353 9220 12462 9240
rect 12324 9211 12462 9220
rect 12649 9236 12686 9315
rect 12727 9302 12837 9315
rect 12801 9246 12832 9247
rect 12649 9216 12658 9236
rect 12678 9216 12686 9236
rect 12203 9184 12210 9211
rect 12229 9210 12266 9211
rect 12325 9210 12362 9211
rect 12174 9159 12210 9184
rect 11645 9157 11686 9158
rect 11481 9150 11686 9157
rect 11481 9139 11655 9150
rect 9811 9084 9848 9085
rect 9761 9075 9848 9084
rect 9761 9055 9819 9075
rect 9839 9055 9848 9075
rect 9761 9045 9848 9055
rect 9907 9075 9944 9085
rect 9907 9055 9915 9075
rect 9935 9055 9944 9075
rect 9761 9044 9792 9045
rect 9756 8976 9866 8989
rect 9907 8976 9944 9055
rect 10218 9034 10283 9110
rect 11481 9106 11489 9139
rect 11482 9097 11489 9106
rect 11538 9130 11655 9139
rect 11675 9130 11686 9150
rect 11538 9122 11686 9130
rect 11753 9154 12112 9158
rect 11753 9149 12075 9154
rect 11753 9125 11866 9149
rect 11890 9130 12075 9149
rect 12099 9130 12112 9154
rect 11890 9125 12112 9130
rect 11753 9122 12112 9125
rect 12174 9122 12209 9159
rect 12277 9156 12377 9159
rect 12277 9152 12344 9156
rect 12277 9126 12289 9152
rect 12315 9130 12344 9152
rect 12370 9130 12377 9156
rect 12315 9126 12377 9130
rect 12277 9122 12377 9126
rect 11538 9106 11549 9122
rect 11538 9097 11546 9106
rect 11753 9101 11784 9122
rect 12174 9101 12210 9122
rect 11596 9100 11633 9101
rect 11261 9057 11326 9076
rect 11261 9039 11286 9057
rect 11304 9039 11326 9057
rect 9694 8974 9944 8976
rect 9694 8971 9795 8974
rect 9694 8952 9759 8971
rect 9756 8944 9759 8952
rect 9788 8944 9795 8971
rect 9823 8947 9833 8974
rect 9862 8952 9944 8974
rect 9967 8999 10284 9034
rect 9862 8947 9866 8952
rect 9823 8944 9866 8947
rect 9756 8930 9866 8944
rect 9182 8912 9523 8913
rect 9107 8910 9523 8912
rect 9967 8910 10007 8999
rect 10218 8972 10283 8999
rect 10218 8954 10241 8972
rect 10259 8954 10283 8972
rect 10218 8934 10283 8954
rect 9104 8907 10007 8910
rect 9104 8887 9110 8907
rect 9130 8887 10007 8907
rect 9104 8883 10007 8887
rect 9967 8880 10007 8883
rect 10219 8873 10284 8894
rect 8437 8865 9098 8866
rect 8437 8858 9371 8865
rect 8437 8857 9343 8858
rect 8437 8837 9288 8857
rect 9320 8838 9343 8857
rect 9368 8838 9371 8858
rect 9320 8837 9371 8838
rect 8437 8830 9371 8837
rect 8036 8788 8204 8789
rect 8439 8788 8478 8830
rect 9267 8828 9371 8830
rect 9336 8826 9371 8828
rect 10219 8855 10243 8873
rect 10261 8855 10284 8873
rect 10219 8808 10284 8855
rect 8036 8762 8480 8788
rect 8036 8760 8204 8762
rect 7841 8483 7905 8502
rect 7841 8444 7858 8483
rect 7892 8444 7905 8483
rect 7841 8425 7905 8444
rect 7646 8396 7741 8422
rect 8036 8409 8063 8760
rect 8439 8756 8480 8762
rect 8103 8549 8167 8561
rect 8443 8557 8480 8756
rect 8942 8783 9014 8800
rect 8942 8744 8950 8783
rect 8995 8744 9014 8783
rect 8708 8646 8819 8661
rect 8708 8644 8750 8646
rect 8708 8624 8715 8644
rect 8734 8624 8750 8644
rect 8708 8616 8750 8624
rect 8778 8644 8819 8646
rect 8778 8624 8792 8644
rect 8811 8624 8819 8644
rect 8778 8616 8819 8624
rect 8708 8610 8819 8616
rect 8651 8588 8900 8610
rect 8651 8557 8688 8588
rect 8864 8586 8900 8588
rect 8864 8557 8901 8586
rect 8103 8548 8138 8549
rect 8080 8543 8138 8548
rect 8080 8523 8083 8543
rect 8103 8529 8138 8543
rect 8158 8529 8167 8549
rect 8103 8521 8167 8529
rect 8129 8520 8167 8521
rect 8130 8519 8167 8520
rect 8233 8553 8269 8554
rect 8341 8553 8377 8554
rect 8233 8545 8377 8553
rect 8233 8525 8241 8545
rect 8261 8525 8349 8545
rect 8369 8525 8377 8545
rect 8233 8519 8377 8525
rect 8443 8549 8481 8557
rect 8549 8553 8585 8554
rect 8443 8529 8452 8549
rect 8472 8529 8481 8549
rect 8443 8520 8481 8529
rect 8500 8546 8585 8553
rect 8500 8526 8507 8546
rect 8528 8545 8585 8546
rect 8528 8526 8557 8545
rect 8500 8525 8557 8526
rect 8577 8525 8585 8545
rect 8443 8519 8480 8520
rect 8500 8519 8585 8525
rect 8651 8549 8689 8557
rect 8762 8553 8798 8554
rect 8651 8529 8660 8549
rect 8680 8529 8689 8549
rect 8651 8520 8689 8529
rect 8713 8545 8798 8553
rect 8713 8525 8770 8545
rect 8790 8525 8798 8545
rect 8651 8519 8688 8520
rect 8713 8519 8798 8525
rect 8864 8549 8902 8557
rect 8864 8529 8873 8549
rect 8893 8529 8902 8549
rect 8864 8520 8902 8529
rect 8942 8534 9014 8744
rect 9084 8778 10284 8808
rect 9084 8777 9528 8778
rect 9084 8775 9252 8777
rect 8942 8520 9025 8534
rect 8864 8519 8901 8520
rect 8287 8498 8323 8519
rect 8713 8498 8744 8519
rect 8942 8498 8959 8520
rect 8120 8494 8220 8498
rect 8120 8490 8182 8494
rect 8120 8464 8127 8490
rect 8153 8468 8182 8490
rect 8208 8468 8220 8494
rect 8153 8464 8220 8468
rect 8120 8461 8220 8464
rect 8288 8461 8323 8498
rect 8385 8495 8744 8498
rect 8385 8490 8607 8495
rect 8385 8466 8398 8490
rect 8422 8471 8607 8490
rect 8631 8471 8744 8495
rect 8422 8466 8744 8471
rect 8385 8462 8744 8466
rect 8811 8490 8959 8498
rect 8811 8470 8822 8490
rect 8842 8487 8959 8490
rect 9012 8487 9025 8520
rect 8842 8470 9025 8487
rect 8811 8463 9025 8470
rect 8811 8462 8852 8463
rect 8942 8462 9025 8463
rect 8287 8436 8323 8461
rect 8135 8409 8172 8410
rect 8231 8409 8268 8410
rect 8287 8409 8294 8436
rect 8035 8400 8173 8409
rect 8035 8380 8144 8400
rect 8164 8380 8173 8400
rect 8035 8373 8173 8380
rect 8231 8406 8294 8409
rect 8315 8409 8323 8436
rect 8342 8409 8379 8410
rect 8315 8406 8379 8409
rect 8231 8400 8379 8406
rect 8231 8380 8240 8400
rect 8260 8380 8350 8400
rect 8370 8380 8379 8400
rect 8035 8371 8131 8373
rect 8231 8370 8379 8380
rect 8438 8400 8475 8410
rect 8550 8409 8587 8410
rect 8531 8407 8587 8409
rect 8438 8380 8446 8400
rect 8466 8380 8475 8400
rect 8287 8369 8323 8370
rect 8135 8238 8172 8239
rect 8438 8238 8475 8380
rect 8500 8400 8587 8407
rect 8500 8397 8558 8400
rect 8500 8377 8505 8397
rect 8526 8380 8558 8397
rect 8578 8380 8587 8400
rect 8526 8377 8587 8380
rect 8500 8370 8587 8377
rect 8646 8400 8683 8410
rect 8646 8380 8654 8400
rect 8674 8380 8683 8400
rect 8500 8369 8531 8370
rect 8646 8301 8683 8380
rect 8713 8409 8744 8462
rect 8950 8429 8964 8462
rect 9017 8429 9025 8462
rect 8950 8423 9025 8429
rect 8950 8418 9020 8423
rect 8763 8409 8800 8410
rect 8713 8400 8800 8409
rect 8713 8380 8771 8400
rect 8791 8380 8800 8400
rect 8713 8370 8800 8380
rect 8859 8400 8896 8410
rect 9084 8405 9111 8775
rect 9151 8545 9215 8557
rect 9491 8553 9528 8777
rect 9999 8758 10063 8760
rect 9995 8746 10063 8758
rect 9995 8713 10006 8746
rect 10046 8713 10063 8746
rect 9995 8703 10063 8713
rect 9756 8642 9867 8657
rect 9756 8640 9798 8642
rect 9756 8620 9763 8640
rect 9782 8620 9798 8640
rect 9756 8612 9798 8620
rect 9826 8640 9867 8642
rect 9826 8620 9840 8640
rect 9859 8620 9867 8640
rect 9826 8612 9867 8620
rect 9756 8606 9867 8612
rect 9699 8584 9948 8606
rect 9699 8553 9736 8584
rect 9912 8582 9948 8584
rect 9912 8553 9949 8582
rect 9151 8544 9186 8545
rect 9128 8539 9186 8544
rect 9128 8519 9131 8539
rect 9151 8525 9186 8539
rect 9206 8525 9215 8545
rect 9151 8517 9215 8525
rect 9177 8516 9215 8517
rect 9178 8515 9215 8516
rect 9281 8549 9317 8550
rect 9389 8549 9425 8550
rect 9281 8541 9425 8549
rect 9281 8521 9289 8541
rect 9309 8521 9397 8541
rect 9417 8521 9425 8541
rect 9281 8515 9425 8521
rect 9491 8545 9529 8553
rect 9597 8549 9633 8550
rect 9491 8525 9500 8545
rect 9520 8525 9529 8545
rect 9491 8516 9529 8525
rect 9548 8542 9633 8549
rect 9548 8522 9555 8542
rect 9576 8541 9633 8542
rect 9576 8522 9605 8541
rect 9548 8521 9605 8522
rect 9625 8521 9633 8541
rect 9491 8515 9528 8516
rect 9548 8515 9633 8521
rect 9699 8545 9737 8553
rect 9810 8549 9846 8550
rect 9699 8525 9708 8545
rect 9728 8525 9737 8545
rect 9699 8516 9737 8525
rect 9761 8541 9846 8549
rect 9761 8521 9818 8541
rect 9838 8521 9846 8541
rect 9699 8515 9736 8516
rect 9761 8515 9846 8521
rect 9912 8545 9950 8553
rect 9912 8525 9921 8545
rect 9941 8525 9950 8545
rect 9912 8516 9950 8525
rect 9999 8519 10063 8703
rect 10219 8577 10284 8778
rect 11261 8838 11326 9039
rect 11482 8913 11546 9097
rect 11595 9091 11633 9100
rect 11595 9071 11604 9091
rect 11624 9071 11633 9091
rect 11595 9063 11633 9071
rect 11699 9095 11784 9101
rect 11809 9100 11846 9101
rect 11699 9075 11707 9095
rect 11727 9075 11784 9095
rect 11699 9067 11784 9075
rect 11808 9091 11846 9100
rect 11808 9071 11817 9091
rect 11837 9071 11846 9091
rect 11699 9066 11735 9067
rect 11808 9063 11846 9071
rect 11912 9095 11997 9101
rect 12017 9100 12054 9101
rect 11912 9075 11920 9095
rect 11940 9094 11997 9095
rect 11940 9075 11969 9094
rect 11912 9074 11969 9075
rect 11990 9074 11997 9094
rect 11912 9067 11997 9074
rect 12016 9091 12054 9100
rect 12016 9071 12025 9091
rect 12045 9071 12054 9091
rect 11912 9066 11948 9067
rect 12016 9063 12054 9071
rect 12120 9095 12264 9101
rect 12120 9075 12128 9095
rect 12148 9075 12236 9095
rect 12256 9075 12264 9095
rect 12120 9067 12264 9075
rect 12120 9066 12156 9067
rect 12228 9066 12264 9067
rect 12330 9100 12367 9101
rect 12330 9099 12368 9100
rect 12330 9091 12394 9099
rect 12330 9071 12339 9091
rect 12359 9077 12394 9091
rect 12414 9077 12417 9097
rect 12359 9072 12417 9077
rect 12359 9071 12394 9072
rect 11596 9034 11633 9063
rect 11597 9032 11633 9034
rect 11809 9032 11846 9063
rect 11597 9010 11846 9032
rect 11678 9004 11789 9010
rect 11678 8996 11719 9004
rect 11678 8976 11686 8996
rect 11705 8976 11719 8996
rect 11678 8974 11719 8976
rect 11747 8996 11789 9004
rect 11747 8976 11763 8996
rect 11782 8976 11789 8996
rect 11747 8974 11789 8976
rect 11678 8959 11789 8974
rect 11482 8903 11550 8913
rect 11482 8870 11499 8903
rect 11539 8870 11550 8903
rect 11482 8858 11550 8870
rect 11482 8856 11546 8858
rect 12017 8839 12054 9063
rect 12330 9059 12394 9071
rect 12434 8841 12461 9211
rect 12649 9206 12686 9216
rect 12745 9236 12832 9246
rect 12745 9216 12754 9236
rect 12774 9216 12832 9236
rect 12745 9207 12832 9216
rect 12745 9206 12782 9207
rect 12525 9193 12595 9198
rect 12520 9187 12595 9193
rect 12520 9154 12528 9187
rect 12581 9154 12595 9187
rect 12801 9154 12832 9207
rect 12862 9236 12899 9315
rect 13014 9246 13045 9247
rect 12862 9216 12871 9236
rect 12891 9216 12899 9236
rect 12862 9206 12899 9216
rect 12958 9239 13045 9246
rect 12958 9236 13019 9239
rect 12958 9216 12967 9236
rect 12987 9219 13019 9236
rect 13040 9219 13045 9239
rect 12987 9216 13045 9219
rect 12958 9209 13045 9216
rect 13070 9236 13107 9378
rect 13373 9377 13410 9378
rect 13222 9246 13258 9247
rect 13070 9216 13079 9236
rect 13099 9216 13107 9236
rect 12958 9207 13014 9209
rect 12958 9206 12995 9207
rect 13070 9206 13107 9216
rect 13166 9236 13314 9246
rect 13414 9243 13510 9245
rect 13166 9216 13175 9236
rect 13195 9216 13285 9236
rect 13305 9216 13314 9236
rect 13166 9210 13314 9216
rect 13166 9207 13230 9210
rect 13166 9206 13203 9207
rect 13222 9180 13230 9207
rect 13251 9207 13314 9210
rect 13372 9236 13510 9243
rect 13372 9216 13381 9236
rect 13401 9216 13510 9236
rect 13372 9207 13510 9216
rect 13251 9180 13258 9207
rect 13277 9206 13314 9207
rect 13373 9206 13410 9207
rect 13222 9155 13258 9180
rect 12520 9153 12603 9154
rect 12693 9153 12734 9154
rect 12520 9146 12734 9153
rect 12520 9129 12703 9146
rect 12520 9096 12533 9129
rect 12586 9126 12703 9129
rect 12723 9126 12734 9146
rect 12586 9118 12734 9126
rect 12801 9150 13160 9154
rect 12801 9145 13123 9150
rect 12801 9121 12914 9145
rect 12938 9126 13123 9145
rect 13147 9126 13160 9150
rect 12938 9121 13160 9126
rect 12801 9118 13160 9121
rect 13222 9118 13257 9155
rect 13325 9152 13425 9155
rect 13325 9148 13392 9152
rect 13325 9122 13337 9148
rect 13363 9126 13392 9148
rect 13418 9126 13425 9152
rect 13363 9122 13425 9126
rect 13325 9118 13425 9122
rect 12586 9096 12603 9118
rect 12801 9097 12832 9118
rect 13222 9097 13258 9118
rect 12644 9096 12681 9097
rect 12520 9082 12603 9096
rect 12293 8839 12461 8841
rect 12017 8838 12461 8839
rect 11261 8808 12461 8838
rect 12531 8872 12603 9082
rect 12643 9087 12681 9096
rect 12643 9067 12652 9087
rect 12672 9067 12681 9087
rect 12643 9059 12681 9067
rect 12747 9091 12832 9097
rect 12857 9096 12894 9097
rect 12747 9071 12755 9091
rect 12775 9071 12832 9091
rect 12747 9063 12832 9071
rect 12856 9087 12894 9096
rect 12856 9067 12865 9087
rect 12885 9067 12894 9087
rect 12747 9062 12783 9063
rect 12856 9059 12894 9067
rect 12960 9091 13045 9097
rect 13065 9096 13102 9097
rect 12960 9071 12968 9091
rect 12988 9090 13045 9091
rect 12988 9071 13017 9090
rect 12960 9070 13017 9071
rect 13038 9070 13045 9090
rect 12960 9063 13045 9070
rect 13064 9087 13102 9096
rect 13064 9067 13073 9087
rect 13093 9067 13102 9087
rect 12960 9062 12996 9063
rect 13064 9059 13102 9067
rect 13168 9091 13312 9097
rect 13168 9071 13176 9091
rect 13196 9071 13284 9091
rect 13304 9071 13312 9091
rect 13168 9063 13312 9071
rect 13168 9062 13204 9063
rect 13276 9062 13312 9063
rect 13378 9096 13415 9097
rect 13378 9095 13416 9096
rect 13378 9087 13442 9095
rect 13378 9067 13387 9087
rect 13407 9073 13442 9087
rect 13462 9073 13465 9093
rect 13407 9068 13465 9073
rect 13407 9067 13442 9068
rect 12644 9030 12681 9059
rect 12645 9028 12681 9030
rect 12857 9028 12894 9059
rect 12645 9006 12894 9028
rect 12726 9000 12837 9006
rect 12726 8992 12767 9000
rect 12726 8972 12734 8992
rect 12753 8972 12767 8992
rect 12726 8970 12767 8972
rect 12795 8992 12837 9000
rect 12795 8972 12811 8992
rect 12830 8972 12837 8992
rect 12795 8970 12837 8972
rect 12726 8955 12837 8970
rect 12531 8833 12550 8872
rect 12595 8833 12603 8872
rect 12531 8816 12603 8833
rect 13065 8860 13102 9059
rect 13378 9055 13442 9067
rect 13065 8854 13106 8860
rect 13482 8856 13509 9207
rect 13341 8854 13509 8856
rect 13065 8828 13509 8854
rect 11261 8761 11326 8808
rect 11261 8743 11284 8761
rect 11302 8743 11326 8761
rect 12174 8788 12209 8790
rect 12174 8786 12278 8788
rect 13067 8786 13106 8828
rect 13341 8827 13509 8828
rect 12174 8779 13108 8786
rect 12174 8778 12225 8779
rect 12174 8758 12177 8778
rect 12202 8759 12225 8778
rect 12257 8759 13108 8779
rect 12202 8758 13108 8759
rect 12174 8751 13108 8758
rect 12447 8750 13108 8751
rect 11261 8722 11326 8743
rect 11538 8733 11578 8736
rect 11538 8729 12441 8733
rect 11538 8709 12415 8729
rect 12435 8709 12441 8729
rect 11538 8706 12441 8709
rect 11262 8662 11327 8682
rect 11262 8644 11286 8662
rect 11304 8644 11327 8662
rect 11262 8617 11327 8644
rect 11538 8617 11578 8706
rect 12022 8704 12438 8706
rect 12022 8703 12363 8704
rect 11679 8672 11789 8686
rect 11679 8669 11722 8672
rect 11679 8664 11683 8669
rect 11261 8582 11578 8617
rect 11601 8642 11683 8664
rect 11712 8642 11722 8669
rect 11750 8645 11757 8672
rect 11786 8664 11789 8672
rect 11786 8645 11851 8664
rect 11750 8642 11851 8645
rect 11601 8640 11851 8642
rect 10219 8559 10241 8577
rect 10259 8559 10284 8577
rect 10219 8540 10284 8559
rect 9912 8515 9949 8516
rect 9335 8494 9371 8515
rect 9761 8494 9792 8515
rect 9999 8510 10007 8519
rect 9996 8494 10007 8510
rect 9168 8490 9268 8494
rect 9168 8486 9230 8490
rect 9168 8460 9175 8486
rect 9201 8464 9230 8486
rect 9256 8464 9268 8490
rect 9201 8460 9268 8464
rect 9168 8457 9268 8460
rect 9336 8457 9371 8494
rect 9433 8491 9792 8494
rect 9433 8486 9655 8491
rect 9433 8462 9446 8486
rect 9470 8467 9655 8486
rect 9679 8467 9792 8491
rect 9470 8462 9792 8467
rect 9433 8458 9792 8462
rect 9859 8486 10007 8494
rect 9859 8466 9870 8486
rect 9890 8477 10007 8486
rect 10056 8510 10063 8519
rect 10056 8477 10064 8510
rect 11262 8506 11327 8582
rect 11601 8561 11638 8640
rect 11679 8627 11789 8640
rect 11753 8571 11784 8572
rect 11601 8541 11610 8561
rect 11630 8541 11638 8561
rect 11601 8531 11638 8541
rect 11697 8561 11784 8571
rect 11697 8541 11706 8561
rect 11726 8541 11784 8561
rect 11697 8532 11784 8541
rect 11697 8531 11734 8532
rect 9890 8466 10064 8477
rect 9859 8459 10064 8466
rect 9859 8458 9900 8459
rect 9335 8432 9371 8457
rect 9183 8405 9220 8406
rect 9279 8405 9316 8406
rect 9335 8405 9342 8432
rect 8859 8380 8867 8400
rect 8887 8380 8896 8400
rect 8713 8369 8744 8370
rect 8708 8301 8818 8314
rect 8859 8301 8896 8380
rect 9083 8396 9221 8405
rect 9083 8376 9192 8396
rect 9212 8376 9221 8396
rect 9083 8369 9221 8376
rect 9279 8402 9342 8405
rect 9363 8405 9371 8432
rect 9390 8405 9427 8406
rect 9363 8402 9427 8405
rect 9279 8396 9427 8402
rect 9279 8376 9288 8396
rect 9308 8376 9398 8396
rect 9418 8376 9427 8396
rect 9083 8367 9179 8369
rect 9279 8366 9427 8376
rect 9486 8396 9523 8406
rect 9598 8405 9635 8406
rect 9579 8403 9635 8405
rect 9486 8376 9494 8396
rect 9514 8376 9523 8396
rect 9335 8365 9371 8366
rect 8646 8299 8896 8301
rect 8646 8296 8747 8299
rect 8646 8277 8711 8296
rect 8708 8269 8711 8277
rect 8740 8269 8747 8296
rect 8775 8272 8785 8299
rect 8814 8277 8896 8299
rect 8814 8272 8818 8277
rect 8775 8269 8818 8272
rect 8708 8255 8818 8269
rect 8134 8237 8475 8238
rect 8059 8232 8475 8237
rect 9183 8234 9220 8235
rect 9486 8234 9523 8376
rect 9548 8396 9635 8403
rect 9548 8393 9606 8396
rect 9548 8373 9553 8393
rect 9574 8376 9606 8393
rect 9626 8376 9635 8396
rect 9574 8373 9635 8376
rect 9548 8366 9635 8373
rect 9694 8396 9731 8406
rect 9694 8376 9702 8396
rect 9722 8376 9731 8396
rect 9548 8365 9579 8366
rect 9694 8297 9731 8376
rect 9761 8405 9792 8458
rect 9996 8456 10064 8459
rect 9996 8414 10008 8456
rect 10057 8414 10064 8456
rect 9811 8405 9848 8406
rect 9761 8396 9848 8405
rect 9761 8376 9819 8396
rect 9839 8376 9848 8396
rect 9761 8366 9848 8376
rect 9907 8396 9944 8406
rect 9996 8401 10064 8414
rect 10219 8478 10284 8495
rect 10219 8460 10243 8478
rect 10261 8460 10284 8478
rect 11262 8488 11284 8506
rect 11302 8488 11327 8506
rect 11262 8467 11327 8488
rect 11475 8486 11540 8495
rect 9907 8376 9915 8396
rect 9935 8376 9944 8396
rect 9761 8365 9792 8366
rect 9756 8297 9866 8310
rect 9907 8297 9944 8376
rect 10219 8321 10284 8460
rect 11475 8449 11485 8486
rect 11525 8478 11540 8486
rect 11753 8479 11784 8532
rect 11814 8561 11851 8640
rect 11966 8571 11997 8572
rect 11814 8541 11823 8561
rect 11843 8541 11851 8561
rect 11814 8531 11851 8541
rect 11910 8564 11997 8571
rect 11910 8561 11971 8564
rect 11910 8541 11919 8561
rect 11939 8544 11971 8561
rect 11992 8544 11997 8564
rect 11939 8541 11997 8544
rect 11910 8534 11997 8541
rect 12022 8561 12059 8703
rect 12325 8702 12362 8703
rect 12174 8571 12210 8572
rect 12022 8541 12031 8561
rect 12051 8541 12059 8561
rect 11910 8532 11966 8534
rect 11910 8531 11947 8532
rect 12022 8531 12059 8541
rect 12118 8561 12266 8571
rect 12366 8568 12462 8570
rect 12118 8541 12127 8561
rect 12147 8541 12237 8561
rect 12257 8541 12266 8561
rect 12118 8535 12266 8541
rect 12118 8532 12182 8535
rect 12118 8531 12155 8532
rect 12174 8505 12182 8532
rect 12203 8532 12266 8535
rect 12324 8561 12462 8568
rect 12324 8541 12333 8561
rect 12353 8541 12462 8561
rect 12324 8532 12462 8541
rect 12203 8505 12210 8532
rect 12229 8531 12266 8532
rect 12325 8531 12362 8532
rect 12174 8480 12210 8505
rect 11645 8478 11686 8479
rect 11525 8471 11686 8478
rect 11525 8451 11655 8471
rect 11675 8451 11686 8471
rect 11525 8449 11686 8451
rect 11475 8443 11686 8449
rect 11753 8475 12112 8479
rect 11753 8470 12075 8475
rect 11753 8446 11866 8470
rect 11890 8451 12075 8470
rect 12099 8451 12112 8475
rect 11890 8446 12112 8451
rect 11753 8443 12112 8446
rect 12174 8443 12209 8480
rect 12277 8477 12377 8480
rect 12277 8473 12344 8477
rect 12277 8447 12289 8473
rect 12315 8451 12344 8473
rect 12370 8451 12377 8477
rect 12315 8447 12377 8451
rect 12277 8443 12377 8447
rect 11475 8430 11542 8443
rect 10219 8315 10241 8321
rect 9694 8295 9944 8297
rect 9694 8292 9795 8295
rect 9694 8273 9759 8292
rect 9756 8265 9759 8273
rect 9788 8265 9795 8292
rect 9823 8268 9833 8295
rect 9862 8273 9944 8295
rect 9973 8303 10241 8315
rect 10259 8303 10284 8321
rect 9973 8280 10284 8303
rect 11267 8407 11323 8427
rect 11267 8389 11286 8407
rect 11304 8389 11323 8407
rect 9973 8279 10028 8280
rect 9862 8268 9866 8273
rect 9823 8265 9866 8268
rect 9756 8251 9866 8265
rect 9182 8233 9523 8234
rect 8059 8212 8062 8232
rect 8082 8212 8475 8232
rect 9107 8232 9523 8233
rect 9973 8232 10016 8279
rect 11267 8276 11323 8389
rect 11475 8409 11489 8430
rect 11525 8409 11542 8430
rect 11753 8422 11784 8443
rect 12174 8422 12210 8443
rect 11596 8421 11633 8422
rect 11475 8402 11542 8409
rect 11595 8412 11633 8421
rect 9107 8228 10016 8232
rect 6982 8177 7693 8179
rect 8232 8177 8321 8180
rect 6982 8168 8321 8177
rect 6982 8130 8244 8168
rect 8269 8133 8288 8168
rect 8313 8133 8321 8168
rect 8426 8179 8471 8212
rect 9107 8208 9110 8228
rect 9130 8208 10016 8228
rect 9484 8203 10016 8208
rect 10224 8222 10283 8244
rect 10224 8204 10243 8222
rect 10261 8204 10283 8222
rect 9272 8179 9371 8181
rect 8426 8169 9371 8179
rect 8426 8143 9294 8169
rect 8427 8142 9294 8143
rect 8269 8130 8321 8133
rect 6982 8122 8321 8130
rect 9272 8131 9294 8142
rect 9319 8134 9338 8169
rect 9363 8134 9371 8169
rect 9319 8131 9371 8134
rect 9272 8123 9371 8131
rect 10224 8130 10283 8204
rect 11267 8169 11322 8276
rect 11475 8250 11540 8402
rect 11595 8392 11604 8412
rect 11624 8392 11633 8412
rect 11595 8384 11633 8392
rect 11699 8416 11784 8422
rect 11809 8421 11846 8422
rect 11699 8396 11707 8416
rect 11727 8396 11784 8416
rect 11699 8388 11784 8396
rect 11808 8412 11846 8421
rect 11808 8392 11817 8412
rect 11837 8392 11846 8412
rect 11699 8387 11735 8388
rect 11808 8384 11846 8392
rect 11912 8416 11997 8422
rect 12017 8421 12054 8422
rect 11912 8396 11920 8416
rect 11940 8415 11997 8416
rect 11940 8396 11969 8415
rect 11912 8395 11969 8396
rect 11990 8395 11997 8415
rect 11912 8388 11997 8395
rect 12016 8412 12054 8421
rect 12016 8392 12025 8412
rect 12045 8392 12054 8412
rect 11912 8387 11948 8388
rect 12016 8384 12054 8392
rect 12120 8416 12264 8422
rect 12120 8396 12128 8416
rect 12148 8396 12236 8416
rect 12256 8396 12264 8416
rect 12120 8388 12264 8396
rect 12120 8387 12156 8388
rect 12228 8387 12264 8388
rect 12330 8421 12367 8422
rect 12330 8420 12368 8421
rect 12330 8412 12394 8420
rect 12330 8392 12339 8412
rect 12359 8398 12394 8412
rect 12414 8398 12417 8418
rect 12359 8393 12417 8398
rect 12359 8392 12394 8393
rect 11596 8355 11633 8384
rect 11597 8353 11633 8355
rect 11809 8353 11846 8384
rect 11597 8331 11846 8353
rect 11678 8325 11789 8331
rect 11678 8317 11719 8325
rect 11678 8297 11686 8317
rect 11705 8297 11719 8317
rect 11678 8295 11719 8297
rect 11747 8317 11789 8325
rect 11747 8297 11763 8317
rect 11782 8297 11789 8317
rect 11747 8295 11789 8297
rect 11678 8280 11789 8295
rect 12017 8285 12054 8384
rect 12330 8380 12394 8392
rect 11680 8277 11784 8280
rect 11468 8240 11589 8250
rect 11468 8238 11537 8240
rect 11468 8197 11481 8238
rect 11518 8199 11537 8238
rect 11574 8199 11589 8240
rect 11518 8197 11589 8199
rect 11468 8179 11589 8197
rect 9298 8122 9370 8123
rect 6982 8121 8320 8122
rect 6982 8119 7693 8121
rect 7842 8080 7906 8084
rect 10217 8082 10283 8130
rect 11260 8135 11325 8169
rect 11680 8135 11784 8137
rect 12015 8135 12056 8285
rect 12434 8277 12461 8532
rect 12523 8522 12603 8533
rect 12523 8496 12540 8522
rect 12580 8496 12603 8522
rect 12523 8469 12603 8496
rect 12523 8443 12544 8469
rect 12584 8443 12603 8469
rect 12523 8424 12603 8443
rect 12523 8398 12547 8424
rect 12587 8398 12603 8424
rect 12523 8347 12603 8398
rect 11260 8132 12056 8135
rect 12435 8146 12461 8277
rect 12525 8147 12595 8347
rect 12435 8132 12463 8146
rect 11260 8097 12463 8132
rect 12524 8125 12596 8147
rect 7842 8071 7916 8080
rect 6357 7588 6471 7592
rect 5562 7584 5662 7588
rect 5562 7580 5624 7584
rect 5562 7554 5569 7580
rect 5595 7558 5624 7580
rect 5650 7558 5662 7584
rect 5595 7554 5662 7558
rect 5562 7551 5662 7554
rect 5730 7551 5765 7588
rect 5827 7585 6186 7588
rect 5827 7580 6049 7585
rect 5827 7556 5840 7580
rect 5864 7561 6049 7580
rect 6073 7561 6186 7585
rect 5864 7556 6186 7561
rect 5827 7552 6186 7556
rect 6253 7585 6471 7588
rect 6253 7584 6436 7585
rect 6253 7580 6379 7584
rect 6253 7560 6264 7580
rect 6284 7560 6379 7580
rect 6403 7561 6436 7584
rect 6460 7561 6471 7585
rect 6403 7560 6471 7561
rect 6253 7553 6471 7560
rect 6253 7552 6294 7553
rect 5729 7526 5765 7551
rect 5577 7499 5614 7500
rect 5673 7499 5710 7500
rect 5729 7499 5736 7526
rect 5477 7490 5615 7499
rect 5477 7470 5586 7490
rect 5606 7470 5615 7490
rect 5477 7463 5615 7470
rect 5673 7496 5736 7499
rect 5757 7499 5765 7526
rect 5784 7499 5821 7500
rect 5757 7496 5821 7499
rect 5673 7490 5821 7496
rect 5673 7470 5682 7490
rect 5702 7470 5792 7490
rect 5812 7470 5821 7490
rect 5477 7461 5573 7463
rect 5673 7460 5821 7470
rect 5880 7490 5917 7500
rect 5992 7499 6029 7500
rect 5973 7497 6029 7499
rect 5880 7470 5888 7490
rect 5908 7470 5917 7490
rect 5729 7459 5765 7460
rect 5577 7328 5614 7329
rect 5880 7328 5917 7470
rect 5942 7490 6029 7497
rect 5942 7487 6000 7490
rect 5942 7467 5947 7487
rect 5968 7470 6000 7487
rect 6020 7470 6029 7490
rect 5968 7467 6029 7470
rect 5942 7460 6029 7467
rect 6088 7490 6125 7500
rect 6088 7470 6096 7490
rect 6116 7470 6125 7490
rect 5942 7459 5973 7460
rect 6088 7391 6125 7470
rect 6155 7499 6186 7552
rect 6357 7550 6471 7553
rect 6400 7518 6471 7550
rect 7646 8029 7730 8054
rect 7646 8001 7661 8029
rect 7705 8001 7730 8029
rect 7646 7972 7730 8001
rect 7842 8023 7856 8071
rect 7893 8023 7916 8071
rect 7842 7995 7916 8023
rect 7646 7944 7658 7972
rect 7702 7944 7730 7972
rect 7646 7923 7730 7944
rect 6205 7499 6242 7500
rect 6155 7490 6242 7499
rect 6155 7470 6213 7490
rect 6233 7470 6242 7490
rect 6155 7460 6242 7470
rect 6301 7490 6338 7500
rect 6301 7470 6309 7490
rect 6329 7470 6338 7490
rect 6155 7459 6186 7460
rect 6150 7391 6260 7404
rect 6301 7391 6338 7470
rect 6088 7389 6338 7391
rect 6088 7386 6189 7389
rect 6088 7367 6153 7386
rect 6150 7359 6153 7367
rect 6182 7359 6189 7386
rect 6217 7362 6227 7389
rect 6256 7367 6338 7389
rect 6256 7362 6260 7367
rect 6217 7359 6260 7362
rect 6150 7345 6260 7359
rect 5576 7327 5917 7328
rect 5501 7324 5917 7327
rect 5501 7322 5924 7324
rect 5501 7302 5504 7322
rect 5524 7302 5924 7322
rect 4692 4961 5332 5049
rect 4692 4610 4776 4961
rect 5258 4930 5302 4936
rect 5258 4904 5266 4930
rect 5291 4904 5302 4930
rect 5258 4855 5302 4904
rect 5258 4835 5655 4855
rect 5675 4835 5678 4855
rect 5258 4830 5678 4835
rect 5258 4829 5603 4830
rect 5258 4825 5302 4829
rect 5565 4828 5602 4829
rect 4919 4798 5029 4812
rect 4919 4795 4962 4798
rect 4919 4790 4923 4795
rect 4841 4768 4923 4790
rect 4952 4768 4962 4795
rect 4990 4771 4997 4798
rect 5026 4790 5029 4798
rect 5026 4771 5091 4790
rect 4990 4768 5091 4771
rect 4841 4766 5091 4768
rect 4841 4687 4878 4766
rect 4919 4753 5029 4766
rect 4993 4697 5024 4698
rect 4841 4667 4850 4687
rect 4870 4667 4878 4687
rect 4841 4657 4878 4667
rect 4937 4687 5024 4697
rect 4937 4667 4946 4687
rect 4966 4667 5024 4687
rect 4937 4658 5024 4667
rect 4937 4657 4974 4658
rect 4692 4604 4801 4610
rect 4993 4605 5024 4658
rect 5054 4687 5091 4766
rect 5206 4697 5237 4698
rect 5054 4667 5063 4687
rect 5083 4667 5091 4687
rect 5054 4657 5091 4667
rect 5150 4690 5237 4697
rect 5150 4687 5211 4690
rect 5150 4667 5159 4687
rect 5179 4670 5211 4687
rect 5232 4670 5237 4690
rect 5179 4667 5237 4670
rect 5150 4660 5237 4667
rect 5262 4687 5299 4825
rect 5414 4697 5450 4698
rect 5262 4667 5271 4687
rect 5291 4667 5299 4687
rect 5150 4658 5206 4660
rect 5150 4657 5187 4658
rect 5262 4657 5299 4667
rect 5358 4687 5506 4697
rect 5606 4694 5702 4696
rect 5358 4667 5367 4687
rect 5387 4667 5477 4687
rect 5497 4667 5506 4687
rect 5358 4661 5506 4667
rect 5358 4658 5422 4661
rect 5358 4657 5395 4658
rect 5414 4631 5422 4658
rect 5443 4658 5506 4661
rect 5564 4687 5702 4694
rect 5564 4667 5573 4687
rect 5593 4667 5702 4687
rect 5564 4658 5702 4667
rect 5443 4631 5450 4658
rect 5469 4657 5506 4658
rect 5565 4657 5602 4658
rect 5414 4606 5450 4631
rect 4885 4604 4926 4605
rect 4692 4597 4926 4604
rect 4692 4577 4895 4597
rect 4915 4577 4926 4597
rect 4692 4569 4926 4577
rect 4993 4601 5352 4605
rect 4993 4596 5315 4601
rect 4993 4572 5106 4596
rect 5130 4577 5315 4596
rect 5339 4577 5352 4601
rect 5130 4572 5352 4577
rect 4993 4569 5352 4572
rect 5414 4569 5449 4606
rect 5517 4603 5617 4606
rect 5517 4599 5584 4603
rect 5517 4573 5529 4599
rect 5555 4577 5584 4599
rect 5610 4577 5617 4603
rect 5555 4573 5617 4577
rect 5517 4569 5617 4573
rect 4692 4551 4801 4569
rect 4993 4548 5024 4569
rect 5414 4548 5450 4569
rect 4836 4547 4873 4548
rect 4835 4538 4873 4547
rect 4835 4518 4844 4538
rect 4864 4518 4873 4538
rect 4835 4510 4873 4518
rect 4939 4542 5024 4548
rect 5049 4547 5086 4548
rect 4939 4522 4947 4542
rect 4967 4522 5024 4542
rect 4939 4514 5024 4522
rect 5048 4538 5086 4547
rect 5048 4518 5057 4538
rect 5077 4518 5086 4538
rect 4939 4513 4975 4514
rect 5048 4510 5086 4518
rect 5152 4542 5237 4548
rect 5257 4547 5294 4548
rect 5152 4522 5160 4542
rect 5180 4541 5237 4542
rect 5180 4522 5209 4541
rect 5152 4521 5209 4522
rect 5230 4521 5237 4541
rect 5152 4514 5237 4521
rect 5256 4538 5294 4547
rect 5256 4518 5265 4538
rect 5285 4518 5294 4538
rect 5152 4513 5188 4514
rect 5256 4510 5294 4518
rect 5360 4543 5504 4548
rect 5360 4542 5413 4543
rect 5360 4522 5368 4542
rect 5388 4523 5413 4542
rect 5446 4542 5504 4543
rect 5446 4523 5476 4542
rect 5388 4522 5476 4523
rect 5496 4522 5504 4542
rect 5360 4514 5504 4522
rect 5360 4513 5396 4514
rect 5468 4513 5504 4514
rect 5570 4547 5607 4548
rect 5570 4546 5608 4547
rect 5570 4538 5634 4546
rect 5570 4518 5579 4538
rect 5599 4524 5634 4538
rect 5654 4524 5657 4544
rect 5599 4519 5657 4524
rect 5599 4518 5634 4519
rect 4836 4481 4873 4510
rect 4837 4479 4873 4481
rect 5049 4479 5086 4510
rect 4837 4457 5086 4479
rect 4918 4451 5029 4457
rect 4918 4443 4959 4451
rect 4918 4423 4926 4443
rect 4945 4423 4959 4443
rect 4918 4421 4959 4423
rect 4987 4443 5029 4451
rect 4987 4423 5003 4443
rect 5022 4423 5029 4443
rect 4987 4421 5029 4423
rect 4918 4406 5029 4421
rect 5257 4389 5294 4510
rect 5570 4506 5634 4518
rect 5674 4395 5701 4658
rect 5728 4404 5764 4411
rect 5728 4395 5734 4404
rect 5652 4391 5734 4395
rect 5533 4389 5734 4391
rect 5257 4366 5734 4389
rect 5757 4366 5764 4404
rect 5257 4363 5764 4366
rect 5533 4362 5701 4363
rect 5728 4360 5764 4363
rect 5846 4262 5924 7302
rect 6980 6555 7039 6565
rect 6980 6527 6993 6555
rect 7021 6527 7039 6555
rect 6980 6478 7039 6527
rect 6586 6343 6754 6344
rect 6990 6343 7037 6478
rect 6586 6317 7037 6343
rect 6586 6315 6754 6317
rect 6586 6048 6613 6315
rect 6990 6311 7037 6317
rect 6653 6188 6717 6200
rect 6993 6196 7030 6311
rect 7258 6285 7369 6300
rect 7258 6283 7300 6285
rect 7258 6263 7265 6283
rect 7284 6263 7300 6283
rect 7258 6255 7300 6263
rect 7328 6283 7369 6285
rect 7328 6263 7342 6283
rect 7361 6263 7369 6283
rect 7328 6255 7369 6263
rect 7258 6249 7369 6255
rect 7201 6227 7450 6249
rect 7201 6196 7238 6227
rect 7414 6225 7450 6227
rect 7414 6196 7451 6225
rect 6653 6187 6688 6188
rect 6630 6182 6688 6187
rect 6630 6162 6633 6182
rect 6653 6168 6688 6182
rect 6708 6168 6717 6188
rect 6653 6160 6717 6168
rect 6679 6159 6717 6160
rect 6680 6158 6717 6159
rect 6783 6192 6819 6193
rect 6891 6192 6927 6193
rect 6783 6184 6927 6192
rect 6783 6164 6791 6184
rect 6811 6164 6899 6184
rect 6919 6164 6927 6184
rect 6783 6158 6927 6164
rect 6993 6188 7031 6196
rect 7099 6192 7135 6193
rect 6993 6168 7002 6188
rect 7022 6168 7031 6188
rect 6993 6159 7031 6168
rect 7050 6185 7135 6192
rect 7050 6165 7057 6185
rect 7078 6184 7135 6185
rect 7078 6165 7107 6184
rect 7050 6164 7107 6165
rect 7127 6164 7135 6184
rect 6993 6158 7030 6159
rect 7050 6158 7135 6164
rect 7201 6188 7239 6196
rect 7312 6192 7348 6193
rect 7201 6168 7210 6188
rect 7230 6168 7239 6188
rect 7201 6159 7239 6168
rect 7263 6184 7348 6192
rect 7263 6164 7320 6184
rect 7340 6164 7348 6184
rect 7201 6158 7238 6159
rect 7263 6158 7348 6164
rect 7414 6188 7452 6196
rect 7414 6168 7423 6188
rect 7443 6168 7452 6188
rect 7414 6159 7452 6168
rect 7414 6158 7451 6159
rect 6837 6137 6873 6158
rect 7263 6137 7294 6158
rect 7474 6143 7531 6151
rect 7474 6137 7482 6143
rect 6670 6133 6770 6137
rect 6670 6129 6732 6133
rect 6670 6103 6677 6129
rect 6703 6107 6732 6129
rect 6758 6107 6770 6133
rect 6703 6103 6770 6107
rect 6670 6100 6770 6103
rect 6838 6100 6873 6137
rect 6935 6134 7294 6137
rect 6935 6129 7157 6134
rect 6935 6105 6948 6129
rect 6972 6110 7157 6129
rect 7181 6110 7294 6134
rect 6972 6105 7294 6110
rect 6935 6101 7294 6105
rect 7361 6129 7482 6137
rect 7361 6109 7372 6129
rect 7392 6120 7482 6129
rect 7508 6120 7531 6143
rect 7392 6109 7531 6120
rect 7361 6107 7531 6109
rect 7361 6102 7482 6107
rect 7361 6101 7402 6102
rect 6837 6075 6873 6100
rect 6685 6048 6722 6049
rect 6781 6048 6818 6049
rect 6837 6048 6844 6075
rect 6585 6039 6723 6048
rect 6585 6019 6694 6039
rect 6714 6019 6723 6039
rect 6585 6012 6723 6019
rect 6781 6045 6844 6048
rect 6865 6048 6873 6075
rect 6892 6048 6929 6049
rect 6865 6045 6929 6048
rect 6781 6039 6929 6045
rect 6781 6019 6790 6039
rect 6810 6019 6900 6039
rect 6920 6019 6929 6039
rect 6585 6010 6681 6012
rect 6781 6009 6929 6019
rect 6988 6039 7025 6049
rect 7100 6048 7137 6049
rect 7081 6046 7137 6048
rect 6988 6019 6996 6039
rect 7016 6019 7025 6039
rect 6837 6008 6873 6009
rect 6685 5877 6722 5878
rect 6988 5877 7025 6019
rect 7050 6039 7137 6046
rect 7050 6036 7108 6039
rect 7050 6016 7055 6036
rect 7076 6019 7108 6036
rect 7128 6019 7137 6039
rect 7076 6016 7137 6019
rect 7050 6009 7137 6016
rect 7196 6039 7233 6049
rect 7196 6019 7204 6039
rect 7224 6019 7233 6039
rect 7050 6008 7081 6009
rect 7196 5940 7233 6019
rect 7263 6048 7294 6101
rect 7313 6048 7350 6049
rect 7263 6039 7350 6048
rect 7263 6019 7321 6039
rect 7341 6019 7350 6039
rect 7263 6009 7350 6019
rect 7409 6039 7446 6049
rect 7409 6019 7417 6039
rect 7437 6019 7446 6039
rect 7263 6008 7294 6009
rect 7258 5940 7368 5953
rect 7409 5940 7446 6019
rect 7196 5938 7446 5940
rect 7196 5935 7297 5938
rect 7196 5916 7261 5935
rect 7258 5908 7261 5916
rect 7290 5908 7297 5935
rect 7325 5911 7335 5938
rect 7364 5916 7446 5938
rect 7364 5911 7368 5916
rect 7325 5908 7368 5911
rect 7258 5894 7368 5908
rect 6684 5876 7025 5877
rect 6609 5871 7025 5876
rect 6609 5851 6612 5871
rect 6632 5851 7026 5871
rect 6835 5818 6872 5828
rect 6835 5781 6844 5818
rect 6861 5781 6872 5818
rect 6835 5760 6872 5781
rect 6544 4821 6712 4822
rect 6841 4821 6870 5760
rect 6983 5146 7026 5851
rect 6984 5138 7026 5146
rect 6984 5127 7029 5138
rect 6984 5089 6994 5127
rect 7019 5089 7029 5127
rect 6984 5080 7029 5089
rect 6544 4795 6988 4821
rect 6544 4793 6712 4795
rect 6544 4526 6571 4793
rect 6841 4791 6870 4795
rect 6611 4666 6675 4678
rect 6951 4674 6988 4795
rect 7216 4763 7327 4778
rect 7216 4761 7258 4763
rect 7216 4741 7223 4761
rect 7242 4741 7258 4761
rect 7216 4733 7258 4741
rect 7286 4761 7327 4763
rect 7286 4741 7300 4761
rect 7319 4741 7327 4761
rect 7286 4733 7327 4741
rect 7216 4727 7327 4733
rect 7159 4705 7408 4727
rect 7159 4674 7196 4705
rect 7372 4703 7408 4705
rect 7372 4674 7409 4703
rect 6611 4665 6646 4666
rect 6588 4660 6646 4665
rect 6588 4640 6591 4660
rect 6611 4646 6646 4660
rect 6666 4646 6675 4666
rect 6611 4638 6675 4646
rect 6637 4637 6675 4638
rect 6638 4636 6675 4637
rect 6741 4670 6777 4671
rect 6849 4670 6885 4671
rect 6741 4662 6885 4670
rect 6741 4642 6749 4662
rect 6769 4642 6857 4662
rect 6877 4642 6885 4662
rect 6741 4636 6885 4642
rect 6951 4666 6989 4674
rect 7057 4670 7093 4671
rect 6951 4646 6960 4666
rect 6980 4646 6989 4666
rect 6951 4637 6989 4646
rect 7008 4663 7093 4670
rect 7008 4643 7015 4663
rect 7036 4662 7093 4663
rect 7036 4643 7065 4662
rect 7008 4642 7065 4643
rect 7085 4642 7093 4662
rect 6951 4636 6988 4637
rect 7008 4636 7093 4642
rect 7159 4666 7197 4674
rect 7270 4670 7306 4671
rect 7159 4646 7168 4666
rect 7188 4646 7197 4666
rect 7159 4637 7197 4646
rect 7221 4662 7306 4670
rect 7221 4642 7278 4662
rect 7298 4642 7306 4662
rect 7159 4636 7196 4637
rect 7221 4636 7306 4642
rect 7372 4666 7410 4674
rect 7372 4646 7381 4666
rect 7401 4646 7410 4666
rect 7372 4637 7410 4646
rect 7372 4636 7409 4637
rect 6795 4615 6831 4636
rect 7221 4615 7252 4636
rect 7646 4619 7738 7923
rect 7844 6156 7916 7995
rect 8946 7945 9018 7962
rect 8946 7897 8958 7945
rect 9004 7897 9018 7945
rect 9486 7925 9527 7927
rect 9758 7925 9862 7927
rect 10217 7925 10282 8082
rect 11260 7940 11325 8097
rect 11680 8095 11784 8097
rect 12015 8095 12056 8097
rect 12524 8077 12538 8125
rect 12584 8077 12596 8125
rect 12524 8060 12596 8077
rect 13626 8027 13698 9866
rect 13804 8099 13896 11403
rect 14290 11386 14321 11407
rect 14711 11386 14747 11407
rect 14133 11385 14170 11386
rect 14132 11376 14170 11385
rect 14132 11356 14141 11376
rect 14161 11356 14170 11376
rect 14132 11348 14170 11356
rect 14236 11380 14321 11386
rect 14346 11385 14383 11386
rect 14236 11360 14244 11380
rect 14264 11360 14321 11380
rect 14236 11352 14321 11360
rect 14345 11376 14383 11385
rect 14345 11356 14354 11376
rect 14374 11356 14383 11376
rect 14236 11351 14272 11352
rect 14345 11348 14383 11356
rect 14449 11380 14534 11386
rect 14554 11385 14591 11386
rect 14449 11360 14457 11380
rect 14477 11379 14534 11380
rect 14477 11360 14506 11379
rect 14449 11359 14506 11360
rect 14527 11359 14534 11379
rect 14449 11352 14534 11359
rect 14553 11376 14591 11385
rect 14553 11356 14562 11376
rect 14582 11356 14591 11376
rect 14449 11351 14485 11352
rect 14553 11348 14591 11356
rect 14657 11380 14801 11386
rect 14657 11360 14665 11380
rect 14685 11360 14773 11380
rect 14793 11360 14801 11380
rect 14657 11352 14801 11360
rect 14657 11351 14693 11352
rect 14765 11351 14801 11352
rect 14867 11385 14904 11386
rect 14867 11384 14905 11385
rect 14867 11376 14931 11384
rect 14867 11356 14876 11376
rect 14896 11362 14931 11376
rect 14951 11362 14954 11382
rect 14896 11357 14954 11362
rect 14896 11356 14931 11357
rect 14133 11319 14170 11348
rect 14134 11317 14170 11319
rect 14346 11317 14383 11348
rect 14134 11295 14383 11317
rect 14215 11289 14326 11295
rect 14215 11281 14256 11289
rect 14215 11261 14223 11281
rect 14242 11261 14256 11281
rect 14215 11259 14256 11261
rect 14284 11281 14326 11289
rect 14284 11261 14300 11281
rect 14319 11261 14326 11281
rect 14284 11259 14326 11261
rect 14215 11244 14326 11259
rect 14554 11227 14591 11348
rect 14867 11344 14931 11356
rect 14672 11227 14701 11231
rect 14971 11229 14998 11496
rect 14830 11227 14998 11229
rect 14554 11201 14998 11227
rect 14513 10933 14558 10942
rect 14513 10895 14523 10933
rect 14548 10895 14558 10933
rect 14513 10884 14558 10895
rect 14516 10876 14558 10884
rect 14516 10171 14559 10876
rect 14672 10262 14701 11201
rect 14830 11200 14998 11201
rect 14670 10241 14707 10262
rect 14670 10204 14681 10241
rect 14698 10204 14707 10241
rect 14670 10194 14707 10204
rect 14516 10151 14910 10171
rect 14930 10151 14933 10171
rect 14517 10146 14933 10151
rect 14517 10145 14858 10146
rect 14174 10114 14284 10128
rect 14174 10111 14217 10114
rect 14174 10106 14178 10111
rect 14096 10084 14178 10106
rect 14207 10084 14217 10111
rect 14245 10087 14252 10114
rect 14281 10106 14284 10114
rect 14281 10087 14346 10106
rect 14245 10084 14346 10087
rect 14096 10082 14346 10084
rect 14096 10003 14133 10082
rect 14174 10069 14284 10082
rect 14248 10013 14279 10014
rect 14096 9983 14105 10003
rect 14125 9983 14133 10003
rect 14096 9973 14133 9983
rect 14192 10003 14279 10013
rect 14192 9983 14201 10003
rect 14221 9983 14279 10003
rect 14192 9974 14279 9983
rect 14192 9973 14229 9974
rect 14248 9921 14279 9974
rect 14309 10003 14346 10082
rect 14461 10013 14492 10014
rect 14309 9983 14318 10003
rect 14338 9983 14346 10003
rect 14309 9973 14346 9983
rect 14405 10006 14492 10013
rect 14405 10003 14466 10006
rect 14405 9983 14414 10003
rect 14434 9986 14466 10003
rect 14487 9986 14492 10006
rect 14434 9983 14492 9986
rect 14405 9976 14492 9983
rect 14517 10003 14554 10145
rect 14820 10144 14857 10145
rect 14669 10013 14705 10014
rect 14517 9983 14526 10003
rect 14546 9983 14554 10003
rect 14405 9974 14461 9976
rect 14405 9973 14442 9974
rect 14517 9973 14554 9983
rect 14613 10003 14761 10013
rect 14861 10010 14957 10012
rect 14613 9983 14622 10003
rect 14642 9983 14732 10003
rect 14752 9983 14761 10003
rect 14613 9977 14761 9983
rect 14613 9974 14677 9977
rect 14613 9973 14650 9974
rect 14669 9947 14677 9974
rect 14698 9974 14761 9977
rect 14819 10003 14957 10010
rect 14819 9983 14828 10003
rect 14848 9983 14957 10003
rect 14819 9974 14957 9983
rect 14698 9947 14705 9974
rect 14724 9973 14761 9974
rect 14820 9973 14857 9974
rect 14669 9922 14705 9947
rect 14140 9920 14181 9921
rect 14060 9915 14181 9920
rect 14011 9913 14181 9915
rect 14011 9902 14150 9913
rect 14011 9879 14034 9902
rect 14060 9893 14150 9902
rect 14170 9893 14181 9913
rect 14060 9885 14181 9893
rect 14248 9917 14607 9921
rect 14248 9912 14570 9917
rect 14248 9888 14361 9912
rect 14385 9893 14570 9912
rect 14594 9893 14607 9917
rect 14385 9888 14607 9893
rect 14248 9885 14607 9888
rect 14669 9885 14704 9922
rect 14772 9919 14872 9922
rect 14772 9915 14839 9919
rect 14772 9889 14784 9915
rect 14810 9893 14839 9915
rect 14865 9893 14872 9919
rect 14810 9889 14872 9893
rect 14772 9885 14872 9889
rect 14060 9879 14068 9885
rect 14011 9871 14068 9879
rect 14248 9864 14279 9885
rect 14669 9864 14705 9885
rect 14091 9863 14128 9864
rect 14090 9854 14128 9863
rect 14090 9834 14099 9854
rect 14119 9834 14128 9854
rect 14090 9826 14128 9834
rect 14194 9858 14279 9864
rect 14304 9863 14341 9864
rect 14194 9838 14202 9858
rect 14222 9838 14279 9858
rect 14194 9830 14279 9838
rect 14303 9854 14341 9863
rect 14303 9834 14312 9854
rect 14332 9834 14341 9854
rect 14194 9829 14230 9830
rect 14303 9826 14341 9834
rect 14407 9858 14492 9864
rect 14512 9863 14549 9864
rect 14407 9838 14415 9858
rect 14435 9857 14492 9858
rect 14435 9838 14464 9857
rect 14407 9837 14464 9838
rect 14485 9837 14492 9857
rect 14407 9830 14492 9837
rect 14511 9854 14549 9863
rect 14511 9834 14520 9854
rect 14540 9834 14549 9854
rect 14407 9829 14443 9830
rect 14511 9826 14549 9834
rect 14615 9858 14759 9864
rect 14615 9838 14623 9858
rect 14643 9838 14731 9858
rect 14751 9838 14759 9858
rect 14615 9830 14759 9838
rect 14615 9829 14651 9830
rect 14723 9829 14759 9830
rect 14825 9863 14862 9864
rect 14825 9862 14863 9863
rect 14825 9854 14889 9862
rect 14825 9834 14834 9854
rect 14854 9840 14889 9854
rect 14909 9840 14912 9860
rect 14854 9835 14912 9840
rect 14854 9834 14889 9835
rect 14091 9797 14128 9826
rect 14092 9795 14128 9797
rect 14304 9795 14341 9826
rect 14092 9773 14341 9795
rect 14173 9767 14284 9773
rect 14173 9759 14214 9767
rect 14173 9739 14181 9759
rect 14200 9739 14214 9759
rect 14173 9737 14214 9739
rect 14242 9759 14284 9767
rect 14242 9739 14258 9759
rect 14277 9739 14284 9759
rect 14242 9737 14284 9739
rect 14173 9722 14284 9737
rect 14512 9711 14549 9826
rect 14825 9822 14889 9834
rect 14505 9705 14552 9711
rect 14929 9707 14956 9974
rect 14788 9705 14956 9707
rect 14505 9679 14956 9705
rect 14505 9544 14552 9679
rect 14788 9678 14956 9679
rect 14503 9495 14562 9544
rect 14503 9467 14521 9495
rect 14549 9467 14562 9495
rect 14503 9457 14562 9467
rect 15618 8720 15696 11760
rect 15618 8700 16018 8720
rect 16038 8700 16041 8720
rect 15618 8698 16041 8700
rect 15625 8695 16041 8698
rect 15625 8694 15966 8695
rect 15282 8663 15392 8677
rect 15282 8660 15325 8663
rect 15282 8655 15286 8660
rect 15204 8633 15286 8655
rect 15315 8633 15325 8660
rect 15353 8636 15360 8663
rect 15389 8655 15392 8663
rect 15389 8636 15454 8655
rect 15353 8633 15454 8636
rect 15204 8631 15454 8633
rect 15204 8552 15241 8631
rect 15282 8618 15392 8631
rect 15356 8562 15387 8563
rect 15204 8532 15213 8552
rect 15233 8532 15241 8552
rect 15204 8522 15241 8532
rect 15300 8552 15387 8562
rect 15300 8532 15309 8552
rect 15329 8532 15387 8552
rect 15300 8523 15387 8532
rect 15300 8522 15337 8523
rect 15074 8469 15185 8472
rect 15356 8470 15387 8523
rect 15417 8552 15454 8631
rect 15569 8562 15600 8563
rect 15417 8532 15426 8552
rect 15446 8532 15454 8552
rect 15417 8522 15454 8532
rect 15513 8555 15600 8562
rect 15513 8552 15574 8555
rect 15513 8532 15522 8552
rect 15542 8535 15574 8552
rect 15595 8535 15600 8555
rect 15542 8532 15600 8535
rect 15513 8525 15600 8532
rect 15625 8552 15662 8694
rect 15928 8693 15965 8694
rect 15777 8562 15813 8563
rect 15625 8532 15634 8552
rect 15654 8532 15662 8552
rect 15513 8523 15569 8525
rect 15513 8522 15550 8523
rect 15625 8522 15662 8532
rect 15721 8552 15869 8562
rect 15969 8559 16065 8561
rect 15721 8532 15730 8552
rect 15750 8532 15840 8552
rect 15860 8532 15869 8552
rect 15721 8526 15869 8532
rect 15721 8523 15785 8526
rect 15721 8522 15758 8523
rect 15777 8496 15785 8523
rect 15806 8523 15869 8526
rect 15927 8552 16065 8559
rect 15927 8532 15936 8552
rect 15956 8532 16065 8552
rect 15927 8523 16065 8532
rect 15806 8496 15813 8523
rect 15832 8522 15869 8523
rect 15928 8522 15965 8523
rect 15777 8471 15813 8496
rect 15248 8469 15289 8470
rect 15074 8462 15289 8469
rect 15074 8461 15139 8462
rect 15074 8437 15082 8461
rect 15106 8438 15139 8461
rect 15163 8442 15258 8462
rect 15278 8442 15289 8462
rect 15163 8438 15289 8442
rect 15106 8437 15289 8438
rect 15074 8434 15289 8437
rect 15356 8466 15715 8470
rect 15356 8461 15678 8466
rect 15356 8437 15469 8461
rect 15493 8442 15678 8461
rect 15702 8442 15715 8466
rect 15493 8437 15715 8442
rect 15356 8434 15715 8437
rect 15777 8434 15812 8471
rect 15880 8468 15980 8471
rect 15880 8464 15947 8468
rect 15880 8438 15892 8464
rect 15918 8442 15947 8464
rect 15973 8442 15980 8468
rect 15918 8438 15980 8442
rect 15880 8434 15980 8438
rect 15074 8430 15185 8434
rect 15356 8413 15387 8434
rect 15777 8413 15813 8434
rect 15199 8412 15236 8413
rect 15198 8403 15236 8412
rect 15198 8383 15207 8403
rect 15227 8383 15236 8403
rect 15198 8375 15236 8383
rect 15302 8407 15387 8413
rect 15412 8412 15449 8413
rect 15302 8387 15310 8407
rect 15330 8387 15387 8407
rect 15302 8379 15387 8387
rect 15411 8403 15449 8412
rect 15411 8383 15420 8403
rect 15440 8383 15449 8403
rect 15302 8378 15338 8379
rect 15411 8375 15449 8383
rect 15515 8407 15600 8413
rect 15620 8412 15657 8413
rect 15515 8387 15523 8407
rect 15543 8406 15600 8407
rect 15543 8387 15572 8406
rect 15515 8386 15572 8387
rect 15593 8386 15600 8406
rect 15515 8379 15600 8386
rect 15619 8403 15657 8412
rect 15619 8383 15628 8403
rect 15648 8383 15657 8403
rect 15515 8378 15551 8379
rect 15619 8375 15657 8383
rect 15723 8407 15867 8413
rect 15723 8387 15731 8407
rect 15751 8406 15839 8407
rect 15751 8387 15785 8406
rect 15723 8384 15785 8387
rect 15809 8387 15839 8406
rect 15859 8387 15867 8407
rect 15809 8384 15867 8387
rect 15723 8379 15867 8384
rect 15723 8378 15759 8379
rect 15831 8378 15867 8379
rect 15933 8412 15970 8413
rect 15933 8411 15971 8412
rect 15933 8403 15997 8411
rect 15933 8383 15942 8403
rect 15962 8389 15997 8403
rect 16017 8389 16020 8409
rect 15962 8384 16020 8389
rect 15962 8383 15997 8384
rect 15199 8346 15236 8375
rect 15200 8344 15236 8346
rect 15412 8344 15449 8375
rect 15200 8322 15449 8344
rect 15281 8316 15392 8322
rect 15281 8308 15322 8316
rect 15281 8288 15289 8308
rect 15308 8288 15322 8308
rect 15281 8286 15322 8288
rect 15350 8308 15392 8316
rect 15350 8288 15366 8308
rect 15385 8288 15392 8308
rect 15350 8286 15392 8288
rect 15281 8271 15392 8286
rect 15620 8260 15657 8375
rect 15933 8371 15997 8383
rect 15616 8254 15671 8260
rect 16037 8256 16064 8523
rect 15896 8254 16064 8256
rect 15616 8229 16064 8254
rect 16377 8314 16483 13567
rect 19649 13555 19668 13581
rect 19708 13555 19729 13581
rect 19649 13528 19729 13555
rect 19649 13502 19672 13528
rect 19712 13502 19729 13528
rect 19649 13491 19729 13502
rect 19791 13492 19818 13747
rect 20196 13739 20237 13889
rect 20468 13885 20572 13889
rect 20924 13850 22285 13889
rect 23138 13903 23237 13911
rect 23138 13900 23190 13903
rect 23138 13865 23146 13900
rect 23171 13865 23190 13900
rect 23215 13892 23237 13903
rect 24188 13904 25527 13912
rect 24188 13901 24240 13904
rect 23215 13891 24082 13892
rect 23215 13865 24083 13891
rect 23138 13855 24083 13865
rect 23138 13853 23237 13855
rect 20663 13827 20784 13845
rect 20663 13825 20734 13827
rect 20663 13784 20678 13825
rect 20715 13786 20734 13825
rect 20771 13786 20784 13827
rect 20715 13784 20784 13786
rect 20663 13774 20784 13784
rect 20468 13744 20572 13746
rect 19858 13632 19922 13644
rect 20198 13640 20235 13739
rect 20463 13729 20574 13744
rect 20463 13727 20505 13729
rect 20463 13707 20470 13727
rect 20489 13707 20505 13727
rect 20463 13699 20505 13707
rect 20533 13727 20574 13729
rect 20533 13707 20547 13727
rect 20566 13707 20574 13727
rect 20533 13699 20574 13707
rect 20463 13693 20574 13699
rect 20406 13671 20655 13693
rect 20406 13640 20443 13671
rect 20619 13669 20655 13671
rect 20619 13640 20656 13669
rect 19858 13631 19893 13632
rect 19835 13626 19893 13631
rect 19835 13606 19838 13626
rect 19858 13612 19893 13626
rect 19913 13612 19922 13632
rect 19858 13604 19922 13612
rect 19884 13603 19922 13604
rect 19885 13602 19922 13603
rect 19988 13636 20024 13637
rect 20096 13636 20132 13637
rect 19988 13628 20132 13636
rect 19988 13608 19996 13628
rect 20016 13608 20104 13628
rect 20124 13608 20132 13628
rect 19988 13602 20132 13608
rect 20198 13632 20236 13640
rect 20304 13636 20340 13637
rect 20198 13612 20207 13632
rect 20227 13612 20236 13632
rect 20198 13603 20236 13612
rect 20255 13629 20340 13636
rect 20255 13609 20262 13629
rect 20283 13628 20340 13629
rect 20283 13609 20312 13628
rect 20255 13608 20312 13609
rect 20332 13608 20340 13628
rect 20198 13602 20235 13603
rect 20255 13602 20340 13608
rect 20406 13632 20444 13640
rect 20517 13636 20553 13637
rect 20406 13612 20415 13632
rect 20435 13612 20444 13632
rect 20406 13603 20444 13612
rect 20468 13628 20553 13636
rect 20468 13608 20525 13628
rect 20545 13608 20553 13628
rect 20406 13602 20443 13603
rect 20468 13602 20553 13608
rect 20619 13632 20657 13640
rect 20619 13612 20628 13632
rect 20648 13612 20657 13632
rect 20712 13622 20777 13774
rect 20930 13748 20985 13850
rect 22226 13830 22285 13850
rect 22226 13812 22248 13830
rect 22266 13812 22285 13830
rect 22226 13790 22285 13812
rect 22493 13826 23025 13831
rect 22493 13806 23379 13826
rect 23399 13806 23402 13826
rect 24038 13822 24083 13855
rect 24188 13866 24196 13901
rect 24221 13866 24240 13901
rect 24265 13866 25527 13904
rect 24188 13857 25527 13866
rect 24188 13854 24277 13857
rect 24816 13855 25527 13857
rect 22493 13802 23402 13806
rect 22493 13755 22536 13802
rect 22986 13801 23402 13802
rect 24034 13802 24427 13822
rect 24447 13802 24450 13822
rect 22986 13800 23327 13801
rect 22643 13769 22753 13783
rect 22643 13766 22686 13769
rect 22643 13761 22647 13766
rect 22481 13754 22536 13755
rect 20619 13603 20657 13612
rect 20710 13615 20777 13622
rect 20619 13602 20656 13603
rect 20042 13581 20078 13602
rect 20468 13581 20499 13602
rect 20710 13594 20727 13615
rect 20763 13594 20777 13615
rect 20929 13635 20985 13748
rect 20929 13617 20948 13635
rect 20966 13617 20985 13635
rect 20929 13597 20985 13617
rect 22225 13731 22536 13754
rect 22225 13713 22250 13731
rect 22268 13719 22536 13731
rect 22565 13739 22647 13761
rect 22676 13739 22686 13766
rect 22714 13742 22721 13769
rect 22750 13761 22753 13769
rect 22750 13742 22815 13761
rect 22714 13739 22815 13742
rect 22565 13737 22815 13739
rect 22268 13713 22290 13719
rect 20710 13581 20777 13594
rect 19875 13577 19975 13581
rect 19875 13573 19937 13577
rect 19875 13547 19882 13573
rect 19908 13551 19937 13573
rect 19963 13551 19975 13577
rect 19908 13547 19975 13551
rect 19875 13544 19975 13547
rect 20043 13544 20078 13581
rect 20140 13578 20499 13581
rect 20140 13573 20362 13578
rect 20140 13549 20153 13573
rect 20177 13554 20362 13573
rect 20386 13554 20499 13578
rect 20177 13549 20499 13554
rect 20140 13545 20499 13549
rect 20566 13575 20777 13581
rect 20566 13573 20727 13575
rect 20566 13553 20577 13573
rect 20597 13553 20727 13573
rect 20566 13546 20727 13553
rect 20566 13545 20607 13546
rect 20042 13519 20078 13544
rect 19890 13492 19927 13493
rect 19986 13492 20023 13493
rect 20042 13492 20049 13519
rect 19790 13483 19928 13492
rect 19790 13463 19899 13483
rect 19919 13463 19928 13483
rect 19790 13456 19928 13463
rect 19986 13489 20049 13492
rect 20070 13492 20078 13519
rect 20097 13492 20134 13493
rect 20070 13489 20134 13492
rect 19986 13483 20134 13489
rect 19986 13463 19995 13483
rect 20015 13463 20105 13483
rect 20125 13463 20134 13483
rect 19790 13454 19886 13456
rect 19986 13453 20134 13463
rect 20193 13483 20230 13493
rect 20305 13492 20342 13493
rect 20286 13490 20342 13492
rect 20193 13463 20201 13483
rect 20221 13463 20230 13483
rect 20042 13452 20078 13453
rect 19890 13321 19927 13322
rect 20193 13321 20230 13463
rect 20255 13483 20342 13490
rect 20255 13480 20313 13483
rect 20255 13460 20260 13480
rect 20281 13463 20313 13480
rect 20333 13463 20342 13483
rect 20281 13460 20342 13463
rect 20255 13453 20342 13460
rect 20401 13483 20438 13493
rect 20401 13463 20409 13483
rect 20429 13463 20438 13483
rect 20255 13452 20286 13453
rect 20401 13384 20438 13463
rect 20468 13492 20499 13545
rect 20712 13538 20727 13546
rect 20767 13538 20777 13575
rect 22225 13574 22290 13713
rect 22565 13658 22602 13737
rect 22643 13724 22753 13737
rect 22717 13668 22748 13669
rect 22565 13638 22574 13658
rect 22594 13638 22602 13658
rect 20712 13529 20777 13538
rect 20925 13536 20990 13557
rect 22225 13556 22248 13574
rect 22266 13556 22290 13574
rect 22225 13539 22290 13556
rect 22445 13620 22513 13633
rect 22565 13628 22602 13638
rect 22661 13658 22748 13668
rect 22661 13638 22670 13658
rect 22690 13638 22748 13658
rect 22661 13629 22748 13638
rect 22661 13628 22698 13629
rect 22445 13578 22452 13620
rect 22501 13578 22513 13620
rect 22445 13575 22513 13578
rect 22717 13576 22748 13629
rect 22778 13658 22815 13737
rect 22930 13668 22961 13669
rect 22778 13638 22787 13658
rect 22807 13638 22815 13658
rect 22778 13628 22815 13638
rect 22874 13661 22961 13668
rect 22874 13658 22935 13661
rect 22874 13638 22883 13658
rect 22903 13641 22935 13658
rect 22956 13641 22961 13661
rect 22903 13638 22961 13641
rect 22874 13631 22961 13638
rect 22986 13658 23023 13800
rect 23289 13799 23326 13800
rect 24034 13797 24450 13802
rect 24034 13796 24375 13797
rect 23691 13765 23801 13779
rect 23691 13762 23734 13765
rect 23691 13757 23695 13762
rect 23613 13735 23695 13757
rect 23724 13735 23734 13762
rect 23762 13738 23769 13765
rect 23798 13757 23801 13765
rect 23798 13738 23863 13757
rect 23762 13735 23863 13738
rect 23613 13733 23863 13735
rect 23138 13668 23174 13669
rect 22986 13638 22995 13658
rect 23015 13638 23023 13658
rect 22874 13629 22930 13631
rect 22874 13628 22911 13629
rect 22986 13628 23023 13638
rect 23082 13658 23230 13668
rect 23330 13665 23426 13667
rect 23082 13638 23091 13658
rect 23111 13638 23201 13658
rect 23221 13638 23230 13658
rect 23082 13632 23230 13638
rect 23082 13629 23146 13632
rect 23082 13628 23119 13629
rect 23138 13602 23146 13629
rect 23167 13629 23230 13632
rect 23288 13658 23426 13665
rect 23288 13638 23297 13658
rect 23317 13638 23426 13658
rect 23288 13629 23426 13638
rect 23613 13654 23650 13733
rect 23691 13720 23801 13733
rect 23765 13664 23796 13665
rect 23613 13634 23622 13654
rect 23642 13634 23650 13654
rect 23167 13602 23174 13629
rect 23193 13628 23230 13629
rect 23289 13628 23326 13629
rect 23138 13577 23174 13602
rect 22609 13575 22650 13576
rect 22445 13568 22650 13575
rect 22445 13557 22619 13568
rect 20925 13518 20950 13536
rect 20968 13518 20990 13536
rect 22445 13524 22453 13557
rect 20518 13492 20555 13493
rect 20468 13483 20555 13492
rect 20468 13463 20526 13483
rect 20546 13463 20555 13483
rect 20468 13453 20555 13463
rect 20614 13483 20651 13493
rect 20614 13463 20622 13483
rect 20642 13463 20651 13483
rect 20468 13452 20499 13453
rect 20463 13384 20573 13397
rect 20614 13384 20651 13463
rect 20925 13442 20990 13518
rect 22446 13515 22453 13524
rect 22502 13548 22619 13557
rect 22639 13548 22650 13568
rect 22502 13540 22650 13548
rect 22717 13572 23076 13576
rect 22717 13567 23039 13572
rect 22717 13543 22830 13567
rect 22854 13548 23039 13567
rect 23063 13548 23076 13572
rect 22854 13543 23076 13548
rect 22717 13540 23076 13543
rect 23138 13540 23173 13577
rect 23241 13574 23341 13577
rect 23241 13570 23308 13574
rect 23241 13544 23253 13570
rect 23279 13548 23308 13570
rect 23334 13548 23341 13574
rect 23279 13544 23341 13548
rect 23241 13540 23341 13544
rect 22502 13524 22513 13540
rect 22502 13515 22510 13524
rect 22717 13519 22748 13540
rect 23138 13519 23174 13540
rect 22560 13518 22597 13519
rect 22225 13475 22290 13494
rect 22225 13457 22250 13475
rect 22268 13457 22290 13475
rect 20401 13382 20651 13384
rect 20401 13379 20502 13382
rect 20401 13360 20466 13379
rect 20463 13352 20466 13360
rect 20495 13352 20502 13379
rect 20530 13355 20540 13382
rect 20569 13360 20651 13382
rect 20674 13407 20991 13442
rect 20569 13355 20573 13360
rect 20530 13352 20573 13355
rect 20463 13338 20573 13352
rect 19889 13320 20230 13321
rect 19814 13318 20230 13320
rect 20674 13318 20714 13407
rect 20925 13380 20990 13407
rect 20925 13362 20948 13380
rect 20966 13362 20990 13380
rect 20925 13342 20990 13362
rect 19811 13315 20714 13318
rect 19811 13295 19817 13315
rect 19837 13295 20714 13315
rect 19811 13291 20714 13295
rect 20674 13288 20714 13291
rect 20926 13281 20991 13302
rect 19144 13273 19805 13274
rect 19144 13266 20078 13273
rect 19144 13265 20050 13266
rect 19144 13245 19995 13265
rect 20027 13246 20050 13265
rect 20075 13246 20078 13266
rect 20027 13245 20078 13246
rect 19144 13238 20078 13245
rect 18743 13196 18911 13197
rect 19146 13196 19185 13238
rect 19974 13236 20078 13238
rect 20043 13234 20078 13236
rect 20926 13263 20950 13281
rect 20968 13263 20991 13281
rect 20926 13216 20991 13263
rect 18743 13170 19187 13196
rect 18743 13168 18911 13170
rect 18743 12817 18770 13168
rect 19146 13164 19187 13170
rect 18810 12957 18874 12969
rect 19150 12965 19187 13164
rect 19649 13191 19721 13208
rect 19649 13152 19657 13191
rect 19702 13152 19721 13191
rect 19415 13054 19526 13069
rect 19415 13052 19457 13054
rect 19415 13032 19422 13052
rect 19441 13032 19457 13052
rect 19415 13024 19457 13032
rect 19485 13052 19526 13054
rect 19485 13032 19499 13052
rect 19518 13032 19526 13052
rect 19485 13024 19526 13032
rect 19415 13018 19526 13024
rect 19358 12996 19607 13018
rect 19358 12965 19395 12996
rect 19571 12994 19607 12996
rect 19571 12965 19608 12994
rect 18810 12956 18845 12957
rect 18787 12951 18845 12956
rect 18787 12931 18790 12951
rect 18810 12937 18845 12951
rect 18865 12937 18874 12957
rect 18810 12929 18874 12937
rect 18836 12928 18874 12929
rect 18837 12927 18874 12928
rect 18940 12961 18976 12962
rect 19048 12961 19084 12962
rect 18940 12953 19084 12961
rect 18940 12933 18948 12953
rect 18968 12933 19056 12953
rect 19076 12933 19084 12953
rect 18940 12927 19084 12933
rect 19150 12957 19188 12965
rect 19256 12961 19292 12962
rect 19150 12937 19159 12957
rect 19179 12937 19188 12957
rect 19150 12928 19188 12937
rect 19207 12954 19292 12961
rect 19207 12934 19214 12954
rect 19235 12953 19292 12954
rect 19235 12934 19264 12953
rect 19207 12933 19264 12934
rect 19284 12933 19292 12953
rect 19150 12927 19187 12928
rect 19207 12927 19292 12933
rect 19358 12957 19396 12965
rect 19469 12961 19505 12962
rect 19358 12937 19367 12957
rect 19387 12937 19396 12957
rect 19358 12928 19396 12937
rect 19420 12953 19505 12961
rect 19420 12933 19477 12953
rect 19497 12933 19505 12953
rect 19358 12927 19395 12928
rect 19420 12927 19505 12933
rect 19571 12957 19609 12965
rect 19571 12937 19580 12957
rect 19600 12937 19609 12957
rect 19571 12928 19609 12937
rect 19649 12942 19721 13152
rect 19791 13186 20991 13216
rect 19791 13185 20235 13186
rect 19791 13183 19959 13185
rect 19649 12928 19732 12942
rect 19571 12927 19608 12928
rect 18994 12906 19030 12927
rect 19420 12906 19451 12927
rect 19649 12906 19666 12928
rect 18827 12902 18927 12906
rect 18827 12898 18889 12902
rect 18827 12872 18834 12898
rect 18860 12876 18889 12898
rect 18915 12876 18927 12902
rect 18860 12872 18927 12876
rect 18827 12869 18927 12872
rect 18995 12869 19030 12906
rect 19092 12903 19451 12906
rect 19092 12898 19314 12903
rect 19092 12874 19105 12898
rect 19129 12879 19314 12898
rect 19338 12879 19451 12903
rect 19129 12874 19451 12879
rect 19092 12870 19451 12874
rect 19518 12898 19666 12906
rect 19518 12878 19529 12898
rect 19549 12895 19666 12898
rect 19719 12895 19732 12928
rect 19549 12878 19732 12895
rect 19518 12871 19732 12878
rect 19518 12870 19559 12871
rect 19649 12870 19732 12871
rect 18994 12844 19030 12869
rect 18842 12817 18879 12818
rect 18938 12817 18975 12818
rect 18994 12817 19001 12844
rect 18742 12808 18880 12817
rect 18742 12788 18851 12808
rect 18871 12788 18880 12808
rect 18742 12781 18880 12788
rect 18938 12814 19001 12817
rect 19022 12817 19030 12844
rect 19049 12817 19086 12818
rect 19022 12814 19086 12817
rect 18938 12808 19086 12814
rect 18938 12788 18947 12808
rect 18967 12788 19057 12808
rect 19077 12788 19086 12808
rect 18742 12779 18838 12781
rect 18938 12778 19086 12788
rect 19145 12808 19182 12818
rect 19257 12817 19294 12818
rect 19238 12815 19294 12817
rect 19145 12788 19153 12808
rect 19173 12788 19182 12808
rect 18994 12777 19030 12778
rect 18842 12646 18879 12647
rect 19145 12646 19182 12788
rect 19207 12808 19294 12815
rect 19207 12805 19265 12808
rect 19207 12785 19212 12805
rect 19233 12788 19265 12805
rect 19285 12788 19294 12808
rect 19233 12785 19294 12788
rect 19207 12778 19294 12785
rect 19353 12808 19390 12818
rect 19353 12788 19361 12808
rect 19381 12788 19390 12808
rect 19207 12777 19238 12778
rect 19353 12709 19390 12788
rect 19420 12817 19451 12870
rect 19657 12837 19671 12870
rect 19724 12837 19732 12870
rect 19657 12831 19732 12837
rect 19657 12826 19727 12831
rect 19470 12817 19507 12818
rect 19420 12808 19507 12817
rect 19420 12788 19478 12808
rect 19498 12788 19507 12808
rect 19420 12778 19507 12788
rect 19566 12808 19603 12818
rect 19791 12813 19818 13183
rect 19858 12953 19922 12965
rect 20198 12961 20235 13185
rect 20706 13166 20770 13168
rect 20702 13154 20770 13166
rect 20702 13121 20713 13154
rect 20753 13121 20770 13154
rect 20702 13111 20770 13121
rect 20463 13050 20574 13065
rect 20463 13048 20505 13050
rect 20463 13028 20470 13048
rect 20489 13028 20505 13048
rect 20463 13020 20505 13028
rect 20533 13048 20574 13050
rect 20533 13028 20547 13048
rect 20566 13028 20574 13048
rect 20533 13020 20574 13028
rect 20463 13014 20574 13020
rect 20406 12992 20655 13014
rect 20406 12961 20443 12992
rect 20619 12990 20655 12992
rect 20619 12961 20656 12990
rect 19858 12952 19893 12953
rect 19835 12947 19893 12952
rect 19835 12927 19838 12947
rect 19858 12933 19893 12947
rect 19913 12933 19922 12953
rect 19858 12925 19922 12933
rect 19884 12924 19922 12925
rect 19885 12923 19922 12924
rect 19988 12957 20024 12958
rect 20096 12957 20132 12958
rect 19988 12949 20132 12957
rect 19988 12929 19996 12949
rect 20016 12929 20104 12949
rect 20124 12929 20132 12949
rect 19988 12923 20132 12929
rect 20198 12953 20236 12961
rect 20304 12957 20340 12958
rect 20198 12933 20207 12953
rect 20227 12933 20236 12953
rect 20198 12924 20236 12933
rect 20255 12950 20340 12957
rect 20255 12930 20262 12950
rect 20283 12949 20340 12950
rect 20283 12930 20312 12949
rect 20255 12929 20312 12930
rect 20332 12929 20340 12949
rect 20198 12923 20235 12924
rect 20255 12923 20340 12929
rect 20406 12953 20444 12961
rect 20517 12957 20553 12958
rect 20406 12933 20415 12953
rect 20435 12933 20444 12953
rect 20406 12924 20444 12933
rect 20468 12949 20553 12957
rect 20468 12929 20525 12949
rect 20545 12929 20553 12949
rect 20406 12923 20443 12924
rect 20468 12923 20553 12929
rect 20619 12953 20657 12961
rect 20619 12933 20628 12953
rect 20648 12933 20657 12953
rect 20619 12924 20657 12933
rect 20706 12927 20770 13111
rect 20926 12985 20991 13186
rect 22225 13256 22290 13457
rect 22446 13331 22510 13515
rect 22559 13509 22597 13518
rect 22559 13489 22568 13509
rect 22588 13489 22597 13509
rect 22559 13481 22597 13489
rect 22663 13513 22748 13519
rect 22773 13518 22810 13519
rect 22663 13493 22671 13513
rect 22691 13493 22748 13513
rect 22663 13485 22748 13493
rect 22772 13509 22810 13518
rect 22772 13489 22781 13509
rect 22801 13489 22810 13509
rect 22663 13484 22699 13485
rect 22772 13481 22810 13489
rect 22876 13513 22961 13519
rect 22981 13518 23018 13519
rect 22876 13493 22884 13513
rect 22904 13512 22961 13513
rect 22904 13493 22933 13512
rect 22876 13492 22933 13493
rect 22954 13492 22961 13512
rect 22876 13485 22961 13492
rect 22980 13509 23018 13518
rect 22980 13489 22989 13509
rect 23009 13489 23018 13509
rect 22876 13484 22912 13485
rect 22980 13481 23018 13489
rect 23084 13513 23228 13519
rect 23084 13493 23092 13513
rect 23112 13493 23200 13513
rect 23220 13493 23228 13513
rect 23084 13485 23228 13493
rect 23084 13484 23120 13485
rect 23192 13484 23228 13485
rect 23294 13518 23331 13519
rect 23294 13517 23332 13518
rect 23294 13509 23358 13517
rect 23294 13489 23303 13509
rect 23323 13495 23358 13509
rect 23378 13495 23381 13515
rect 23323 13490 23381 13495
rect 23323 13489 23358 13490
rect 22560 13452 22597 13481
rect 22561 13450 22597 13452
rect 22773 13450 22810 13481
rect 22561 13428 22810 13450
rect 22642 13422 22753 13428
rect 22642 13414 22683 13422
rect 22642 13394 22650 13414
rect 22669 13394 22683 13414
rect 22642 13392 22683 13394
rect 22711 13414 22753 13422
rect 22711 13394 22727 13414
rect 22746 13394 22753 13414
rect 22711 13392 22753 13394
rect 22642 13377 22753 13392
rect 22446 13321 22514 13331
rect 22446 13288 22463 13321
rect 22503 13288 22514 13321
rect 22446 13276 22514 13288
rect 22446 13274 22510 13276
rect 22981 13257 23018 13481
rect 23294 13477 23358 13489
rect 23398 13259 23425 13629
rect 23613 13624 23650 13634
rect 23709 13654 23796 13664
rect 23709 13634 23718 13654
rect 23738 13634 23796 13654
rect 23709 13625 23796 13634
rect 23709 13624 23746 13625
rect 23489 13611 23559 13616
rect 23484 13605 23559 13611
rect 23484 13572 23492 13605
rect 23545 13572 23559 13605
rect 23765 13572 23796 13625
rect 23826 13654 23863 13733
rect 23978 13664 24009 13665
rect 23826 13634 23835 13654
rect 23855 13634 23863 13654
rect 23826 13624 23863 13634
rect 23922 13657 24009 13664
rect 23922 13654 23983 13657
rect 23922 13634 23931 13654
rect 23951 13637 23983 13654
rect 24004 13637 24009 13657
rect 23951 13634 24009 13637
rect 23922 13627 24009 13634
rect 24034 13654 24071 13796
rect 24337 13795 24374 13796
rect 24186 13664 24222 13665
rect 24034 13634 24043 13654
rect 24063 13634 24071 13654
rect 23922 13625 23978 13627
rect 23922 13624 23959 13625
rect 24034 13624 24071 13634
rect 24130 13654 24278 13664
rect 24378 13661 24474 13663
rect 24130 13634 24139 13654
rect 24159 13634 24249 13654
rect 24269 13634 24278 13654
rect 24130 13628 24278 13634
rect 24130 13625 24194 13628
rect 24130 13624 24167 13625
rect 24186 13598 24194 13625
rect 24215 13625 24278 13628
rect 24336 13654 24474 13661
rect 24336 13634 24345 13654
rect 24365 13634 24474 13654
rect 24336 13625 24474 13634
rect 24215 13598 24222 13625
rect 24241 13624 24278 13625
rect 24337 13624 24374 13625
rect 24186 13573 24222 13598
rect 23484 13571 23567 13572
rect 23657 13571 23698 13572
rect 23484 13564 23698 13571
rect 23484 13547 23667 13564
rect 23484 13514 23497 13547
rect 23550 13544 23667 13547
rect 23687 13544 23698 13564
rect 23550 13536 23698 13544
rect 23765 13568 24124 13572
rect 23765 13563 24087 13568
rect 23765 13539 23878 13563
rect 23902 13544 24087 13563
rect 24111 13544 24124 13568
rect 23902 13539 24124 13544
rect 23765 13536 24124 13539
rect 24186 13536 24221 13573
rect 24289 13570 24389 13573
rect 24289 13566 24356 13570
rect 24289 13540 24301 13566
rect 24327 13544 24356 13566
rect 24382 13544 24389 13570
rect 24327 13540 24389 13544
rect 24289 13536 24389 13540
rect 23550 13514 23567 13536
rect 23765 13515 23796 13536
rect 24186 13515 24222 13536
rect 23608 13514 23645 13515
rect 23484 13500 23567 13514
rect 23257 13257 23425 13259
rect 22981 13256 23425 13257
rect 22225 13226 23425 13256
rect 23495 13290 23567 13500
rect 23607 13505 23645 13514
rect 23607 13485 23616 13505
rect 23636 13485 23645 13505
rect 23607 13477 23645 13485
rect 23711 13509 23796 13515
rect 23821 13514 23858 13515
rect 23711 13489 23719 13509
rect 23739 13489 23796 13509
rect 23711 13481 23796 13489
rect 23820 13505 23858 13514
rect 23820 13485 23829 13505
rect 23849 13485 23858 13505
rect 23711 13480 23747 13481
rect 23820 13477 23858 13485
rect 23924 13509 24009 13515
rect 24029 13514 24066 13515
rect 23924 13489 23932 13509
rect 23952 13508 24009 13509
rect 23952 13489 23981 13508
rect 23924 13488 23981 13489
rect 24002 13488 24009 13508
rect 23924 13481 24009 13488
rect 24028 13505 24066 13514
rect 24028 13485 24037 13505
rect 24057 13485 24066 13505
rect 23924 13480 23960 13481
rect 24028 13477 24066 13485
rect 24132 13509 24276 13515
rect 24132 13489 24140 13509
rect 24160 13489 24248 13509
rect 24268 13489 24276 13509
rect 24132 13481 24276 13489
rect 24132 13480 24168 13481
rect 24240 13480 24276 13481
rect 24342 13514 24379 13515
rect 24342 13513 24380 13514
rect 24342 13505 24406 13513
rect 24342 13485 24351 13505
rect 24371 13491 24406 13505
rect 24426 13491 24429 13511
rect 24371 13486 24429 13491
rect 24371 13485 24406 13486
rect 23608 13448 23645 13477
rect 23609 13446 23645 13448
rect 23821 13446 23858 13477
rect 23609 13424 23858 13446
rect 23690 13418 23801 13424
rect 23690 13410 23731 13418
rect 23690 13390 23698 13410
rect 23717 13390 23731 13410
rect 23690 13388 23731 13390
rect 23759 13410 23801 13418
rect 23759 13390 23775 13410
rect 23794 13390 23801 13410
rect 23759 13388 23801 13390
rect 23690 13373 23801 13388
rect 23495 13251 23514 13290
rect 23559 13251 23567 13290
rect 23495 13234 23567 13251
rect 24029 13278 24066 13477
rect 24342 13473 24406 13485
rect 24029 13272 24070 13278
rect 24446 13274 24473 13625
rect 24768 13612 24863 13638
rect 24604 13590 24668 13609
rect 24604 13551 24617 13590
rect 24651 13551 24668 13590
rect 24604 13532 24668 13551
rect 24305 13272 24473 13274
rect 24029 13246 24473 13272
rect 22225 13179 22290 13226
rect 22225 13161 22248 13179
rect 22266 13161 22290 13179
rect 23138 13206 23173 13208
rect 23138 13204 23242 13206
rect 24031 13204 24070 13246
rect 24305 13245 24473 13246
rect 23138 13197 24072 13204
rect 23138 13196 23189 13197
rect 23138 13176 23141 13196
rect 23166 13177 23189 13196
rect 23221 13177 24072 13197
rect 23166 13176 24072 13177
rect 23138 13169 24072 13176
rect 23411 13168 24072 13169
rect 22225 13140 22290 13161
rect 22502 13151 22542 13154
rect 22502 13147 23405 13151
rect 22502 13127 23379 13147
rect 23399 13127 23405 13147
rect 22502 13124 23405 13127
rect 22226 13080 22291 13100
rect 22226 13062 22250 13080
rect 22268 13062 22291 13080
rect 22226 13035 22291 13062
rect 22502 13035 22542 13124
rect 22986 13122 23402 13124
rect 22986 13121 23327 13122
rect 22643 13090 22753 13104
rect 22643 13087 22686 13090
rect 22643 13082 22647 13087
rect 22225 13000 22542 13035
rect 22565 13060 22647 13082
rect 22676 13060 22686 13087
rect 22714 13063 22721 13090
rect 22750 13082 22753 13090
rect 22750 13063 22815 13082
rect 22714 13060 22815 13063
rect 22565 13058 22815 13060
rect 20926 12967 20948 12985
rect 20966 12967 20991 12985
rect 20926 12948 20991 12967
rect 20619 12923 20656 12924
rect 20042 12902 20078 12923
rect 20468 12902 20499 12923
rect 20706 12918 20714 12927
rect 20703 12902 20714 12918
rect 19875 12898 19975 12902
rect 19875 12894 19937 12898
rect 19875 12868 19882 12894
rect 19908 12872 19937 12894
rect 19963 12872 19975 12898
rect 19908 12868 19975 12872
rect 19875 12865 19975 12868
rect 20043 12865 20078 12902
rect 20140 12899 20499 12902
rect 20140 12894 20362 12899
rect 20140 12870 20153 12894
rect 20177 12875 20362 12894
rect 20386 12875 20499 12899
rect 20177 12870 20499 12875
rect 20140 12866 20499 12870
rect 20566 12894 20714 12902
rect 20566 12874 20577 12894
rect 20597 12885 20714 12894
rect 20763 12918 20770 12927
rect 22226 12924 22291 13000
rect 22565 12979 22602 13058
rect 22643 13045 22753 13058
rect 22717 12989 22748 12990
rect 22565 12959 22574 12979
rect 22594 12959 22602 12979
rect 22565 12949 22602 12959
rect 22661 12979 22748 12989
rect 22661 12959 22670 12979
rect 22690 12959 22748 12979
rect 22661 12950 22748 12959
rect 22661 12949 22698 12950
rect 20763 12885 20771 12918
rect 22226 12906 22248 12924
rect 22266 12906 22291 12924
rect 20597 12874 20771 12885
rect 20566 12867 20771 12874
rect 20566 12866 20607 12867
rect 20042 12840 20078 12865
rect 19890 12813 19927 12814
rect 19986 12813 20023 12814
rect 20042 12813 20049 12840
rect 19566 12788 19574 12808
rect 19594 12788 19603 12808
rect 19420 12777 19451 12778
rect 19415 12709 19525 12722
rect 19566 12709 19603 12788
rect 19790 12804 19928 12813
rect 19790 12784 19899 12804
rect 19919 12784 19928 12804
rect 19790 12777 19928 12784
rect 19986 12810 20049 12813
rect 20070 12813 20078 12840
rect 20097 12813 20134 12814
rect 20070 12810 20134 12813
rect 19986 12804 20134 12810
rect 19986 12784 19995 12804
rect 20015 12784 20105 12804
rect 20125 12784 20134 12804
rect 19790 12775 19886 12777
rect 19986 12774 20134 12784
rect 20193 12804 20230 12814
rect 20305 12813 20342 12814
rect 20286 12811 20342 12813
rect 20193 12784 20201 12804
rect 20221 12784 20230 12804
rect 20042 12773 20078 12774
rect 19353 12707 19603 12709
rect 19353 12704 19454 12707
rect 19353 12685 19418 12704
rect 19415 12677 19418 12685
rect 19447 12677 19454 12704
rect 19482 12680 19492 12707
rect 19521 12685 19603 12707
rect 19521 12680 19525 12685
rect 19482 12677 19525 12680
rect 19415 12663 19525 12677
rect 18841 12645 19182 12646
rect 18766 12640 19182 12645
rect 19890 12642 19927 12643
rect 20193 12642 20230 12784
rect 20255 12804 20342 12811
rect 20255 12801 20313 12804
rect 20255 12781 20260 12801
rect 20281 12784 20313 12801
rect 20333 12784 20342 12804
rect 20281 12781 20342 12784
rect 20255 12774 20342 12781
rect 20401 12804 20438 12814
rect 20401 12784 20409 12804
rect 20429 12784 20438 12804
rect 20255 12773 20286 12774
rect 20401 12705 20438 12784
rect 20468 12813 20499 12866
rect 20703 12864 20771 12867
rect 20703 12822 20715 12864
rect 20764 12822 20771 12864
rect 20518 12813 20555 12814
rect 20468 12804 20555 12813
rect 20468 12784 20526 12804
rect 20546 12784 20555 12804
rect 20468 12774 20555 12784
rect 20614 12804 20651 12814
rect 20703 12809 20771 12822
rect 20926 12886 20991 12903
rect 20926 12868 20950 12886
rect 20968 12868 20991 12886
rect 22226 12885 22291 12906
rect 22439 12904 22504 12913
rect 20614 12784 20622 12804
rect 20642 12784 20651 12804
rect 20468 12773 20499 12774
rect 20463 12705 20573 12718
rect 20614 12705 20651 12784
rect 20926 12729 20991 12868
rect 22439 12867 22449 12904
rect 22489 12896 22504 12904
rect 22717 12897 22748 12950
rect 22778 12979 22815 13058
rect 22930 12989 22961 12990
rect 22778 12959 22787 12979
rect 22807 12959 22815 12979
rect 22778 12949 22815 12959
rect 22874 12982 22961 12989
rect 22874 12979 22935 12982
rect 22874 12959 22883 12979
rect 22903 12962 22935 12979
rect 22956 12962 22961 12982
rect 22903 12959 22961 12962
rect 22874 12952 22961 12959
rect 22986 12979 23023 13121
rect 23289 13120 23326 13121
rect 24606 13061 24668 13532
rect 24768 13571 24794 13612
rect 24830 13571 24863 13612
rect 24768 13275 24863 13571
rect 24768 13231 24783 13275
rect 24843 13231 24863 13275
rect 24768 13211 24863 13231
rect 25480 13142 25523 13855
rect 26556 13745 27449 13785
rect 26556 13678 26589 13745
rect 26675 13678 27457 13745
rect 30622 13681 30692 13934
rect 31161 13931 31202 13933
rect 31433 13931 31537 13933
rect 31873 13931 32996 13964
rect 30754 13896 32996 13931
rect 35524 13907 36235 13909
rect 33847 13905 33919 13906
rect 35405 13905 36235 13907
rect 30754 13882 30782 13896
rect 30756 13751 30782 13882
rect 31161 13894 32996 13896
rect 31161 13893 31304 13894
rect 31562 13893 32996 13894
rect 26556 13610 27457 13678
rect 26565 13609 26671 13610
rect 27340 13516 27457 13610
rect 30614 13630 30694 13681
rect 30614 13604 30630 13630
rect 30670 13604 30694 13630
rect 30614 13585 30694 13604
rect 30614 13559 30633 13585
rect 30673 13559 30694 13585
rect 30614 13532 30694 13559
rect 25480 13122 25874 13142
rect 25894 13122 25897 13142
rect 25481 13117 25897 13122
rect 25481 13116 25822 13117
rect 25138 13085 25248 13099
rect 25138 13082 25181 13085
rect 25138 13077 25142 13082
rect 24601 13009 24676 13061
rect 25060 13055 25142 13077
rect 25171 13055 25181 13082
rect 25209 13058 25216 13085
rect 25245 13077 25248 13085
rect 25245 13058 25310 13077
rect 25209 13055 25310 13058
rect 25060 13053 25310 13055
rect 24970 13009 25016 13010
rect 23138 12989 23174 12990
rect 22986 12959 22995 12979
rect 23015 12959 23023 12979
rect 22874 12950 22930 12952
rect 22874 12949 22911 12950
rect 22986 12949 23023 12959
rect 23082 12979 23230 12989
rect 23330 12986 23426 12988
rect 23082 12959 23091 12979
rect 23111 12959 23201 12979
rect 23221 12959 23230 12979
rect 23082 12953 23230 12959
rect 23082 12950 23146 12953
rect 23082 12949 23119 12950
rect 23138 12923 23146 12950
rect 23167 12950 23230 12953
rect 23288 12979 23426 12986
rect 23288 12959 23297 12979
rect 23317 12959 23426 12979
rect 23288 12950 23426 12959
rect 24601 12974 25016 13009
rect 23167 12923 23174 12950
rect 23193 12949 23230 12950
rect 23289 12949 23326 12950
rect 23138 12898 23174 12923
rect 22609 12896 22650 12897
rect 22489 12889 22650 12896
rect 22489 12869 22619 12889
rect 22639 12869 22650 12889
rect 22489 12867 22650 12869
rect 22439 12861 22650 12867
rect 22717 12893 23076 12897
rect 22717 12888 23039 12893
rect 22717 12864 22830 12888
rect 22854 12869 23039 12888
rect 23063 12869 23076 12893
rect 22854 12864 23076 12869
rect 22717 12861 23076 12864
rect 23138 12861 23173 12898
rect 23241 12895 23341 12898
rect 23241 12891 23308 12895
rect 23241 12865 23253 12891
rect 23279 12869 23308 12891
rect 23334 12869 23341 12895
rect 23279 12865 23341 12869
rect 23241 12861 23341 12865
rect 22439 12848 22506 12861
rect 20926 12723 20948 12729
rect 20401 12703 20651 12705
rect 20401 12700 20502 12703
rect 20401 12681 20466 12700
rect 20463 12673 20466 12681
rect 20495 12673 20502 12700
rect 20530 12676 20540 12703
rect 20569 12681 20651 12703
rect 20680 12711 20948 12723
rect 20966 12711 20991 12729
rect 20680 12688 20991 12711
rect 22231 12825 22287 12845
rect 22231 12807 22250 12825
rect 22268 12807 22287 12825
rect 22231 12694 22287 12807
rect 22439 12827 22453 12848
rect 22489 12827 22506 12848
rect 22717 12840 22748 12861
rect 23138 12840 23174 12861
rect 22560 12839 22597 12840
rect 22439 12820 22506 12827
rect 22559 12830 22597 12839
rect 20680 12687 20735 12688
rect 20569 12676 20573 12681
rect 20530 12673 20573 12676
rect 20463 12659 20573 12673
rect 19889 12641 20230 12642
rect 18766 12620 18769 12640
rect 18789 12620 19182 12640
rect 19814 12640 20230 12641
rect 20680 12640 20723 12687
rect 19814 12636 20723 12640
rect 19133 12587 19178 12620
rect 19814 12616 19817 12636
rect 19837 12616 20723 12636
rect 20191 12611 20723 12616
rect 20931 12630 20990 12652
rect 20931 12612 20950 12630
rect 20968 12612 20990 12630
rect 19979 12587 20078 12589
rect 19133 12577 20078 12587
rect 17690 12557 17749 12567
rect 17690 12529 17703 12557
rect 17731 12529 17749 12557
rect 19133 12551 20001 12577
rect 19134 12550 20001 12551
rect 19979 12539 20001 12550
rect 20026 12542 20045 12577
rect 20070 12542 20078 12577
rect 20026 12539 20078 12542
rect 20931 12541 20990 12612
rect 22231 12556 22286 12694
rect 22439 12668 22504 12820
rect 22559 12810 22568 12830
rect 22588 12810 22597 12830
rect 22559 12802 22597 12810
rect 22663 12834 22748 12840
rect 22773 12839 22810 12840
rect 22663 12814 22671 12834
rect 22691 12814 22748 12834
rect 22663 12806 22748 12814
rect 22772 12830 22810 12839
rect 22772 12810 22781 12830
rect 22801 12810 22810 12830
rect 22663 12805 22699 12806
rect 22772 12802 22810 12810
rect 22876 12834 22961 12840
rect 22981 12839 23018 12840
rect 22876 12814 22884 12834
rect 22904 12833 22961 12834
rect 22904 12814 22933 12833
rect 22876 12813 22933 12814
rect 22954 12813 22961 12833
rect 22876 12806 22961 12813
rect 22980 12830 23018 12839
rect 22980 12810 22989 12830
rect 23009 12810 23018 12830
rect 22876 12805 22912 12806
rect 22980 12802 23018 12810
rect 23084 12834 23228 12840
rect 23084 12814 23092 12834
rect 23112 12814 23200 12834
rect 23220 12814 23228 12834
rect 23084 12806 23228 12814
rect 23084 12805 23120 12806
rect 23192 12805 23228 12806
rect 23294 12839 23331 12840
rect 23294 12838 23332 12839
rect 23294 12830 23358 12838
rect 23294 12810 23303 12830
rect 23323 12816 23358 12830
rect 23378 12816 23381 12836
rect 23323 12811 23381 12816
rect 23323 12810 23358 12811
rect 22560 12773 22597 12802
rect 22561 12771 22597 12773
rect 22773 12771 22810 12802
rect 22561 12749 22810 12771
rect 22642 12743 22753 12749
rect 22642 12735 22683 12743
rect 22642 12715 22650 12735
rect 22669 12715 22683 12735
rect 22642 12713 22683 12715
rect 22711 12735 22753 12743
rect 22711 12715 22727 12735
rect 22746 12715 22753 12735
rect 22711 12713 22753 12715
rect 22642 12700 22753 12713
rect 22981 12703 23018 12802
rect 23294 12798 23358 12810
rect 22432 12658 22553 12668
rect 22432 12656 22501 12658
rect 22432 12615 22445 12656
rect 22482 12617 22501 12656
rect 22538 12617 22553 12658
rect 22482 12615 22553 12617
rect 22432 12597 22553 12615
rect 22224 12553 22288 12556
rect 22644 12553 22748 12559
rect 22979 12553 23020 12703
rect 23398 12695 23425 12950
rect 23487 12940 23567 12951
rect 23487 12914 23504 12940
rect 23544 12914 23567 12940
rect 23487 12887 23567 12914
rect 23487 12861 23508 12887
rect 23548 12861 23567 12887
rect 23487 12842 23567 12861
rect 23487 12816 23511 12842
rect 23551 12816 23567 12842
rect 23487 12765 23567 12816
rect 22224 12550 23020 12553
rect 23399 12564 23425 12695
rect 23399 12550 23427 12564
rect 19979 12531 20078 12539
rect 20005 12530 20077 12531
rect 17690 12480 17749 12529
rect 19659 12504 19726 12523
rect 19659 12483 19676 12504
rect 17296 12345 17464 12346
rect 17700 12345 17747 12480
rect 17296 12319 17747 12345
rect 17296 12317 17464 12319
rect 17296 12050 17323 12317
rect 17700 12313 17747 12319
rect 19657 12438 19676 12483
rect 19706 12483 19726 12504
rect 19706 12438 19727 12483
rect 20196 12480 20237 12482
rect 20468 12480 20572 12482
rect 20928 12480 20992 12541
rect 17363 12190 17427 12202
rect 17703 12198 17740 12313
rect 17968 12287 18079 12302
rect 17968 12285 18010 12287
rect 17968 12265 17975 12285
rect 17994 12265 18010 12285
rect 17968 12257 18010 12265
rect 18038 12285 18079 12287
rect 18038 12265 18052 12285
rect 18071 12265 18079 12285
rect 18038 12257 18079 12265
rect 17968 12251 18079 12257
rect 17911 12229 18160 12251
rect 19657 12230 19727 12438
rect 19789 12445 20992 12480
rect 22224 12515 23427 12550
rect 23489 12557 23559 12765
rect 24601 12690 24676 12974
rect 24970 12891 25016 12974
rect 25060 12974 25097 13053
rect 25138 13040 25248 13053
rect 25212 12984 25243 12985
rect 25060 12954 25069 12974
rect 25089 12954 25097 12974
rect 25060 12944 25097 12954
rect 25156 12974 25243 12984
rect 25156 12954 25165 12974
rect 25185 12954 25243 12974
rect 25156 12945 25243 12954
rect 25156 12944 25193 12945
rect 25212 12892 25243 12945
rect 25273 12974 25310 13053
rect 25425 12984 25456 12985
rect 25273 12954 25282 12974
rect 25302 12954 25310 12974
rect 25273 12944 25310 12954
rect 25369 12977 25456 12984
rect 25369 12974 25430 12977
rect 25369 12954 25378 12974
rect 25398 12957 25430 12974
rect 25451 12957 25456 12977
rect 25398 12954 25456 12957
rect 25369 12947 25456 12954
rect 25481 12974 25518 13116
rect 25784 13115 25821 13116
rect 25633 12984 25669 12985
rect 25481 12954 25490 12974
rect 25510 12954 25518 12974
rect 25369 12945 25425 12947
rect 25369 12944 25406 12945
rect 25481 12944 25518 12954
rect 25577 12974 25725 12984
rect 25825 12981 25921 12983
rect 25577 12954 25586 12974
rect 25606 12954 25696 12974
rect 25716 12954 25725 12974
rect 25577 12948 25725 12954
rect 25577 12945 25641 12948
rect 25577 12944 25614 12945
rect 25633 12918 25641 12945
rect 25662 12945 25725 12948
rect 25783 12974 25921 12981
rect 25783 12954 25792 12974
rect 25812 12954 25921 12974
rect 25783 12945 25921 12954
rect 25662 12918 25669 12945
rect 25688 12944 25725 12945
rect 25784 12944 25821 12945
rect 25633 12893 25669 12918
rect 25104 12891 25145 12892
rect 24970 12884 25145 12891
rect 24768 12858 24854 12877
rect 24768 12817 24783 12858
rect 24837 12817 24854 12858
rect 24970 12864 25114 12884
rect 25134 12864 25145 12884
rect 24970 12856 25145 12864
rect 25212 12888 25571 12892
rect 25212 12883 25534 12888
rect 25212 12859 25325 12883
rect 25349 12864 25534 12883
rect 25558 12864 25571 12888
rect 25349 12859 25571 12864
rect 25212 12856 25571 12859
rect 25633 12856 25668 12893
rect 25736 12890 25836 12893
rect 25736 12886 25803 12890
rect 25736 12860 25748 12886
rect 25774 12864 25803 12886
rect 25829 12864 25836 12890
rect 25774 12860 25836 12864
rect 25736 12856 25836 12860
rect 24970 12852 25016 12856
rect 25212 12835 25243 12856
rect 25633 12835 25669 12856
rect 25055 12834 25092 12835
rect 24768 12781 24854 12817
rect 25054 12825 25092 12834
rect 25054 12805 25063 12825
rect 25083 12805 25092 12825
rect 25054 12797 25092 12805
rect 25158 12829 25243 12835
rect 25268 12834 25305 12835
rect 25158 12809 25166 12829
rect 25186 12809 25243 12829
rect 25158 12801 25243 12809
rect 25267 12825 25305 12834
rect 25267 12805 25276 12825
rect 25296 12805 25305 12825
rect 25158 12800 25194 12801
rect 25267 12797 25305 12805
rect 25371 12829 25456 12835
rect 25476 12834 25513 12835
rect 25371 12809 25379 12829
rect 25399 12828 25456 12829
rect 25399 12809 25428 12828
rect 25371 12808 25428 12809
rect 25449 12808 25456 12828
rect 25371 12801 25456 12808
rect 25475 12825 25513 12834
rect 25475 12805 25484 12825
rect 25504 12805 25513 12825
rect 25371 12800 25407 12801
rect 25475 12797 25513 12805
rect 25579 12829 25723 12835
rect 25579 12809 25587 12829
rect 25607 12809 25695 12829
rect 25715 12809 25723 12829
rect 25579 12801 25723 12809
rect 25579 12800 25615 12801
rect 22224 12454 22288 12515
rect 22644 12513 22748 12515
rect 22979 12513 23020 12515
rect 23489 12512 23510 12557
rect 23490 12491 23510 12512
rect 23540 12512 23559 12557
rect 24596 12648 24676 12690
rect 23540 12491 23557 12512
rect 23490 12472 23557 12491
rect 23139 12464 23211 12465
rect 23138 12456 23237 12464
rect 19789 12431 19817 12445
rect 19791 12300 19817 12431
rect 20196 12442 20992 12445
rect 17911 12198 17948 12229
rect 18124 12227 18160 12229
rect 18124 12198 18161 12227
rect 17363 12189 17398 12190
rect 17340 12184 17398 12189
rect 17340 12164 17343 12184
rect 17363 12170 17398 12184
rect 17418 12170 17427 12190
rect 17363 12162 17427 12170
rect 17389 12161 17427 12162
rect 17390 12160 17427 12161
rect 17493 12194 17529 12195
rect 17601 12194 17637 12195
rect 17493 12186 17637 12194
rect 17493 12166 17501 12186
rect 17521 12166 17609 12186
rect 17629 12166 17637 12186
rect 17493 12160 17637 12166
rect 17703 12190 17741 12198
rect 17809 12194 17845 12195
rect 17703 12170 17712 12190
rect 17732 12170 17741 12190
rect 17703 12161 17741 12170
rect 17760 12187 17845 12194
rect 17760 12167 17767 12187
rect 17788 12186 17845 12187
rect 17788 12167 17817 12186
rect 17760 12166 17817 12167
rect 17837 12166 17845 12186
rect 17703 12160 17740 12161
rect 17760 12160 17845 12166
rect 17911 12190 17949 12198
rect 18022 12194 18058 12195
rect 17911 12170 17920 12190
rect 17940 12170 17949 12190
rect 17911 12161 17949 12170
rect 17973 12186 18058 12194
rect 17973 12166 18030 12186
rect 18050 12166 18058 12186
rect 17911 12160 17948 12161
rect 17973 12160 18058 12166
rect 18124 12190 18162 12198
rect 18124 12170 18133 12190
rect 18153 12170 18162 12190
rect 18124 12161 18162 12170
rect 19649 12179 19729 12230
rect 18124 12160 18161 12161
rect 17547 12139 17583 12160
rect 17973 12139 18004 12160
rect 18184 12145 18241 12153
rect 18184 12139 18192 12145
rect 17380 12135 17480 12139
rect 17380 12131 17442 12135
rect 17380 12105 17387 12131
rect 17413 12109 17442 12131
rect 17468 12109 17480 12135
rect 17413 12105 17480 12109
rect 17380 12102 17480 12105
rect 17548 12102 17583 12139
rect 17645 12136 18004 12139
rect 17645 12131 17867 12136
rect 17645 12107 17658 12131
rect 17682 12112 17867 12131
rect 17891 12112 18004 12136
rect 17682 12107 18004 12112
rect 17645 12103 18004 12107
rect 18071 12131 18192 12139
rect 18071 12111 18082 12131
rect 18102 12122 18192 12131
rect 18218 12122 18241 12145
rect 18102 12111 18241 12122
rect 18071 12109 18241 12111
rect 18544 12138 18616 12158
rect 18544 12115 18572 12138
rect 18598 12115 18616 12138
rect 18071 12104 18192 12109
rect 18071 12103 18112 12104
rect 17547 12077 17583 12102
rect 17395 12050 17432 12051
rect 17491 12050 17528 12051
rect 17547 12050 17554 12077
rect 17295 12041 17433 12050
rect 17295 12021 17404 12041
rect 17424 12021 17433 12041
rect 17295 12014 17433 12021
rect 17491 12047 17554 12050
rect 17575 12050 17583 12077
rect 17602 12050 17639 12051
rect 17575 12047 17639 12050
rect 17491 12041 17639 12047
rect 17491 12021 17500 12041
rect 17520 12021 17610 12041
rect 17630 12021 17639 12041
rect 17295 12012 17391 12014
rect 17491 12011 17639 12021
rect 17698 12041 17735 12051
rect 17810 12050 17847 12051
rect 17791 12048 17847 12050
rect 17698 12021 17706 12041
rect 17726 12021 17735 12041
rect 17547 12010 17583 12011
rect 17395 11879 17432 11880
rect 17698 11879 17735 12021
rect 17760 12041 17847 12048
rect 17760 12038 17818 12041
rect 17760 12018 17765 12038
rect 17786 12021 17818 12038
rect 17838 12021 17847 12041
rect 17786 12018 17847 12021
rect 17760 12011 17847 12018
rect 17906 12041 17943 12051
rect 17906 12021 17914 12041
rect 17934 12021 17943 12041
rect 17760 12010 17791 12011
rect 17906 11942 17943 12021
rect 17973 12050 18004 12103
rect 18544 12053 18616 12115
rect 19649 12153 19665 12179
rect 19705 12153 19729 12179
rect 19649 12134 19729 12153
rect 19649 12108 19668 12134
rect 19708 12108 19729 12134
rect 19649 12081 19729 12108
rect 19649 12055 19672 12081
rect 19712 12055 19729 12081
rect 18023 12050 18060 12051
rect 17973 12041 18060 12050
rect 17973 12021 18031 12041
rect 18051 12021 18060 12041
rect 17973 12011 18060 12021
rect 18119 12041 18156 12051
rect 18119 12021 18127 12041
rect 18147 12021 18156 12041
rect 17973 12010 18004 12011
rect 17968 11942 18078 11955
rect 18119 11942 18156 12021
rect 17906 11940 18156 11942
rect 17906 11937 18007 11940
rect 17906 11918 17971 11937
rect 17968 11910 17971 11918
rect 18000 11910 18007 11937
rect 18035 11913 18045 11940
rect 18074 11918 18156 11940
rect 18074 11913 18078 11918
rect 18035 11910 18078 11913
rect 17968 11896 18078 11910
rect 17394 11878 17735 11879
rect 17319 11873 17735 11878
rect 17319 11853 17322 11873
rect 17342 11853 17736 11873
rect 17545 11820 17582 11830
rect 17545 11783 17554 11820
rect 17571 11783 17582 11820
rect 17545 11762 17582 11783
rect 17254 10823 17422 10824
rect 17551 10823 17580 11762
rect 17693 11148 17736 11853
rect 18548 11502 18610 12053
rect 19649 12044 19729 12055
rect 19791 12045 19818 12300
rect 20196 12292 20237 12442
rect 20468 12436 20572 12442
rect 20928 12439 20992 12442
rect 20663 12380 20784 12398
rect 20663 12378 20734 12380
rect 20663 12337 20678 12378
rect 20715 12339 20734 12378
rect 20771 12339 20784 12380
rect 20715 12337 20784 12339
rect 20663 12327 20784 12337
rect 19858 12185 19922 12197
rect 20198 12193 20235 12292
rect 20463 12282 20574 12295
rect 20463 12280 20505 12282
rect 20463 12260 20470 12280
rect 20489 12260 20505 12280
rect 20463 12252 20505 12260
rect 20533 12280 20574 12282
rect 20533 12260 20547 12280
rect 20566 12260 20574 12280
rect 20533 12252 20574 12260
rect 20463 12246 20574 12252
rect 20406 12224 20655 12246
rect 20406 12193 20443 12224
rect 20619 12222 20655 12224
rect 20619 12193 20656 12222
rect 19858 12184 19893 12185
rect 19835 12179 19893 12184
rect 19835 12159 19838 12179
rect 19858 12165 19893 12179
rect 19913 12165 19922 12185
rect 19858 12157 19922 12165
rect 19884 12156 19922 12157
rect 19885 12155 19922 12156
rect 19988 12189 20024 12190
rect 20096 12189 20132 12190
rect 19988 12181 20132 12189
rect 19988 12161 19996 12181
rect 20016 12161 20104 12181
rect 20124 12161 20132 12181
rect 19988 12155 20132 12161
rect 20198 12185 20236 12193
rect 20304 12189 20340 12190
rect 20198 12165 20207 12185
rect 20227 12165 20236 12185
rect 20198 12156 20236 12165
rect 20255 12182 20340 12189
rect 20255 12162 20262 12182
rect 20283 12181 20340 12182
rect 20283 12162 20312 12181
rect 20255 12161 20312 12162
rect 20332 12161 20340 12181
rect 20198 12155 20235 12156
rect 20255 12155 20340 12161
rect 20406 12185 20444 12193
rect 20517 12189 20553 12190
rect 20406 12165 20415 12185
rect 20435 12165 20444 12185
rect 20406 12156 20444 12165
rect 20468 12181 20553 12189
rect 20468 12161 20525 12181
rect 20545 12161 20553 12181
rect 20406 12155 20443 12156
rect 20468 12155 20553 12161
rect 20619 12185 20657 12193
rect 20619 12165 20628 12185
rect 20648 12165 20657 12185
rect 20712 12175 20777 12327
rect 20930 12301 20985 12439
rect 22226 12383 22285 12454
rect 23138 12453 23190 12456
rect 23138 12418 23146 12453
rect 23171 12418 23190 12453
rect 23215 12445 23237 12456
rect 23215 12444 24082 12445
rect 23215 12418 24083 12444
rect 23138 12408 24083 12418
rect 23138 12406 23237 12408
rect 22226 12365 22248 12383
rect 22266 12365 22285 12383
rect 22226 12343 22285 12365
rect 22493 12379 23025 12384
rect 22493 12359 23379 12379
rect 23399 12359 23402 12379
rect 24038 12375 24083 12408
rect 22493 12355 23402 12359
rect 22493 12308 22536 12355
rect 22986 12354 23402 12355
rect 24034 12355 24427 12375
rect 24447 12355 24450 12375
rect 22986 12353 23327 12354
rect 22643 12322 22753 12336
rect 22643 12319 22686 12322
rect 22643 12314 22647 12319
rect 22481 12307 22536 12308
rect 20619 12156 20657 12165
rect 20710 12168 20777 12175
rect 20619 12155 20656 12156
rect 20042 12134 20078 12155
rect 20468 12134 20499 12155
rect 20710 12147 20727 12168
rect 20763 12147 20777 12168
rect 20929 12188 20985 12301
rect 20929 12170 20948 12188
rect 20966 12170 20985 12188
rect 20929 12150 20985 12170
rect 22225 12284 22536 12307
rect 22225 12266 22250 12284
rect 22268 12272 22536 12284
rect 22565 12292 22647 12314
rect 22676 12292 22686 12319
rect 22714 12295 22721 12322
rect 22750 12314 22753 12322
rect 22750 12295 22815 12314
rect 22714 12292 22815 12295
rect 22565 12290 22815 12292
rect 22268 12266 22290 12272
rect 20710 12134 20777 12147
rect 19875 12130 19975 12134
rect 19875 12126 19937 12130
rect 19875 12100 19882 12126
rect 19908 12104 19937 12126
rect 19963 12104 19975 12130
rect 19908 12100 19975 12104
rect 19875 12097 19975 12100
rect 20043 12097 20078 12134
rect 20140 12131 20499 12134
rect 20140 12126 20362 12131
rect 20140 12102 20153 12126
rect 20177 12107 20362 12126
rect 20386 12107 20499 12131
rect 20177 12102 20499 12107
rect 20140 12098 20499 12102
rect 20566 12128 20777 12134
rect 20566 12126 20727 12128
rect 20566 12106 20577 12126
rect 20597 12106 20727 12126
rect 20566 12099 20727 12106
rect 20566 12098 20607 12099
rect 20042 12072 20078 12097
rect 19890 12045 19927 12046
rect 19986 12045 20023 12046
rect 20042 12045 20049 12072
rect 19790 12036 19928 12045
rect 19790 12016 19899 12036
rect 19919 12016 19928 12036
rect 19790 12009 19928 12016
rect 19986 12042 20049 12045
rect 20070 12045 20078 12072
rect 20097 12045 20134 12046
rect 20070 12042 20134 12045
rect 19986 12036 20134 12042
rect 19986 12016 19995 12036
rect 20015 12016 20105 12036
rect 20125 12016 20134 12036
rect 19790 12007 19886 12009
rect 19986 12006 20134 12016
rect 20193 12036 20230 12046
rect 20305 12045 20342 12046
rect 20286 12043 20342 12045
rect 20193 12016 20201 12036
rect 20221 12016 20230 12036
rect 20042 12005 20078 12006
rect 19890 11874 19927 11875
rect 20193 11874 20230 12016
rect 20255 12036 20342 12043
rect 20255 12033 20313 12036
rect 20255 12013 20260 12033
rect 20281 12016 20313 12033
rect 20333 12016 20342 12036
rect 20281 12013 20342 12016
rect 20255 12006 20342 12013
rect 20401 12036 20438 12046
rect 20401 12016 20409 12036
rect 20429 12016 20438 12036
rect 20255 12005 20286 12006
rect 20401 11937 20438 12016
rect 20468 12045 20499 12098
rect 20712 12091 20727 12099
rect 20767 12091 20777 12128
rect 22225 12127 22290 12266
rect 22565 12211 22602 12290
rect 22643 12277 22753 12290
rect 22717 12221 22748 12222
rect 22565 12191 22574 12211
rect 22594 12191 22602 12211
rect 20712 12082 20777 12091
rect 20925 12089 20990 12110
rect 22225 12109 22248 12127
rect 22266 12109 22290 12127
rect 22225 12092 22290 12109
rect 22445 12173 22513 12186
rect 22565 12181 22602 12191
rect 22661 12211 22748 12221
rect 22661 12191 22670 12211
rect 22690 12191 22748 12211
rect 22661 12182 22748 12191
rect 22661 12181 22698 12182
rect 22445 12131 22452 12173
rect 22501 12131 22513 12173
rect 22445 12128 22513 12131
rect 22717 12129 22748 12182
rect 22778 12211 22815 12290
rect 22930 12221 22961 12222
rect 22778 12191 22787 12211
rect 22807 12191 22815 12211
rect 22778 12181 22815 12191
rect 22874 12214 22961 12221
rect 22874 12211 22935 12214
rect 22874 12191 22883 12211
rect 22903 12194 22935 12211
rect 22956 12194 22961 12214
rect 22903 12191 22961 12194
rect 22874 12184 22961 12191
rect 22986 12211 23023 12353
rect 23289 12352 23326 12353
rect 24034 12350 24450 12355
rect 24034 12349 24375 12350
rect 23691 12318 23801 12332
rect 23691 12315 23734 12318
rect 23691 12310 23695 12315
rect 23613 12288 23695 12310
rect 23724 12288 23734 12315
rect 23762 12291 23769 12318
rect 23798 12310 23801 12318
rect 23798 12291 23863 12310
rect 23762 12288 23863 12291
rect 23613 12286 23863 12288
rect 23138 12221 23174 12222
rect 22986 12191 22995 12211
rect 23015 12191 23023 12211
rect 22874 12182 22930 12184
rect 22874 12181 22911 12182
rect 22986 12181 23023 12191
rect 23082 12211 23230 12221
rect 23330 12218 23426 12220
rect 23082 12191 23091 12211
rect 23111 12191 23201 12211
rect 23221 12191 23230 12211
rect 23082 12185 23230 12191
rect 23082 12182 23146 12185
rect 23082 12181 23119 12182
rect 23138 12155 23146 12182
rect 23167 12182 23230 12185
rect 23288 12211 23426 12218
rect 23288 12191 23297 12211
rect 23317 12191 23426 12211
rect 23288 12182 23426 12191
rect 23613 12207 23650 12286
rect 23691 12273 23801 12286
rect 23765 12217 23796 12218
rect 23613 12187 23622 12207
rect 23642 12187 23650 12207
rect 23167 12155 23174 12182
rect 23193 12181 23230 12182
rect 23289 12181 23326 12182
rect 23138 12130 23174 12155
rect 22609 12128 22650 12129
rect 22445 12121 22650 12128
rect 22445 12110 22619 12121
rect 20925 12071 20950 12089
rect 20968 12071 20990 12089
rect 22445 12077 22453 12110
rect 20518 12045 20555 12046
rect 20468 12036 20555 12045
rect 20468 12016 20526 12036
rect 20546 12016 20555 12036
rect 20468 12006 20555 12016
rect 20614 12036 20651 12046
rect 20614 12016 20622 12036
rect 20642 12016 20651 12036
rect 20468 12005 20499 12006
rect 20463 11937 20573 11950
rect 20614 11937 20651 12016
rect 20925 11995 20990 12071
rect 22446 12068 22453 12077
rect 22502 12101 22619 12110
rect 22639 12101 22650 12121
rect 22502 12093 22650 12101
rect 22717 12125 23076 12129
rect 22717 12120 23039 12125
rect 22717 12096 22830 12120
rect 22854 12101 23039 12120
rect 23063 12101 23076 12125
rect 22854 12096 23076 12101
rect 22717 12093 23076 12096
rect 23138 12093 23173 12130
rect 23241 12127 23341 12130
rect 23241 12123 23308 12127
rect 23241 12097 23253 12123
rect 23279 12101 23308 12123
rect 23334 12101 23341 12127
rect 23279 12097 23341 12101
rect 23241 12093 23341 12097
rect 22502 12077 22513 12093
rect 22502 12068 22510 12077
rect 22717 12072 22748 12093
rect 23138 12072 23174 12093
rect 22560 12071 22597 12072
rect 22225 12028 22290 12047
rect 22225 12010 22250 12028
rect 22268 12010 22290 12028
rect 20401 11935 20651 11937
rect 20401 11932 20502 11935
rect 20401 11913 20466 11932
rect 20463 11905 20466 11913
rect 20495 11905 20502 11932
rect 20530 11908 20540 11935
rect 20569 11913 20651 11935
rect 20674 11960 20991 11995
rect 20569 11908 20573 11913
rect 20530 11905 20573 11908
rect 20463 11891 20573 11905
rect 19889 11873 20230 11874
rect 19814 11871 20230 11873
rect 20674 11871 20714 11960
rect 20925 11933 20990 11960
rect 20925 11915 20948 11933
rect 20966 11915 20990 11933
rect 20925 11895 20990 11915
rect 19811 11868 20714 11871
rect 19811 11848 19817 11868
rect 19837 11848 20714 11868
rect 19811 11844 20714 11848
rect 20674 11841 20714 11844
rect 20926 11834 20991 11855
rect 19144 11826 19805 11827
rect 19144 11819 20078 11826
rect 19144 11818 20050 11819
rect 19144 11798 19995 11818
rect 20027 11799 20050 11818
rect 20075 11799 20078 11819
rect 20027 11798 20078 11799
rect 19144 11791 20078 11798
rect 18743 11749 18911 11750
rect 19146 11749 19185 11791
rect 19974 11789 20078 11791
rect 20043 11787 20078 11789
rect 20926 11816 20950 11834
rect 20968 11816 20991 11834
rect 20926 11769 20991 11816
rect 18743 11723 19187 11749
rect 18743 11721 18911 11723
rect 18545 11418 18614 11502
rect 17694 11140 17736 11148
rect 17694 11129 17739 11140
rect 17694 11091 17704 11129
rect 17729 11091 17739 11129
rect 17694 11082 17739 11091
rect 18543 10939 18614 11418
rect 18743 11370 18770 11721
rect 19146 11717 19187 11723
rect 18810 11510 18874 11522
rect 19150 11518 19187 11717
rect 19649 11744 19721 11761
rect 19649 11705 19657 11744
rect 19702 11705 19721 11744
rect 19415 11607 19526 11622
rect 19415 11605 19457 11607
rect 19415 11585 19422 11605
rect 19441 11585 19457 11605
rect 19415 11577 19457 11585
rect 19485 11605 19526 11607
rect 19485 11585 19499 11605
rect 19518 11585 19526 11605
rect 19485 11577 19526 11585
rect 19415 11571 19526 11577
rect 19358 11549 19607 11571
rect 19358 11518 19395 11549
rect 19571 11547 19607 11549
rect 19571 11518 19608 11547
rect 18810 11509 18845 11510
rect 18787 11504 18845 11509
rect 18787 11484 18790 11504
rect 18810 11490 18845 11504
rect 18865 11490 18874 11510
rect 18810 11482 18874 11490
rect 18836 11481 18874 11482
rect 18837 11480 18874 11481
rect 18940 11514 18976 11515
rect 19048 11514 19084 11515
rect 18940 11506 19084 11514
rect 18940 11486 18948 11506
rect 18968 11486 19056 11506
rect 19076 11486 19084 11506
rect 18940 11480 19084 11486
rect 19150 11510 19188 11518
rect 19256 11514 19292 11515
rect 19150 11490 19159 11510
rect 19179 11490 19188 11510
rect 19150 11481 19188 11490
rect 19207 11507 19292 11514
rect 19207 11487 19214 11507
rect 19235 11506 19292 11507
rect 19235 11487 19264 11506
rect 19207 11486 19264 11487
rect 19284 11486 19292 11506
rect 19150 11480 19187 11481
rect 19207 11480 19292 11486
rect 19358 11510 19396 11518
rect 19469 11514 19505 11515
rect 19358 11490 19367 11510
rect 19387 11490 19396 11510
rect 19358 11481 19396 11490
rect 19420 11506 19505 11514
rect 19420 11486 19477 11506
rect 19497 11486 19505 11506
rect 19358 11480 19395 11481
rect 19420 11480 19505 11486
rect 19571 11510 19609 11518
rect 19571 11490 19580 11510
rect 19600 11490 19609 11510
rect 19571 11481 19609 11490
rect 19649 11495 19721 11705
rect 19791 11739 20991 11769
rect 19791 11738 20235 11739
rect 19791 11736 19959 11738
rect 19649 11481 19732 11495
rect 19571 11480 19608 11481
rect 18994 11459 19030 11480
rect 19420 11459 19451 11480
rect 19649 11459 19666 11481
rect 18827 11455 18927 11459
rect 18827 11451 18889 11455
rect 18827 11425 18834 11451
rect 18860 11429 18889 11451
rect 18915 11429 18927 11455
rect 18860 11425 18927 11429
rect 18827 11422 18927 11425
rect 18995 11422 19030 11459
rect 19092 11456 19451 11459
rect 19092 11451 19314 11456
rect 19092 11427 19105 11451
rect 19129 11432 19314 11451
rect 19338 11432 19451 11456
rect 19129 11427 19451 11432
rect 19092 11423 19451 11427
rect 19518 11451 19666 11459
rect 19518 11431 19529 11451
rect 19549 11448 19666 11451
rect 19719 11448 19732 11481
rect 19549 11431 19732 11448
rect 19518 11424 19732 11431
rect 19518 11423 19559 11424
rect 19649 11423 19732 11424
rect 18994 11397 19030 11422
rect 18842 11370 18879 11371
rect 18938 11370 18975 11371
rect 18994 11370 19001 11397
rect 18742 11361 18880 11370
rect 18742 11341 18851 11361
rect 18871 11341 18880 11361
rect 18742 11334 18880 11341
rect 18938 11367 19001 11370
rect 19022 11370 19030 11397
rect 19049 11370 19086 11371
rect 19022 11367 19086 11370
rect 18938 11361 19086 11367
rect 18938 11341 18947 11361
rect 18967 11341 19057 11361
rect 19077 11341 19086 11361
rect 18742 11332 18838 11334
rect 18938 11331 19086 11341
rect 19145 11361 19182 11371
rect 19257 11370 19294 11371
rect 19238 11368 19294 11370
rect 19145 11341 19153 11361
rect 19173 11341 19182 11361
rect 18994 11330 19030 11331
rect 18842 11199 18879 11200
rect 19145 11199 19182 11341
rect 19207 11361 19294 11368
rect 19207 11358 19265 11361
rect 19207 11338 19212 11358
rect 19233 11341 19265 11358
rect 19285 11341 19294 11361
rect 19233 11338 19294 11341
rect 19207 11331 19294 11338
rect 19353 11361 19390 11371
rect 19353 11341 19361 11361
rect 19381 11341 19390 11361
rect 19207 11330 19238 11331
rect 19353 11262 19390 11341
rect 19420 11370 19451 11423
rect 19657 11390 19671 11423
rect 19724 11390 19732 11423
rect 19657 11384 19732 11390
rect 19657 11379 19727 11384
rect 19470 11370 19507 11371
rect 19420 11361 19507 11370
rect 19420 11341 19478 11361
rect 19498 11341 19507 11361
rect 19420 11331 19507 11341
rect 19566 11361 19603 11371
rect 19791 11366 19818 11736
rect 19858 11506 19922 11518
rect 20198 11514 20235 11738
rect 20706 11719 20770 11721
rect 20702 11707 20770 11719
rect 20702 11674 20713 11707
rect 20753 11674 20770 11707
rect 20702 11664 20770 11674
rect 20463 11603 20574 11618
rect 20463 11601 20505 11603
rect 20463 11581 20470 11601
rect 20489 11581 20505 11601
rect 20463 11573 20505 11581
rect 20533 11601 20574 11603
rect 20533 11581 20547 11601
rect 20566 11581 20574 11601
rect 20533 11573 20574 11581
rect 20463 11567 20574 11573
rect 20406 11545 20655 11567
rect 20406 11514 20443 11545
rect 20619 11543 20655 11545
rect 20619 11514 20656 11543
rect 19858 11505 19893 11506
rect 19835 11500 19893 11505
rect 19835 11480 19838 11500
rect 19858 11486 19893 11500
rect 19913 11486 19922 11506
rect 19858 11478 19922 11486
rect 19884 11477 19922 11478
rect 19885 11476 19922 11477
rect 19988 11510 20024 11511
rect 20096 11510 20132 11511
rect 19988 11502 20132 11510
rect 19988 11482 19996 11502
rect 20016 11482 20104 11502
rect 20124 11482 20132 11502
rect 19988 11476 20132 11482
rect 20198 11506 20236 11514
rect 20304 11510 20340 11511
rect 20198 11486 20207 11506
rect 20227 11486 20236 11506
rect 20198 11477 20236 11486
rect 20255 11503 20340 11510
rect 20255 11483 20262 11503
rect 20283 11502 20340 11503
rect 20283 11483 20312 11502
rect 20255 11482 20312 11483
rect 20332 11482 20340 11502
rect 20198 11476 20235 11477
rect 20255 11476 20340 11482
rect 20406 11506 20444 11514
rect 20517 11510 20553 11511
rect 20406 11486 20415 11506
rect 20435 11486 20444 11506
rect 20406 11477 20444 11486
rect 20468 11502 20553 11510
rect 20468 11482 20525 11502
rect 20545 11482 20553 11502
rect 20406 11476 20443 11477
rect 20468 11476 20553 11482
rect 20619 11506 20657 11514
rect 20619 11486 20628 11506
rect 20648 11486 20657 11506
rect 20619 11477 20657 11486
rect 20706 11480 20770 11664
rect 20926 11538 20991 11739
rect 22225 11809 22290 12010
rect 22446 11884 22510 12068
rect 22559 12062 22597 12071
rect 22559 12042 22568 12062
rect 22588 12042 22597 12062
rect 22559 12034 22597 12042
rect 22663 12066 22748 12072
rect 22773 12071 22810 12072
rect 22663 12046 22671 12066
rect 22691 12046 22748 12066
rect 22663 12038 22748 12046
rect 22772 12062 22810 12071
rect 22772 12042 22781 12062
rect 22801 12042 22810 12062
rect 22663 12037 22699 12038
rect 22772 12034 22810 12042
rect 22876 12066 22961 12072
rect 22981 12071 23018 12072
rect 22876 12046 22884 12066
rect 22904 12065 22961 12066
rect 22904 12046 22933 12065
rect 22876 12045 22933 12046
rect 22954 12045 22961 12065
rect 22876 12038 22961 12045
rect 22980 12062 23018 12071
rect 22980 12042 22989 12062
rect 23009 12042 23018 12062
rect 22876 12037 22912 12038
rect 22980 12034 23018 12042
rect 23084 12066 23228 12072
rect 23084 12046 23092 12066
rect 23112 12046 23200 12066
rect 23220 12046 23228 12066
rect 23084 12038 23228 12046
rect 23084 12037 23120 12038
rect 23192 12037 23228 12038
rect 23294 12071 23331 12072
rect 23294 12070 23332 12071
rect 23294 12062 23358 12070
rect 23294 12042 23303 12062
rect 23323 12048 23358 12062
rect 23378 12048 23381 12068
rect 23323 12043 23381 12048
rect 23323 12042 23358 12043
rect 22560 12005 22597 12034
rect 22561 12003 22597 12005
rect 22773 12003 22810 12034
rect 22561 11981 22810 12003
rect 22642 11975 22753 11981
rect 22642 11967 22683 11975
rect 22642 11947 22650 11967
rect 22669 11947 22683 11967
rect 22642 11945 22683 11947
rect 22711 11967 22753 11975
rect 22711 11947 22727 11967
rect 22746 11947 22753 11967
rect 22711 11945 22753 11947
rect 22642 11930 22753 11945
rect 22446 11874 22514 11884
rect 22446 11841 22463 11874
rect 22503 11841 22514 11874
rect 22446 11829 22514 11841
rect 22446 11827 22510 11829
rect 22981 11810 23018 12034
rect 23294 12030 23358 12042
rect 23398 11812 23425 12182
rect 23613 12177 23650 12187
rect 23709 12207 23796 12217
rect 23709 12187 23718 12207
rect 23738 12187 23796 12207
rect 23709 12178 23796 12187
rect 23709 12177 23746 12178
rect 23489 12164 23559 12169
rect 23484 12158 23559 12164
rect 23484 12125 23492 12158
rect 23545 12125 23559 12158
rect 23765 12125 23796 12178
rect 23826 12207 23863 12286
rect 23978 12217 24009 12218
rect 23826 12187 23835 12207
rect 23855 12187 23863 12207
rect 23826 12177 23863 12187
rect 23922 12210 24009 12217
rect 23922 12207 23983 12210
rect 23922 12187 23931 12207
rect 23951 12190 23983 12207
rect 24004 12190 24009 12210
rect 23951 12187 24009 12190
rect 23922 12180 24009 12187
rect 24034 12207 24071 12349
rect 24337 12348 24374 12349
rect 24186 12217 24222 12218
rect 24034 12187 24043 12207
rect 24063 12187 24071 12207
rect 23922 12178 23978 12180
rect 23922 12177 23959 12178
rect 24034 12177 24071 12187
rect 24130 12207 24278 12217
rect 24378 12214 24474 12216
rect 24130 12187 24139 12207
rect 24159 12187 24249 12207
rect 24269 12187 24278 12207
rect 24130 12181 24278 12187
rect 24130 12178 24194 12181
rect 24130 12177 24167 12178
rect 24186 12151 24194 12178
rect 24215 12178 24278 12181
rect 24336 12207 24474 12214
rect 24336 12187 24345 12207
rect 24365 12187 24474 12207
rect 24336 12178 24474 12187
rect 24215 12151 24222 12178
rect 24241 12177 24278 12178
rect 24337 12177 24374 12178
rect 24186 12126 24222 12151
rect 23484 12124 23567 12125
rect 23657 12124 23698 12125
rect 23484 12117 23698 12124
rect 23484 12100 23667 12117
rect 23484 12067 23497 12100
rect 23550 12097 23667 12100
rect 23687 12097 23698 12117
rect 23550 12089 23698 12097
rect 23765 12121 24124 12125
rect 23765 12116 24087 12121
rect 23765 12092 23878 12116
rect 23902 12097 24087 12116
rect 24111 12097 24124 12121
rect 23902 12092 24124 12097
rect 23765 12089 24124 12092
rect 24186 12089 24221 12126
rect 24289 12123 24389 12126
rect 24289 12119 24356 12123
rect 24289 12093 24301 12119
rect 24327 12097 24356 12119
rect 24382 12097 24389 12123
rect 24327 12093 24389 12097
rect 24289 12089 24389 12093
rect 23550 12067 23567 12089
rect 23765 12068 23796 12089
rect 24186 12068 24222 12089
rect 23608 12067 23645 12068
rect 23484 12053 23567 12067
rect 23257 11810 23425 11812
rect 22981 11809 23425 11810
rect 22225 11779 23425 11809
rect 23495 11843 23567 12053
rect 23607 12058 23645 12067
rect 23607 12038 23616 12058
rect 23636 12038 23645 12058
rect 23607 12030 23645 12038
rect 23711 12062 23796 12068
rect 23821 12067 23858 12068
rect 23711 12042 23719 12062
rect 23739 12042 23796 12062
rect 23711 12034 23796 12042
rect 23820 12058 23858 12067
rect 23820 12038 23829 12058
rect 23849 12038 23858 12058
rect 23711 12033 23747 12034
rect 23820 12030 23858 12038
rect 23924 12062 24009 12068
rect 24029 12067 24066 12068
rect 23924 12042 23932 12062
rect 23952 12061 24009 12062
rect 23952 12042 23981 12061
rect 23924 12041 23981 12042
rect 24002 12041 24009 12061
rect 23924 12034 24009 12041
rect 24028 12058 24066 12067
rect 24028 12038 24037 12058
rect 24057 12038 24066 12058
rect 23924 12033 23960 12034
rect 24028 12030 24066 12038
rect 24132 12062 24276 12068
rect 24132 12042 24140 12062
rect 24160 12042 24248 12062
rect 24268 12042 24276 12062
rect 24132 12034 24276 12042
rect 24132 12033 24168 12034
rect 24240 12033 24276 12034
rect 24342 12067 24379 12068
rect 24342 12066 24380 12067
rect 24342 12058 24406 12066
rect 24342 12038 24351 12058
rect 24371 12044 24406 12058
rect 24426 12044 24429 12064
rect 24371 12039 24429 12044
rect 24371 12038 24406 12039
rect 23608 12001 23645 12030
rect 23609 11999 23645 12001
rect 23821 11999 23858 12030
rect 23609 11977 23858 11999
rect 23690 11971 23801 11977
rect 23690 11963 23731 11971
rect 23690 11943 23698 11963
rect 23717 11943 23731 11963
rect 23690 11941 23731 11943
rect 23759 11963 23801 11971
rect 23759 11943 23775 11963
rect 23794 11943 23801 11963
rect 23759 11941 23801 11943
rect 23690 11926 23801 11941
rect 23495 11804 23514 11843
rect 23559 11804 23567 11843
rect 23495 11787 23567 11804
rect 24029 11831 24066 12030
rect 24342 12026 24406 12038
rect 24029 11825 24070 11831
rect 24446 11827 24473 12178
rect 24596 12048 24675 12648
rect 24772 12196 24851 12781
rect 25055 12768 25092 12797
rect 25056 12766 25092 12768
rect 25268 12766 25305 12797
rect 25056 12744 25305 12766
rect 25137 12738 25248 12744
rect 25137 12730 25178 12738
rect 25137 12710 25145 12730
rect 25164 12710 25178 12730
rect 25137 12708 25178 12710
rect 25206 12730 25248 12738
rect 25206 12710 25222 12730
rect 25241 12710 25248 12730
rect 25206 12708 25248 12710
rect 25137 12693 25248 12708
rect 25476 12682 25513 12797
rect 25469 12570 25516 12682
rect 25637 12642 25667 12801
rect 25687 12800 25723 12801
rect 25789 12834 25826 12835
rect 25789 12833 25827 12834
rect 25789 12825 25853 12833
rect 25789 12805 25798 12825
rect 25818 12811 25853 12825
rect 25873 12811 25876 12831
rect 25818 12806 25876 12811
rect 25818 12805 25853 12806
rect 25789 12793 25853 12805
rect 25637 12638 25723 12642
rect 25637 12620 25652 12638
rect 25704 12620 25723 12638
rect 25637 12611 25723 12620
rect 25893 12572 25920 12945
rect 25752 12570 25920 12572
rect 25469 12544 25920 12570
rect 25469 12466 25516 12544
rect 25752 12543 25920 12544
rect 25414 12465 25516 12466
rect 25413 12457 25516 12465
rect 25413 12454 25465 12457
rect 25413 12419 25421 12454
rect 25446 12419 25465 12454
rect 25490 12419 25516 12457
rect 25413 12413 25516 12419
rect 25676 12458 25712 12462
rect 25676 12435 25684 12458
rect 25708 12435 25712 12458
rect 25676 12414 25712 12435
rect 25413 12409 25512 12413
rect 25676 12391 25684 12414
rect 25708 12391 25712 12414
rect 24305 11825 24473 11827
rect 24029 11799 24473 11825
rect 22225 11732 22290 11779
rect 22225 11714 22248 11732
rect 22266 11714 22290 11732
rect 23138 11759 23173 11761
rect 23138 11757 23242 11759
rect 24031 11757 24070 11799
rect 24305 11798 24473 11799
rect 23138 11750 24072 11757
rect 23138 11749 23189 11750
rect 23138 11729 23141 11749
rect 23166 11730 23189 11749
rect 23221 11730 24072 11750
rect 23166 11729 24072 11730
rect 23138 11722 24072 11729
rect 23411 11721 24072 11722
rect 22225 11693 22290 11714
rect 22502 11704 22542 11707
rect 22502 11700 23405 11704
rect 22502 11680 23379 11700
rect 23399 11680 23405 11700
rect 22502 11677 23405 11680
rect 22226 11633 22291 11653
rect 22226 11615 22250 11633
rect 22268 11615 22291 11633
rect 22226 11588 22291 11615
rect 22502 11588 22542 11677
rect 22986 11675 23402 11677
rect 22986 11674 23327 11675
rect 22643 11643 22753 11657
rect 22643 11640 22686 11643
rect 22643 11635 22647 11640
rect 22225 11553 22542 11588
rect 22565 11613 22647 11635
rect 22676 11613 22686 11640
rect 22714 11616 22721 11643
rect 22750 11635 22753 11643
rect 22750 11616 22815 11635
rect 22714 11613 22815 11616
rect 22565 11611 22815 11613
rect 20926 11520 20948 11538
rect 20966 11520 20991 11538
rect 20926 11501 20991 11520
rect 20619 11476 20656 11477
rect 20042 11455 20078 11476
rect 20468 11455 20499 11476
rect 20706 11471 20714 11480
rect 20703 11455 20714 11471
rect 19875 11451 19975 11455
rect 19875 11447 19937 11451
rect 19875 11421 19882 11447
rect 19908 11425 19937 11447
rect 19963 11425 19975 11451
rect 19908 11421 19975 11425
rect 19875 11418 19975 11421
rect 20043 11418 20078 11455
rect 20140 11452 20499 11455
rect 20140 11447 20362 11452
rect 20140 11423 20153 11447
rect 20177 11428 20362 11447
rect 20386 11428 20499 11452
rect 20177 11423 20499 11428
rect 20140 11419 20499 11423
rect 20566 11447 20714 11455
rect 20566 11427 20577 11447
rect 20597 11438 20714 11447
rect 20763 11471 20770 11480
rect 22226 11477 22291 11553
rect 22565 11532 22602 11611
rect 22643 11598 22753 11611
rect 22717 11542 22748 11543
rect 22565 11512 22574 11532
rect 22594 11512 22602 11532
rect 22565 11502 22602 11512
rect 22661 11532 22748 11542
rect 22661 11512 22670 11532
rect 22690 11512 22748 11532
rect 22661 11503 22748 11512
rect 22661 11502 22698 11503
rect 20763 11438 20771 11471
rect 22226 11459 22248 11477
rect 22266 11459 22291 11477
rect 20597 11427 20771 11438
rect 20566 11420 20771 11427
rect 20566 11419 20607 11420
rect 20042 11393 20078 11418
rect 19890 11366 19927 11367
rect 19986 11366 20023 11367
rect 20042 11366 20049 11393
rect 19566 11341 19574 11361
rect 19594 11341 19603 11361
rect 19420 11330 19451 11331
rect 19415 11262 19525 11275
rect 19566 11262 19603 11341
rect 19790 11357 19928 11366
rect 19790 11337 19899 11357
rect 19919 11337 19928 11357
rect 19790 11330 19928 11337
rect 19986 11363 20049 11366
rect 20070 11366 20078 11393
rect 20097 11366 20134 11367
rect 20070 11363 20134 11366
rect 19986 11357 20134 11363
rect 19986 11337 19995 11357
rect 20015 11337 20105 11357
rect 20125 11337 20134 11357
rect 19790 11328 19886 11330
rect 19986 11327 20134 11337
rect 20193 11357 20230 11367
rect 20305 11366 20342 11367
rect 20286 11364 20342 11366
rect 20193 11337 20201 11357
rect 20221 11337 20230 11357
rect 20042 11326 20078 11327
rect 19353 11260 19603 11262
rect 19353 11257 19454 11260
rect 19353 11238 19418 11257
rect 19415 11230 19418 11238
rect 19447 11230 19454 11257
rect 19482 11233 19492 11260
rect 19521 11238 19603 11260
rect 19521 11233 19525 11238
rect 19482 11230 19525 11233
rect 19415 11216 19525 11230
rect 18841 11198 19182 11199
rect 18766 11193 19182 11198
rect 19890 11195 19927 11196
rect 20193 11195 20230 11337
rect 20255 11357 20342 11364
rect 20255 11354 20313 11357
rect 20255 11334 20260 11354
rect 20281 11337 20313 11354
rect 20333 11337 20342 11357
rect 20281 11334 20342 11337
rect 20255 11327 20342 11334
rect 20401 11357 20438 11367
rect 20401 11337 20409 11357
rect 20429 11337 20438 11357
rect 20255 11326 20286 11327
rect 20401 11258 20438 11337
rect 20468 11366 20499 11419
rect 20703 11417 20771 11420
rect 20703 11375 20715 11417
rect 20764 11375 20771 11417
rect 20518 11366 20555 11367
rect 20468 11357 20555 11366
rect 20468 11337 20526 11357
rect 20546 11337 20555 11357
rect 20468 11327 20555 11337
rect 20614 11357 20651 11367
rect 20703 11362 20771 11375
rect 20926 11439 20991 11456
rect 20926 11421 20950 11439
rect 20968 11421 20991 11439
rect 22226 11438 22291 11459
rect 22439 11457 22504 11466
rect 20614 11337 20622 11357
rect 20642 11337 20651 11357
rect 20468 11326 20499 11327
rect 20463 11258 20573 11271
rect 20614 11258 20651 11337
rect 20926 11282 20991 11421
rect 22439 11420 22449 11457
rect 22489 11449 22504 11457
rect 22717 11450 22748 11503
rect 22778 11532 22815 11611
rect 22930 11542 22961 11543
rect 22778 11512 22787 11532
rect 22807 11512 22815 11532
rect 22778 11502 22815 11512
rect 22874 11535 22961 11542
rect 22874 11532 22935 11535
rect 22874 11512 22883 11532
rect 22903 11515 22935 11532
rect 22956 11515 22961 11535
rect 22903 11512 22961 11515
rect 22874 11505 22961 11512
rect 22986 11532 23023 11674
rect 23289 11673 23326 11674
rect 23138 11542 23174 11543
rect 22986 11512 22995 11532
rect 23015 11512 23023 11532
rect 22874 11503 22930 11505
rect 22874 11502 22911 11503
rect 22986 11502 23023 11512
rect 23082 11532 23230 11542
rect 23330 11539 23426 11541
rect 23082 11512 23091 11532
rect 23111 11512 23201 11532
rect 23221 11512 23230 11532
rect 23082 11506 23230 11512
rect 23082 11503 23146 11506
rect 23082 11502 23119 11503
rect 23138 11476 23146 11503
rect 23167 11503 23230 11506
rect 23288 11532 23426 11539
rect 23288 11512 23297 11532
rect 23317 11512 23426 11532
rect 23288 11503 23426 11512
rect 23167 11476 23174 11503
rect 23193 11502 23230 11503
rect 23289 11502 23326 11503
rect 23138 11451 23174 11476
rect 22609 11449 22650 11450
rect 22489 11442 22650 11449
rect 22489 11422 22619 11442
rect 22639 11422 22650 11442
rect 22489 11420 22650 11422
rect 22439 11414 22650 11420
rect 22717 11446 23076 11450
rect 22717 11441 23039 11446
rect 22717 11417 22830 11441
rect 22854 11422 23039 11441
rect 23063 11422 23076 11446
rect 22854 11417 23076 11422
rect 22717 11414 23076 11417
rect 23138 11414 23173 11451
rect 23241 11448 23341 11451
rect 23241 11444 23308 11448
rect 23241 11418 23253 11444
rect 23279 11422 23308 11444
rect 23334 11422 23341 11448
rect 23279 11418 23341 11422
rect 23241 11414 23341 11418
rect 22439 11401 22506 11414
rect 20926 11276 20948 11282
rect 20401 11256 20651 11258
rect 20401 11253 20502 11256
rect 20401 11234 20466 11253
rect 20463 11226 20466 11234
rect 20495 11226 20502 11253
rect 20530 11229 20540 11256
rect 20569 11234 20651 11256
rect 20680 11264 20948 11276
rect 20966 11264 20991 11282
rect 20680 11241 20991 11264
rect 22231 11378 22287 11398
rect 22231 11360 22250 11378
rect 22268 11360 22287 11378
rect 22231 11247 22287 11360
rect 22439 11380 22453 11401
rect 22489 11380 22506 11401
rect 22717 11393 22748 11414
rect 23138 11393 23174 11414
rect 22560 11392 22597 11393
rect 22439 11373 22506 11380
rect 22559 11383 22597 11392
rect 20680 11240 20735 11241
rect 20569 11229 20573 11234
rect 20530 11226 20573 11229
rect 20463 11212 20573 11226
rect 19889 11194 20230 11195
rect 18766 11173 18769 11193
rect 18789 11173 19182 11193
rect 19814 11193 20230 11194
rect 20680 11193 20723 11240
rect 19814 11189 20723 11193
rect 19133 11140 19178 11173
rect 19814 11169 19817 11189
rect 19837 11169 20723 11189
rect 20191 11164 20723 11169
rect 20931 11183 20990 11205
rect 20931 11165 20950 11183
rect 20968 11165 20990 11183
rect 19979 11140 20078 11142
rect 19133 11130 20078 11140
rect 19133 11104 20001 11130
rect 19134 11103 20001 11104
rect 19979 11092 20001 11103
rect 20026 11095 20045 11130
rect 20070 11095 20078 11130
rect 20026 11092 20078 11095
rect 19979 11084 20078 11092
rect 20005 11083 20077 11084
rect 20931 11035 20990 11165
rect 22231 11118 22286 11247
rect 22439 11221 22504 11373
rect 22559 11363 22568 11383
rect 22588 11363 22597 11383
rect 22559 11355 22597 11363
rect 22663 11387 22748 11393
rect 22773 11392 22810 11393
rect 22663 11367 22671 11387
rect 22691 11367 22748 11387
rect 22663 11359 22748 11367
rect 22772 11383 22810 11392
rect 22772 11363 22781 11383
rect 22801 11363 22810 11383
rect 22663 11358 22699 11359
rect 22772 11355 22810 11363
rect 22876 11387 22961 11393
rect 22981 11392 23018 11393
rect 22876 11367 22884 11387
rect 22904 11386 22961 11387
rect 22904 11367 22933 11386
rect 22876 11366 22933 11367
rect 22954 11366 22961 11386
rect 22876 11359 22961 11366
rect 22980 11383 23018 11392
rect 22980 11363 22989 11383
rect 23009 11363 23018 11383
rect 22876 11358 22912 11359
rect 22980 11355 23018 11363
rect 23084 11387 23228 11393
rect 23084 11367 23092 11387
rect 23112 11367 23200 11387
rect 23220 11367 23228 11387
rect 23084 11359 23228 11367
rect 23084 11358 23120 11359
rect 23192 11358 23228 11359
rect 23294 11392 23331 11393
rect 23294 11391 23332 11392
rect 23294 11383 23358 11391
rect 23294 11363 23303 11383
rect 23323 11369 23358 11383
rect 23378 11369 23381 11389
rect 23323 11364 23381 11369
rect 23323 11363 23358 11364
rect 22560 11326 22597 11355
rect 22561 11324 22597 11326
rect 22773 11324 22810 11355
rect 22561 11302 22810 11324
rect 22642 11296 22753 11302
rect 22642 11288 22683 11296
rect 22642 11268 22650 11288
rect 22669 11268 22683 11288
rect 22642 11266 22683 11268
rect 22711 11288 22753 11296
rect 22711 11268 22727 11288
rect 22746 11268 22753 11288
rect 22711 11266 22753 11268
rect 22642 11251 22753 11266
rect 22981 11256 23018 11355
rect 23294 11351 23358 11363
rect 22644 11242 22748 11251
rect 22432 11211 22553 11221
rect 22432 11209 22501 11211
rect 22432 11168 22445 11209
rect 22482 11170 22501 11209
rect 22538 11170 22553 11211
rect 22482 11168 22553 11170
rect 22432 11150 22553 11168
rect 22225 11106 22286 11118
rect 22979 11106 23020 11256
rect 23398 11248 23425 11503
rect 23487 11493 23567 11504
rect 23487 11467 23504 11493
rect 23544 11467 23567 11493
rect 23487 11440 23567 11467
rect 23487 11414 23508 11440
rect 23548 11414 23567 11440
rect 23487 11395 23567 11414
rect 23487 11369 23511 11395
rect 23551 11369 23567 11395
rect 23487 11318 23567 11369
rect 22225 11103 23020 11106
rect 23399 11117 23425 11248
rect 23489 11162 23559 11318
rect 23488 11146 23564 11162
rect 23399 11103 23427 11117
rect 22225 11068 23427 11103
rect 23488 11109 23503 11146
rect 23547 11109 23564 11146
rect 23488 11089 23564 11109
rect 24602 11139 24672 12048
rect 24771 11483 24852 12196
rect 25676 12082 25712 12391
rect 25600 12053 25713 12082
rect 25600 11697 25631 12053
rect 25670 11798 26661 11823
rect 25670 11793 25730 11798
rect 25670 11772 25689 11793
rect 25709 11777 25730 11793
rect 25750 11777 26661 11798
rect 25709 11772 26661 11777
rect 25670 11764 26661 11772
rect 25675 11741 25781 11764
rect 25675 11738 25780 11741
rect 25524 11677 25917 11697
rect 25937 11677 25940 11697
rect 25524 11672 25940 11677
rect 25524 11671 25865 11672
rect 25181 11640 25291 11654
rect 25181 11637 25224 11640
rect 25181 11632 25185 11637
rect 25103 11610 25185 11632
rect 25214 11610 25224 11637
rect 25252 11613 25259 11640
rect 25288 11632 25291 11640
rect 25288 11613 25353 11632
rect 25252 11610 25353 11613
rect 25103 11608 25353 11610
rect 25103 11529 25140 11608
rect 25181 11595 25291 11608
rect 25255 11539 25286 11540
rect 25103 11509 25112 11529
rect 25132 11509 25140 11529
rect 25103 11499 25140 11509
rect 25199 11529 25286 11539
rect 25199 11509 25208 11529
rect 25228 11509 25286 11529
rect 25199 11500 25286 11509
rect 25199 11499 25236 11500
rect 24769 11447 24861 11483
rect 25255 11447 25286 11500
rect 25316 11529 25353 11608
rect 25468 11539 25499 11540
rect 25316 11509 25325 11529
rect 25345 11509 25353 11529
rect 25316 11499 25353 11509
rect 25412 11532 25499 11539
rect 25412 11529 25473 11532
rect 25412 11509 25421 11529
rect 25441 11512 25473 11529
rect 25494 11512 25499 11532
rect 25441 11509 25499 11512
rect 25412 11502 25499 11509
rect 25524 11529 25561 11671
rect 25827 11670 25864 11671
rect 25676 11539 25712 11540
rect 25524 11509 25533 11529
rect 25553 11509 25561 11529
rect 25412 11500 25468 11502
rect 25412 11499 25449 11500
rect 25524 11499 25561 11509
rect 25620 11529 25768 11539
rect 25868 11536 25964 11538
rect 25620 11509 25629 11529
rect 25649 11509 25739 11529
rect 25759 11509 25768 11529
rect 25620 11503 25768 11509
rect 25620 11500 25684 11503
rect 25620 11499 25657 11500
rect 25676 11473 25684 11500
rect 25705 11500 25768 11503
rect 25826 11529 25964 11536
rect 25826 11509 25835 11529
rect 25855 11509 25964 11529
rect 25826 11500 25964 11509
rect 25705 11473 25712 11500
rect 25731 11499 25768 11500
rect 25827 11499 25864 11500
rect 25676 11448 25712 11473
rect 24769 11446 25105 11447
rect 25147 11446 25188 11447
rect 24769 11439 25188 11446
rect 24769 11419 25157 11439
rect 25177 11419 25188 11439
rect 24769 11411 25188 11419
rect 25255 11443 25614 11447
rect 25255 11438 25577 11443
rect 25255 11414 25368 11438
rect 25392 11419 25577 11438
rect 25601 11419 25614 11443
rect 25392 11414 25614 11419
rect 25255 11411 25614 11414
rect 25676 11411 25711 11448
rect 25779 11445 25879 11448
rect 25779 11441 25846 11445
rect 25779 11415 25791 11441
rect 25817 11419 25846 11441
rect 25872 11419 25879 11445
rect 25817 11415 25879 11419
rect 25779 11411 25879 11415
rect 24769 11407 25105 11411
rect 24602 11089 24674 11139
rect 19653 11005 19729 11029
rect 19653 10939 19665 11005
rect 19719 10939 19729 11005
rect 20197 10960 20238 10962
rect 20469 10960 20573 10962
rect 20931 10960 20992 11035
rect 22225 10993 22286 11068
rect 22644 11066 22748 11068
rect 22979 11066 23020 11068
rect 23488 11023 23498 11089
rect 23552 11023 23564 11089
rect 23488 10999 23564 11023
rect 18543 10889 18615 10939
rect 17254 10797 17698 10823
rect 17254 10795 17422 10797
rect 17254 10528 17281 10795
rect 17551 10793 17580 10797
rect 17321 10668 17385 10680
rect 17661 10676 17698 10797
rect 17926 10765 18037 10780
rect 17926 10763 17968 10765
rect 17926 10743 17933 10763
rect 17952 10743 17968 10763
rect 17926 10735 17968 10743
rect 17996 10763 18037 10765
rect 17996 10743 18010 10763
rect 18029 10743 18037 10763
rect 17996 10735 18037 10743
rect 17926 10729 18037 10735
rect 17869 10707 18118 10729
rect 17869 10676 17906 10707
rect 18082 10705 18118 10707
rect 18082 10676 18119 10705
rect 17321 10667 17356 10668
rect 17298 10662 17356 10667
rect 17298 10642 17301 10662
rect 17321 10648 17356 10662
rect 17376 10648 17385 10668
rect 17321 10640 17385 10648
rect 17347 10639 17385 10640
rect 17348 10638 17385 10639
rect 17451 10672 17487 10673
rect 17559 10672 17595 10673
rect 17451 10664 17595 10672
rect 17451 10644 17459 10664
rect 17479 10644 17567 10664
rect 17587 10644 17595 10664
rect 17451 10638 17595 10644
rect 17661 10668 17699 10676
rect 17767 10672 17803 10673
rect 17661 10648 17670 10668
rect 17690 10648 17699 10668
rect 17661 10639 17699 10648
rect 17718 10665 17803 10672
rect 17718 10645 17725 10665
rect 17746 10664 17803 10665
rect 17746 10645 17775 10664
rect 17718 10644 17775 10645
rect 17795 10644 17803 10664
rect 17661 10638 17698 10639
rect 17718 10638 17803 10644
rect 17869 10668 17907 10676
rect 17980 10672 18016 10673
rect 17869 10648 17878 10668
rect 17898 10648 17907 10668
rect 17869 10639 17907 10648
rect 17931 10664 18016 10672
rect 17931 10644 17988 10664
rect 18008 10644 18016 10664
rect 17869 10638 17906 10639
rect 17931 10638 18016 10644
rect 18082 10668 18120 10676
rect 18082 10648 18091 10668
rect 18111 10648 18120 10668
rect 18082 10639 18120 10648
rect 18082 10638 18119 10639
rect 17505 10617 17541 10638
rect 17931 10617 17962 10638
rect 18112 10617 18446 10621
rect 17338 10613 17438 10617
rect 17338 10609 17400 10613
rect 17338 10583 17345 10609
rect 17371 10587 17400 10609
rect 17426 10587 17438 10613
rect 17371 10583 17438 10587
rect 17338 10580 17438 10583
rect 17506 10580 17541 10617
rect 17603 10614 17962 10617
rect 17603 10609 17825 10614
rect 17603 10585 17616 10609
rect 17640 10590 17825 10609
rect 17849 10590 17962 10614
rect 17640 10585 17962 10590
rect 17603 10581 17962 10585
rect 18029 10609 18446 10617
rect 18029 10589 18040 10609
rect 18060 10589 18446 10609
rect 18029 10582 18446 10589
rect 18029 10581 18070 10582
rect 18112 10581 18446 10582
rect 17505 10555 17541 10580
rect 17353 10528 17390 10529
rect 17449 10528 17486 10529
rect 17505 10528 17512 10555
rect 17253 10519 17391 10528
rect 17253 10499 17362 10519
rect 17382 10499 17391 10519
rect 17253 10492 17391 10499
rect 17449 10525 17512 10528
rect 17533 10528 17541 10555
rect 17560 10528 17597 10529
rect 17533 10525 17597 10528
rect 17449 10519 17597 10525
rect 17449 10499 17458 10519
rect 17478 10499 17568 10519
rect 17588 10499 17597 10519
rect 17253 10490 17349 10492
rect 17449 10489 17597 10499
rect 17656 10519 17693 10529
rect 17768 10528 17805 10529
rect 17749 10526 17805 10528
rect 17656 10499 17664 10519
rect 17684 10499 17693 10519
rect 17505 10488 17541 10489
rect 17353 10357 17390 10358
rect 17656 10357 17693 10499
rect 17718 10519 17805 10526
rect 17718 10516 17776 10519
rect 17718 10496 17723 10516
rect 17744 10499 17776 10516
rect 17796 10499 17805 10519
rect 17744 10496 17805 10499
rect 17718 10489 17805 10496
rect 17864 10519 17901 10529
rect 17864 10499 17872 10519
rect 17892 10499 17901 10519
rect 17718 10488 17749 10489
rect 17864 10420 17901 10499
rect 17931 10528 17962 10581
rect 17981 10528 18018 10529
rect 17931 10519 18018 10528
rect 17931 10499 17989 10519
rect 18009 10499 18018 10519
rect 17931 10489 18018 10499
rect 18077 10519 18114 10529
rect 18077 10499 18085 10519
rect 18105 10499 18114 10519
rect 17931 10488 17962 10489
rect 17926 10420 18036 10433
rect 18077 10420 18114 10499
rect 17864 10418 18114 10420
rect 17864 10415 17965 10418
rect 17864 10396 17929 10415
rect 17926 10388 17929 10396
rect 17958 10388 17965 10415
rect 17993 10391 18003 10418
rect 18032 10396 18114 10418
rect 18032 10391 18036 10396
rect 17993 10388 18036 10391
rect 17926 10374 18036 10388
rect 17352 10356 17693 10357
rect 17277 10351 17693 10356
rect 17277 10331 17280 10351
rect 17300 10331 17693 10351
rect 17586 9966 17617 10331
rect 17504 9937 17617 9966
rect 17505 9637 17541 9937
rect 18365 9832 18446 10581
rect 18545 9980 18615 10889
rect 19653 10919 19729 10939
rect 19653 10882 19670 10919
rect 19714 10882 19729 10919
rect 19790 10925 20992 10960
rect 19790 10911 19818 10925
rect 19653 10866 19729 10882
rect 19658 10710 19728 10866
rect 19792 10780 19818 10911
rect 20197 10922 20992 10925
rect 19650 10659 19730 10710
rect 19650 10633 19666 10659
rect 19706 10633 19730 10659
rect 19650 10614 19730 10633
rect 19650 10588 19669 10614
rect 19709 10588 19730 10614
rect 19650 10561 19730 10588
rect 19650 10535 19673 10561
rect 19713 10535 19730 10561
rect 19650 10524 19730 10535
rect 19792 10525 19819 10780
rect 20197 10772 20238 10922
rect 20931 10910 20992 10922
rect 20664 10860 20785 10878
rect 20664 10858 20735 10860
rect 20664 10817 20679 10858
rect 20716 10819 20735 10858
rect 20772 10819 20785 10860
rect 20716 10817 20785 10819
rect 20664 10807 20785 10817
rect 20469 10777 20573 10786
rect 19859 10665 19923 10677
rect 20199 10673 20236 10772
rect 20464 10762 20575 10777
rect 20464 10760 20506 10762
rect 20464 10740 20471 10760
rect 20490 10740 20506 10760
rect 20464 10732 20506 10740
rect 20534 10760 20575 10762
rect 20534 10740 20548 10760
rect 20567 10740 20575 10760
rect 20534 10732 20575 10740
rect 20464 10726 20575 10732
rect 20407 10704 20656 10726
rect 20407 10673 20444 10704
rect 20620 10702 20656 10704
rect 20620 10673 20657 10702
rect 19859 10664 19894 10665
rect 19836 10659 19894 10664
rect 19836 10639 19839 10659
rect 19859 10645 19894 10659
rect 19914 10645 19923 10665
rect 19859 10637 19923 10645
rect 19885 10636 19923 10637
rect 19886 10635 19923 10636
rect 19989 10669 20025 10670
rect 20097 10669 20133 10670
rect 19989 10661 20133 10669
rect 19989 10641 19997 10661
rect 20017 10641 20105 10661
rect 20125 10641 20133 10661
rect 19989 10635 20133 10641
rect 20199 10665 20237 10673
rect 20305 10669 20341 10670
rect 20199 10645 20208 10665
rect 20228 10645 20237 10665
rect 20199 10636 20237 10645
rect 20256 10662 20341 10669
rect 20256 10642 20263 10662
rect 20284 10661 20341 10662
rect 20284 10642 20313 10661
rect 20256 10641 20313 10642
rect 20333 10641 20341 10661
rect 20199 10635 20236 10636
rect 20256 10635 20341 10641
rect 20407 10665 20445 10673
rect 20518 10669 20554 10670
rect 20407 10645 20416 10665
rect 20436 10645 20445 10665
rect 20407 10636 20445 10645
rect 20469 10661 20554 10669
rect 20469 10641 20526 10661
rect 20546 10641 20554 10661
rect 20407 10635 20444 10636
rect 20469 10635 20554 10641
rect 20620 10665 20658 10673
rect 20620 10645 20629 10665
rect 20649 10645 20658 10665
rect 20713 10655 20778 10807
rect 20931 10781 20986 10910
rect 22227 10863 22286 10993
rect 23140 10944 23212 10945
rect 23139 10936 23238 10944
rect 23139 10933 23191 10936
rect 23139 10898 23147 10933
rect 23172 10898 23191 10933
rect 23216 10925 23238 10936
rect 23216 10924 24083 10925
rect 23216 10898 24084 10924
rect 23139 10888 24084 10898
rect 23139 10886 23238 10888
rect 22227 10845 22249 10863
rect 22267 10845 22286 10863
rect 22227 10823 22286 10845
rect 22494 10859 23026 10864
rect 22494 10839 23380 10859
rect 23400 10839 23403 10859
rect 24039 10855 24084 10888
rect 22494 10835 23403 10839
rect 22494 10788 22537 10835
rect 22987 10834 23403 10835
rect 24035 10835 24428 10855
rect 24448 10835 24451 10855
rect 22987 10833 23328 10834
rect 22644 10802 22754 10816
rect 22644 10799 22687 10802
rect 22644 10794 22648 10799
rect 22482 10787 22537 10788
rect 20620 10636 20658 10645
rect 20711 10648 20778 10655
rect 20620 10635 20657 10636
rect 20043 10614 20079 10635
rect 20469 10614 20500 10635
rect 20711 10627 20728 10648
rect 20764 10627 20778 10648
rect 20930 10668 20986 10781
rect 20930 10650 20949 10668
rect 20967 10650 20986 10668
rect 20930 10630 20986 10650
rect 22226 10764 22537 10787
rect 22226 10746 22251 10764
rect 22269 10752 22537 10764
rect 22566 10772 22648 10794
rect 22677 10772 22687 10799
rect 22715 10775 22722 10802
rect 22751 10794 22754 10802
rect 22751 10775 22816 10794
rect 22715 10772 22816 10775
rect 22566 10770 22816 10772
rect 22269 10746 22291 10752
rect 20711 10614 20778 10627
rect 19876 10610 19976 10614
rect 19876 10606 19938 10610
rect 19876 10580 19883 10606
rect 19909 10584 19938 10606
rect 19964 10584 19976 10610
rect 19909 10580 19976 10584
rect 19876 10577 19976 10580
rect 20044 10577 20079 10614
rect 20141 10611 20500 10614
rect 20141 10606 20363 10611
rect 20141 10582 20154 10606
rect 20178 10587 20363 10606
rect 20387 10587 20500 10611
rect 20178 10582 20500 10587
rect 20141 10578 20500 10582
rect 20567 10608 20778 10614
rect 20567 10606 20728 10608
rect 20567 10586 20578 10606
rect 20598 10586 20728 10606
rect 20567 10579 20728 10586
rect 20567 10578 20608 10579
rect 20043 10552 20079 10577
rect 19891 10525 19928 10526
rect 19987 10525 20024 10526
rect 20043 10525 20050 10552
rect 19791 10516 19929 10525
rect 19791 10496 19900 10516
rect 19920 10496 19929 10516
rect 19791 10489 19929 10496
rect 19987 10522 20050 10525
rect 20071 10525 20079 10552
rect 20098 10525 20135 10526
rect 20071 10522 20135 10525
rect 19987 10516 20135 10522
rect 19987 10496 19996 10516
rect 20016 10496 20106 10516
rect 20126 10496 20135 10516
rect 19791 10487 19887 10489
rect 19987 10486 20135 10496
rect 20194 10516 20231 10526
rect 20306 10525 20343 10526
rect 20287 10523 20343 10525
rect 20194 10496 20202 10516
rect 20222 10496 20231 10516
rect 20043 10485 20079 10486
rect 19891 10354 19928 10355
rect 20194 10354 20231 10496
rect 20256 10516 20343 10523
rect 20256 10513 20314 10516
rect 20256 10493 20261 10513
rect 20282 10496 20314 10513
rect 20334 10496 20343 10516
rect 20282 10493 20343 10496
rect 20256 10486 20343 10493
rect 20402 10516 20439 10526
rect 20402 10496 20410 10516
rect 20430 10496 20439 10516
rect 20256 10485 20287 10486
rect 20402 10417 20439 10496
rect 20469 10525 20500 10578
rect 20713 10571 20728 10579
rect 20768 10571 20778 10608
rect 22226 10607 22291 10746
rect 22566 10691 22603 10770
rect 22644 10757 22754 10770
rect 22718 10701 22749 10702
rect 22566 10671 22575 10691
rect 22595 10671 22603 10691
rect 20713 10562 20778 10571
rect 20926 10569 20991 10590
rect 22226 10589 22249 10607
rect 22267 10589 22291 10607
rect 22226 10572 22291 10589
rect 22446 10653 22514 10666
rect 22566 10661 22603 10671
rect 22662 10691 22749 10701
rect 22662 10671 22671 10691
rect 22691 10671 22749 10691
rect 22662 10662 22749 10671
rect 22662 10661 22699 10662
rect 22446 10611 22453 10653
rect 22502 10611 22514 10653
rect 22446 10608 22514 10611
rect 22718 10609 22749 10662
rect 22779 10691 22816 10770
rect 22931 10701 22962 10702
rect 22779 10671 22788 10691
rect 22808 10671 22816 10691
rect 22779 10661 22816 10671
rect 22875 10694 22962 10701
rect 22875 10691 22936 10694
rect 22875 10671 22884 10691
rect 22904 10674 22936 10691
rect 22957 10674 22962 10694
rect 22904 10671 22962 10674
rect 22875 10664 22962 10671
rect 22987 10691 23024 10833
rect 23290 10832 23327 10833
rect 24035 10830 24451 10835
rect 24035 10829 24376 10830
rect 23692 10798 23802 10812
rect 23692 10795 23735 10798
rect 23692 10790 23696 10795
rect 23614 10768 23696 10790
rect 23725 10768 23735 10795
rect 23763 10771 23770 10798
rect 23799 10790 23802 10798
rect 23799 10771 23864 10790
rect 23763 10768 23864 10771
rect 23614 10766 23864 10768
rect 23139 10701 23175 10702
rect 22987 10671 22996 10691
rect 23016 10671 23024 10691
rect 22875 10662 22931 10664
rect 22875 10661 22912 10662
rect 22987 10661 23024 10671
rect 23083 10691 23231 10701
rect 23331 10698 23427 10700
rect 23083 10671 23092 10691
rect 23112 10671 23202 10691
rect 23222 10671 23231 10691
rect 23083 10665 23231 10671
rect 23083 10662 23147 10665
rect 23083 10661 23120 10662
rect 23139 10635 23147 10662
rect 23168 10662 23231 10665
rect 23289 10691 23427 10698
rect 23289 10671 23298 10691
rect 23318 10671 23427 10691
rect 23289 10662 23427 10671
rect 23614 10687 23651 10766
rect 23692 10753 23802 10766
rect 23766 10697 23797 10698
rect 23614 10667 23623 10687
rect 23643 10667 23651 10687
rect 23168 10635 23175 10662
rect 23194 10661 23231 10662
rect 23290 10661 23327 10662
rect 23139 10610 23175 10635
rect 22610 10608 22651 10609
rect 22446 10601 22651 10608
rect 22446 10590 22620 10601
rect 20926 10551 20951 10569
rect 20969 10551 20991 10569
rect 22446 10557 22454 10590
rect 20519 10525 20556 10526
rect 20469 10516 20556 10525
rect 20469 10496 20527 10516
rect 20547 10496 20556 10516
rect 20469 10486 20556 10496
rect 20615 10516 20652 10526
rect 20615 10496 20623 10516
rect 20643 10496 20652 10516
rect 20469 10485 20500 10486
rect 20464 10417 20574 10430
rect 20615 10417 20652 10496
rect 20926 10475 20991 10551
rect 22447 10548 22454 10557
rect 22503 10581 22620 10590
rect 22640 10581 22651 10601
rect 22503 10573 22651 10581
rect 22718 10605 23077 10609
rect 22718 10600 23040 10605
rect 22718 10576 22831 10600
rect 22855 10581 23040 10600
rect 23064 10581 23077 10605
rect 22855 10576 23077 10581
rect 22718 10573 23077 10576
rect 23139 10573 23174 10610
rect 23242 10607 23342 10610
rect 23242 10603 23309 10607
rect 23242 10577 23254 10603
rect 23280 10581 23309 10603
rect 23335 10581 23342 10607
rect 23280 10577 23342 10581
rect 23242 10573 23342 10577
rect 22503 10557 22514 10573
rect 22503 10548 22511 10557
rect 22718 10552 22749 10573
rect 23139 10552 23175 10573
rect 22561 10551 22598 10552
rect 22226 10508 22291 10527
rect 22226 10490 22251 10508
rect 22269 10490 22291 10508
rect 20402 10415 20652 10417
rect 20402 10412 20503 10415
rect 20402 10393 20467 10412
rect 20464 10385 20467 10393
rect 20496 10385 20503 10412
rect 20531 10388 20541 10415
rect 20570 10393 20652 10415
rect 20675 10440 20992 10475
rect 20570 10388 20574 10393
rect 20531 10385 20574 10388
rect 20464 10371 20574 10385
rect 19890 10353 20231 10354
rect 19815 10351 20231 10353
rect 20675 10351 20715 10440
rect 20926 10413 20991 10440
rect 20926 10395 20949 10413
rect 20967 10395 20991 10413
rect 20926 10375 20991 10395
rect 19812 10348 20715 10351
rect 19812 10328 19818 10348
rect 19838 10328 20715 10348
rect 19812 10324 20715 10328
rect 20675 10321 20715 10324
rect 20927 10314 20992 10335
rect 19145 10306 19806 10307
rect 19145 10299 20079 10306
rect 19145 10298 20051 10299
rect 19145 10278 19996 10298
rect 20028 10279 20051 10298
rect 20076 10279 20079 10299
rect 20028 10278 20079 10279
rect 19145 10271 20079 10278
rect 18744 10229 18912 10230
rect 19147 10229 19186 10271
rect 19975 10269 20079 10271
rect 20044 10267 20079 10269
rect 20927 10296 20951 10314
rect 20969 10296 20992 10314
rect 20927 10249 20992 10296
rect 18744 10203 19188 10229
rect 18744 10201 18912 10203
rect 17505 9614 17509 9637
rect 17533 9614 17541 9637
rect 17705 9615 17804 9619
rect 17505 9593 17541 9614
rect 17505 9570 17509 9593
rect 17533 9570 17541 9593
rect 17505 9566 17541 9570
rect 17701 9609 17804 9615
rect 17701 9571 17727 9609
rect 17752 9574 17771 9609
rect 17796 9574 17804 9609
rect 17752 9571 17804 9574
rect 17701 9563 17804 9571
rect 17701 9562 17803 9563
rect 17297 9484 17465 9485
rect 17701 9484 17748 9562
rect 17297 9458 17748 9484
rect 17297 9456 17465 9458
rect 17297 9083 17324 9456
rect 17494 9408 17580 9417
rect 17494 9390 17513 9408
rect 17565 9390 17580 9408
rect 17494 9386 17580 9390
rect 17364 9223 17428 9235
rect 17364 9222 17399 9223
rect 17341 9217 17399 9222
rect 17341 9197 17344 9217
rect 17364 9203 17399 9217
rect 17419 9203 17428 9223
rect 17364 9195 17428 9203
rect 17390 9194 17428 9195
rect 17391 9193 17428 9194
rect 17494 9227 17530 9228
rect 17550 9227 17580 9386
rect 17701 9346 17748 9458
rect 17704 9231 17741 9346
rect 17969 9320 18080 9335
rect 17969 9318 18011 9320
rect 17969 9298 17976 9318
rect 17995 9298 18011 9318
rect 17969 9290 18011 9298
rect 18039 9318 18080 9320
rect 18039 9298 18053 9318
rect 18072 9298 18080 9318
rect 18039 9290 18080 9298
rect 17969 9284 18080 9290
rect 17912 9262 18161 9284
rect 17912 9231 17949 9262
rect 18125 9260 18161 9262
rect 18125 9231 18162 9260
rect 18366 9247 18445 9832
rect 18542 9380 18621 9980
rect 18744 9850 18771 10201
rect 19147 10197 19188 10203
rect 18811 9990 18875 10002
rect 19151 9998 19188 10197
rect 19650 10224 19722 10241
rect 19650 10185 19658 10224
rect 19703 10185 19722 10224
rect 19416 10087 19527 10102
rect 19416 10085 19458 10087
rect 19416 10065 19423 10085
rect 19442 10065 19458 10085
rect 19416 10057 19458 10065
rect 19486 10085 19527 10087
rect 19486 10065 19500 10085
rect 19519 10065 19527 10085
rect 19486 10057 19527 10065
rect 19416 10051 19527 10057
rect 19359 10029 19608 10051
rect 19359 9998 19396 10029
rect 19572 10027 19608 10029
rect 19572 9998 19609 10027
rect 18811 9989 18846 9990
rect 18788 9984 18846 9989
rect 18788 9964 18791 9984
rect 18811 9970 18846 9984
rect 18866 9970 18875 9990
rect 18811 9962 18875 9970
rect 18837 9961 18875 9962
rect 18838 9960 18875 9961
rect 18941 9994 18977 9995
rect 19049 9994 19085 9995
rect 18941 9986 19085 9994
rect 18941 9966 18949 9986
rect 18969 9966 19057 9986
rect 19077 9966 19085 9986
rect 18941 9960 19085 9966
rect 19151 9990 19189 9998
rect 19257 9994 19293 9995
rect 19151 9970 19160 9990
rect 19180 9970 19189 9990
rect 19151 9961 19189 9970
rect 19208 9987 19293 9994
rect 19208 9967 19215 9987
rect 19236 9986 19293 9987
rect 19236 9967 19265 9986
rect 19208 9966 19265 9967
rect 19285 9966 19293 9986
rect 19151 9960 19188 9961
rect 19208 9960 19293 9966
rect 19359 9990 19397 9998
rect 19470 9994 19506 9995
rect 19359 9970 19368 9990
rect 19388 9970 19397 9990
rect 19359 9961 19397 9970
rect 19421 9986 19506 9994
rect 19421 9966 19478 9986
rect 19498 9966 19506 9986
rect 19359 9960 19396 9961
rect 19421 9960 19506 9966
rect 19572 9990 19610 9998
rect 19572 9970 19581 9990
rect 19601 9970 19610 9990
rect 19572 9961 19610 9970
rect 19650 9975 19722 10185
rect 19792 10219 20992 10249
rect 19792 10218 20236 10219
rect 19792 10216 19960 10218
rect 19650 9961 19733 9975
rect 19572 9960 19609 9961
rect 18995 9939 19031 9960
rect 19421 9939 19452 9960
rect 19650 9939 19667 9961
rect 18828 9935 18928 9939
rect 18828 9931 18890 9935
rect 18828 9905 18835 9931
rect 18861 9909 18890 9931
rect 18916 9909 18928 9935
rect 18861 9905 18928 9909
rect 18828 9902 18928 9905
rect 18996 9902 19031 9939
rect 19093 9936 19452 9939
rect 19093 9931 19315 9936
rect 19093 9907 19106 9931
rect 19130 9912 19315 9931
rect 19339 9912 19452 9936
rect 19130 9907 19452 9912
rect 19093 9903 19452 9907
rect 19519 9931 19667 9939
rect 19519 9911 19530 9931
rect 19550 9928 19667 9931
rect 19720 9928 19733 9961
rect 19550 9911 19733 9928
rect 19519 9904 19733 9911
rect 19519 9903 19560 9904
rect 19650 9903 19733 9904
rect 18995 9877 19031 9902
rect 18843 9850 18880 9851
rect 18939 9850 18976 9851
rect 18995 9850 19002 9877
rect 18743 9841 18881 9850
rect 18743 9821 18852 9841
rect 18872 9821 18881 9841
rect 18743 9814 18881 9821
rect 18939 9847 19002 9850
rect 19023 9850 19031 9877
rect 19050 9850 19087 9851
rect 19023 9847 19087 9850
rect 18939 9841 19087 9847
rect 18939 9821 18948 9841
rect 18968 9821 19058 9841
rect 19078 9821 19087 9841
rect 18743 9812 18839 9814
rect 18939 9811 19087 9821
rect 19146 9841 19183 9851
rect 19258 9850 19295 9851
rect 19239 9848 19295 9850
rect 19146 9821 19154 9841
rect 19174 9821 19183 9841
rect 18995 9810 19031 9811
rect 18843 9679 18880 9680
rect 19146 9679 19183 9821
rect 19208 9841 19295 9848
rect 19208 9838 19266 9841
rect 19208 9818 19213 9838
rect 19234 9821 19266 9838
rect 19286 9821 19295 9841
rect 19234 9818 19295 9821
rect 19208 9811 19295 9818
rect 19354 9841 19391 9851
rect 19354 9821 19362 9841
rect 19382 9821 19391 9841
rect 19208 9810 19239 9811
rect 19354 9742 19391 9821
rect 19421 9850 19452 9903
rect 19658 9870 19672 9903
rect 19725 9870 19733 9903
rect 19658 9864 19733 9870
rect 19658 9859 19728 9864
rect 19471 9850 19508 9851
rect 19421 9841 19508 9850
rect 19421 9821 19479 9841
rect 19499 9821 19508 9841
rect 19421 9811 19508 9821
rect 19567 9841 19604 9851
rect 19792 9846 19819 10216
rect 19859 9986 19923 9998
rect 20199 9994 20236 10218
rect 20707 10199 20771 10201
rect 20703 10187 20771 10199
rect 20703 10154 20714 10187
rect 20754 10154 20771 10187
rect 20703 10144 20771 10154
rect 20464 10083 20575 10098
rect 20464 10081 20506 10083
rect 20464 10061 20471 10081
rect 20490 10061 20506 10081
rect 20464 10053 20506 10061
rect 20534 10081 20575 10083
rect 20534 10061 20548 10081
rect 20567 10061 20575 10081
rect 20534 10053 20575 10061
rect 20464 10047 20575 10053
rect 20407 10025 20656 10047
rect 20407 9994 20444 10025
rect 20620 10023 20656 10025
rect 20620 9994 20657 10023
rect 19859 9985 19894 9986
rect 19836 9980 19894 9985
rect 19836 9960 19839 9980
rect 19859 9966 19894 9980
rect 19914 9966 19923 9986
rect 19859 9958 19923 9966
rect 19885 9957 19923 9958
rect 19886 9956 19923 9957
rect 19989 9990 20025 9991
rect 20097 9990 20133 9991
rect 19989 9982 20133 9990
rect 19989 9962 19997 9982
rect 20017 9962 20105 9982
rect 20125 9962 20133 9982
rect 19989 9956 20133 9962
rect 20199 9986 20237 9994
rect 20305 9990 20341 9991
rect 20199 9966 20208 9986
rect 20228 9966 20237 9986
rect 20199 9957 20237 9966
rect 20256 9983 20341 9990
rect 20256 9963 20263 9983
rect 20284 9982 20341 9983
rect 20284 9963 20313 9982
rect 20256 9962 20313 9963
rect 20333 9962 20341 9982
rect 20199 9956 20236 9957
rect 20256 9956 20341 9962
rect 20407 9986 20445 9994
rect 20518 9990 20554 9991
rect 20407 9966 20416 9986
rect 20436 9966 20445 9986
rect 20407 9957 20445 9966
rect 20469 9982 20554 9990
rect 20469 9962 20526 9982
rect 20546 9962 20554 9982
rect 20407 9956 20444 9957
rect 20469 9956 20554 9962
rect 20620 9986 20658 9994
rect 20620 9966 20629 9986
rect 20649 9966 20658 9986
rect 20620 9957 20658 9966
rect 20707 9960 20771 10144
rect 20927 10018 20992 10219
rect 22226 10289 22291 10490
rect 22447 10364 22511 10548
rect 22560 10542 22598 10551
rect 22560 10522 22569 10542
rect 22589 10522 22598 10542
rect 22560 10514 22598 10522
rect 22664 10546 22749 10552
rect 22774 10551 22811 10552
rect 22664 10526 22672 10546
rect 22692 10526 22749 10546
rect 22664 10518 22749 10526
rect 22773 10542 22811 10551
rect 22773 10522 22782 10542
rect 22802 10522 22811 10542
rect 22664 10517 22700 10518
rect 22773 10514 22811 10522
rect 22877 10546 22962 10552
rect 22982 10551 23019 10552
rect 22877 10526 22885 10546
rect 22905 10545 22962 10546
rect 22905 10526 22934 10545
rect 22877 10525 22934 10526
rect 22955 10525 22962 10545
rect 22877 10518 22962 10525
rect 22981 10542 23019 10551
rect 22981 10522 22990 10542
rect 23010 10522 23019 10542
rect 22877 10517 22913 10518
rect 22981 10514 23019 10522
rect 23085 10546 23229 10552
rect 23085 10526 23093 10546
rect 23113 10526 23201 10546
rect 23221 10526 23229 10546
rect 23085 10518 23229 10526
rect 23085 10517 23121 10518
rect 23193 10517 23229 10518
rect 23295 10551 23332 10552
rect 23295 10550 23333 10551
rect 23295 10542 23359 10550
rect 23295 10522 23304 10542
rect 23324 10528 23359 10542
rect 23379 10528 23382 10548
rect 23324 10523 23382 10528
rect 23324 10522 23359 10523
rect 22561 10485 22598 10514
rect 22562 10483 22598 10485
rect 22774 10483 22811 10514
rect 22562 10461 22811 10483
rect 22643 10455 22754 10461
rect 22643 10447 22684 10455
rect 22643 10427 22651 10447
rect 22670 10427 22684 10447
rect 22643 10425 22684 10427
rect 22712 10447 22754 10455
rect 22712 10427 22728 10447
rect 22747 10427 22754 10447
rect 22712 10425 22754 10427
rect 22643 10410 22754 10425
rect 22447 10354 22515 10364
rect 22447 10321 22464 10354
rect 22504 10321 22515 10354
rect 22447 10309 22515 10321
rect 22447 10307 22511 10309
rect 22982 10290 23019 10514
rect 23295 10510 23359 10522
rect 23399 10292 23426 10662
rect 23614 10657 23651 10667
rect 23710 10687 23797 10697
rect 23710 10667 23719 10687
rect 23739 10667 23797 10687
rect 23710 10658 23797 10667
rect 23710 10657 23747 10658
rect 23490 10644 23560 10649
rect 23485 10638 23560 10644
rect 23485 10605 23493 10638
rect 23546 10605 23560 10638
rect 23766 10605 23797 10658
rect 23827 10687 23864 10766
rect 23979 10697 24010 10698
rect 23827 10667 23836 10687
rect 23856 10667 23864 10687
rect 23827 10657 23864 10667
rect 23923 10690 24010 10697
rect 23923 10687 23984 10690
rect 23923 10667 23932 10687
rect 23952 10670 23984 10687
rect 24005 10670 24010 10690
rect 23952 10667 24010 10670
rect 23923 10660 24010 10667
rect 24035 10687 24072 10829
rect 24338 10828 24375 10829
rect 24187 10697 24223 10698
rect 24035 10667 24044 10687
rect 24064 10667 24072 10687
rect 23923 10658 23979 10660
rect 23923 10657 23960 10658
rect 24035 10657 24072 10667
rect 24131 10687 24279 10697
rect 24379 10694 24475 10696
rect 24131 10667 24140 10687
rect 24160 10667 24250 10687
rect 24270 10667 24279 10687
rect 24131 10661 24279 10667
rect 24131 10658 24195 10661
rect 24131 10657 24168 10658
rect 24187 10631 24195 10658
rect 24216 10658 24279 10661
rect 24337 10687 24475 10694
rect 24337 10667 24346 10687
rect 24366 10667 24475 10687
rect 24337 10658 24475 10667
rect 24216 10631 24223 10658
rect 24242 10657 24279 10658
rect 24338 10657 24375 10658
rect 24187 10606 24223 10631
rect 23485 10604 23568 10605
rect 23658 10604 23699 10605
rect 23485 10597 23699 10604
rect 23485 10580 23668 10597
rect 23485 10547 23498 10580
rect 23551 10577 23668 10580
rect 23688 10577 23699 10597
rect 23551 10569 23699 10577
rect 23766 10601 24125 10605
rect 23766 10596 24088 10601
rect 23766 10572 23879 10596
rect 23903 10577 24088 10596
rect 24112 10577 24125 10601
rect 23903 10572 24125 10577
rect 23766 10569 24125 10572
rect 24187 10569 24222 10606
rect 24290 10603 24390 10606
rect 24290 10599 24357 10603
rect 24290 10573 24302 10599
rect 24328 10577 24357 10599
rect 24383 10577 24390 10603
rect 24328 10573 24390 10577
rect 24290 10569 24390 10573
rect 23551 10547 23568 10569
rect 23766 10548 23797 10569
rect 24187 10548 24223 10569
rect 23609 10547 23646 10548
rect 23485 10533 23568 10547
rect 23258 10290 23426 10292
rect 22982 10289 23426 10290
rect 22226 10259 23426 10289
rect 23496 10323 23568 10533
rect 23608 10538 23646 10547
rect 23608 10518 23617 10538
rect 23637 10518 23646 10538
rect 23608 10510 23646 10518
rect 23712 10542 23797 10548
rect 23822 10547 23859 10548
rect 23712 10522 23720 10542
rect 23740 10522 23797 10542
rect 23712 10514 23797 10522
rect 23821 10538 23859 10547
rect 23821 10518 23830 10538
rect 23850 10518 23859 10538
rect 23712 10513 23748 10514
rect 23821 10510 23859 10518
rect 23925 10542 24010 10548
rect 24030 10547 24067 10548
rect 23925 10522 23933 10542
rect 23953 10541 24010 10542
rect 23953 10522 23982 10541
rect 23925 10521 23982 10522
rect 24003 10521 24010 10541
rect 23925 10514 24010 10521
rect 24029 10538 24067 10547
rect 24029 10518 24038 10538
rect 24058 10518 24067 10538
rect 23925 10513 23961 10514
rect 24029 10510 24067 10518
rect 24133 10542 24277 10548
rect 24133 10522 24141 10542
rect 24161 10522 24249 10542
rect 24269 10522 24277 10542
rect 24133 10514 24277 10522
rect 24133 10513 24169 10514
rect 24241 10513 24277 10514
rect 24343 10547 24380 10548
rect 24343 10546 24381 10547
rect 24343 10538 24407 10546
rect 24343 10518 24352 10538
rect 24372 10524 24407 10538
rect 24427 10524 24430 10544
rect 24372 10519 24430 10524
rect 24372 10518 24407 10519
rect 23609 10481 23646 10510
rect 23610 10479 23646 10481
rect 23822 10479 23859 10510
rect 23610 10457 23859 10479
rect 23691 10451 23802 10457
rect 23691 10443 23732 10451
rect 23691 10423 23699 10443
rect 23718 10423 23732 10443
rect 23691 10421 23732 10423
rect 23760 10443 23802 10451
rect 23760 10423 23776 10443
rect 23795 10423 23802 10443
rect 23760 10421 23802 10423
rect 23691 10406 23802 10421
rect 23496 10284 23515 10323
rect 23560 10284 23568 10323
rect 23496 10267 23568 10284
rect 24030 10311 24067 10510
rect 24343 10506 24407 10518
rect 24030 10305 24071 10311
rect 24447 10307 24474 10658
rect 24603 10610 24674 11089
rect 24603 10526 24672 10610
rect 24306 10305 24474 10307
rect 24030 10279 24474 10305
rect 22226 10212 22291 10259
rect 22226 10194 22249 10212
rect 22267 10194 22291 10212
rect 23139 10239 23174 10241
rect 23139 10237 23243 10239
rect 24032 10237 24071 10279
rect 24306 10278 24474 10279
rect 23139 10230 24073 10237
rect 23139 10229 23190 10230
rect 23139 10209 23142 10229
rect 23167 10210 23190 10229
rect 23222 10210 24073 10230
rect 23167 10209 24073 10210
rect 23139 10202 24073 10209
rect 23412 10201 24073 10202
rect 22226 10173 22291 10194
rect 22503 10184 22543 10187
rect 22503 10180 23406 10184
rect 22503 10160 23380 10180
rect 23400 10160 23406 10180
rect 22503 10157 23406 10160
rect 22227 10113 22292 10133
rect 22227 10095 22251 10113
rect 22269 10095 22292 10113
rect 22227 10068 22292 10095
rect 22503 10068 22543 10157
rect 22987 10155 23403 10157
rect 22987 10154 23328 10155
rect 22644 10123 22754 10137
rect 22644 10120 22687 10123
rect 22644 10115 22648 10120
rect 22226 10033 22543 10068
rect 22566 10093 22648 10115
rect 22677 10093 22687 10120
rect 22715 10096 22722 10123
rect 22751 10115 22754 10123
rect 22751 10096 22816 10115
rect 22715 10093 22816 10096
rect 22566 10091 22816 10093
rect 20927 10000 20949 10018
rect 20967 10000 20992 10018
rect 20927 9981 20992 10000
rect 20620 9956 20657 9957
rect 20043 9935 20079 9956
rect 20469 9935 20500 9956
rect 20707 9951 20715 9960
rect 20704 9935 20715 9951
rect 19876 9931 19976 9935
rect 19876 9927 19938 9931
rect 19876 9901 19883 9927
rect 19909 9905 19938 9927
rect 19964 9905 19976 9931
rect 19909 9901 19976 9905
rect 19876 9898 19976 9901
rect 20044 9898 20079 9935
rect 20141 9932 20500 9935
rect 20141 9927 20363 9932
rect 20141 9903 20154 9927
rect 20178 9908 20363 9927
rect 20387 9908 20500 9932
rect 20178 9903 20500 9908
rect 20141 9899 20500 9903
rect 20567 9927 20715 9935
rect 20567 9907 20578 9927
rect 20598 9918 20715 9927
rect 20764 9951 20771 9960
rect 22227 9957 22292 10033
rect 22566 10012 22603 10091
rect 22644 10078 22754 10091
rect 22718 10022 22749 10023
rect 22566 9992 22575 10012
rect 22595 9992 22603 10012
rect 22566 9982 22603 9992
rect 22662 10012 22749 10022
rect 22662 9992 22671 10012
rect 22691 9992 22749 10012
rect 22662 9983 22749 9992
rect 22662 9982 22699 9983
rect 20764 9918 20772 9951
rect 22227 9939 22249 9957
rect 22267 9939 22292 9957
rect 20598 9907 20772 9918
rect 20567 9900 20772 9907
rect 20567 9899 20608 9900
rect 20043 9873 20079 9898
rect 19891 9846 19928 9847
rect 19987 9846 20024 9847
rect 20043 9846 20050 9873
rect 19567 9821 19575 9841
rect 19595 9821 19604 9841
rect 19421 9810 19452 9811
rect 19416 9742 19526 9755
rect 19567 9742 19604 9821
rect 19791 9837 19929 9846
rect 19791 9817 19900 9837
rect 19920 9817 19929 9837
rect 19791 9810 19929 9817
rect 19987 9843 20050 9846
rect 20071 9846 20079 9873
rect 20098 9846 20135 9847
rect 20071 9843 20135 9846
rect 19987 9837 20135 9843
rect 19987 9817 19996 9837
rect 20016 9817 20106 9837
rect 20126 9817 20135 9837
rect 19791 9808 19887 9810
rect 19987 9807 20135 9817
rect 20194 9837 20231 9847
rect 20306 9846 20343 9847
rect 20287 9844 20343 9846
rect 20194 9817 20202 9837
rect 20222 9817 20231 9837
rect 20043 9806 20079 9807
rect 19354 9740 19604 9742
rect 19354 9737 19455 9740
rect 19354 9718 19419 9737
rect 19416 9710 19419 9718
rect 19448 9710 19455 9737
rect 19483 9713 19493 9740
rect 19522 9718 19604 9740
rect 19522 9713 19526 9718
rect 19483 9710 19526 9713
rect 19416 9696 19526 9710
rect 18842 9678 19183 9679
rect 18767 9673 19183 9678
rect 19891 9675 19928 9676
rect 20194 9675 20231 9817
rect 20256 9837 20343 9844
rect 20256 9834 20314 9837
rect 20256 9814 20261 9834
rect 20282 9817 20314 9834
rect 20334 9817 20343 9837
rect 20282 9814 20343 9817
rect 20256 9807 20343 9814
rect 20402 9837 20439 9847
rect 20402 9817 20410 9837
rect 20430 9817 20439 9837
rect 20256 9806 20287 9807
rect 20402 9738 20439 9817
rect 20469 9846 20500 9899
rect 20704 9897 20772 9900
rect 20704 9855 20716 9897
rect 20765 9855 20772 9897
rect 20519 9846 20556 9847
rect 20469 9837 20556 9846
rect 20469 9817 20527 9837
rect 20547 9817 20556 9837
rect 20469 9807 20556 9817
rect 20615 9837 20652 9847
rect 20704 9842 20772 9855
rect 20927 9919 20992 9936
rect 20927 9901 20951 9919
rect 20969 9901 20992 9919
rect 22227 9918 22292 9939
rect 22440 9937 22505 9946
rect 20615 9817 20623 9837
rect 20643 9817 20652 9837
rect 20469 9806 20500 9807
rect 20464 9738 20574 9751
rect 20615 9738 20652 9817
rect 20927 9762 20992 9901
rect 22440 9900 22450 9937
rect 22490 9929 22505 9937
rect 22718 9930 22749 9983
rect 22779 10012 22816 10091
rect 22931 10022 22962 10023
rect 22779 9992 22788 10012
rect 22808 9992 22816 10012
rect 22779 9982 22816 9992
rect 22875 10015 22962 10022
rect 22875 10012 22936 10015
rect 22875 9992 22884 10012
rect 22904 9995 22936 10012
rect 22957 9995 22962 10015
rect 22904 9992 22962 9995
rect 22875 9985 22962 9992
rect 22987 10012 23024 10154
rect 23290 10153 23327 10154
rect 23139 10022 23175 10023
rect 22987 9992 22996 10012
rect 23016 9992 23024 10012
rect 22875 9983 22931 9985
rect 22875 9982 22912 9983
rect 22987 9982 23024 9992
rect 23083 10012 23231 10022
rect 23331 10019 23427 10021
rect 23083 9992 23092 10012
rect 23112 9992 23202 10012
rect 23222 9992 23231 10012
rect 23083 9986 23231 9992
rect 23083 9983 23147 9986
rect 23083 9982 23120 9983
rect 23139 9956 23147 9983
rect 23168 9983 23231 9986
rect 23289 10012 23427 10019
rect 23289 9992 23298 10012
rect 23318 9992 23427 10012
rect 24607 10010 24669 10526
rect 23289 9983 23427 9992
rect 23168 9956 23175 9983
rect 23194 9982 23231 9983
rect 23290 9982 23327 9983
rect 23139 9931 23175 9956
rect 22610 9929 22651 9930
rect 22490 9922 22651 9929
rect 22490 9902 22620 9922
rect 22640 9902 22651 9922
rect 22490 9900 22651 9902
rect 22440 9894 22651 9900
rect 22718 9926 23077 9930
rect 22718 9921 23040 9926
rect 22718 9897 22831 9921
rect 22855 9902 23040 9921
rect 23064 9902 23077 9926
rect 22855 9897 23077 9902
rect 22718 9894 23077 9897
rect 23139 9894 23174 9931
rect 23242 9928 23342 9931
rect 23242 9924 23309 9928
rect 23242 9898 23254 9924
rect 23280 9902 23309 9924
rect 23335 9902 23342 9928
rect 23280 9898 23342 9902
rect 23242 9894 23342 9898
rect 22440 9881 22507 9894
rect 20927 9756 20949 9762
rect 20402 9736 20652 9738
rect 20402 9733 20503 9736
rect 20402 9714 20467 9733
rect 20464 9706 20467 9714
rect 20496 9706 20503 9733
rect 20531 9709 20541 9736
rect 20570 9714 20652 9736
rect 20681 9744 20949 9756
rect 20967 9744 20992 9762
rect 20681 9721 20992 9744
rect 22232 9858 22288 9878
rect 22232 9840 22251 9858
rect 22269 9840 22288 9858
rect 22232 9727 22288 9840
rect 22440 9860 22454 9881
rect 22490 9860 22507 9881
rect 22718 9873 22749 9894
rect 23139 9873 23175 9894
rect 22561 9872 22598 9873
rect 22440 9853 22507 9860
rect 22560 9863 22598 9872
rect 20681 9720 20736 9721
rect 20570 9709 20574 9714
rect 20531 9706 20574 9709
rect 20464 9692 20574 9706
rect 19890 9674 20231 9675
rect 18767 9653 18770 9673
rect 18790 9653 19183 9673
rect 19815 9673 20231 9674
rect 20681 9673 20724 9720
rect 19815 9669 20724 9673
rect 19134 9620 19179 9653
rect 19815 9649 19818 9669
rect 19838 9649 20724 9669
rect 20192 9644 20724 9649
rect 20932 9663 20991 9685
rect 20932 9645 20951 9663
rect 20969 9645 20991 9663
rect 19980 9620 20079 9622
rect 19134 9610 20079 9620
rect 19134 9584 20002 9610
rect 19135 9583 20002 9584
rect 19980 9572 20002 9583
rect 20027 9575 20046 9610
rect 20071 9575 20079 9610
rect 20027 9572 20079 9575
rect 20932 9574 20991 9645
rect 22232 9589 22287 9727
rect 22440 9701 22505 9853
rect 22560 9843 22569 9863
rect 22589 9843 22598 9863
rect 22560 9835 22598 9843
rect 22664 9867 22749 9873
rect 22774 9872 22811 9873
rect 22664 9847 22672 9867
rect 22692 9847 22749 9867
rect 22664 9839 22749 9847
rect 22773 9863 22811 9872
rect 22773 9843 22782 9863
rect 22802 9843 22811 9863
rect 22664 9838 22700 9839
rect 22773 9835 22811 9843
rect 22877 9867 22962 9873
rect 22982 9872 23019 9873
rect 22877 9847 22885 9867
rect 22905 9866 22962 9867
rect 22905 9847 22934 9866
rect 22877 9846 22934 9847
rect 22955 9846 22962 9866
rect 22877 9839 22962 9846
rect 22981 9863 23019 9872
rect 22981 9843 22990 9863
rect 23010 9843 23019 9863
rect 22877 9838 22913 9839
rect 22981 9835 23019 9843
rect 23085 9867 23229 9873
rect 23085 9847 23093 9867
rect 23113 9847 23201 9867
rect 23221 9847 23229 9867
rect 23085 9839 23229 9847
rect 23085 9838 23121 9839
rect 23193 9838 23229 9839
rect 23295 9872 23332 9873
rect 23295 9871 23333 9872
rect 23295 9863 23359 9871
rect 23295 9843 23304 9863
rect 23324 9849 23359 9863
rect 23379 9849 23382 9869
rect 23324 9844 23382 9849
rect 23324 9843 23359 9844
rect 22561 9806 22598 9835
rect 22562 9804 22598 9806
rect 22774 9804 22811 9835
rect 22562 9782 22811 9804
rect 22643 9776 22754 9782
rect 22643 9768 22684 9776
rect 22643 9748 22651 9768
rect 22670 9748 22684 9768
rect 22643 9746 22684 9748
rect 22712 9768 22754 9776
rect 22712 9748 22728 9768
rect 22747 9748 22754 9768
rect 22712 9746 22754 9748
rect 22643 9733 22754 9746
rect 22982 9736 23019 9835
rect 23295 9831 23359 9843
rect 22433 9691 22554 9701
rect 22433 9689 22502 9691
rect 22433 9648 22446 9689
rect 22483 9650 22502 9689
rect 22539 9650 22554 9691
rect 22483 9648 22554 9650
rect 22433 9630 22554 9648
rect 22225 9586 22289 9589
rect 22645 9586 22749 9592
rect 22980 9586 23021 9736
rect 23399 9728 23426 9983
rect 23488 9973 23568 9984
rect 23488 9947 23505 9973
rect 23545 9947 23568 9973
rect 23488 9920 23568 9947
rect 23488 9894 23509 9920
rect 23549 9894 23568 9920
rect 23488 9875 23568 9894
rect 23488 9849 23512 9875
rect 23552 9849 23568 9875
rect 23488 9798 23568 9849
rect 24591 9975 24669 10010
rect 24591 9913 24673 9975
rect 24591 9890 24619 9913
rect 24645 9890 24673 9913
rect 24591 9870 24673 9890
rect 22225 9583 23021 9586
rect 23400 9597 23426 9728
rect 23400 9583 23428 9597
rect 19980 9564 20079 9572
rect 20006 9563 20078 9564
rect 19660 9537 19727 9556
rect 19660 9516 19677 9537
rect 18541 9338 18621 9380
rect 19658 9471 19677 9516
rect 19707 9516 19727 9537
rect 19707 9471 19728 9516
rect 20197 9513 20238 9515
rect 20469 9513 20573 9515
rect 20929 9513 20993 9574
rect 17602 9227 17638 9228
rect 17494 9219 17638 9227
rect 17494 9199 17502 9219
rect 17522 9199 17610 9219
rect 17630 9199 17638 9219
rect 17494 9193 17638 9199
rect 17704 9223 17742 9231
rect 17810 9227 17846 9228
rect 17704 9203 17713 9223
rect 17733 9203 17742 9223
rect 17704 9194 17742 9203
rect 17761 9220 17846 9227
rect 17761 9200 17768 9220
rect 17789 9219 17846 9220
rect 17789 9200 17818 9219
rect 17761 9199 17818 9200
rect 17838 9199 17846 9219
rect 17704 9193 17741 9194
rect 17761 9193 17846 9199
rect 17912 9223 17950 9231
rect 18023 9227 18059 9228
rect 17912 9203 17921 9223
rect 17941 9203 17950 9223
rect 17912 9194 17950 9203
rect 17974 9219 18059 9227
rect 17974 9199 18031 9219
rect 18051 9199 18059 9219
rect 17912 9193 17949 9194
rect 17974 9193 18059 9199
rect 18125 9223 18163 9231
rect 18125 9203 18134 9223
rect 18154 9203 18163 9223
rect 18125 9194 18163 9203
rect 18363 9211 18449 9247
rect 18125 9193 18162 9194
rect 17548 9172 17584 9193
rect 17974 9172 18005 9193
rect 18201 9172 18247 9176
rect 17381 9168 17481 9172
rect 17381 9164 17443 9168
rect 17381 9138 17388 9164
rect 17414 9142 17443 9164
rect 17469 9142 17481 9168
rect 17414 9138 17481 9142
rect 17381 9135 17481 9138
rect 17549 9135 17584 9172
rect 17646 9169 18005 9172
rect 17646 9164 17868 9169
rect 17646 9140 17659 9164
rect 17683 9145 17868 9164
rect 17892 9145 18005 9169
rect 17683 9140 18005 9145
rect 17646 9136 18005 9140
rect 18072 9164 18247 9172
rect 18072 9144 18083 9164
rect 18103 9144 18247 9164
rect 18363 9170 18380 9211
rect 18434 9170 18449 9211
rect 18363 9151 18449 9170
rect 18072 9137 18247 9144
rect 18072 9136 18113 9137
rect 17548 9110 17584 9135
rect 17396 9083 17433 9084
rect 17492 9083 17529 9084
rect 17548 9083 17555 9110
rect 17296 9074 17434 9083
rect 17296 9054 17405 9074
rect 17425 9054 17434 9074
rect 17296 9047 17434 9054
rect 17492 9080 17555 9083
rect 17576 9083 17584 9110
rect 17603 9083 17640 9084
rect 17576 9080 17640 9083
rect 17492 9074 17640 9080
rect 17492 9054 17501 9074
rect 17521 9054 17611 9074
rect 17631 9054 17640 9074
rect 17296 9045 17392 9047
rect 17492 9044 17640 9054
rect 17699 9074 17736 9084
rect 17811 9083 17848 9084
rect 17792 9081 17848 9083
rect 17699 9054 17707 9074
rect 17727 9054 17736 9074
rect 17548 9043 17584 9044
rect 17396 8912 17433 8913
rect 17699 8912 17736 9054
rect 17761 9074 17848 9081
rect 17761 9071 17819 9074
rect 17761 9051 17766 9071
rect 17787 9054 17819 9071
rect 17839 9054 17848 9074
rect 17787 9051 17848 9054
rect 17761 9044 17848 9051
rect 17907 9074 17944 9084
rect 17907 9054 17915 9074
rect 17935 9054 17944 9074
rect 17761 9043 17792 9044
rect 17907 8975 17944 9054
rect 17974 9083 18005 9136
rect 18024 9083 18061 9084
rect 17974 9074 18061 9083
rect 17974 9054 18032 9074
rect 18052 9054 18061 9074
rect 17974 9044 18061 9054
rect 18120 9074 18157 9084
rect 18120 9054 18128 9074
rect 18148 9054 18157 9074
rect 17974 9043 18005 9044
rect 17969 8975 18079 8988
rect 18120 8975 18157 9054
rect 18201 9054 18247 9137
rect 18541 9054 18616 9338
rect 19658 9263 19728 9471
rect 19790 9478 20993 9513
rect 22225 9548 23428 9583
rect 23490 9590 23560 9798
rect 22225 9487 22289 9548
rect 22645 9546 22749 9548
rect 22980 9546 23021 9548
rect 23490 9545 23511 9590
rect 23491 9524 23511 9545
rect 23541 9545 23560 9590
rect 23541 9524 23558 9545
rect 23491 9505 23558 9524
rect 23140 9497 23212 9498
rect 23139 9489 23238 9497
rect 19790 9464 19818 9478
rect 19792 9333 19818 9464
rect 20197 9475 20993 9478
rect 19650 9212 19730 9263
rect 19650 9186 19666 9212
rect 19706 9186 19730 9212
rect 19650 9167 19730 9186
rect 19650 9141 19669 9167
rect 19709 9141 19730 9167
rect 19650 9114 19730 9141
rect 19650 9088 19673 9114
rect 19713 9088 19730 9114
rect 19650 9077 19730 9088
rect 19792 9078 19819 9333
rect 20197 9325 20238 9475
rect 20469 9469 20573 9475
rect 20929 9472 20993 9475
rect 20664 9413 20785 9431
rect 20664 9411 20735 9413
rect 20664 9370 20679 9411
rect 20716 9372 20735 9411
rect 20772 9372 20785 9413
rect 20716 9370 20785 9372
rect 20664 9360 20785 9370
rect 19859 9218 19923 9230
rect 20199 9226 20236 9325
rect 20464 9315 20575 9328
rect 20464 9313 20506 9315
rect 20464 9293 20471 9313
rect 20490 9293 20506 9313
rect 20464 9285 20506 9293
rect 20534 9313 20575 9315
rect 20534 9293 20548 9313
rect 20567 9293 20575 9313
rect 20534 9285 20575 9293
rect 20464 9279 20575 9285
rect 20407 9257 20656 9279
rect 20407 9226 20444 9257
rect 20620 9255 20656 9257
rect 20620 9226 20657 9255
rect 19859 9217 19894 9218
rect 19836 9212 19894 9217
rect 19836 9192 19839 9212
rect 19859 9198 19894 9212
rect 19914 9198 19923 9218
rect 19859 9190 19923 9198
rect 19885 9189 19923 9190
rect 19886 9188 19923 9189
rect 19989 9222 20025 9223
rect 20097 9222 20133 9223
rect 19989 9214 20133 9222
rect 19989 9194 19997 9214
rect 20017 9194 20105 9214
rect 20125 9194 20133 9214
rect 19989 9188 20133 9194
rect 20199 9218 20237 9226
rect 20305 9222 20341 9223
rect 20199 9198 20208 9218
rect 20228 9198 20237 9218
rect 20199 9189 20237 9198
rect 20256 9215 20341 9222
rect 20256 9195 20263 9215
rect 20284 9214 20341 9215
rect 20284 9195 20313 9214
rect 20256 9194 20313 9195
rect 20333 9194 20341 9214
rect 20199 9188 20236 9189
rect 20256 9188 20341 9194
rect 20407 9218 20445 9226
rect 20518 9222 20554 9223
rect 20407 9198 20416 9218
rect 20436 9198 20445 9218
rect 20407 9189 20445 9198
rect 20469 9214 20554 9222
rect 20469 9194 20526 9214
rect 20546 9194 20554 9214
rect 20407 9188 20444 9189
rect 20469 9188 20554 9194
rect 20620 9218 20658 9226
rect 20620 9198 20629 9218
rect 20649 9198 20658 9218
rect 20713 9208 20778 9360
rect 20931 9334 20986 9472
rect 22227 9416 22286 9487
rect 23139 9486 23191 9489
rect 23139 9451 23147 9486
rect 23172 9451 23191 9486
rect 23216 9478 23238 9489
rect 23216 9477 24083 9478
rect 23216 9451 24084 9477
rect 23139 9441 24084 9451
rect 23139 9439 23238 9441
rect 22227 9398 22249 9416
rect 22267 9398 22286 9416
rect 22227 9376 22286 9398
rect 22494 9412 23026 9417
rect 22494 9392 23380 9412
rect 23400 9392 23403 9412
rect 24039 9408 24084 9441
rect 22494 9388 23403 9392
rect 22494 9341 22537 9388
rect 22987 9387 23403 9388
rect 24035 9388 24428 9408
rect 24448 9388 24451 9408
rect 22987 9386 23328 9387
rect 22644 9355 22754 9369
rect 22644 9352 22687 9355
rect 22644 9347 22648 9352
rect 22482 9340 22537 9341
rect 20620 9189 20658 9198
rect 20711 9201 20778 9208
rect 20620 9188 20657 9189
rect 20043 9167 20079 9188
rect 20469 9167 20500 9188
rect 20711 9180 20728 9201
rect 20764 9180 20778 9201
rect 20930 9221 20986 9334
rect 20930 9203 20949 9221
rect 20967 9203 20986 9221
rect 20930 9183 20986 9203
rect 22226 9317 22537 9340
rect 22226 9299 22251 9317
rect 22269 9305 22537 9317
rect 22566 9325 22648 9347
rect 22677 9325 22687 9352
rect 22715 9328 22722 9355
rect 22751 9347 22754 9355
rect 22751 9328 22816 9347
rect 22715 9325 22816 9328
rect 22566 9323 22816 9325
rect 22269 9299 22291 9305
rect 20711 9167 20778 9180
rect 19876 9163 19976 9167
rect 19876 9159 19938 9163
rect 19876 9133 19883 9159
rect 19909 9137 19938 9159
rect 19964 9137 19976 9163
rect 19909 9133 19976 9137
rect 19876 9130 19976 9133
rect 20044 9130 20079 9167
rect 20141 9164 20500 9167
rect 20141 9159 20363 9164
rect 20141 9135 20154 9159
rect 20178 9140 20363 9159
rect 20387 9140 20500 9164
rect 20178 9135 20500 9140
rect 20141 9131 20500 9135
rect 20567 9161 20778 9167
rect 20567 9159 20728 9161
rect 20567 9139 20578 9159
rect 20598 9139 20728 9159
rect 20567 9132 20728 9139
rect 20567 9131 20608 9132
rect 20043 9105 20079 9130
rect 19891 9078 19928 9079
rect 19987 9078 20024 9079
rect 20043 9078 20050 9105
rect 18201 9019 18616 9054
rect 19791 9069 19929 9078
rect 19791 9049 19900 9069
rect 19920 9049 19929 9069
rect 19791 9042 19929 9049
rect 19987 9075 20050 9078
rect 20071 9078 20079 9105
rect 20098 9078 20135 9079
rect 20071 9075 20135 9078
rect 19987 9069 20135 9075
rect 19987 9049 19996 9069
rect 20016 9049 20106 9069
rect 20126 9049 20135 9069
rect 19791 9040 19887 9042
rect 19987 9039 20135 9049
rect 20194 9069 20231 9079
rect 20306 9078 20343 9079
rect 20287 9076 20343 9078
rect 20194 9049 20202 9069
rect 20222 9049 20231 9069
rect 20043 9038 20079 9039
rect 18201 9018 18247 9019
rect 17907 8973 18157 8975
rect 17907 8970 18008 8973
rect 17907 8951 17972 8970
rect 17969 8943 17972 8951
rect 18001 8943 18008 8970
rect 18036 8946 18046 8973
rect 18075 8951 18157 8973
rect 18541 8967 18616 9019
rect 18075 8946 18079 8951
rect 18036 8943 18079 8946
rect 17969 8929 18079 8943
rect 17395 8911 17736 8912
rect 17320 8906 17736 8911
rect 17320 8886 17323 8906
rect 17343 8886 17737 8906
rect 16377 8239 17183 8314
rect 15616 8195 15625 8229
rect 15654 8228 16064 8229
rect 15654 8195 15671 8228
rect 15896 8227 16064 8228
rect 15616 8169 15671 8195
rect 15616 8135 15624 8169
rect 15653 8135 15671 8169
rect 15616 8123 15671 8135
rect 13812 8078 13896 8099
rect 13812 8050 13840 8078
rect 13884 8050 13896 8078
rect 13626 7999 13700 8027
rect 13626 7951 13649 7999
rect 13686 7951 13700 7999
rect 13812 8021 13896 8050
rect 13812 7993 13837 8021
rect 13881 7993 13896 8021
rect 13812 7968 13896 7993
rect 15952 7982 16040 7986
rect 13626 7942 13700 7951
rect 8946 7875 9018 7897
rect 9079 7890 10282 7925
rect 9079 7876 9107 7890
rect 8947 7675 9017 7875
rect 9081 7745 9107 7876
rect 9486 7887 10282 7890
rect 8939 7624 9019 7675
rect 8939 7598 8955 7624
rect 8995 7598 9019 7624
rect 8939 7579 9019 7598
rect 8939 7553 8958 7579
rect 8998 7553 9019 7579
rect 8939 7526 9019 7553
rect 8939 7500 8962 7526
rect 9002 7500 9019 7526
rect 8939 7489 9019 7500
rect 9081 7490 9108 7745
rect 9486 7737 9527 7887
rect 9758 7885 9862 7887
rect 10217 7853 10282 7887
rect 11259 7892 11325 7940
rect 13636 7938 13700 7942
rect 15952 7965 16216 7982
rect 15952 7911 16132 7965
rect 16195 7911 16216 7965
rect 13849 7901 14560 7903
rect 13222 7900 14560 7901
rect 12172 7899 12244 7900
rect 9953 7825 10074 7843
rect 9953 7823 10024 7825
rect 9953 7782 9968 7823
rect 10005 7784 10024 7823
rect 10061 7784 10074 7825
rect 10005 7782 10074 7784
rect 9953 7772 10074 7782
rect 9758 7742 9862 7745
rect 9148 7630 9212 7642
rect 9488 7638 9525 7737
rect 9753 7727 9864 7742
rect 9753 7725 9795 7727
rect 9753 7705 9760 7725
rect 9779 7705 9795 7725
rect 9753 7697 9795 7705
rect 9823 7725 9864 7727
rect 9823 7705 9837 7725
rect 9856 7705 9864 7725
rect 9823 7697 9864 7705
rect 9753 7691 9864 7697
rect 9696 7669 9945 7691
rect 9696 7638 9733 7669
rect 9909 7667 9945 7669
rect 9909 7638 9946 7667
rect 9148 7629 9183 7630
rect 9125 7624 9183 7629
rect 9125 7604 9128 7624
rect 9148 7610 9183 7624
rect 9203 7610 9212 7630
rect 9148 7602 9212 7610
rect 9174 7601 9212 7602
rect 9175 7600 9212 7601
rect 9278 7634 9314 7635
rect 9386 7634 9422 7635
rect 9278 7626 9422 7634
rect 9278 7606 9286 7626
rect 9306 7606 9394 7626
rect 9414 7606 9422 7626
rect 9278 7600 9422 7606
rect 9488 7630 9526 7638
rect 9594 7634 9630 7635
rect 9488 7610 9497 7630
rect 9517 7610 9526 7630
rect 9488 7601 9526 7610
rect 9545 7627 9630 7634
rect 9545 7607 9552 7627
rect 9573 7626 9630 7627
rect 9573 7607 9602 7626
rect 9545 7606 9602 7607
rect 9622 7606 9630 7626
rect 9488 7600 9525 7601
rect 9545 7600 9630 7606
rect 9696 7630 9734 7638
rect 9807 7634 9843 7635
rect 9696 7610 9705 7630
rect 9725 7610 9734 7630
rect 9696 7601 9734 7610
rect 9758 7626 9843 7634
rect 9758 7606 9815 7626
rect 9835 7606 9843 7626
rect 9696 7600 9733 7601
rect 9758 7600 9843 7606
rect 9909 7630 9947 7638
rect 9909 7610 9918 7630
rect 9938 7610 9947 7630
rect 10002 7620 10067 7772
rect 10220 7746 10275 7853
rect 11259 7818 11318 7892
rect 12171 7891 12270 7899
rect 12171 7888 12223 7891
rect 12171 7853 12179 7888
rect 12204 7853 12223 7888
rect 12248 7880 12270 7891
rect 13221 7892 14560 7900
rect 13221 7889 13273 7892
rect 12248 7879 13115 7880
rect 12248 7853 13116 7879
rect 12171 7843 13116 7853
rect 12171 7841 12270 7843
rect 11259 7800 11281 7818
rect 11299 7800 11318 7818
rect 11259 7778 11318 7800
rect 11526 7814 12058 7819
rect 11526 7794 12412 7814
rect 12432 7794 12435 7814
rect 13071 7810 13116 7843
rect 13221 7854 13229 7889
rect 13254 7854 13273 7889
rect 13298 7854 14560 7892
rect 13221 7845 14560 7854
rect 13221 7842 13310 7845
rect 13849 7843 14560 7845
rect 15952 7894 16216 7911
rect 11526 7790 12435 7794
rect 9909 7601 9947 7610
rect 10000 7613 10067 7620
rect 9909 7600 9946 7601
rect 9332 7579 9368 7600
rect 9758 7579 9789 7600
rect 10000 7592 10017 7613
rect 10053 7592 10067 7613
rect 10219 7633 10275 7746
rect 11526 7743 11569 7790
rect 12019 7789 12435 7790
rect 13067 7790 13460 7810
rect 13480 7790 13483 7810
rect 12019 7788 12360 7789
rect 11676 7757 11786 7771
rect 11676 7754 11719 7757
rect 11676 7749 11680 7754
rect 11514 7742 11569 7743
rect 10219 7615 10238 7633
rect 10256 7615 10275 7633
rect 10219 7595 10275 7615
rect 11258 7719 11569 7742
rect 11258 7701 11283 7719
rect 11301 7707 11569 7719
rect 11598 7727 11680 7749
rect 11709 7727 11719 7754
rect 11747 7730 11754 7757
rect 11783 7749 11786 7757
rect 11783 7730 11848 7749
rect 11747 7727 11848 7730
rect 11598 7725 11848 7727
rect 11301 7701 11323 7707
rect 10000 7579 10067 7592
rect 9165 7575 9265 7579
rect 9165 7571 9227 7575
rect 9165 7545 9172 7571
rect 9198 7549 9227 7571
rect 9253 7549 9265 7575
rect 9198 7545 9265 7549
rect 9165 7542 9265 7545
rect 9333 7542 9368 7579
rect 9430 7576 9789 7579
rect 9430 7571 9652 7576
rect 9430 7547 9443 7571
rect 9467 7552 9652 7571
rect 9676 7552 9789 7576
rect 9467 7547 9789 7552
rect 9430 7543 9789 7547
rect 9856 7573 10067 7579
rect 9856 7571 10017 7573
rect 9856 7551 9867 7571
rect 9887 7551 10017 7571
rect 9856 7544 10017 7551
rect 9856 7543 9897 7544
rect 9332 7517 9368 7542
rect 9180 7490 9217 7491
rect 9276 7490 9313 7491
rect 9332 7490 9339 7517
rect 9080 7481 9218 7490
rect 9080 7461 9189 7481
rect 9209 7461 9218 7481
rect 9080 7454 9218 7461
rect 9276 7487 9339 7490
rect 9360 7490 9368 7517
rect 9387 7490 9424 7491
rect 9360 7487 9424 7490
rect 9276 7481 9424 7487
rect 9276 7461 9285 7481
rect 9305 7461 9395 7481
rect 9415 7461 9424 7481
rect 9080 7452 9176 7454
rect 9276 7451 9424 7461
rect 9483 7481 9520 7491
rect 9595 7490 9632 7491
rect 9576 7488 9632 7490
rect 9483 7461 9491 7481
rect 9511 7461 9520 7481
rect 9332 7450 9368 7451
rect 9180 7319 9217 7320
rect 9483 7319 9520 7461
rect 9545 7481 9632 7488
rect 9545 7478 9603 7481
rect 9545 7458 9550 7478
rect 9571 7461 9603 7478
rect 9623 7461 9632 7481
rect 9571 7458 9632 7461
rect 9545 7451 9632 7458
rect 9691 7481 9728 7491
rect 9691 7461 9699 7481
rect 9719 7461 9728 7481
rect 9545 7450 9576 7451
rect 9691 7382 9728 7461
rect 9758 7490 9789 7543
rect 10002 7536 10017 7544
rect 10057 7536 10067 7573
rect 11258 7562 11323 7701
rect 11598 7646 11635 7725
rect 11676 7712 11786 7725
rect 11750 7656 11781 7657
rect 11598 7626 11607 7646
rect 11627 7626 11635 7646
rect 10002 7527 10067 7536
rect 10215 7534 10280 7555
rect 10215 7516 10240 7534
rect 10258 7516 10280 7534
rect 11258 7544 11281 7562
rect 11299 7544 11323 7562
rect 11258 7527 11323 7544
rect 11478 7608 11546 7621
rect 11598 7616 11635 7626
rect 11694 7646 11781 7656
rect 11694 7626 11703 7646
rect 11723 7626 11781 7646
rect 11694 7617 11781 7626
rect 11694 7616 11731 7617
rect 11478 7566 11485 7608
rect 11534 7566 11546 7608
rect 11478 7563 11546 7566
rect 11750 7564 11781 7617
rect 11811 7646 11848 7725
rect 11963 7656 11994 7657
rect 11811 7626 11820 7646
rect 11840 7626 11848 7646
rect 11811 7616 11848 7626
rect 11907 7649 11994 7656
rect 11907 7646 11968 7649
rect 11907 7626 11916 7646
rect 11936 7629 11968 7646
rect 11989 7629 11994 7649
rect 11936 7626 11994 7629
rect 11907 7619 11994 7626
rect 12019 7646 12056 7788
rect 12322 7787 12359 7788
rect 13067 7785 13483 7790
rect 13067 7784 13408 7785
rect 12724 7753 12834 7767
rect 12724 7750 12767 7753
rect 12724 7745 12728 7750
rect 12646 7723 12728 7745
rect 12757 7723 12767 7750
rect 12795 7726 12802 7753
rect 12831 7745 12834 7753
rect 12831 7726 12896 7745
rect 12795 7723 12896 7726
rect 12646 7721 12896 7723
rect 12171 7656 12207 7657
rect 12019 7626 12028 7646
rect 12048 7626 12056 7646
rect 11907 7617 11963 7619
rect 11907 7616 11944 7617
rect 12019 7616 12056 7626
rect 12115 7646 12263 7656
rect 12363 7653 12459 7655
rect 12115 7626 12124 7646
rect 12144 7626 12234 7646
rect 12254 7626 12263 7646
rect 12115 7620 12263 7626
rect 12115 7617 12179 7620
rect 12115 7616 12152 7617
rect 12171 7590 12179 7617
rect 12200 7617 12263 7620
rect 12321 7646 12459 7653
rect 12321 7626 12330 7646
rect 12350 7626 12459 7646
rect 12321 7617 12459 7626
rect 12646 7642 12683 7721
rect 12724 7708 12834 7721
rect 12798 7652 12829 7653
rect 12646 7622 12655 7642
rect 12675 7622 12683 7642
rect 12200 7590 12207 7617
rect 12226 7616 12263 7617
rect 12322 7616 12359 7617
rect 12171 7565 12207 7590
rect 11642 7563 11683 7564
rect 11478 7556 11683 7563
rect 11478 7545 11652 7556
rect 9808 7490 9845 7491
rect 9758 7481 9845 7490
rect 9758 7461 9816 7481
rect 9836 7461 9845 7481
rect 9758 7451 9845 7461
rect 9904 7481 9941 7491
rect 9904 7461 9912 7481
rect 9932 7461 9941 7481
rect 9758 7450 9789 7451
rect 9753 7382 9863 7395
rect 9904 7382 9941 7461
rect 10215 7440 10280 7516
rect 11478 7512 11486 7545
rect 11479 7503 11486 7512
rect 11535 7536 11652 7545
rect 11672 7536 11683 7556
rect 11535 7528 11683 7536
rect 11750 7560 12109 7564
rect 11750 7555 12072 7560
rect 11750 7531 11863 7555
rect 11887 7536 12072 7555
rect 12096 7536 12109 7560
rect 11887 7531 12109 7536
rect 11750 7528 12109 7531
rect 12171 7528 12206 7565
rect 12274 7562 12374 7565
rect 12274 7558 12341 7562
rect 12274 7532 12286 7558
rect 12312 7536 12341 7558
rect 12367 7536 12374 7562
rect 12312 7532 12374 7536
rect 12274 7528 12374 7532
rect 11535 7512 11546 7528
rect 11535 7503 11543 7512
rect 11750 7507 11781 7528
rect 12171 7507 12207 7528
rect 11593 7506 11630 7507
rect 11258 7463 11323 7482
rect 11258 7445 11283 7463
rect 11301 7445 11323 7463
rect 9691 7380 9941 7382
rect 9691 7377 9792 7380
rect 9691 7358 9756 7377
rect 9753 7350 9756 7358
rect 9785 7350 9792 7377
rect 9820 7353 9830 7380
rect 9859 7358 9941 7380
rect 9964 7405 10281 7440
rect 9859 7353 9863 7358
rect 9820 7350 9863 7353
rect 9753 7336 9863 7350
rect 9179 7318 9520 7319
rect 9104 7316 9520 7318
rect 9964 7316 10004 7405
rect 10215 7378 10280 7405
rect 10215 7360 10238 7378
rect 10256 7360 10280 7378
rect 10215 7340 10280 7360
rect 9101 7313 10004 7316
rect 9101 7293 9107 7313
rect 9127 7293 10004 7313
rect 9101 7289 10004 7293
rect 9964 7286 10004 7289
rect 10216 7279 10281 7300
rect 8434 7271 9095 7272
rect 8434 7264 9368 7271
rect 8434 7263 9340 7264
rect 8434 7243 9285 7263
rect 9317 7244 9340 7263
rect 9365 7244 9368 7264
rect 9317 7243 9368 7244
rect 8434 7236 9368 7243
rect 8033 7194 8201 7195
rect 8436 7194 8475 7236
rect 9264 7234 9368 7236
rect 9333 7232 9368 7234
rect 10216 7261 10240 7279
rect 10258 7261 10281 7279
rect 10216 7214 10281 7261
rect 8033 7168 8477 7194
rect 8033 7166 8201 7168
rect 8033 6815 8060 7166
rect 8436 7162 8477 7168
rect 8100 6955 8164 6967
rect 8440 6963 8477 7162
rect 8939 7189 9011 7206
rect 8939 7150 8947 7189
rect 8992 7150 9011 7189
rect 8705 7052 8816 7067
rect 8705 7050 8747 7052
rect 8705 7030 8712 7050
rect 8731 7030 8747 7050
rect 8705 7022 8747 7030
rect 8775 7050 8816 7052
rect 8775 7030 8789 7050
rect 8808 7030 8816 7050
rect 8775 7022 8816 7030
rect 8705 7016 8816 7022
rect 8648 6994 8897 7016
rect 8648 6963 8685 6994
rect 8861 6992 8897 6994
rect 8861 6963 8898 6992
rect 8100 6954 8135 6955
rect 8077 6949 8135 6954
rect 8077 6929 8080 6949
rect 8100 6935 8135 6949
rect 8155 6935 8164 6955
rect 8100 6927 8164 6935
rect 8126 6926 8164 6927
rect 8127 6925 8164 6926
rect 8230 6959 8266 6960
rect 8338 6959 8374 6960
rect 8230 6951 8374 6959
rect 8230 6931 8238 6951
rect 8258 6931 8346 6951
rect 8366 6931 8374 6951
rect 8230 6925 8374 6931
rect 8440 6955 8478 6963
rect 8546 6959 8582 6960
rect 8440 6935 8449 6955
rect 8469 6935 8478 6955
rect 8440 6926 8478 6935
rect 8497 6952 8582 6959
rect 8497 6932 8504 6952
rect 8525 6951 8582 6952
rect 8525 6932 8554 6951
rect 8497 6931 8554 6932
rect 8574 6931 8582 6951
rect 8440 6925 8477 6926
rect 8497 6925 8582 6931
rect 8648 6955 8686 6963
rect 8759 6959 8795 6960
rect 8648 6935 8657 6955
rect 8677 6935 8686 6955
rect 8648 6926 8686 6935
rect 8710 6951 8795 6959
rect 8710 6931 8767 6951
rect 8787 6931 8795 6951
rect 8648 6925 8685 6926
rect 8710 6925 8795 6931
rect 8861 6955 8899 6963
rect 8861 6935 8870 6955
rect 8890 6935 8899 6955
rect 8861 6926 8899 6935
rect 8939 6940 9011 7150
rect 9081 7184 10281 7214
rect 9081 7183 9525 7184
rect 9081 7181 9249 7183
rect 8939 6926 9022 6940
rect 8861 6925 8898 6926
rect 8284 6904 8320 6925
rect 8710 6904 8741 6925
rect 8939 6904 8956 6926
rect 8117 6900 8217 6904
rect 8117 6896 8179 6900
rect 8117 6870 8124 6896
rect 8150 6874 8179 6896
rect 8205 6874 8217 6900
rect 8150 6870 8217 6874
rect 8117 6867 8217 6870
rect 8285 6867 8320 6904
rect 8382 6901 8741 6904
rect 8382 6896 8604 6901
rect 8382 6872 8395 6896
rect 8419 6877 8604 6896
rect 8628 6877 8741 6901
rect 8419 6872 8741 6877
rect 8382 6868 8741 6872
rect 8808 6896 8956 6904
rect 8808 6876 8819 6896
rect 8839 6893 8956 6896
rect 9009 6893 9022 6926
rect 8839 6876 9022 6893
rect 8808 6869 9022 6876
rect 8808 6868 8849 6869
rect 8939 6868 9022 6869
rect 8284 6842 8320 6867
rect 8132 6815 8169 6816
rect 8228 6815 8265 6816
rect 8284 6815 8291 6842
rect 8032 6806 8170 6815
rect 8032 6786 8141 6806
rect 8161 6786 8170 6806
rect 8032 6779 8170 6786
rect 8228 6812 8291 6815
rect 8312 6815 8320 6842
rect 8339 6815 8376 6816
rect 8312 6812 8376 6815
rect 8228 6806 8376 6812
rect 8228 6786 8237 6806
rect 8257 6786 8347 6806
rect 8367 6786 8376 6806
rect 8032 6777 8128 6779
rect 8228 6776 8376 6786
rect 8435 6806 8472 6816
rect 8547 6815 8584 6816
rect 8528 6813 8584 6815
rect 8435 6786 8443 6806
rect 8463 6786 8472 6806
rect 8284 6775 8320 6776
rect 8132 6644 8169 6645
rect 8435 6644 8472 6786
rect 8497 6806 8584 6813
rect 8497 6803 8555 6806
rect 8497 6783 8502 6803
rect 8523 6786 8555 6803
rect 8575 6786 8584 6806
rect 8523 6783 8584 6786
rect 8497 6776 8584 6783
rect 8643 6806 8680 6816
rect 8643 6786 8651 6806
rect 8671 6786 8680 6806
rect 8497 6775 8528 6776
rect 8643 6707 8680 6786
rect 8710 6815 8741 6868
rect 8947 6835 8961 6868
rect 9014 6835 9022 6868
rect 8947 6829 9022 6835
rect 8947 6824 9017 6829
rect 8760 6815 8797 6816
rect 8710 6806 8797 6815
rect 8710 6786 8768 6806
rect 8788 6786 8797 6806
rect 8710 6776 8797 6786
rect 8856 6806 8893 6816
rect 9081 6811 9108 7181
rect 9148 6951 9212 6963
rect 9488 6959 9525 7183
rect 9996 7164 10060 7166
rect 9992 7152 10060 7164
rect 9992 7119 10003 7152
rect 10043 7119 10060 7152
rect 9992 7109 10060 7119
rect 9753 7048 9864 7063
rect 9753 7046 9795 7048
rect 9753 7026 9760 7046
rect 9779 7026 9795 7046
rect 9753 7018 9795 7026
rect 9823 7046 9864 7048
rect 9823 7026 9837 7046
rect 9856 7026 9864 7046
rect 9823 7018 9864 7026
rect 9753 7012 9864 7018
rect 9696 6990 9945 7012
rect 9696 6959 9733 6990
rect 9909 6988 9945 6990
rect 9909 6959 9946 6988
rect 9148 6950 9183 6951
rect 9125 6945 9183 6950
rect 9125 6925 9128 6945
rect 9148 6931 9183 6945
rect 9203 6931 9212 6951
rect 9148 6923 9212 6931
rect 9174 6922 9212 6923
rect 9175 6921 9212 6922
rect 9278 6955 9314 6956
rect 9386 6955 9422 6956
rect 9278 6947 9422 6955
rect 9278 6927 9286 6947
rect 9306 6927 9394 6947
rect 9414 6927 9422 6947
rect 9278 6921 9422 6927
rect 9488 6951 9526 6959
rect 9594 6955 9630 6956
rect 9488 6931 9497 6951
rect 9517 6931 9526 6951
rect 9488 6922 9526 6931
rect 9545 6948 9630 6955
rect 9545 6928 9552 6948
rect 9573 6947 9630 6948
rect 9573 6928 9602 6947
rect 9545 6927 9602 6928
rect 9622 6927 9630 6947
rect 9488 6921 9525 6922
rect 9545 6921 9630 6927
rect 9696 6951 9734 6959
rect 9807 6955 9843 6956
rect 9696 6931 9705 6951
rect 9725 6931 9734 6951
rect 9696 6922 9734 6931
rect 9758 6947 9843 6955
rect 9758 6927 9815 6947
rect 9835 6927 9843 6947
rect 9696 6921 9733 6922
rect 9758 6921 9843 6927
rect 9909 6951 9947 6959
rect 9909 6931 9918 6951
rect 9938 6931 9947 6951
rect 9909 6922 9947 6931
rect 9996 6925 10060 7109
rect 10216 6983 10281 7184
rect 11258 7244 11323 7445
rect 11479 7319 11543 7503
rect 11592 7497 11630 7506
rect 11592 7477 11601 7497
rect 11621 7477 11630 7497
rect 11592 7469 11630 7477
rect 11696 7501 11781 7507
rect 11806 7506 11843 7507
rect 11696 7481 11704 7501
rect 11724 7481 11781 7501
rect 11696 7473 11781 7481
rect 11805 7497 11843 7506
rect 11805 7477 11814 7497
rect 11834 7477 11843 7497
rect 11696 7472 11732 7473
rect 11805 7469 11843 7477
rect 11909 7501 11994 7507
rect 12014 7506 12051 7507
rect 11909 7481 11917 7501
rect 11937 7500 11994 7501
rect 11937 7481 11966 7500
rect 11909 7480 11966 7481
rect 11987 7480 11994 7500
rect 11909 7473 11994 7480
rect 12013 7497 12051 7506
rect 12013 7477 12022 7497
rect 12042 7477 12051 7497
rect 11909 7472 11945 7473
rect 12013 7469 12051 7477
rect 12117 7501 12261 7507
rect 12117 7481 12125 7501
rect 12145 7481 12233 7501
rect 12253 7481 12261 7501
rect 12117 7473 12261 7481
rect 12117 7472 12153 7473
rect 12225 7472 12261 7473
rect 12327 7506 12364 7507
rect 12327 7505 12365 7506
rect 12327 7497 12391 7505
rect 12327 7477 12336 7497
rect 12356 7483 12391 7497
rect 12411 7483 12414 7503
rect 12356 7478 12414 7483
rect 12356 7477 12391 7478
rect 11593 7440 11630 7469
rect 11594 7438 11630 7440
rect 11806 7438 11843 7469
rect 11594 7416 11843 7438
rect 11675 7410 11786 7416
rect 11675 7402 11716 7410
rect 11675 7382 11683 7402
rect 11702 7382 11716 7402
rect 11675 7380 11716 7382
rect 11744 7402 11786 7410
rect 11744 7382 11760 7402
rect 11779 7382 11786 7402
rect 11744 7380 11786 7382
rect 11675 7365 11786 7380
rect 11479 7309 11547 7319
rect 11479 7276 11496 7309
rect 11536 7276 11547 7309
rect 11479 7264 11547 7276
rect 11479 7262 11543 7264
rect 12014 7245 12051 7469
rect 12327 7465 12391 7477
rect 12431 7247 12458 7617
rect 12646 7612 12683 7622
rect 12742 7642 12829 7652
rect 12742 7622 12751 7642
rect 12771 7622 12829 7642
rect 12742 7613 12829 7622
rect 12742 7612 12779 7613
rect 12522 7599 12592 7604
rect 12517 7593 12592 7599
rect 12517 7560 12525 7593
rect 12578 7560 12592 7593
rect 12798 7560 12829 7613
rect 12859 7642 12896 7721
rect 13011 7652 13042 7653
rect 12859 7622 12868 7642
rect 12888 7622 12896 7642
rect 12859 7612 12896 7622
rect 12955 7645 13042 7652
rect 12955 7642 13016 7645
rect 12955 7622 12964 7642
rect 12984 7625 13016 7642
rect 13037 7625 13042 7645
rect 12984 7622 13042 7625
rect 12955 7615 13042 7622
rect 13067 7642 13104 7784
rect 13370 7783 13407 7784
rect 13219 7652 13255 7653
rect 13067 7622 13076 7642
rect 13096 7622 13104 7642
rect 12955 7613 13011 7615
rect 12955 7612 12992 7613
rect 13067 7612 13104 7622
rect 13163 7642 13311 7652
rect 13411 7649 13507 7651
rect 13163 7622 13172 7642
rect 13192 7622 13282 7642
rect 13302 7622 13311 7642
rect 13163 7616 13311 7622
rect 13163 7613 13227 7616
rect 13163 7612 13200 7613
rect 13219 7586 13227 7613
rect 13248 7613 13311 7616
rect 13369 7642 13507 7649
rect 13369 7622 13378 7642
rect 13398 7622 13507 7642
rect 13369 7613 13507 7622
rect 13248 7586 13255 7613
rect 13274 7612 13311 7613
rect 13370 7612 13407 7613
rect 13219 7561 13255 7586
rect 12517 7559 12600 7560
rect 12690 7559 12731 7560
rect 12517 7552 12731 7559
rect 12517 7535 12700 7552
rect 12517 7502 12530 7535
rect 12583 7532 12700 7535
rect 12720 7532 12731 7552
rect 12583 7524 12731 7532
rect 12798 7556 13157 7560
rect 12798 7551 13120 7556
rect 12798 7527 12911 7551
rect 12935 7532 13120 7551
rect 13144 7532 13157 7556
rect 12935 7527 13157 7532
rect 12798 7524 13157 7527
rect 13219 7524 13254 7561
rect 13322 7558 13422 7561
rect 13322 7554 13389 7558
rect 13322 7528 13334 7554
rect 13360 7532 13389 7554
rect 13415 7532 13422 7558
rect 13360 7528 13422 7532
rect 13322 7524 13422 7528
rect 12583 7502 12600 7524
rect 12798 7503 12829 7524
rect 13219 7503 13255 7524
rect 12641 7502 12678 7503
rect 12517 7488 12600 7502
rect 12290 7245 12458 7247
rect 12014 7244 12458 7245
rect 11258 7214 12458 7244
rect 12528 7278 12600 7488
rect 12640 7493 12678 7502
rect 12640 7473 12649 7493
rect 12669 7473 12678 7493
rect 12640 7465 12678 7473
rect 12744 7497 12829 7503
rect 12854 7502 12891 7503
rect 12744 7477 12752 7497
rect 12772 7477 12829 7497
rect 12744 7469 12829 7477
rect 12853 7493 12891 7502
rect 12853 7473 12862 7493
rect 12882 7473 12891 7493
rect 12744 7468 12780 7469
rect 12853 7465 12891 7473
rect 12957 7497 13042 7503
rect 13062 7502 13099 7503
rect 12957 7477 12965 7497
rect 12985 7496 13042 7497
rect 12985 7477 13014 7496
rect 12957 7476 13014 7477
rect 13035 7476 13042 7496
rect 12957 7469 13042 7476
rect 13061 7493 13099 7502
rect 13061 7473 13070 7493
rect 13090 7473 13099 7493
rect 12957 7468 12993 7469
rect 13061 7465 13099 7473
rect 13165 7497 13309 7503
rect 13165 7477 13173 7497
rect 13193 7477 13281 7497
rect 13301 7477 13309 7497
rect 13165 7469 13309 7477
rect 13165 7468 13201 7469
rect 13273 7468 13309 7469
rect 13375 7502 13412 7503
rect 13375 7501 13413 7502
rect 13375 7493 13439 7501
rect 13375 7473 13384 7493
rect 13404 7479 13439 7493
rect 13459 7479 13462 7499
rect 13404 7474 13462 7479
rect 13404 7473 13439 7474
rect 12641 7436 12678 7465
rect 12642 7434 12678 7436
rect 12854 7434 12891 7465
rect 12642 7412 12891 7434
rect 12723 7406 12834 7412
rect 12723 7398 12764 7406
rect 12723 7378 12731 7398
rect 12750 7378 12764 7398
rect 12723 7376 12764 7378
rect 12792 7398 12834 7406
rect 12792 7378 12808 7398
rect 12827 7378 12834 7398
rect 12792 7376 12834 7378
rect 12723 7361 12834 7376
rect 12528 7239 12547 7278
rect 12592 7239 12600 7278
rect 12528 7222 12600 7239
rect 13062 7266 13099 7465
rect 13375 7461 13439 7473
rect 13062 7260 13103 7266
rect 13479 7262 13506 7613
rect 13801 7600 13896 7626
rect 13637 7578 13701 7597
rect 13637 7539 13650 7578
rect 13684 7539 13701 7578
rect 13637 7520 13701 7539
rect 13338 7260 13506 7262
rect 13062 7234 13506 7260
rect 11258 7167 11323 7214
rect 11258 7149 11281 7167
rect 11299 7149 11323 7167
rect 12171 7194 12206 7196
rect 12171 7192 12275 7194
rect 13064 7192 13103 7234
rect 13338 7233 13506 7234
rect 12171 7185 13105 7192
rect 12171 7184 12222 7185
rect 12171 7164 12174 7184
rect 12199 7165 12222 7184
rect 12254 7165 13105 7185
rect 12199 7164 13105 7165
rect 12171 7157 13105 7164
rect 12444 7156 13105 7157
rect 11258 7128 11323 7149
rect 11535 7139 11575 7142
rect 11535 7135 12438 7139
rect 11535 7115 12412 7135
rect 12432 7115 12438 7135
rect 11535 7112 12438 7115
rect 11259 7068 11324 7088
rect 11259 7050 11283 7068
rect 11301 7050 11324 7068
rect 11259 7023 11324 7050
rect 11535 7023 11575 7112
rect 12019 7110 12435 7112
rect 12019 7109 12360 7110
rect 11676 7078 11786 7092
rect 11676 7075 11719 7078
rect 11676 7070 11680 7075
rect 11258 6988 11575 7023
rect 11598 7048 11680 7070
rect 11709 7048 11719 7075
rect 11747 7051 11754 7078
rect 11783 7070 11786 7078
rect 11783 7051 11848 7070
rect 11747 7048 11848 7051
rect 11598 7046 11848 7048
rect 10216 6965 10238 6983
rect 10256 6965 10281 6983
rect 10216 6946 10281 6965
rect 9909 6921 9946 6922
rect 9332 6900 9368 6921
rect 9758 6900 9789 6921
rect 9996 6916 10004 6925
rect 9993 6900 10004 6916
rect 9165 6896 9265 6900
rect 9165 6892 9227 6896
rect 9165 6866 9172 6892
rect 9198 6870 9227 6892
rect 9253 6870 9265 6896
rect 9198 6866 9265 6870
rect 9165 6863 9265 6866
rect 9333 6863 9368 6900
rect 9430 6897 9789 6900
rect 9430 6892 9652 6897
rect 9430 6868 9443 6892
rect 9467 6873 9652 6892
rect 9676 6873 9789 6897
rect 9467 6868 9789 6873
rect 9430 6864 9789 6868
rect 9856 6892 10004 6900
rect 9856 6872 9867 6892
rect 9887 6883 10004 6892
rect 10053 6916 10060 6925
rect 10053 6883 10061 6916
rect 11259 6912 11324 6988
rect 11598 6967 11635 7046
rect 11676 7033 11786 7046
rect 11750 6977 11781 6978
rect 11598 6947 11607 6967
rect 11627 6947 11635 6967
rect 11598 6937 11635 6947
rect 11694 6967 11781 6977
rect 11694 6947 11703 6967
rect 11723 6947 11781 6967
rect 11694 6938 11781 6947
rect 11694 6937 11731 6938
rect 9887 6872 10061 6883
rect 9856 6865 10061 6872
rect 9856 6864 9897 6865
rect 9332 6838 9368 6863
rect 9180 6811 9217 6812
rect 9276 6811 9313 6812
rect 9332 6811 9339 6838
rect 8856 6786 8864 6806
rect 8884 6786 8893 6806
rect 8710 6775 8741 6776
rect 8705 6707 8815 6720
rect 8856 6707 8893 6786
rect 9080 6802 9218 6811
rect 9080 6782 9189 6802
rect 9209 6782 9218 6802
rect 9080 6775 9218 6782
rect 9276 6808 9339 6811
rect 9360 6811 9368 6838
rect 9387 6811 9424 6812
rect 9360 6808 9424 6811
rect 9276 6802 9424 6808
rect 9276 6782 9285 6802
rect 9305 6782 9395 6802
rect 9415 6782 9424 6802
rect 9080 6773 9176 6775
rect 9276 6772 9424 6782
rect 9483 6802 9520 6812
rect 9595 6811 9632 6812
rect 9576 6809 9632 6811
rect 9483 6782 9491 6802
rect 9511 6782 9520 6802
rect 9332 6771 9368 6772
rect 8643 6705 8893 6707
rect 8643 6702 8744 6705
rect 8643 6683 8708 6702
rect 8705 6675 8708 6683
rect 8737 6675 8744 6702
rect 8772 6678 8782 6705
rect 8811 6683 8893 6705
rect 8811 6678 8815 6683
rect 8772 6675 8815 6678
rect 8705 6661 8815 6675
rect 8131 6643 8472 6644
rect 8056 6638 8472 6643
rect 9180 6640 9217 6641
rect 9483 6640 9520 6782
rect 9545 6802 9632 6809
rect 9545 6799 9603 6802
rect 9545 6779 9550 6799
rect 9571 6782 9603 6799
rect 9623 6782 9632 6802
rect 9571 6779 9632 6782
rect 9545 6772 9632 6779
rect 9691 6802 9728 6812
rect 9691 6782 9699 6802
rect 9719 6782 9728 6802
rect 9545 6771 9576 6772
rect 9691 6703 9728 6782
rect 9758 6811 9789 6864
rect 9993 6862 10061 6865
rect 9993 6820 10005 6862
rect 10054 6820 10061 6862
rect 9808 6811 9845 6812
rect 9758 6802 9845 6811
rect 9758 6782 9816 6802
rect 9836 6782 9845 6802
rect 9758 6772 9845 6782
rect 9904 6802 9941 6812
rect 9993 6807 10061 6820
rect 10216 6884 10281 6901
rect 10216 6866 10240 6884
rect 10258 6866 10281 6884
rect 11259 6894 11281 6912
rect 11299 6894 11324 6912
rect 11259 6873 11324 6894
rect 11472 6892 11537 6901
rect 9904 6782 9912 6802
rect 9932 6782 9941 6802
rect 9758 6771 9789 6772
rect 9753 6703 9863 6716
rect 9904 6703 9941 6782
rect 10216 6727 10281 6866
rect 11472 6855 11482 6892
rect 11522 6884 11537 6892
rect 11750 6885 11781 6938
rect 11811 6967 11848 7046
rect 11963 6977 11994 6978
rect 11811 6947 11820 6967
rect 11840 6947 11848 6967
rect 11811 6937 11848 6947
rect 11907 6970 11994 6977
rect 11907 6967 11968 6970
rect 11907 6947 11916 6967
rect 11936 6950 11968 6967
rect 11989 6950 11994 6970
rect 11936 6947 11994 6950
rect 11907 6940 11994 6947
rect 12019 6967 12056 7109
rect 12322 7108 12359 7109
rect 13639 7049 13701 7520
rect 13801 7559 13827 7600
rect 13863 7559 13896 7600
rect 13801 7263 13896 7559
rect 13801 7219 13816 7263
rect 13876 7219 13896 7263
rect 13801 7199 13896 7219
rect 14513 7130 14556 7843
rect 14513 7110 14907 7130
rect 14927 7110 14930 7130
rect 14514 7105 14930 7110
rect 14514 7104 14855 7105
rect 14171 7073 14281 7087
rect 14171 7070 14214 7073
rect 14171 7065 14175 7070
rect 13634 6997 13709 7049
rect 14093 7043 14175 7065
rect 14204 7043 14214 7070
rect 14242 7046 14249 7073
rect 14278 7065 14281 7073
rect 14278 7046 14343 7065
rect 14242 7043 14343 7046
rect 14093 7041 14343 7043
rect 14003 6997 14049 6998
rect 12171 6977 12207 6978
rect 12019 6947 12028 6967
rect 12048 6947 12056 6967
rect 11907 6938 11963 6940
rect 11907 6937 11944 6938
rect 12019 6937 12056 6947
rect 12115 6967 12263 6977
rect 12363 6974 12459 6976
rect 12115 6947 12124 6967
rect 12144 6947 12234 6967
rect 12254 6947 12263 6967
rect 12115 6941 12263 6947
rect 12115 6938 12179 6941
rect 12115 6937 12152 6938
rect 12171 6911 12179 6938
rect 12200 6938 12263 6941
rect 12321 6967 12459 6974
rect 12321 6947 12330 6967
rect 12350 6947 12459 6967
rect 12321 6938 12459 6947
rect 13634 6962 14049 6997
rect 12200 6911 12207 6938
rect 12226 6937 12263 6938
rect 12322 6937 12359 6938
rect 12171 6886 12207 6911
rect 11642 6884 11683 6885
rect 11522 6877 11683 6884
rect 11522 6857 11652 6877
rect 11672 6857 11683 6877
rect 11522 6855 11683 6857
rect 11472 6849 11683 6855
rect 11750 6881 12109 6885
rect 11750 6876 12072 6881
rect 11750 6852 11863 6876
rect 11887 6857 12072 6876
rect 12096 6857 12109 6881
rect 11887 6852 12109 6857
rect 11750 6849 12109 6852
rect 12171 6849 12206 6886
rect 12274 6883 12374 6886
rect 12274 6879 12341 6883
rect 12274 6853 12286 6879
rect 12312 6857 12341 6879
rect 12367 6857 12374 6883
rect 12312 6853 12374 6857
rect 12274 6849 12374 6853
rect 11472 6836 11539 6849
rect 10216 6721 10238 6727
rect 9691 6701 9941 6703
rect 9691 6698 9792 6701
rect 9691 6679 9756 6698
rect 9753 6671 9756 6679
rect 9785 6671 9792 6698
rect 9820 6674 9830 6701
rect 9859 6679 9941 6701
rect 9970 6709 10238 6721
rect 10256 6709 10281 6727
rect 9970 6686 10281 6709
rect 11264 6813 11320 6833
rect 11264 6795 11283 6813
rect 11301 6795 11320 6813
rect 9970 6685 10025 6686
rect 9859 6674 9863 6679
rect 9820 6671 9863 6674
rect 9753 6657 9863 6671
rect 9179 6639 9520 6640
rect 8056 6618 8059 6638
rect 8079 6618 8472 6638
rect 9104 6638 9520 6639
rect 9970 6638 10013 6685
rect 11264 6682 11320 6795
rect 11472 6815 11486 6836
rect 11522 6815 11539 6836
rect 11750 6828 11781 6849
rect 12171 6828 12207 6849
rect 11593 6827 11630 6828
rect 11472 6808 11539 6815
rect 11592 6818 11630 6827
rect 9104 6634 10013 6638
rect 8423 6585 8468 6618
rect 9104 6614 9107 6634
rect 9127 6614 10013 6634
rect 9481 6609 10013 6614
rect 10221 6628 10280 6650
rect 10221 6610 10240 6628
rect 10258 6610 10280 6628
rect 9269 6585 9368 6587
rect 8423 6575 9368 6585
rect 8423 6549 9291 6575
rect 8424 6548 9291 6549
rect 9269 6537 9291 6548
rect 9316 6540 9335 6575
rect 9360 6540 9368 6575
rect 9316 6537 9368 6540
rect 10221 6539 10280 6610
rect 11264 6544 11319 6682
rect 11472 6656 11537 6808
rect 11592 6798 11601 6818
rect 11621 6798 11630 6818
rect 11592 6790 11630 6798
rect 11696 6822 11781 6828
rect 11806 6827 11843 6828
rect 11696 6802 11704 6822
rect 11724 6802 11781 6822
rect 11696 6794 11781 6802
rect 11805 6818 11843 6827
rect 11805 6798 11814 6818
rect 11834 6798 11843 6818
rect 11696 6793 11732 6794
rect 11805 6790 11843 6798
rect 11909 6822 11994 6828
rect 12014 6827 12051 6828
rect 11909 6802 11917 6822
rect 11937 6821 11994 6822
rect 11937 6802 11966 6821
rect 11909 6801 11966 6802
rect 11987 6801 11994 6821
rect 11909 6794 11994 6801
rect 12013 6818 12051 6827
rect 12013 6798 12022 6818
rect 12042 6798 12051 6818
rect 11909 6793 11945 6794
rect 12013 6790 12051 6798
rect 12117 6822 12261 6828
rect 12117 6802 12125 6822
rect 12145 6802 12233 6822
rect 12253 6802 12261 6822
rect 12117 6794 12261 6802
rect 12117 6793 12153 6794
rect 12225 6793 12261 6794
rect 12327 6827 12364 6828
rect 12327 6826 12365 6827
rect 12327 6818 12391 6826
rect 12327 6798 12336 6818
rect 12356 6804 12391 6818
rect 12411 6804 12414 6824
rect 12356 6799 12414 6804
rect 12356 6798 12391 6799
rect 11593 6761 11630 6790
rect 11594 6759 11630 6761
rect 11806 6759 11843 6790
rect 11594 6737 11843 6759
rect 11675 6731 11786 6737
rect 11675 6723 11716 6731
rect 11675 6703 11683 6723
rect 11702 6703 11716 6723
rect 11675 6701 11716 6703
rect 11744 6723 11786 6731
rect 11744 6703 11760 6723
rect 11779 6703 11786 6723
rect 11744 6701 11786 6703
rect 11675 6688 11786 6701
rect 12014 6691 12051 6790
rect 12327 6786 12391 6798
rect 11465 6646 11586 6656
rect 11465 6644 11534 6646
rect 11465 6603 11478 6644
rect 11515 6605 11534 6644
rect 11571 6605 11586 6646
rect 11515 6603 11586 6605
rect 11465 6585 11586 6603
rect 11257 6541 11321 6544
rect 11677 6541 11781 6547
rect 12012 6541 12053 6691
rect 12431 6683 12458 6938
rect 12520 6928 12600 6939
rect 12520 6902 12537 6928
rect 12577 6902 12600 6928
rect 12520 6875 12600 6902
rect 12520 6849 12541 6875
rect 12581 6849 12600 6875
rect 12520 6830 12600 6849
rect 12520 6804 12544 6830
rect 12584 6804 12600 6830
rect 12520 6753 12600 6804
rect 9269 6529 9368 6537
rect 9295 6528 9367 6529
rect 8949 6502 9016 6521
rect 8949 6481 8966 6502
rect 8947 6436 8966 6481
rect 8996 6481 9016 6502
rect 8996 6436 9017 6481
rect 9486 6478 9527 6480
rect 9758 6478 9862 6480
rect 10218 6478 10282 6539
rect 8947 6228 9017 6436
rect 9079 6443 10282 6478
rect 9079 6429 9107 6443
rect 9081 6298 9107 6429
rect 9486 6440 10282 6443
rect 11257 6538 12053 6541
rect 12432 6552 12458 6683
rect 12432 6538 12460 6552
rect 11257 6503 12460 6538
rect 12522 6545 12592 6753
rect 13634 6678 13709 6962
rect 14003 6879 14049 6962
rect 14093 6962 14130 7041
rect 14171 7028 14281 7041
rect 14245 6972 14276 6973
rect 14093 6942 14102 6962
rect 14122 6942 14130 6962
rect 14093 6932 14130 6942
rect 14189 6962 14276 6972
rect 14189 6942 14198 6962
rect 14218 6942 14276 6962
rect 14189 6933 14276 6942
rect 14189 6932 14226 6933
rect 14245 6880 14276 6933
rect 14306 6962 14343 7041
rect 14458 6972 14489 6973
rect 14306 6942 14315 6962
rect 14335 6942 14343 6962
rect 14306 6932 14343 6942
rect 14402 6965 14489 6972
rect 14402 6962 14463 6965
rect 14402 6942 14411 6962
rect 14431 6945 14463 6962
rect 14484 6945 14489 6965
rect 14431 6942 14489 6945
rect 14402 6935 14489 6942
rect 14514 6962 14551 7104
rect 14817 7103 14854 7104
rect 14666 6972 14702 6973
rect 14514 6942 14523 6962
rect 14543 6942 14551 6962
rect 14402 6933 14458 6935
rect 14402 6932 14439 6933
rect 14514 6932 14551 6942
rect 14610 6962 14758 6972
rect 14858 6969 14954 6971
rect 14610 6942 14619 6962
rect 14639 6942 14729 6962
rect 14749 6942 14758 6962
rect 14610 6936 14758 6942
rect 14610 6933 14674 6936
rect 14610 6932 14647 6933
rect 14666 6906 14674 6933
rect 14695 6933 14758 6936
rect 14816 6962 14954 6969
rect 14816 6942 14825 6962
rect 14845 6942 14954 6962
rect 14816 6933 14954 6942
rect 14695 6906 14702 6933
rect 14721 6932 14758 6933
rect 14817 6932 14854 6933
rect 14666 6881 14702 6906
rect 14137 6879 14178 6880
rect 14003 6872 14178 6879
rect 13801 6846 13887 6865
rect 13801 6805 13816 6846
rect 13870 6805 13887 6846
rect 14003 6852 14147 6872
rect 14167 6852 14178 6872
rect 14003 6844 14178 6852
rect 14245 6876 14604 6880
rect 14245 6871 14567 6876
rect 14245 6847 14358 6871
rect 14382 6852 14567 6871
rect 14591 6852 14604 6876
rect 14382 6847 14604 6852
rect 14245 6844 14604 6847
rect 14666 6844 14701 6881
rect 14769 6878 14869 6881
rect 14769 6874 14836 6878
rect 14769 6848 14781 6874
rect 14807 6852 14836 6874
rect 14862 6852 14869 6878
rect 14807 6848 14869 6852
rect 14769 6844 14869 6848
rect 14003 6840 14049 6844
rect 14245 6823 14276 6844
rect 14666 6823 14702 6844
rect 14088 6822 14125 6823
rect 13801 6769 13887 6805
rect 14087 6813 14125 6822
rect 14087 6793 14096 6813
rect 14116 6793 14125 6813
rect 14087 6785 14125 6793
rect 14191 6817 14276 6823
rect 14301 6822 14338 6823
rect 14191 6797 14199 6817
rect 14219 6797 14276 6817
rect 14191 6789 14276 6797
rect 14300 6813 14338 6822
rect 14300 6793 14309 6813
rect 14329 6793 14338 6813
rect 14191 6788 14227 6789
rect 14300 6785 14338 6793
rect 14404 6817 14489 6823
rect 14509 6822 14546 6823
rect 14404 6797 14412 6817
rect 14432 6816 14489 6817
rect 14432 6797 14461 6816
rect 14404 6796 14461 6797
rect 14482 6796 14489 6816
rect 14404 6789 14489 6796
rect 14508 6813 14546 6822
rect 14508 6793 14517 6813
rect 14537 6793 14546 6813
rect 14404 6788 14440 6789
rect 14508 6785 14546 6793
rect 14612 6817 14756 6823
rect 14612 6797 14620 6817
rect 14640 6797 14728 6817
rect 14748 6797 14756 6817
rect 14612 6789 14756 6797
rect 14612 6788 14648 6789
rect 11257 6442 11321 6503
rect 11677 6501 11781 6503
rect 12012 6501 12053 6503
rect 12522 6500 12543 6545
rect 12523 6479 12543 6500
rect 12573 6500 12592 6545
rect 13629 6636 13709 6678
rect 12573 6479 12590 6500
rect 12523 6460 12590 6479
rect 12172 6452 12244 6453
rect 12171 6444 12270 6452
rect 7834 6136 7916 6156
rect 7834 6113 7862 6136
rect 7888 6113 7916 6136
rect 7834 6051 7916 6113
rect 7838 6016 7916 6051
rect 8939 6177 9019 6228
rect 8939 6151 8955 6177
rect 8995 6151 9019 6177
rect 8939 6132 9019 6151
rect 8939 6106 8958 6132
rect 8998 6106 9019 6132
rect 8939 6079 9019 6106
rect 8939 6053 8962 6079
rect 9002 6053 9019 6079
rect 8939 6042 9019 6053
rect 9081 6043 9108 6298
rect 9486 6290 9527 6440
rect 9758 6434 9862 6440
rect 10218 6437 10282 6440
rect 9953 6378 10074 6396
rect 9953 6376 10024 6378
rect 9953 6335 9968 6376
rect 10005 6337 10024 6376
rect 10061 6337 10074 6378
rect 10005 6335 10074 6337
rect 9953 6325 10074 6335
rect 9148 6183 9212 6195
rect 9488 6191 9525 6290
rect 9753 6280 9864 6293
rect 9753 6278 9795 6280
rect 9753 6258 9760 6278
rect 9779 6258 9795 6278
rect 9753 6250 9795 6258
rect 9823 6278 9864 6280
rect 9823 6258 9837 6278
rect 9856 6258 9864 6278
rect 9823 6250 9864 6258
rect 9753 6244 9864 6250
rect 9696 6222 9945 6244
rect 9696 6191 9733 6222
rect 9909 6220 9945 6222
rect 9909 6191 9946 6220
rect 9148 6182 9183 6183
rect 9125 6177 9183 6182
rect 9125 6157 9128 6177
rect 9148 6163 9183 6177
rect 9203 6163 9212 6183
rect 9148 6155 9212 6163
rect 9174 6154 9212 6155
rect 9175 6153 9212 6154
rect 9278 6187 9314 6188
rect 9386 6187 9422 6188
rect 9278 6179 9422 6187
rect 9278 6159 9286 6179
rect 9306 6159 9394 6179
rect 9414 6159 9422 6179
rect 9278 6153 9422 6159
rect 9488 6183 9526 6191
rect 9594 6187 9630 6188
rect 9488 6163 9497 6183
rect 9517 6163 9526 6183
rect 9488 6154 9526 6163
rect 9545 6180 9630 6187
rect 9545 6160 9552 6180
rect 9573 6179 9630 6180
rect 9573 6160 9602 6179
rect 9545 6159 9602 6160
rect 9622 6159 9630 6179
rect 9488 6153 9525 6154
rect 9545 6153 9630 6159
rect 9696 6183 9734 6191
rect 9807 6187 9843 6188
rect 9696 6163 9705 6183
rect 9725 6163 9734 6183
rect 9696 6154 9734 6163
rect 9758 6179 9843 6187
rect 9758 6159 9815 6179
rect 9835 6159 9843 6179
rect 9696 6153 9733 6154
rect 9758 6153 9843 6159
rect 9909 6183 9947 6191
rect 9909 6163 9918 6183
rect 9938 6163 9947 6183
rect 10002 6173 10067 6325
rect 10220 6299 10275 6437
rect 11259 6371 11318 6442
rect 12171 6441 12223 6444
rect 12171 6406 12179 6441
rect 12204 6406 12223 6441
rect 12248 6433 12270 6444
rect 12248 6432 13115 6433
rect 12248 6406 13116 6432
rect 12171 6396 13116 6406
rect 12171 6394 12270 6396
rect 11259 6353 11281 6371
rect 11299 6353 11318 6371
rect 11259 6331 11318 6353
rect 11526 6367 12058 6372
rect 11526 6347 12412 6367
rect 12432 6347 12435 6367
rect 13071 6363 13116 6396
rect 11526 6343 12435 6347
rect 9909 6154 9947 6163
rect 10000 6166 10067 6173
rect 9909 6153 9946 6154
rect 9332 6132 9368 6153
rect 9758 6132 9789 6153
rect 10000 6145 10017 6166
rect 10053 6145 10067 6166
rect 10219 6186 10275 6299
rect 11526 6296 11569 6343
rect 12019 6342 12435 6343
rect 13067 6343 13460 6363
rect 13480 6343 13483 6363
rect 12019 6341 12360 6342
rect 11676 6310 11786 6324
rect 11676 6307 11719 6310
rect 11676 6302 11680 6307
rect 11514 6295 11569 6296
rect 10219 6168 10238 6186
rect 10256 6168 10275 6186
rect 10219 6148 10275 6168
rect 11258 6272 11569 6295
rect 11258 6254 11283 6272
rect 11301 6260 11569 6272
rect 11598 6280 11680 6302
rect 11709 6280 11719 6307
rect 11747 6283 11754 6310
rect 11783 6302 11786 6310
rect 11783 6283 11848 6302
rect 11747 6280 11848 6283
rect 11598 6278 11848 6280
rect 11301 6254 11323 6260
rect 10000 6132 10067 6145
rect 9165 6128 9265 6132
rect 9165 6124 9227 6128
rect 9165 6098 9172 6124
rect 9198 6102 9227 6124
rect 9253 6102 9265 6128
rect 9198 6098 9265 6102
rect 9165 6095 9265 6098
rect 9333 6095 9368 6132
rect 9430 6129 9789 6132
rect 9430 6124 9652 6129
rect 9430 6100 9443 6124
rect 9467 6105 9652 6124
rect 9676 6105 9789 6129
rect 9467 6100 9789 6105
rect 9430 6096 9789 6100
rect 9856 6126 10067 6132
rect 9856 6124 10017 6126
rect 9856 6104 9867 6124
rect 9887 6104 10017 6124
rect 9856 6097 10017 6104
rect 9856 6096 9897 6097
rect 9332 6070 9368 6095
rect 9180 6043 9217 6044
rect 9276 6043 9313 6044
rect 9332 6043 9339 6070
rect 9080 6034 9218 6043
rect 7838 5500 7900 6016
rect 9080 6014 9189 6034
rect 9209 6014 9218 6034
rect 9080 6007 9218 6014
rect 9276 6040 9339 6043
rect 9360 6043 9368 6070
rect 9387 6043 9424 6044
rect 9360 6040 9424 6043
rect 9276 6034 9424 6040
rect 9276 6014 9285 6034
rect 9305 6014 9395 6034
rect 9415 6014 9424 6034
rect 9080 6005 9176 6007
rect 9276 6004 9424 6014
rect 9483 6034 9520 6044
rect 9595 6043 9632 6044
rect 9576 6041 9632 6043
rect 9483 6014 9491 6034
rect 9511 6014 9520 6034
rect 9332 6003 9368 6004
rect 9180 5872 9217 5873
rect 9483 5872 9520 6014
rect 9545 6034 9632 6041
rect 9545 6031 9603 6034
rect 9545 6011 9550 6031
rect 9571 6014 9603 6031
rect 9623 6014 9632 6034
rect 9571 6011 9632 6014
rect 9545 6004 9632 6011
rect 9691 6034 9728 6044
rect 9691 6014 9699 6034
rect 9719 6014 9728 6034
rect 9545 6003 9576 6004
rect 9691 5935 9728 6014
rect 9758 6043 9789 6096
rect 10002 6089 10017 6097
rect 10057 6089 10067 6126
rect 11258 6115 11323 6254
rect 11598 6199 11635 6278
rect 11676 6265 11786 6278
rect 11750 6209 11781 6210
rect 11598 6179 11607 6199
rect 11627 6179 11635 6199
rect 10002 6080 10067 6089
rect 10215 6087 10280 6108
rect 10215 6069 10240 6087
rect 10258 6069 10280 6087
rect 11258 6097 11281 6115
rect 11299 6097 11323 6115
rect 11258 6080 11323 6097
rect 11478 6161 11546 6174
rect 11598 6169 11635 6179
rect 11694 6199 11781 6209
rect 11694 6179 11703 6199
rect 11723 6179 11781 6199
rect 11694 6170 11781 6179
rect 11694 6169 11731 6170
rect 11478 6119 11485 6161
rect 11534 6119 11546 6161
rect 11478 6116 11546 6119
rect 11750 6117 11781 6170
rect 11811 6199 11848 6278
rect 11963 6209 11994 6210
rect 11811 6179 11820 6199
rect 11840 6179 11848 6199
rect 11811 6169 11848 6179
rect 11907 6202 11994 6209
rect 11907 6199 11968 6202
rect 11907 6179 11916 6199
rect 11936 6182 11968 6199
rect 11989 6182 11994 6202
rect 11936 6179 11994 6182
rect 11907 6172 11994 6179
rect 12019 6199 12056 6341
rect 12322 6340 12359 6341
rect 13067 6338 13483 6343
rect 13067 6337 13408 6338
rect 12724 6306 12834 6320
rect 12724 6303 12767 6306
rect 12724 6298 12728 6303
rect 12646 6276 12728 6298
rect 12757 6276 12767 6303
rect 12795 6279 12802 6306
rect 12831 6298 12834 6306
rect 12831 6279 12896 6298
rect 12795 6276 12896 6279
rect 12646 6274 12896 6276
rect 12171 6209 12207 6210
rect 12019 6179 12028 6199
rect 12048 6179 12056 6199
rect 11907 6170 11963 6172
rect 11907 6169 11944 6170
rect 12019 6169 12056 6179
rect 12115 6199 12263 6209
rect 12363 6206 12459 6208
rect 12115 6179 12124 6199
rect 12144 6179 12234 6199
rect 12254 6179 12263 6199
rect 12115 6173 12263 6179
rect 12115 6170 12179 6173
rect 12115 6169 12152 6170
rect 12171 6143 12179 6170
rect 12200 6170 12263 6173
rect 12321 6199 12459 6206
rect 12321 6179 12330 6199
rect 12350 6179 12459 6199
rect 12321 6170 12459 6179
rect 12646 6195 12683 6274
rect 12724 6261 12834 6274
rect 12798 6205 12829 6206
rect 12646 6175 12655 6195
rect 12675 6175 12683 6195
rect 12200 6143 12207 6170
rect 12226 6169 12263 6170
rect 12322 6169 12359 6170
rect 12171 6118 12207 6143
rect 11642 6116 11683 6117
rect 11478 6109 11683 6116
rect 11478 6098 11652 6109
rect 9808 6043 9845 6044
rect 9758 6034 9845 6043
rect 9758 6014 9816 6034
rect 9836 6014 9845 6034
rect 9758 6004 9845 6014
rect 9904 6034 9941 6044
rect 9904 6014 9912 6034
rect 9932 6014 9941 6034
rect 9758 6003 9789 6004
rect 9753 5935 9863 5948
rect 9904 5935 9941 6014
rect 10215 5993 10280 6069
rect 11478 6065 11486 6098
rect 11479 6056 11486 6065
rect 11535 6089 11652 6098
rect 11672 6089 11683 6109
rect 11535 6081 11683 6089
rect 11750 6113 12109 6117
rect 11750 6108 12072 6113
rect 11750 6084 11863 6108
rect 11887 6089 12072 6108
rect 12096 6089 12109 6113
rect 11887 6084 12109 6089
rect 11750 6081 12109 6084
rect 12171 6081 12206 6118
rect 12274 6115 12374 6118
rect 12274 6111 12341 6115
rect 12274 6085 12286 6111
rect 12312 6089 12341 6111
rect 12367 6089 12374 6115
rect 12312 6085 12374 6089
rect 12274 6081 12374 6085
rect 11535 6065 11546 6081
rect 11535 6056 11543 6065
rect 11750 6060 11781 6081
rect 12171 6060 12207 6081
rect 11593 6059 11630 6060
rect 11258 6016 11323 6035
rect 11258 5998 11283 6016
rect 11301 5998 11323 6016
rect 9691 5933 9941 5935
rect 9691 5930 9792 5933
rect 9691 5911 9756 5930
rect 9753 5903 9756 5911
rect 9785 5903 9792 5930
rect 9820 5906 9830 5933
rect 9859 5911 9941 5933
rect 9964 5958 10281 5993
rect 9859 5906 9863 5911
rect 9820 5903 9863 5906
rect 9753 5889 9863 5903
rect 9179 5871 9520 5872
rect 9104 5869 9520 5871
rect 9964 5869 10004 5958
rect 10215 5931 10280 5958
rect 10215 5913 10238 5931
rect 10256 5913 10280 5931
rect 10215 5893 10280 5913
rect 9101 5866 10004 5869
rect 9101 5846 9107 5866
rect 9127 5846 10004 5866
rect 9101 5842 10004 5846
rect 9964 5839 10004 5842
rect 10216 5832 10281 5853
rect 8434 5824 9095 5825
rect 8434 5817 9368 5824
rect 8434 5816 9340 5817
rect 8434 5796 9285 5816
rect 9317 5797 9340 5816
rect 9365 5797 9368 5817
rect 9317 5796 9368 5797
rect 8434 5789 9368 5796
rect 8033 5747 8201 5748
rect 8436 5747 8475 5789
rect 9264 5787 9368 5789
rect 9333 5785 9368 5787
rect 10216 5814 10240 5832
rect 10258 5814 10281 5832
rect 10216 5767 10281 5814
rect 8033 5721 8477 5747
rect 8033 5719 8201 5721
rect 7835 5416 7904 5500
rect 7833 4937 7904 5416
rect 8033 5368 8060 5719
rect 8436 5715 8477 5721
rect 8100 5508 8164 5520
rect 8440 5516 8477 5715
rect 8939 5742 9011 5759
rect 8939 5703 8947 5742
rect 8992 5703 9011 5742
rect 8705 5605 8816 5620
rect 8705 5603 8747 5605
rect 8705 5583 8712 5603
rect 8731 5583 8747 5603
rect 8705 5575 8747 5583
rect 8775 5603 8816 5605
rect 8775 5583 8789 5603
rect 8808 5583 8816 5603
rect 8775 5575 8816 5583
rect 8705 5569 8816 5575
rect 8648 5547 8897 5569
rect 8648 5516 8685 5547
rect 8861 5545 8897 5547
rect 8861 5516 8898 5545
rect 8100 5507 8135 5508
rect 8077 5502 8135 5507
rect 8077 5482 8080 5502
rect 8100 5488 8135 5502
rect 8155 5488 8164 5508
rect 8100 5480 8164 5488
rect 8126 5479 8164 5480
rect 8127 5478 8164 5479
rect 8230 5512 8266 5513
rect 8338 5512 8374 5513
rect 8230 5504 8374 5512
rect 8230 5484 8238 5504
rect 8258 5484 8346 5504
rect 8366 5484 8374 5504
rect 8230 5478 8374 5484
rect 8440 5508 8478 5516
rect 8546 5512 8582 5513
rect 8440 5488 8449 5508
rect 8469 5488 8478 5508
rect 8440 5479 8478 5488
rect 8497 5505 8582 5512
rect 8497 5485 8504 5505
rect 8525 5504 8582 5505
rect 8525 5485 8554 5504
rect 8497 5484 8554 5485
rect 8574 5484 8582 5504
rect 8440 5478 8477 5479
rect 8497 5478 8582 5484
rect 8648 5508 8686 5516
rect 8759 5512 8795 5513
rect 8648 5488 8657 5508
rect 8677 5488 8686 5508
rect 8648 5479 8686 5488
rect 8710 5504 8795 5512
rect 8710 5484 8767 5504
rect 8787 5484 8795 5504
rect 8648 5478 8685 5479
rect 8710 5478 8795 5484
rect 8861 5508 8899 5516
rect 8861 5488 8870 5508
rect 8890 5488 8899 5508
rect 8861 5479 8899 5488
rect 8939 5493 9011 5703
rect 9081 5737 10281 5767
rect 9081 5736 9525 5737
rect 9081 5734 9249 5736
rect 8939 5479 9022 5493
rect 8861 5478 8898 5479
rect 8284 5457 8320 5478
rect 8710 5457 8741 5478
rect 8939 5457 8956 5479
rect 8117 5453 8217 5457
rect 8117 5449 8179 5453
rect 8117 5423 8124 5449
rect 8150 5427 8179 5449
rect 8205 5427 8217 5453
rect 8150 5423 8217 5427
rect 8117 5420 8217 5423
rect 8285 5420 8320 5457
rect 8382 5454 8741 5457
rect 8382 5449 8604 5454
rect 8382 5425 8395 5449
rect 8419 5430 8604 5449
rect 8628 5430 8741 5454
rect 8419 5425 8741 5430
rect 8382 5421 8741 5425
rect 8808 5449 8956 5457
rect 8808 5429 8819 5449
rect 8839 5446 8956 5449
rect 9009 5446 9022 5479
rect 8839 5429 9022 5446
rect 8808 5422 9022 5429
rect 8808 5421 8849 5422
rect 8939 5421 9022 5422
rect 8284 5395 8320 5420
rect 8132 5368 8169 5369
rect 8228 5368 8265 5369
rect 8284 5368 8291 5395
rect 8032 5359 8170 5368
rect 8032 5339 8141 5359
rect 8161 5339 8170 5359
rect 8032 5332 8170 5339
rect 8228 5365 8291 5368
rect 8312 5368 8320 5395
rect 8339 5368 8376 5369
rect 8312 5365 8376 5368
rect 8228 5359 8376 5365
rect 8228 5339 8237 5359
rect 8257 5339 8347 5359
rect 8367 5339 8376 5359
rect 8032 5330 8128 5332
rect 8228 5329 8376 5339
rect 8435 5359 8472 5369
rect 8547 5368 8584 5369
rect 8528 5366 8584 5368
rect 8435 5339 8443 5359
rect 8463 5339 8472 5359
rect 8284 5328 8320 5329
rect 8132 5197 8169 5198
rect 8435 5197 8472 5339
rect 8497 5359 8584 5366
rect 8497 5356 8555 5359
rect 8497 5336 8502 5356
rect 8523 5339 8555 5356
rect 8575 5339 8584 5359
rect 8523 5336 8584 5339
rect 8497 5329 8584 5336
rect 8643 5359 8680 5369
rect 8643 5339 8651 5359
rect 8671 5339 8680 5359
rect 8497 5328 8528 5329
rect 8643 5260 8680 5339
rect 8710 5368 8741 5421
rect 8947 5388 8961 5421
rect 9014 5388 9022 5421
rect 8947 5382 9022 5388
rect 8947 5377 9017 5382
rect 8760 5368 8797 5369
rect 8710 5359 8797 5368
rect 8710 5339 8768 5359
rect 8788 5339 8797 5359
rect 8710 5329 8797 5339
rect 8856 5359 8893 5369
rect 9081 5364 9108 5734
rect 9148 5504 9212 5516
rect 9488 5512 9525 5736
rect 9996 5717 10060 5719
rect 9992 5705 10060 5717
rect 9992 5672 10003 5705
rect 10043 5672 10060 5705
rect 9992 5662 10060 5672
rect 9753 5601 9864 5616
rect 9753 5599 9795 5601
rect 9753 5579 9760 5599
rect 9779 5579 9795 5599
rect 9753 5571 9795 5579
rect 9823 5599 9864 5601
rect 9823 5579 9837 5599
rect 9856 5579 9864 5599
rect 9823 5571 9864 5579
rect 9753 5565 9864 5571
rect 9696 5543 9945 5565
rect 9696 5512 9733 5543
rect 9909 5541 9945 5543
rect 9909 5512 9946 5541
rect 9148 5503 9183 5504
rect 9125 5498 9183 5503
rect 9125 5478 9128 5498
rect 9148 5484 9183 5498
rect 9203 5484 9212 5504
rect 9148 5476 9212 5484
rect 9174 5475 9212 5476
rect 9175 5474 9212 5475
rect 9278 5508 9314 5509
rect 9386 5508 9422 5509
rect 9278 5500 9422 5508
rect 9278 5480 9286 5500
rect 9306 5480 9394 5500
rect 9414 5480 9422 5500
rect 9278 5474 9422 5480
rect 9488 5504 9526 5512
rect 9594 5508 9630 5509
rect 9488 5484 9497 5504
rect 9517 5484 9526 5504
rect 9488 5475 9526 5484
rect 9545 5501 9630 5508
rect 9545 5481 9552 5501
rect 9573 5500 9630 5501
rect 9573 5481 9602 5500
rect 9545 5480 9602 5481
rect 9622 5480 9630 5500
rect 9488 5474 9525 5475
rect 9545 5474 9630 5480
rect 9696 5504 9734 5512
rect 9807 5508 9843 5509
rect 9696 5484 9705 5504
rect 9725 5484 9734 5504
rect 9696 5475 9734 5484
rect 9758 5500 9843 5508
rect 9758 5480 9815 5500
rect 9835 5480 9843 5500
rect 9696 5474 9733 5475
rect 9758 5474 9843 5480
rect 9909 5504 9947 5512
rect 9909 5484 9918 5504
rect 9938 5484 9947 5504
rect 9909 5475 9947 5484
rect 9996 5478 10060 5662
rect 10216 5536 10281 5737
rect 11258 5797 11323 5998
rect 11479 5872 11543 6056
rect 11592 6050 11630 6059
rect 11592 6030 11601 6050
rect 11621 6030 11630 6050
rect 11592 6022 11630 6030
rect 11696 6054 11781 6060
rect 11806 6059 11843 6060
rect 11696 6034 11704 6054
rect 11724 6034 11781 6054
rect 11696 6026 11781 6034
rect 11805 6050 11843 6059
rect 11805 6030 11814 6050
rect 11834 6030 11843 6050
rect 11696 6025 11732 6026
rect 11805 6022 11843 6030
rect 11909 6054 11994 6060
rect 12014 6059 12051 6060
rect 11909 6034 11917 6054
rect 11937 6053 11994 6054
rect 11937 6034 11966 6053
rect 11909 6033 11966 6034
rect 11987 6033 11994 6053
rect 11909 6026 11994 6033
rect 12013 6050 12051 6059
rect 12013 6030 12022 6050
rect 12042 6030 12051 6050
rect 11909 6025 11945 6026
rect 12013 6022 12051 6030
rect 12117 6054 12261 6060
rect 12117 6034 12125 6054
rect 12145 6034 12233 6054
rect 12253 6034 12261 6054
rect 12117 6026 12261 6034
rect 12117 6025 12153 6026
rect 12225 6025 12261 6026
rect 12327 6059 12364 6060
rect 12327 6058 12365 6059
rect 12327 6050 12391 6058
rect 12327 6030 12336 6050
rect 12356 6036 12391 6050
rect 12411 6036 12414 6056
rect 12356 6031 12414 6036
rect 12356 6030 12391 6031
rect 11593 5993 11630 6022
rect 11594 5991 11630 5993
rect 11806 5991 11843 6022
rect 11594 5969 11843 5991
rect 11675 5963 11786 5969
rect 11675 5955 11716 5963
rect 11675 5935 11683 5955
rect 11702 5935 11716 5955
rect 11675 5933 11716 5935
rect 11744 5955 11786 5963
rect 11744 5935 11760 5955
rect 11779 5935 11786 5955
rect 11744 5933 11786 5935
rect 11675 5918 11786 5933
rect 11479 5862 11547 5872
rect 11479 5829 11496 5862
rect 11536 5829 11547 5862
rect 11479 5817 11547 5829
rect 11479 5815 11543 5817
rect 12014 5798 12051 6022
rect 12327 6018 12391 6030
rect 12431 5800 12458 6170
rect 12646 6165 12683 6175
rect 12742 6195 12829 6205
rect 12742 6175 12751 6195
rect 12771 6175 12829 6195
rect 12742 6166 12829 6175
rect 12742 6165 12779 6166
rect 12522 6152 12592 6157
rect 12517 6146 12592 6152
rect 12517 6113 12525 6146
rect 12578 6113 12592 6146
rect 12798 6113 12829 6166
rect 12859 6195 12896 6274
rect 13011 6205 13042 6206
rect 12859 6175 12868 6195
rect 12888 6175 12896 6195
rect 12859 6165 12896 6175
rect 12955 6198 13042 6205
rect 12955 6195 13016 6198
rect 12955 6175 12964 6195
rect 12984 6178 13016 6195
rect 13037 6178 13042 6198
rect 12984 6175 13042 6178
rect 12955 6168 13042 6175
rect 13067 6195 13104 6337
rect 13370 6336 13407 6337
rect 13219 6205 13255 6206
rect 13067 6175 13076 6195
rect 13096 6175 13104 6195
rect 12955 6166 13011 6168
rect 12955 6165 12992 6166
rect 13067 6165 13104 6175
rect 13163 6195 13311 6205
rect 13411 6202 13507 6204
rect 13163 6175 13172 6195
rect 13192 6175 13282 6195
rect 13302 6175 13311 6195
rect 13163 6169 13311 6175
rect 13163 6166 13227 6169
rect 13163 6165 13200 6166
rect 13219 6139 13227 6166
rect 13248 6166 13311 6169
rect 13369 6195 13507 6202
rect 13369 6175 13378 6195
rect 13398 6175 13507 6195
rect 13369 6166 13507 6175
rect 13248 6139 13255 6166
rect 13274 6165 13311 6166
rect 13370 6165 13407 6166
rect 13219 6114 13255 6139
rect 12517 6112 12600 6113
rect 12690 6112 12731 6113
rect 12517 6105 12731 6112
rect 12517 6088 12700 6105
rect 12517 6055 12530 6088
rect 12583 6085 12700 6088
rect 12720 6085 12731 6105
rect 12583 6077 12731 6085
rect 12798 6109 13157 6113
rect 12798 6104 13120 6109
rect 12798 6080 12911 6104
rect 12935 6085 13120 6104
rect 13144 6085 13157 6109
rect 12935 6080 13157 6085
rect 12798 6077 13157 6080
rect 13219 6077 13254 6114
rect 13322 6111 13422 6114
rect 13322 6107 13389 6111
rect 13322 6081 13334 6107
rect 13360 6085 13389 6107
rect 13415 6085 13422 6111
rect 13360 6081 13422 6085
rect 13322 6077 13422 6081
rect 12583 6055 12600 6077
rect 12798 6056 12829 6077
rect 13219 6056 13255 6077
rect 12641 6055 12678 6056
rect 12517 6041 12600 6055
rect 12290 5798 12458 5800
rect 12014 5797 12458 5798
rect 11258 5767 12458 5797
rect 12528 5831 12600 6041
rect 12640 6046 12678 6055
rect 12640 6026 12649 6046
rect 12669 6026 12678 6046
rect 12640 6018 12678 6026
rect 12744 6050 12829 6056
rect 12854 6055 12891 6056
rect 12744 6030 12752 6050
rect 12772 6030 12829 6050
rect 12744 6022 12829 6030
rect 12853 6046 12891 6055
rect 12853 6026 12862 6046
rect 12882 6026 12891 6046
rect 12744 6021 12780 6022
rect 12853 6018 12891 6026
rect 12957 6050 13042 6056
rect 13062 6055 13099 6056
rect 12957 6030 12965 6050
rect 12985 6049 13042 6050
rect 12985 6030 13014 6049
rect 12957 6029 13014 6030
rect 13035 6029 13042 6049
rect 12957 6022 13042 6029
rect 13061 6046 13099 6055
rect 13061 6026 13070 6046
rect 13090 6026 13099 6046
rect 12957 6021 12993 6022
rect 13061 6018 13099 6026
rect 13165 6050 13309 6056
rect 13165 6030 13173 6050
rect 13193 6030 13281 6050
rect 13301 6030 13309 6050
rect 13165 6022 13309 6030
rect 13165 6021 13201 6022
rect 13273 6021 13309 6022
rect 13375 6055 13412 6056
rect 13375 6054 13413 6055
rect 13375 6046 13439 6054
rect 13375 6026 13384 6046
rect 13404 6032 13439 6046
rect 13459 6032 13462 6052
rect 13404 6027 13462 6032
rect 13404 6026 13439 6027
rect 12641 5989 12678 6018
rect 12642 5987 12678 5989
rect 12854 5987 12891 6018
rect 12642 5965 12891 5987
rect 12723 5959 12834 5965
rect 12723 5951 12764 5959
rect 12723 5931 12731 5951
rect 12750 5931 12764 5951
rect 12723 5929 12764 5931
rect 12792 5951 12834 5959
rect 12792 5931 12808 5951
rect 12827 5931 12834 5951
rect 12792 5929 12834 5931
rect 12723 5914 12834 5929
rect 12528 5792 12547 5831
rect 12592 5792 12600 5831
rect 12528 5775 12600 5792
rect 13062 5819 13099 6018
rect 13375 6014 13439 6026
rect 13062 5813 13103 5819
rect 13479 5815 13506 6166
rect 13629 6036 13708 6636
rect 13805 6184 13884 6769
rect 14088 6756 14125 6785
rect 14089 6754 14125 6756
rect 14301 6754 14338 6785
rect 14089 6732 14338 6754
rect 14170 6726 14281 6732
rect 14170 6718 14211 6726
rect 14170 6698 14178 6718
rect 14197 6698 14211 6718
rect 14170 6696 14211 6698
rect 14239 6718 14281 6726
rect 14239 6698 14255 6718
rect 14274 6698 14281 6718
rect 14239 6696 14281 6698
rect 14170 6681 14281 6696
rect 14509 6670 14546 6785
rect 14502 6558 14549 6670
rect 14670 6630 14700 6789
rect 14720 6788 14756 6789
rect 14822 6822 14859 6823
rect 14822 6821 14860 6822
rect 14822 6813 14886 6821
rect 14822 6793 14831 6813
rect 14851 6799 14886 6813
rect 14906 6799 14909 6819
rect 14851 6794 14909 6799
rect 14851 6793 14886 6794
rect 14822 6781 14886 6793
rect 14670 6626 14756 6630
rect 14670 6608 14685 6626
rect 14737 6608 14756 6626
rect 14670 6599 14756 6608
rect 14926 6560 14953 6933
rect 14785 6558 14953 6560
rect 14502 6532 14953 6558
rect 14502 6454 14549 6532
rect 14785 6531 14953 6532
rect 14447 6453 14549 6454
rect 14446 6445 14549 6453
rect 14446 6442 14498 6445
rect 14446 6407 14454 6442
rect 14479 6407 14498 6442
rect 14523 6407 14549 6445
rect 14446 6401 14549 6407
rect 14709 6446 14745 6450
rect 14709 6423 14717 6446
rect 14741 6423 14745 6446
rect 14709 6402 14745 6423
rect 14446 6397 14545 6401
rect 14709 6379 14717 6402
rect 14741 6379 14745 6402
rect 13338 5813 13506 5815
rect 13062 5787 13506 5813
rect 11258 5720 11323 5767
rect 11258 5702 11281 5720
rect 11299 5702 11323 5720
rect 12171 5747 12206 5749
rect 12171 5745 12275 5747
rect 13064 5745 13103 5787
rect 13338 5786 13506 5787
rect 12171 5738 13105 5745
rect 12171 5737 12222 5738
rect 12171 5717 12174 5737
rect 12199 5718 12222 5737
rect 12254 5718 13105 5738
rect 12199 5717 13105 5718
rect 12171 5710 13105 5717
rect 12444 5709 13105 5710
rect 11258 5681 11323 5702
rect 11535 5692 11575 5695
rect 11535 5688 12438 5692
rect 11535 5668 12412 5688
rect 12432 5668 12438 5688
rect 11535 5665 12438 5668
rect 11259 5621 11324 5641
rect 11259 5603 11283 5621
rect 11301 5603 11324 5621
rect 11259 5576 11324 5603
rect 11535 5576 11575 5665
rect 12019 5663 12435 5665
rect 12019 5662 12360 5663
rect 11676 5631 11786 5645
rect 11676 5628 11719 5631
rect 11676 5623 11680 5628
rect 11258 5541 11575 5576
rect 11598 5601 11680 5623
rect 11709 5601 11719 5628
rect 11747 5604 11754 5631
rect 11783 5623 11786 5631
rect 11783 5604 11848 5623
rect 11747 5601 11848 5604
rect 11598 5599 11848 5601
rect 10216 5518 10238 5536
rect 10256 5518 10281 5536
rect 10216 5499 10281 5518
rect 9909 5474 9946 5475
rect 9332 5453 9368 5474
rect 9758 5453 9789 5474
rect 9996 5469 10004 5478
rect 9993 5453 10004 5469
rect 9165 5449 9265 5453
rect 9165 5445 9227 5449
rect 9165 5419 9172 5445
rect 9198 5423 9227 5445
rect 9253 5423 9265 5449
rect 9198 5419 9265 5423
rect 9165 5416 9265 5419
rect 9333 5416 9368 5453
rect 9430 5450 9789 5453
rect 9430 5445 9652 5450
rect 9430 5421 9443 5445
rect 9467 5426 9652 5445
rect 9676 5426 9789 5450
rect 9467 5421 9789 5426
rect 9430 5417 9789 5421
rect 9856 5445 10004 5453
rect 9856 5425 9867 5445
rect 9887 5436 10004 5445
rect 10053 5469 10060 5478
rect 10053 5436 10061 5469
rect 11259 5465 11324 5541
rect 11598 5520 11635 5599
rect 11676 5586 11786 5599
rect 11750 5530 11781 5531
rect 11598 5500 11607 5520
rect 11627 5500 11635 5520
rect 11598 5490 11635 5500
rect 11694 5520 11781 5530
rect 11694 5500 11703 5520
rect 11723 5500 11781 5520
rect 11694 5491 11781 5500
rect 11694 5490 11731 5491
rect 9887 5425 10061 5436
rect 9856 5418 10061 5425
rect 9856 5417 9897 5418
rect 9332 5391 9368 5416
rect 9180 5364 9217 5365
rect 9276 5364 9313 5365
rect 9332 5364 9339 5391
rect 8856 5339 8864 5359
rect 8884 5339 8893 5359
rect 8710 5328 8741 5329
rect 8705 5260 8815 5273
rect 8856 5260 8893 5339
rect 9080 5355 9218 5364
rect 9080 5335 9189 5355
rect 9209 5335 9218 5355
rect 9080 5328 9218 5335
rect 9276 5361 9339 5364
rect 9360 5364 9368 5391
rect 9387 5364 9424 5365
rect 9360 5361 9424 5364
rect 9276 5355 9424 5361
rect 9276 5335 9285 5355
rect 9305 5335 9395 5355
rect 9415 5335 9424 5355
rect 9080 5326 9176 5328
rect 9276 5325 9424 5335
rect 9483 5355 9520 5365
rect 9595 5364 9632 5365
rect 9576 5362 9632 5364
rect 9483 5335 9491 5355
rect 9511 5335 9520 5355
rect 9332 5324 9368 5325
rect 8643 5258 8893 5260
rect 8643 5255 8744 5258
rect 8643 5236 8708 5255
rect 8705 5228 8708 5236
rect 8737 5228 8744 5255
rect 8772 5231 8782 5258
rect 8811 5236 8893 5258
rect 8811 5231 8815 5236
rect 8772 5228 8815 5231
rect 8705 5214 8815 5228
rect 8131 5196 8472 5197
rect 8056 5191 8472 5196
rect 9180 5193 9217 5194
rect 9483 5193 9520 5335
rect 9545 5355 9632 5362
rect 9545 5352 9603 5355
rect 9545 5332 9550 5352
rect 9571 5335 9603 5352
rect 9623 5335 9632 5355
rect 9571 5332 9632 5335
rect 9545 5325 9632 5332
rect 9691 5355 9728 5365
rect 9691 5335 9699 5355
rect 9719 5335 9728 5355
rect 9545 5324 9576 5325
rect 9691 5256 9728 5335
rect 9758 5364 9789 5417
rect 9993 5415 10061 5418
rect 9993 5373 10005 5415
rect 10054 5373 10061 5415
rect 9808 5364 9845 5365
rect 9758 5355 9845 5364
rect 9758 5335 9816 5355
rect 9836 5335 9845 5355
rect 9758 5325 9845 5335
rect 9904 5355 9941 5365
rect 9993 5360 10061 5373
rect 10216 5437 10281 5454
rect 10216 5419 10240 5437
rect 10258 5419 10281 5437
rect 11259 5447 11281 5465
rect 11299 5447 11324 5465
rect 11259 5426 11324 5447
rect 11472 5445 11537 5454
rect 9904 5335 9912 5355
rect 9932 5335 9941 5355
rect 9758 5324 9789 5325
rect 9753 5256 9863 5269
rect 9904 5256 9941 5335
rect 10216 5280 10281 5419
rect 11472 5408 11482 5445
rect 11522 5437 11537 5445
rect 11750 5438 11781 5491
rect 11811 5520 11848 5599
rect 11963 5530 11994 5531
rect 11811 5500 11820 5520
rect 11840 5500 11848 5520
rect 11811 5490 11848 5500
rect 11907 5523 11994 5530
rect 11907 5520 11968 5523
rect 11907 5500 11916 5520
rect 11936 5503 11968 5520
rect 11989 5503 11994 5523
rect 11936 5500 11994 5503
rect 11907 5493 11994 5500
rect 12019 5520 12056 5662
rect 12322 5661 12359 5662
rect 12171 5530 12207 5531
rect 12019 5500 12028 5520
rect 12048 5500 12056 5520
rect 11907 5491 11963 5493
rect 11907 5490 11944 5491
rect 12019 5490 12056 5500
rect 12115 5520 12263 5530
rect 12363 5527 12459 5529
rect 12115 5500 12124 5520
rect 12144 5500 12234 5520
rect 12254 5500 12263 5520
rect 12115 5494 12263 5500
rect 12115 5491 12179 5494
rect 12115 5490 12152 5491
rect 12171 5464 12179 5491
rect 12200 5491 12263 5494
rect 12321 5520 12459 5527
rect 12321 5500 12330 5520
rect 12350 5500 12459 5520
rect 12321 5491 12459 5500
rect 12200 5464 12207 5491
rect 12226 5490 12263 5491
rect 12322 5490 12359 5491
rect 12171 5439 12207 5464
rect 11642 5437 11683 5438
rect 11522 5430 11683 5437
rect 11522 5410 11652 5430
rect 11672 5410 11683 5430
rect 11522 5408 11683 5410
rect 11472 5402 11683 5408
rect 11750 5434 12109 5438
rect 11750 5429 12072 5434
rect 11750 5405 11863 5429
rect 11887 5410 12072 5429
rect 12096 5410 12109 5434
rect 11887 5405 12109 5410
rect 11750 5402 12109 5405
rect 12171 5402 12206 5439
rect 12274 5436 12374 5439
rect 12274 5432 12341 5436
rect 12274 5406 12286 5432
rect 12312 5410 12341 5432
rect 12367 5410 12374 5436
rect 12312 5406 12374 5410
rect 12274 5402 12374 5406
rect 11472 5389 11539 5402
rect 10216 5274 10238 5280
rect 9691 5254 9941 5256
rect 9691 5251 9792 5254
rect 9691 5232 9756 5251
rect 9753 5224 9756 5232
rect 9785 5224 9792 5251
rect 9820 5227 9830 5254
rect 9859 5232 9941 5254
rect 9970 5262 10238 5274
rect 10256 5262 10281 5280
rect 9970 5239 10281 5262
rect 11264 5366 11320 5386
rect 11264 5348 11283 5366
rect 11301 5348 11320 5366
rect 9970 5238 10025 5239
rect 9859 5227 9863 5232
rect 9820 5224 9863 5227
rect 9753 5210 9863 5224
rect 9179 5192 9520 5193
rect 8056 5171 8059 5191
rect 8079 5171 8472 5191
rect 9104 5191 9520 5192
rect 9970 5191 10013 5238
rect 11264 5235 11320 5348
rect 11472 5368 11486 5389
rect 11522 5368 11539 5389
rect 11750 5381 11781 5402
rect 12171 5381 12207 5402
rect 11593 5380 11630 5381
rect 11472 5361 11539 5368
rect 11592 5371 11630 5380
rect 9104 5187 10013 5191
rect 8423 5138 8468 5171
rect 9104 5167 9107 5187
rect 9127 5167 10013 5187
rect 9481 5162 10013 5167
rect 10221 5181 10280 5203
rect 10221 5163 10240 5181
rect 10258 5163 10280 5181
rect 9269 5138 9368 5140
rect 8423 5128 9368 5138
rect 8423 5102 9291 5128
rect 8424 5101 9291 5102
rect 9269 5090 9291 5101
rect 9316 5093 9335 5128
rect 9360 5093 9368 5128
rect 9316 5090 9368 5093
rect 9269 5082 9368 5090
rect 9295 5081 9367 5082
rect 10221 5033 10280 5163
rect 11264 5106 11319 5235
rect 11472 5209 11537 5361
rect 11592 5351 11601 5371
rect 11621 5351 11630 5371
rect 11592 5343 11630 5351
rect 11696 5375 11781 5381
rect 11806 5380 11843 5381
rect 11696 5355 11704 5375
rect 11724 5355 11781 5375
rect 11696 5347 11781 5355
rect 11805 5371 11843 5380
rect 11805 5351 11814 5371
rect 11834 5351 11843 5371
rect 11696 5346 11732 5347
rect 11805 5343 11843 5351
rect 11909 5375 11994 5381
rect 12014 5380 12051 5381
rect 11909 5355 11917 5375
rect 11937 5374 11994 5375
rect 11937 5355 11966 5374
rect 11909 5354 11966 5355
rect 11987 5354 11994 5374
rect 11909 5347 11994 5354
rect 12013 5371 12051 5380
rect 12013 5351 12022 5371
rect 12042 5351 12051 5371
rect 11909 5346 11945 5347
rect 12013 5343 12051 5351
rect 12117 5375 12261 5381
rect 12117 5355 12125 5375
rect 12145 5355 12233 5375
rect 12253 5355 12261 5375
rect 12117 5347 12261 5355
rect 12117 5346 12153 5347
rect 12225 5346 12261 5347
rect 12327 5380 12364 5381
rect 12327 5379 12365 5380
rect 12327 5371 12391 5379
rect 12327 5351 12336 5371
rect 12356 5357 12391 5371
rect 12411 5357 12414 5377
rect 12356 5352 12414 5357
rect 12356 5351 12391 5352
rect 11593 5314 11630 5343
rect 11594 5312 11630 5314
rect 11806 5312 11843 5343
rect 11594 5290 11843 5312
rect 11675 5284 11786 5290
rect 11675 5276 11716 5284
rect 11675 5256 11683 5276
rect 11702 5256 11716 5276
rect 11675 5254 11716 5256
rect 11744 5276 11786 5284
rect 11744 5256 11760 5276
rect 11779 5256 11786 5276
rect 11744 5254 11786 5256
rect 11675 5239 11786 5254
rect 12014 5244 12051 5343
rect 12327 5339 12391 5351
rect 11677 5230 11781 5239
rect 11465 5199 11586 5209
rect 11465 5197 11534 5199
rect 11465 5156 11478 5197
rect 11515 5158 11534 5197
rect 11571 5158 11586 5199
rect 11515 5156 11586 5158
rect 11465 5138 11586 5156
rect 11258 5094 11319 5106
rect 12012 5094 12053 5244
rect 12431 5236 12458 5491
rect 12520 5481 12600 5492
rect 12520 5455 12537 5481
rect 12577 5455 12600 5481
rect 12520 5428 12600 5455
rect 12520 5402 12541 5428
rect 12581 5402 12600 5428
rect 12520 5383 12600 5402
rect 12520 5357 12544 5383
rect 12584 5357 12600 5383
rect 12520 5306 12600 5357
rect 11258 5091 12053 5094
rect 12432 5105 12458 5236
rect 12522 5150 12592 5306
rect 12521 5134 12597 5150
rect 12432 5091 12460 5105
rect 11258 5056 12460 5091
rect 12521 5097 12536 5134
rect 12580 5097 12597 5134
rect 12521 5077 12597 5097
rect 13635 5127 13705 6036
rect 13804 5515 13885 6184
rect 14709 6079 14745 6379
rect 14633 6050 14746 6079
rect 14633 5685 14664 6050
rect 14557 5665 14950 5685
rect 14970 5665 14973 5685
rect 14557 5660 14973 5665
rect 14557 5659 14898 5660
rect 14214 5628 14324 5642
rect 14214 5625 14257 5628
rect 14214 5620 14218 5625
rect 14136 5598 14218 5620
rect 14247 5598 14257 5625
rect 14285 5601 14292 5628
rect 14321 5620 14324 5628
rect 14321 5601 14386 5620
rect 14285 5598 14386 5601
rect 14136 5596 14386 5598
rect 14136 5517 14173 5596
rect 14214 5583 14324 5596
rect 14288 5527 14319 5528
rect 13798 5435 13897 5515
rect 14136 5497 14145 5517
rect 14165 5497 14173 5517
rect 14136 5487 14173 5497
rect 14232 5517 14319 5527
rect 14232 5497 14241 5517
rect 14261 5497 14319 5517
rect 14232 5488 14319 5497
rect 14232 5487 14269 5488
rect 14288 5435 14319 5488
rect 14349 5517 14386 5596
rect 14501 5527 14532 5528
rect 14349 5497 14358 5517
rect 14378 5497 14386 5517
rect 14349 5487 14386 5497
rect 14445 5520 14532 5527
rect 14445 5517 14506 5520
rect 14445 5497 14454 5517
rect 14474 5500 14506 5517
rect 14527 5500 14532 5520
rect 14474 5497 14532 5500
rect 14445 5490 14532 5497
rect 14557 5517 14594 5659
rect 14860 5658 14897 5659
rect 14709 5527 14745 5528
rect 14557 5497 14566 5517
rect 14586 5497 14594 5517
rect 14445 5488 14501 5490
rect 14445 5487 14482 5488
rect 14557 5487 14594 5497
rect 14653 5517 14801 5527
rect 14901 5524 14997 5526
rect 14653 5497 14662 5517
rect 14682 5497 14772 5517
rect 14792 5497 14801 5517
rect 14653 5491 14801 5497
rect 14653 5488 14717 5491
rect 14653 5487 14690 5488
rect 14709 5461 14717 5488
rect 14738 5488 14801 5491
rect 14859 5517 14997 5524
rect 14859 5497 14868 5517
rect 14888 5497 14997 5517
rect 14859 5488 14997 5497
rect 14738 5461 14745 5488
rect 14764 5487 14801 5488
rect 14860 5487 14897 5488
rect 14709 5436 14745 5461
rect 13798 5434 14138 5435
rect 14180 5434 14221 5435
rect 13798 5427 14221 5434
rect 13798 5407 14190 5427
rect 14210 5407 14221 5427
rect 13798 5399 14221 5407
rect 14288 5431 14647 5435
rect 14288 5426 14610 5431
rect 14288 5402 14401 5426
rect 14425 5407 14610 5426
rect 14634 5407 14647 5431
rect 14425 5402 14647 5407
rect 14288 5399 14647 5402
rect 14709 5399 14744 5436
rect 14812 5433 14912 5436
rect 14812 5429 14879 5433
rect 14812 5403 14824 5429
rect 14850 5407 14879 5429
rect 14905 5407 14912 5433
rect 14850 5403 14912 5407
rect 14812 5399 14912 5403
rect 13798 5395 14138 5399
rect 13635 5077 13707 5127
rect 8943 5003 9019 5027
rect 8943 4937 8955 5003
rect 9009 4937 9019 5003
rect 9487 4958 9528 4960
rect 9759 4958 9863 4960
rect 10221 4958 10282 5033
rect 11258 4981 11319 5056
rect 11677 5054 11781 5056
rect 12012 5054 12053 5056
rect 12521 5011 12531 5077
rect 12585 5011 12597 5077
rect 12521 4987 12597 5011
rect 7833 4887 7905 4937
rect 7402 4615 7738 4619
rect 6628 4611 6728 4615
rect 6628 4607 6690 4611
rect 6628 4581 6635 4607
rect 6661 4585 6690 4607
rect 6716 4585 6728 4611
rect 6661 4581 6728 4585
rect 6628 4578 6728 4581
rect 6796 4578 6831 4615
rect 6893 4612 7252 4615
rect 6893 4607 7115 4612
rect 6893 4583 6906 4607
rect 6930 4588 7115 4607
rect 7139 4588 7252 4612
rect 6930 4583 7252 4588
rect 6893 4579 7252 4583
rect 7319 4607 7738 4615
rect 7319 4587 7330 4607
rect 7350 4587 7738 4607
rect 7319 4580 7738 4587
rect 7319 4579 7360 4580
rect 7402 4579 7738 4580
rect 6795 4553 6831 4578
rect 6643 4526 6680 4527
rect 6739 4526 6776 4527
rect 6795 4526 6802 4553
rect 6543 4517 6681 4526
rect 6543 4497 6652 4517
rect 6672 4497 6681 4517
rect 6543 4490 6681 4497
rect 6739 4523 6802 4526
rect 6823 4526 6831 4553
rect 6850 4526 6887 4527
rect 6823 4523 6887 4526
rect 6739 4517 6887 4523
rect 6739 4497 6748 4517
rect 6768 4497 6858 4517
rect 6878 4497 6887 4517
rect 6543 4488 6639 4490
rect 6739 4487 6887 4497
rect 6946 4517 6983 4527
rect 7058 4526 7095 4527
rect 7039 4524 7095 4526
rect 6946 4497 6954 4517
rect 6974 4497 6983 4517
rect 6795 4486 6831 4487
rect 6643 4355 6680 4356
rect 6946 4355 6983 4497
rect 7008 4517 7095 4524
rect 7008 4514 7066 4517
rect 7008 4494 7013 4514
rect 7034 4497 7066 4514
rect 7086 4497 7095 4517
rect 7034 4494 7095 4497
rect 7008 4487 7095 4494
rect 7154 4517 7191 4527
rect 7154 4497 7162 4517
rect 7182 4497 7191 4517
rect 7008 4486 7039 4487
rect 7154 4418 7191 4497
rect 7221 4526 7252 4579
rect 7646 4543 7738 4579
rect 7271 4526 7308 4527
rect 7221 4517 7308 4526
rect 7221 4497 7279 4517
rect 7299 4497 7308 4517
rect 7221 4487 7308 4497
rect 7367 4517 7404 4527
rect 7367 4497 7375 4517
rect 7395 4497 7404 4517
rect 7221 4486 7252 4487
rect 7216 4418 7326 4431
rect 7367 4418 7404 4497
rect 7154 4416 7404 4418
rect 7154 4413 7255 4416
rect 7154 4394 7219 4413
rect 7216 4386 7219 4394
rect 7248 4386 7255 4413
rect 7283 4389 7293 4416
rect 7322 4394 7404 4416
rect 7322 4389 7326 4394
rect 7283 4386 7326 4389
rect 7216 4372 7326 4386
rect 6642 4354 6983 4355
rect 6567 4349 6983 4354
rect 6567 4329 6570 4349
rect 6590 4329 6983 4349
rect 6727 4285 6832 4288
rect 6726 4262 6832 4285
rect 5846 4260 6347 4262
rect 6488 4260 6837 4262
rect 3960 4239 3997 4260
rect 3960 4202 3971 4239
rect 3988 4202 3997 4239
rect 5846 4254 6837 4260
rect 5846 4249 6798 4254
rect 5846 4228 6757 4249
rect 6777 4233 6798 4249
rect 6818 4233 6837 4254
rect 6777 4228 6837 4233
rect 5846 4203 6837 4228
rect 6322 4202 6504 4203
rect 3960 4192 3997 4202
rect 3806 4149 4200 4169
rect 4220 4149 4223 4169
rect 3807 4144 4223 4149
rect 3807 4143 4148 4144
rect 3464 4112 3574 4126
rect 3464 4109 3507 4112
rect 3464 4104 3468 4109
rect 3386 4082 3468 4104
rect 3497 4082 3507 4109
rect 3535 4085 3542 4112
rect 3571 4104 3574 4112
rect 3571 4085 3636 4104
rect 3535 4082 3636 4085
rect 3386 4080 3636 4082
rect 3386 4001 3423 4080
rect 3464 4067 3574 4080
rect 3538 4011 3569 4012
rect 3386 3981 3395 4001
rect 3415 3981 3423 4001
rect 3386 3971 3423 3981
rect 3482 4001 3569 4011
rect 3482 3981 3491 4001
rect 3511 3981 3569 4001
rect 3482 3972 3569 3981
rect 3482 3971 3519 3972
rect 3538 3919 3569 3972
rect 3599 4001 3636 4080
rect 3751 4011 3782 4012
rect 3599 3981 3608 4001
rect 3628 3981 3636 4001
rect 3599 3971 3636 3981
rect 3695 4004 3782 4011
rect 3695 4001 3756 4004
rect 3695 3981 3704 4001
rect 3724 3984 3756 4001
rect 3777 3984 3782 4004
rect 3724 3981 3782 3984
rect 3695 3974 3782 3981
rect 3807 4001 3844 4143
rect 4110 4142 4147 4143
rect 3959 4011 3995 4012
rect 3807 3981 3816 4001
rect 3836 3981 3844 4001
rect 3695 3972 3751 3974
rect 3695 3971 3732 3972
rect 3807 3971 3844 3981
rect 3903 4001 4051 4011
rect 4151 4008 4247 4010
rect 3903 3981 3912 4001
rect 3932 3981 4022 4001
rect 4042 3981 4051 4001
rect 3903 3975 4051 3981
rect 3903 3972 3967 3975
rect 3903 3971 3940 3972
rect 3959 3945 3967 3972
rect 3988 3972 4051 3975
rect 4109 4001 4247 4008
rect 4109 3981 4118 4001
rect 4138 3981 4247 4001
rect 4109 3972 4247 3981
rect 6876 3973 6907 4329
rect 3988 3945 3995 3972
rect 4014 3971 4051 3972
rect 4110 3971 4147 3972
rect 3959 3920 3995 3945
rect 3430 3918 3471 3919
rect 3350 3913 3471 3918
rect 3301 3911 3471 3913
rect 3301 3900 3440 3911
rect 3301 3877 3324 3900
rect 3350 3891 3440 3900
rect 3460 3891 3471 3911
rect 3350 3883 3471 3891
rect 3538 3915 3897 3919
rect 3538 3910 3860 3915
rect 3538 3886 3651 3910
rect 3675 3891 3860 3910
rect 3884 3891 3897 3915
rect 3675 3886 3897 3891
rect 3538 3883 3897 3886
rect 3959 3883 3994 3920
rect 4062 3917 4162 3920
rect 4062 3913 4129 3917
rect 4062 3887 4074 3913
rect 4100 3891 4129 3913
rect 4155 3891 4162 3917
rect 4100 3887 4162 3891
rect 4062 3883 4162 3887
rect 3350 3877 3358 3883
rect 3301 3869 3358 3877
rect 3538 3862 3569 3883
rect 3959 3862 3995 3883
rect 3381 3861 3418 3862
rect 3380 3852 3418 3861
rect 3380 3832 3389 3852
rect 3409 3832 3418 3852
rect 3380 3824 3418 3832
rect 3484 3856 3569 3862
rect 3594 3861 3631 3862
rect 3484 3836 3492 3856
rect 3512 3836 3569 3856
rect 3484 3828 3569 3836
rect 3593 3852 3631 3861
rect 3593 3832 3602 3852
rect 3622 3832 3631 3852
rect 3484 3827 3520 3828
rect 3593 3824 3631 3832
rect 3697 3856 3782 3862
rect 3802 3861 3839 3862
rect 3697 3836 3705 3856
rect 3725 3855 3782 3856
rect 3725 3836 3754 3855
rect 3697 3835 3754 3836
rect 3775 3835 3782 3855
rect 3697 3828 3782 3835
rect 3801 3852 3839 3861
rect 3801 3832 3810 3852
rect 3830 3832 3839 3852
rect 3697 3827 3733 3828
rect 3801 3824 3839 3832
rect 3905 3856 4049 3862
rect 3905 3836 3913 3856
rect 3933 3836 4021 3856
rect 4041 3836 4049 3856
rect 3905 3828 4049 3836
rect 3905 3827 3941 3828
rect 4013 3827 4049 3828
rect 4115 3861 4152 3862
rect 4115 3860 4153 3861
rect 4115 3852 4179 3860
rect 4115 3832 4124 3852
rect 4144 3838 4179 3852
rect 4199 3838 4202 3858
rect 4144 3833 4202 3838
rect 4144 3832 4179 3833
rect 3381 3795 3418 3824
rect 3382 3793 3418 3795
rect 3594 3793 3631 3824
rect 3382 3771 3631 3793
rect 3463 3765 3574 3771
rect 3463 3757 3504 3765
rect 3463 3737 3471 3757
rect 3490 3737 3504 3757
rect 3463 3735 3504 3737
rect 3532 3757 3574 3765
rect 3532 3737 3548 3757
rect 3567 3737 3574 3757
rect 3532 3735 3574 3737
rect 3463 3720 3574 3735
rect 3802 3709 3839 3824
rect 4115 3820 4179 3832
rect 3795 3703 3842 3709
rect 4219 3705 4246 3972
rect 6794 3944 6907 3973
rect 4078 3703 4246 3705
rect 3795 3677 4246 3703
rect 3795 3542 3842 3677
rect 4078 3676 4246 3677
rect 6795 3635 6831 3944
rect 7655 3830 7736 4543
rect 7835 3978 7905 4887
rect 8943 4917 9019 4937
rect 8943 4880 8960 4917
rect 9004 4880 9019 4917
rect 9080 4923 10282 4958
rect 9080 4909 9108 4923
rect 8943 4864 9019 4880
rect 8948 4708 9018 4864
rect 9082 4778 9108 4909
rect 9487 4920 10282 4923
rect 8940 4657 9020 4708
rect 8940 4631 8956 4657
rect 8996 4631 9020 4657
rect 8940 4612 9020 4631
rect 8940 4586 8959 4612
rect 8999 4586 9020 4612
rect 8940 4559 9020 4586
rect 8940 4533 8963 4559
rect 9003 4533 9020 4559
rect 8940 4522 9020 4533
rect 9082 4523 9109 4778
rect 9487 4770 9528 4920
rect 10221 4908 10282 4920
rect 9954 4858 10075 4876
rect 9954 4856 10025 4858
rect 9954 4815 9969 4856
rect 10006 4817 10025 4856
rect 10062 4817 10075 4858
rect 10006 4815 10075 4817
rect 9954 4805 10075 4815
rect 9759 4775 9863 4784
rect 9149 4663 9213 4675
rect 9489 4671 9526 4770
rect 9754 4760 9865 4775
rect 9754 4758 9796 4760
rect 9754 4738 9761 4758
rect 9780 4738 9796 4758
rect 9754 4730 9796 4738
rect 9824 4758 9865 4760
rect 9824 4738 9838 4758
rect 9857 4738 9865 4758
rect 9824 4730 9865 4738
rect 9754 4724 9865 4730
rect 9697 4702 9946 4724
rect 9697 4671 9734 4702
rect 9910 4700 9946 4702
rect 9910 4671 9947 4700
rect 9149 4662 9184 4663
rect 9126 4657 9184 4662
rect 9126 4637 9129 4657
rect 9149 4643 9184 4657
rect 9204 4643 9213 4663
rect 9149 4635 9213 4643
rect 9175 4634 9213 4635
rect 9176 4633 9213 4634
rect 9279 4667 9315 4668
rect 9387 4667 9423 4668
rect 9279 4659 9423 4667
rect 9279 4639 9287 4659
rect 9307 4639 9395 4659
rect 9415 4639 9423 4659
rect 9279 4633 9423 4639
rect 9489 4663 9527 4671
rect 9595 4667 9631 4668
rect 9489 4643 9498 4663
rect 9518 4643 9527 4663
rect 9489 4634 9527 4643
rect 9546 4660 9631 4667
rect 9546 4640 9553 4660
rect 9574 4659 9631 4660
rect 9574 4640 9603 4659
rect 9546 4639 9603 4640
rect 9623 4639 9631 4659
rect 9489 4633 9526 4634
rect 9546 4633 9631 4639
rect 9697 4663 9735 4671
rect 9808 4667 9844 4668
rect 9697 4643 9706 4663
rect 9726 4643 9735 4663
rect 9697 4634 9735 4643
rect 9759 4659 9844 4667
rect 9759 4639 9816 4659
rect 9836 4639 9844 4659
rect 9697 4633 9734 4634
rect 9759 4633 9844 4639
rect 9910 4663 9948 4671
rect 9910 4643 9919 4663
rect 9939 4643 9948 4663
rect 10003 4653 10068 4805
rect 10221 4779 10276 4908
rect 11260 4851 11319 4981
rect 12173 4932 12245 4933
rect 12172 4924 12271 4932
rect 12172 4921 12224 4924
rect 12172 4886 12180 4921
rect 12205 4886 12224 4921
rect 12249 4913 12271 4924
rect 12249 4912 13116 4913
rect 12249 4886 13117 4912
rect 12172 4876 13117 4886
rect 12172 4874 12271 4876
rect 11260 4833 11282 4851
rect 11300 4833 11319 4851
rect 11260 4811 11319 4833
rect 11527 4847 12059 4852
rect 11527 4827 12413 4847
rect 12433 4827 12436 4847
rect 13072 4843 13117 4876
rect 11527 4823 12436 4827
rect 9910 4634 9948 4643
rect 10001 4646 10068 4653
rect 9910 4633 9947 4634
rect 9333 4612 9369 4633
rect 9759 4612 9790 4633
rect 10001 4625 10018 4646
rect 10054 4625 10068 4646
rect 10220 4666 10276 4779
rect 11527 4776 11570 4823
rect 12020 4822 12436 4823
rect 13068 4823 13461 4843
rect 13481 4823 13484 4843
rect 12020 4821 12361 4822
rect 11677 4790 11787 4804
rect 11677 4787 11720 4790
rect 11677 4782 11681 4787
rect 11515 4775 11570 4776
rect 10220 4648 10239 4666
rect 10257 4648 10276 4666
rect 10220 4628 10276 4648
rect 11259 4752 11570 4775
rect 11259 4734 11284 4752
rect 11302 4740 11570 4752
rect 11599 4760 11681 4782
rect 11710 4760 11720 4787
rect 11748 4763 11755 4790
rect 11784 4782 11787 4790
rect 11784 4763 11849 4782
rect 11748 4760 11849 4763
rect 11599 4758 11849 4760
rect 11302 4734 11324 4740
rect 10001 4612 10068 4625
rect 9166 4608 9266 4612
rect 9166 4604 9228 4608
rect 9166 4578 9173 4604
rect 9199 4582 9228 4604
rect 9254 4582 9266 4608
rect 9199 4578 9266 4582
rect 9166 4575 9266 4578
rect 9334 4575 9369 4612
rect 9431 4609 9790 4612
rect 9431 4604 9653 4609
rect 9431 4580 9444 4604
rect 9468 4585 9653 4604
rect 9677 4585 9790 4609
rect 9468 4580 9790 4585
rect 9431 4576 9790 4580
rect 9857 4606 10068 4612
rect 9857 4604 10018 4606
rect 9857 4584 9868 4604
rect 9888 4584 10018 4604
rect 9857 4577 10018 4584
rect 9857 4576 9898 4577
rect 9333 4550 9369 4575
rect 9181 4523 9218 4524
rect 9277 4523 9314 4524
rect 9333 4523 9340 4550
rect 9081 4514 9219 4523
rect 9081 4494 9190 4514
rect 9210 4494 9219 4514
rect 9081 4487 9219 4494
rect 9277 4520 9340 4523
rect 9361 4523 9369 4550
rect 9388 4523 9425 4524
rect 9361 4520 9425 4523
rect 9277 4514 9425 4520
rect 9277 4494 9286 4514
rect 9306 4494 9396 4514
rect 9416 4494 9425 4514
rect 9081 4485 9177 4487
rect 9277 4484 9425 4494
rect 9484 4514 9521 4524
rect 9596 4523 9633 4524
rect 9577 4521 9633 4523
rect 9484 4494 9492 4514
rect 9512 4494 9521 4514
rect 9333 4483 9369 4484
rect 9181 4352 9218 4353
rect 9484 4352 9521 4494
rect 9546 4514 9633 4521
rect 9546 4511 9604 4514
rect 9546 4491 9551 4511
rect 9572 4494 9604 4511
rect 9624 4494 9633 4514
rect 9572 4491 9633 4494
rect 9546 4484 9633 4491
rect 9692 4514 9729 4524
rect 9692 4494 9700 4514
rect 9720 4494 9729 4514
rect 9546 4483 9577 4484
rect 9692 4415 9729 4494
rect 9759 4523 9790 4576
rect 10003 4569 10018 4577
rect 10058 4569 10068 4606
rect 11259 4595 11324 4734
rect 11599 4679 11636 4758
rect 11677 4745 11787 4758
rect 11751 4689 11782 4690
rect 11599 4659 11608 4679
rect 11628 4659 11636 4679
rect 10003 4560 10068 4569
rect 10216 4567 10281 4588
rect 10216 4549 10241 4567
rect 10259 4549 10281 4567
rect 11259 4577 11282 4595
rect 11300 4577 11324 4595
rect 11259 4560 11324 4577
rect 11479 4641 11547 4654
rect 11599 4649 11636 4659
rect 11695 4679 11782 4689
rect 11695 4659 11704 4679
rect 11724 4659 11782 4679
rect 11695 4650 11782 4659
rect 11695 4649 11732 4650
rect 11479 4599 11486 4641
rect 11535 4599 11547 4641
rect 11479 4596 11547 4599
rect 11751 4597 11782 4650
rect 11812 4679 11849 4758
rect 11964 4689 11995 4690
rect 11812 4659 11821 4679
rect 11841 4659 11849 4679
rect 11812 4649 11849 4659
rect 11908 4682 11995 4689
rect 11908 4679 11969 4682
rect 11908 4659 11917 4679
rect 11937 4662 11969 4679
rect 11990 4662 11995 4682
rect 11937 4659 11995 4662
rect 11908 4652 11995 4659
rect 12020 4679 12057 4821
rect 12323 4820 12360 4821
rect 13068 4818 13484 4823
rect 13068 4817 13409 4818
rect 12725 4786 12835 4800
rect 12725 4783 12768 4786
rect 12725 4778 12729 4783
rect 12647 4756 12729 4778
rect 12758 4756 12768 4783
rect 12796 4759 12803 4786
rect 12832 4778 12835 4786
rect 12832 4759 12897 4778
rect 12796 4756 12897 4759
rect 12647 4754 12897 4756
rect 12172 4689 12208 4690
rect 12020 4659 12029 4679
rect 12049 4659 12057 4679
rect 11908 4650 11964 4652
rect 11908 4649 11945 4650
rect 12020 4649 12057 4659
rect 12116 4679 12264 4689
rect 12364 4686 12460 4688
rect 12116 4659 12125 4679
rect 12145 4659 12235 4679
rect 12255 4659 12264 4679
rect 12116 4653 12264 4659
rect 12116 4650 12180 4653
rect 12116 4649 12153 4650
rect 12172 4623 12180 4650
rect 12201 4650 12264 4653
rect 12322 4679 12460 4686
rect 12322 4659 12331 4679
rect 12351 4659 12460 4679
rect 12322 4650 12460 4659
rect 12647 4675 12684 4754
rect 12725 4741 12835 4754
rect 12799 4685 12830 4686
rect 12647 4655 12656 4675
rect 12676 4655 12684 4675
rect 12201 4623 12208 4650
rect 12227 4649 12264 4650
rect 12323 4649 12360 4650
rect 12172 4598 12208 4623
rect 11643 4596 11684 4597
rect 11479 4589 11684 4596
rect 11479 4578 11653 4589
rect 9809 4523 9846 4524
rect 9759 4514 9846 4523
rect 9759 4494 9817 4514
rect 9837 4494 9846 4514
rect 9759 4484 9846 4494
rect 9905 4514 9942 4524
rect 9905 4494 9913 4514
rect 9933 4494 9942 4514
rect 9759 4483 9790 4484
rect 9754 4415 9864 4428
rect 9905 4415 9942 4494
rect 10216 4473 10281 4549
rect 11479 4545 11487 4578
rect 11480 4536 11487 4545
rect 11536 4569 11653 4578
rect 11673 4569 11684 4589
rect 11536 4561 11684 4569
rect 11751 4593 12110 4597
rect 11751 4588 12073 4593
rect 11751 4564 11864 4588
rect 11888 4569 12073 4588
rect 12097 4569 12110 4593
rect 11888 4564 12110 4569
rect 11751 4561 12110 4564
rect 12172 4561 12207 4598
rect 12275 4595 12375 4598
rect 12275 4591 12342 4595
rect 12275 4565 12287 4591
rect 12313 4569 12342 4591
rect 12368 4569 12375 4595
rect 12313 4565 12375 4569
rect 12275 4561 12375 4565
rect 11536 4545 11547 4561
rect 11536 4536 11544 4545
rect 11751 4540 11782 4561
rect 12172 4540 12208 4561
rect 11594 4539 11631 4540
rect 11259 4496 11324 4515
rect 11259 4478 11284 4496
rect 11302 4478 11324 4496
rect 9692 4413 9942 4415
rect 9692 4410 9793 4413
rect 9692 4391 9757 4410
rect 9754 4383 9757 4391
rect 9786 4383 9793 4410
rect 9821 4386 9831 4413
rect 9860 4391 9942 4413
rect 9965 4438 10282 4473
rect 9860 4386 9864 4391
rect 9821 4383 9864 4386
rect 9754 4369 9864 4383
rect 9180 4351 9521 4352
rect 9105 4349 9521 4351
rect 9965 4349 10005 4438
rect 10216 4411 10281 4438
rect 10216 4393 10239 4411
rect 10257 4393 10281 4411
rect 10216 4373 10281 4393
rect 9102 4346 10005 4349
rect 9102 4326 9108 4346
rect 9128 4326 10005 4346
rect 9102 4322 10005 4326
rect 9965 4319 10005 4322
rect 10217 4312 10282 4333
rect 8435 4304 9096 4305
rect 8435 4297 9369 4304
rect 8435 4296 9341 4297
rect 8435 4276 9286 4296
rect 9318 4277 9341 4296
rect 9366 4277 9369 4297
rect 9318 4276 9369 4277
rect 8435 4269 9369 4276
rect 8034 4227 8202 4228
rect 8437 4227 8476 4269
rect 9265 4267 9369 4269
rect 9334 4265 9369 4267
rect 10217 4294 10241 4312
rect 10259 4294 10282 4312
rect 10217 4247 10282 4294
rect 8034 4201 8478 4227
rect 8034 4199 8202 4201
rect 6795 3612 6799 3635
rect 6823 3612 6831 3635
rect 6995 3613 7094 3617
rect 6795 3591 6831 3612
rect 6795 3568 6799 3591
rect 6823 3568 6831 3591
rect 6795 3564 6831 3568
rect 6991 3607 7094 3613
rect 6991 3569 7017 3607
rect 7042 3572 7061 3607
rect 7086 3572 7094 3607
rect 7042 3569 7094 3572
rect 6991 3561 7094 3569
rect 6991 3560 7093 3561
rect 3793 3493 3852 3542
rect 3793 3465 3811 3493
rect 3839 3465 3852 3493
rect 3793 3455 3852 3465
rect 6587 3482 6755 3483
rect 6991 3482 7038 3560
rect 6587 3456 7038 3482
rect 6587 3454 6755 3456
rect 6587 3081 6614 3454
rect 6784 3406 6870 3415
rect 6784 3388 6803 3406
rect 6855 3388 6870 3406
rect 6784 3384 6870 3388
rect 6654 3221 6718 3233
rect 6654 3220 6689 3221
rect 6631 3215 6689 3220
rect 6631 3195 6634 3215
rect 6654 3201 6689 3215
rect 6709 3201 6718 3221
rect 6654 3193 6718 3201
rect 6680 3192 6718 3193
rect 6681 3191 6718 3192
rect 6784 3225 6820 3226
rect 6840 3225 6870 3384
rect 6991 3344 7038 3456
rect 6994 3229 7031 3344
rect 7259 3318 7370 3333
rect 7259 3316 7301 3318
rect 7259 3296 7266 3316
rect 7285 3296 7301 3316
rect 7259 3288 7301 3296
rect 7329 3316 7370 3318
rect 7329 3296 7343 3316
rect 7362 3296 7370 3316
rect 7329 3288 7370 3296
rect 7259 3282 7370 3288
rect 7202 3260 7451 3282
rect 7202 3229 7239 3260
rect 7415 3258 7451 3260
rect 7415 3229 7452 3258
rect 7656 3245 7735 3830
rect 7832 3378 7911 3978
rect 8034 3848 8061 4199
rect 8437 4195 8478 4201
rect 8101 3988 8165 4000
rect 8441 3996 8478 4195
rect 8940 4222 9012 4239
rect 8940 4183 8948 4222
rect 8993 4183 9012 4222
rect 8706 4085 8817 4100
rect 8706 4083 8748 4085
rect 8706 4063 8713 4083
rect 8732 4063 8748 4083
rect 8706 4055 8748 4063
rect 8776 4083 8817 4085
rect 8776 4063 8790 4083
rect 8809 4063 8817 4083
rect 8776 4055 8817 4063
rect 8706 4049 8817 4055
rect 8649 4027 8898 4049
rect 8649 3996 8686 4027
rect 8862 4025 8898 4027
rect 8862 3996 8899 4025
rect 8101 3987 8136 3988
rect 8078 3982 8136 3987
rect 8078 3962 8081 3982
rect 8101 3968 8136 3982
rect 8156 3968 8165 3988
rect 8101 3960 8165 3968
rect 8127 3959 8165 3960
rect 8128 3958 8165 3959
rect 8231 3992 8267 3993
rect 8339 3992 8375 3993
rect 8231 3984 8375 3992
rect 8231 3964 8239 3984
rect 8259 3964 8347 3984
rect 8367 3964 8375 3984
rect 8231 3958 8375 3964
rect 8441 3988 8479 3996
rect 8547 3992 8583 3993
rect 8441 3968 8450 3988
rect 8470 3968 8479 3988
rect 8441 3959 8479 3968
rect 8498 3985 8583 3992
rect 8498 3965 8505 3985
rect 8526 3984 8583 3985
rect 8526 3965 8555 3984
rect 8498 3964 8555 3965
rect 8575 3964 8583 3984
rect 8441 3958 8478 3959
rect 8498 3958 8583 3964
rect 8649 3988 8687 3996
rect 8760 3992 8796 3993
rect 8649 3968 8658 3988
rect 8678 3968 8687 3988
rect 8649 3959 8687 3968
rect 8711 3984 8796 3992
rect 8711 3964 8768 3984
rect 8788 3964 8796 3984
rect 8649 3958 8686 3959
rect 8711 3958 8796 3964
rect 8862 3988 8900 3996
rect 8862 3968 8871 3988
rect 8891 3968 8900 3988
rect 8862 3959 8900 3968
rect 8940 3973 9012 4183
rect 9082 4217 10282 4247
rect 9082 4216 9526 4217
rect 9082 4214 9250 4216
rect 8940 3959 9023 3973
rect 8862 3958 8899 3959
rect 8285 3937 8321 3958
rect 8711 3937 8742 3958
rect 8940 3937 8957 3959
rect 8118 3933 8218 3937
rect 8118 3929 8180 3933
rect 8118 3903 8125 3929
rect 8151 3907 8180 3929
rect 8206 3907 8218 3933
rect 8151 3903 8218 3907
rect 8118 3900 8218 3903
rect 8286 3900 8321 3937
rect 8383 3934 8742 3937
rect 8383 3929 8605 3934
rect 8383 3905 8396 3929
rect 8420 3910 8605 3929
rect 8629 3910 8742 3934
rect 8420 3905 8742 3910
rect 8383 3901 8742 3905
rect 8809 3929 8957 3937
rect 8809 3909 8820 3929
rect 8840 3926 8957 3929
rect 9010 3926 9023 3959
rect 8840 3909 9023 3926
rect 8809 3902 9023 3909
rect 8809 3901 8850 3902
rect 8940 3901 9023 3902
rect 8285 3875 8321 3900
rect 8133 3848 8170 3849
rect 8229 3848 8266 3849
rect 8285 3848 8292 3875
rect 8033 3839 8171 3848
rect 8033 3819 8142 3839
rect 8162 3819 8171 3839
rect 8033 3812 8171 3819
rect 8229 3845 8292 3848
rect 8313 3848 8321 3875
rect 8340 3848 8377 3849
rect 8313 3845 8377 3848
rect 8229 3839 8377 3845
rect 8229 3819 8238 3839
rect 8258 3819 8348 3839
rect 8368 3819 8377 3839
rect 8033 3810 8129 3812
rect 8229 3809 8377 3819
rect 8436 3839 8473 3849
rect 8548 3848 8585 3849
rect 8529 3846 8585 3848
rect 8436 3819 8444 3839
rect 8464 3819 8473 3839
rect 8285 3808 8321 3809
rect 8133 3677 8170 3678
rect 8436 3677 8473 3819
rect 8498 3839 8585 3846
rect 8498 3836 8556 3839
rect 8498 3816 8503 3836
rect 8524 3819 8556 3836
rect 8576 3819 8585 3839
rect 8524 3816 8585 3819
rect 8498 3809 8585 3816
rect 8644 3839 8681 3849
rect 8644 3819 8652 3839
rect 8672 3819 8681 3839
rect 8498 3808 8529 3809
rect 8644 3740 8681 3819
rect 8711 3848 8742 3901
rect 8948 3868 8962 3901
rect 9015 3868 9023 3901
rect 8948 3862 9023 3868
rect 8948 3857 9018 3862
rect 8761 3848 8798 3849
rect 8711 3839 8798 3848
rect 8711 3819 8769 3839
rect 8789 3819 8798 3839
rect 8711 3809 8798 3819
rect 8857 3839 8894 3849
rect 9082 3844 9109 4214
rect 9149 3984 9213 3996
rect 9489 3992 9526 4216
rect 9997 4197 10061 4199
rect 9993 4185 10061 4197
rect 9993 4152 10004 4185
rect 10044 4152 10061 4185
rect 9993 4142 10061 4152
rect 9754 4081 9865 4096
rect 9754 4079 9796 4081
rect 9754 4059 9761 4079
rect 9780 4059 9796 4079
rect 9754 4051 9796 4059
rect 9824 4079 9865 4081
rect 9824 4059 9838 4079
rect 9857 4059 9865 4079
rect 9824 4051 9865 4059
rect 9754 4045 9865 4051
rect 9697 4023 9946 4045
rect 9697 3992 9734 4023
rect 9910 4021 9946 4023
rect 9910 3992 9947 4021
rect 9149 3983 9184 3984
rect 9126 3978 9184 3983
rect 9126 3958 9129 3978
rect 9149 3964 9184 3978
rect 9204 3964 9213 3984
rect 9149 3956 9213 3964
rect 9175 3955 9213 3956
rect 9176 3954 9213 3955
rect 9279 3988 9315 3989
rect 9387 3988 9423 3989
rect 9279 3980 9423 3988
rect 9279 3960 9287 3980
rect 9307 3960 9395 3980
rect 9415 3960 9423 3980
rect 9279 3954 9423 3960
rect 9489 3984 9527 3992
rect 9595 3988 9631 3989
rect 9489 3964 9498 3984
rect 9518 3964 9527 3984
rect 9489 3955 9527 3964
rect 9546 3981 9631 3988
rect 9546 3961 9553 3981
rect 9574 3980 9631 3981
rect 9574 3961 9603 3980
rect 9546 3960 9603 3961
rect 9623 3960 9631 3980
rect 9489 3954 9526 3955
rect 9546 3954 9631 3960
rect 9697 3984 9735 3992
rect 9808 3988 9844 3989
rect 9697 3964 9706 3984
rect 9726 3964 9735 3984
rect 9697 3955 9735 3964
rect 9759 3980 9844 3988
rect 9759 3960 9816 3980
rect 9836 3960 9844 3980
rect 9697 3954 9734 3955
rect 9759 3954 9844 3960
rect 9910 3984 9948 3992
rect 9910 3964 9919 3984
rect 9939 3964 9948 3984
rect 9910 3955 9948 3964
rect 9997 3958 10061 4142
rect 10217 4016 10282 4217
rect 11259 4277 11324 4478
rect 11480 4352 11544 4536
rect 11593 4530 11631 4539
rect 11593 4510 11602 4530
rect 11622 4510 11631 4530
rect 11593 4502 11631 4510
rect 11697 4534 11782 4540
rect 11807 4539 11844 4540
rect 11697 4514 11705 4534
rect 11725 4514 11782 4534
rect 11697 4506 11782 4514
rect 11806 4530 11844 4539
rect 11806 4510 11815 4530
rect 11835 4510 11844 4530
rect 11697 4505 11733 4506
rect 11806 4502 11844 4510
rect 11910 4534 11995 4540
rect 12015 4539 12052 4540
rect 11910 4514 11918 4534
rect 11938 4533 11995 4534
rect 11938 4514 11967 4533
rect 11910 4513 11967 4514
rect 11988 4513 11995 4533
rect 11910 4506 11995 4513
rect 12014 4530 12052 4539
rect 12014 4510 12023 4530
rect 12043 4510 12052 4530
rect 11910 4505 11946 4506
rect 12014 4502 12052 4510
rect 12118 4534 12262 4540
rect 12118 4514 12126 4534
rect 12146 4514 12234 4534
rect 12254 4514 12262 4534
rect 12118 4506 12262 4514
rect 12118 4505 12154 4506
rect 12226 4505 12262 4506
rect 12328 4539 12365 4540
rect 12328 4538 12366 4539
rect 12328 4530 12392 4538
rect 12328 4510 12337 4530
rect 12357 4516 12392 4530
rect 12412 4516 12415 4536
rect 12357 4511 12415 4516
rect 12357 4510 12392 4511
rect 11594 4473 11631 4502
rect 11595 4471 11631 4473
rect 11807 4471 11844 4502
rect 11595 4449 11844 4471
rect 11676 4443 11787 4449
rect 11676 4435 11717 4443
rect 11676 4415 11684 4435
rect 11703 4415 11717 4435
rect 11676 4413 11717 4415
rect 11745 4435 11787 4443
rect 11745 4415 11761 4435
rect 11780 4415 11787 4435
rect 11745 4413 11787 4415
rect 11676 4398 11787 4413
rect 11480 4342 11548 4352
rect 11480 4309 11497 4342
rect 11537 4309 11548 4342
rect 11480 4297 11548 4309
rect 11480 4295 11544 4297
rect 12015 4278 12052 4502
rect 12328 4498 12392 4510
rect 12432 4280 12459 4650
rect 12647 4645 12684 4655
rect 12743 4675 12830 4685
rect 12743 4655 12752 4675
rect 12772 4655 12830 4675
rect 12743 4646 12830 4655
rect 12743 4645 12780 4646
rect 12523 4632 12593 4637
rect 12518 4626 12593 4632
rect 12518 4593 12526 4626
rect 12579 4593 12593 4626
rect 12799 4593 12830 4646
rect 12860 4675 12897 4754
rect 13012 4685 13043 4686
rect 12860 4655 12869 4675
rect 12889 4655 12897 4675
rect 12860 4645 12897 4655
rect 12956 4678 13043 4685
rect 12956 4675 13017 4678
rect 12956 4655 12965 4675
rect 12985 4658 13017 4675
rect 13038 4658 13043 4678
rect 12985 4655 13043 4658
rect 12956 4648 13043 4655
rect 13068 4675 13105 4817
rect 13371 4816 13408 4817
rect 13220 4685 13256 4686
rect 13068 4655 13077 4675
rect 13097 4655 13105 4675
rect 12956 4646 13012 4648
rect 12956 4645 12993 4646
rect 13068 4645 13105 4655
rect 13164 4675 13312 4685
rect 13412 4682 13508 4684
rect 13164 4655 13173 4675
rect 13193 4655 13283 4675
rect 13303 4655 13312 4675
rect 13164 4649 13312 4655
rect 13164 4646 13228 4649
rect 13164 4645 13201 4646
rect 13220 4619 13228 4646
rect 13249 4646 13312 4649
rect 13370 4675 13508 4682
rect 13370 4655 13379 4675
rect 13399 4655 13508 4675
rect 13370 4646 13508 4655
rect 13249 4619 13256 4646
rect 13275 4645 13312 4646
rect 13371 4645 13408 4646
rect 13220 4594 13256 4619
rect 12518 4592 12601 4593
rect 12691 4592 12732 4593
rect 12518 4585 12732 4592
rect 12518 4568 12701 4585
rect 12518 4535 12531 4568
rect 12584 4565 12701 4568
rect 12721 4565 12732 4585
rect 12584 4557 12732 4565
rect 12799 4589 13158 4593
rect 12799 4584 13121 4589
rect 12799 4560 12912 4584
rect 12936 4565 13121 4584
rect 13145 4565 13158 4589
rect 12936 4560 13158 4565
rect 12799 4557 13158 4560
rect 13220 4557 13255 4594
rect 13323 4591 13423 4594
rect 13323 4587 13390 4591
rect 13323 4561 13335 4587
rect 13361 4565 13390 4587
rect 13416 4565 13423 4591
rect 13361 4561 13423 4565
rect 13323 4557 13423 4561
rect 12584 4535 12601 4557
rect 12799 4536 12830 4557
rect 13220 4536 13256 4557
rect 12642 4535 12679 4536
rect 12518 4521 12601 4535
rect 12291 4278 12459 4280
rect 12015 4277 12459 4278
rect 11259 4247 12459 4277
rect 12529 4311 12601 4521
rect 12641 4526 12679 4535
rect 12641 4506 12650 4526
rect 12670 4506 12679 4526
rect 12641 4498 12679 4506
rect 12745 4530 12830 4536
rect 12855 4535 12892 4536
rect 12745 4510 12753 4530
rect 12773 4510 12830 4530
rect 12745 4502 12830 4510
rect 12854 4526 12892 4535
rect 12854 4506 12863 4526
rect 12883 4506 12892 4526
rect 12745 4501 12781 4502
rect 12854 4498 12892 4506
rect 12958 4530 13043 4536
rect 13063 4535 13100 4536
rect 12958 4510 12966 4530
rect 12986 4529 13043 4530
rect 12986 4510 13015 4529
rect 12958 4509 13015 4510
rect 13036 4509 13043 4529
rect 12958 4502 13043 4509
rect 13062 4526 13100 4535
rect 13062 4506 13071 4526
rect 13091 4506 13100 4526
rect 12958 4501 12994 4502
rect 13062 4498 13100 4506
rect 13166 4530 13310 4536
rect 13166 4510 13174 4530
rect 13194 4510 13282 4530
rect 13302 4510 13310 4530
rect 13166 4502 13310 4510
rect 13166 4501 13202 4502
rect 13274 4501 13310 4502
rect 13376 4535 13413 4536
rect 13376 4534 13414 4535
rect 13376 4526 13440 4534
rect 13376 4506 13385 4526
rect 13405 4512 13440 4526
rect 13460 4512 13463 4532
rect 13405 4507 13463 4512
rect 13405 4506 13440 4507
rect 12642 4469 12679 4498
rect 12643 4467 12679 4469
rect 12855 4467 12892 4498
rect 12643 4445 12892 4467
rect 12724 4439 12835 4445
rect 12724 4431 12765 4439
rect 12724 4411 12732 4431
rect 12751 4411 12765 4431
rect 12724 4409 12765 4411
rect 12793 4431 12835 4439
rect 12793 4411 12809 4431
rect 12828 4411 12835 4431
rect 12793 4409 12835 4411
rect 12724 4394 12835 4409
rect 12529 4272 12548 4311
rect 12593 4272 12601 4311
rect 12529 4255 12601 4272
rect 13063 4299 13100 4498
rect 13376 4494 13440 4506
rect 13063 4293 13104 4299
rect 13480 4295 13507 4646
rect 13636 4598 13707 5077
rect 13636 4514 13705 4598
rect 13339 4293 13507 4295
rect 13063 4267 13507 4293
rect 11259 4200 11324 4247
rect 11259 4182 11282 4200
rect 11300 4182 11324 4200
rect 12172 4227 12207 4229
rect 12172 4225 12276 4227
rect 13065 4225 13104 4267
rect 13339 4266 13507 4267
rect 12172 4218 13106 4225
rect 12172 4217 12223 4218
rect 12172 4197 12175 4217
rect 12200 4198 12223 4217
rect 12255 4198 13106 4218
rect 12200 4197 13106 4198
rect 12172 4190 13106 4197
rect 12445 4189 13106 4190
rect 11259 4161 11324 4182
rect 11536 4172 11576 4175
rect 11536 4168 12439 4172
rect 11536 4148 12413 4168
rect 12433 4148 12439 4168
rect 11536 4145 12439 4148
rect 11260 4101 11325 4121
rect 11260 4083 11284 4101
rect 11302 4083 11325 4101
rect 11260 4056 11325 4083
rect 11536 4056 11576 4145
rect 12020 4143 12436 4145
rect 12020 4142 12361 4143
rect 11677 4111 11787 4125
rect 11677 4108 11720 4111
rect 11677 4103 11681 4108
rect 11259 4021 11576 4056
rect 11599 4081 11681 4103
rect 11710 4081 11720 4108
rect 11748 4084 11755 4111
rect 11784 4103 11787 4111
rect 11784 4084 11849 4103
rect 11748 4081 11849 4084
rect 11599 4079 11849 4081
rect 10217 3998 10239 4016
rect 10257 3998 10282 4016
rect 10217 3979 10282 3998
rect 9910 3954 9947 3955
rect 9333 3933 9369 3954
rect 9759 3933 9790 3954
rect 9997 3949 10005 3958
rect 9994 3933 10005 3949
rect 9166 3929 9266 3933
rect 9166 3925 9228 3929
rect 9166 3899 9173 3925
rect 9199 3903 9228 3925
rect 9254 3903 9266 3929
rect 9199 3899 9266 3903
rect 9166 3896 9266 3899
rect 9334 3896 9369 3933
rect 9431 3930 9790 3933
rect 9431 3925 9653 3930
rect 9431 3901 9444 3925
rect 9468 3906 9653 3925
rect 9677 3906 9790 3930
rect 9468 3901 9790 3906
rect 9431 3897 9790 3901
rect 9857 3925 10005 3933
rect 9857 3905 9868 3925
rect 9888 3916 10005 3925
rect 10054 3949 10061 3958
rect 10054 3916 10062 3949
rect 11260 3945 11325 4021
rect 11599 4000 11636 4079
rect 11677 4066 11787 4079
rect 11751 4010 11782 4011
rect 11599 3980 11608 4000
rect 11628 3980 11636 4000
rect 11599 3970 11636 3980
rect 11695 4000 11782 4010
rect 11695 3980 11704 4000
rect 11724 3980 11782 4000
rect 11695 3971 11782 3980
rect 11695 3970 11732 3971
rect 9888 3905 10062 3916
rect 9857 3898 10062 3905
rect 9857 3897 9898 3898
rect 9333 3871 9369 3896
rect 9181 3844 9218 3845
rect 9277 3844 9314 3845
rect 9333 3844 9340 3871
rect 8857 3819 8865 3839
rect 8885 3819 8894 3839
rect 8711 3808 8742 3809
rect 8706 3740 8816 3753
rect 8857 3740 8894 3819
rect 9081 3835 9219 3844
rect 9081 3815 9190 3835
rect 9210 3815 9219 3835
rect 9081 3808 9219 3815
rect 9277 3841 9340 3844
rect 9361 3844 9369 3871
rect 9388 3844 9425 3845
rect 9361 3841 9425 3844
rect 9277 3835 9425 3841
rect 9277 3815 9286 3835
rect 9306 3815 9396 3835
rect 9416 3815 9425 3835
rect 9081 3806 9177 3808
rect 9277 3805 9425 3815
rect 9484 3835 9521 3845
rect 9596 3844 9633 3845
rect 9577 3842 9633 3844
rect 9484 3815 9492 3835
rect 9512 3815 9521 3835
rect 9333 3804 9369 3805
rect 8644 3738 8894 3740
rect 8644 3735 8745 3738
rect 8644 3716 8709 3735
rect 8706 3708 8709 3716
rect 8738 3708 8745 3735
rect 8773 3711 8783 3738
rect 8812 3716 8894 3738
rect 8812 3711 8816 3716
rect 8773 3708 8816 3711
rect 8706 3694 8816 3708
rect 8132 3676 8473 3677
rect 8057 3671 8473 3676
rect 9181 3673 9218 3674
rect 9484 3673 9521 3815
rect 9546 3835 9633 3842
rect 9546 3832 9604 3835
rect 9546 3812 9551 3832
rect 9572 3815 9604 3832
rect 9624 3815 9633 3835
rect 9572 3812 9633 3815
rect 9546 3805 9633 3812
rect 9692 3835 9729 3845
rect 9692 3815 9700 3835
rect 9720 3815 9729 3835
rect 9546 3804 9577 3805
rect 9692 3736 9729 3815
rect 9759 3844 9790 3897
rect 9994 3895 10062 3898
rect 9994 3853 10006 3895
rect 10055 3853 10062 3895
rect 9809 3844 9846 3845
rect 9759 3835 9846 3844
rect 9759 3815 9817 3835
rect 9837 3815 9846 3835
rect 9759 3805 9846 3815
rect 9905 3835 9942 3845
rect 9994 3840 10062 3853
rect 10217 3917 10282 3934
rect 10217 3899 10241 3917
rect 10259 3899 10282 3917
rect 11260 3927 11282 3945
rect 11300 3927 11325 3945
rect 11260 3906 11325 3927
rect 11473 3925 11538 3934
rect 9905 3815 9913 3835
rect 9933 3815 9942 3835
rect 9759 3804 9790 3805
rect 9754 3736 9864 3749
rect 9905 3736 9942 3815
rect 10217 3760 10282 3899
rect 11473 3888 11483 3925
rect 11523 3917 11538 3925
rect 11751 3918 11782 3971
rect 11812 4000 11849 4079
rect 11964 4010 11995 4011
rect 11812 3980 11821 4000
rect 11841 3980 11849 4000
rect 11812 3970 11849 3980
rect 11908 4003 11995 4010
rect 11908 4000 11969 4003
rect 11908 3980 11917 4000
rect 11937 3983 11969 4000
rect 11990 3983 11995 4003
rect 11937 3980 11995 3983
rect 11908 3973 11995 3980
rect 12020 4000 12057 4142
rect 12323 4141 12360 4142
rect 12172 4010 12208 4011
rect 12020 3980 12029 4000
rect 12049 3980 12057 4000
rect 11908 3971 11964 3973
rect 11908 3970 11945 3971
rect 12020 3970 12057 3980
rect 12116 4000 12264 4010
rect 12364 4007 12460 4009
rect 12116 3980 12125 4000
rect 12145 3980 12235 4000
rect 12255 3980 12264 4000
rect 12116 3974 12264 3980
rect 12116 3971 12180 3974
rect 12116 3970 12153 3971
rect 12172 3944 12180 3971
rect 12201 3971 12264 3974
rect 12322 4000 12460 4007
rect 13640 4002 13702 4514
rect 12322 3980 12331 4000
rect 12351 3980 12460 4000
rect 12322 3971 12460 3980
rect 12201 3944 12208 3971
rect 12227 3970 12264 3971
rect 12323 3970 12360 3971
rect 12172 3919 12208 3944
rect 11643 3917 11684 3918
rect 11523 3910 11684 3917
rect 11523 3890 11653 3910
rect 11673 3890 11684 3910
rect 11523 3888 11684 3890
rect 11473 3882 11684 3888
rect 11751 3914 12110 3918
rect 11751 3909 12073 3914
rect 11751 3885 11864 3909
rect 11888 3890 12073 3909
rect 12097 3890 12110 3914
rect 11888 3885 12110 3890
rect 11751 3882 12110 3885
rect 12172 3882 12207 3919
rect 12275 3916 12375 3919
rect 12275 3912 12342 3916
rect 12275 3886 12287 3912
rect 12313 3890 12342 3912
rect 12368 3890 12375 3916
rect 12313 3886 12375 3890
rect 12275 3882 12375 3886
rect 11473 3869 11540 3882
rect 10217 3754 10239 3760
rect 9692 3734 9942 3736
rect 9692 3731 9793 3734
rect 9692 3712 9757 3731
rect 9754 3704 9757 3712
rect 9786 3704 9793 3731
rect 9821 3707 9831 3734
rect 9860 3712 9942 3734
rect 9971 3742 10239 3754
rect 10257 3742 10282 3760
rect 9971 3719 10282 3742
rect 11265 3846 11321 3866
rect 11265 3828 11284 3846
rect 11302 3828 11321 3846
rect 9971 3718 10026 3719
rect 9860 3707 9864 3712
rect 9821 3704 9864 3707
rect 9754 3690 9864 3704
rect 9180 3672 9521 3673
rect 8057 3651 8060 3671
rect 8080 3651 8473 3671
rect 9105 3671 9521 3672
rect 9971 3671 10014 3718
rect 11265 3715 11321 3828
rect 11473 3848 11487 3869
rect 11523 3848 11540 3869
rect 11751 3861 11782 3882
rect 12172 3861 12208 3882
rect 11594 3860 11631 3861
rect 11473 3841 11540 3848
rect 11593 3851 11631 3860
rect 9105 3667 10014 3671
rect 8424 3618 8469 3651
rect 9105 3647 9108 3667
rect 9128 3647 10014 3667
rect 9482 3642 10014 3647
rect 10222 3661 10281 3683
rect 10222 3643 10241 3661
rect 10259 3643 10281 3661
rect 9270 3618 9369 3620
rect 8424 3608 9369 3618
rect 8424 3582 9292 3608
rect 8425 3581 9292 3582
rect 9270 3570 9292 3581
rect 9317 3573 9336 3608
rect 9361 3573 9369 3608
rect 9317 3570 9369 3573
rect 10222 3572 10281 3643
rect 11265 3577 11320 3715
rect 11473 3689 11538 3841
rect 11593 3831 11602 3851
rect 11622 3831 11631 3851
rect 11593 3823 11631 3831
rect 11697 3855 11782 3861
rect 11807 3860 11844 3861
rect 11697 3835 11705 3855
rect 11725 3835 11782 3855
rect 11697 3827 11782 3835
rect 11806 3851 11844 3860
rect 11806 3831 11815 3851
rect 11835 3831 11844 3851
rect 11697 3826 11733 3827
rect 11806 3823 11844 3831
rect 11910 3855 11995 3861
rect 12015 3860 12052 3861
rect 11910 3835 11918 3855
rect 11938 3854 11995 3855
rect 11938 3835 11967 3854
rect 11910 3834 11967 3835
rect 11988 3834 11995 3854
rect 11910 3827 11995 3834
rect 12014 3851 12052 3860
rect 12014 3831 12023 3851
rect 12043 3831 12052 3851
rect 11910 3826 11946 3827
rect 12014 3823 12052 3831
rect 12118 3855 12262 3861
rect 12118 3835 12126 3855
rect 12146 3835 12234 3855
rect 12254 3835 12262 3855
rect 12118 3827 12262 3835
rect 12118 3826 12154 3827
rect 12226 3826 12262 3827
rect 12328 3860 12365 3861
rect 12328 3859 12366 3860
rect 12328 3851 12392 3859
rect 12328 3831 12337 3851
rect 12357 3837 12392 3851
rect 12412 3837 12415 3857
rect 12357 3832 12415 3837
rect 12357 3831 12392 3832
rect 11594 3794 11631 3823
rect 11595 3792 11631 3794
rect 11807 3792 11844 3823
rect 11595 3770 11844 3792
rect 11676 3764 11787 3770
rect 11676 3756 11717 3764
rect 11676 3736 11684 3756
rect 11703 3736 11717 3756
rect 11676 3734 11717 3736
rect 11745 3756 11787 3764
rect 11745 3736 11761 3756
rect 11780 3736 11787 3756
rect 11745 3734 11787 3736
rect 11676 3721 11787 3734
rect 12015 3724 12052 3823
rect 12328 3819 12392 3831
rect 11466 3679 11587 3689
rect 11466 3677 11535 3679
rect 11466 3636 11479 3677
rect 11516 3638 11535 3677
rect 11572 3638 11587 3679
rect 11516 3636 11587 3638
rect 11466 3618 11587 3636
rect 11258 3574 11322 3577
rect 11678 3574 11782 3580
rect 12013 3574 12054 3724
rect 12432 3716 12459 3971
rect 12521 3961 12601 3972
rect 12521 3935 12538 3961
rect 12578 3935 12601 3961
rect 12521 3908 12601 3935
rect 13644 3963 13702 4002
rect 13644 3928 13706 3963
rect 12521 3882 12542 3908
rect 12582 3882 12601 3908
rect 12521 3863 12601 3882
rect 12521 3837 12545 3863
rect 12585 3837 12601 3863
rect 12521 3786 12601 3837
rect 13593 3901 13706 3928
rect 13593 3899 13652 3901
rect 13593 3868 13607 3899
rect 13632 3878 13652 3899
rect 13678 3878 13706 3901
rect 13632 3868 13706 3878
rect 13593 3858 13706 3868
rect 9270 3562 9369 3570
rect 9296 3561 9368 3562
rect 8950 3535 9017 3554
rect 8950 3514 8967 3535
rect 7831 3336 7911 3378
rect 8948 3469 8967 3514
rect 8997 3514 9017 3535
rect 8997 3469 9018 3514
rect 9487 3511 9528 3513
rect 9759 3511 9863 3513
rect 10219 3511 10283 3572
rect 6892 3225 6928 3226
rect 6784 3217 6928 3225
rect 6784 3197 6792 3217
rect 6812 3197 6900 3217
rect 6920 3197 6928 3217
rect 6784 3191 6928 3197
rect 6994 3221 7032 3229
rect 7100 3225 7136 3226
rect 6994 3201 7003 3221
rect 7023 3201 7032 3221
rect 6994 3192 7032 3201
rect 7051 3218 7136 3225
rect 7051 3198 7058 3218
rect 7079 3217 7136 3218
rect 7079 3198 7108 3217
rect 7051 3197 7108 3198
rect 7128 3197 7136 3217
rect 6994 3191 7031 3192
rect 7051 3191 7136 3197
rect 7202 3221 7240 3229
rect 7313 3225 7349 3226
rect 7202 3201 7211 3221
rect 7231 3201 7240 3221
rect 7202 3192 7240 3201
rect 7264 3217 7349 3225
rect 7264 3197 7321 3217
rect 7341 3197 7349 3217
rect 7202 3191 7239 3192
rect 7264 3191 7349 3197
rect 7415 3221 7453 3229
rect 7415 3201 7424 3221
rect 7444 3201 7453 3221
rect 7415 3192 7453 3201
rect 7653 3209 7739 3245
rect 7415 3191 7452 3192
rect 6838 3170 6874 3191
rect 7264 3170 7295 3191
rect 7491 3170 7537 3174
rect 6671 3166 6771 3170
rect 6671 3162 6733 3166
rect 6671 3136 6678 3162
rect 6704 3140 6733 3162
rect 6759 3140 6771 3166
rect 6704 3136 6771 3140
rect 6671 3133 6771 3136
rect 6839 3133 6874 3170
rect 6936 3167 7295 3170
rect 6936 3162 7158 3167
rect 6936 3138 6949 3162
rect 6973 3143 7158 3162
rect 7182 3143 7295 3167
rect 6973 3138 7295 3143
rect 6936 3134 7295 3138
rect 7362 3162 7537 3170
rect 7362 3142 7373 3162
rect 7393 3142 7537 3162
rect 7653 3168 7670 3209
rect 7724 3168 7739 3209
rect 7653 3149 7739 3168
rect 7362 3135 7537 3142
rect 7362 3134 7403 3135
rect 6838 3108 6874 3133
rect 6686 3081 6723 3082
rect 6782 3081 6819 3082
rect 6838 3081 6845 3108
rect 6586 3072 6724 3081
rect 6586 3052 6695 3072
rect 6715 3052 6724 3072
rect 6586 3045 6724 3052
rect 6782 3078 6845 3081
rect 6866 3081 6874 3108
rect 6893 3081 6930 3082
rect 6866 3078 6930 3081
rect 6782 3072 6930 3078
rect 6782 3052 6791 3072
rect 6811 3052 6901 3072
rect 6921 3052 6930 3072
rect 6586 3043 6682 3045
rect 6782 3042 6930 3052
rect 6989 3072 7026 3082
rect 7101 3081 7138 3082
rect 7082 3079 7138 3081
rect 6989 3052 6997 3072
rect 7017 3052 7026 3072
rect 6838 3041 6874 3042
rect 6686 2910 6723 2911
rect 6989 2910 7026 3052
rect 7051 3072 7138 3079
rect 7051 3069 7109 3072
rect 7051 3049 7056 3069
rect 7077 3052 7109 3069
rect 7129 3052 7138 3072
rect 7077 3049 7138 3052
rect 7051 3042 7138 3049
rect 7197 3072 7234 3082
rect 7197 3052 7205 3072
rect 7225 3052 7234 3072
rect 7051 3041 7082 3042
rect 7197 2973 7234 3052
rect 7264 3081 7295 3134
rect 7314 3081 7351 3082
rect 7264 3072 7351 3081
rect 7264 3052 7322 3072
rect 7342 3052 7351 3072
rect 7264 3042 7351 3052
rect 7410 3072 7447 3082
rect 7410 3052 7418 3072
rect 7438 3052 7447 3072
rect 7264 3041 7295 3042
rect 7259 2973 7369 2986
rect 7410 2973 7447 3052
rect 7491 3052 7537 3135
rect 7831 3052 7906 3336
rect 8948 3261 9018 3469
rect 9080 3476 10283 3511
rect 9080 3462 9108 3476
rect 9082 3331 9108 3462
rect 9487 3473 10283 3476
rect 11258 3571 12054 3574
rect 12433 3585 12459 3716
rect 12433 3571 12461 3585
rect 11258 3536 12461 3571
rect 12523 3578 12593 3786
rect 11258 3475 11322 3536
rect 11678 3534 11782 3536
rect 12013 3534 12054 3536
rect 12523 3533 12544 3578
rect 12524 3512 12544 3533
rect 12574 3533 12593 3578
rect 12574 3512 12591 3533
rect 12524 3493 12591 3512
rect 12173 3485 12245 3486
rect 12172 3477 12271 3485
rect 8940 3210 9020 3261
rect 8940 3184 8956 3210
rect 8996 3184 9020 3210
rect 8940 3165 9020 3184
rect 8940 3139 8959 3165
rect 8999 3139 9020 3165
rect 8940 3112 9020 3139
rect 8940 3086 8963 3112
rect 9003 3086 9020 3112
rect 8940 3075 9020 3086
rect 9082 3076 9109 3331
rect 9487 3323 9528 3473
rect 9759 3467 9863 3473
rect 10219 3470 10283 3473
rect 9954 3411 10075 3429
rect 9954 3409 10025 3411
rect 9954 3368 9969 3409
rect 10006 3370 10025 3409
rect 10062 3370 10075 3411
rect 10006 3368 10075 3370
rect 9954 3358 10075 3368
rect 9149 3216 9213 3228
rect 9489 3224 9526 3323
rect 9754 3313 9865 3326
rect 9754 3311 9796 3313
rect 9754 3291 9761 3311
rect 9780 3291 9796 3311
rect 9754 3283 9796 3291
rect 9824 3311 9865 3313
rect 9824 3291 9838 3311
rect 9857 3291 9865 3311
rect 9824 3283 9865 3291
rect 9754 3277 9865 3283
rect 9697 3255 9946 3277
rect 9697 3224 9734 3255
rect 9910 3253 9946 3255
rect 9910 3224 9947 3253
rect 9149 3215 9184 3216
rect 9126 3210 9184 3215
rect 9126 3190 9129 3210
rect 9149 3196 9184 3210
rect 9204 3196 9213 3216
rect 9149 3188 9213 3196
rect 9175 3187 9213 3188
rect 9176 3186 9213 3187
rect 9279 3220 9315 3221
rect 9387 3220 9423 3221
rect 9279 3212 9423 3220
rect 9279 3192 9287 3212
rect 9307 3192 9395 3212
rect 9415 3192 9423 3212
rect 9279 3186 9423 3192
rect 9489 3216 9527 3224
rect 9595 3220 9631 3221
rect 9489 3196 9498 3216
rect 9518 3196 9527 3216
rect 9489 3187 9527 3196
rect 9546 3213 9631 3220
rect 9546 3193 9553 3213
rect 9574 3212 9631 3213
rect 9574 3193 9603 3212
rect 9546 3192 9603 3193
rect 9623 3192 9631 3212
rect 9489 3186 9526 3187
rect 9546 3186 9631 3192
rect 9697 3216 9735 3224
rect 9808 3220 9844 3221
rect 9697 3196 9706 3216
rect 9726 3196 9735 3216
rect 9697 3187 9735 3196
rect 9759 3212 9844 3220
rect 9759 3192 9816 3212
rect 9836 3192 9844 3212
rect 9697 3186 9734 3187
rect 9759 3186 9844 3192
rect 9910 3216 9948 3224
rect 9910 3196 9919 3216
rect 9939 3196 9948 3216
rect 10003 3206 10068 3358
rect 10221 3332 10276 3470
rect 11260 3404 11319 3475
rect 12172 3474 12224 3477
rect 12172 3439 12180 3474
rect 12205 3439 12224 3474
rect 12249 3466 12271 3477
rect 12249 3465 13116 3466
rect 12249 3439 13117 3465
rect 12172 3429 13117 3439
rect 12172 3427 12271 3429
rect 11260 3386 11282 3404
rect 11300 3386 11319 3404
rect 11260 3364 11319 3386
rect 11527 3400 12059 3405
rect 11527 3380 12413 3400
rect 12433 3380 12436 3400
rect 13072 3396 13117 3429
rect 11527 3376 12436 3380
rect 9910 3187 9948 3196
rect 10001 3199 10068 3206
rect 9910 3186 9947 3187
rect 9333 3165 9369 3186
rect 9759 3165 9790 3186
rect 10001 3178 10018 3199
rect 10054 3178 10068 3199
rect 10220 3219 10276 3332
rect 11527 3329 11570 3376
rect 12020 3375 12436 3376
rect 13068 3376 13461 3396
rect 13481 3376 13484 3396
rect 12020 3374 12361 3375
rect 11677 3343 11787 3357
rect 11677 3340 11720 3343
rect 11677 3335 11681 3340
rect 11515 3328 11570 3329
rect 10220 3201 10239 3219
rect 10257 3201 10276 3219
rect 10220 3181 10276 3201
rect 11259 3305 11570 3328
rect 11259 3287 11284 3305
rect 11302 3293 11570 3305
rect 11599 3313 11681 3335
rect 11710 3313 11720 3340
rect 11748 3316 11755 3343
rect 11784 3335 11787 3343
rect 11784 3316 11849 3335
rect 11748 3313 11849 3316
rect 11599 3311 11849 3313
rect 11302 3287 11324 3293
rect 10001 3165 10068 3178
rect 9166 3161 9266 3165
rect 9166 3157 9228 3161
rect 9166 3131 9173 3157
rect 9199 3135 9228 3157
rect 9254 3135 9266 3161
rect 9199 3131 9266 3135
rect 9166 3128 9266 3131
rect 9334 3128 9369 3165
rect 9431 3162 9790 3165
rect 9431 3157 9653 3162
rect 9431 3133 9444 3157
rect 9468 3138 9653 3157
rect 9677 3138 9790 3162
rect 9468 3133 9790 3138
rect 9431 3129 9790 3133
rect 9857 3159 10068 3165
rect 9857 3157 10018 3159
rect 9857 3137 9868 3157
rect 9888 3137 10018 3157
rect 9857 3130 10018 3137
rect 9857 3129 9898 3130
rect 9333 3103 9369 3128
rect 9181 3076 9218 3077
rect 9277 3076 9314 3077
rect 9333 3076 9340 3103
rect 7491 3017 7906 3052
rect 9081 3067 9219 3076
rect 9081 3047 9190 3067
rect 9210 3047 9219 3067
rect 9081 3040 9219 3047
rect 9277 3073 9340 3076
rect 9361 3076 9369 3103
rect 9388 3076 9425 3077
rect 9361 3073 9425 3076
rect 9277 3067 9425 3073
rect 9277 3047 9286 3067
rect 9306 3047 9396 3067
rect 9416 3047 9425 3067
rect 9081 3038 9177 3040
rect 9277 3037 9425 3047
rect 9484 3067 9521 3077
rect 9596 3076 9633 3077
rect 9577 3074 9633 3076
rect 9484 3047 9492 3067
rect 9512 3047 9521 3067
rect 9333 3036 9369 3037
rect 7491 3016 7537 3017
rect 7197 2971 7447 2973
rect 7197 2968 7298 2971
rect 7197 2949 7262 2968
rect 7259 2941 7262 2949
rect 7291 2941 7298 2968
rect 7326 2944 7336 2971
rect 7365 2949 7447 2971
rect 7831 2965 7906 3017
rect 7365 2944 7369 2949
rect 7326 2941 7369 2944
rect 7259 2927 7369 2941
rect 6685 2909 7026 2910
rect 6610 2904 7026 2909
rect 6610 2884 6613 2904
rect 6633 2884 7027 2904
rect 3090 2475 6158 2500
rect 3090 2410 5953 2475
rect 6084 2410 6158 2475
rect 3090 2393 6158 2410
rect 6984 2380 7027 2884
rect 7644 2795 7739 2815
rect 7644 2751 7664 2795
rect 7724 2751 7739 2795
rect 7644 2455 7739 2751
rect 7644 2414 7677 2455
rect 7713 2414 7739 2455
rect 7839 2494 7901 2965
rect 9181 2905 9218 2906
rect 9484 2905 9521 3047
rect 9546 3067 9633 3074
rect 9546 3064 9604 3067
rect 9546 3044 9551 3064
rect 9572 3047 9604 3064
rect 9624 3047 9633 3067
rect 9572 3044 9633 3047
rect 9546 3037 9633 3044
rect 9692 3067 9729 3077
rect 9692 3047 9700 3067
rect 9720 3047 9729 3067
rect 9546 3036 9577 3037
rect 9692 2968 9729 3047
rect 9759 3076 9790 3129
rect 10003 3122 10018 3130
rect 10058 3122 10068 3159
rect 11259 3148 11324 3287
rect 11599 3232 11636 3311
rect 11677 3298 11787 3311
rect 11751 3242 11782 3243
rect 11599 3212 11608 3232
rect 11628 3212 11636 3232
rect 10003 3113 10068 3122
rect 10216 3120 10281 3141
rect 10216 3102 10241 3120
rect 10259 3102 10281 3120
rect 11259 3130 11282 3148
rect 11300 3130 11324 3148
rect 11259 3113 11324 3130
rect 11479 3194 11547 3207
rect 11599 3202 11636 3212
rect 11695 3232 11782 3242
rect 11695 3212 11704 3232
rect 11724 3212 11782 3232
rect 11695 3203 11782 3212
rect 11695 3202 11732 3203
rect 11479 3152 11486 3194
rect 11535 3152 11547 3194
rect 11479 3149 11547 3152
rect 11751 3150 11782 3203
rect 11812 3232 11849 3311
rect 11964 3242 11995 3243
rect 11812 3212 11821 3232
rect 11841 3212 11849 3232
rect 11812 3202 11849 3212
rect 11908 3235 11995 3242
rect 11908 3232 11969 3235
rect 11908 3212 11917 3232
rect 11937 3215 11969 3232
rect 11990 3215 11995 3235
rect 11937 3212 11995 3215
rect 11908 3205 11995 3212
rect 12020 3232 12057 3374
rect 12323 3373 12360 3374
rect 13068 3371 13484 3376
rect 13068 3370 13409 3371
rect 12725 3339 12835 3353
rect 12725 3336 12768 3339
rect 12725 3331 12729 3336
rect 12647 3309 12729 3331
rect 12758 3309 12768 3336
rect 12796 3312 12803 3339
rect 12832 3331 12835 3339
rect 12832 3312 12897 3331
rect 12796 3309 12897 3312
rect 12647 3307 12897 3309
rect 12172 3242 12208 3243
rect 12020 3212 12029 3232
rect 12049 3212 12057 3232
rect 11908 3203 11964 3205
rect 11908 3202 11945 3203
rect 12020 3202 12057 3212
rect 12116 3232 12264 3242
rect 12364 3239 12460 3241
rect 12116 3212 12125 3232
rect 12145 3212 12235 3232
rect 12255 3212 12264 3232
rect 12116 3206 12264 3212
rect 12116 3203 12180 3206
rect 12116 3202 12153 3203
rect 12172 3176 12180 3203
rect 12201 3203 12264 3206
rect 12322 3232 12460 3239
rect 12322 3212 12331 3232
rect 12351 3212 12460 3232
rect 12322 3203 12460 3212
rect 12647 3228 12684 3307
rect 12725 3294 12835 3307
rect 12799 3238 12830 3239
rect 12647 3208 12656 3228
rect 12676 3208 12684 3228
rect 12201 3176 12208 3203
rect 12227 3202 12264 3203
rect 12323 3202 12360 3203
rect 12172 3151 12208 3176
rect 11643 3149 11684 3150
rect 11479 3142 11684 3149
rect 11479 3131 11653 3142
rect 9809 3076 9846 3077
rect 9759 3067 9846 3076
rect 9759 3047 9817 3067
rect 9837 3047 9846 3067
rect 9759 3037 9846 3047
rect 9905 3067 9942 3077
rect 9905 3047 9913 3067
rect 9933 3047 9942 3067
rect 9759 3036 9790 3037
rect 9754 2968 9864 2981
rect 9905 2968 9942 3047
rect 10216 3026 10281 3102
rect 11479 3098 11487 3131
rect 11480 3089 11487 3098
rect 11536 3122 11653 3131
rect 11673 3122 11684 3142
rect 11536 3114 11684 3122
rect 11751 3146 12110 3150
rect 11751 3141 12073 3146
rect 11751 3117 11864 3141
rect 11888 3122 12073 3141
rect 12097 3122 12110 3146
rect 11888 3117 12110 3122
rect 11751 3114 12110 3117
rect 12172 3114 12207 3151
rect 12275 3148 12375 3151
rect 12275 3144 12342 3148
rect 12275 3118 12287 3144
rect 12313 3122 12342 3144
rect 12368 3122 12375 3148
rect 12313 3118 12375 3122
rect 12275 3114 12375 3118
rect 11536 3098 11547 3114
rect 11536 3089 11544 3098
rect 11751 3093 11782 3114
rect 12172 3093 12208 3114
rect 11594 3092 11631 3093
rect 11259 3049 11324 3068
rect 11259 3031 11284 3049
rect 11302 3031 11324 3049
rect 9692 2966 9942 2968
rect 9692 2963 9793 2966
rect 9692 2944 9757 2963
rect 9754 2936 9757 2944
rect 9786 2936 9793 2963
rect 9821 2939 9831 2966
rect 9860 2944 9942 2966
rect 9965 2991 10282 3026
rect 9860 2939 9864 2944
rect 9821 2936 9864 2939
rect 9754 2922 9864 2936
rect 9180 2904 9521 2905
rect 9105 2902 9521 2904
rect 9965 2902 10005 2991
rect 10216 2964 10281 2991
rect 10216 2946 10239 2964
rect 10257 2946 10281 2964
rect 10216 2926 10281 2946
rect 9102 2899 10005 2902
rect 9102 2879 9108 2899
rect 9128 2879 10005 2899
rect 9102 2875 10005 2879
rect 9965 2872 10005 2875
rect 10217 2865 10282 2886
rect 8435 2857 9096 2858
rect 8435 2850 9369 2857
rect 8435 2849 9341 2850
rect 8435 2829 9286 2849
rect 9318 2830 9341 2849
rect 9366 2830 9369 2850
rect 9318 2829 9369 2830
rect 8435 2822 9369 2829
rect 8034 2780 8202 2781
rect 8437 2780 8476 2822
rect 9265 2820 9369 2822
rect 9334 2818 9369 2820
rect 10217 2847 10241 2865
rect 10259 2847 10282 2865
rect 10217 2800 10282 2847
rect 8034 2754 8478 2780
rect 8034 2752 8202 2754
rect 7839 2475 7903 2494
rect 7839 2436 7856 2475
rect 7890 2436 7903 2475
rect 7839 2417 7903 2436
rect 7644 2388 7739 2414
rect 8034 2401 8061 2752
rect 8437 2748 8478 2754
rect 8101 2541 8165 2553
rect 8441 2549 8478 2748
rect 8940 2775 9012 2792
rect 8940 2736 8948 2775
rect 8993 2736 9012 2775
rect 8706 2638 8817 2653
rect 8706 2636 8748 2638
rect 8706 2616 8713 2636
rect 8732 2616 8748 2636
rect 8706 2608 8748 2616
rect 8776 2636 8817 2638
rect 8776 2616 8790 2636
rect 8809 2616 8817 2636
rect 8776 2608 8817 2616
rect 8706 2602 8817 2608
rect 8649 2580 8898 2602
rect 8649 2549 8686 2580
rect 8862 2578 8898 2580
rect 8862 2549 8899 2578
rect 8101 2540 8136 2541
rect 8078 2535 8136 2540
rect 8078 2515 8081 2535
rect 8101 2521 8136 2535
rect 8156 2521 8165 2541
rect 8101 2513 8165 2521
rect 8127 2512 8165 2513
rect 8128 2511 8165 2512
rect 8231 2545 8267 2546
rect 8339 2545 8375 2546
rect 8231 2537 8375 2545
rect 8231 2517 8239 2537
rect 8259 2517 8347 2537
rect 8367 2517 8375 2537
rect 8231 2511 8375 2517
rect 8441 2541 8479 2549
rect 8547 2545 8583 2546
rect 8441 2521 8450 2541
rect 8470 2521 8479 2541
rect 8441 2512 8479 2521
rect 8498 2538 8583 2545
rect 8498 2518 8505 2538
rect 8526 2537 8583 2538
rect 8526 2518 8555 2537
rect 8498 2517 8555 2518
rect 8575 2517 8583 2537
rect 8441 2511 8478 2512
rect 8498 2511 8583 2517
rect 8649 2541 8687 2549
rect 8760 2545 8796 2546
rect 8649 2521 8658 2541
rect 8678 2521 8687 2541
rect 8649 2512 8687 2521
rect 8711 2537 8796 2545
rect 8711 2517 8768 2537
rect 8788 2517 8796 2537
rect 8649 2511 8686 2512
rect 8711 2511 8796 2517
rect 8862 2541 8900 2549
rect 8862 2521 8871 2541
rect 8891 2521 8900 2541
rect 8862 2512 8900 2521
rect 8940 2526 9012 2736
rect 9082 2770 10282 2800
rect 9082 2769 9526 2770
rect 9082 2767 9250 2769
rect 8940 2512 9023 2526
rect 8862 2511 8899 2512
rect 8285 2490 8321 2511
rect 8711 2490 8742 2511
rect 8940 2490 8957 2512
rect 8118 2486 8218 2490
rect 8118 2482 8180 2486
rect 8118 2456 8125 2482
rect 8151 2460 8180 2482
rect 8206 2460 8218 2486
rect 8151 2456 8218 2460
rect 8118 2453 8218 2456
rect 8286 2453 8321 2490
rect 8383 2487 8742 2490
rect 8383 2482 8605 2487
rect 8383 2458 8396 2482
rect 8420 2463 8605 2482
rect 8629 2463 8742 2487
rect 8420 2458 8742 2463
rect 8383 2454 8742 2458
rect 8809 2482 8957 2490
rect 8809 2462 8820 2482
rect 8840 2479 8957 2482
rect 9010 2479 9023 2512
rect 8840 2462 9023 2479
rect 8809 2455 9023 2462
rect 8809 2454 8850 2455
rect 8940 2454 9023 2455
rect 8285 2428 8321 2453
rect 8133 2401 8170 2402
rect 8229 2401 8266 2402
rect 8285 2401 8292 2428
rect 8033 2392 8171 2401
rect 2845 2294 3002 2307
rect 2845 2290 3006 2294
rect 1725 2144 1751 2249
rect 2845 2183 2886 2290
rect 2986 2183 3006 2290
rect 2845 2154 3006 2183
rect 6982 2171 7031 2380
rect 8033 2372 8142 2392
rect 8162 2372 8171 2392
rect 8033 2365 8171 2372
rect 8229 2398 8292 2401
rect 8313 2401 8321 2428
rect 8340 2401 8377 2402
rect 8313 2398 8377 2401
rect 8229 2392 8377 2398
rect 8229 2372 8238 2392
rect 8258 2372 8348 2392
rect 8368 2372 8377 2392
rect 8033 2363 8129 2365
rect 8229 2362 8377 2372
rect 8436 2392 8473 2402
rect 8548 2401 8585 2402
rect 8529 2399 8585 2401
rect 8436 2372 8444 2392
rect 8464 2372 8473 2392
rect 8285 2361 8321 2362
rect 8133 2230 8170 2231
rect 8436 2230 8473 2372
rect 8498 2392 8585 2399
rect 8498 2389 8556 2392
rect 8498 2369 8503 2389
rect 8524 2372 8556 2389
rect 8576 2372 8585 2392
rect 8524 2369 8585 2372
rect 8498 2362 8585 2369
rect 8644 2392 8681 2402
rect 8644 2372 8652 2392
rect 8672 2372 8681 2392
rect 8498 2361 8529 2362
rect 8644 2293 8681 2372
rect 8711 2401 8742 2454
rect 8948 2421 8962 2454
rect 9015 2421 9023 2454
rect 8948 2415 9023 2421
rect 8948 2410 9018 2415
rect 8761 2401 8798 2402
rect 8711 2392 8798 2401
rect 8711 2372 8769 2392
rect 8789 2372 8798 2392
rect 8711 2362 8798 2372
rect 8857 2392 8894 2402
rect 9082 2397 9109 2767
rect 9149 2537 9213 2549
rect 9489 2545 9526 2769
rect 9997 2750 10061 2752
rect 9993 2738 10061 2750
rect 9993 2705 10004 2738
rect 10044 2705 10061 2738
rect 9993 2695 10061 2705
rect 9754 2634 9865 2649
rect 9754 2632 9796 2634
rect 9754 2612 9761 2632
rect 9780 2612 9796 2632
rect 9754 2604 9796 2612
rect 9824 2632 9865 2634
rect 9824 2612 9838 2632
rect 9857 2612 9865 2632
rect 9824 2604 9865 2612
rect 9754 2598 9865 2604
rect 9697 2576 9946 2598
rect 9697 2545 9734 2576
rect 9910 2574 9946 2576
rect 9910 2545 9947 2574
rect 9149 2536 9184 2537
rect 9126 2531 9184 2536
rect 9126 2511 9129 2531
rect 9149 2517 9184 2531
rect 9204 2517 9213 2537
rect 9149 2509 9213 2517
rect 9175 2508 9213 2509
rect 9176 2507 9213 2508
rect 9279 2541 9315 2542
rect 9387 2541 9423 2542
rect 9279 2533 9423 2541
rect 9279 2513 9287 2533
rect 9307 2513 9395 2533
rect 9415 2513 9423 2533
rect 9279 2507 9423 2513
rect 9489 2537 9527 2545
rect 9595 2541 9631 2542
rect 9489 2517 9498 2537
rect 9518 2517 9527 2537
rect 9489 2508 9527 2517
rect 9546 2534 9631 2541
rect 9546 2514 9553 2534
rect 9574 2533 9631 2534
rect 9574 2514 9603 2533
rect 9546 2513 9603 2514
rect 9623 2513 9631 2533
rect 9489 2507 9526 2508
rect 9546 2507 9631 2513
rect 9697 2537 9735 2545
rect 9808 2541 9844 2542
rect 9697 2517 9706 2537
rect 9726 2517 9735 2537
rect 9697 2508 9735 2517
rect 9759 2533 9844 2541
rect 9759 2513 9816 2533
rect 9836 2513 9844 2533
rect 9697 2507 9734 2508
rect 9759 2507 9844 2513
rect 9910 2537 9948 2545
rect 9910 2517 9919 2537
rect 9939 2517 9948 2537
rect 9910 2508 9948 2517
rect 9997 2511 10061 2695
rect 10217 2569 10282 2770
rect 11259 2830 11324 3031
rect 11480 2905 11544 3089
rect 11593 3083 11631 3092
rect 11593 3063 11602 3083
rect 11622 3063 11631 3083
rect 11593 3055 11631 3063
rect 11697 3087 11782 3093
rect 11807 3092 11844 3093
rect 11697 3067 11705 3087
rect 11725 3067 11782 3087
rect 11697 3059 11782 3067
rect 11806 3083 11844 3092
rect 11806 3063 11815 3083
rect 11835 3063 11844 3083
rect 11697 3058 11733 3059
rect 11806 3055 11844 3063
rect 11910 3087 11995 3093
rect 12015 3092 12052 3093
rect 11910 3067 11918 3087
rect 11938 3086 11995 3087
rect 11938 3067 11967 3086
rect 11910 3066 11967 3067
rect 11988 3066 11995 3086
rect 11910 3059 11995 3066
rect 12014 3083 12052 3092
rect 12014 3063 12023 3083
rect 12043 3063 12052 3083
rect 11910 3058 11946 3059
rect 12014 3055 12052 3063
rect 12118 3087 12262 3093
rect 12118 3067 12126 3087
rect 12146 3067 12234 3087
rect 12254 3067 12262 3087
rect 12118 3059 12262 3067
rect 12118 3058 12154 3059
rect 12226 3058 12262 3059
rect 12328 3092 12365 3093
rect 12328 3091 12366 3092
rect 12328 3083 12392 3091
rect 12328 3063 12337 3083
rect 12357 3069 12392 3083
rect 12412 3069 12415 3089
rect 12357 3064 12415 3069
rect 12357 3063 12392 3064
rect 11594 3026 11631 3055
rect 11595 3024 11631 3026
rect 11807 3024 11844 3055
rect 11595 3002 11844 3024
rect 11676 2996 11787 3002
rect 11676 2988 11717 2996
rect 11676 2968 11684 2988
rect 11703 2968 11717 2988
rect 11676 2966 11717 2968
rect 11745 2988 11787 2996
rect 11745 2968 11761 2988
rect 11780 2968 11787 2988
rect 11745 2966 11787 2968
rect 11676 2951 11787 2966
rect 11480 2895 11548 2905
rect 11480 2862 11497 2895
rect 11537 2862 11548 2895
rect 11480 2850 11548 2862
rect 11480 2848 11544 2850
rect 12015 2831 12052 3055
rect 12328 3051 12392 3063
rect 12432 2833 12459 3203
rect 12647 3198 12684 3208
rect 12743 3228 12830 3238
rect 12743 3208 12752 3228
rect 12772 3208 12830 3228
rect 12743 3199 12830 3208
rect 12743 3198 12780 3199
rect 12523 3185 12593 3190
rect 12518 3179 12593 3185
rect 12518 3146 12526 3179
rect 12579 3146 12593 3179
rect 12799 3146 12830 3199
rect 12860 3228 12897 3307
rect 13012 3238 13043 3239
rect 12860 3208 12869 3228
rect 12889 3208 12897 3228
rect 12860 3198 12897 3208
rect 12956 3231 13043 3238
rect 12956 3228 13017 3231
rect 12956 3208 12965 3228
rect 12985 3211 13017 3228
rect 13038 3211 13043 3231
rect 12985 3208 13043 3211
rect 12956 3201 13043 3208
rect 13068 3228 13105 3370
rect 13371 3369 13408 3370
rect 13220 3238 13256 3239
rect 13068 3208 13077 3228
rect 13097 3208 13105 3228
rect 12956 3199 13012 3201
rect 12956 3198 12993 3199
rect 13068 3198 13105 3208
rect 13164 3228 13312 3238
rect 13412 3235 13508 3237
rect 13164 3208 13173 3228
rect 13193 3208 13283 3228
rect 13303 3208 13312 3228
rect 13164 3202 13312 3208
rect 13164 3199 13228 3202
rect 13164 3198 13201 3199
rect 13220 3172 13228 3199
rect 13249 3199 13312 3202
rect 13370 3228 13508 3235
rect 13370 3208 13379 3228
rect 13399 3208 13508 3228
rect 13370 3199 13508 3208
rect 13249 3172 13256 3199
rect 13275 3198 13312 3199
rect 13371 3198 13408 3199
rect 13220 3147 13256 3172
rect 12518 3145 12601 3146
rect 12691 3145 12732 3146
rect 12518 3138 12732 3145
rect 12518 3121 12701 3138
rect 12518 3088 12531 3121
rect 12584 3118 12701 3121
rect 12721 3118 12732 3138
rect 12584 3110 12732 3118
rect 12799 3142 13158 3146
rect 12799 3137 13121 3142
rect 12799 3113 12912 3137
rect 12936 3118 13121 3137
rect 13145 3118 13158 3142
rect 12936 3113 13158 3118
rect 12799 3110 13158 3113
rect 13220 3110 13255 3147
rect 13323 3144 13423 3147
rect 13323 3140 13390 3144
rect 13323 3114 13335 3140
rect 13361 3118 13390 3140
rect 13416 3118 13423 3144
rect 13361 3114 13423 3118
rect 13323 3110 13423 3114
rect 12584 3088 12601 3110
rect 12799 3089 12830 3110
rect 13220 3089 13256 3110
rect 12642 3088 12679 3089
rect 12518 3074 12601 3088
rect 12291 2831 12459 2833
rect 12015 2830 12459 2831
rect 11259 2800 12459 2830
rect 12529 2864 12601 3074
rect 12641 3079 12679 3088
rect 12641 3059 12650 3079
rect 12670 3059 12679 3079
rect 12641 3051 12679 3059
rect 12745 3083 12830 3089
rect 12855 3088 12892 3089
rect 12745 3063 12753 3083
rect 12773 3063 12830 3083
rect 12745 3055 12830 3063
rect 12854 3079 12892 3088
rect 12854 3059 12863 3079
rect 12883 3059 12892 3079
rect 12745 3054 12781 3055
rect 12854 3051 12892 3059
rect 12958 3083 13043 3089
rect 13063 3088 13100 3089
rect 12958 3063 12966 3083
rect 12986 3082 13043 3083
rect 12986 3063 13015 3082
rect 12958 3062 13015 3063
rect 13036 3062 13043 3082
rect 12958 3055 13043 3062
rect 13062 3079 13100 3088
rect 13062 3059 13071 3079
rect 13091 3059 13100 3079
rect 12958 3054 12994 3055
rect 13062 3051 13100 3059
rect 13166 3083 13310 3089
rect 13166 3063 13174 3083
rect 13194 3063 13282 3083
rect 13302 3063 13310 3083
rect 13166 3055 13310 3063
rect 13166 3054 13202 3055
rect 13274 3054 13310 3055
rect 13376 3088 13413 3089
rect 13376 3087 13414 3088
rect 13376 3079 13440 3087
rect 13376 3059 13385 3079
rect 13405 3065 13440 3079
rect 13460 3065 13463 3085
rect 13405 3060 13463 3065
rect 13405 3059 13440 3060
rect 12642 3022 12679 3051
rect 12643 3020 12679 3022
rect 12855 3020 12892 3051
rect 12643 2998 12892 3020
rect 12724 2992 12835 2998
rect 12724 2984 12765 2992
rect 12724 2964 12732 2984
rect 12751 2964 12765 2984
rect 12724 2962 12765 2964
rect 12793 2984 12835 2992
rect 12793 2964 12809 2984
rect 12828 2964 12835 2984
rect 12793 2962 12835 2964
rect 12724 2947 12835 2962
rect 12529 2825 12548 2864
rect 12593 2825 12601 2864
rect 12529 2808 12601 2825
rect 13063 2852 13100 3051
rect 13376 3047 13440 3059
rect 13063 2846 13104 2852
rect 13480 2848 13507 3199
rect 13339 2846 13507 2848
rect 13063 2820 13507 2846
rect 11259 2753 11324 2800
rect 11259 2735 11282 2753
rect 11300 2735 11324 2753
rect 12172 2780 12207 2782
rect 12172 2778 12276 2780
rect 13065 2778 13104 2820
rect 13339 2819 13507 2820
rect 12172 2771 13106 2778
rect 12172 2770 12223 2771
rect 12172 2750 12175 2770
rect 12200 2751 12223 2770
rect 12255 2751 13106 2771
rect 12200 2750 13106 2751
rect 12172 2743 13106 2750
rect 12445 2742 13106 2743
rect 11259 2714 11324 2735
rect 11536 2725 11576 2728
rect 11536 2721 12439 2725
rect 11536 2701 12413 2721
rect 12433 2701 12439 2721
rect 11536 2698 12439 2701
rect 11260 2654 11325 2674
rect 11260 2636 11284 2654
rect 11302 2636 11325 2654
rect 11260 2609 11325 2636
rect 11536 2609 11576 2698
rect 12020 2696 12436 2698
rect 12020 2695 12361 2696
rect 11677 2664 11787 2678
rect 11677 2661 11720 2664
rect 11677 2656 11681 2661
rect 11259 2574 11576 2609
rect 11599 2634 11681 2656
rect 11710 2634 11720 2661
rect 11748 2637 11755 2664
rect 11784 2656 11787 2664
rect 11784 2637 11849 2656
rect 11748 2634 11849 2637
rect 11599 2632 11849 2634
rect 10217 2551 10239 2569
rect 10257 2551 10282 2569
rect 10217 2532 10282 2551
rect 9910 2507 9947 2508
rect 9333 2486 9369 2507
rect 9759 2486 9790 2507
rect 9997 2502 10005 2511
rect 9994 2486 10005 2502
rect 9166 2482 9266 2486
rect 9166 2478 9228 2482
rect 9166 2452 9173 2478
rect 9199 2456 9228 2478
rect 9254 2456 9266 2482
rect 9199 2452 9266 2456
rect 9166 2449 9266 2452
rect 9334 2449 9369 2486
rect 9431 2483 9790 2486
rect 9431 2478 9653 2483
rect 9431 2454 9444 2478
rect 9468 2459 9653 2478
rect 9677 2459 9790 2483
rect 9468 2454 9790 2459
rect 9431 2450 9790 2454
rect 9857 2478 10005 2486
rect 9857 2458 9868 2478
rect 9888 2469 10005 2478
rect 10054 2502 10061 2511
rect 10054 2469 10062 2502
rect 11260 2498 11325 2574
rect 11599 2553 11636 2632
rect 11677 2619 11787 2632
rect 11751 2563 11782 2564
rect 11599 2533 11608 2553
rect 11628 2533 11636 2553
rect 11599 2523 11636 2533
rect 11695 2553 11782 2563
rect 11695 2533 11704 2553
rect 11724 2533 11782 2553
rect 11695 2524 11782 2533
rect 11695 2523 11732 2524
rect 9888 2458 10062 2469
rect 9857 2451 10062 2458
rect 9857 2450 9898 2451
rect 9333 2424 9369 2449
rect 9181 2397 9218 2398
rect 9277 2397 9314 2398
rect 9333 2397 9340 2424
rect 8857 2372 8865 2392
rect 8885 2372 8894 2392
rect 8711 2361 8742 2362
rect 8706 2293 8816 2306
rect 8857 2293 8894 2372
rect 9081 2388 9219 2397
rect 9081 2368 9190 2388
rect 9210 2368 9219 2388
rect 9081 2361 9219 2368
rect 9277 2394 9340 2397
rect 9361 2397 9369 2424
rect 9388 2397 9425 2398
rect 9361 2394 9425 2397
rect 9277 2388 9425 2394
rect 9277 2368 9286 2388
rect 9306 2368 9396 2388
rect 9416 2368 9425 2388
rect 9081 2359 9177 2361
rect 9277 2358 9425 2368
rect 9484 2388 9521 2398
rect 9596 2397 9633 2398
rect 9577 2395 9633 2397
rect 9484 2368 9492 2388
rect 9512 2368 9521 2388
rect 9333 2357 9369 2358
rect 8644 2291 8894 2293
rect 8644 2288 8745 2291
rect 8644 2269 8709 2288
rect 8706 2261 8709 2269
rect 8738 2261 8745 2288
rect 8773 2264 8783 2291
rect 8812 2269 8894 2291
rect 8812 2264 8816 2269
rect 8773 2261 8816 2264
rect 8706 2247 8816 2261
rect 8132 2229 8473 2230
rect 8057 2224 8473 2229
rect 9181 2226 9218 2227
rect 9484 2226 9521 2368
rect 9546 2388 9633 2395
rect 9546 2385 9604 2388
rect 9546 2365 9551 2385
rect 9572 2368 9604 2385
rect 9624 2368 9633 2388
rect 9572 2365 9633 2368
rect 9546 2358 9633 2365
rect 9692 2388 9729 2398
rect 9692 2368 9700 2388
rect 9720 2368 9729 2388
rect 9546 2357 9577 2358
rect 9692 2289 9729 2368
rect 9759 2397 9790 2450
rect 9994 2448 10062 2451
rect 9994 2406 10006 2448
rect 10055 2406 10062 2448
rect 9809 2397 9846 2398
rect 9759 2388 9846 2397
rect 9759 2368 9817 2388
rect 9837 2368 9846 2388
rect 9759 2358 9846 2368
rect 9905 2388 9942 2398
rect 9994 2393 10062 2406
rect 10217 2470 10282 2487
rect 10217 2452 10241 2470
rect 10259 2452 10282 2470
rect 11260 2480 11282 2498
rect 11300 2480 11325 2498
rect 11260 2459 11325 2480
rect 11473 2478 11538 2487
rect 9905 2368 9913 2388
rect 9933 2368 9942 2388
rect 9759 2357 9790 2358
rect 9754 2289 9864 2302
rect 9905 2289 9942 2368
rect 10217 2313 10282 2452
rect 11473 2441 11483 2478
rect 11523 2470 11538 2478
rect 11751 2471 11782 2524
rect 11812 2553 11849 2632
rect 11964 2563 11995 2564
rect 11812 2533 11821 2553
rect 11841 2533 11849 2553
rect 11812 2523 11849 2533
rect 11908 2556 11995 2563
rect 11908 2553 11969 2556
rect 11908 2533 11917 2553
rect 11937 2536 11969 2553
rect 11990 2536 11995 2556
rect 11937 2533 11995 2536
rect 11908 2526 11995 2533
rect 12020 2553 12057 2695
rect 12323 2694 12360 2695
rect 12172 2563 12208 2564
rect 12020 2533 12029 2553
rect 12049 2533 12057 2553
rect 11908 2524 11964 2526
rect 11908 2523 11945 2524
rect 12020 2523 12057 2533
rect 12116 2553 12264 2563
rect 12364 2560 12460 2562
rect 12116 2533 12125 2553
rect 12145 2533 12235 2553
rect 12255 2533 12264 2553
rect 12116 2527 12264 2533
rect 12116 2524 12180 2527
rect 12116 2523 12153 2524
rect 12172 2497 12180 2524
rect 12201 2524 12264 2527
rect 12322 2553 12460 2560
rect 12322 2533 12331 2553
rect 12351 2533 12460 2553
rect 12322 2524 12460 2533
rect 12201 2497 12208 2524
rect 12227 2523 12264 2524
rect 12323 2523 12360 2524
rect 12172 2472 12208 2497
rect 11643 2470 11684 2471
rect 11523 2463 11684 2470
rect 11523 2443 11653 2463
rect 11673 2443 11684 2463
rect 11523 2441 11684 2443
rect 11473 2435 11684 2441
rect 11751 2467 12110 2471
rect 11751 2462 12073 2467
rect 11751 2438 11864 2462
rect 11888 2443 12073 2462
rect 12097 2443 12110 2467
rect 11888 2438 12110 2443
rect 11751 2435 12110 2438
rect 12172 2435 12207 2472
rect 12275 2469 12375 2472
rect 12275 2465 12342 2469
rect 12275 2439 12287 2465
rect 12313 2443 12342 2465
rect 12368 2443 12375 2469
rect 12313 2439 12375 2443
rect 12275 2435 12375 2439
rect 11473 2422 11540 2435
rect 11265 2399 11321 2419
rect 11265 2381 11284 2399
rect 11302 2381 11321 2399
rect 11265 2346 11321 2381
rect 10217 2307 10239 2313
rect 9692 2287 9942 2289
rect 9692 2284 9793 2287
rect 9692 2265 9757 2284
rect 9754 2257 9757 2265
rect 9786 2257 9793 2284
rect 9821 2260 9831 2287
rect 9860 2265 9942 2287
rect 9971 2295 10239 2307
rect 10257 2295 10282 2313
rect 9971 2272 10282 2295
rect 9971 2271 10026 2272
rect 9860 2260 9864 2265
rect 9821 2257 9864 2260
rect 9754 2243 9864 2257
rect 9180 2225 9521 2226
rect 8057 2204 8060 2224
rect 8080 2204 8473 2224
rect 9105 2224 9521 2225
rect 9971 2224 10014 2271
rect 11227 2268 11321 2346
rect 11473 2401 11487 2422
rect 11523 2401 11540 2422
rect 11751 2414 11782 2435
rect 12172 2414 12208 2435
rect 11594 2413 11631 2414
rect 11473 2394 11540 2401
rect 11593 2404 11631 2413
rect 9105 2220 10014 2224
rect 1725 2130 1753 2144
rect 2849 2141 3006 2154
rect 6980 2169 7797 2171
rect 8230 2169 8319 2172
rect 6980 2160 8319 2169
rect 527 2095 1753 2130
rect 6980 2122 8242 2160
rect 8267 2125 8286 2160
rect 8311 2125 8319 2160
rect 8424 2171 8469 2204
rect 9105 2200 9108 2220
rect 9128 2200 10014 2220
rect 9482 2195 10014 2200
rect 10222 2214 10281 2236
rect 10222 2196 10241 2214
rect 10259 2196 10281 2214
rect 9270 2171 9369 2173
rect 8424 2161 9369 2171
rect 8424 2135 9292 2161
rect 8425 2134 9292 2135
rect 8267 2122 8319 2125
rect 6980 2114 8319 2122
rect 9270 2123 9292 2134
rect 9317 2126 9336 2161
rect 9361 2126 9369 2161
rect 9317 2123 9369 2126
rect 9270 2115 9369 2123
rect 9296 2114 9368 2115
rect 6980 2113 8318 2114
rect 6980 2111 7797 2113
rect 7571 2107 7797 2111
rect 527 2019 612 2095
rect 970 2093 1074 2095
rect 1305 2093 1346 2095
rect 10222 2019 10281 2196
rect 11227 2127 11320 2268
rect 11473 2242 11538 2394
rect 11593 2384 11602 2404
rect 11622 2384 11631 2404
rect 11593 2376 11631 2384
rect 11697 2408 11782 2414
rect 11807 2413 11844 2414
rect 11697 2388 11705 2408
rect 11725 2388 11782 2408
rect 11697 2380 11782 2388
rect 11806 2404 11844 2413
rect 11806 2384 11815 2404
rect 11835 2384 11844 2404
rect 11697 2379 11733 2380
rect 11806 2376 11844 2384
rect 11910 2408 11995 2414
rect 12015 2413 12052 2414
rect 11910 2388 11918 2408
rect 11938 2407 11995 2408
rect 11938 2388 11967 2407
rect 11910 2387 11967 2388
rect 11988 2387 11995 2407
rect 11910 2380 11995 2387
rect 12014 2404 12052 2413
rect 12014 2384 12023 2404
rect 12043 2384 12052 2404
rect 11910 2379 11946 2380
rect 12014 2376 12052 2384
rect 12118 2408 12262 2414
rect 12118 2388 12126 2408
rect 12146 2388 12234 2408
rect 12254 2388 12262 2408
rect 12118 2380 12262 2388
rect 12118 2379 12154 2380
rect 12226 2379 12262 2380
rect 12328 2413 12365 2414
rect 12328 2412 12366 2413
rect 12328 2404 12392 2412
rect 12328 2384 12337 2404
rect 12357 2390 12392 2404
rect 12412 2390 12415 2410
rect 12357 2385 12415 2390
rect 12357 2384 12392 2385
rect 11594 2347 11631 2376
rect 11595 2345 11631 2347
rect 11807 2345 11844 2376
rect 11595 2323 11844 2345
rect 11676 2317 11787 2323
rect 11676 2309 11717 2317
rect 11676 2289 11684 2309
rect 11703 2289 11717 2309
rect 11676 2287 11717 2289
rect 11745 2309 11787 2317
rect 11745 2289 11761 2309
rect 11780 2289 11787 2309
rect 11745 2287 11787 2289
rect 11676 2272 11787 2287
rect 12015 2277 12052 2376
rect 12328 2372 12392 2384
rect 12432 2333 12459 2524
rect 11678 2263 11782 2272
rect 11466 2232 11587 2242
rect 11466 2230 11535 2232
rect 11466 2189 11479 2230
rect 11516 2191 11535 2230
rect 11572 2191 11587 2232
rect 11516 2189 11587 2191
rect 11466 2171 11587 2189
rect 11678 2127 11782 2136
rect 12013 2127 12054 2277
rect 11227 2125 12054 2127
rect 11235 2124 12054 2125
rect 12433 2243 12458 2333
rect 13593 2301 13692 3858
rect 13798 2494 13897 5395
rect 14288 5378 14319 5399
rect 14709 5378 14745 5399
rect 14131 5377 14168 5378
rect 14130 5368 14168 5377
rect 14130 5348 14139 5368
rect 14159 5348 14168 5368
rect 14130 5340 14168 5348
rect 14234 5372 14319 5378
rect 14344 5377 14381 5378
rect 14234 5352 14242 5372
rect 14262 5352 14319 5372
rect 14234 5344 14319 5352
rect 14343 5368 14381 5377
rect 14343 5348 14352 5368
rect 14372 5348 14381 5368
rect 14234 5343 14270 5344
rect 14343 5340 14381 5348
rect 14447 5372 14532 5378
rect 14552 5377 14589 5378
rect 14447 5352 14455 5372
rect 14475 5371 14532 5372
rect 14475 5352 14504 5371
rect 14447 5351 14504 5352
rect 14525 5351 14532 5371
rect 14447 5344 14532 5351
rect 14551 5368 14589 5377
rect 14551 5348 14560 5368
rect 14580 5348 14589 5368
rect 14447 5343 14483 5344
rect 14551 5340 14589 5348
rect 14655 5372 14799 5378
rect 14655 5352 14663 5372
rect 14683 5352 14771 5372
rect 14791 5352 14799 5372
rect 14655 5344 14799 5352
rect 14655 5343 14691 5344
rect 14763 5343 14799 5344
rect 14865 5377 14902 5378
rect 14865 5376 14903 5377
rect 14865 5368 14929 5376
rect 14865 5348 14874 5368
rect 14894 5354 14929 5368
rect 14949 5354 14952 5374
rect 14894 5349 14952 5354
rect 14894 5348 14929 5349
rect 14131 5311 14168 5340
rect 14132 5309 14168 5311
rect 14344 5309 14381 5340
rect 14132 5287 14381 5309
rect 14213 5281 14324 5287
rect 14213 5273 14254 5281
rect 14213 5253 14221 5273
rect 14240 5253 14254 5273
rect 14213 5251 14254 5253
rect 14282 5273 14324 5281
rect 14282 5253 14298 5273
rect 14317 5253 14324 5273
rect 14282 5251 14324 5253
rect 14213 5236 14324 5251
rect 14552 5219 14589 5340
rect 14865 5336 14929 5348
rect 14670 5219 14699 5223
rect 14969 5221 14996 5488
rect 14828 5219 14996 5221
rect 14552 5193 14996 5219
rect 14511 4925 14556 4934
rect 14511 4887 14521 4925
rect 14546 4887 14556 4925
rect 14511 4876 14556 4887
rect 14514 4868 14556 4876
rect 14514 4163 14557 4868
rect 14670 4254 14699 5193
rect 14828 5192 14996 5193
rect 15400 5043 15484 5047
rect 15952 5043 16040 7894
rect 16579 7881 16634 7893
rect 16579 7847 16597 7881
rect 16626 7847 16634 7881
rect 16579 7821 16634 7847
rect 16186 7788 16354 7789
rect 16579 7788 16596 7821
rect 16186 7787 16596 7788
rect 16625 7787 16634 7821
rect 16186 7762 16634 7787
rect 16186 7760 16354 7762
rect 16186 7493 16213 7760
rect 16579 7756 16634 7762
rect 16253 7633 16317 7645
rect 16593 7641 16630 7756
rect 16858 7730 16969 7745
rect 16858 7728 16900 7730
rect 16858 7708 16865 7728
rect 16884 7708 16900 7728
rect 16858 7700 16900 7708
rect 16928 7728 16969 7730
rect 16928 7708 16942 7728
rect 16961 7708 16969 7728
rect 16928 7700 16969 7708
rect 16858 7694 16969 7700
rect 16801 7672 17050 7694
rect 16801 7641 16838 7672
rect 17014 7670 17050 7672
rect 17014 7641 17051 7670
rect 16253 7632 16288 7633
rect 16230 7627 16288 7632
rect 16230 7607 16233 7627
rect 16253 7613 16288 7627
rect 16308 7613 16317 7633
rect 16253 7605 16317 7613
rect 16279 7604 16317 7605
rect 16280 7603 16317 7604
rect 16383 7637 16419 7638
rect 16491 7637 16527 7638
rect 16383 7629 16527 7637
rect 16383 7609 16391 7629
rect 16411 7609 16499 7629
rect 16519 7609 16527 7629
rect 16383 7603 16527 7609
rect 16593 7633 16631 7641
rect 16699 7637 16735 7638
rect 16593 7613 16602 7633
rect 16622 7613 16631 7633
rect 16593 7604 16631 7613
rect 16650 7630 16735 7637
rect 16650 7610 16657 7630
rect 16678 7629 16735 7630
rect 16678 7610 16707 7629
rect 16650 7609 16707 7610
rect 16727 7609 16735 7629
rect 16593 7603 16630 7604
rect 16650 7603 16735 7609
rect 16801 7633 16839 7641
rect 16912 7637 16948 7638
rect 16801 7613 16810 7633
rect 16830 7613 16839 7633
rect 16801 7604 16839 7613
rect 16863 7629 16948 7637
rect 16863 7609 16920 7629
rect 16940 7609 16948 7629
rect 16801 7603 16838 7604
rect 16863 7603 16948 7609
rect 17014 7633 17052 7641
rect 17014 7613 17023 7633
rect 17043 7613 17052 7633
rect 17014 7604 17052 7613
rect 17014 7603 17051 7604
rect 16437 7582 16473 7603
rect 16863 7582 16894 7603
rect 17108 7586 17179 8239
rect 17694 8173 17737 8886
rect 18354 8797 18449 8817
rect 18354 8753 18374 8797
rect 18434 8753 18449 8797
rect 18354 8457 18449 8753
rect 18354 8416 18387 8457
rect 18423 8416 18449 8457
rect 18549 8496 18611 8967
rect 19891 8907 19928 8908
rect 20194 8907 20231 9049
rect 20256 9069 20343 9076
rect 20256 9066 20314 9069
rect 20256 9046 20261 9066
rect 20282 9049 20314 9066
rect 20334 9049 20343 9069
rect 20282 9046 20343 9049
rect 20256 9039 20343 9046
rect 20402 9069 20439 9079
rect 20402 9049 20410 9069
rect 20430 9049 20439 9069
rect 20256 9038 20287 9039
rect 20402 8970 20439 9049
rect 20469 9078 20500 9131
rect 20713 9124 20728 9132
rect 20768 9124 20778 9161
rect 22226 9160 22291 9299
rect 22566 9244 22603 9323
rect 22644 9310 22754 9323
rect 22718 9254 22749 9255
rect 22566 9224 22575 9244
rect 22595 9224 22603 9244
rect 20713 9115 20778 9124
rect 20926 9122 20991 9143
rect 22226 9142 22249 9160
rect 22267 9142 22291 9160
rect 22226 9125 22291 9142
rect 22446 9206 22514 9219
rect 22566 9214 22603 9224
rect 22662 9244 22749 9254
rect 22662 9224 22671 9244
rect 22691 9224 22749 9244
rect 22662 9215 22749 9224
rect 22662 9214 22699 9215
rect 22446 9164 22453 9206
rect 22502 9164 22514 9206
rect 22446 9161 22514 9164
rect 22718 9162 22749 9215
rect 22779 9244 22816 9323
rect 22931 9254 22962 9255
rect 22779 9224 22788 9244
rect 22808 9224 22816 9244
rect 22779 9214 22816 9224
rect 22875 9247 22962 9254
rect 22875 9244 22936 9247
rect 22875 9224 22884 9244
rect 22904 9227 22936 9244
rect 22957 9227 22962 9247
rect 22904 9224 22962 9227
rect 22875 9217 22962 9224
rect 22987 9244 23024 9386
rect 23290 9385 23327 9386
rect 24035 9383 24451 9388
rect 24035 9382 24376 9383
rect 23692 9351 23802 9365
rect 23692 9348 23735 9351
rect 23692 9343 23696 9348
rect 23614 9321 23696 9343
rect 23725 9321 23735 9348
rect 23763 9324 23770 9351
rect 23799 9343 23802 9351
rect 23799 9324 23864 9343
rect 23763 9321 23864 9324
rect 23614 9319 23864 9321
rect 23139 9254 23175 9255
rect 22987 9224 22996 9244
rect 23016 9224 23024 9244
rect 22875 9215 22931 9217
rect 22875 9214 22912 9215
rect 22987 9214 23024 9224
rect 23083 9244 23231 9254
rect 23331 9251 23427 9253
rect 23083 9224 23092 9244
rect 23112 9224 23202 9244
rect 23222 9224 23231 9244
rect 23083 9218 23231 9224
rect 23083 9215 23147 9218
rect 23083 9214 23120 9215
rect 23139 9188 23147 9215
rect 23168 9215 23231 9218
rect 23289 9244 23427 9251
rect 23289 9224 23298 9244
rect 23318 9224 23427 9244
rect 23289 9215 23427 9224
rect 23614 9240 23651 9319
rect 23692 9306 23802 9319
rect 23766 9250 23797 9251
rect 23614 9220 23623 9240
rect 23643 9220 23651 9240
rect 23168 9188 23175 9215
rect 23194 9214 23231 9215
rect 23290 9214 23327 9215
rect 23139 9163 23175 9188
rect 22610 9161 22651 9162
rect 22446 9154 22651 9161
rect 22446 9143 22620 9154
rect 20926 9104 20951 9122
rect 20969 9104 20991 9122
rect 22446 9110 22454 9143
rect 20519 9078 20556 9079
rect 20469 9069 20556 9078
rect 20469 9049 20527 9069
rect 20547 9049 20556 9069
rect 20469 9039 20556 9049
rect 20615 9069 20652 9079
rect 20615 9049 20623 9069
rect 20643 9049 20652 9069
rect 20469 9038 20500 9039
rect 20464 8970 20574 8983
rect 20615 8970 20652 9049
rect 20926 9028 20991 9104
rect 22447 9101 22454 9110
rect 22503 9134 22620 9143
rect 22640 9134 22651 9154
rect 22503 9126 22651 9134
rect 22718 9158 23077 9162
rect 22718 9153 23040 9158
rect 22718 9129 22831 9153
rect 22855 9134 23040 9153
rect 23064 9134 23077 9158
rect 22855 9129 23077 9134
rect 22718 9126 23077 9129
rect 23139 9126 23174 9163
rect 23242 9160 23342 9163
rect 23242 9156 23309 9160
rect 23242 9130 23254 9156
rect 23280 9134 23309 9156
rect 23335 9134 23342 9160
rect 23280 9130 23342 9134
rect 23242 9126 23342 9130
rect 22503 9110 22514 9126
rect 22503 9101 22511 9110
rect 22718 9105 22749 9126
rect 23139 9105 23175 9126
rect 22561 9104 22598 9105
rect 22226 9061 22291 9080
rect 22226 9043 22251 9061
rect 22269 9043 22291 9061
rect 20402 8968 20652 8970
rect 20402 8965 20503 8968
rect 20402 8946 20467 8965
rect 20464 8938 20467 8946
rect 20496 8938 20503 8965
rect 20531 8941 20541 8968
rect 20570 8946 20652 8968
rect 20675 8993 20992 9028
rect 20570 8941 20574 8946
rect 20531 8938 20574 8941
rect 20464 8924 20574 8938
rect 19890 8906 20231 8907
rect 19815 8904 20231 8906
rect 20675 8904 20715 8993
rect 20926 8966 20991 8993
rect 20926 8948 20949 8966
rect 20967 8948 20991 8966
rect 20926 8928 20991 8948
rect 19812 8901 20715 8904
rect 19812 8881 19818 8901
rect 19838 8881 20715 8901
rect 19812 8877 20715 8881
rect 20675 8874 20715 8877
rect 20927 8867 20992 8888
rect 19145 8859 19806 8860
rect 19145 8852 20079 8859
rect 19145 8851 20051 8852
rect 19145 8831 19996 8851
rect 20028 8832 20051 8851
rect 20076 8832 20079 8852
rect 20028 8831 20079 8832
rect 19145 8824 20079 8831
rect 18744 8782 18912 8783
rect 19147 8782 19186 8824
rect 19975 8822 20079 8824
rect 20044 8820 20079 8822
rect 20927 8849 20951 8867
rect 20969 8849 20992 8867
rect 20927 8802 20992 8849
rect 18744 8756 19188 8782
rect 18744 8754 18912 8756
rect 18549 8477 18613 8496
rect 18549 8438 18566 8477
rect 18600 8438 18613 8477
rect 18549 8419 18613 8438
rect 18354 8390 18449 8416
rect 18744 8403 18771 8754
rect 19147 8750 19188 8756
rect 18811 8543 18875 8555
rect 19151 8551 19188 8750
rect 19650 8777 19722 8794
rect 19650 8738 19658 8777
rect 19703 8738 19722 8777
rect 19416 8640 19527 8655
rect 19416 8638 19458 8640
rect 19416 8618 19423 8638
rect 19442 8618 19458 8638
rect 19416 8610 19458 8618
rect 19486 8638 19527 8640
rect 19486 8618 19500 8638
rect 19519 8618 19527 8638
rect 19486 8610 19527 8618
rect 19416 8604 19527 8610
rect 19359 8582 19608 8604
rect 19359 8551 19396 8582
rect 19572 8580 19608 8582
rect 19572 8551 19609 8580
rect 18811 8542 18846 8543
rect 18788 8537 18846 8542
rect 18788 8517 18791 8537
rect 18811 8523 18846 8537
rect 18866 8523 18875 8543
rect 18811 8515 18875 8523
rect 18837 8514 18875 8515
rect 18838 8513 18875 8514
rect 18941 8547 18977 8548
rect 19049 8547 19085 8548
rect 18941 8539 19085 8547
rect 18941 8519 18949 8539
rect 18969 8519 19057 8539
rect 19077 8519 19085 8539
rect 18941 8513 19085 8519
rect 19151 8543 19189 8551
rect 19257 8547 19293 8548
rect 19151 8523 19160 8543
rect 19180 8523 19189 8543
rect 19151 8514 19189 8523
rect 19208 8540 19293 8547
rect 19208 8520 19215 8540
rect 19236 8539 19293 8540
rect 19236 8520 19265 8539
rect 19208 8519 19265 8520
rect 19285 8519 19293 8539
rect 19151 8513 19188 8514
rect 19208 8513 19293 8519
rect 19359 8543 19397 8551
rect 19470 8547 19506 8548
rect 19359 8523 19368 8543
rect 19388 8523 19397 8543
rect 19359 8514 19397 8523
rect 19421 8539 19506 8547
rect 19421 8519 19478 8539
rect 19498 8519 19506 8539
rect 19359 8513 19396 8514
rect 19421 8513 19506 8519
rect 19572 8543 19610 8551
rect 19572 8523 19581 8543
rect 19601 8523 19610 8543
rect 19572 8514 19610 8523
rect 19650 8528 19722 8738
rect 19792 8772 20992 8802
rect 19792 8771 20236 8772
rect 19792 8769 19960 8771
rect 19650 8514 19733 8528
rect 19572 8513 19609 8514
rect 18995 8492 19031 8513
rect 19421 8492 19452 8513
rect 19650 8492 19667 8514
rect 18828 8488 18928 8492
rect 18828 8484 18890 8488
rect 18828 8458 18835 8484
rect 18861 8462 18890 8484
rect 18916 8462 18928 8488
rect 18861 8458 18928 8462
rect 18828 8455 18928 8458
rect 18996 8455 19031 8492
rect 19093 8489 19452 8492
rect 19093 8484 19315 8489
rect 19093 8460 19106 8484
rect 19130 8465 19315 8484
rect 19339 8465 19452 8489
rect 19130 8460 19452 8465
rect 19093 8456 19452 8460
rect 19519 8484 19667 8492
rect 19519 8464 19530 8484
rect 19550 8481 19667 8484
rect 19720 8481 19733 8514
rect 19550 8464 19733 8481
rect 19519 8457 19733 8464
rect 19519 8456 19560 8457
rect 19650 8456 19733 8457
rect 18995 8430 19031 8455
rect 18843 8403 18880 8404
rect 18939 8403 18976 8404
rect 18995 8403 19002 8430
rect 18743 8394 18881 8403
rect 18743 8374 18852 8394
rect 18872 8374 18881 8394
rect 18743 8367 18881 8374
rect 18939 8400 19002 8403
rect 19023 8403 19031 8430
rect 19050 8403 19087 8404
rect 19023 8400 19087 8403
rect 18939 8394 19087 8400
rect 18939 8374 18948 8394
rect 18968 8374 19058 8394
rect 19078 8374 19087 8394
rect 18743 8365 18839 8367
rect 18939 8364 19087 8374
rect 19146 8394 19183 8404
rect 19258 8403 19295 8404
rect 19239 8401 19295 8403
rect 19146 8374 19154 8394
rect 19174 8374 19183 8394
rect 18995 8363 19031 8364
rect 18843 8232 18880 8233
rect 19146 8232 19183 8374
rect 19208 8394 19295 8401
rect 19208 8391 19266 8394
rect 19208 8371 19213 8391
rect 19234 8374 19266 8391
rect 19286 8374 19295 8394
rect 19234 8371 19295 8374
rect 19208 8364 19295 8371
rect 19354 8394 19391 8404
rect 19354 8374 19362 8394
rect 19382 8374 19391 8394
rect 19208 8363 19239 8364
rect 19354 8295 19391 8374
rect 19421 8403 19452 8456
rect 19658 8423 19672 8456
rect 19725 8423 19733 8456
rect 19658 8417 19733 8423
rect 19658 8412 19728 8417
rect 19471 8403 19508 8404
rect 19421 8394 19508 8403
rect 19421 8374 19479 8394
rect 19499 8374 19508 8394
rect 19421 8364 19508 8374
rect 19567 8394 19604 8404
rect 19792 8399 19819 8769
rect 19859 8539 19923 8551
rect 20199 8547 20236 8771
rect 20707 8752 20771 8754
rect 20703 8740 20771 8752
rect 20703 8707 20714 8740
rect 20754 8707 20771 8740
rect 20703 8697 20771 8707
rect 20464 8636 20575 8651
rect 20464 8634 20506 8636
rect 20464 8614 20471 8634
rect 20490 8614 20506 8634
rect 20464 8606 20506 8614
rect 20534 8634 20575 8636
rect 20534 8614 20548 8634
rect 20567 8614 20575 8634
rect 20534 8606 20575 8614
rect 20464 8600 20575 8606
rect 20407 8578 20656 8600
rect 20407 8547 20444 8578
rect 20620 8576 20656 8578
rect 20620 8547 20657 8576
rect 19859 8538 19894 8539
rect 19836 8533 19894 8538
rect 19836 8513 19839 8533
rect 19859 8519 19894 8533
rect 19914 8519 19923 8539
rect 19859 8511 19923 8519
rect 19885 8510 19923 8511
rect 19886 8509 19923 8510
rect 19989 8543 20025 8544
rect 20097 8543 20133 8544
rect 19989 8535 20133 8543
rect 19989 8515 19997 8535
rect 20017 8515 20105 8535
rect 20125 8515 20133 8535
rect 19989 8509 20133 8515
rect 20199 8539 20237 8547
rect 20305 8543 20341 8544
rect 20199 8519 20208 8539
rect 20228 8519 20237 8539
rect 20199 8510 20237 8519
rect 20256 8536 20341 8543
rect 20256 8516 20263 8536
rect 20284 8535 20341 8536
rect 20284 8516 20313 8535
rect 20256 8515 20313 8516
rect 20333 8515 20341 8535
rect 20199 8509 20236 8510
rect 20256 8509 20341 8515
rect 20407 8539 20445 8547
rect 20518 8543 20554 8544
rect 20407 8519 20416 8539
rect 20436 8519 20445 8539
rect 20407 8510 20445 8519
rect 20469 8535 20554 8543
rect 20469 8515 20526 8535
rect 20546 8515 20554 8535
rect 20407 8509 20444 8510
rect 20469 8509 20554 8515
rect 20620 8539 20658 8547
rect 20620 8519 20629 8539
rect 20649 8519 20658 8539
rect 20620 8510 20658 8519
rect 20707 8513 20771 8697
rect 20927 8571 20992 8772
rect 22226 8842 22291 9043
rect 22447 8917 22511 9101
rect 22560 9095 22598 9104
rect 22560 9075 22569 9095
rect 22589 9075 22598 9095
rect 22560 9067 22598 9075
rect 22664 9099 22749 9105
rect 22774 9104 22811 9105
rect 22664 9079 22672 9099
rect 22692 9079 22749 9099
rect 22664 9071 22749 9079
rect 22773 9095 22811 9104
rect 22773 9075 22782 9095
rect 22802 9075 22811 9095
rect 22664 9070 22700 9071
rect 22773 9067 22811 9075
rect 22877 9099 22962 9105
rect 22982 9104 23019 9105
rect 22877 9079 22885 9099
rect 22905 9098 22962 9099
rect 22905 9079 22934 9098
rect 22877 9078 22934 9079
rect 22955 9078 22962 9098
rect 22877 9071 22962 9078
rect 22981 9095 23019 9104
rect 22981 9075 22990 9095
rect 23010 9075 23019 9095
rect 22877 9070 22913 9071
rect 22981 9067 23019 9075
rect 23085 9099 23229 9105
rect 23085 9079 23093 9099
rect 23113 9079 23201 9099
rect 23221 9079 23229 9099
rect 23085 9071 23229 9079
rect 23085 9070 23121 9071
rect 23193 9070 23229 9071
rect 23295 9104 23332 9105
rect 23295 9103 23333 9104
rect 23295 9095 23359 9103
rect 23295 9075 23304 9095
rect 23324 9081 23359 9095
rect 23379 9081 23382 9101
rect 23324 9076 23382 9081
rect 23324 9075 23359 9076
rect 22561 9038 22598 9067
rect 22562 9036 22598 9038
rect 22774 9036 22811 9067
rect 22562 9014 22811 9036
rect 22643 9008 22754 9014
rect 22643 9000 22684 9008
rect 22643 8980 22651 9000
rect 22670 8980 22684 9000
rect 22643 8978 22684 8980
rect 22712 9000 22754 9008
rect 22712 8980 22728 9000
rect 22747 8980 22754 9000
rect 22712 8978 22754 8980
rect 22643 8963 22754 8978
rect 22447 8907 22515 8917
rect 22447 8874 22464 8907
rect 22504 8874 22515 8907
rect 22447 8862 22515 8874
rect 22447 8860 22511 8862
rect 22982 8843 23019 9067
rect 23295 9063 23359 9075
rect 23399 8845 23426 9215
rect 23614 9210 23651 9220
rect 23710 9240 23797 9250
rect 23710 9220 23719 9240
rect 23739 9220 23797 9240
rect 23710 9211 23797 9220
rect 23710 9210 23747 9211
rect 23490 9197 23560 9202
rect 23485 9191 23560 9197
rect 23485 9158 23493 9191
rect 23546 9158 23560 9191
rect 23766 9158 23797 9211
rect 23827 9240 23864 9319
rect 23979 9250 24010 9251
rect 23827 9220 23836 9240
rect 23856 9220 23864 9240
rect 23827 9210 23864 9220
rect 23923 9243 24010 9250
rect 23923 9240 23984 9243
rect 23923 9220 23932 9240
rect 23952 9223 23984 9240
rect 24005 9223 24010 9243
rect 23952 9220 24010 9223
rect 23923 9213 24010 9220
rect 24035 9240 24072 9382
rect 24338 9381 24375 9382
rect 24187 9250 24223 9251
rect 24035 9220 24044 9240
rect 24064 9220 24072 9240
rect 23923 9211 23979 9213
rect 23923 9210 23960 9211
rect 24035 9210 24072 9220
rect 24131 9240 24279 9250
rect 24379 9247 24475 9249
rect 24131 9220 24140 9240
rect 24160 9220 24250 9240
rect 24270 9220 24279 9240
rect 24131 9214 24279 9220
rect 24131 9211 24195 9214
rect 24131 9210 24168 9211
rect 24187 9184 24195 9211
rect 24216 9211 24279 9214
rect 24337 9240 24475 9247
rect 24337 9220 24346 9240
rect 24366 9220 24475 9240
rect 24337 9211 24475 9220
rect 24216 9184 24223 9211
rect 24242 9210 24279 9211
rect 24338 9210 24375 9211
rect 24187 9159 24223 9184
rect 23485 9157 23568 9158
rect 23658 9157 23699 9158
rect 23485 9150 23699 9157
rect 23485 9133 23668 9150
rect 23485 9100 23498 9133
rect 23551 9130 23668 9133
rect 23688 9130 23699 9150
rect 23551 9122 23699 9130
rect 23766 9154 24125 9158
rect 23766 9149 24088 9154
rect 23766 9125 23879 9149
rect 23903 9130 24088 9149
rect 24112 9130 24125 9154
rect 23903 9125 24125 9130
rect 23766 9122 24125 9125
rect 24187 9122 24222 9159
rect 24290 9156 24390 9159
rect 24290 9152 24357 9156
rect 24290 9126 24302 9152
rect 24328 9130 24357 9152
rect 24383 9130 24390 9156
rect 24328 9126 24390 9130
rect 24290 9122 24390 9126
rect 23551 9100 23568 9122
rect 23766 9101 23797 9122
rect 24187 9101 24223 9122
rect 23609 9100 23646 9101
rect 23485 9086 23568 9100
rect 23258 8843 23426 8845
rect 22982 8842 23426 8843
rect 22226 8812 23426 8842
rect 23496 8876 23568 9086
rect 23608 9091 23646 9100
rect 23608 9071 23617 9091
rect 23637 9071 23646 9091
rect 23608 9063 23646 9071
rect 23712 9095 23797 9101
rect 23822 9100 23859 9101
rect 23712 9075 23720 9095
rect 23740 9075 23797 9095
rect 23712 9067 23797 9075
rect 23821 9091 23859 9100
rect 23821 9071 23830 9091
rect 23850 9071 23859 9091
rect 23712 9066 23748 9067
rect 23821 9063 23859 9071
rect 23925 9095 24010 9101
rect 24030 9100 24067 9101
rect 23925 9075 23933 9095
rect 23953 9094 24010 9095
rect 23953 9075 23982 9094
rect 23925 9074 23982 9075
rect 24003 9074 24010 9094
rect 23925 9067 24010 9074
rect 24029 9091 24067 9100
rect 24029 9071 24038 9091
rect 24058 9071 24067 9091
rect 23925 9066 23961 9067
rect 24029 9063 24067 9071
rect 24133 9095 24277 9101
rect 24133 9075 24141 9095
rect 24161 9075 24249 9095
rect 24269 9075 24277 9095
rect 24133 9067 24277 9075
rect 24133 9066 24169 9067
rect 24241 9066 24277 9067
rect 24343 9100 24380 9101
rect 24343 9099 24381 9100
rect 24343 9091 24407 9099
rect 24343 9071 24352 9091
rect 24372 9077 24407 9091
rect 24427 9077 24430 9097
rect 24372 9072 24430 9077
rect 24372 9071 24407 9072
rect 23609 9034 23646 9063
rect 23610 9032 23646 9034
rect 23822 9032 23859 9063
rect 23610 9010 23859 9032
rect 23691 9004 23802 9010
rect 23691 8996 23732 9004
rect 23691 8976 23699 8996
rect 23718 8976 23732 8996
rect 23691 8974 23732 8976
rect 23760 8996 23802 9004
rect 23760 8976 23776 8996
rect 23795 8976 23802 8996
rect 23760 8974 23802 8976
rect 23691 8959 23802 8974
rect 23496 8837 23515 8876
rect 23560 8837 23568 8876
rect 23496 8820 23568 8837
rect 24030 8864 24067 9063
rect 24343 9059 24407 9071
rect 24030 8858 24071 8864
rect 24447 8860 24474 9211
rect 24306 8858 24474 8860
rect 24030 8832 24474 8858
rect 22226 8765 22291 8812
rect 22226 8747 22249 8765
rect 22267 8747 22291 8765
rect 23139 8792 23174 8794
rect 23139 8790 23243 8792
rect 24032 8790 24071 8832
rect 24306 8831 24474 8832
rect 23139 8783 24073 8790
rect 23139 8782 23190 8783
rect 23139 8762 23142 8782
rect 23167 8763 23190 8782
rect 23222 8763 24073 8783
rect 23167 8762 24073 8763
rect 23139 8755 24073 8762
rect 23412 8754 24073 8755
rect 22226 8726 22291 8747
rect 22503 8737 22543 8740
rect 22503 8733 23406 8737
rect 22503 8713 23380 8733
rect 23400 8713 23406 8733
rect 22503 8710 23406 8713
rect 22227 8666 22292 8686
rect 22227 8648 22251 8666
rect 22269 8648 22292 8666
rect 22227 8621 22292 8648
rect 22503 8621 22543 8710
rect 22987 8708 23403 8710
rect 22987 8707 23328 8708
rect 22644 8676 22754 8690
rect 22644 8673 22687 8676
rect 22644 8668 22648 8673
rect 22226 8586 22543 8621
rect 22566 8646 22648 8668
rect 22677 8646 22687 8673
rect 22715 8649 22722 8676
rect 22751 8668 22754 8676
rect 22751 8649 22816 8668
rect 22715 8646 22816 8649
rect 22566 8644 22816 8646
rect 20927 8553 20949 8571
rect 20967 8553 20992 8571
rect 20927 8534 20992 8553
rect 20620 8509 20657 8510
rect 20043 8488 20079 8509
rect 20469 8488 20500 8509
rect 20707 8504 20715 8513
rect 20704 8488 20715 8504
rect 19876 8484 19976 8488
rect 19876 8480 19938 8484
rect 19876 8454 19883 8480
rect 19909 8458 19938 8480
rect 19964 8458 19976 8484
rect 19909 8454 19976 8458
rect 19876 8451 19976 8454
rect 20044 8451 20079 8488
rect 20141 8485 20500 8488
rect 20141 8480 20363 8485
rect 20141 8456 20154 8480
rect 20178 8461 20363 8480
rect 20387 8461 20500 8485
rect 20178 8456 20500 8461
rect 20141 8452 20500 8456
rect 20567 8480 20715 8488
rect 20567 8460 20578 8480
rect 20598 8471 20715 8480
rect 20764 8504 20771 8513
rect 22227 8510 22292 8586
rect 22566 8565 22603 8644
rect 22644 8631 22754 8644
rect 22718 8575 22749 8576
rect 22566 8545 22575 8565
rect 22595 8545 22603 8565
rect 22566 8535 22603 8545
rect 22662 8565 22749 8575
rect 22662 8545 22671 8565
rect 22691 8545 22749 8565
rect 22662 8536 22749 8545
rect 22662 8535 22699 8536
rect 20764 8471 20772 8504
rect 22227 8492 22249 8510
rect 22267 8492 22292 8510
rect 20598 8460 20772 8471
rect 20567 8453 20772 8460
rect 20567 8452 20608 8453
rect 20043 8426 20079 8451
rect 19891 8399 19928 8400
rect 19987 8399 20024 8400
rect 20043 8399 20050 8426
rect 19567 8374 19575 8394
rect 19595 8374 19604 8394
rect 19421 8363 19452 8364
rect 19416 8295 19526 8308
rect 19567 8295 19604 8374
rect 19791 8390 19929 8399
rect 19791 8370 19900 8390
rect 19920 8370 19929 8390
rect 19791 8363 19929 8370
rect 19987 8396 20050 8399
rect 20071 8399 20079 8426
rect 20098 8399 20135 8400
rect 20071 8396 20135 8399
rect 19987 8390 20135 8396
rect 19987 8370 19996 8390
rect 20016 8370 20106 8390
rect 20126 8370 20135 8390
rect 19791 8361 19887 8363
rect 19987 8360 20135 8370
rect 20194 8390 20231 8400
rect 20306 8399 20343 8400
rect 20287 8397 20343 8399
rect 20194 8370 20202 8390
rect 20222 8370 20231 8390
rect 20043 8359 20079 8360
rect 19354 8293 19604 8295
rect 19354 8290 19455 8293
rect 19354 8271 19419 8290
rect 19416 8263 19419 8271
rect 19448 8263 19455 8290
rect 19483 8266 19493 8293
rect 19522 8271 19604 8293
rect 19522 8266 19526 8271
rect 19483 8263 19526 8266
rect 19416 8249 19526 8263
rect 18842 8231 19183 8232
rect 18767 8226 19183 8231
rect 19891 8228 19928 8229
rect 20194 8228 20231 8370
rect 20256 8390 20343 8397
rect 20256 8387 20314 8390
rect 20256 8367 20261 8387
rect 20282 8370 20314 8387
rect 20334 8370 20343 8390
rect 20282 8367 20343 8370
rect 20256 8360 20343 8367
rect 20402 8390 20439 8400
rect 20402 8370 20410 8390
rect 20430 8370 20439 8390
rect 20256 8359 20287 8360
rect 20402 8291 20439 8370
rect 20469 8399 20500 8452
rect 20704 8450 20772 8453
rect 20704 8408 20716 8450
rect 20765 8408 20772 8450
rect 20519 8399 20556 8400
rect 20469 8390 20556 8399
rect 20469 8370 20527 8390
rect 20547 8370 20556 8390
rect 20469 8360 20556 8370
rect 20615 8390 20652 8400
rect 20704 8395 20772 8408
rect 20927 8472 20992 8489
rect 20927 8454 20951 8472
rect 20969 8454 20992 8472
rect 22227 8471 22292 8492
rect 22440 8490 22505 8499
rect 20615 8370 20623 8390
rect 20643 8370 20652 8390
rect 20469 8359 20500 8360
rect 20464 8291 20574 8304
rect 20615 8291 20652 8370
rect 20927 8315 20992 8454
rect 22440 8453 22450 8490
rect 22490 8482 22505 8490
rect 22718 8483 22749 8536
rect 22779 8565 22816 8644
rect 22931 8575 22962 8576
rect 22779 8545 22788 8565
rect 22808 8545 22816 8565
rect 22779 8535 22816 8545
rect 22875 8568 22962 8575
rect 22875 8565 22936 8568
rect 22875 8545 22884 8565
rect 22904 8548 22936 8565
rect 22957 8548 22962 8568
rect 22904 8545 22962 8548
rect 22875 8538 22962 8545
rect 22987 8565 23024 8707
rect 23290 8706 23327 8707
rect 23139 8575 23175 8576
rect 22987 8545 22996 8565
rect 23016 8545 23024 8565
rect 22875 8536 22931 8538
rect 22875 8535 22912 8536
rect 22987 8535 23024 8545
rect 23083 8565 23231 8575
rect 23331 8572 23427 8574
rect 23083 8545 23092 8565
rect 23112 8545 23202 8565
rect 23222 8545 23231 8565
rect 23083 8539 23231 8545
rect 23083 8536 23147 8539
rect 23083 8535 23120 8536
rect 23139 8509 23147 8536
rect 23168 8536 23231 8539
rect 23289 8565 23427 8572
rect 23289 8545 23298 8565
rect 23318 8545 23427 8565
rect 23289 8536 23427 8545
rect 23168 8509 23175 8536
rect 23194 8535 23231 8536
rect 23290 8535 23327 8536
rect 23139 8484 23175 8509
rect 22610 8482 22651 8483
rect 22490 8475 22651 8482
rect 22490 8455 22620 8475
rect 22640 8455 22651 8475
rect 22490 8453 22651 8455
rect 22440 8447 22651 8453
rect 22718 8479 23077 8483
rect 22718 8474 23040 8479
rect 22718 8450 22831 8474
rect 22855 8455 23040 8474
rect 23064 8455 23077 8479
rect 22855 8450 23077 8455
rect 22718 8447 23077 8450
rect 23139 8447 23174 8484
rect 23242 8481 23342 8484
rect 23242 8477 23309 8481
rect 23242 8451 23254 8477
rect 23280 8455 23309 8477
rect 23335 8455 23342 8481
rect 23280 8451 23342 8455
rect 23242 8447 23342 8451
rect 22440 8434 22507 8447
rect 20927 8309 20949 8315
rect 20402 8289 20652 8291
rect 20402 8286 20503 8289
rect 20402 8267 20467 8286
rect 20464 8259 20467 8267
rect 20496 8259 20503 8286
rect 20531 8262 20541 8289
rect 20570 8267 20652 8289
rect 20681 8297 20949 8309
rect 20967 8297 20992 8315
rect 20681 8274 20992 8297
rect 22232 8411 22288 8431
rect 22232 8393 22251 8411
rect 22269 8393 22288 8411
rect 22232 8280 22288 8393
rect 22440 8413 22454 8434
rect 22490 8413 22507 8434
rect 22718 8426 22749 8447
rect 23139 8426 23175 8447
rect 22561 8425 22598 8426
rect 22440 8406 22507 8413
rect 22560 8416 22598 8425
rect 20681 8273 20736 8274
rect 20570 8262 20574 8267
rect 20531 8259 20574 8262
rect 20464 8245 20574 8259
rect 19890 8227 20231 8228
rect 18767 8206 18770 8226
rect 18790 8206 19183 8226
rect 19815 8226 20231 8227
rect 20681 8226 20724 8273
rect 19815 8222 20724 8226
rect 17690 8171 18401 8173
rect 18940 8171 19029 8174
rect 17690 8162 19029 8171
rect 17690 8124 18952 8162
rect 18977 8127 18996 8162
rect 19021 8127 19029 8162
rect 19134 8173 19179 8206
rect 19815 8202 19818 8222
rect 19838 8202 20724 8222
rect 20192 8197 20724 8202
rect 20932 8216 20991 8238
rect 20932 8198 20951 8216
rect 20969 8198 20991 8216
rect 19980 8173 20079 8175
rect 19134 8163 20079 8173
rect 19134 8137 20002 8163
rect 19135 8136 20002 8137
rect 18977 8124 19029 8127
rect 17690 8116 19029 8124
rect 19980 8125 20002 8136
rect 20027 8128 20046 8163
rect 20071 8128 20079 8163
rect 20027 8125 20079 8128
rect 19980 8117 20079 8125
rect 20932 8124 20991 8198
rect 22232 8173 22287 8280
rect 22440 8254 22505 8406
rect 22560 8396 22569 8416
rect 22589 8396 22598 8416
rect 22560 8388 22598 8396
rect 22664 8420 22749 8426
rect 22774 8425 22811 8426
rect 22664 8400 22672 8420
rect 22692 8400 22749 8420
rect 22664 8392 22749 8400
rect 22773 8416 22811 8425
rect 22773 8396 22782 8416
rect 22802 8396 22811 8416
rect 22664 8391 22700 8392
rect 22773 8388 22811 8396
rect 22877 8420 22962 8426
rect 22982 8425 23019 8426
rect 22877 8400 22885 8420
rect 22905 8419 22962 8420
rect 22905 8400 22934 8419
rect 22877 8399 22934 8400
rect 22955 8399 22962 8419
rect 22877 8392 22962 8399
rect 22981 8416 23019 8425
rect 22981 8396 22990 8416
rect 23010 8396 23019 8416
rect 22877 8391 22913 8392
rect 22981 8388 23019 8396
rect 23085 8420 23229 8426
rect 23085 8400 23093 8420
rect 23113 8400 23201 8420
rect 23221 8400 23229 8420
rect 23085 8392 23229 8400
rect 23085 8391 23121 8392
rect 23193 8391 23229 8392
rect 23295 8425 23332 8426
rect 23295 8424 23333 8425
rect 23295 8416 23359 8424
rect 23295 8396 23304 8416
rect 23324 8402 23359 8416
rect 23379 8402 23382 8422
rect 23324 8397 23382 8402
rect 23324 8396 23359 8397
rect 22561 8359 22598 8388
rect 22562 8357 22598 8359
rect 22774 8357 22811 8388
rect 22562 8335 22811 8357
rect 22643 8329 22754 8335
rect 22643 8321 22684 8329
rect 22643 8301 22651 8321
rect 22670 8301 22684 8321
rect 22643 8299 22684 8301
rect 22712 8321 22754 8329
rect 22712 8301 22728 8321
rect 22747 8301 22754 8321
rect 22712 8299 22754 8301
rect 22643 8284 22754 8299
rect 22982 8289 23019 8388
rect 23295 8384 23359 8396
rect 22645 8281 22749 8284
rect 22433 8244 22554 8254
rect 22433 8242 22502 8244
rect 22433 8201 22446 8242
rect 22483 8203 22502 8242
rect 22539 8203 22554 8244
rect 22483 8201 22554 8203
rect 22433 8183 22554 8201
rect 20006 8116 20078 8117
rect 17690 8115 19028 8116
rect 17690 8113 18401 8115
rect 18550 8074 18614 8078
rect 20925 8076 20991 8124
rect 22225 8139 22290 8173
rect 22645 8139 22749 8141
rect 22980 8139 23021 8289
rect 23399 8281 23426 8536
rect 23488 8526 23568 8537
rect 23488 8500 23505 8526
rect 23545 8500 23568 8526
rect 23488 8473 23568 8500
rect 23488 8447 23509 8473
rect 23549 8447 23568 8473
rect 23488 8428 23568 8447
rect 23488 8402 23512 8428
rect 23552 8402 23568 8428
rect 23488 8351 23568 8402
rect 22225 8136 23021 8139
rect 23400 8150 23426 8281
rect 23490 8151 23560 8351
rect 23400 8136 23428 8150
rect 22225 8101 23428 8136
rect 23489 8129 23561 8151
rect 18550 8065 18624 8074
rect 17065 7582 17179 7586
rect 16270 7578 16370 7582
rect 16270 7574 16332 7578
rect 16270 7548 16277 7574
rect 16303 7552 16332 7574
rect 16358 7552 16370 7578
rect 16303 7548 16370 7552
rect 16270 7545 16370 7548
rect 16438 7545 16473 7582
rect 16535 7579 16894 7582
rect 16535 7574 16757 7579
rect 16535 7550 16548 7574
rect 16572 7555 16757 7574
rect 16781 7555 16894 7579
rect 16572 7550 16894 7555
rect 16535 7546 16894 7550
rect 16961 7579 17179 7582
rect 16961 7578 17144 7579
rect 16961 7574 17087 7578
rect 16961 7554 16972 7574
rect 16992 7554 17087 7574
rect 17111 7555 17144 7578
rect 17168 7555 17179 7579
rect 17111 7554 17179 7555
rect 16961 7547 17179 7554
rect 16961 7546 17002 7547
rect 16437 7520 16473 7545
rect 16285 7493 16322 7494
rect 16381 7493 16418 7494
rect 16437 7493 16444 7520
rect 16185 7484 16323 7493
rect 16185 7464 16294 7484
rect 16314 7464 16323 7484
rect 16185 7457 16323 7464
rect 16381 7490 16444 7493
rect 16465 7493 16473 7520
rect 16492 7493 16529 7494
rect 16465 7490 16529 7493
rect 16381 7484 16529 7490
rect 16381 7464 16390 7484
rect 16410 7464 16500 7484
rect 16520 7464 16529 7484
rect 16185 7455 16281 7457
rect 16381 7454 16529 7464
rect 16588 7484 16625 7494
rect 16700 7493 16737 7494
rect 16681 7491 16737 7493
rect 16588 7464 16596 7484
rect 16616 7464 16625 7484
rect 16437 7453 16473 7454
rect 16285 7322 16322 7323
rect 16588 7322 16625 7464
rect 16650 7484 16737 7491
rect 16650 7481 16708 7484
rect 16650 7461 16655 7481
rect 16676 7464 16708 7481
rect 16728 7464 16737 7484
rect 16676 7461 16737 7464
rect 16650 7454 16737 7461
rect 16796 7484 16833 7494
rect 16796 7464 16804 7484
rect 16824 7464 16833 7484
rect 16650 7453 16681 7454
rect 16796 7385 16833 7464
rect 16863 7493 16894 7546
rect 17065 7544 17179 7547
rect 17108 7512 17179 7544
rect 18354 8023 18438 8048
rect 18354 7995 18369 8023
rect 18413 7995 18438 8023
rect 18354 7966 18438 7995
rect 18550 8017 18564 8065
rect 18601 8017 18624 8065
rect 18550 7989 18624 8017
rect 18354 7938 18366 7966
rect 18410 7938 18438 7966
rect 18354 7917 18438 7938
rect 16913 7493 16950 7494
rect 16863 7484 16950 7493
rect 16863 7464 16921 7484
rect 16941 7464 16950 7484
rect 16863 7454 16950 7464
rect 17009 7484 17046 7494
rect 17009 7464 17017 7484
rect 17037 7464 17046 7484
rect 16863 7453 16894 7454
rect 16858 7385 16968 7398
rect 17009 7385 17046 7464
rect 16796 7383 17046 7385
rect 16796 7380 16897 7383
rect 16796 7361 16861 7380
rect 16858 7353 16861 7361
rect 16890 7353 16897 7380
rect 16925 7356 16935 7383
rect 16964 7361 17046 7383
rect 16964 7356 16968 7361
rect 16925 7353 16968 7356
rect 16858 7339 16968 7353
rect 16284 7321 16625 7322
rect 16209 7318 16625 7321
rect 16209 7316 16632 7318
rect 16209 7296 16212 7316
rect 16232 7296 16632 7316
rect 15400 4955 16040 5043
rect 15400 4604 15484 4955
rect 15966 4924 16010 4930
rect 15966 4898 15974 4924
rect 15999 4898 16010 4924
rect 15966 4849 16010 4898
rect 15966 4829 16363 4849
rect 16383 4829 16386 4849
rect 15966 4824 16386 4829
rect 15966 4823 16311 4824
rect 15966 4819 16010 4823
rect 16273 4822 16310 4823
rect 15627 4792 15737 4806
rect 15627 4789 15670 4792
rect 15627 4784 15631 4789
rect 15549 4762 15631 4784
rect 15660 4762 15670 4789
rect 15698 4765 15705 4792
rect 15734 4784 15737 4792
rect 15734 4765 15799 4784
rect 15698 4762 15799 4765
rect 15549 4760 15799 4762
rect 15549 4681 15586 4760
rect 15627 4747 15737 4760
rect 15701 4691 15732 4692
rect 15549 4661 15558 4681
rect 15578 4661 15586 4681
rect 15549 4651 15586 4661
rect 15645 4681 15732 4691
rect 15645 4661 15654 4681
rect 15674 4661 15732 4681
rect 15645 4652 15732 4661
rect 15645 4651 15682 4652
rect 15400 4598 15509 4604
rect 15701 4599 15732 4652
rect 15762 4681 15799 4760
rect 15914 4691 15945 4692
rect 15762 4661 15771 4681
rect 15791 4661 15799 4681
rect 15762 4651 15799 4661
rect 15858 4684 15945 4691
rect 15858 4681 15919 4684
rect 15858 4661 15867 4681
rect 15887 4664 15919 4681
rect 15940 4664 15945 4684
rect 15887 4661 15945 4664
rect 15858 4654 15945 4661
rect 15970 4681 16007 4819
rect 16122 4691 16158 4692
rect 15970 4661 15979 4681
rect 15999 4661 16007 4681
rect 15858 4652 15914 4654
rect 15858 4651 15895 4652
rect 15970 4651 16007 4661
rect 16066 4681 16214 4691
rect 16314 4688 16410 4690
rect 16066 4661 16075 4681
rect 16095 4661 16185 4681
rect 16205 4661 16214 4681
rect 16066 4655 16214 4661
rect 16066 4652 16130 4655
rect 16066 4651 16103 4652
rect 16122 4625 16130 4652
rect 16151 4652 16214 4655
rect 16272 4681 16410 4688
rect 16272 4661 16281 4681
rect 16301 4661 16410 4681
rect 16272 4652 16410 4661
rect 16151 4625 16158 4652
rect 16177 4651 16214 4652
rect 16273 4651 16310 4652
rect 16122 4600 16158 4625
rect 15593 4598 15634 4599
rect 15400 4591 15634 4598
rect 15400 4571 15603 4591
rect 15623 4571 15634 4591
rect 15400 4563 15634 4571
rect 15701 4595 16060 4599
rect 15701 4590 16023 4595
rect 15701 4566 15814 4590
rect 15838 4571 16023 4590
rect 16047 4571 16060 4595
rect 15838 4566 16060 4571
rect 15701 4563 16060 4566
rect 16122 4563 16157 4600
rect 16225 4597 16325 4600
rect 16225 4593 16292 4597
rect 16225 4567 16237 4593
rect 16263 4571 16292 4593
rect 16318 4571 16325 4597
rect 16263 4567 16325 4571
rect 16225 4563 16325 4567
rect 15400 4545 15509 4563
rect 15701 4542 15732 4563
rect 16122 4542 16158 4563
rect 15544 4541 15581 4542
rect 15543 4532 15581 4541
rect 15543 4512 15552 4532
rect 15572 4512 15581 4532
rect 15543 4504 15581 4512
rect 15647 4536 15732 4542
rect 15757 4541 15794 4542
rect 15647 4516 15655 4536
rect 15675 4516 15732 4536
rect 15647 4508 15732 4516
rect 15756 4532 15794 4541
rect 15756 4512 15765 4532
rect 15785 4512 15794 4532
rect 15647 4507 15683 4508
rect 15756 4504 15794 4512
rect 15860 4536 15945 4542
rect 15965 4541 16002 4542
rect 15860 4516 15868 4536
rect 15888 4535 15945 4536
rect 15888 4516 15917 4535
rect 15860 4515 15917 4516
rect 15938 4515 15945 4535
rect 15860 4508 15945 4515
rect 15964 4532 16002 4541
rect 15964 4512 15973 4532
rect 15993 4512 16002 4532
rect 15860 4507 15896 4508
rect 15964 4504 16002 4512
rect 16068 4537 16212 4542
rect 16068 4536 16121 4537
rect 16068 4516 16076 4536
rect 16096 4517 16121 4536
rect 16154 4536 16212 4537
rect 16154 4517 16184 4536
rect 16096 4516 16184 4517
rect 16204 4516 16212 4536
rect 16068 4508 16212 4516
rect 16068 4507 16104 4508
rect 16176 4507 16212 4508
rect 16278 4541 16315 4542
rect 16278 4540 16316 4541
rect 16278 4532 16342 4540
rect 16278 4512 16287 4532
rect 16307 4518 16342 4532
rect 16362 4518 16365 4538
rect 16307 4513 16365 4518
rect 16307 4512 16342 4513
rect 15544 4475 15581 4504
rect 15545 4473 15581 4475
rect 15757 4473 15794 4504
rect 15545 4451 15794 4473
rect 15626 4445 15737 4451
rect 15626 4437 15667 4445
rect 15626 4417 15634 4437
rect 15653 4417 15667 4437
rect 15626 4415 15667 4417
rect 15695 4437 15737 4445
rect 15695 4417 15711 4437
rect 15730 4417 15737 4437
rect 15695 4415 15737 4417
rect 15626 4400 15737 4415
rect 15965 4383 16002 4504
rect 16278 4500 16342 4512
rect 16382 4389 16409 4652
rect 16436 4398 16472 4405
rect 16436 4389 16442 4398
rect 16360 4385 16442 4389
rect 16241 4383 16442 4385
rect 15965 4360 16442 4383
rect 16465 4360 16472 4398
rect 15965 4357 16472 4360
rect 16241 4356 16409 4357
rect 16436 4354 16472 4357
rect 16554 4256 16632 7296
rect 17688 6549 17747 6559
rect 17688 6521 17701 6549
rect 17729 6521 17747 6549
rect 17688 6472 17747 6521
rect 17294 6337 17462 6338
rect 17698 6337 17745 6472
rect 17294 6311 17745 6337
rect 17294 6309 17462 6311
rect 17294 6042 17321 6309
rect 17698 6305 17745 6311
rect 17361 6182 17425 6194
rect 17701 6190 17738 6305
rect 17966 6279 18077 6294
rect 17966 6277 18008 6279
rect 17966 6257 17973 6277
rect 17992 6257 18008 6277
rect 17966 6249 18008 6257
rect 18036 6277 18077 6279
rect 18036 6257 18050 6277
rect 18069 6257 18077 6277
rect 18036 6249 18077 6257
rect 17966 6243 18077 6249
rect 17909 6221 18158 6243
rect 17909 6190 17946 6221
rect 18122 6219 18158 6221
rect 18122 6190 18159 6219
rect 17361 6181 17396 6182
rect 17338 6176 17396 6181
rect 17338 6156 17341 6176
rect 17361 6162 17396 6176
rect 17416 6162 17425 6182
rect 17361 6154 17425 6162
rect 17387 6153 17425 6154
rect 17388 6152 17425 6153
rect 17491 6186 17527 6187
rect 17599 6186 17635 6187
rect 17491 6178 17635 6186
rect 17491 6158 17499 6178
rect 17519 6158 17607 6178
rect 17627 6158 17635 6178
rect 17491 6152 17635 6158
rect 17701 6182 17739 6190
rect 17807 6186 17843 6187
rect 17701 6162 17710 6182
rect 17730 6162 17739 6182
rect 17701 6153 17739 6162
rect 17758 6179 17843 6186
rect 17758 6159 17765 6179
rect 17786 6178 17843 6179
rect 17786 6159 17815 6178
rect 17758 6158 17815 6159
rect 17835 6158 17843 6178
rect 17701 6152 17738 6153
rect 17758 6152 17843 6158
rect 17909 6182 17947 6190
rect 18020 6186 18056 6187
rect 17909 6162 17918 6182
rect 17938 6162 17947 6182
rect 17909 6153 17947 6162
rect 17971 6178 18056 6186
rect 17971 6158 18028 6178
rect 18048 6158 18056 6178
rect 17909 6152 17946 6153
rect 17971 6152 18056 6158
rect 18122 6182 18160 6190
rect 18122 6162 18131 6182
rect 18151 6162 18160 6182
rect 18122 6153 18160 6162
rect 18122 6152 18159 6153
rect 17545 6131 17581 6152
rect 17971 6131 18002 6152
rect 18182 6137 18239 6145
rect 18182 6131 18190 6137
rect 17378 6127 17478 6131
rect 17378 6123 17440 6127
rect 17378 6097 17385 6123
rect 17411 6101 17440 6123
rect 17466 6101 17478 6127
rect 17411 6097 17478 6101
rect 17378 6094 17478 6097
rect 17546 6094 17581 6131
rect 17643 6128 18002 6131
rect 17643 6123 17865 6128
rect 17643 6099 17656 6123
rect 17680 6104 17865 6123
rect 17889 6104 18002 6128
rect 17680 6099 18002 6104
rect 17643 6095 18002 6099
rect 18069 6123 18190 6131
rect 18069 6103 18080 6123
rect 18100 6114 18190 6123
rect 18216 6114 18239 6137
rect 18100 6103 18239 6114
rect 18069 6101 18239 6103
rect 18069 6096 18190 6101
rect 18069 6095 18110 6096
rect 17545 6069 17581 6094
rect 17393 6042 17430 6043
rect 17489 6042 17526 6043
rect 17545 6042 17552 6069
rect 17293 6033 17431 6042
rect 17293 6013 17402 6033
rect 17422 6013 17431 6033
rect 17293 6006 17431 6013
rect 17489 6039 17552 6042
rect 17573 6042 17581 6069
rect 17600 6042 17637 6043
rect 17573 6039 17637 6042
rect 17489 6033 17637 6039
rect 17489 6013 17498 6033
rect 17518 6013 17608 6033
rect 17628 6013 17637 6033
rect 17293 6004 17389 6006
rect 17489 6003 17637 6013
rect 17696 6033 17733 6043
rect 17808 6042 17845 6043
rect 17789 6040 17845 6042
rect 17696 6013 17704 6033
rect 17724 6013 17733 6033
rect 17545 6002 17581 6003
rect 17393 5871 17430 5872
rect 17696 5871 17733 6013
rect 17758 6033 17845 6040
rect 17758 6030 17816 6033
rect 17758 6010 17763 6030
rect 17784 6013 17816 6030
rect 17836 6013 17845 6033
rect 17784 6010 17845 6013
rect 17758 6003 17845 6010
rect 17904 6033 17941 6043
rect 17904 6013 17912 6033
rect 17932 6013 17941 6033
rect 17758 6002 17789 6003
rect 17904 5934 17941 6013
rect 17971 6042 18002 6095
rect 18021 6042 18058 6043
rect 17971 6033 18058 6042
rect 17971 6013 18029 6033
rect 18049 6013 18058 6033
rect 17971 6003 18058 6013
rect 18117 6033 18154 6043
rect 18117 6013 18125 6033
rect 18145 6013 18154 6033
rect 17971 6002 18002 6003
rect 17966 5934 18076 5947
rect 18117 5934 18154 6013
rect 17904 5932 18154 5934
rect 17904 5929 18005 5932
rect 17904 5910 17969 5929
rect 17966 5902 17969 5910
rect 17998 5902 18005 5929
rect 18033 5905 18043 5932
rect 18072 5910 18154 5932
rect 18072 5905 18076 5910
rect 18033 5902 18076 5905
rect 17966 5888 18076 5902
rect 17392 5870 17733 5871
rect 17317 5865 17733 5870
rect 17317 5845 17320 5865
rect 17340 5845 17734 5865
rect 17543 5812 17580 5822
rect 17543 5775 17552 5812
rect 17569 5775 17580 5812
rect 17543 5754 17580 5775
rect 17252 4815 17420 4816
rect 17549 4815 17578 5754
rect 17691 5140 17734 5845
rect 17692 5132 17734 5140
rect 17692 5121 17737 5132
rect 17692 5083 17702 5121
rect 17727 5083 17737 5121
rect 17692 5074 17737 5083
rect 17252 4789 17696 4815
rect 17252 4787 17420 4789
rect 17252 4520 17279 4787
rect 17549 4785 17578 4789
rect 17319 4660 17383 4672
rect 17659 4668 17696 4789
rect 17924 4757 18035 4772
rect 17924 4755 17966 4757
rect 17924 4735 17931 4755
rect 17950 4735 17966 4755
rect 17924 4727 17966 4735
rect 17994 4755 18035 4757
rect 17994 4735 18008 4755
rect 18027 4735 18035 4755
rect 17994 4727 18035 4735
rect 17924 4721 18035 4727
rect 17867 4699 18116 4721
rect 17867 4668 17904 4699
rect 18080 4697 18116 4699
rect 18080 4668 18117 4697
rect 17319 4659 17354 4660
rect 17296 4654 17354 4659
rect 17296 4634 17299 4654
rect 17319 4640 17354 4654
rect 17374 4640 17383 4660
rect 17319 4632 17383 4640
rect 17345 4631 17383 4632
rect 17346 4630 17383 4631
rect 17449 4664 17485 4665
rect 17557 4664 17593 4665
rect 17449 4656 17593 4664
rect 17449 4636 17457 4656
rect 17477 4636 17565 4656
rect 17585 4636 17593 4656
rect 17449 4630 17593 4636
rect 17659 4660 17697 4668
rect 17765 4664 17801 4665
rect 17659 4640 17668 4660
rect 17688 4640 17697 4660
rect 17659 4631 17697 4640
rect 17716 4657 17801 4664
rect 17716 4637 17723 4657
rect 17744 4656 17801 4657
rect 17744 4637 17773 4656
rect 17716 4636 17773 4637
rect 17793 4636 17801 4656
rect 17659 4630 17696 4631
rect 17716 4630 17801 4636
rect 17867 4660 17905 4668
rect 17978 4664 18014 4665
rect 17867 4640 17876 4660
rect 17896 4640 17905 4660
rect 17867 4631 17905 4640
rect 17929 4656 18014 4664
rect 17929 4636 17986 4656
rect 18006 4636 18014 4656
rect 17867 4630 17904 4631
rect 17929 4630 18014 4636
rect 18080 4660 18118 4668
rect 18080 4640 18089 4660
rect 18109 4640 18118 4660
rect 18080 4631 18118 4640
rect 18080 4630 18117 4631
rect 17503 4609 17539 4630
rect 17929 4609 17960 4630
rect 18354 4613 18446 7917
rect 18552 6150 18624 7989
rect 19654 7939 19726 7956
rect 19654 7891 19666 7939
rect 19712 7891 19726 7939
rect 20194 7919 20235 7921
rect 20466 7919 20570 7921
rect 20925 7919 20990 8076
rect 22225 7944 22290 8101
rect 22645 8099 22749 8101
rect 22980 8099 23021 8101
rect 23489 8081 23503 8129
rect 23549 8081 23561 8129
rect 23489 8064 23561 8081
rect 24591 8031 24663 9870
rect 24769 8103 24861 11407
rect 25255 11390 25286 11411
rect 25676 11390 25712 11411
rect 25098 11389 25135 11390
rect 25097 11380 25135 11389
rect 25097 11360 25106 11380
rect 25126 11360 25135 11380
rect 25097 11352 25135 11360
rect 25201 11384 25286 11390
rect 25311 11389 25348 11390
rect 25201 11364 25209 11384
rect 25229 11364 25286 11384
rect 25201 11356 25286 11364
rect 25310 11380 25348 11389
rect 25310 11360 25319 11380
rect 25339 11360 25348 11380
rect 25201 11355 25237 11356
rect 25310 11352 25348 11360
rect 25414 11384 25499 11390
rect 25519 11389 25556 11390
rect 25414 11364 25422 11384
rect 25442 11383 25499 11384
rect 25442 11364 25471 11383
rect 25414 11363 25471 11364
rect 25492 11363 25499 11383
rect 25414 11356 25499 11363
rect 25518 11380 25556 11389
rect 25518 11360 25527 11380
rect 25547 11360 25556 11380
rect 25414 11355 25450 11356
rect 25518 11352 25556 11360
rect 25622 11384 25766 11390
rect 25622 11364 25630 11384
rect 25650 11364 25738 11384
rect 25758 11364 25766 11384
rect 25622 11356 25766 11364
rect 25622 11355 25658 11356
rect 25730 11355 25766 11356
rect 25832 11389 25869 11390
rect 25832 11388 25870 11389
rect 25832 11380 25896 11388
rect 25832 11360 25841 11380
rect 25861 11366 25896 11380
rect 25916 11366 25919 11386
rect 25861 11361 25919 11366
rect 25861 11360 25896 11361
rect 25098 11323 25135 11352
rect 25099 11321 25135 11323
rect 25311 11321 25348 11352
rect 25099 11299 25348 11321
rect 25180 11293 25291 11299
rect 25180 11285 25221 11293
rect 25180 11265 25188 11285
rect 25207 11265 25221 11285
rect 25180 11263 25221 11265
rect 25249 11285 25291 11293
rect 25249 11265 25265 11285
rect 25284 11265 25291 11285
rect 25249 11263 25291 11265
rect 25180 11248 25291 11263
rect 25519 11231 25556 11352
rect 25832 11348 25896 11360
rect 25637 11231 25666 11235
rect 25936 11233 25963 11500
rect 25795 11231 25963 11233
rect 25519 11205 25963 11231
rect 25478 10937 25523 10946
rect 25478 10899 25488 10937
rect 25513 10899 25523 10937
rect 25478 10888 25523 10899
rect 25481 10880 25523 10888
rect 25481 10175 25524 10880
rect 25637 10266 25666 11205
rect 25795 11204 25963 11205
rect 25635 10245 25672 10266
rect 25635 10208 25646 10245
rect 25663 10208 25672 10245
rect 25635 10198 25672 10208
rect 25481 10155 25875 10175
rect 25895 10155 25898 10175
rect 25482 10150 25898 10155
rect 25482 10149 25823 10150
rect 25139 10118 25249 10132
rect 25139 10115 25182 10118
rect 25139 10110 25143 10115
rect 25061 10088 25143 10110
rect 25172 10088 25182 10115
rect 25210 10091 25217 10118
rect 25246 10110 25249 10118
rect 25246 10091 25311 10110
rect 25210 10088 25311 10091
rect 25061 10086 25311 10088
rect 25061 10007 25098 10086
rect 25139 10073 25249 10086
rect 25213 10017 25244 10018
rect 25061 9987 25070 10007
rect 25090 9987 25098 10007
rect 25061 9977 25098 9987
rect 25157 10007 25244 10017
rect 25157 9987 25166 10007
rect 25186 9987 25244 10007
rect 25157 9978 25244 9987
rect 25157 9977 25194 9978
rect 25213 9925 25244 9978
rect 25274 10007 25311 10086
rect 25426 10017 25457 10018
rect 25274 9987 25283 10007
rect 25303 9987 25311 10007
rect 25274 9977 25311 9987
rect 25370 10010 25457 10017
rect 25370 10007 25431 10010
rect 25370 9987 25379 10007
rect 25399 9990 25431 10007
rect 25452 9990 25457 10010
rect 25399 9987 25457 9990
rect 25370 9980 25457 9987
rect 25482 10007 25519 10149
rect 25785 10148 25822 10149
rect 25634 10017 25670 10018
rect 25482 9987 25491 10007
rect 25511 9987 25519 10007
rect 25370 9978 25426 9980
rect 25370 9977 25407 9978
rect 25482 9977 25519 9987
rect 25578 10007 25726 10017
rect 25826 10014 25922 10016
rect 25578 9987 25587 10007
rect 25607 9987 25697 10007
rect 25717 9987 25726 10007
rect 25578 9981 25726 9987
rect 25578 9978 25642 9981
rect 25578 9977 25615 9978
rect 25634 9951 25642 9978
rect 25663 9978 25726 9981
rect 25784 10007 25922 10014
rect 25784 9987 25793 10007
rect 25813 9987 25922 10007
rect 25784 9978 25922 9987
rect 25663 9951 25670 9978
rect 25689 9977 25726 9978
rect 25785 9977 25822 9978
rect 25634 9926 25670 9951
rect 25105 9924 25146 9925
rect 25025 9919 25146 9924
rect 24976 9917 25146 9919
rect 24976 9906 25115 9917
rect 24976 9883 24999 9906
rect 25025 9897 25115 9906
rect 25135 9897 25146 9917
rect 25025 9889 25146 9897
rect 25213 9921 25572 9925
rect 25213 9916 25535 9921
rect 25213 9892 25326 9916
rect 25350 9897 25535 9916
rect 25559 9897 25572 9921
rect 25350 9892 25572 9897
rect 25213 9889 25572 9892
rect 25634 9889 25669 9926
rect 25737 9923 25837 9926
rect 25737 9919 25804 9923
rect 25737 9893 25749 9919
rect 25775 9897 25804 9919
rect 25830 9897 25837 9923
rect 25775 9893 25837 9897
rect 25737 9889 25837 9893
rect 25025 9883 25033 9889
rect 24976 9875 25033 9883
rect 25213 9868 25244 9889
rect 25634 9868 25670 9889
rect 25056 9867 25093 9868
rect 25055 9858 25093 9867
rect 25055 9838 25064 9858
rect 25084 9838 25093 9858
rect 25055 9830 25093 9838
rect 25159 9862 25244 9868
rect 25269 9867 25306 9868
rect 25159 9842 25167 9862
rect 25187 9842 25244 9862
rect 25159 9834 25244 9842
rect 25268 9858 25306 9867
rect 25268 9838 25277 9858
rect 25297 9838 25306 9858
rect 25159 9833 25195 9834
rect 25268 9830 25306 9838
rect 25372 9862 25457 9868
rect 25477 9867 25514 9868
rect 25372 9842 25380 9862
rect 25400 9861 25457 9862
rect 25400 9842 25429 9861
rect 25372 9841 25429 9842
rect 25450 9841 25457 9861
rect 25372 9834 25457 9841
rect 25476 9858 25514 9867
rect 25476 9838 25485 9858
rect 25505 9838 25514 9858
rect 25372 9833 25408 9834
rect 25476 9830 25514 9838
rect 25580 9862 25724 9868
rect 25580 9842 25588 9862
rect 25608 9842 25696 9862
rect 25716 9842 25724 9862
rect 25580 9834 25724 9842
rect 25580 9833 25616 9834
rect 25688 9833 25724 9834
rect 25790 9867 25827 9868
rect 25790 9866 25828 9867
rect 25790 9858 25854 9866
rect 25790 9838 25799 9858
rect 25819 9844 25854 9858
rect 25874 9844 25877 9864
rect 25819 9839 25877 9844
rect 25819 9838 25854 9839
rect 25056 9801 25093 9830
rect 25057 9799 25093 9801
rect 25269 9799 25306 9830
rect 25057 9777 25306 9799
rect 25138 9771 25249 9777
rect 25138 9763 25179 9771
rect 25138 9743 25146 9763
rect 25165 9743 25179 9763
rect 25138 9741 25179 9743
rect 25207 9763 25249 9771
rect 25207 9743 25223 9763
rect 25242 9743 25249 9763
rect 25207 9741 25249 9743
rect 25138 9726 25249 9741
rect 25477 9715 25514 9830
rect 25790 9826 25854 9838
rect 25470 9709 25517 9715
rect 25894 9711 25921 9978
rect 25753 9709 25921 9711
rect 25470 9683 25921 9709
rect 25470 9548 25517 9683
rect 25753 9682 25921 9683
rect 25468 9499 25527 9548
rect 25468 9471 25486 9499
rect 25514 9471 25527 9499
rect 25468 9461 25527 9471
rect 26583 8724 26661 11764
rect 26583 8704 26983 8724
rect 27003 8704 27006 8724
rect 26583 8702 27006 8704
rect 26590 8699 27006 8702
rect 26590 8698 26931 8699
rect 26247 8667 26357 8681
rect 26247 8664 26290 8667
rect 26247 8659 26251 8664
rect 26169 8637 26251 8659
rect 26280 8637 26290 8664
rect 26318 8640 26325 8667
rect 26354 8659 26357 8667
rect 26354 8640 26419 8659
rect 26318 8637 26419 8640
rect 26169 8635 26419 8637
rect 26169 8556 26206 8635
rect 26247 8622 26357 8635
rect 26321 8566 26352 8567
rect 26169 8536 26178 8556
rect 26198 8536 26206 8556
rect 26169 8526 26206 8536
rect 26265 8556 26352 8566
rect 26265 8536 26274 8556
rect 26294 8536 26352 8556
rect 26265 8527 26352 8536
rect 26265 8526 26302 8527
rect 26039 8473 26150 8476
rect 26321 8474 26352 8527
rect 26382 8556 26419 8635
rect 26534 8566 26565 8567
rect 26382 8536 26391 8556
rect 26411 8536 26419 8556
rect 26382 8526 26419 8536
rect 26478 8559 26565 8566
rect 26478 8556 26539 8559
rect 26478 8536 26487 8556
rect 26507 8539 26539 8556
rect 26560 8539 26565 8559
rect 26507 8536 26565 8539
rect 26478 8529 26565 8536
rect 26590 8556 26627 8698
rect 26893 8697 26930 8698
rect 26742 8566 26778 8567
rect 26590 8536 26599 8556
rect 26619 8536 26627 8556
rect 26478 8527 26534 8529
rect 26478 8526 26515 8527
rect 26590 8526 26627 8536
rect 26686 8556 26834 8566
rect 26934 8563 27030 8565
rect 26686 8536 26695 8556
rect 26715 8536 26805 8556
rect 26825 8536 26834 8556
rect 26686 8530 26834 8536
rect 26686 8527 26750 8530
rect 26686 8526 26723 8527
rect 26742 8500 26750 8527
rect 26771 8527 26834 8530
rect 26892 8556 27030 8563
rect 26892 8536 26901 8556
rect 26921 8536 27030 8556
rect 26892 8527 27030 8536
rect 26771 8500 26778 8527
rect 26797 8526 26834 8527
rect 26893 8526 26930 8527
rect 26742 8475 26778 8500
rect 26213 8473 26254 8474
rect 26039 8466 26254 8473
rect 26039 8465 26104 8466
rect 26039 8441 26047 8465
rect 26071 8442 26104 8465
rect 26128 8446 26223 8466
rect 26243 8446 26254 8466
rect 26128 8442 26254 8446
rect 26071 8441 26254 8442
rect 26039 8438 26254 8441
rect 26321 8470 26680 8474
rect 26321 8465 26643 8470
rect 26321 8441 26434 8465
rect 26458 8446 26643 8465
rect 26667 8446 26680 8470
rect 26458 8441 26680 8446
rect 26321 8438 26680 8441
rect 26742 8438 26777 8475
rect 26845 8472 26945 8475
rect 26845 8468 26912 8472
rect 26845 8442 26857 8468
rect 26883 8446 26912 8468
rect 26938 8446 26945 8472
rect 26883 8442 26945 8446
rect 26845 8438 26945 8442
rect 26039 8434 26150 8438
rect 26321 8417 26352 8438
rect 26742 8417 26778 8438
rect 26164 8416 26201 8417
rect 26163 8407 26201 8416
rect 26163 8387 26172 8407
rect 26192 8387 26201 8407
rect 26163 8379 26201 8387
rect 26267 8411 26352 8417
rect 26377 8416 26414 8417
rect 26267 8391 26275 8411
rect 26295 8391 26352 8411
rect 26267 8383 26352 8391
rect 26376 8407 26414 8416
rect 26376 8387 26385 8407
rect 26405 8387 26414 8407
rect 26267 8382 26303 8383
rect 26376 8379 26414 8387
rect 26480 8411 26565 8417
rect 26585 8416 26622 8417
rect 26480 8391 26488 8411
rect 26508 8410 26565 8411
rect 26508 8391 26537 8410
rect 26480 8390 26537 8391
rect 26558 8390 26565 8410
rect 26480 8383 26565 8390
rect 26584 8407 26622 8416
rect 26584 8387 26593 8407
rect 26613 8387 26622 8407
rect 26480 8382 26516 8383
rect 26584 8379 26622 8387
rect 26688 8411 26832 8417
rect 26688 8391 26696 8411
rect 26716 8410 26804 8411
rect 26716 8391 26750 8410
rect 26688 8388 26750 8391
rect 26774 8391 26804 8410
rect 26824 8391 26832 8411
rect 26774 8388 26832 8391
rect 26688 8383 26832 8388
rect 26688 8382 26724 8383
rect 26796 8382 26832 8383
rect 26898 8416 26935 8417
rect 26898 8415 26936 8416
rect 26898 8407 26962 8415
rect 26898 8387 26907 8407
rect 26927 8393 26962 8407
rect 26982 8393 26985 8413
rect 26927 8388 26985 8393
rect 26927 8387 26962 8388
rect 26164 8350 26201 8379
rect 26165 8348 26201 8350
rect 26377 8348 26414 8379
rect 26165 8326 26414 8348
rect 26246 8320 26357 8326
rect 26246 8312 26287 8320
rect 26246 8292 26254 8312
rect 26273 8292 26287 8312
rect 26246 8290 26287 8292
rect 26315 8312 26357 8320
rect 26315 8292 26331 8312
rect 26350 8292 26357 8312
rect 26315 8290 26357 8292
rect 26246 8275 26357 8290
rect 26585 8264 26622 8379
rect 26898 8375 26962 8387
rect 26581 8258 26636 8264
rect 27002 8260 27029 8527
rect 26861 8258 27029 8260
rect 26581 8233 27029 8258
rect 27342 8318 27448 13516
rect 30614 13506 30637 13532
rect 30677 13506 30694 13532
rect 30614 13495 30694 13506
rect 30756 13496 30783 13751
rect 31161 13743 31202 13893
rect 31873 13862 32996 13893
rect 33846 13897 33945 13905
rect 33846 13894 33898 13897
rect 31628 13831 31749 13849
rect 31628 13829 31699 13831
rect 31628 13788 31643 13829
rect 31680 13790 31699 13829
rect 31736 13790 31749 13831
rect 31680 13788 31749 13790
rect 31628 13778 31749 13788
rect 30823 13636 30887 13648
rect 31163 13644 31200 13743
rect 31428 13733 31539 13744
rect 31428 13731 31470 13733
rect 31428 13711 31435 13731
rect 31454 13711 31470 13731
rect 31428 13703 31470 13711
rect 31498 13731 31539 13733
rect 31498 13711 31512 13731
rect 31531 13711 31539 13731
rect 31498 13703 31539 13711
rect 31428 13697 31539 13703
rect 31371 13675 31620 13697
rect 31371 13644 31408 13675
rect 31584 13673 31620 13675
rect 31584 13644 31621 13673
rect 30823 13635 30858 13636
rect 30800 13630 30858 13635
rect 30800 13610 30803 13630
rect 30823 13616 30858 13630
rect 30878 13616 30887 13636
rect 30823 13608 30887 13616
rect 30849 13607 30887 13608
rect 30850 13606 30887 13607
rect 30953 13640 30989 13641
rect 31061 13640 31097 13641
rect 30953 13632 31097 13640
rect 30953 13612 30961 13632
rect 30981 13612 31069 13632
rect 31089 13612 31097 13632
rect 30953 13606 31097 13612
rect 31163 13636 31201 13644
rect 31269 13640 31305 13641
rect 31163 13616 31172 13636
rect 31192 13616 31201 13636
rect 31163 13607 31201 13616
rect 31220 13633 31305 13640
rect 31220 13613 31227 13633
rect 31248 13632 31305 13633
rect 31248 13613 31277 13632
rect 31220 13612 31277 13613
rect 31297 13612 31305 13632
rect 31163 13606 31200 13607
rect 31220 13606 31305 13612
rect 31371 13636 31409 13644
rect 31482 13640 31518 13641
rect 31371 13616 31380 13636
rect 31400 13616 31409 13636
rect 31371 13607 31409 13616
rect 31433 13632 31518 13640
rect 31433 13612 31490 13632
rect 31510 13612 31518 13632
rect 31371 13606 31408 13607
rect 31433 13606 31518 13612
rect 31584 13636 31622 13644
rect 31584 13616 31593 13636
rect 31613 13616 31622 13636
rect 31677 13626 31742 13778
rect 31895 13752 31950 13862
rect 32934 13824 32993 13862
rect 33846 13859 33854 13894
rect 33879 13859 33898 13894
rect 33923 13886 33945 13897
rect 34896 13898 36235 13905
rect 34896 13895 34948 13898
rect 33923 13885 34790 13886
rect 33923 13859 34791 13885
rect 33846 13849 34791 13859
rect 33846 13847 33945 13849
rect 32934 13806 32956 13824
rect 32974 13806 32993 13824
rect 32934 13784 32993 13806
rect 33201 13820 33733 13825
rect 33201 13800 34087 13820
rect 34107 13800 34110 13820
rect 34746 13816 34791 13849
rect 34896 13860 34904 13895
rect 34929 13860 34948 13895
rect 34973 13860 36235 13898
rect 34896 13851 36235 13860
rect 34896 13848 34985 13851
rect 35524 13849 36235 13851
rect 33201 13796 34110 13800
rect 31584 13607 31622 13616
rect 31675 13619 31742 13626
rect 31584 13606 31621 13607
rect 31007 13585 31043 13606
rect 31433 13585 31464 13606
rect 31675 13598 31692 13619
rect 31728 13598 31742 13619
rect 31894 13639 31950 13752
rect 33201 13749 33244 13796
rect 33694 13795 34110 13796
rect 34742 13796 35135 13816
rect 35155 13796 35158 13816
rect 33694 13794 34035 13795
rect 33351 13763 33461 13777
rect 33351 13760 33394 13763
rect 33351 13755 33355 13760
rect 33189 13748 33244 13749
rect 31894 13621 31913 13639
rect 31931 13621 31950 13639
rect 31894 13601 31950 13621
rect 32933 13725 33244 13748
rect 32933 13707 32958 13725
rect 32976 13713 33244 13725
rect 33273 13733 33355 13755
rect 33384 13733 33394 13760
rect 33422 13736 33429 13763
rect 33458 13755 33461 13763
rect 33458 13736 33523 13755
rect 33422 13733 33523 13736
rect 33273 13731 33523 13733
rect 32976 13707 32998 13713
rect 31675 13585 31742 13598
rect 30840 13581 30940 13585
rect 30840 13577 30902 13581
rect 30840 13551 30847 13577
rect 30873 13555 30902 13577
rect 30928 13555 30940 13581
rect 30873 13551 30940 13555
rect 30840 13548 30940 13551
rect 31008 13548 31043 13585
rect 31105 13582 31464 13585
rect 31105 13577 31327 13582
rect 31105 13553 31118 13577
rect 31142 13558 31327 13577
rect 31351 13558 31464 13582
rect 31142 13553 31464 13558
rect 31105 13549 31464 13553
rect 31531 13579 31742 13585
rect 31531 13577 31692 13579
rect 31531 13557 31542 13577
rect 31562 13557 31692 13577
rect 31531 13550 31692 13557
rect 31531 13549 31572 13550
rect 31007 13523 31043 13548
rect 30855 13496 30892 13497
rect 30951 13496 30988 13497
rect 31007 13496 31014 13523
rect 30755 13487 30893 13496
rect 30755 13467 30864 13487
rect 30884 13467 30893 13487
rect 30755 13460 30893 13467
rect 30951 13493 31014 13496
rect 31035 13496 31043 13523
rect 31062 13496 31099 13497
rect 31035 13493 31099 13496
rect 30951 13487 31099 13493
rect 30951 13467 30960 13487
rect 30980 13467 31070 13487
rect 31090 13467 31099 13487
rect 30755 13458 30851 13460
rect 30951 13457 31099 13467
rect 31158 13487 31195 13497
rect 31270 13496 31307 13497
rect 31251 13494 31307 13496
rect 31158 13467 31166 13487
rect 31186 13467 31195 13487
rect 31007 13456 31043 13457
rect 30855 13325 30892 13326
rect 31158 13325 31195 13467
rect 31220 13487 31307 13494
rect 31220 13484 31278 13487
rect 31220 13464 31225 13484
rect 31246 13467 31278 13484
rect 31298 13467 31307 13487
rect 31246 13464 31307 13467
rect 31220 13457 31307 13464
rect 31366 13487 31403 13497
rect 31366 13467 31374 13487
rect 31394 13467 31403 13487
rect 31220 13456 31251 13457
rect 31366 13388 31403 13467
rect 31433 13496 31464 13549
rect 31677 13542 31692 13550
rect 31732 13542 31742 13579
rect 32933 13568 32998 13707
rect 33273 13652 33310 13731
rect 33351 13718 33461 13731
rect 33425 13662 33456 13663
rect 33273 13632 33282 13652
rect 33302 13632 33310 13652
rect 31677 13533 31742 13542
rect 31890 13540 31955 13561
rect 31890 13522 31915 13540
rect 31933 13522 31955 13540
rect 32933 13550 32956 13568
rect 32974 13550 32998 13568
rect 32933 13533 32998 13550
rect 33153 13614 33221 13627
rect 33273 13622 33310 13632
rect 33369 13652 33456 13662
rect 33369 13632 33378 13652
rect 33398 13632 33456 13652
rect 33369 13623 33456 13632
rect 33369 13622 33406 13623
rect 33153 13572 33160 13614
rect 33209 13572 33221 13614
rect 33153 13569 33221 13572
rect 33425 13570 33456 13623
rect 33486 13652 33523 13731
rect 33638 13662 33669 13663
rect 33486 13632 33495 13652
rect 33515 13632 33523 13652
rect 33486 13622 33523 13632
rect 33582 13655 33669 13662
rect 33582 13652 33643 13655
rect 33582 13632 33591 13652
rect 33611 13635 33643 13652
rect 33664 13635 33669 13655
rect 33611 13632 33669 13635
rect 33582 13625 33669 13632
rect 33694 13652 33731 13794
rect 33997 13793 34034 13794
rect 34742 13791 35158 13796
rect 34742 13790 35083 13791
rect 34399 13759 34509 13773
rect 34399 13756 34442 13759
rect 34399 13751 34403 13756
rect 34321 13729 34403 13751
rect 34432 13729 34442 13756
rect 34470 13732 34477 13759
rect 34506 13751 34509 13759
rect 34506 13732 34571 13751
rect 34470 13729 34571 13732
rect 34321 13727 34571 13729
rect 33846 13662 33882 13663
rect 33694 13632 33703 13652
rect 33723 13632 33731 13652
rect 33582 13623 33638 13625
rect 33582 13622 33619 13623
rect 33694 13622 33731 13632
rect 33790 13652 33938 13662
rect 34038 13659 34134 13661
rect 33790 13632 33799 13652
rect 33819 13632 33909 13652
rect 33929 13632 33938 13652
rect 33790 13626 33938 13632
rect 33790 13623 33854 13626
rect 33790 13622 33827 13623
rect 33846 13596 33854 13623
rect 33875 13623 33938 13626
rect 33996 13652 34134 13659
rect 33996 13632 34005 13652
rect 34025 13632 34134 13652
rect 33996 13623 34134 13632
rect 34321 13648 34358 13727
rect 34399 13714 34509 13727
rect 34473 13658 34504 13659
rect 34321 13628 34330 13648
rect 34350 13628 34358 13648
rect 33875 13596 33882 13623
rect 33901 13622 33938 13623
rect 33997 13622 34034 13623
rect 33846 13571 33882 13596
rect 33317 13569 33358 13570
rect 33153 13562 33358 13569
rect 33153 13551 33327 13562
rect 31483 13496 31520 13497
rect 31433 13487 31520 13496
rect 31433 13467 31491 13487
rect 31511 13467 31520 13487
rect 31433 13457 31520 13467
rect 31579 13487 31616 13497
rect 31579 13467 31587 13487
rect 31607 13467 31616 13487
rect 31433 13456 31464 13457
rect 31428 13388 31538 13401
rect 31579 13388 31616 13467
rect 31890 13446 31955 13522
rect 33153 13518 33161 13551
rect 33154 13509 33161 13518
rect 33210 13542 33327 13551
rect 33347 13542 33358 13562
rect 33210 13534 33358 13542
rect 33425 13566 33784 13570
rect 33425 13561 33747 13566
rect 33425 13537 33538 13561
rect 33562 13542 33747 13561
rect 33771 13542 33784 13566
rect 33562 13537 33784 13542
rect 33425 13534 33784 13537
rect 33846 13534 33881 13571
rect 33949 13568 34049 13571
rect 33949 13564 34016 13568
rect 33949 13538 33961 13564
rect 33987 13542 34016 13564
rect 34042 13542 34049 13568
rect 33987 13538 34049 13542
rect 33949 13534 34049 13538
rect 33210 13518 33221 13534
rect 33210 13509 33218 13518
rect 33425 13513 33456 13534
rect 33846 13513 33882 13534
rect 33268 13512 33305 13513
rect 32933 13469 32998 13488
rect 32933 13451 32958 13469
rect 32976 13451 32998 13469
rect 31366 13386 31616 13388
rect 31366 13383 31467 13386
rect 31366 13364 31431 13383
rect 31428 13356 31431 13364
rect 31460 13356 31467 13383
rect 31495 13359 31505 13386
rect 31534 13364 31616 13386
rect 31639 13411 31956 13446
rect 31534 13359 31538 13364
rect 31495 13356 31538 13359
rect 31428 13342 31538 13356
rect 30854 13324 31195 13325
rect 30779 13322 31195 13324
rect 31639 13322 31679 13411
rect 31890 13384 31955 13411
rect 31890 13366 31913 13384
rect 31931 13366 31955 13384
rect 31890 13346 31955 13366
rect 30776 13319 31679 13322
rect 30776 13299 30782 13319
rect 30802 13299 31679 13319
rect 30776 13295 31679 13299
rect 31639 13292 31679 13295
rect 31891 13285 31956 13306
rect 30109 13277 30770 13278
rect 30109 13270 31043 13277
rect 30109 13269 31015 13270
rect 30109 13249 30960 13269
rect 30992 13250 31015 13269
rect 31040 13250 31043 13270
rect 30992 13249 31043 13250
rect 30109 13242 31043 13249
rect 29708 13200 29876 13201
rect 30111 13200 30150 13242
rect 30939 13240 31043 13242
rect 31008 13238 31043 13240
rect 31891 13267 31915 13285
rect 31933 13267 31956 13285
rect 31891 13220 31956 13267
rect 29708 13174 30152 13200
rect 29708 13172 29876 13174
rect 29708 12821 29735 13172
rect 30111 13168 30152 13174
rect 29775 12961 29839 12973
rect 30115 12969 30152 13168
rect 30614 13195 30686 13212
rect 30614 13156 30622 13195
rect 30667 13156 30686 13195
rect 30380 13058 30491 13073
rect 30380 13056 30422 13058
rect 30380 13036 30387 13056
rect 30406 13036 30422 13056
rect 30380 13028 30422 13036
rect 30450 13056 30491 13058
rect 30450 13036 30464 13056
rect 30483 13036 30491 13056
rect 30450 13028 30491 13036
rect 30380 13022 30491 13028
rect 30323 13000 30572 13022
rect 30323 12969 30360 13000
rect 30536 12998 30572 13000
rect 30536 12969 30573 12998
rect 29775 12960 29810 12961
rect 29752 12955 29810 12960
rect 29752 12935 29755 12955
rect 29775 12941 29810 12955
rect 29830 12941 29839 12961
rect 29775 12933 29839 12941
rect 29801 12932 29839 12933
rect 29802 12931 29839 12932
rect 29905 12965 29941 12966
rect 30013 12965 30049 12966
rect 29905 12957 30049 12965
rect 29905 12937 29913 12957
rect 29933 12937 30021 12957
rect 30041 12937 30049 12957
rect 29905 12931 30049 12937
rect 30115 12961 30153 12969
rect 30221 12965 30257 12966
rect 30115 12941 30124 12961
rect 30144 12941 30153 12961
rect 30115 12932 30153 12941
rect 30172 12958 30257 12965
rect 30172 12938 30179 12958
rect 30200 12957 30257 12958
rect 30200 12938 30229 12957
rect 30172 12937 30229 12938
rect 30249 12937 30257 12957
rect 30115 12931 30152 12932
rect 30172 12931 30257 12937
rect 30323 12961 30361 12969
rect 30434 12965 30470 12966
rect 30323 12941 30332 12961
rect 30352 12941 30361 12961
rect 30323 12932 30361 12941
rect 30385 12957 30470 12965
rect 30385 12937 30442 12957
rect 30462 12937 30470 12957
rect 30323 12931 30360 12932
rect 30385 12931 30470 12937
rect 30536 12961 30574 12969
rect 30536 12941 30545 12961
rect 30565 12941 30574 12961
rect 30536 12932 30574 12941
rect 30614 12946 30686 13156
rect 30756 13190 31956 13220
rect 30756 13189 31200 13190
rect 30756 13187 30924 13189
rect 30614 12932 30697 12946
rect 30536 12931 30573 12932
rect 29959 12910 29995 12931
rect 30385 12910 30416 12931
rect 30614 12910 30631 12932
rect 29792 12906 29892 12910
rect 29792 12902 29854 12906
rect 29792 12876 29799 12902
rect 29825 12880 29854 12902
rect 29880 12880 29892 12906
rect 29825 12876 29892 12880
rect 29792 12873 29892 12876
rect 29960 12873 29995 12910
rect 30057 12907 30416 12910
rect 30057 12902 30279 12907
rect 30057 12878 30070 12902
rect 30094 12883 30279 12902
rect 30303 12883 30416 12907
rect 30094 12878 30416 12883
rect 30057 12874 30416 12878
rect 30483 12902 30631 12910
rect 30483 12882 30494 12902
rect 30514 12899 30631 12902
rect 30684 12899 30697 12932
rect 30514 12882 30697 12899
rect 30483 12875 30697 12882
rect 30483 12874 30524 12875
rect 30614 12874 30697 12875
rect 29959 12848 29995 12873
rect 29807 12821 29844 12822
rect 29903 12821 29940 12822
rect 29959 12821 29966 12848
rect 29707 12812 29845 12821
rect 29707 12792 29816 12812
rect 29836 12792 29845 12812
rect 29707 12785 29845 12792
rect 29903 12818 29966 12821
rect 29987 12821 29995 12848
rect 30014 12821 30051 12822
rect 29987 12818 30051 12821
rect 29903 12812 30051 12818
rect 29903 12792 29912 12812
rect 29932 12792 30022 12812
rect 30042 12792 30051 12812
rect 29707 12783 29803 12785
rect 29903 12782 30051 12792
rect 30110 12812 30147 12822
rect 30222 12821 30259 12822
rect 30203 12819 30259 12821
rect 30110 12792 30118 12812
rect 30138 12792 30147 12812
rect 29959 12781 29995 12782
rect 29807 12650 29844 12651
rect 30110 12650 30147 12792
rect 30172 12812 30259 12819
rect 30172 12809 30230 12812
rect 30172 12789 30177 12809
rect 30198 12792 30230 12809
rect 30250 12792 30259 12812
rect 30198 12789 30259 12792
rect 30172 12782 30259 12789
rect 30318 12812 30355 12822
rect 30318 12792 30326 12812
rect 30346 12792 30355 12812
rect 30172 12781 30203 12782
rect 30318 12713 30355 12792
rect 30385 12821 30416 12874
rect 30622 12841 30636 12874
rect 30689 12841 30697 12874
rect 30622 12835 30697 12841
rect 30622 12830 30692 12835
rect 30435 12821 30472 12822
rect 30385 12812 30472 12821
rect 30385 12792 30443 12812
rect 30463 12792 30472 12812
rect 30385 12782 30472 12792
rect 30531 12812 30568 12822
rect 30756 12817 30783 13187
rect 30823 12957 30887 12969
rect 31163 12965 31200 13189
rect 31671 13170 31735 13172
rect 31667 13158 31735 13170
rect 31667 13125 31678 13158
rect 31718 13125 31735 13158
rect 31667 13115 31735 13125
rect 31428 13054 31539 13069
rect 31428 13052 31470 13054
rect 31428 13032 31435 13052
rect 31454 13032 31470 13052
rect 31428 13024 31470 13032
rect 31498 13052 31539 13054
rect 31498 13032 31512 13052
rect 31531 13032 31539 13052
rect 31498 13024 31539 13032
rect 31428 13018 31539 13024
rect 31371 12996 31620 13018
rect 31371 12965 31408 12996
rect 31584 12994 31620 12996
rect 31584 12965 31621 12994
rect 30823 12956 30858 12957
rect 30800 12951 30858 12956
rect 30800 12931 30803 12951
rect 30823 12937 30858 12951
rect 30878 12937 30887 12957
rect 30823 12929 30887 12937
rect 30849 12928 30887 12929
rect 30850 12927 30887 12928
rect 30953 12961 30989 12962
rect 31061 12961 31097 12962
rect 30953 12953 31097 12961
rect 30953 12933 30961 12953
rect 30981 12933 31069 12953
rect 31089 12933 31097 12953
rect 30953 12927 31097 12933
rect 31163 12957 31201 12965
rect 31269 12961 31305 12962
rect 31163 12937 31172 12957
rect 31192 12937 31201 12957
rect 31163 12928 31201 12937
rect 31220 12954 31305 12961
rect 31220 12934 31227 12954
rect 31248 12953 31305 12954
rect 31248 12934 31277 12953
rect 31220 12933 31277 12934
rect 31297 12933 31305 12953
rect 31163 12927 31200 12928
rect 31220 12927 31305 12933
rect 31371 12957 31409 12965
rect 31482 12961 31518 12962
rect 31371 12937 31380 12957
rect 31400 12937 31409 12957
rect 31371 12928 31409 12937
rect 31433 12953 31518 12961
rect 31433 12933 31490 12953
rect 31510 12933 31518 12953
rect 31371 12927 31408 12928
rect 31433 12927 31518 12933
rect 31584 12957 31622 12965
rect 31584 12937 31593 12957
rect 31613 12937 31622 12957
rect 31584 12928 31622 12937
rect 31671 12931 31735 13115
rect 31891 12989 31956 13190
rect 32933 13250 32998 13451
rect 33154 13325 33218 13509
rect 33267 13503 33305 13512
rect 33267 13483 33276 13503
rect 33296 13483 33305 13503
rect 33267 13475 33305 13483
rect 33371 13507 33456 13513
rect 33481 13512 33518 13513
rect 33371 13487 33379 13507
rect 33399 13487 33456 13507
rect 33371 13479 33456 13487
rect 33480 13503 33518 13512
rect 33480 13483 33489 13503
rect 33509 13483 33518 13503
rect 33371 13478 33407 13479
rect 33480 13475 33518 13483
rect 33584 13507 33669 13513
rect 33689 13512 33726 13513
rect 33584 13487 33592 13507
rect 33612 13506 33669 13507
rect 33612 13487 33641 13506
rect 33584 13486 33641 13487
rect 33662 13486 33669 13506
rect 33584 13479 33669 13486
rect 33688 13503 33726 13512
rect 33688 13483 33697 13503
rect 33717 13483 33726 13503
rect 33584 13478 33620 13479
rect 33688 13475 33726 13483
rect 33792 13507 33936 13513
rect 33792 13487 33800 13507
rect 33820 13487 33908 13507
rect 33928 13487 33936 13507
rect 33792 13479 33936 13487
rect 33792 13478 33828 13479
rect 33900 13478 33936 13479
rect 34002 13512 34039 13513
rect 34002 13511 34040 13512
rect 34002 13503 34066 13511
rect 34002 13483 34011 13503
rect 34031 13489 34066 13503
rect 34086 13489 34089 13509
rect 34031 13484 34089 13489
rect 34031 13483 34066 13484
rect 33268 13446 33305 13475
rect 33269 13444 33305 13446
rect 33481 13444 33518 13475
rect 33269 13422 33518 13444
rect 33350 13416 33461 13422
rect 33350 13408 33391 13416
rect 33350 13388 33358 13408
rect 33377 13388 33391 13408
rect 33350 13386 33391 13388
rect 33419 13408 33461 13416
rect 33419 13388 33435 13408
rect 33454 13388 33461 13408
rect 33419 13386 33461 13388
rect 33350 13371 33461 13386
rect 33154 13315 33222 13325
rect 33154 13282 33171 13315
rect 33211 13282 33222 13315
rect 33154 13270 33222 13282
rect 33154 13268 33218 13270
rect 33689 13251 33726 13475
rect 34002 13471 34066 13483
rect 34106 13253 34133 13623
rect 34321 13618 34358 13628
rect 34417 13648 34504 13658
rect 34417 13628 34426 13648
rect 34446 13628 34504 13648
rect 34417 13619 34504 13628
rect 34417 13618 34454 13619
rect 34197 13605 34267 13610
rect 34192 13599 34267 13605
rect 34192 13566 34200 13599
rect 34253 13566 34267 13599
rect 34473 13566 34504 13619
rect 34534 13648 34571 13727
rect 34686 13658 34717 13659
rect 34534 13628 34543 13648
rect 34563 13628 34571 13648
rect 34534 13618 34571 13628
rect 34630 13651 34717 13658
rect 34630 13648 34691 13651
rect 34630 13628 34639 13648
rect 34659 13631 34691 13648
rect 34712 13631 34717 13651
rect 34659 13628 34717 13631
rect 34630 13621 34717 13628
rect 34742 13648 34779 13790
rect 35045 13789 35082 13790
rect 34894 13658 34930 13659
rect 34742 13628 34751 13648
rect 34771 13628 34779 13648
rect 34630 13619 34686 13621
rect 34630 13618 34667 13619
rect 34742 13618 34779 13628
rect 34838 13648 34986 13658
rect 35086 13655 35182 13657
rect 34838 13628 34847 13648
rect 34867 13628 34957 13648
rect 34977 13628 34986 13648
rect 34838 13622 34986 13628
rect 34838 13619 34902 13622
rect 34838 13618 34875 13619
rect 34894 13592 34902 13619
rect 34923 13619 34986 13622
rect 35044 13648 35182 13655
rect 35044 13628 35053 13648
rect 35073 13628 35182 13648
rect 35044 13619 35182 13628
rect 34923 13592 34930 13619
rect 34949 13618 34986 13619
rect 35045 13618 35082 13619
rect 34894 13567 34930 13592
rect 34192 13565 34275 13566
rect 34365 13565 34406 13566
rect 34192 13558 34406 13565
rect 34192 13541 34375 13558
rect 34192 13508 34205 13541
rect 34258 13538 34375 13541
rect 34395 13538 34406 13558
rect 34258 13530 34406 13538
rect 34473 13562 34832 13566
rect 34473 13557 34795 13562
rect 34473 13533 34586 13557
rect 34610 13538 34795 13557
rect 34819 13538 34832 13562
rect 34610 13533 34832 13538
rect 34473 13530 34832 13533
rect 34894 13530 34929 13567
rect 34997 13564 35097 13567
rect 34997 13560 35064 13564
rect 34997 13534 35009 13560
rect 35035 13538 35064 13560
rect 35090 13538 35097 13564
rect 35035 13534 35097 13538
rect 34997 13530 35097 13534
rect 34258 13508 34275 13530
rect 34473 13509 34504 13530
rect 34894 13509 34930 13530
rect 34316 13508 34353 13509
rect 34192 13494 34275 13508
rect 33965 13251 34133 13253
rect 33689 13250 34133 13251
rect 32933 13220 34133 13250
rect 34203 13284 34275 13494
rect 34315 13499 34353 13508
rect 34315 13479 34324 13499
rect 34344 13479 34353 13499
rect 34315 13471 34353 13479
rect 34419 13503 34504 13509
rect 34529 13508 34566 13509
rect 34419 13483 34427 13503
rect 34447 13483 34504 13503
rect 34419 13475 34504 13483
rect 34528 13499 34566 13508
rect 34528 13479 34537 13499
rect 34557 13479 34566 13499
rect 34419 13474 34455 13475
rect 34528 13471 34566 13479
rect 34632 13503 34717 13509
rect 34737 13508 34774 13509
rect 34632 13483 34640 13503
rect 34660 13502 34717 13503
rect 34660 13483 34689 13502
rect 34632 13482 34689 13483
rect 34710 13482 34717 13502
rect 34632 13475 34717 13482
rect 34736 13499 34774 13508
rect 34736 13479 34745 13499
rect 34765 13479 34774 13499
rect 34632 13474 34668 13475
rect 34736 13471 34774 13479
rect 34840 13503 34984 13509
rect 34840 13483 34848 13503
rect 34868 13483 34956 13503
rect 34976 13483 34984 13503
rect 34840 13475 34984 13483
rect 34840 13474 34876 13475
rect 34948 13474 34984 13475
rect 35050 13508 35087 13509
rect 35050 13507 35088 13508
rect 35050 13499 35114 13507
rect 35050 13479 35059 13499
rect 35079 13485 35114 13499
rect 35134 13485 35137 13505
rect 35079 13480 35137 13485
rect 35079 13479 35114 13480
rect 34316 13442 34353 13471
rect 34317 13440 34353 13442
rect 34529 13440 34566 13471
rect 34317 13418 34566 13440
rect 34398 13412 34509 13418
rect 34398 13404 34439 13412
rect 34398 13384 34406 13404
rect 34425 13384 34439 13404
rect 34398 13382 34439 13384
rect 34467 13404 34509 13412
rect 34467 13384 34483 13404
rect 34502 13384 34509 13404
rect 34467 13382 34509 13384
rect 34398 13367 34509 13382
rect 34203 13245 34222 13284
rect 34267 13245 34275 13284
rect 34203 13228 34275 13245
rect 34737 13272 34774 13471
rect 35050 13467 35114 13479
rect 34737 13266 34778 13272
rect 35154 13268 35181 13619
rect 35476 13606 35571 13632
rect 35312 13584 35376 13603
rect 35312 13545 35325 13584
rect 35359 13545 35376 13584
rect 35312 13526 35376 13545
rect 35013 13266 35181 13268
rect 34737 13240 35181 13266
rect 32933 13173 32998 13220
rect 32933 13155 32956 13173
rect 32974 13155 32998 13173
rect 33846 13200 33881 13202
rect 33846 13198 33950 13200
rect 34739 13198 34778 13240
rect 35013 13239 35181 13240
rect 33846 13191 34780 13198
rect 33846 13190 33897 13191
rect 33846 13170 33849 13190
rect 33874 13171 33897 13190
rect 33929 13171 34780 13191
rect 33874 13170 34780 13171
rect 33846 13163 34780 13170
rect 34119 13162 34780 13163
rect 32933 13134 32998 13155
rect 33210 13145 33250 13148
rect 33210 13141 34113 13145
rect 33210 13121 34087 13141
rect 34107 13121 34113 13141
rect 33210 13118 34113 13121
rect 32934 13074 32999 13094
rect 32934 13056 32958 13074
rect 32976 13056 32999 13074
rect 32934 13029 32999 13056
rect 33210 13029 33250 13118
rect 33694 13116 34110 13118
rect 33694 13115 34035 13116
rect 33351 13084 33461 13098
rect 33351 13081 33394 13084
rect 33351 13076 33355 13081
rect 32933 12994 33250 13029
rect 33273 13054 33355 13076
rect 33384 13054 33394 13081
rect 33422 13057 33429 13084
rect 33458 13076 33461 13084
rect 33458 13057 33523 13076
rect 33422 13054 33523 13057
rect 33273 13052 33523 13054
rect 31891 12971 31913 12989
rect 31931 12971 31956 12989
rect 31891 12952 31956 12971
rect 31584 12927 31621 12928
rect 31007 12906 31043 12927
rect 31433 12906 31464 12927
rect 31671 12922 31679 12931
rect 31668 12906 31679 12922
rect 30840 12902 30940 12906
rect 30840 12898 30902 12902
rect 30840 12872 30847 12898
rect 30873 12876 30902 12898
rect 30928 12876 30940 12902
rect 30873 12872 30940 12876
rect 30840 12869 30940 12872
rect 31008 12869 31043 12906
rect 31105 12903 31464 12906
rect 31105 12898 31327 12903
rect 31105 12874 31118 12898
rect 31142 12879 31327 12898
rect 31351 12879 31464 12903
rect 31142 12874 31464 12879
rect 31105 12870 31464 12874
rect 31531 12898 31679 12906
rect 31531 12878 31542 12898
rect 31562 12889 31679 12898
rect 31728 12922 31735 12931
rect 31728 12889 31736 12922
rect 32934 12918 32999 12994
rect 33273 12973 33310 13052
rect 33351 13039 33461 13052
rect 33425 12983 33456 12984
rect 33273 12953 33282 12973
rect 33302 12953 33310 12973
rect 33273 12943 33310 12953
rect 33369 12973 33456 12983
rect 33369 12953 33378 12973
rect 33398 12953 33456 12973
rect 33369 12944 33456 12953
rect 33369 12943 33406 12944
rect 31562 12878 31736 12889
rect 31531 12871 31736 12878
rect 31531 12870 31572 12871
rect 31007 12844 31043 12869
rect 30855 12817 30892 12818
rect 30951 12817 30988 12818
rect 31007 12817 31014 12844
rect 30531 12792 30539 12812
rect 30559 12792 30568 12812
rect 30385 12781 30416 12782
rect 30380 12713 30490 12726
rect 30531 12713 30568 12792
rect 30755 12808 30893 12817
rect 30755 12788 30864 12808
rect 30884 12788 30893 12808
rect 30755 12781 30893 12788
rect 30951 12814 31014 12817
rect 31035 12817 31043 12844
rect 31062 12817 31099 12818
rect 31035 12814 31099 12817
rect 30951 12808 31099 12814
rect 30951 12788 30960 12808
rect 30980 12788 31070 12808
rect 31090 12788 31099 12808
rect 30755 12779 30851 12781
rect 30951 12778 31099 12788
rect 31158 12808 31195 12818
rect 31270 12817 31307 12818
rect 31251 12815 31307 12817
rect 31158 12788 31166 12808
rect 31186 12788 31195 12808
rect 31007 12777 31043 12778
rect 30318 12711 30568 12713
rect 30318 12708 30419 12711
rect 30318 12689 30383 12708
rect 30380 12681 30383 12689
rect 30412 12681 30419 12708
rect 30447 12684 30457 12711
rect 30486 12689 30568 12711
rect 30486 12684 30490 12689
rect 30447 12681 30490 12684
rect 30380 12667 30490 12681
rect 29806 12649 30147 12650
rect 29731 12644 30147 12649
rect 30855 12646 30892 12647
rect 31158 12646 31195 12788
rect 31220 12808 31307 12815
rect 31220 12805 31278 12808
rect 31220 12785 31225 12805
rect 31246 12788 31278 12805
rect 31298 12788 31307 12808
rect 31246 12785 31307 12788
rect 31220 12778 31307 12785
rect 31366 12808 31403 12818
rect 31366 12788 31374 12808
rect 31394 12788 31403 12808
rect 31220 12777 31251 12778
rect 31366 12709 31403 12788
rect 31433 12817 31464 12870
rect 31668 12868 31736 12871
rect 31668 12826 31680 12868
rect 31729 12826 31736 12868
rect 31483 12817 31520 12818
rect 31433 12808 31520 12817
rect 31433 12788 31491 12808
rect 31511 12788 31520 12808
rect 31433 12778 31520 12788
rect 31579 12808 31616 12818
rect 31668 12813 31736 12826
rect 31891 12890 31956 12907
rect 31891 12872 31915 12890
rect 31933 12872 31956 12890
rect 32934 12900 32956 12918
rect 32974 12900 32999 12918
rect 32934 12879 32999 12900
rect 33147 12898 33212 12907
rect 31579 12788 31587 12808
rect 31607 12788 31616 12808
rect 31433 12777 31464 12778
rect 31428 12709 31538 12722
rect 31579 12709 31616 12788
rect 31891 12733 31956 12872
rect 33147 12861 33157 12898
rect 33197 12890 33212 12898
rect 33425 12891 33456 12944
rect 33486 12973 33523 13052
rect 33638 12983 33669 12984
rect 33486 12953 33495 12973
rect 33515 12953 33523 12973
rect 33486 12943 33523 12953
rect 33582 12976 33669 12983
rect 33582 12973 33643 12976
rect 33582 12953 33591 12973
rect 33611 12956 33643 12973
rect 33664 12956 33669 12976
rect 33611 12953 33669 12956
rect 33582 12946 33669 12953
rect 33694 12973 33731 13115
rect 33997 13114 34034 13115
rect 35314 13055 35376 13526
rect 35476 13565 35502 13606
rect 35538 13565 35571 13606
rect 35476 13269 35571 13565
rect 35476 13225 35491 13269
rect 35551 13225 35571 13269
rect 35476 13205 35571 13225
rect 36188 13136 36231 13849
rect 36771 13791 36917 13802
rect 36771 13775 38153 13791
rect 36771 13770 38180 13775
rect 36771 13764 36863 13770
rect 36771 13667 36803 13764
rect 36841 13673 36863 13764
rect 36901 13673 38180 13770
rect 41330 13675 41400 13928
rect 41869 13925 41910 13927
rect 42141 13925 42245 13927
rect 41462 13923 42656 13925
rect 41462 13890 42658 13923
rect 41462 13876 41490 13890
rect 41464 13745 41490 13876
rect 41869 13887 42658 13890
rect 36841 13667 38180 13673
rect 36771 13640 38180 13667
rect 38050 13565 38180 13640
rect 41322 13624 41402 13675
rect 41322 13598 41338 13624
rect 41378 13598 41402 13624
rect 41322 13579 41402 13598
rect 36188 13116 36582 13136
rect 36602 13116 36605 13136
rect 36189 13111 36605 13116
rect 36189 13110 36530 13111
rect 35846 13079 35956 13093
rect 35846 13076 35889 13079
rect 35846 13071 35850 13076
rect 35309 13003 35384 13055
rect 35768 13049 35850 13071
rect 35879 13049 35889 13076
rect 35917 13052 35924 13079
rect 35953 13071 35956 13079
rect 35953 13052 36018 13071
rect 35917 13049 36018 13052
rect 35768 13047 36018 13049
rect 35678 13003 35724 13004
rect 33846 12983 33882 12984
rect 33694 12953 33703 12973
rect 33723 12953 33731 12973
rect 33582 12944 33638 12946
rect 33582 12943 33619 12944
rect 33694 12943 33731 12953
rect 33790 12973 33938 12983
rect 34038 12980 34134 12982
rect 33790 12953 33799 12973
rect 33819 12953 33909 12973
rect 33929 12953 33938 12973
rect 33790 12947 33938 12953
rect 33790 12944 33854 12947
rect 33790 12943 33827 12944
rect 33846 12917 33854 12944
rect 33875 12944 33938 12947
rect 33996 12973 34134 12980
rect 33996 12953 34005 12973
rect 34025 12953 34134 12973
rect 33996 12944 34134 12953
rect 35309 12968 35724 13003
rect 33875 12917 33882 12944
rect 33901 12943 33938 12944
rect 33997 12943 34034 12944
rect 33846 12892 33882 12917
rect 33317 12890 33358 12891
rect 33197 12883 33358 12890
rect 33197 12863 33327 12883
rect 33347 12863 33358 12883
rect 33197 12861 33358 12863
rect 33147 12855 33358 12861
rect 33425 12887 33784 12891
rect 33425 12882 33747 12887
rect 33425 12858 33538 12882
rect 33562 12863 33747 12882
rect 33771 12863 33784 12887
rect 33562 12858 33784 12863
rect 33425 12855 33784 12858
rect 33846 12855 33881 12892
rect 33949 12889 34049 12892
rect 33949 12885 34016 12889
rect 33949 12859 33961 12885
rect 33987 12863 34016 12885
rect 34042 12863 34049 12889
rect 33987 12859 34049 12863
rect 33949 12855 34049 12859
rect 33147 12842 33214 12855
rect 31891 12727 31913 12733
rect 31366 12707 31616 12709
rect 31366 12704 31467 12707
rect 31366 12685 31431 12704
rect 31428 12677 31431 12685
rect 31460 12677 31467 12704
rect 31495 12680 31505 12707
rect 31534 12685 31616 12707
rect 31645 12715 31913 12727
rect 31931 12715 31956 12733
rect 31645 12692 31956 12715
rect 32939 12819 32995 12839
rect 32939 12801 32958 12819
rect 32976 12801 32995 12819
rect 31645 12691 31700 12692
rect 31534 12680 31538 12685
rect 31495 12677 31538 12680
rect 31428 12663 31538 12677
rect 30854 12645 31195 12646
rect 29731 12624 29734 12644
rect 29754 12624 30147 12644
rect 30779 12644 31195 12645
rect 31645 12644 31688 12691
rect 32939 12688 32995 12801
rect 33147 12821 33161 12842
rect 33197 12821 33214 12842
rect 33425 12834 33456 12855
rect 33846 12834 33882 12855
rect 33268 12833 33305 12834
rect 33147 12814 33214 12821
rect 33267 12824 33305 12833
rect 30779 12640 31688 12644
rect 30098 12591 30143 12624
rect 30779 12620 30782 12640
rect 30802 12620 31688 12640
rect 31156 12615 31688 12620
rect 31896 12634 31955 12656
rect 31896 12616 31915 12634
rect 31933 12616 31955 12634
rect 30944 12591 31043 12593
rect 30098 12581 31043 12591
rect 28655 12561 28714 12571
rect 28655 12533 28668 12561
rect 28696 12533 28714 12561
rect 30098 12555 30966 12581
rect 30099 12554 30966 12555
rect 30944 12543 30966 12554
rect 30991 12546 31010 12581
rect 31035 12546 31043 12581
rect 30991 12543 31043 12546
rect 31896 12545 31955 12616
rect 32939 12550 32994 12688
rect 33147 12662 33212 12814
rect 33267 12804 33276 12824
rect 33296 12804 33305 12824
rect 33267 12796 33305 12804
rect 33371 12828 33456 12834
rect 33481 12833 33518 12834
rect 33371 12808 33379 12828
rect 33399 12808 33456 12828
rect 33371 12800 33456 12808
rect 33480 12824 33518 12833
rect 33480 12804 33489 12824
rect 33509 12804 33518 12824
rect 33371 12799 33407 12800
rect 33480 12796 33518 12804
rect 33584 12828 33669 12834
rect 33689 12833 33726 12834
rect 33584 12808 33592 12828
rect 33612 12827 33669 12828
rect 33612 12808 33641 12827
rect 33584 12807 33641 12808
rect 33662 12807 33669 12827
rect 33584 12800 33669 12807
rect 33688 12824 33726 12833
rect 33688 12804 33697 12824
rect 33717 12804 33726 12824
rect 33584 12799 33620 12800
rect 33688 12796 33726 12804
rect 33792 12828 33936 12834
rect 33792 12808 33800 12828
rect 33820 12808 33908 12828
rect 33928 12808 33936 12828
rect 33792 12800 33936 12808
rect 33792 12799 33828 12800
rect 33900 12799 33936 12800
rect 34002 12833 34039 12834
rect 34002 12832 34040 12833
rect 34002 12824 34066 12832
rect 34002 12804 34011 12824
rect 34031 12810 34066 12824
rect 34086 12810 34089 12830
rect 34031 12805 34089 12810
rect 34031 12804 34066 12805
rect 33268 12767 33305 12796
rect 33269 12765 33305 12767
rect 33481 12765 33518 12796
rect 33269 12743 33518 12765
rect 33350 12737 33461 12743
rect 33350 12729 33391 12737
rect 33350 12709 33358 12729
rect 33377 12709 33391 12729
rect 33350 12707 33391 12709
rect 33419 12729 33461 12737
rect 33419 12709 33435 12729
rect 33454 12709 33461 12729
rect 33419 12707 33461 12709
rect 33350 12694 33461 12707
rect 33689 12697 33726 12796
rect 34002 12792 34066 12804
rect 33140 12652 33261 12662
rect 33140 12650 33209 12652
rect 33140 12609 33153 12650
rect 33190 12611 33209 12650
rect 33246 12611 33261 12652
rect 33190 12609 33261 12611
rect 33140 12591 33261 12609
rect 32932 12547 32996 12550
rect 33352 12547 33456 12553
rect 33687 12547 33728 12697
rect 34106 12689 34133 12944
rect 34195 12934 34275 12945
rect 34195 12908 34212 12934
rect 34252 12908 34275 12934
rect 34195 12881 34275 12908
rect 34195 12855 34216 12881
rect 34256 12855 34275 12881
rect 34195 12836 34275 12855
rect 34195 12810 34219 12836
rect 34259 12810 34275 12836
rect 34195 12759 34275 12810
rect 30944 12535 31043 12543
rect 30970 12534 31042 12535
rect 28655 12484 28714 12533
rect 30624 12508 30691 12527
rect 30624 12487 30641 12508
rect 28261 12349 28429 12350
rect 28665 12349 28712 12484
rect 28261 12323 28712 12349
rect 28261 12321 28429 12323
rect 28261 12054 28288 12321
rect 28665 12317 28712 12323
rect 30622 12442 30641 12487
rect 30671 12487 30691 12508
rect 30671 12442 30692 12487
rect 31161 12484 31202 12486
rect 31433 12484 31537 12486
rect 31893 12484 31957 12545
rect 28328 12194 28392 12206
rect 28668 12202 28705 12317
rect 28933 12291 29044 12306
rect 28933 12289 28975 12291
rect 28933 12269 28940 12289
rect 28959 12269 28975 12289
rect 28933 12261 28975 12269
rect 29003 12289 29044 12291
rect 29003 12269 29017 12289
rect 29036 12269 29044 12289
rect 29003 12261 29044 12269
rect 28933 12255 29044 12261
rect 28876 12233 29125 12255
rect 30622 12234 30692 12442
rect 30754 12449 31957 12484
rect 30754 12435 30782 12449
rect 30756 12304 30782 12435
rect 31161 12446 31957 12449
rect 32932 12544 33728 12547
rect 34107 12558 34133 12689
rect 34107 12544 34135 12558
rect 32932 12509 34135 12544
rect 34197 12551 34267 12759
rect 35309 12684 35384 12968
rect 35678 12885 35724 12968
rect 35768 12968 35805 13047
rect 35846 13034 35956 13047
rect 35920 12978 35951 12979
rect 35768 12948 35777 12968
rect 35797 12948 35805 12968
rect 35768 12938 35805 12948
rect 35864 12968 35951 12978
rect 35864 12948 35873 12968
rect 35893 12948 35951 12968
rect 35864 12939 35951 12948
rect 35864 12938 35901 12939
rect 35920 12886 35951 12939
rect 35981 12968 36018 13047
rect 36133 12978 36164 12979
rect 35981 12948 35990 12968
rect 36010 12948 36018 12968
rect 35981 12938 36018 12948
rect 36077 12971 36164 12978
rect 36077 12968 36138 12971
rect 36077 12948 36086 12968
rect 36106 12951 36138 12968
rect 36159 12951 36164 12971
rect 36106 12948 36164 12951
rect 36077 12941 36164 12948
rect 36189 12968 36226 13110
rect 36492 13109 36529 13110
rect 36341 12978 36377 12979
rect 36189 12948 36198 12968
rect 36218 12948 36226 12968
rect 36077 12939 36133 12941
rect 36077 12938 36114 12939
rect 36189 12938 36226 12948
rect 36285 12968 36433 12978
rect 36533 12975 36629 12977
rect 36285 12948 36294 12968
rect 36314 12948 36404 12968
rect 36424 12948 36433 12968
rect 36285 12942 36433 12948
rect 36285 12939 36349 12942
rect 36285 12938 36322 12939
rect 36341 12912 36349 12939
rect 36370 12939 36433 12942
rect 36491 12968 36629 12975
rect 36491 12948 36500 12968
rect 36520 12948 36629 12968
rect 36491 12939 36629 12948
rect 36370 12912 36377 12939
rect 36396 12938 36433 12939
rect 36492 12938 36529 12939
rect 36341 12887 36377 12912
rect 35812 12885 35853 12886
rect 35678 12878 35853 12885
rect 35476 12852 35562 12871
rect 35476 12811 35491 12852
rect 35545 12811 35562 12852
rect 35678 12858 35822 12878
rect 35842 12858 35853 12878
rect 35678 12850 35853 12858
rect 35920 12882 36279 12886
rect 35920 12877 36242 12882
rect 35920 12853 36033 12877
rect 36057 12858 36242 12877
rect 36266 12858 36279 12882
rect 36057 12853 36279 12858
rect 35920 12850 36279 12853
rect 36341 12850 36376 12887
rect 36444 12884 36544 12887
rect 36444 12880 36511 12884
rect 36444 12854 36456 12880
rect 36482 12858 36511 12880
rect 36537 12858 36544 12884
rect 36482 12854 36544 12858
rect 36444 12850 36544 12854
rect 35678 12846 35724 12850
rect 35920 12829 35951 12850
rect 36341 12829 36377 12850
rect 35763 12828 35800 12829
rect 35476 12775 35562 12811
rect 35762 12819 35800 12828
rect 35762 12799 35771 12819
rect 35791 12799 35800 12819
rect 35762 12791 35800 12799
rect 35866 12823 35951 12829
rect 35976 12828 36013 12829
rect 35866 12803 35874 12823
rect 35894 12803 35951 12823
rect 35866 12795 35951 12803
rect 35975 12819 36013 12828
rect 35975 12799 35984 12819
rect 36004 12799 36013 12819
rect 35866 12794 35902 12795
rect 35975 12791 36013 12799
rect 36079 12823 36164 12829
rect 36184 12828 36221 12829
rect 36079 12803 36087 12823
rect 36107 12822 36164 12823
rect 36107 12803 36136 12822
rect 36079 12802 36136 12803
rect 36157 12802 36164 12822
rect 36079 12795 36164 12802
rect 36183 12819 36221 12828
rect 36183 12799 36192 12819
rect 36212 12799 36221 12819
rect 36079 12794 36115 12795
rect 36183 12791 36221 12799
rect 36287 12823 36431 12829
rect 36287 12803 36295 12823
rect 36315 12803 36403 12823
rect 36423 12803 36431 12823
rect 36287 12795 36431 12803
rect 36287 12794 36323 12795
rect 32932 12448 32996 12509
rect 33352 12507 33456 12509
rect 33687 12507 33728 12509
rect 34197 12506 34218 12551
rect 34198 12485 34218 12506
rect 34248 12506 34267 12551
rect 35304 12642 35384 12684
rect 34248 12485 34265 12506
rect 34198 12466 34265 12485
rect 33847 12458 33919 12459
rect 33846 12450 33945 12458
rect 28876 12202 28913 12233
rect 29089 12231 29125 12233
rect 29089 12202 29126 12231
rect 28328 12193 28363 12194
rect 28305 12188 28363 12193
rect 28305 12168 28308 12188
rect 28328 12174 28363 12188
rect 28383 12174 28392 12194
rect 28328 12166 28392 12174
rect 28354 12165 28392 12166
rect 28355 12164 28392 12165
rect 28458 12198 28494 12199
rect 28566 12198 28602 12199
rect 28458 12190 28602 12198
rect 28458 12170 28466 12190
rect 28486 12170 28574 12190
rect 28594 12170 28602 12190
rect 28458 12164 28602 12170
rect 28668 12194 28706 12202
rect 28774 12198 28810 12199
rect 28668 12174 28677 12194
rect 28697 12174 28706 12194
rect 28668 12165 28706 12174
rect 28725 12191 28810 12198
rect 28725 12171 28732 12191
rect 28753 12190 28810 12191
rect 28753 12171 28782 12190
rect 28725 12170 28782 12171
rect 28802 12170 28810 12190
rect 28668 12164 28705 12165
rect 28725 12164 28810 12170
rect 28876 12194 28914 12202
rect 28987 12198 29023 12199
rect 28876 12174 28885 12194
rect 28905 12174 28914 12194
rect 28876 12165 28914 12174
rect 28938 12190 29023 12198
rect 28938 12170 28995 12190
rect 29015 12170 29023 12190
rect 28876 12164 28913 12165
rect 28938 12164 29023 12170
rect 29089 12194 29127 12202
rect 29089 12174 29098 12194
rect 29118 12174 29127 12194
rect 29089 12165 29127 12174
rect 30614 12183 30694 12234
rect 29089 12164 29126 12165
rect 28512 12143 28548 12164
rect 28938 12143 28969 12164
rect 29149 12149 29206 12157
rect 29149 12143 29157 12149
rect 28345 12139 28445 12143
rect 28345 12135 28407 12139
rect 28345 12109 28352 12135
rect 28378 12113 28407 12135
rect 28433 12113 28445 12139
rect 28378 12109 28445 12113
rect 28345 12106 28445 12109
rect 28513 12106 28548 12143
rect 28610 12140 28969 12143
rect 28610 12135 28832 12140
rect 28610 12111 28623 12135
rect 28647 12116 28832 12135
rect 28856 12116 28969 12140
rect 28647 12111 28969 12116
rect 28610 12107 28969 12111
rect 29036 12135 29157 12143
rect 29036 12115 29047 12135
rect 29067 12126 29157 12135
rect 29183 12126 29206 12149
rect 29067 12115 29206 12126
rect 29036 12113 29206 12115
rect 29509 12142 29581 12162
rect 29509 12119 29537 12142
rect 29563 12119 29581 12142
rect 29036 12108 29157 12113
rect 29036 12107 29077 12108
rect 28512 12081 28548 12106
rect 28360 12054 28397 12055
rect 28456 12054 28493 12055
rect 28512 12054 28519 12081
rect 28260 12045 28398 12054
rect 28260 12025 28369 12045
rect 28389 12025 28398 12045
rect 28260 12018 28398 12025
rect 28456 12051 28519 12054
rect 28540 12054 28548 12081
rect 28567 12054 28604 12055
rect 28540 12051 28604 12054
rect 28456 12045 28604 12051
rect 28456 12025 28465 12045
rect 28485 12025 28575 12045
rect 28595 12025 28604 12045
rect 28260 12016 28356 12018
rect 28456 12015 28604 12025
rect 28663 12045 28700 12055
rect 28775 12054 28812 12055
rect 28756 12052 28812 12054
rect 28663 12025 28671 12045
rect 28691 12025 28700 12045
rect 28512 12014 28548 12015
rect 28360 11883 28397 11884
rect 28663 11883 28700 12025
rect 28725 12045 28812 12052
rect 28725 12042 28783 12045
rect 28725 12022 28730 12042
rect 28751 12025 28783 12042
rect 28803 12025 28812 12045
rect 28751 12022 28812 12025
rect 28725 12015 28812 12022
rect 28871 12045 28908 12055
rect 28871 12025 28879 12045
rect 28899 12025 28908 12045
rect 28725 12014 28756 12015
rect 28871 11946 28908 12025
rect 28938 12054 28969 12107
rect 29509 12057 29581 12119
rect 30614 12157 30630 12183
rect 30670 12157 30694 12183
rect 30614 12138 30694 12157
rect 30614 12112 30633 12138
rect 30673 12112 30694 12138
rect 30614 12085 30694 12112
rect 30614 12059 30637 12085
rect 30677 12059 30694 12085
rect 28988 12054 29025 12055
rect 28938 12045 29025 12054
rect 28938 12025 28996 12045
rect 29016 12025 29025 12045
rect 28938 12015 29025 12025
rect 29084 12045 29121 12055
rect 29084 12025 29092 12045
rect 29112 12025 29121 12045
rect 28938 12014 28969 12015
rect 28933 11946 29043 11959
rect 29084 11946 29121 12025
rect 28871 11944 29121 11946
rect 28871 11941 28972 11944
rect 28871 11922 28936 11941
rect 28933 11914 28936 11922
rect 28965 11914 28972 11941
rect 29000 11917 29010 11944
rect 29039 11922 29121 11944
rect 29039 11917 29043 11922
rect 29000 11914 29043 11917
rect 28933 11900 29043 11914
rect 28359 11882 28700 11883
rect 28284 11877 28700 11882
rect 28284 11857 28287 11877
rect 28307 11857 28701 11877
rect 28510 11824 28547 11834
rect 28510 11787 28519 11824
rect 28536 11787 28547 11824
rect 28510 11766 28547 11787
rect 28219 10827 28387 10828
rect 28516 10827 28545 11766
rect 28658 11152 28701 11857
rect 29513 11506 29575 12057
rect 30614 12048 30694 12059
rect 30756 12049 30783 12304
rect 31161 12296 31202 12446
rect 31433 12440 31537 12446
rect 31893 12443 31957 12446
rect 31628 12384 31749 12402
rect 31628 12382 31699 12384
rect 31628 12341 31643 12382
rect 31680 12343 31699 12382
rect 31736 12343 31749 12384
rect 31680 12341 31749 12343
rect 31628 12331 31749 12341
rect 30823 12189 30887 12201
rect 31163 12197 31200 12296
rect 31428 12286 31539 12299
rect 31428 12284 31470 12286
rect 31428 12264 31435 12284
rect 31454 12264 31470 12284
rect 31428 12256 31470 12264
rect 31498 12284 31539 12286
rect 31498 12264 31512 12284
rect 31531 12264 31539 12284
rect 31498 12256 31539 12264
rect 31428 12250 31539 12256
rect 31371 12228 31620 12250
rect 31371 12197 31408 12228
rect 31584 12226 31620 12228
rect 31584 12197 31621 12226
rect 30823 12188 30858 12189
rect 30800 12183 30858 12188
rect 30800 12163 30803 12183
rect 30823 12169 30858 12183
rect 30878 12169 30887 12189
rect 30823 12161 30887 12169
rect 30849 12160 30887 12161
rect 30850 12159 30887 12160
rect 30953 12193 30989 12194
rect 31061 12193 31097 12194
rect 30953 12185 31097 12193
rect 30953 12165 30961 12185
rect 30981 12165 31069 12185
rect 31089 12165 31097 12185
rect 30953 12159 31097 12165
rect 31163 12189 31201 12197
rect 31269 12193 31305 12194
rect 31163 12169 31172 12189
rect 31192 12169 31201 12189
rect 31163 12160 31201 12169
rect 31220 12186 31305 12193
rect 31220 12166 31227 12186
rect 31248 12185 31305 12186
rect 31248 12166 31277 12185
rect 31220 12165 31277 12166
rect 31297 12165 31305 12185
rect 31163 12159 31200 12160
rect 31220 12159 31305 12165
rect 31371 12189 31409 12197
rect 31482 12193 31518 12194
rect 31371 12169 31380 12189
rect 31400 12169 31409 12189
rect 31371 12160 31409 12169
rect 31433 12185 31518 12193
rect 31433 12165 31490 12185
rect 31510 12165 31518 12185
rect 31371 12159 31408 12160
rect 31433 12159 31518 12165
rect 31584 12189 31622 12197
rect 31584 12169 31593 12189
rect 31613 12169 31622 12189
rect 31677 12179 31742 12331
rect 31895 12305 31950 12443
rect 32934 12377 32993 12448
rect 33846 12447 33898 12450
rect 33846 12412 33854 12447
rect 33879 12412 33898 12447
rect 33923 12439 33945 12450
rect 33923 12438 34790 12439
rect 33923 12412 34791 12438
rect 33846 12402 34791 12412
rect 33846 12400 33945 12402
rect 32934 12359 32956 12377
rect 32974 12359 32993 12377
rect 32934 12337 32993 12359
rect 33201 12373 33733 12378
rect 33201 12353 34087 12373
rect 34107 12353 34110 12373
rect 34746 12369 34791 12402
rect 33201 12349 34110 12353
rect 31584 12160 31622 12169
rect 31675 12172 31742 12179
rect 31584 12159 31621 12160
rect 31007 12138 31043 12159
rect 31433 12138 31464 12159
rect 31675 12151 31692 12172
rect 31728 12151 31742 12172
rect 31894 12192 31950 12305
rect 33201 12302 33244 12349
rect 33694 12348 34110 12349
rect 34742 12349 35135 12369
rect 35155 12349 35158 12369
rect 33694 12347 34035 12348
rect 33351 12316 33461 12330
rect 33351 12313 33394 12316
rect 33351 12308 33355 12313
rect 33189 12301 33244 12302
rect 31894 12174 31913 12192
rect 31931 12174 31950 12192
rect 31894 12154 31950 12174
rect 32933 12278 33244 12301
rect 32933 12260 32958 12278
rect 32976 12266 33244 12278
rect 33273 12286 33355 12308
rect 33384 12286 33394 12313
rect 33422 12289 33429 12316
rect 33458 12308 33461 12316
rect 33458 12289 33523 12308
rect 33422 12286 33523 12289
rect 33273 12284 33523 12286
rect 32976 12260 32998 12266
rect 31675 12138 31742 12151
rect 30840 12134 30940 12138
rect 30840 12130 30902 12134
rect 30840 12104 30847 12130
rect 30873 12108 30902 12130
rect 30928 12108 30940 12134
rect 30873 12104 30940 12108
rect 30840 12101 30940 12104
rect 31008 12101 31043 12138
rect 31105 12135 31464 12138
rect 31105 12130 31327 12135
rect 31105 12106 31118 12130
rect 31142 12111 31327 12130
rect 31351 12111 31464 12135
rect 31142 12106 31464 12111
rect 31105 12102 31464 12106
rect 31531 12132 31742 12138
rect 31531 12130 31692 12132
rect 31531 12110 31542 12130
rect 31562 12110 31692 12130
rect 31531 12103 31692 12110
rect 31531 12102 31572 12103
rect 31007 12076 31043 12101
rect 30855 12049 30892 12050
rect 30951 12049 30988 12050
rect 31007 12049 31014 12076
rect 30755 12040 30893 12049
rect 30755 12020 30864 12040
rect 30884 12020 30893 12040
rect 30755 12013 30893 12020
rect 30951 12046 31014 12049
rect 31035 12049 31043 12076
rect 31062 12049 31099 12050
rect 31035 12046 31099 12049
rect 30951 12040 31099 12046
rect 30951 12020 30960 12040
rect 30980 12020 31070 12040
rect 31090 12020 31099 12040
rect 30755 12011 30851 12013
rect 30951 12010 31099 12020
rect 31158 12040 31195 12050
rect 31270 12049 31307 12050
rect 31251 12047 31307 12049
rect 31158 12020 31166 12040
rect 31186 12020 31195 12040
rect 31007 12009 31043 12010
rect 30855 11878 30892 11879
rect 31158 11878 31195 12020
rect 31220 12040 31307 12047
rect 31220 12037 31278 12040
rect 31220 12017 31225 12037
rect 31246 12020 31278 12037
rect 31298 12020 31307 12040
rect 31246 12017 31307 12020
rect 31220 12010 31307 12017
rect 31366 12040 31403 12050
rect 31366 12020 31374 12040
rect 31394 12020 31403 12040
rect 31220 12009 31251 12010
rect 31366 11941 31403 12020
rect 31433 12049 31464 12102
rect 31677 12095 31692 12103
rect 31732 12095 31742 12132
rect 32933 12121 32998 12260
rect 33273 12205 33310 12284
rect 33351 12271 33461 12284
rect 33425 12215 33456 12216
rect 33273 12185 33282 12205
rect 33302 12185 33310 12205
rect 31677 12086 31742 12095
rect 31890 12093 31955 12114
rect 31890 12075 31915 12093
rect 31933 12075 31955 12093
rect 32933 12103 32956 12121
rect 32974 12103 32998 12121
rect 32933 12086 32998 12103
rect 33153 12167 33221 12180
rect 33273 12175 33310 12185
rect 33369 12205 33456 12215
rect 33369 12185 33378 12205
rect 33398 12185 33456 12205
rect 33369 12176 33456 12185
rect 33369 12175 33406 12176
rect 33153 12125 33160 12167
rect 33209 12125 33221 12167
rect 33153 12122 33221 12125
rect 33425 12123 33456 12176
rect 33486 12205 33523 12284
rect 33638 12215 33669 12216
rect 33486 12185 33495 12205
rect 33515 12185 33523 12205
rect 33486 12175 33523 12185
rect 33582 12208 33669 12215
rect 33582 12205 33643 12208
rect 33582 12185 33591 12205
rect 33611 12188 33643 12205
rect 33664 12188 33669 12208
rect 33611 12185 33669 12188
rect 33582 12178 33669 12185
rect 33694 12205 33731 12347
rect 33997 12346 34034 12347
rect 34742 12344 35158 12349
rect 34742 12343 35083 12344
rect 34399 12312 34509 12326
rect 34399 12309 34442 12312
rect 34399 12304 34403 12309
rect 34321 12282 34403 12304
rect 34432 12282 34442 12309
rect 34470 12285 34477 12312
rect 34506 12304 34509 12312
rect 34506 12285 34571 12304
rect 34470 12282 34571 12285
rect 34321 12280 34571 12282
rect 33846 12215 33882 12216
rect 33694 12185 33703 12205
rect 33723 12185 33731 12205
rect 33582 12176 33638 12178
rect 33582 12175 33619 12176
rect 33694 12175 33731 12185
rect 33790 12205 33938 12215
rect 34038 12212 34134 12214
rect 33790 12185 33799 12205
rect 33819 12185 33909 12205
rect 33929 12185 33938 12205
rect 33790 12179 33938 12185
rect 33790 12176 33854 12179
rect 33790 12175 33827 12176
rect 33846 12149 33854 12176
rect 33875 12176 33938 12179
rect 33996 12205 34134 12212
rect 33996 12185 34005 12205
rect 34025 12185 34134 12205
rect 33996 12176 34134 12185
rect 34321 12201 34358 12280
rect 34399 12267 34509 12280
rect 34473 12211 34504 12212
rect 34321 12181 34330 12201
rect 34350 12181 34358 12201
rect 33875 12149 33882 12176
rect 33901 12175 33938 12176
rect 33997 12175 34034 12176
rect 33846 12124 33882 12149
rect 33317 12122 33358 12123
rect 33153 12115 33358 12122
rect 33153 12104 33327 12115
rect 31483 12049 31520 12050
rect 31433 12040 31520 12049
rect 31433 12020 31491 12040
rect 31511 12020 31520 12040
rect 31433 12010 31520 12020
rect 31579 12040 31616 12050
rect 31579 12020 31587 12040
rect 31607 12020 31616 12040
rect 31433 12009 31464 12010
rect 31428 11941 31538 11954
rect 31579 11941 31616 12020
rect 31890 11999 31955 12075
rect 33153 12071 33161 12104
rect 33154 12062 33161 12071
rect 33210 12095 33327 12104
rect 33347 12095 33358 12115
rect 33210 12087 33358 12095
rect 33425 12119 33784 12123
rect 33425 12114 33747 12119
rect 33425 12090 33538 12114
rect 33562 12095 33747 12114
rect 33771 12095 33784 12119
rect 33562 12090 33784 12095
rect 33425 12087 33784 12090
rect 33846 12087 33881 12124
rect 33949 12121 34049 12124
rect 33949 12117 34016 12121
rect 33949 12091 33961 12117
rect 33987 12095 34016 12117
rect 34042 12095 34049 12121
rect 33987 12091 34049 12095
rect 33949 12087 34049 12091
rect 33210 12071 33221 12087
rect 33210 12062 33218 12071
rect 33425 12066 33456 12087
rect 33846 12066 33882 12087
rect 33268 12065 33305 12066
rect 32933 12022 32998 12041
rect 32933 12004 32958 12022
rect 32976 12004 32998 12022
rect 31366 11939 31616 11941
rect 31366 11936 31467 11939
rect 31366 11917 31431 11936
rect 31428 11909 31431 11917
rect 31460 11909 31467 11936
rect 31495 11912 31505 11939
rect 31534 11917 31616 11939
rect 31639 11964 31956 11999
rect 31534 11912 31538 11917
rect 31495 11909 31538 11912
rect 31428 11895 31538 11909
rect 30854 11877 31195 11878
rect 30779 11875 31195 11877
rect 31639 11875 31679 11964
rect 31890 11937 31955 11964
rect 31890 11919 31913 11937
rect 31931 11919 31955 11937
rect 31890 11899 31955 11919
rect 30776 11872 31679 11875
rect 30776 11852 30782 11872
rect 30802 11852 31679 11872
rect 30776 11848 31679 11852
rect 31639 11845 31679 11848
rect 31891 11838 31956 11859
rect 30109 11830 30770 11831
rect 30109 11823 31043 11830
rect 30109 11822 31015 11823
rect 30109 11802 30960 11822
rect 30992 11803 31015 11822
rect 31040 11803 31043 11823
rect 30992 11802 31043 11803
rect 30109 11795 31043 11802
rect 29708 11753 29876 11754
rect 30111 11753 30150 11795
rect 30939 11793 31043 11795
rect 31008 11791 31043 11793
rect 31891 11820 31915 11838
rect 31933 11820 31956 11838
rect 31891 11773 31956 11820
rect 29708 11727 30152 11753
rect 29708 11725 29876 11727
rect 29510 11422 29579 11506
rect 28659 11144 28701 11152
rect 28659 11133 28704 11144
rect 28659 11095 28669 11133
rect 28694 11095 28704 11133
rect 28659 11086 28704 11095
rect 29508 10943 29579 11422
rect 29708 11374 29735 11725
rect 30111 11721 30152 11727
rect 29775 11514 29839 11526
rect 30115 11522 30152 11721
rect 30614 11748 30686 11765
rect 30614 11709 30622 11748
rect 30667 11709 30686 11748
rect 30380 11611 30491 11626
rect 30380 11609 30422 11611
rect 30380 11589 30387 11609
rect 30406 11589 30422 11609
rect 30380 11581 30422 11589
rect 30450 11609 30491 11611
rect 30450 11589 30464 11609
rect 30483 11589 30491 11609
rect 30450 11581 30491 11589
rect 30380 11575 30491 11581
rect 30323 11553 30572 11575
rect 30323 11522 30360 11553
rect 30536 11551 30572 11553
rect 30536 11522 30573 11551
rect 29775 11513 29810 11514
rect 29752 11508 29810 11513
rect 29752 11488 29755 11508
rect 29775 11494 29810 11508
rect 29830 11494 29839 11514
rect 29775 11486 29839 11494
rect 29801 11485 29839 11486
rect 29802 11484 29839 11485
rect 29905 11518 29941 11519
rect 30013 11518 30049 11519
rect 29905 11510 30049 11518
rect 29905 11490 29913 11510
rect 29933 11490 30021 11510
rect 30041 11490 30049 11510
rect 29905 11484 30049 11490
rect 30115 11514 30153 11522
rect 30221 11518 30257 11519
rect 30115 11494 30124 11514
rect 30144 11494 30153 11514
rect 30115 11485 30153 11494
rect 30172 11511 30257 11518
rect 30172 11491 30179 11511
rect 30200 11510 30257 11511
rect 30200 11491 30229 11510
rect 30172 11490 30229 11491
rect 30249 11490 30257 11510
rect 30115 11484 30152 11485
rect 30172 11484 30257 11490
rect 30323 11514 30361 11522
rect 30434 11518 30470 11519
rect 30323 11494 30332 11514
rect 30352 11494 30361 11514
rect 30323 11485 30361 11494
rect 30385 11510 30470 11518
rect 30385 11490 30442 11510
rect 30462 11490 30470 11510
rect 30323 11484 30360 11485
rect 30385 11484 30470 11490
rect 30536 11514 30574 11522
rect 30536 11494 30545 11514
rect 30565 11494 30574 11514
rect 30536 11485 30574 11494
rect 30614 11499 30686 11709
rect 30756 11743 31956 11773
rect 30756 11742 31200 11743
rect 30756 11740 30924 11742
rect 30614 11485 30697 11499
rect 30536 11484 30573 11485
rect 29959 11463 29995 11484
rect 30385 11463 30416 11484
rect 30614 11463 30631 11485
rect 29792 11459 29892 11463
rect 29792 11455 29854 11459
rect 29792 11429 29799 11455
rect 29825 11433 29854 11455
rect 29880 11433 29892 11459
rect 29825 11429 29892 11433
rect 29792 11426 29892 11429
rect 29960 11426 29995 11463
rect 30057 11460 30416 11463
rect 30057 11455 30279 11460
rect 30057 11431 30070 11455
rect 30094 11436 30279 11455
rect 30303 11436 30416 11460
rect 30094 11431 30416 11436
rect 30057 11427 30416 11431
rect 30483 11455 30631 11463
rect 30483 11435 30494 11455
rect 30514 11452 30631 11455
rect 30684 11452 30697 11485
rect 30514 11435 30697 11452
rect 30483 11428 30697 11435
rect 30483 11427 30524 11428
rect 30614 11427 30697 11428
rect 29959 11401 29995 11426
rect 29807 11374 29844 11375
rect 29903 11374 29940 11375
rect 29959 11374 29966 11401
rect 29707 11365 29845 11374
rect 29707 11345 29816 11365
rect 29836 11345 29845 11365
rect 29707 11338 29845 11345
rect 29903 11371 29966 11374
rect 29987 11374 29995 11401
rect 30014 11374 30051 11375
rect 29987 11371 30051 11374
rect 29903 11365 30051 11371
rect 29903 11345 29912 11365
rect 29932 11345 30022 11365
rect 30042 11345 30051 11365
rect 29707 11336 29803 11338
rect 29903 11335 30051 11345
rect 30110 11365 30147 11375
rect 30222 11374 30259 11375
rect 30203 11372 30259 11374
rect 30110 11345 30118 11365
rect 30138 11345 30147 11365
rect 29959 11334 29995 11335
rect 29807 11203 29844 11204
rect 30110 11203 30147 11345
rect 30172 11365 30259 11372
rect 30172 11362 30230 11365
rect 30172 11342 30177 11362
rect 30198 11345 30230 11362
rect 30250 11345 30259 11365
rect 30198 11342 30259 11345
rect 30172 11335 30259 11342
rect 30318 11365 30355 11375
rect 30318 11345 30326 11365
rect 30346 11345 30355 11365
rect 30172 11334 30203 11335
rect 30318 11266 30355 11345
rect 30385 11374 30416 11427
rect 30622 11394 30636 11427
rect 30689 11394 30697 11427
rect 30622 11388 30697 11394
rect 30622 11383 30692 11388
rect 30435 11374 30472 11375
rect 30385 11365 30472 11374
rect 30385 11345 30443 11365
rect 30463 11345 30472 11365
rect 30385 11335 30472 11345
rect 30531 11365 30568 11375
rect 30756 11370 30783 11740
rect 30823 11510 30887 11522
rect 31163 11518 31200 11742
rect 31671 11723 31735 11725
rect 31667 11711 31735 11723
rect 31667 11678 31678 11711
rect 31718 11678 31735 11711
rect 31667 11668 31735 11678
rect 31428 11607 31539 11622
rect 31428 11605 31470 11607
rect 31428 11585 31435 11605
rect 31454 11585 31470 11605
rect 31428 11577 31470 11585
rect 31498 11605 31539 11607
rect 31498 11585 31512 11605
rect 31531 11585 31539 11605
rect 31498 11577 31539 11585
rect 31428 11571 31539 11577
rect 31371 11549 31620 11571
rect 31371 11518 31408 11549
rect 31584 11547 31620 11549
rect 31584 11518 31621 11547
rect 30823 11509 30858 11510
rect 30800 11504 30858 11509
rect 30800 11484 30803 11504
rect 30823 11490 30858 11504
rect 30878 11490 30887 11510
rect 30823 11482 30887 11490
rect 30849 11481 30887 11482
rect 30850 11480 30887 11481
rect 30953 11514 30989 11515
rect 31061 11514 31097 11515
rect 30953 11506 31097 11514
rect 30953 11486 30961 11506
rect 30981 11486 31069 11506
rect 31089 11486 31097 11506
rect 30953 11480 31097 11486
rect 31163 11510 31201 11518
rect 31269 11514 31305 11515
rect 31163 11490 31172 11510
rect 31192 11490 31201 11510
rect 31163 11481 31201 11490
rect 31220 11507 31305 11514
rect 31220 11487 31227 11507
rect 31248 11506 31305 11507
rect 31248 11487 31277 11506
rect 31220 11486 31277 11487
rect 31297 11486 31305 11506
rect 31163 11480 31200 11481
rect 31220 11480 31305 11486
rect 31371 11510 31409 11518
rect 31482 11514 31518 11515
rect 31371 11490 31380 11510
rect 31400 11490 31409 11510
rect 31371 11481 31409 11490
rect 31433 11506 31518 11514
rect 31433 11486 31490 11506
rect 31510 11486 31518 11506
rect 31371 11480 31408 11481
rect 31433 11480 31518 11486
rect 31584 11510 31622 11518
rect 31584 11490 31593 11510
rect 31613 11490 31622 11510
rect 31584 11481 31622 11490
rect 31671 11484 31735 11668
rect 31891 11542 31956 11743
rect 32933 11803 32998 12004
rect 33154 11878 33218 12062
rect 33267 12056 33305 12065
rect 33267 12036 33276 12056
rect 33296 12036 33305 12056
rect 33267 12028 33305 12036
rect 33371 12060 33456 12066
rect 33481 12065 33518 12066
rect 33371 12040 33379 12060
rect 33399 12040 33456 12060
rect 33371 12032 33456 12040
rect 33480 12056 33518 12065
rect 33480 12036 33489 12056
rect 33509 12036 33518 12056
rect 33371 12031 33407 12032
rect 33480 12028 33518 12036
rect 33584 12060 33669 12066
rect 33689 12065 33726 12066
rect 33584 12040 33592 12060
rect 33612 12059 33669 12060
rect 33612 12040 33641 12059
rect 33584 12039 33641 12040
rect 33662 12039 33669 12059
rect 33584 12032 33669 12039
rect 33688 12056 33726 12065
rect 33688 12036 33697 12056
rect 33717 12036 33726 12056
rect 33584 12031 33620 12032
rect 33688 12028 33726 12036
rect 33792 12060 33936 12066
rect 33792 12040 33800 12060
rect 33820 12040 33908 12060
rect 33928 12040 33936 12060
rect 33792 12032 33936 12040
rect 33792 12031 33828 12032
rect 33900 12031 33936 12032
rect 34002 12065 34039 12066
rect 34002 12064 34040 12065
rect 34002 12056 34066 12064
rect 34002 12036 34011 12056
rect 34031 12042 34066 12056
rect 34086 12042 34089 12062
rect 34031 12037 34089 12042
rect 34031 12036 34066 12037
rect 33268 11999 33305 12028
rect 33269 11997 33305 11999
rect 33481 11997 33518 12028
rect 33269 11975 33518 11997
rect 33350 11969 33461 11975
rect 33350 11961 33391 11969
rect 33350 11941 33358 11961
rect 33377 11941 33391 11961
rect 33350 11939 33391 11941
rect 33419 11961 33461 11969
rect 33419 11941 33435 11961
rect 33454 11941 33461 11961
rect 33419 11939 33461 11941
rect 33350 11924 33461 11939
rect 33154 11868 33222 11878
rect 33154 11835 33171 11868
rect 33211 11835 33222 11868
rect 33154 11823 33222 11835
rect 33154 11821 33218 11823
rect 33689 11804 33726 12028
rect 34002 12024 34066 12036
rect 34106 11806 34133 12176
rect 34321 12171 34358 12181
rect 34417 12201 34504 12211
rect 34417 12181 34426 12201
rect 34446 12181 34504 12201
rect 34417 12172 34504 12181
rect 34417 12171 34454 12172
rect 34197 12158 34267 12163
rect 34192 12152 34267 12158
rect 34192 12119 34200 12152
rect 34253 12119 34267 12152
rect 34473 12119 34504 12172
rect 34534 12201 34571 12280
rect 34686 12211 34717 12212
rect 34534 12181 34543 12201
rect 34563 12181 34571 12201
rect 34534 12171 34571 12181
rect 34630 12204 34717 12211
rect 34630 12201 34691 12204
rect 34630 12181 34639 12201
rect 34659 12184 34691 12201
rect 34712 12184 34717 12204
rect 34659 12181 34717 12184
rect 34630 12174 34717 12181
rect 34742 12201 34779 12343
rect 35045 12342 35082 12343
rect 34894 12211 34930 12212
rect 34742 12181 34751 12201
rect 34771 12181 34779 12201
rect 34630 12172 34686 12174
rect 34630 12171 34667 12172
rect 34742 12171 34779 12181
rect 34838 12201 34986 12211
rect 35086 12208 35182 12210
rect 34838 12181 34847 12201
rect 34867 12181 34957 12201
rect 34977 12181 34986 12201
rect 34838 12175 34986 12181
rect 34838 12172 34902 12175
rect 34838 12171 34875 12172
rect 34894 12145 34902 12172
rect 34923 12172 34986 12175
rect 35044 12201 35182 12208
rect 35044 12181 35053 12201
rect 35073 12181 35182 12201
rect 35044 12172 35182 12181
rect 34923 12145 34930 12172
rect 34949 12171 34986 12172
rect 35045 12171 35082 12172
rect 34894 12120 34930 12145
rect 34192 12118 34275 12119
rect 34365 12118 34406 12119
rect 34192 12111 34406 12118
rect 34192 12094 34375 12111
rect 34192 12061 34205 12094
rect 34258 12091 34375 12094
rect 34395 12091 34406 12111
rect 34258 12083 34406 12091
rect 34473 12115 34832 12119
rect 34473 12110 34795 12115
rect 34473 12086 34586 12110
rect 34610 12091 34795 12110
rect 34819 12091 34832 12115
rect 34610 12086 34832 12091
rect 34473 12083 34832 12086
rect 34894 12083 34929 12120
rect 34997 12117 35097 12120
rect 34997 12113 35064 12117
rect 34997 12087 35009 12113
rect 35035 12091 35064 12113
rect 35090 12091 35097 12117
rect 35035 12087 35097 12091
rect 34997 12083 35097 12087
rect 34258 12061 34275 12083
rect 34473 12062 34504 12083
rect 34894 12062 34930 12083
rect 34316 12061 34353 12062
rect 34192 12047 34275 12061
rect 33965 11804 34133 11806
rect 33689 11803 34133 11804
rect 32933 11773 34133 11803
rect 34203 11837 34275 12047
rect 34315 12052 34353 12061
rect 34315 12032 34324 12052
rect 34344 12032 34353 12052
rect 34315 12024 34353 12032
rect 34419 12056 34504 12062
rect 34529 12061 34566 12062
rect 34419 12036 34427 12056
rect 34447 12036 34504 12056
rect 34419 12028 34504 12036
rect 34528 12052 34566 12061
rect 34528 12032 34537 12052
rect 34557 12032 34566 12052
rect 34419 12027 34455 12028
rect 34528 12024 34566 12032
rect 34632 12056 34717 12062
rect 34737 12061 34774 12062
rect 34632 12036 34640 12056
rect 34660 12055 34717 12056
rect 34660 12036 34689 12055
rect 34632 12035 34689 12036
rect 34710 12035 34717 12055
rect 34632 12028 34717 12035
rect 34736 12052 34774 12061
rect 34736 12032 34745 12052
rect 34765 12032 34774 12052
rect 34632 12027 34668 12028
rect 34736 12024 34774 12032
rect 34840 12056 34984 12062
rect 34840 12036 34848 12056
rect 34868 12036 34956 12056
rect 34976 12036 34984 12056
rect 34840 12028 34984 12036
rect 34840 12027 34876 12028
rect 34948 12027 34984 12028
rect 35050 12061 35087 12062
rect 35050 12060 35088 12061
rect 35050 12052 35114 12060
rect 35050 12032 35059 12052
rect 35079 12038 35114 12052
rect 35134 12038 35137 12058
rect 35079 12033 35137 12038
rect 35079 12032 35114 12033
rect 34316 11995 34353 12024
rect 34317 11993 34353 11995
rect 34529 11993 34566 12024
rect 34317 11971 34566 11993
rect 34398 11965 34509 11971
rect 34398 11957 34439 11965
rect 34398 11937 34406 11957
rect 34425 11937 34439 11957
rect 34398 11935 34439 11937
rect 34467 11957 34509 11965
rect 34467 11937 34483 11957
rect 34502 11937 34509 11957
rect 34467 11935 34509 11937
rect 34398 11920 34509 11935
rect 34203 11798 34222 11837
rect 34267 11798 34275 11837
rect 34203 11781 34275 11798
rect 34737 11825 34774 12024
rect 35050 12020 35114 12032
rect 34737 11819 34778 11825
rect 35154 11821 35181 12172
rect 35304 12042 35383 12642
rect 35480 12190 35559 12775
rect 35763 12762 35800 12791
rect 35764 12760 35800 12762
rect 35976 12760 36013 12791
rect 35764 12738 36013 12760
rect 35845 12732 35956 12738
rect 35845 12724 35886 12732
rect 35845 12704 35853 12724
rect 35872 12704 35886 12724
rect 35845 12702 35886 12704
rect 35914 12724 35956 12732
rect 35914 12704 35930 12724
rect 35949 12704 35956 12724
rect 35914 12702 35956 12704
rect 35845 12687 35956 12702
rect 36184 12676 36221 12791
rect 36177 12564 36224 12676
rect 36345 12636 36375 12795
rect 36395 12794 36431 12795
rect 36497 12828 36534 12829
rect 36497 12827 36535 12828
rect 36497 12819 36561 12827
rect 36497 12799 36506 12819
rect 36526 12805 36561 12819
rect 36581 12805 36584 12825
rect 36526 12800 36584 12805
rect 36526 12799 36561 12800
rect 36497 12787 36561 12799
rect 36345 12632 36431 12636
rect 36345 12614 36360 12632
rect 36412 12614 36431 12632
rect 36345 12605 36431 12614
rect 36601 12566 36628 12939
rect 36460 12564 36628 12566
rect 36177 12538 36628 12564
rect 36177 12460 36224 12538
rect 36460 12537 36628 12538
rect 36122 12459 36224 12460
rect 36121 12451 36224 12459
rect 36121 12448 36173 12451
rect 36121 12413 36129 12448
rect 36154 12413 36173 12448
rect 36198 12413 36224 12451
rect 36121 12407 36224 12413
rect 36384 12452 36420 12456
rect 36384 12429 36392 12452
rect 36416 12429 36420 12452
rect 36384 12408 36420 12429
rect 36121 12403 36220 12407
rect 36384 12385 36392 12408
rect 36416 12385 36420 12408
rect 35013 11819 35181 11821
rect 34737 11793 35181 11819
rect 32933 11726 32998 11773
rect 32933 11708 32956 11726
rect 32974 11708 32998 11726
rect 33846 11753 33881 11755
rect 33846 11751 33950 11753
rect 34739 11751 34778 11793
rect 35013 11792 35181 11793
rect 33846 11744 34780 11751
rect 33846 11743 33897 11744
rect 33846 11723 33849 11743
rect 33874 11724 33897 11743
rect 33929 11724 34780 11744
rect 33874 11723 34780 11724
rect 33846 11716 34780 11723
rect 34119 11715 34780 11716
rect 32933 11687 32998 11708
rect 33210 11698 33250 11701
rect 33210 11694 34113 11698
rect 33210 11674 34087 11694
rect 34107 11674 34113 11694
rect 33210 11671 34113 11674
rect 32934 11627 32999 11647
rect 32934 11609 32958 11627
rect 32976 11609 32999 11627
rect 32934 11582 32999 11609
rect 33210 11582 33250 11671
rect 33694 11669 34110 11671
rect 33694 11668 34035 11669
rect 33351 11637 33461 11651
rect 33351 11634 33394 11637
rect 33351 11629 33355 11634
rect 32933 11547 33250 11582
rect 33273 11607 33355 11629
rect 33384 11607 33394 11634
rect 33422 11610 33429 11637
rect 33458 11629 33461 11637
rect 33458 11610 33523 11629
rect 33422 11607 33523 11610
rect 33273 11605 33523 11607
rect 31891 11524 31913 11542
rect 31931 11524 31956 11542
rect 31891 11505 31956 11524
rect 31584 11480 31621 11481
rect 31007 11459 31043 11480
rect 31433 11459 31464 11480
rect 31671 11475 31679 11484
rect 31668 11459 31679 11475
rect 30840 11455 30940 11459
rect 30840 11451 30902 11455
rect 30840 11425 30847 11451
rect 30873 11429 30902 11451
rect 30928 11429 30940 11455
rect 30873 11425 30940 11429
rect 30840 11422 30940 11425
rect 31008 11422 31043 11459
rect 31105 11456 31464 11459
rect 31105 11451 31327 11456
rect 31105 11427 31118 11451
rect 31142 11432 31327 11451
rect 31351 11432 31464 11456
rect 31142 11427 31464 11432
rect 31105 11423 31464 11427
rect 31531 11451 31679 11459
rect 31531 11431 31542 11451
rect 31562 11442 31679 11451
rect 31728 11475 31735 11484
rect 31728 11442 31736 11475
rect 32934 11471 32999 11547
rect 33273 11526 33310 11605
rect 33351 11592 33461 11605
rect 33425 11536 33456 11537
rect 33273 11506 33282 11526
rect 33302 11506 33310 11526
rect 33273 11496 33310 11506
rect 33369 11526 33456 11536
rect 33369 11506 33378 11526
rect 33398 11506 33456 11526
rect 33369 11497 33456 11506
rect 33369 11496 33406 11497
rect 31562 11431 31736 11442
rect 31531 11424 31736 11431
rect 31531 11423 31572 11424
rect 31007 11397 31043 11422
rect 30855 11370 30892 11371
rect 30951 11370 30988 11371
rect 31007 11370 31014 11397
rect 30531 11345 30539 11365
rect 30559 11345 30568 11365
rect 30385 11334 30416 11335
rect 30380 11266 30490 11279
rect 30531 11266 30568 11345
rect 30755 11361 30893 11370
rect 30755 11341 30864 11361
rect 30884 11341 30893 11361
rect 30755 11334 30893 11341
rect 30951 11367 31014 11370
rect 31035 11370 31043 11397
rect 31062 11370 31099 11371
rect 31035 11367 31099 11370
rect 30951 11361 31099 11367
rect 30951 11341 30960 11361
rect 30980 11341 31070 11361
rect 31090 11341 31099 11361
rect 30755 11332 30851 11334
rect 30951 11331 31099 11341
rect 31158 11361 31195 11371
rect 31270 11370 31307 11371
rect 31251 11368 31307 11370
rect 31158 11341 31166 11361
rect 31186 11341 31195 11361
rect 31007 11330 31043 11331
rect 30318 11264 30568 11266
rect 30318 11261 30419 11264
rect 30318 11242 30383 11261
rect 30380 11234 30383 11242
rect 30412 11234 30419 11261
rect 30447 11237 30457 11264
rect 30486 11242 30568 11264
rect 30486 11237 30490 11242
rect 30447 11234 30490 11237
rect 30380 11220 30490 11234
rect 29806 11202 30147 11203
rect 29731 11197 30147 11202
rect 30855 11199 30892 11200
rect 31158 11199 31195 11341
rect 31220 11361 31307 11368
rect 31220 11358 31278 11361
rect 31220 11338 31225 11358
rect 31246 11341 31278 11358
rect 31298 11341 31307 11361
rect 31246 11338 31307 11341
rect 31220 11331 31307 11338
rect 31366 11361 31403 11371
rect 31366 11341 31374 11361
rect 31394 11341 31403 11361
rect 31220 11330 31251 11331
rect 31366 11262 31403 11341
rect 31433 11370 31464 11423
rect 31668 11421 31736 11424
rect 31668 11379 31680 11421
rect 31729 11379 31736 11421
rect 31483 11370 31520 11371
rect 31433 11361 31520 11370
rect 31433 11341 31491 11361
rect 31511 11341 31520 11361
rect 31433 11331 31520 11341
rect 31579 11361 31616 11371
rect 31668 11366 31736 11379
rect 31891 11443 31956 11460
rect 31891 11425 31915 11443
rect 31933 11425 31956 11443
rect 32934 11453 32956 11471
rect 32974 11453 32999 11471
rect 32934 11432 32999 11453
rect 33147 11451 33212 11460
rect 31579 11341 31587 11361
rect 31607 11341 31616 11361
rect 31433 11330 31464 11331
rect 31428 11262 31538 11275
rect 31579 11262 31616 11341
rect 31891 11286 31956 11425
rect 33147 11414 33157 11451
rect 33197 11443 33212 11451
rect 33425 11444 33456 11497
rect 33486 11526 33523 11605
rect 33638 11536 33669 11537
rect 33486 11506 33495 11526
rect 33515 11506 33523 11526
rect 33486 11496 33523 11506
rect 33582 11529 33669 11536
rect 33582 11526 33643 11529
rect 33582 11506 33591 11526
rect 33611 11509 33643 11526
rect 33664 11509 33669 11529
rect 33611 11506 33669 11509
rect 33582 11499 33669 11506
rect 33694 11526 33731 11668
rect 33997 11667 34034 11668
rect 33846 11536 33882 11537
rect 33694 11506 33703 11526
rect 33723 11506 33731 11526
rect 33582 11497 33638 11499
rect 33582 11496 33619 11497
rect 33694 11496 33731 11506
rect 33790 11526 33938 11536
rect 34038 11533 34134 11535
rect 33790 11506 33799 11526
rect 33819 11506 33909 11526
rect 33929 11506 33938 11526
rect 33790 11500 33938 11506
rect 33790 11497 33854 11500
rect 33790 11496 33827 11497
rect 33846 11470 33854 11497
rect 33875 11497 33938 11500
rect 33996 11526 34134 11533
rect 33996 11506 34005 11526
rect 34025 11506 34134 11526
rect 33996 11497 34134 11506
rect 33875 11470 33882 11497
rect 33901 11496 33938 11497
rect 33997 11496 34034 11497
rect 33846 11445 33882 11470
rect 33317 11443 33358 11444
rect 33197 11436 33358 11443
rect 33197 11416 33327 11436
rect 33347 11416 33358 11436
rect 33197 11414 33358 11416
rect 33147 11408 33358 11414
rect 33425 11440 33784 11444
rect 33425 11435 33747 11440
rect 33425 11411 33538 11435
rect 33562 11416 33747 11435
rect 33771 11416 33784 11440
rect 33562 11411 33784 11416
rect 33425 11408 33784 11411
rect 33846 11408 33881 11445
rect 33949 11442 34049 11445
rect 33949 11438 34016 11442
rect 33949 11412 33961 11438
rect 33987 11416 34016 11438
rect 34042 11416 34049 11442
rect 33987 11412 34049 11416
rect 33949 11408 34049 11412
rect 33147 11395 33214 11408
rect 31891 11280 31913 11286
rect 31366 11260 31616 11262
rect 31366 11257 31467 11260
rect 31366 11238 31431 11257
rect 31428 11230 31431 11238
rect 31460 11230 31467 11257
rect 31495 11233 31505 11260
rect 31534 11238 31616 11260
rect 31645 11268 31913 11280
rect 31931 11268 31956 11286
rect 31645 11245 31956 11268
rect 32939 11372 32995 11392
rect 32939 11354 32958 11372
rect 32976 11354 32995 11372
rect 31645 11244 31700 11245
rect 31534 11233 31538 11238
rect 31495 11230 31538 11233
rect 31428 11216 31538 11230
rect 30854 11198 31195 11199
rect 29731 11177 29734 11197
rect 29754 11177 30147 11197
rect 30779 11197 31195 11198
rect 31645 11197 31688 11244
rect 32939 11241 32995 11354
rect 33147 11374 33161 11395
rect 33197 11374 33214 11395
rect 33425 11387 33456 11408
rect 33846 11387 33882 11408
rect 33268 11386 33305 11387
rect 33147 11367 33214 11374
rect 33267 11377 33305 11386
rect 30779 11193 31688 11197
rect 30098 11144 30143 11177
rect 30779 11173 30782 11193
rect 30802 11173 31688 11193
rect 31156 11168 31688 11173
rect 31896 11187 31955 11209
rect 31896 11169 31915 11187
rect 31933 11169 31955 11187
rect 30944 11144 31043 11146
rect 30098 11134 31043 11144
rect 30098 11108 30966 11134
rect 30099 11107 30966 11108
rect 30944 11096 30966 11107
rect 30991 11099 31010 11134
rect 31035 11099 31043 11134
rect 30991 11096 31043 11099
rect 30944 11088 31043 11096
rect 30970 11087 31042 11088
rect 31896 11039 31955 11169
rect 32939 11112 32994 11241
rect 33147 11215 33212 11367
rect 33267 11357 33276 11377
rect 33296 11357 33305 11377
rect 33267 11349 33305 11357
rect 33371 11381 33456 11387
rect 33481 11386 33518 11387
rect 33371 11361 33379 11381
rect 33399 11361 33456 11381
rect 33371 11353 33456 11361
rect 33480 11377 33518 11386
rect 33480 11357 33489 11377
rect 33509 11357 33518 11377
rect 33371 11352 33407 11353
rect 33480 11349 33518 11357
rect 33584 11381 33669 11387
rect 33689 11386 33726 11387
rect 33584 11361 33592 11381
rect 33612 11380 33669 11381
rect 33612 11361 33641 11380
rect 33584 11360 33641 11361
rect 33662 11360 33669 11380
rect 33584 11353 33669 11360
rect 33688 11377 33726 11386
rect 33688 11357 33697 11377
rect 33717 11357 33726 11377
rect 33584 11352 33620 11353
rect 33688 11349 33726 11357
rect 33792 11381 33936 11387
rect 33792 11361 33800 11381
rect 33820 11361 33908 11381
rect 33928 11361 33936 11381
rect 33792 11353 33936 11361
rect 33792 11352 33828 11353
rect 33900 11352 33936 11353
rect 34002 11386 34039 11387
rect 34002 11385 34040 11386
rect 34002 11377 34066 11385
rect 34002 11357 34011 11377
rect 34031 11363 34066 11377
rect 34086 11363 34089 11383
rect 34031 11358 34089 11363
rect 34031 11357 34066 11358
rect 33268 11320 33305 11349
rect 33269 11318 33305 11320
rect 33481 11318 33518 11349
rect 33269 11296 33518 11318
rect 33350 11290 33461 11296
rect 33350 11282 33391 11290
rect 33350 11262 33358 11282
rect 33377 11262 33391 11282
rect 33350 11260 33391 11262
rect 33419 11282 33461 11290
rect 33419 11262 33435 11282
rect 33454 11262 33461 11282
rect 33419 11260 33461 11262
rect 33350 11245 33461 11260
rect 33689 11250 33726 11349
rect 34002 11345 34066 11357
rect 33352 11236 33456 11245
rect 33140 11205 33261 11215
rect 33140 11203 33209 11205
rect 33140 11162 33153 11203
rect 33190 11164 33209 11203
rect 33246 11164 33261 11205
rect 33190 11162 33261 11164
rect 33140 11144 33261 11162
rect 32933 11100 32994 11112
rect 33687 11100 33728 11250
rect 34106 11242 34133 11497
rect 34195 11487 34275 11498
rect 34195 11461 34212 11487
rect 34252 11461 34275 11487
rect 34195 11434 34275 11461
rect 34195 11408 34216 11434
rect 34256 11408 34275 11434
rect 34195 11389 34275 11408
rect 34195 11363 34219 11389
rect 34259 11363 34275 11389
rect 34195 11312 34275 11363
rect 32933 11097 33728 11100
rect 34107 11111 34133 11242
rect 34197 11156 34267 11312
rect 34196 11140 34272 11156
rect 34107 11097 34135 11111
rect 32933 11062 34135 11097
rect 34196 11103 34211 11140
rect 34255 11103 34272 11140
rect 34196 11083 34272 11103
rect 35310 11133 35380 12042
rect 35479 11477 35560 12190
rect 36384 12076 36420 12385
rect 36308 12047 36421 12076
rect 36308 11691 36339 12047
rect 36378 11792 37369 11817
rect 36378 11787 36438 11792
rect 36378 11766 36397 11787
rect 36417 11771 36438 11787
rect 36458 11771 37369 11792
rect 36417 11766 37369 11771
rect 36378 11758 37369 11766
rect 36383 11735 36489 11758
rect 36383 11732 36488 11735
rect 36232 11671 36625 11691
rect 36645 11671 36648 11691
rect 36232 11666 36648 11671
rect 36232 11665 36573 11666
rect 35889 11634 35999 11648
rect 35889 11631 35932 11634
rect 35889 11626 35893 11631
rect 35811 11604 35893 11626
rect 35922 11604 35932 11631
rect 35960 11607 35967 11634
rect 35996 11626 35999 11634
rect 35996 11607 36061 11626
rect 35960 11604 36061 11607
rect 35811 11602 36061 11604
rect 35811 11523 35848 11602
rect 35889 11589 35999 11602
rect 35963 11533 35994 11534
rect 35811 11503 35820 11523
rect 35840 11503 35848 11523
rect 35811 11493 35848 11503
rect 35907 11523 35994 11533
rect 35907 11503 35916 11523
rect 35936 11503 35994 11523
rect 35907 11494 35994 11503
rect 35907 11493 35944 11494
rect 35477 11441 35569 11477
rect 35963 11441 35994 11494
rect 36024 11523 36061 11602
rect 36176 11533 36207 11534
rect 36024 11503 36033 11523
rect 36053 11503 36061 11523
rect 36024 11493 36061 11503
rect 36120 11526 36207 11533
rect 36120 11523 36181 11526
rect 36120 11503 36129 11523
rect 36149 11506 36181 11523
rect 36202 11506 36207 11526
rect 36149 11503 36207 11506
rect 36120 11496 36207 11503
rect 36232 11523 36269 11665
rect 36535 11664 36572 11665
rect 36384 11533 36420 11534
rect 36232 11503 36241 11523
rect 36261 11503 36269 11523
rect 36120 11494 36176 11496
rect 36120 11493 36157 11494
rect 36232 11493 36269 11503
rect 36328 11523 36476 11533
rect 36576 11530 36672 11532
rect 36328 11503 36337 11523
rect 36357 11503 36447 11523
rect 36467 11503 36476 11523
rect 36328 11497 36476 11503
rect 36328 11494 36392 11497
rect 36328 11493 36365 11494
rect 36384 11467 36392 11494
rect 36413 11494 36476 11497
rect 36534 11523 36672 11530
rect 36534 11503 36543 11523
rect 36563 11503 36672 11523
rect 36534 11494 36672 11503
rect 36413 11467 36420 11494
rect 36439 11493 36476 11494
rect 36535 11493 36572 11494
rect 36384 11442 36420 11467
rect 35477 11440 35813 11441
rect 35855 11440 35896 11441
rect 35477 11433 35896 11440
rect 35477 11413 35865 11433
rect 35885 11413 35896 11433
rect 35477 11405 35896 11413
rect 35963 11437 36322 11441
rect 35963 11432 36285 11437
rect 35963 11408 36076 11432
rect 36100 11413 36285 11432
rect 36309 11413 36322 11437
rect 36100 11408 36322 11413
rect 35963 11405 36322 11408
rect 36384 11405 36419 11442
rect 36487 11439 36587 11442
rect 36487 11435 36554 11439
rect 36487 11409 36499 11435
rect 36525 11413 36554 11435
rect 36580 11413 36587 11439
rect 36525 11409 36587 11413
rect 36487 11405 36587 11409
rect 35477 11401 35813 11405
rect 35310 11083 35382 11133
rect 30618 11009 30694 11033
rect 30618 10943 30630 11009
rect 30684 10943 30694 11009
rect 31162 10964 31203 10966
rect 31434 10964 31538 10966
rect 31896 10964 31957 11039
rect 32933 10987 32994 11062
rect 33352 11060 33456 11062
rect 33687 11060 33728 11062
rect 34196 11017 34206 11083
rect 34260 11017 34272 11083
rect 34196 10993 34272 11017
rect 29508 10893 29580 10943
rect 28219 10801 28663 10827
rect 28219 10799 28387 10801
rect 28219 10532 28246 10799
rect 28516 10797 28545 10801
rect 28286 10672 28350 10684
rect 28626 10680 28663 10801
rect 28891 10769 29002 10784
rect 28891 10767 28933 10769
rect 28891 10747 28898 10767
rect 28917 10747 28933 10767
rect 28891 10739 28933 10747
rect 28961 10767 29002 10769
rect 28961 10747 28975 10767
rect 28994 10747 29002 10767
rect 28961 10739 29002 10747
rect 28891 10733 29002 10739
rect 28834 10711 29083 10733
rect 28834 10680 28871 10711
rect 29047 10709 29083 10711
rect 29047 10680 29084 10709
rect 28286 10671 28321 10672
rect 28263 10666 28321 10671
rect 28263 10646 28266 10666
rect 28286 10652 28321 10666
rect 28341 10652 28350 10672
rect 28286 10644 28350 10652
rect 28312 10643 28350 10644
rect 28313 10642 28350 10643
rect 28416 10676 28452 10677
rect 28524 10676 28560 10677
rect 28416 10668 28560 10676
rect 28416 10648 28424 10668
rect 28444 10648 28532 10668
rect 28552 10648 28560 10668
rect 28416 10642 28560 10648
rect 28626 10672 28664 10680
rect 28732 10676 28768 10677
rect 28626 10652 28635 10672
rect 28655 10652 28664 10672
rect 28626 10643 28664 10652
rect 28683 10669 28768 10676
rect 28683 10649 28690 10669
rect 28711 10668 28768 10669
rect 28711 10649 28740 10668
rect 28683 10648 28740 10649
rect 28760 10648 28768 10668
rect 28626 10642 28663 10643
rect 28683 10642 28768 10648
rect 28834 10672 28872 10680
rect 28945 10676 28981 10677
rect 28834 10652 28843 10672
rect 28863 10652 28872 10672
rect 28834 10643 28872 10652
rect 28896 10668 28981 10676
rect 28896 10648 28953 10668
rect 28973 10648 28981 10668
rect 28834 10642 28871 10643
rect 28896 10642 28981 10648
rect 29047 10672 29085 10680
rect 29047 10652 29056 10672
rect 29076 10652 29085 10672
rect 29047 10643 29085 10652
rect 29047 10642 29084 10643
rect 28470 10621 28506 10642
rect 28896 10621 28927 10642
rect 29077 10621 29411 10625
rect 28303 10617 28403 10621
rect 28303 10613 28365 10617
rect 28303 10587 28310 10613
rect 28336 10591 28365 10613
rect 28391 10591 28403 10617
rect 28336 10587 28403 10591
rect 28303 10584 28403 10587
rect 28471 10584 28506 10621
rect 28568 10618 28927 10621
rect 28568 10613 28790 10618
rect 28568 10589 28581 10613
rect 28605 10594 28790 10613
rect 28814 10594 28927 10618
rect 28605 10589 28927 10594
rect 28568 10585 28927 10589
rect 28994 10613 29411 10621
rect 28994 10593 29005 10613
rect 29025 10593 29411 10613
rect 28994 10586 29411 10593
rect 28994 10585 29035 10586
rect 29077 10585 29411 10586
rect 28470 10559 28506 10584
rect 28318 10532 28355 10533
rect 28414 10532 28451 10533
rect 28470 10532 28477 10559
rect 28218 10523 28356 10532
rect 28218 10503 28327 10523
rect 28347 10503 28356 10523
rect 28218 10496 28356 10503
rect 28414 10529 28477 10532
rect 28498 10532 28506 10559
rect 28525 10532 28562 10533
rect 28498 10529 28562 10532
rect 28414 10523 28562 10529
rect 28414 10503 28423 10523
rect 28443 10503 28533 10523
rect 28553 10503 28562 10523
rect 28218 10494 28314 10496
rect 28414 10493 28562 10503
rect 28621 10523 28658 10533
rect 28733 10532 28770 10533
rect 28714 10530 28770 10532
rect 28621 10503 28629 10523
rect 28649 10503 28658 10523
rect 28470 10492 28506 10493
rect 28318 10361 28355 10362
rect 28621 10361 28658 10503
rect 28683 10523 28770 10530
rect 28683 10520 28741 10523
rect 28683 10500 28688 10520
rect 28709 10503 28741 10520
rect 28761 10503 28770 10523
rect 28709 10500 28770 10503
rect 28683 10493 28770 10500
rect 28829 10523 28866 10533
rect 28829 10503 28837 10523
rect 28857 10503 28866 10523
rect 28683 10492 28714 10493
rect 28829 10424 28866 10503
rect 28896 10532 28927 10585
rect 28946 10532 28983 10533
rect 28896 10523 28983 10532
rect 28896 10503 28954 10523
rect 28974 10503 28983 10523
rect 28896 10493 28983 10503
rect 29042 10523 29079 10533
rect 29042 10503 29050 10523
rect 29070 10503 29079 10523
rect 28896 10492 28927 10493
rect 28891 10424 29001 10437
rect 29042 10424 29079 10503
rect 28829 10422 29079 10424
rect 28829 10419 28930 10422
rect 28829 10400 28894 10419
rect 28891 10392 28894 10400
rect 28923 10392 28930 10419
rect 28958 10395 28968 10422
rect 28997 10400 29079 10422
rect 28997 10395 29001 10400
rect 28958 10392 29001 10395
rect 28891 10378 29001 10392
rect 28317 10360 28658 10361
rect 28242 10355 28658 10360
rect 28242 10335 28245 10355
rect 28265 10335 28658 10355
rect 28551 9970 28582 10335
rect 28469 9941 28582 9970
rect 28470 9641 28506 9941
rect 29330 9836 29411 10585
rect 29510 9984 29580 10893
rect 30618 10923 30694 10943
rect 30618 10886 30635 10923
rect 30679 10886 30694 10923
rect 30755 10929 31957 10964
rect 30755 10915 30783 10929
rect 30618 10870 30694 10886
rect 30623 10714 30693 10870
rect 30757 10784 30783 10915
rect 31162 10926 31957 10929
rect 30615 10663 30695 10714
rect 30615 10637 30631 10663
rect 30671 10637 30695 10663
rect 30615 10618 30695 10637
rect 30615 10592 30634 10618
rect 30674 10592 30695 10618
rect 30615 10565 30695 10592
rect 30615 10539 30638 10565
rect 30678 10539 30695 10565
rect 30615 10528 30695 10539
rect 30757 10529 30784 10784
rect 31162 10776 31203 10926
rect 31896 10914 31957 10926
rect 31629 10864 31750 10882
rect 31629 10862 31700 10864
rect 31629 10821 31644 10862
rect 31681 10823 31700 10862
rect 31737 10823 31750 10864
rect 31681 10821 31750 10823
rect 31629 10811 31750 10821
rect 31434 10781 31538 10790
rect 30824 10669 30888 10681
rect 31164 10677 31201 10776
rect 31429 10766 31540 10781
rect 31429 10764 31471 10766
rect 31429 10744 31436 10764
rect 31455 10744 31471 10764
rect 31429 10736 31471 10744
rect 31499 10764 31540 10766
rect 31499 10744 31513 10764
rect 31532 10744 31540 10764
rect 31499 10736 31540 10744
rect 31429 10730 31540 10736
rect 31372 10708 31621 10730
rect 31372 10677 31409 10708
rect 31585 10706 31621 10708
rect 31585 10677 31622 10706
rect 30824 10668 30859 10669
rect 30801 10663 30859 10668
rect 30801 10643 30804 10663
rect 30824 10649 30859 10663
rect 30879 10649 30888 10669
rect 30824 10641 30888 10649
rect 30850 10640 30888 10641
rect 30851 10639 30888 10640
rect 30954 10673 30990 10674
rect 31062 10673 31098 10674
rect 30954 10665 31098 10673
rect 30954 10645 30962 10665
rect 30982 10645 31070 10665
rect 31090 10645 31098 10665
rect 30954 10639 31098 10645
rect 31164 10669 31202 10677
rect 31270 10673 31306 10674
rect 31164 10649 31173 10669
rect 31193 10649 31202 10669
rect 31164 10640 31202 10649
rect 31221 10666 31306 10673
rect 31221 10646 31228 10666
rect 31249 10665 31306 10666
rect 31249 10646 31278 10665
rect 31221 10645 31278 10646
rect 31298 10645 31306 10665
rect 31164 10639 31201 10640
rect 31221 10639 31306 10645
rect 31372 10669 31410 10677
rect 31483 10673 31519 10674
rect 31372 10649 31381 10669
rect 31401 10649 31410 10669
rect 31372 10640 31410 10649
rect 31434 10665 31519 10673
rect 31434 10645 31491 10665
rect 31511 10645 31519 10665
rect 31372 10639 31409 10640
rect 31434 10639 31519 10645
rect 31585 10669 31623 10677
rect 31585 10649 31594 10669
rect 31614 10649 31623 10669
rect 31678 10659 31743 10811
rect 31896 10785 31951 10914
rect 32935 10857 32994 10987
rect 33848 10938 33920 10939
rect 33847 10930 33946 10938
rect 33847 10927 33899 10930
rect 33847 10892 33855 10927
rect 33880 10892 33899 10927
rect 33924 10919 33946 10930
rect 33924 10918 34791 10919
rect 33924 10892 34792 10918
rect 33847 10882 34792 10892
rect 33847 10880 33946 10882
rect 32935 10839 32957 10857
rect 32975 10839 32994 10857
rect 32935 10817 32994 10839
rect 33202 10853 33734 10858
rect 33202 10833 34088 10853
rect 34108 10833 34111 10853
rect 34747 10849 34792 10882
rect 33202 10829 34111 10833
rect 31585 10640 31623 10649
rect 31676 10652 31743 10659
rect 31585 10639 31622 10640
rect 31008 10618 31044 10639
rect 31434 10618 31465 10639
rect 31676 10631 31693 10652
rect 31729 10631 31743 10652
rect 31895 10672 31951 10785
rect 33202 10782 33245 10829
rect 33695 10828 34111 10829
rect 34743 10829 35136 10849
rect 35156 10829 35159 10849
rect 33695 10827 34036 10828
rect 33352 10796 33462 10810
rect 33352 10793 33395 10796
rect 33352 10788 33356 10793
rect 33190 10781 33245 10782
rect 31895 10654 31914 10672
rect 31932 10654 31951 10672
rect 31895 10634 31951 10654
rect 32934 10758 33245 10781
rect 32934 10740 32959 10758
rect 32977 10746 33245 10758
rect 33274 10766 33356 10788
rect 33385 10766 33395 10793
rect 33423 10769 33430 10796
rect 33459 10788 33462 10796
rect 33459 10769 33524 10788
rect 33423 10766 33524 10769
rect 33274 10764 33524 10766
rect 32977 10740 32999 10746
rect 31676 10618 31743 10631
rect 30841 10614 30941 10618
rect 30841 10610 30903 10614
rect 30841 10584 30848 10610
rect 30874 10588 30903 10610
rect 30929 10588 30941 10614
rect 30874 10584 30941 10588
rect 30841 10581 30941 10584
rect 31009 10581 31044 10618
rect 31106 10615 31465 10618
rect 31106 10610 31328 10615
rect 31106 10586 31119 10610
rect 31143 10591 31328 10610
rect 31352 10591 31465 10615
rect 31143 10586 31465 10591
rect 31106 10582 31465 10586
rect 31532 10612 31743 10618
rect 31532 10610 31693 10612
rect 31532 10590 31543 10610
rect 31563 10590 31693 10610
rect 31532 10583 31693 10590
rect 31532 10582 31573 10583
rect 31008 10556 31044 10581
rect 30856 10529 30893 10530
rect 30952 10529 30989 10530
rect 31008 10529 31015 10556
rect 30756 10520 30894 10529
rect 30756 10500 30865 10520
rect 30885 10500 30894 10520
rect 30756 10493 30894 10500
rect 30952 10526 31015 10529
rect 31036 10529 31044 10556
rect 31063 10529 31100 10530
rect 31036 10526 31100 10529
rect 30952 10520 31100 10526
rect 30952 10500 30961 10520
rect 30981 10500 31071 10520
rect 31091 10500 31100 10520
rect 30756 10491 30852 10493
rect 30952 10490 31100 10500
rect 31159 10520 31196 10530
rect 31271 10529 31308 10530
rect 31252 10527 31308 10529
rect 31159 10500 31167 10520
rect 31187 10500 31196 10520
rect 31008 10489 31044 10490
rect 30856 10358 30893 10359
rect 31159 10358 31196 10500
rect 31221 10520 31308 10527
rect 31221 10517 31279 10520
rect 31221 10497 31226 10517
rect 31247 10500 31279 10517
rect 31299 10500 31308 10520
rect 31247 10497 31308 10500
rect 31221 10490 31308 10497
rect 31367 10520 31404 10530
rect 31367 10500 31375 10520
rect 31395 10500 31404 10520
rect 31221 10489 31252 10490
rect 31367 10421 31404 10500
rect 31434 10529 31465 10582
rect 31678 10575 31693 10583
rect 31733 10575 31743 10612
rect 32934 10601 32999 10740
rect 33274 10685 33311 10764
rect 33352 10751 33462 10764
rect 33426 10695 33457 10696
rect 33274 10665 33283 10685
rect 33303 10665 33311 10685
rect 31678 10566 31743 10575
rect 31891 10573 31956 10594
rect 31891 10555 31916 10573
rect 31934 10555 31956 10573
rect 32934 10583 32957 10601
rect 32975 10583 32999 10601
rect 32934 10566 32999 10583
rect 33154 10647 33222 10660
rect 33274 10655 33311 10665
rect 33370 10685 33457 10695
rect 33370 10665 33379 10685
rect 33399 10665 33457 10685
rect 33370 10656 33457 10665
rect 33370 10655 33407 10656
rect 33154 10605 33161 10647
rect 33210 10605 33222 10647
rect 33154 10602 33222 10605
rect 33426 10603 33457 10656
rect 33487 10685 33524 10764
rect 33639 10695 33670 10696
rect 33487 10665 33496 10685
rect 33516 10665 33524 10685
rect 33487 10655 33524 10665
rect 33583 10688 33670 10695
rect 33583 10685 33644 10688
rect 33583 10665 33592 10685
rect 33612 10668 33644 10685
rect 33665 10668 33670 10688
rect 33612 10665 33670 10668
rect 33583 10658 33670 10665
rect 33695 10685 33732 10827
rect 33998 10826 34035 10827
rect 34743 10824 35159 10829
rect 34743 10823 35084 10824
rect 34400 10792 34510 10806
rect 34400 10789 34443 10792
rect 34400 10784 34404 10789
rect 34322 10762 34404 10784
rect 34433 10762 34443 10789
rect 34471 10765 34478 10792
rect 34507 10784 34510 10792
rect 34507 10765 34572 10784
rect 34471 10762 34572 10765
rect 34322 10760 34572 10762
rect 33847 10695 33883 10696
rect 33695 10665 33704 10685
rect 33724 10665 33732 10685
rect 33583 10656 33639 10658
rect 33583 10655 33620 10656
rect 33695 10655 33732 10665
rect 33791 10685 33939 10695
rect 34039 10692 34135 10694
rect 33791 10665 33800 10685
rect 33820 10665 33910 10685
rect 33930 10665 33939 10685
rect 33791 10659 33939 10665
rect 33791 10656 33855 10659
rect 33791 10655 33828 10656
rect 33847 10629 33855 10656
rect 33876 10656 33939 10659
rect 33997 10685 34135 10692
rect 33997 10665 34006 10685
rect 34026 10665 34135 10685
rect 33997 10656 34135 10665
rect 34322 10681 34359 10760
rect 34400 10747 34510 10760
rect 34474 10691 34505 10692
rect 34322 10661 34331 10681
rect 34351 10661 34359 10681
rect 33876 10629 33883 10656
rect 33902 10655 33939 10656
rect 33998 10655 34035 10656
rect 33847 10604 33883 10629
rect 33318 10602 33359 10603
rect 33154 10595 33359 10602
rect 33154 10584 33328 10595
rect 31484 10529 31521 10530
rect 31434 10520 31521 10529
rect 31434 10500 31492 10520
rect 31512 10500 31521 10520
rect 31434 10490 31521 10500
rect 31580 10520 31617 10530
rect 31580 10500 31588 10520
rect 31608 10500 31617 10520
rect 31434 10489 31465 10490
rect 31429 10421 31539 10434
rect 31580 10421 31617 10500
rect 31891 10479 31956 10555
rect 33154 10551 33162 10584
rect 33155 10542 33162 10551
rect 33211 10575 33328 10584
rect 33348 10575 33359 10595
rect 33211 10567 33359 10575
rect 33426 10599 33785 10603
rect 33426 10594 33748 10599
rect 33426 10570 33539 10594
rect 33563 10575 33748 10594
rect 33772 10575 33785 10599
rect 33563 10570 33785 10575
rect 33426 10567 33785 10570
rect 33847 10567 33882 10604
rect 33950 10601 34050 10604
rect 33950 10597 34017 10601
rect 33950 10571 33962 10597
rect 33988 10575 34017 10597
rect 34043 10575 34050 10601
rect 33988 10571 34050 10575
rect 33950 10567 34050 10571
rect 33211 10551 33222 10567
rect 33211 10542 33219 10551
rect 33426 10546 33457 10567
rect 33847 10546 33883 10567
rect 33269 10545 33306 10546
rect 32934 10502 32999 10521
rect 32934 10484 32959 10502
rect 32977 10484 32999 10502
rect 31367 10419 31617 10421
rect 31367 10416 31468 10419
rect 31367 10397 31432 10416
rect 31429 10389 31432 10397
rect 31461 10389 31468 10416
rect 31496 10392 31506 10419
rect 31535 10397 31617 10419
rect 31640 10444 31957 10479
rect 31535 10392 31539 10397
rect 31496 10389 31539 10392
rect 31429 10375 31539 10389
rect 30855 10357 31196 10358
rect 30780 10355 31196 10357
rect 31640 10355 31680 10444
rect 31891 10417 31956 10444
rect 31891 10399 31914 10417
rect 31932 10399 31956 10417
rect 31891 10379 31956 10399
rect 30777 10352 31680 10355
rect 30777 10332 30783 10352
rect 30803 10332 31680 10352
rect 30777 10328 31680 10332
rect 31640 10325 31680 10328
rect 31892 10318 31957 10339
rect 30110 10310 30771 10311
rect 30110 10303 31044 10310
rect 30110 10302 31016 10303
rect 30110 10282 30961 10302
rect 30993 10283 31016 10302
rect 31041 10283 31044 10303
rect 30993 10282 31044 10283
rect 30110 10275 31044 10282
rect 29709 10233 29877 10234
rect 30112 10233 30151 10275
rect 30940 10273 31044 10275
rect 31009 10271 31044 10273
rect 31892 10300 31916 10318
rect 31934 10300 31957 10318
rect 31892 10253 31957 10300
rect 29709 10207 30153 10233
rect 29709 10205 29877 10207
rect 28470 9618 28474 9641
rect 28498 9618 28506 9641
rect 28670 9619 28769 9623
rect 28470 9597 28506 9618
rect 28470 9574 28474 9597
rect 28498 9574 28506 9597
rect 28470 9570 28506 9574
rect 28666 9613 28769 9619
rect 28666 9575 28692 9613
rect 28717 9578 28736 9613
rect 28761 9578 28769 9613
rect 28717 9575 28769 9578
rect 28666 9567 28769 9575
rect 28666 9566 28768 9567
rect 28262 9488 28430 9489
rect 28666 9488 28713 9566
rect 28262 9462 28713 9488
rect 28262 9460 28430 9462
rect 28262 9087 28289 9460
rect 28459 9412 28545 9421
rect 28459 9394 28478 9412
rect 28530 9394 28545 9412
rect 28459 9390 28545 9394
rect 28329 9227 28393 9239
rect 28329 9226 28364 9227
rect 28306 9221 28364 9226
rect 28306 9201 28309 9221
rect 28329 9207 28364 9221
rect 28384 9207 28393 9227
rect 28329 9199 28393 9207
rect 28355 9198 28393 9199
rect 28356 9197 28393 9198
rect 28459 9231 28495 9232
rect 28515 9231 28545 9390
rect 28666 9350 28713 9462
rect 28669 9235 28706 9350
rect 28934 9324 29045 9339
rect 28934 9322 28976 9324
rect 28934 9302 28941 9322
rect 28960 9302 28976 9322
rect 28934 9294 28976 9302
rect 29004 9322 29045 9324
rect 29004 9302 29018 9322
rect 29037 9302 29045 9322
rect 29004 9294 29045 9302
rect 28934 9288 29045 9294
rect 28877 9266 29126 9288
rect 28877 9235 28914 9266
rect 29090 9264 29126 9266
rect 29090 9235 29127 9264
rect 29331 9251 29410 9836
rect 29507 9384 29586 9984
rect 29709 9854 29736 10205
rect 30112 10201 30153 10207
rect 29776 9994 29840 10006
rect 30116 10002 30153 10201
rect 30615 10228 30687 10245
rect 30615 10189 30623 10228
rect 30668 10189 30687 10228
rect 30381 10091 30492 10106
rect 30381 10089 30423 10091
rect 30381 10069 30388 10089
rect 30407 10069 30423 10089
rect 30381 10061 30423 10069
rect 30451 10089 30492 10091
rect 30451 10069 30465 10089
rect 30484 10069 30492 10089
rect 30451 10061 30492 10069
rect 30381 10055 30492 10061
rect 30324 10033 30573 10055
rect 30324 10002 30361 10033
rect 30537 10031 30573 10033
rect 30537 10002 30574 10031
rect 29776 9993 29811 9994
rect 29753 9988 29811 9993
rect 29753 9968 29756 9988
rect 29776 9974 29811 9988
rect 29831 9974 29840 9994
rect 29776 9966 29840 9974
rect 29802 9965 29840 9966
rect 29803 9964 29840 9965
rect 29906 9998 29942 9999
rect 30014 9998 30050 9999
rect 29906 9990 30050 9998
rect 29906 9970 29914 9990
rect 29934 9970 30022 9990
rect 30042 9970 30050 9990
rect 29906 9964 30050 9970
rect 30116 9994 30154 10002
rect 30222 9998 30258 9999
rect 30116 9974 30125 9994
rect 30145 9974 30154 9994
rect 30116 9965 30154 9974
rect 30173 9991 30258 9998
rect 30173 9971 30180 9991
rect 30201 9990 30258 9991
rect 30201 9971 30230 9990
rect 30173 9970 30230 9971
rect 30250 9970 30258 9990
rect 30116 9964 30153 9965
rect 30173 9964 30258 9970
rect 30324 9994 30362 10002
rect 30435 9998 30471 9999
rect 30324 9974 30333 9994
rect 30353 9974 30362 9994
rect 30324 9965 30362 9974
rect 30386 9990 30471 9998
rect 30386 9970 30443 9990
rect 30463 9970 30471 9990
rect 30324 9964 30361 9965
rect 30386 9964 30471 9970
rect 30537 9994 30575 10002
rect 30537 9974 30546 9994
rect 30566 9974 30575 9994
rect 30537 9965 30575 9974
rect 30615 9979 30687 10189
rect 30757 10223 31957 10253
rect 30757 10222 31201 10223
rect 30757 10220 30925 10222
rect 30615 9965 30698 9979
rect 30537 9964 30574 9965
rect 29960 9943 29996 9964
rect 30386 9943 30417 9964
rect 30615 9943 30632 9965
rect 29793 9939 29893 9943
rect 29793 9935 29855 9939
rect 29793 9909 29800 9935
rect 29826 9913 29855 9935
rect 29881 9913 29893 9939
rect 29826 9909 29893 9913
rect 29793 9906 29893 9909
rect 29961 9906 29996 9943
rect 30058 9940 30417 9943
rect 30058 9935 30280 9940
rect 30058 9911 30071 9935
rect 30095 9916 30280 9935
rect 30304 9916 30417 9940
rect 30095 9911 30417 9916
rect 30058 9907 30417 9911
rect 30484 9935 30632 9943
rect 30484 9915 30495 9935
rect 30515 9932 30632 9935
rect 30685 9932 30698 9965
rect 30515 9915 30698 9932
rect 30484 9908 30698 9915
rect 30484 9907 30525 9908
rect 30615 9907 30698 9908
rect 29960 9881 29996 9906
rect 29808 9854 29845 9855
rect 29904 9854 29941 9855
rect 29960 9854 29967 9881
rect 29708 9845 29846 9854
rect 29708 9825 29817 9845
rect 29837 9825 29846 9845
rect 29708 9818 29846 9825
rect 29904 9851 29967 9854
rect 29988 9854 29996 9881
rect 30015 9854 30052 9855
rect 29988 9851 30052 9854
rect 29904 9845 30052 9851
rect 29904 9825 29913 9845
rect 29933 9825 30023 9845
rect 30043 9825 30052 9845
rect 29708 9816 29804 9818
rect 29904 9815 30052 9825
rect 30111 9845 30148 9855
rect 30223 9854 30260 9855
rect 30204 9852 30260 9854
rect 30111 9825 30119 9845
rect 30139 9825 30148 9845
rect 29960 9814 29996 9815
rect 29808 9683 29845 9684
rect 30111 9683 30148 9825
rect 30173 9845 30260 9852
rect 30173 9842 30231 9845
rect 30173 9822 30178 9842
rect 30199 9825 30231 9842
rect 30251 9825 30260 9845
rect 30199 9822 30260 9825
rect 30173 9815 30260 9822
rect 30319 9845 30356 9855
rect 30319 9825 30327 9845
rect 30347 9825 30356 9845
rect 30173 9814 30204 9815
rect 30319 9746 30356 9825
rect 30386 9854 30417 9907
rect 30623 9874 30637 9907
rect 30690 9874 30698 9907
rect 30623 9868 30698 9874
rect 30623 9863 30693 9868
rect 30436 9854 30473 9855
rect 30386 9845 30473 9854
rect 30386 9825 30444 9845
rect 30464 9825 30473 9845
rect 30386 9815 30473 9825
rect 30532 9845 30569 9855
rect 30757 9850 30784 10220
rect 30824 9990 30888 10002
rect 31164 9998 31201 10222
rect 31672 10203 31736 10205
rect 31668 10191 31736 10203
rect 31668 10158 31679 10191
rect 31719 10158 31736 10191
rect 31668 10148 31736 10158
rect 31429 10087 31540 10102
rect 31429 10085 31471 10087
rect 31429 10065 31436 10085
rect 31455 10065 31471 10085
rect 31429 10057 31471 10065
rect 31499 10085 31540 10087
rect 31499 10065 31513 10085
rect 31532 10065 31540 10085
rect 31499 10057 31540 10065
rect 31429 10051 31540 10057
rect 31372 10029 31621 10051
rect 31372 9998 31409 10029
rect 31585 10027 31621 10029
rect 31585 9998 31622 10027
rect 30824 9989 30859 9990
rect 30801 9984 30859 9989
rect 30801 9964 30804 9984
rect 30824 9970 30859 9984
rect 30879 9970 30888 9990
rect 30824 9962 30888 9970
rect 30850 9961 30888 9962
rect 30851 9960 30888 9961
rect 30954 9994 30990 9995
rect 31062 9994 31098 9995
rect 30954 9986 31098 9994
rect 30954 9966 30962 9986
rect 30982 9966 31070 9986
rect 31090 9966 31098 9986
rect 30954 9960 31098 9966
rect 31164 9990 31202 9998
rect 31270 9994 31306 9995
rect 31164 9970 31173 9990
rect 31193 9970 31202 9990
rect 31164 9961 31202 9970
rect 31221 9987 31306 9994
rect 31221 9967 31228 9987
rect 31249 9986 31306 9987
rect 31249 9967 31278 9986
rect 31221 9966 31278 9967
rect 31298 9966 31306 9986
rect 31164 9960 31201 9961
rect 31221 9960 31306 9966
rect 31372 9990 31410 9998
rect 31483 9994 31519 9995
rect 31372 9970 31381 9990
rect 31401 9970 31410 9990
rect 31372 9961 31410 9970
rect 31434 9986 31519 9994
rect 31434 9966 31491 9986
rect 31511 9966 31519 9986
rect 31372 9960 31409 9961
rect 31434 9960 31519 9966
rect 31585 9990 31623 9998
rect 31585 9970 31594 9990
rect 31614 9970 31623 9990
rect 31585 9961 31623 9970
rect 31672 9964 31736 10148
rect 31892 10022 31957 10223
rect 32934 10283 32999 10484
rect 33155 10358 33219 10542
rect 33268 10536 33306 10545
rect 33268 10516 33277 10536
rect 33297 10516 33306 10536
rect 33268 10508 33306 10516
rect 33372 10540 33457 10546
rect 33482 10545 33519 10546
rect 33372 10520 33380 10540
rect 33400 10520 33457 10540
rect 33372 10512 33457 10520
rect 33481 10536 33519 10545
rect 33481 10516 33490 10536
rect 33510 10516 33519 10536
rect 33372 10511 33408 10512
rect 33481 10508 33519 10516
rect 33585 10540 33670 10546
rect 33690 10545 33727 10546
rect 33585 10520 33593 10540
rect 33613 10539 33670 10540
rect 33613 10520 33642 10539
rect 33585 10519 33642 10520
rect 33663 10519 33670 10539
rect 33585 10512 33670 10519
rect 33689 10536 33727 10545
rect 33689 10516 33698 10536
rect 33718 10516 33727 10536
rect 33585 10511 33621 10512
rect 33689 10508 33727 10516
rect 33793 10540 33937 10546
rect 33793 10520 33801 10540
rect 33821 10520 33909 10540
rect 33929 10520 33937 10540
rect 33793 10512 33937 10520
rect 33793 10511 33829 10512
rect 33901 10511 33937 10512
rect 34003 10545 34040 10546
rect 34003 10544 34041 10545
rect 34003 10536 34067 10544
rect 34003 10516 34012 10536
rect 34032 10522 34067 10536
rect 34087 10522 34090 10542
rect 34032 10517 34090 10522
rect 34032 10516 34067 10517
rect 33269 10479 33306 10508
rect 33270 10477 33306 10479
rect 33482 10477 33519 10508
rect 33270 10455 33519 10477
rect 33351 10449 33462 10455
rect 33351 10441 33392 10449
rect 33351 10421 33359 10441
rect 33378 10421 33392 10441
rect 33351 10419 33392 10421
rect 33420 10441 33462 10449
rect 33420 10421 33436 10441
rect 33455 10421 33462 10441
rect 33420 10419 33462 10421
rect 33351 10404 33462 10419
rect 33155 10348 33223 10358
rect 33155 10315 33172 10348
rect 33212 10315 33223 10348
rect 33155 10303 33223 10315
rect 33155 10301 33219 10303
rect 33690 10284 33727 10508
rect 34003 10504 34067 10516
rect 34107 10286 34134 10656
rect 34322 10651 34359 10661
rect 34418 10681 34505 10691
rect 34418 10661 34427 10681
rect 34447 10661 34505 10681
rect 34418 10652 34505 10661
rect 34418 10651 34455 10652
rect 34198 10638 34268 10643
rect 34193 10632 34268 10638
rect 34193 10599 34201 10632
rect 34254 10599 34268 10632
rect 34474 10599 34505 10652
rect 34535 10681 34572 10760
rect 34687 10691 34718 10692
rect 34535 10661 34544 10681
rect 34564 10661 34572 10681
rect 34535 10651 34572 10661
rect 34631 10684 34718 10691
rect 34631 10681 34692 10684
rect 34631 10661 34640 10681
rect 34660 10664 34692 10681
rect 34713 10664 34718 10684
rect 34660 10661 34718 10664
rect 34631 10654 34718 10661
rect 34743 10681 34780 10823
rect 35046 10822 35083 10823
rect 34895 10691 34931 10692
rect 34743 10661 34752 10681
rect 34772 10661 34780 10681
rect 34631 10652 34687 10654
rect 34631 10651 34668 10652
rect 34743 10651 34780 10661
rect 34839 10681 34987 10691
rect 35087 10688 35183 10690
rect 34839 10661 34848 10681
rect 34868 10661 34958 10681
rect 34978 10661 34987 10681
rect 34839 10655 34987 10661
rect 34839 10652 34903 10655
rect 34839 10651 34876 10652
rect 34895 10625 34903 10652
rect 34924 10652 34987 10655
rect 35045 10681 35183 10688
rect 35045 10661 35054 10681
rect 35074 10661 35183 10681
rect 35045 10652 35183 10661
rect 34924 10625 34931 10652
rect 34950 10651 34987 10652
rect 35046 10651 35083 10652
rect 34895 10600 34931 10625
rect 34193 10598 34276 10599
rect 34366 10598 34407 10599
rect 34193 10591 34407 10598
rect 34193 10574 34376 10591
rect 34193 10541 34206 10574
rect 34259 10571 34376 10574
rect 34396 10571 34407 10591
rect 34259 10563 34407 10571
rect 34474 10595 34833 10599
rect 34474 10590 34796 10595
rect 34474 10566 34587 10590
rect 34611 10571 34796 10590
rect 34820 10571 34833 10595
rect 34611 10566 34833 10571
rect 34474 10563 34833 10566
rect 34895 10563 34930 10600
rect 34998 10597 35098 10600
rect 34998 10593 35065 10597
rect 34998 10567 35010 10593
rect 35036 10571 35065 10593
rect 35091 10571 35098 10597
rect 35036 10567 35098 10571
rect 34998 10563 35098 10567
rect 34259 10541 34276 10563
rect 34474 10542 34505 10563
rect 34895 10542 34931 10563
rect 34317 10541 34354 10542
rect 34193 10527 34276 10541
rect 33966 10284 34134 10286
rect 33690 10283 34134 10284
rect 32934 10253 34134 10283
rect 34204 10317 34276 10527
rect 34316 10532 34354 10541
rect 34316 10512 34325 10532
rect 34345 10512 34354 10532
rect 34316 10504 34354 10512
rect 34420 10536 34505 10542
rect 34530 10541 34567 10542
rect 34420 10516 34428 10536
rect 34448 10516 34505 10536
rect 34420 10508 34505 10516
rect 34529 10532 34567 10541
rect 34529 10512 34538 10532
rect 34558 10512 34567 10532
rect 34420 10507 34456 10508
rect 34529 10504 34567 10512
rect 34633 10536 34718 10542
rect 34738 10541 34775 10542
rect 34633 10516 34641 10536
rect 34661 10535 34718 10536
rect 34661 10516 34690 10535
rect 34633 10515 34690 10516
rect 34711 10515 34718 10535
rect 34633 10508 34718 10515
rect 34737 10532 34775 10541
rect 34737 10512 34746 10532
rect 34766 10512 34775 10532
rect 34633 10507 34669 10508
rect 34737 10504 34775 10512
rect 34841 10536 34985 10542
rect 34841 10516 34849 10536
rect 34869 10516 34957 10536
rect 34977 10516 34985 10536
rect 34841 10508 34985 10516
rect 34841 10507 34877 10508
rect 34949 10507 34985 10508
rect 35051 10541 35088 10542
rect 35051 10540 35089 10541
rect 35051 10532 35115 10540
rect 35051 10512 35060 10532
rect 35080 10518 35115 10532
rect 35135 10518 35138 10538
rect 35080 10513 35138 10518
rect 35080 10512 35115 10513
rect 34317 10475 34354 10504
rect 34318 10473 34354 10475
rect 34530 10473 34567 10504
rect 34318 10451 34567 10473
rect 34399 10445 34510 10451
rect 34399 10437 34440 10445
rect 34399 10417 34407 10437
rect 34426 10417 34440 10437
rect 34399 10415 34440 10417
rect 34468 10437 34510 10445
rect 34468 10417 34484 10437
rect 34503 10417 34510 10437
rect 34468 10415 34510 10417
rect 34399 10400 34510 10415
rect 34204 10278 34223 10317
rect 34268 10278 34276 10317
rect 34204 10261 34276 10278
rect 34738 10305 34775 10504
rect 35051 10500 35115 10512
rect 34738 10299 34779 10305
rect 35155 10301 35182 10652
rect 35311 10604 35382 11083
rect 35311 10520 35380 10604
rect 35014 10299 35182 10301
rect 34738 10273 35182 10299
rect 32934 10206 32999 10253
rect 32934 10188 32957 10206
rect 32975 10188 32999 10206
rect 33847 10233 33882 10235
rect 33847 10231 33951 10233
rect 34740 10231 34779 10273
rect 35014 10272 35182 10273
rect 33847 10224 34781 10231
rect 33847 10223 33898 10224
rect 33847 10203 33850 10223
rect 33875 10204 33898 10223
rect 33930 10204 34781 10224
rect 33875 10203 34781 10204
rect 33847 10196 34781 10203
rect 34120 10195 34781 10196
rect 32934 10167 32999 10188
rect 33211 10178 33251 10181
rect 33211 10174 34114 10178
rect 33211 10154 34088 10174
rect 34108 10154 34114 10174
rect 33211 10151 34114 10154
rect 32935 10107 33000 10127
rect 32935 10089 32959 10107
rect 32977 10089 33000 10107
rect 32935 10062 33000 10089
rect 33211 10062 33251 10151
rect 33695 10149 34111 10151
rect 33695 10148 34036 10149
rect 33352 10117 33462 10131
rect 33352 10114 33395 10117
rect 33352 10109 33356 10114
rect 32934 10027 33251 10062
rect 33274 10087 33356 10109
rect 33385 10087 33395 10114
rect 33423 10090 33430 10117
rect 33459 10109 33462 10117
rect 33459 10090 33524 10109
rect 33423 10087 33524 10090
rect 33274 10085 33524 10087
rect 31892 10004 31914 10022
rect 31932 10004 31957 10022
rect 31892 9985 31957 10004
rect 31585 9960 31622 9961
rect 31008 9939 31044 9960
rect 31434 9939 31465 9960
rect 31672 9955 31680 9964
rect 31669 9939 31680 9955
rect 30841 9935 30941 9939
rect 30841 9931 30903 9935
rect 30841 9905 30848 9931
rect 30874 9909 30903 9931
rect 30929 9909 30941 9935
rect 30874 9905 30941 9909
rect 30841 9902 30941 9905
rect 31009 9902 31044 9939
rect 31106 9936 31465 9939
rect 31106 9931 31328 9936
rect 31106 9907 31119 9931
rect 31143 9912 31328 9931
rect 31352 9912 31465 9936
rect 31143 9907 31465 9912
rect 31106 9903 31465 9907
rect 31532 9931 31680 9939
rect 31532 9911 31543 9931
rect 31563 9922 31680 9931
rect 31729 9955 31736 9964
rect 31729 9922 31737 9955
rect 32935 9951 33000 10027
rect 33274 10006 33311 10085
rect 33352 10072 33462 10085
rect 33426 10016 33457 10017
rect 33274 9986 33283 10006
rect 33303 9986 33311 10006
rect 33274 9976 33311 9986
rect 33370 10006 33457 10016
rect 33370 9986 33379 10006
rect 33399 9986 33457 10006
rect 33370 9977 33457 9986
rect 33370 9976 33407 9977
rect 31563 9911 31737 9922
rect 31532 9904 31737 9911
rect 31532 9903 31573 9904
rect 31008 9877 31044 9902
rect 30856 9850 30893 9851
rect 30952 9850 30989 9851
rect 31008 9850 31015 9877
rect 30532 9825 30540 9845
rect 30560 9825 30569 9845
rect 30386 9814 30417 9815
rect 30381 9746 30491 9759
rect 30532 9746 30569 9825
rect 30756 9841 30894 9850
rect 30756 9821 30865 9841
rect 30885 9821 30894 9841
rect 30756 9814 30894 9821
rect 30952 9847 31015 9850
rect 31036 9850 31044 9877
rect 31063 9850 31100 9851
rect 31036 9847 31100 9850
rect 30952 9841 31100 9847
rect 30952 9821 30961 9841
rect 30981 9821 31071 9841
rect 31091 9821 31100 9841
rect 30756 9812 30852 9814
rect 30952 9811 31100 9821
rect 31159 9841 31196 9851
rect 31271 9850 31308 9851
rect 31252 9848 31308 9850
rect 31159 9821 31167 9841
rect 31187 9821 31196 9841
rect 31008 9810 31044 9811
rect 30319 9744 30569 9746
rect 30319 9741 30420 9744
rect 30319 9722 30384 9741
rect 30381 9714 30384 9722
rect 30413 9714 30420 9741
rect 30448 9717 30458 9744
rect 30487 9722 30569 9744
rect 30487 9717 30491 9722
rect 30448 9714 30491 9717
rect 30381 9700 30491 9714
rect 29807 9682 30148 9683
rect 29732 9677 30148 9682
rect 30856 9679 30893 9680
rect 31159 9679 31196 9821
rect 31221 9841 31308 9848
rect 31221 9838 31279 9841
rect 31221 9818 31226 9838
rect 31247 9821 31279 9838
rect 31299 9821 31308 9841
rect 31247 9818 31308 9821
rect 31221 9811 31308 9818
rect 31367 9841 31404 9851
rect 31367 9821 31375 9841
rect 31395 9821 31404 9841
rect 31221 9810 31252 9811
rect 31367 9742 31404 9821
rect 31434 9850 31465 9903
rect 31669 9901 31737 9904
rect 31669 9859 31681 9901
rect 31730 9859 31737 9901
rect 31484 9850 31521 9851
rect 31434 9841 31521 9850
rect 31434 9821 31492 9841
rect 31512 9821 31521 9841
rect 31434 9811 31521 9821
rect 31580 9841 31617 9851
rect 31669 9846 31737 9859
rect 31892 9923 31957 9940
rect 31892 9905 31916 9923
rect 31934 9905 31957 9923
rect 32935 9933 32957 9951
rect 32975 9933 33000 9951
rect 32935 9912 33000 9933
rect 33148 9931 33213 9940
rect 31580 9821 31588 9841
rect 31608 9821 31617 9841
rect 31434 9810 31465 9811
rect 31429 9742 31539 9755
rect 31580 9742 31617 9821
rect 31892 9766 31957 9905
rect 33148 9894 33158 9931
rect 33198 9923 33213 9931
rect 33426 9924 33457 9977
rect 33487 10006 33524 10085
rect 33639 10016 33670 10017
rect 33487 9986 33496 10006
rect 33516 9986 33524 10006
rect 33487 9976 33524 9986
rect 33583 10009 33670 10016
rect 33583 10006 33644 10009
rect 33583 9986 33592 10006
rect 33612 9989 33644 10006
rect 33665 9989 33670 10009
rect 33612 9986 33670 9989
rect 33583 9979 33670 9986
rect 33695 10006 33732 10148
rect 33998 10147 34035 10148
rect 33847 10016 33883 10017
rect 33695 9986 33704 10006
rect 33724 9986 33732 10006
rect 33583 9977 33639 9979
rect 33583 9976 33620 9977
rect 33695 9976 33732 9986
rect 33791 10006 33939 10016
rect 34039 10013 34135 10015
rect 33791 9986 33800 10006
rect 33820 9986 33910 10006
rect 33930 9986 33939 10006
rect 33791 9980 33939 9986
rect 33791 9977 33855 9980
rect 33791 9976 33828 9977
rect 33847 9950 33855 9977
rect 33876 9977 33939 9980
rect 33997 10006 34135 10013
rect 33997 9986 34006 10006
rect 34026 9986 34135 10006
rect 35315 10004 35377 10520
rect 33997 9977 34135 9986
rect 33876 9950 33883 9977
rect 33902 9976 33939 9977
rect 33998 9976 34035 9977
rect 33847 9925 33883 9950
rect 33318 9923 33359 9924
rect 33198 9916 33359 9923
rect 33198 9896 33328 9916
rect 33348 9896 33359 9916
rect 33198 9894 33359 9896
rect 33148 9888 33359 9894
rect 33426 9920 33785 9924
rect 33426 9915 33748 9920
rect 33426 9891 33539 9915
rect 33563 9896 33748 9915
rect 33772 9896 33785 9920
rect 33563 9891 33785 9896
rect 33426 9888 33785 9891
rect 33847 9888 33882 9925
rect 33950 9922 34050 9925
rect 33950 9918 34017 9922
rect 33950 9892 33962 9918
rect 33988 9896 34017 9918
rect 34043 9896 34050 9922
rect 33988 9892 34050 9896
rect 33950 9888 34050 9892
rect 33148 9875 33215 9888
rect 31892 9760 31914 9766
rect 31367 9740 31617 9742
rect 31367 9737 31468 9740
rect 31367 9718 31432 9737
rect 31429 9710 31432 9718
rect 31461 9710 31468 9737
rect 31496 9713 31506 9740
rect 31535 9718 31617 9740
rect 31646 9748 31914 9760
rect 31932 9748 31957 9766
rect 31646 9725 31957 9748
rect 32940 9852 32996 9872
rect 32940 9834 32959 9852
rect 32977 9834 32996 9852
rect 31646 9724 31701 9725
rect 31535 9713 31539 9718
rect 31496 9710 31539 9713
rect 31429 9696 31539 9710
rect 30855 9678 31196 9679
rect 29732 9657 29735 9677
rect 29755 9657 30148 9677
rect 30780 9677 31196 9678
rect 31646 9677 31689 9724
rect 32940 9721 32996 9834
rect 33148 9854 33162 9875
rect 33198 9854 33215 9875
rect 33426 9867 33457 9888
rect 33847 9867 33883 9888
rect 33269 9866 33306 9867
rect 33148 9847 33215 9854
rect 33268 9857 33306 9866
rect 30780 9673 31689 9677
rect 30099 9624 30144 9657
rect 30780 9653 30783 9673
rect 30803 9653 31689 9673
rect 31157 9648 31689 9653
rect 31897 9667 31956 9689
rect 31897 9649 31916 9667
rect 31934 9649 31956 9667
rect 30945 9624 31044 9626
rect 30099 9614 31044 9624
rect 30099 9588 30967 9614
rect 30100 9587 30967 9588
rect 30945 9576 30967 9587
rect 30992 9579 31011 9614
rect 31036 9579 31044 9614
rect 30992 9576 31044 9579
rect 31897 9578 31956 9649
rect 32940 9583 32995 9721
rect 33148 9695 33213 9847
rect 33268 9837 33277 9857
rect 33297 9837 33306 9857
rect 33268 9829 33306 9837
rect 33372 9861 33457 9867
rect 33482 9866 33519 9867
rect 33372 9841 33380 9861
rect 33400 9841 33457 9861
rect 33372 9833 33457 9841
rect 33481 9857 33519 9866
rect 33481 9837 33490 9857
rect 33510 9837 33519 9857
rect 33372 9832 33408 9833
rect 33481 9829 33519 9837
rect 33585 9861 33670 9867
rect 33690 9866 33727 9867
rect 33585 9841 33593 9861
rect 33613 9860 33670 9861
rect 33613 9841 33642 9860
rect 33585 9840 33642 9841
rect 33663 9840 33670 9860
rect 33585 9833 33670 9840
rect 33689 9857 33727 9866
rect 33689 9837 33698 9857
rect 33718 9837 33727 9857
rect 33585 9832 33621 9833
rect 33689 9829 33727 9837
rect 33793 9861 33937 9867
rect 33793 9841 33801 9861
rect 33821 9841 33909 9861
rect 33929 9841 33937 9861
rect 33793 9833 33937 9841
rect 33793 9832 33829 9833
rect 33901 9832 33937 9833
rect 34003 9866 34040 9867
rect 34003 9865 34041 9866
rect 34003 9857 34067 9865
rect 34003 9837 34012 9857
rect 34032 9843 34067 9857
rect 34087 9843 34090 9863
rect 34032 9838 34090 9843
rect 34032 9837 34067 9838
rect 33269 9800 33306 9829
rect 33270 9798 33306 9800
rect 33482 9798 33519 9829
rect 33270 9776 33519 9798
rect 33351 9770 33462 9776
rect 33351 9762 33392 9770
rect 33351 9742 33359 9762
rect 33378 9742 33392 9762
rect 33351 9740 33392 9742
rect 33420 9762 33462 9770
rect 33420 9742 33436 9762
rect 33455 9742 33462 9762
rect 33420 9740 33462 9742
rect 33351 9727 33462 9740
rect 33690 9730 33727 9829
rect 34003 9825 34067 9837
rect 33141 9685 33262 9695
rect 33141 9683 33210 9685
rect 33141 9642 33154 9683
rect 33191 9644 33210 9683
rect 33247 9644 33262 9685
rect 33191 9642 33262 9644
rect 33141 9624 33262 9642
rect 32933 9580 32997 9583
rect 33353 9580 33457 9586
rect 33688 9580 33729 9730
rect 34107 9722 34134 9977
rect 34196 9967 34276 9978
rect 34196 9941 34213 9967
rect 34253 9941 34276 9967
rect 34196 9914 34276 9941
rect 34196 9888 34217 9914
rect 34257 9888 34276 9914
rect 34196 9869 34276 9888
rect 34196 9843 34220 9869
rect 34260 9843 34276 9869
rect 34196 9792 34276 9843
rect 35299 9969 35377 10004
rect 35299 9907 35381 9969
rect 35299 9884 35327 9907
rect 35353 9884 35381 9907
rect 35299 9864 35381 9884
rect 30945 9568 31044 9576
rect 30971 9567 31043 9568
rect 30625 9541 30692 9560
rect 30625 9520 30642 9541
rect 29506 9342 29586 9384
rect 30623 9475 30642 9520
rect 30672 9520 30692 9541
rect 30672 9475 30693 9520
rect 31162 9517 31203 9519
rect 31434 9517 31538 9519
rect 31894 9517 31958 9578
rect 28567 9231 28603 9232
rect 28459 9223 28603 9231
rect 28459 9203 28467 9223
rect 28487 9203 28575 9223
rect 28595 9203 28603 9223
rect 28459 9197 28603 9203
rect 28669 9227 28707 9235
rect 28775 9231 28811 9232
rect 28669 9207 28678 9227
rect 28698 9207 28707 9227
rect 28669 9198 28707 9207
rect 28726 9224 28811 9231
rect 28726 9204 28733 9224
rect 28754 9223 28811 9224
rect 28754 9204 28783 9223
rect 28726 9203 28783 9204
rect 28803 9203 28811 9223
rect 28669 9197 28706 9198
rect 28726 9197 28811 9203
rect 28877 9227 28915 9235
rect 28988 9231 29024 9232
rect 28877 9207 28886 9227
rect 28906 9207 28915 9227
rect 28877 9198 28915 9207
rect 28939 9223 29024 9231
rect 28939 9203 28996 9223
rect 29016 9203 29024 9223
rect 28877 9197 28914 9198
rect 28939 9197 29024 9203
rect 29090 9227 29128 9235
rect 29090 9207 29099 9227
rect 29119 9207 29128 9227
rect 29090 9198 29128 9207
rect 29328 9215 29414 9251
rect 29090 9197 29127 9198
rect 28513 9176 28549 9197
rect 28939 9176 28970 9197
rect 29166 9176 29212 9180
rect 28346 9172 28446 9176
rect 28346 9168 28408 9172
rect 28346 9142 28353 9168
rect 28379 9146 28408 9168
rect 28434 9146 28446 9172
rect 28379 9142 28446 9146
rect 28346 9139 28446 9142
rect 28514 9139 28549 9176
rect 28611 9173 28970 9176
rect 28611 9168 28833 9173
rect 28611 9144 28624 9168
rect 28648 9149 28833 9168
rect 28857 9149 28970 9173
rect 28648 9144 28970 9149
rect 28611 9140 28970 9144
rect 29037 9168 29212 9176
rect 29037 9148 29048 9168
rect 29068 9148 29212 9168
rect 29328 9174 29345 9215
rect 29399 9174 29414 9215
rect 29328 9155 29414 9174
rect 29037 9141 29212 9148
rect 29037 9140 29078 9141
rect 28513 9114 28549 9139
rect 28361 9087 28398 9088
rect 28457 9087 28494 9088
rect 28513 9087 28520 9114
rect 28261 9078 28399 9087
rect 28261 9058 28370 9078
rect 28390 9058 28399 9078
rect 28261 9051 28399 9058
rect 28457 9084 28520 9087
rect 28541 9087 28549 9114
rect 28568 9087 28605 9088
rect 28541 9084 28605 9087
rect 28457 9078 28605 9084
rect 28457 9058 28466 9078
rect 28486 9058 28576 9078
rect 28596 9058 28605 9078
rect 28261 9049 28357 9051
rect 28457 9048 28605 9058
rect 28664 9078 28701 9088
rect 28776 9087 28813 9088
rect 28757 9085 28813 9087
rect 28664 9058 28672 9078
rect 28692 9058 28701 9078
rect 28513 9047 28549 9048
rect 28361 8916 28398 8917
rect 28664 8916 28701 9058
rect 28726 9078 28813 9085
rect 28726 9075 28784 9078
rect 28726 9055 28731 9075
rect 28752 9058 28784 9075
rect 28804 9058 28813 9078
rect 28752 9055 28813 9058
rect 28726 9048 28813 9055
rect 28872 9078 28909 9088
rect 28872 9058 28880 9078
rect 28900 9058 28909 9078
rect 28726 9047 28757 9048
rect 28872 8979 28909 9058
rect 28939 9087 28970 9140
rect 28989 9087 29026 9088
rect 28939 9078 29026 9087
rect 28939 9058 28997 9078
rect 29017 9058 29026 9078
rect 28939 9048 29026 9058
rect 29085 9078 29122 9088
rect 29085 9058 29093 9078
rect 29113 9058 29122 9078
rect 28939 9047 28970 9048
rect 28934 8979 29044 8992
rect 29085 8979 29122 9058
rect 29166 9058 29212 9141
rect 29506 9058 29581 9342
rect 30623 9267 30693 9475
rect 30755 9482 31958 9517
rect 30755 9468 30783 9482
rect 30757 9337 30783 9468
rect 31162 9479 31958 9482
rect 32933 9577 33729 9580
rect 34108 9591 34134 9722
rect 34108 9577 34136 9591
rect 32933 9542 34136 9577
rect 34198 9584 34268 9792
rect 32933 9481 32997 9542
rect 33353 9540 33457 9542
rect 33688 9540 33729 9542
rect 34198 9539 34219 9584
rect 34199 9518 34219 9539
rect 34249 9539 34268 9584
rect 34249 9518 34266 9539
rect 34199 9499 34266 9518
rect 33848 9491 33920 9492
rect 33847 9483 33946 9491
rect 30615 9216 30695 9267
rect 30615 9190 30631 9216
rect 30671 9190 30695 9216
rect 30615 9171 30695 9190
rect 30615 9145 30634 9171
rect 30674 9145 30695 9171
rect 30615 9118 30695 9145
rect 30615 9092 30638 9118
rect 30678 9092 30695 9118
rect 30615 9081 30695 9092
rect 30757 9082 30784 9337
rect 31162 9329 31203 9479
rect 31434 9473 31538 9479
rect 31894 9476 31958 9479
rect 31629 9417 31750 9435
rect 31629 9415 31700 9417
rect 31629 9374 31644 9415
rect 31681 9376 31700 9415
rect 31737 9376 31750 9417
rect 31681 9374 31750 9376
rect 31629 9364 31750 9374
rect 30824 9222 30888 9234
rect 31164 9230 31201 9329
rect 31429 9319 31540 9332
rect 31429 9317 31471 9319
rect 31429 9297 31436 9317
rect 31455 9297 31471 9317
rect 31429 9289 31471 9297
rect 31499 9317 31540 9319
rect 31499 9297 31513 9317
rect 31532 9297 31540 9317
rect 31499 9289 31540 9297
rect 31429 9283 31540 9289
rect 31372 9261 31621 9283
rect 31372 9230 31409 9261
rect 31585 9259 31621 9261
rect 31585 9230 31622 9259
rect 30824 9221 30859 9222
rect 30801 9216 30859 9221
rect 30801 9196 30804 9216
rect 30824 9202 30859 9216
rect 30879 9202 30888 9222
rect 30824 9194 30888 9202
rect 30850 9193 30888 9194
rect 30851 9192 30888 9193
rect 30954 9226 30990 9227
rect 31062 9226 31098 9227
rect 30954 9218 31098 9226
rect 30954 9198 30962 9218
rect 30982 9198 31070 9218
rect 31090 9198 31098 9218
rect 30954 9192 31098 9198
rect 31164 9222 31202 9230
rect 31270 9226 31306 9227
rect 31164 9202 31173 9222
rect 31193 9202 31202 9222
rect 31164 9193 31202 9202
rect 31221 9219 31306 9226
rect 31221 9199 31228 9219
rect 31249 9218 31306 9219
rect 31249 9199 31278 9218
rect 31221 9198 31278 9199
rect 31298 9198 31306 9218
rect 31164 9192 31201 9193
rect 31221 9192 31306 9198
rect 31372 9222 31410 9230
rect 31483 9226 31519 9227
rect 31372 9202 31381 9222
rect 31401 9202 31410 9222
rect 31372 9193 31410 9202
rect 31434 9218 31519 9226
rect 31434 9198 31491 9218
rect 31511 9198 31519 9218
rect 31372 9192 31409 9193
rect 31434 9192 31519 9198
rect 31585 9222 31623 9230
rect 31585 9202 31594 9222
rect 31614 9202 31623 9222
rect 31678 9212 31743 9364
rect 31896 9338 31951 9476
rect 32935 9410 32994 9481
rect 33847 9480 33899 9483
rect 33847 9445 33855 9480
rect 33880 9445 33899 9480
rect 33924 9472 33946 9483
rect 33924 9471 34791 9472
rect 33924 9445 34792 9471
rect 33847 9435 34792 9445
rect 33847 9433 33946 9435
rect 32935 9392 32957 9410
rect 32975 9392 32994 9410
rect 32935 9370 32994 9392
rect 33202 9406 33734 9411
rect 33202 9386 34088 9406
rect 34108 9386 34111 9406
rect 34747 9402 34792 9435
rect 33202 9382 34111 9386
rect 31585 9193 31623 9202
rect 31676 9205 31743 9212
rect 31585 9192 31622 9193
rect 31008 9171 31044 9192
rect 31434 9171 31465 9192
rect 31676 9184 31693 9205
rect 31729 9184 31743 9205
rect 31895 9225 31951 9338
rect 33202 9335 33245 9382
rect 33695 9381 34111 9382
rect 34743 9382 35136 9402
rect 35156 9382 35159 9402
rect 33695 9380 34036 9381
rect 33352 9349 33462 9363
rect 33352 9346 33395 9349
rect 33352 9341 33356 9346
rect 33190 9334 33245 9335
rect 31895 9207 31914 9225
rect 31932 9207 31951 9225
rect 31895 9187 31951 9207
rect 32934 9311 33245 9334
rect 32934 9293 32959 9311
rect 32977 9299 33245 9311
rect 33274 9319 33356 9341
rect 33385 9319 33395 9346
rect 33423 9322 33430 9349
rect 33459 9341 33462 9349
rect 33459 9322 33524 9341
rect 33423 9319 33524 9322
rect 33274 9317 33524 9319
rect 32977 9293 32999 9299
rect 31676 9171 31743 9184
rect 30841 9167 30941 9171
rect 30841 9163 30903 9167
rect 30841 9137 30848 9163
rect 30874 9141 30903 9163
rect 30929 9141 30941 9167
rect 30874 9137 30941 9141
rect 30841 9134 30941 9137
rect 31009 9134 31044 9171
rect 31106 9168 31465 9171
rect 31106 9163 31328 9168
rect 31106 9139 31119 9163
rect 31143 9144 31328 9163
rect 31352 9144 31465 9168
rect 31143 9139 31465 9144
rect 31106 9135 31465 9139
rect 31532 9165 31743 9171
rect 31532 9163 31693 9165
rect 31532 9143 31543 9163
rect 31563 9143 31693 9163
rect 31532 9136 31693 9143
rect 31532 9135 31573 9136
rect 31008 9109 31044 9134
rect 30856 9082 30893 9083
rect 30952 9082 30989 9083
rect 31008 9082 31015 9109
rect 29166 9023 29581 9058
rect 30756 9073 30894 9082
rect 30756 9053 30865 9073
rect 30885 9053 30894 9073
rect 30756 9046 30894 9053
rect 30952 9079 31015 9082
rect 31036 9082 31044 9109
rect 31063 9082 31100 9083
rect 31036 9079 31100 9082
rect 30952 9073 31100 9079
rect 30952 9053 30961 9073
rect 30981 9053 31071 9073
rect 31091 9053 31100 9073
rect 30756 9044 30852 9046
rect 30952 9043 31100 9053
rect 31159 9073 31196 9083
rect 31271 9082 31308 9083
rect 31252 9080 31308 9082
rect 31159 9053 31167 9073
rect 31187 9053 31196 9073
rect 31008 9042 31044 9043
rect 29166 9022 29212 9023
rect 28872 8977 29122 8979
rect 28872 8974 28973 8977
rect 28872 8955 28937 8974
rect 28934 8947 28937 8955
rect 28966 8947 28973 8974
rect 29001 8950 29011 8977
rect 29040 8955 29122 8977
rect 29506 8971 29581 9023
rect 29040 8950 29044 8955
rect 29001 8947 29044 8950
rect 28934 8933 29044 8947
rect 28360 8915 28701 8916
rect 28285 8910 28701 8915
rect 28285 8890 28288 8910
rect 28308 8890 28702 8910
rect 27342 8243 28148 8318
rect 26581 8199 26590 8233
rect 26619 8232 27029 8233
rect 26619 8199 26636 8232
rect 26861 8231 27029 8232
rect 26581 8173 26636 8199
rect 26581 8139 26589 8173
rect 26618 8139 26636 8173
rect 26581 8127 26636 8139
rect 24777 8082 24861 8103
rect 24777 8054 24805 8082
rect 24849 8054 24861 8082
rect 24591 8003 24665 8031
rect 24591 7955 24614 8003
rect 24651 7955 24665 8003
rect 24777 8025 24861 8054
rect 24777 7997 24802 8025
rect 24846 7997 24861 8025
rect 24777 7972 24861 7997
rect 26917 7986 27005 7990
rect 24591 7946 24665 7955
rect 19654 7869 19726 7891
rect 19787 7884 20990 7919
rect 19787 7870 19815 7884
rect 19655 7669 19725 7869
rect 19789 7739 19815 7870
rect 20194 7881 20990 7884
rect 19647 7618 19727 7669
rect 19647 7592 19663 7618
rect 19703 7592 19727 7618
rect 19647 7573 19727 7592
rect 19647 7547 19666 7573
rect 19706 7547 19727 7573
rect 19647 7520 19727 7547
rect 19647 7494 19670 7520
rect 19710 7494 19727 7520
rect 19647 7483 19727 7494
rect 19789 7484 19816 7739
rect 20194 7731 20235 7881
rect 20466 7879 20570 7881
rect 20925 7847 20990 7881
rect 22224 7896 22290 7944
rect 24601 7942 24665 7946
rect 26917 7969 27181 7986
rect 26917 7915 27097 7969
rect 27160 7915 27181 7969
rect 24814 7905 25525 7907
rect 24187 7904 25525 7905
rect 23137 7903 23209 7904
rect 20661 7819 20782 7837
rect 20661 7817 20732 7819
rect 20661 7776 20676 7817
rect 20713 7778 20732 7817
rect 20769 7778 20782 7819
rect 20713 7776 20782 7778
rect 20661 7766 20782 7776
rect 20466 7736 20570 7739
rect 19856 7624 19920 7636
rect 20196 7632 20233 7731
rect 20461 7721 20572 7736
rect 20461 7719 20503 7721
rect 20461 7699 20468 7719
rect 20487 7699 20503 7719
rect 20461 7691 20503 7699
rect 20531 7719 20572 7721
rect 20531 7699 20545 7719
rect 20564 7699 20572 7719
rect 20531 7691 20572 7699
rect 20461 7685 20572 7691
rect 20404 7663 20653 7685
rect 20404 7632 20441 7663
rect 20617 7661 20653 7663
rect 20617 7632 20654 7661
rect 19856 7623 19891 7624
rect 19833 7618 19891 7623
rect 19833 7598 19836 7618
rect 19856 7604 19891 7618
rect 19911 7604 19920 7624
rect 19856 7596 19920 7604
rect 19882 7595 19920 7596
rect 19883 7594 19920 7595
rect 19986 7628 20022 7629
rect 20094 7628 20130 7629
rect 19986 7620 20130 7628
rect 19986 7600 19994 7620
rect 20014 7600 20102 7620
rect 20122 7600 20130 7620
rect 19986 7594 20130 7600
rect 20196 7624 20234 7632
rect 20302 7628 20338 7629
rect 20196 7604 20205 7624
rect 20225 7604 20234 7624
rect 20196 7595 20234 7604
rect 20253 7621 20338 7628
rect 20253 7601 20260 7621
rect 20281 7620 20338 7621
rect 20281 7601 20310 7620
rect 20253 7600 20310 7601
rect 20330 7600 20338 7620
rect 20196 7594 20233 7595
rect 20253 7594 20338 7600
rect 20404 7624 20442 7632
rect 20515 7628 20551 7629
rect 20404 7604 20413 7624
rect 20433 7604 20442 7624
rect 20404 7595 20442 7604
rect 20466 7620 20551 7628
rect 20466 7600 20523 7620
rect 20543 7600 20551 7620
rect 20404 7594 20441 7595
rect 20466 7594 20551 7600
rect 20617 7624 20655 7632
rect 20617 7604 20626 7624
rect 20646 7604 20655 7624
rect 20710 7614 20775 7766
rect 20928 7740 20983 7847
rect 22224 7822 22283 7896
rect 23136 7895 23235 7903
rect 23136 7892 23188 7895
rect 23136 7857 23144 7892
rect 23169 7857 23188 7892
rect 23213 7884 23235 7895
rect 24186 7896 25525 7904
rect 24186 7893 24238 7896
rect 23213 7883 24080 7884
rect 23213 7857 24081 7883
rect 23136 7847 24081 7857
rect 23136 7845 23235 7847
rect 22224 7804 22246 7822
rect 22264 7804 22283 7822
rect 22224 7782 22283 7804
rect 22491 7818 23023 7823
rect 22491 7798 23377 7818
rect 23397 7798 23400 7818
rect 24036 7814 24081 7847
rect 24186 7858 24194 7893
rect 24219 7858 24238 7893
rect 24263 7858 25525 7896
rect 24186 7849 25525 7858
rect 24186 7846 24275 7849
rect 24814 7847 25525 7849
rect 26917 7898 27181 7915
rect 22491 7794 23400 7798
rect 22491 7747 22534 7794
rect 22984 7793 23400 7794
rect 24032 7794 24425 7814
rect 24445 7794 24448 7814
rect 22984 7792 23325 7793
rect 22641 7761 22751 7775
rect 22641 7758 22684 7761
rect 22641 7753 22645 7758
rect 22479 7746 22534 7747
rect 20617 7595 20655 7604
rect 20708 7607 20775 7614
rect 20617 7594 20654 7595
rect 20040 7573 20076 7594
rect 20466 7573 20497 7594
rect 20708 7586 20725 7607
rect 20761 7586 20775 7607
rect 20927 7627 20983 7740
rect 20927 7609 20946 7627
rect 20964 7609 20983 7627
rect 20927 7589 20983 7609
rect 22223 7723 22534 7746
rect 22223 7705 22248 7723
rect 22266 7711 22534 7723
rect 22563 7731 22645 7753
rect 22674 7731 22684 7758
rect 22712 7734 22719 7761
rect 22748 7753 22751 7761
rect 22748 7734 22813 7753
rect 22712 7731 22813 7734
rect 22563 7729 22813 7731
rect 22266 7705 22288 7711
rect 20708 7573 20775 7586
rect 19873 7569 19973 7573
rect 19873 7565 19935 7569
rect 19873 7539 19880 7565
rect 19906 7543 19935 7565
rect 19961 7543 19973 7569
rect 19906 7539 19973 7543
rect 19873 7536 19973 7539
rect 20041 7536 20076 7573
rect 20138 7570 20497 7573
rect 20138 7565 20360 7570
rect 20138 7541 20151 7565
rect 20175 7546 20360 7565
rect 20384 7546 20497 7570
rect 20175 7541 20497 7546
rect 20138 7537 20497 7541
rect 20564 7567 20775 7573
rect 20564 7565 20725 7567
rect 20564 7545 20575 7565
rect 20595 7545 20725 7565
rect 20564 7538 20725 7545
rect 20564 7537 20605 7538
rect 20040 7511 20076 7536
rect 19888 7484 19925 7485
rect 19984 7484 20021 7485
rect 20040 7484 20047 7511
rect 19788 7475 19926 7484
rect 19788 7455 19897 7475
rect 19917 7455 19926 7475
rect 19788 7448 19926 7455
rect 19984 7481 20047 7484
rect 20068 7484 20076 7511
rect 20095 7484 20132 7485
rect 20068 7481 20132 7484
rect 19984 7475 20132 7481
rect 19984 7455 19993 7475
rect 20013 7455 20103 7475
rect 20123 7455 20132 7475
rect 19788 7446 19884 7448
rect 19984 7445 20132 7455
rect 20191 7475 20228 7485
rect 20303 7484 20340 7485
rect 20284 7482 20340 7484
rect 20191 7455 20199 7475
rect 20219 7455 20228 7475
rect 20040 7444 20076 7445
rect 19888 7313 19925 7314
rect 20191 7313 20228 7455
rect 20253 7475 20340 7482
rect 20253 7472 20311 7475
rect 20253 7452 20258 7472
rect 20279 7455 20311 7472
rect 20331 7455 20340 7475
rect 20279 7452 20340 7455
rect 20253 7445 20340 7452
rect 20399 7475 20436 7485
rect 20399 7455 20407 7475
rect 20427 7455 20436 7475
rect 20253 7444 20284 7445
rect 20399 7376 20436 7455
rect 20466 7484 20497 7537
rect 20710 7530 20725 7538
rect 20765 7530 20775 7567
rect 22223 7566 22288 7705
rect 22563 7650 22600 7729
rect 22641 7716 22751 7729
rect 22715 7660 22746 7661
rect 22563 7630 22572 7650
rect 22592 7630 22600 7650
rect 20710 7521 20775 7530
rect 20923 7528 20988 7549
rect 22223 7548 22246 7566
rect 22264 7548 22288 7566
rect 22223 7531 22288 7548
rect 22443 7612 22511 7625
rect 22563 7620 22600 7630
rect 22659 7650 22746 7660
rect 22659 7630 22668 7650
rect 22688 7630 22746 7650
rect 22659 7621 22746 7630
rect 22659 7620 22696 7621
rect 22443 7570 22450 7612
rect 22499 7570 22511 7612
rect 22443 7567 22511 7570
rect 22715 7568 22746 7621
rect 22776 7650 22813 7729
rect 22928 7660 22959 7661
rect 22776 7630 22785 7650
rect 22805 7630 22813 7650
rect 22776 7620 22813 7630
rect 22872 7653 22959 7660
rect 22872 7650 22933 7653
rect 22872 7630 22881 7650
rect 22901 7633 22933 7650
rect 22954 7633 22959 7653
rect 22901 7630 22959 7633
rect 22872 7623 22959 7630
rect 22984 7650 23021 7792
rect 23287 7791 23324 7792
rect 24032 7789 24448 7794
rect 24032 7788 24373 7789
rect 23689 7757 23799 7771
rect 23689 7754 23732 7757
rect 23689 7749 23693 7754
rect 23611 7727 23693 7749
rect 23722 7727 23732 7754
rect 23760 7730 23767 7757
rect 23796 7749 23799 7757
rect 23796 7730 23861 7749
rect 23760 7727 23861 7730
rect 23611 7725 23861 7727
rect 23136 7660 23172 7661
rect 22984 7630 22993 7650
rect 23013 7630 23021 7650
rect 22872 7621 22928 7623
rect 22872 7620 22909 7621
rect 22984 7620 23021 7630
rect 23080 7650 23228 7660
rect 23328 7657 23424 7659
rect 23080 7630 23089 7650
rect 23109 7630 23199 7650
rect 23219 7630 23228 7650
rect 23080 7624 23228 7630
rect 23080 7621 23144 7624
rect 23080 7620 23117 7621
rect 23136 7594 23144 7621
rect 23165 7621 23228 7624
rect 23286 7650 23424 7657
rect 23286 7630 23295 7650
rect 23315 7630 23424 7650
rect 23286 7621 23424 7630
rect 23611 7646 23648 7725
rect 23689 7712 23799 7725
rect 23763 7656 23794 7657
rect 23611 7626 23620 7646
rect 23640 7626 23648 7646
rect 23165 7594 23172 7621
rect 23191 7620 23228 7621
rect 23287 7620 23324 7621
rect 23136 7569 23172 7594
rect 22607 7567 22648 7568
rect 22443 7560 22648 7567
rect 22443 7549 22617 7560
rect 20923 7510 20948 7528
rect 20966 7510 20988 7528
rect 22443 7516 22451 7549
rect 20516 7484 20553 7485
rect 20466 7475 20553 7484
rect 20466 7455 20524 7475
rect 20544 7455 20553 7475
rect 20466 7445 20553 7455
rect 20612 7475 20649 7485
rect 20612 7455 20620 7475
rect 20640 7455 20649 7475
rect 20466 7444 20497 7445
rect 20461 7376 20571 7389
rect 20612 7376 20649 7455
rect 20923 7434 20988 7510
rect 22444 7507 22451 7516
rect 22500 7540 22617 7549
rect 22637 7540 22648 7560
rect 22500 7532 22648 7540
rect 22715 7564 23074 7568
rect 22715 7559 23037 7564
rect 22715 7535 22828 7559
rect 22852 7540 23037 7559
rect 23061 7540 23074 7564
rect 22852 7535 23074 7540
rect 22715 7532 23074 7535
rect 23136 7532 23171 7569
rect 23239 7566 23339 7569
rect 23239 7562 23306 7566
rect 23239 7536 23251 7562
rect 23277 7540 23306 7562
rect 23332 7540 23339 7566
rect 23277 7536 23339 7540
rect 23239 7532 23339 7536
rect 22500 7516 22511 7532
rect 22500 7507 22508 7516
rect 22715 7511 22746 7532
rect 23136 7511 23172 7532
rect 22558 7510 22595 7511
rect 22223 7467 22288 7486
rect 22223 7449 22248 7467
rect 22266 7449 22288 7467
rect 20399 7374 20649 7376
rect 20399 7371 20500 7374
rect 20399 7352 20464 7371
rect 20461 7344 20464 7352
rect 20493 7344 20500 7371
rect 20528 7347 20538 7374
rect 20567 7352 20649 7374
rect 20672 7399 20989 7434
rect 20567 7347 20571 7352
rect 20528 7344 20571 7347
rect 20461 7330 20571 7344
rect 19887 7312 20228 7313
rect 19812 7310 20228 7312
rect 20672 7310 20712 7399
rect 20923 7372 20988 7399
rect 20923 7354 20946 7372
rect 20964 7354 20988 7372
rect 20923 7334 20988 7354
rect 19809 7307 20712 7310
rect 19809 7287 19815 7307
rect 19835 7287 20712 7307
rect 19809 7283 20712 7287
rect 20672 7280 20712 7283
rect 20924 7273 20989 7294
rect 19142 7265 19803 7266
rect 19142 7258 20076 7265
rect 19142 7257 20048 7258
rect 19142 7237 19993 7257
rect 20025 7238 20048 7257
rect 20073 7238 20076 7258
rect 20025 7237 20076 7238
rect 19142 7230 20076 7237
rect 18741 7188 18909 7189
rect 19144 7188 19183 7230
rect 19972 7228 20076 7230
rect 20041 7226 20076 7228
rect 20924 7255 20948 7273
rect 20966 7255 20989 7273
rect 20924 7208 20989 7255
rect 18741 7162 19185 7188
rect 18741 7160 18909 7162
rect 18741 6809 18768 7160
rect 19144 7156 19185 7162
rect 18808 6949 18872 6961
rect 19148 6957 19185 7156
rect 19647 7183 19719 7200
rect 19647 7144 19655 7183
rect 19700 7144 19719 7183
rect 19413 7046 19524 7061
rect 19413 7044 19455 7046
rect 19413 7024 19420 7044
rect 19439 7024 19455 7044
rect 19413 7016 19455 7024
rect 19483 7044 19524 7046
rect 19483 7024 19497 7044
rect 19516 7024 19524 7044
rect 19483 7016 19524 7024
rect 19413 7010 19524 7016
rect 19356 6988 19605 7010
rect 19356 6957 19393 6988
rect 19569 6986 19605 6988
rect 19569 6957 19606 6986
rect 18808 6948 18843 6949
rect 18785 6943 18843 6948
rect 18785 6923 18788 6943
rect 18808 6929 18843 6943
rect 18863 6929 18872 6949
rect 18808 6921 18872 6929
rect 18834 6920 18872 6921
rect 18835 6919 18872 6920
rect 18938 6953 18974 6954
rect 19046 6953 19082 6954
rect 18938 6945 19082 6953
rect 18938 6925 18946 6945
rect 18966 6925 19054 6945
rect 19074 6925 19082 6945
rect 18938 6919 19082 6925
rect 19148 6949 19186 6957
rect 19254 6953 19290 6954
rect 19148 6929 19157 6949
rect 19177 6929 19186 6949
rect 19148 6920 19186 6929
rect 19205 6946 19290 6953
rect 19205 6926 19212 6946
rect 19233 6945 19290 6946
rect 19233 6926 19262 6945
rect 19205 6925 19262 6926
rect 19282 6925 19290 6945
rect 19148 6919 19185 6920
rect 19205 6919 19290 6925
rect 19356 6949 19394 6957
rect 19467 6953 19503 6954
rect 19356 6929 19365 6949
rect 19385 6929 19394 6949
rect 19356 6920 19394 6929
rect 19418 6945 19503 6953
rect 19418 6925 19475 6945
rect 19495 6925 19503 6945
rect 19356 6919 19393 6920
rect 19418 6919 19503 6925
rect 19569 6949 19607 6957
rect 19569 6929 19578 6949
rect 19598 6929 19607 6949
rect 19569 6920 19607 6929
rect 19647 6934 19719 7144
rect 19789 7178 20989 7208
rect 19789 7177 20233 7178
rect 19789 7175 19957 7177
rect 19647 6920 19730 6934
rect 19569 6919 19606 6920
rect 18992 6898 19028 6919
rect 19418 6898 19449 6919
rect 19647 6898 19664 6920
rect 18825 6894 18925 6898
rect 18825 6890 18887 6894
rect 18825 6864 18832 6890
rect 18858 6868 18887 6890
rect 18913 6868 18925 6894
rect 18858 6864 18925 6868
rect 18825 6861 18925 6864
rect 18993 6861 19028 6898
rect 19090 6895 19449 6898
rect 19090 6890 19312 6895
rect 19090 6866 19103 6890
rect 19127 6871 19312 6890
rect 19336 6871 19449 6895
rect 19127 6866 19449 6871
rect 19090 6862 19449 6866
rect 19516 6890 19664 6898
rect 19516 6870 19527 6890
rect 19547 6887 19664 6890
rect 19717 6887 19730 6920
rect 19547 6870 19730 6887
rect 19516 6863 19730 6870
rect 19516 6862 19557 6863
rect 19647 6862 19730 6863
rect 18992 6836 19028 6861
rect 18840 6809 18877 6810
rect 18936 6809 18973 6810
rect 18992 6809 18999 6836
rect 18740 6800 18878 6809
rect 18740 6780 18849 6800
rect 18869 6780 18878 6800
rect 18740 6773 18878 6780
rect 18936 6806 18999 6809
rect 19020 6809 19028 6836
rect 19047 6809 19084 6810
rect 19020 6806 19084 6809
rect 18936 6800 19084 6806
rect 18936 6780 18945 6800
rect 18965 6780 19055 6800
rect 19075 6780 19084 6800
rect 18740 6771 18836 6773
rect 18936 6770 19084 6780
rect 19143 6800 19180 6810
rect 19255 6809 19292 6810
rect 19236 6807 19292 6809
rect 19143 6780 19151 6800
rect 19171 6780 19180 6800
rect 18992 6769 19028 6770
rect 18840 6638 18877 6639
rect 19143 6638 19180 6780
rect 19205 6800 19292 6807
rect 19205 6797 19263 6800
rect 19205 6777 19210 6797
rect 19231 6780 19263 6797
rect 19283 6780 19292 6800
rect 19231 6777 19292 6780
rect 19205 6770 19292 6777
rect 19351 6800 19388 6810
rect 19351 6780 19359 6800
rect 19379 6780 19388 6800
rect 19205 6769 19236 6770
rect 19351 6701 19388 6780
rect 19418 6809 19449 6862
rect 19655 6829 19669 6862
rect 19722 6829 19730 6862
rect 19655 6823 19730 6829
rect 19655 6818 19725 6823
rect 19468 6809 19505 6810
rect 19418 6800 19505 6809
rect 19418 6780 19476 6800
rect 19496 6780 19505 6800
rect 19418 6770 19505 6780
rect 19564 6800 19601 6810
rect 19789 6805 19816 7175
rect 19856 6945 19920 6957
rect 20196 6953 20233 7177
rect 20704 7158 20768 7160
rect 20700 7146 20768 7158
rect 20700 7113 20711 7146
rect 20751 7113 20768 7146
rect 20700 7103 20768 7113
rect 20461 7042 20572 7057
rect 20461 7040 20503 7042
rect 20461 7020 20468 7040
rect 20487 7020 20503 7040
rect 20461 7012 20503 7020
rect 20531 7040 20572 7042
rect 20531 7020 20545 7040
rect 20564 7020 20572 7040
rect 20531 7012 20572 7020
rect 20461 7006 20572 7012
rect 20404 6984 20653 7006
rect 20404 6953 20441 6984
rect 20617 6982 20653 6984
rect 20617 6953 20654 6982
rect 19856 6944 19891 6945
rect 19833 6939 19891 6944
rect 19833 6919 19836 6939
rect 19856 6925 19891 6939
rect 19911 6925 19920 6945
rect 19856 6917 19920 6925
rect 19882 6916 19920 6917
rect 19883 6915 19920 6916
rect 19986 6949 20022 6950
rect 20094 6949 20130 6950
rect 19986 6941 20130 6949
rect 19986 6921 19994 6941
rect 20014 6921 20102 6941
rect 20122 6921 20130 6941
rect 19986 6915 20130 6921
rect 20196 6945 20234 6953
rect 20302 6949 20338 6950
rect 20196 6925 20205 6945
rect 20225 6925 20234 6945
rect 20196 6916 20234 6925
rect 20253 6942 20338 6949
rect 20253 6922 20260 6942
rect 20281 6941 20338 6942
rect 20281 6922 20310 6941
rect 20253 6921 20310 6922
rect 20330 6921 20338 6941
rect 20196 6915 20233 6916
rect 20253 6915 20338 6921
rect 20404 6945 20442 6953
rect 20515 6949 20551 6950
rect 20404 6925 20413 6945
rect 20433 6925 20442 6945
rect 20404 6916 20442 6925
rect 20466 6941 20551 6949
rect 20466 6921 20523 6941
rect 20543 6921 20551 6941
rect 20404 6915 20441 6916
rect 20466 6915 20551 6921
rect 20617 6945 20655 6953
rect 20617 6925 20626 6945
rect 20646 6925 20655 6945
rect 20617 6916 20655 6925
rect 20704 6919 20768 7103
rect 20924 6977 20989 7178
rect 22223 7248 22288 7449
rect 22444 7323 22508 7507
rect 22557 7501 22595 7510
rect 22557 7481 22566 7501
rect 22586 7481 22595 7501
rect 22557 7473 22595 7481
rect 22661 7505 22746 7511
rect 22771 7510 22808 7511
rect 22661 7485 22669 7505
rect 22689 7485 22746 7505
rect 22661 7477 22746 7485
rect 22770 7501 22808 7510
rect 22770 7481 22779 7501
rect 22799 7481 22808 7501
rect 22661 7476 22697 7477
rect 22770 7473 22808 7481
rect 22874 7505 22959 7511
rect 22979 7510 23016 7511
rect 22874 7485 22882 7505
rect 22902 7504 22959 7505
rect 22902 7485 22931 7504
rect 22874 7484 22931 7485
rect 22952 7484 22959 7504
rect 22874 7477 22959 7484
rect 22978 7501 23016 7510
rect 22978 7481 22987 7501
rect 23007 7481 23016 7501
rect 22874 7476 22910 7477
rect 22978 7473 23016 7481
rect 23082 7505 23226 7511
rect 23082 7485 23090 7505
rect 23110 7485 23198 7505
rect 23218 7485 23226 7505
rect 23082 7477 23226 7485
rect 23082 7476 23118 7477
rect 23190 7476 23226 7477
rect 23292 7510 23329 7511
rect 23292 7509 23330 7510
rect 23292 7501 23356 7509
rect 23292 7481 23301 7501
rect 23321 7487 23356 7501
rect 23376 7487 23379 7507
rect 23321 7482 23379 7487
rect 23321 7481 23356 7482
rect 22558 7444 22595 7473
rect 22559 7442 22595 7444
rect 22771 7442 22808 7473
rect 22559 7420 22808 7442
rect 22640 7414 22751 7420
rect 22640 7406 22681 7414
rect 22640 7386 22648 7406
rect 22667 7386 22681 7406
rect 22640 7384 22681 7386
rect 22709 7406 22751 7414
rect 22709 7386 22725 7406
rect 22744 7386 22751 7406
rect 22709 7384 22751 7386
rect 22640 7369 22751 7384
rect 22444 7313 22512 7323
rect 22444 7280 22461 7313
rect 22501 7280 22512 7313
rect 22444 7268 22512 7280
rect 22444 7266 22508 7268
rect 22979 7249 23016 7473
rect 23292 7469 23356 7481
rect 23396 7251 23423 7621
rect 23611 7616 23648 7626
rect 23707 7646 23794 7656
rect 23707 7626 23716 7646
rect 23736 7626 23794 7646
rect 23707 7617 23794 7626
rect 23707 7616 23744 7617
rect 23487 7603 23557 7608
rect 23482 7597 23557 7603
rect 23482 7564 23490 7597
rect 23543 7564 23557 7597
rect 23763 7564 23794 7617
rect 23824 7646 23861 7725
rect 23976 7656 24007 7657
rect 23824 7626 23833 7646
rect 23853 7626 23861 7646
rect 23824 7616 23861 7626
rect 23920 7649 24007 7656
rect 23920 7646 23981 7649
rect 23920 7626 23929 7646
rect 23949 7629 23981 7646
rect 24002 7629 24007 7649
rect 23949 7626 24007 7629
rect 23920 7619 24007 7626
rect 24032 7646 24069 7788
rect 24335 7787 24372 7788
rect 24184 7656 24220 7657
rect 24032 7626 24041 7646
rect 24061 7626 24069 7646
rect 23920 7617 23976 7619
rect 23920 7616 23957 7617
rect 24032 7616 24069 7626
rect 24128 7646 24276 7656
rect 24376 7653 24472 7655
rect 24128 7626 24137 7646
rect 24157 7626 24247 7646
rect 24267 7626 24276 7646
rect 24128 7620 24276 7626
rect 24128 7617 24192 7620
rect 24128 7616 24165 7617
rect 24184 7590 24192 7617
rect 24213 7617 24276 7620
rect 24334 7646 24472 7653
rect 24334 7626 24343 7646
rect 24363 7626 24472 7646
rect 24334 7617 24472 7626
rect 24213 7590 24220 7617
rect 24239 7616 24276 7617
rect 24335 7616 24372 7617
rect 24184 7565 24220 7590
rect 23482 7563 23565 7564
rect 23655 7563 23696 7564
rect 23482 7556 23696 7563
rect 23482 7539 23665 7556
rect 23482 7506 23495 7539
rect 23548 7536 23665 7539
rect 23685 7536 23696 7556
rect 23548 7528 23696 7536
rect 23763 7560 24122 7564
rect 23763 7555 24085 7560
rect 23763 7531 23876 7555
rect 23900 7536 24085 7555
rect 24109 7536 24122 7560
rect 23900 7531 24122 7536
rect 23763 7528 24122 7531
rect 24184 7528 24219 7565
rect 24287 7562 24387 7565
rect 24287 7558 24354 7562
rect 24287 7532 24299 7558
rect 24325 7536 24354 7558
rect 24380 7536 24387 7562
rect 24325 7532 24387 7536
rect 24287 7528 24387 7532
rect 23548 7506 23565 7528
rect 23763 7507 23794 7528
rect 24184 7507 24220 7528
rect 23606 7506 23643 7507
rect 23482 7492 23565 7506
rect 23255 7249 23423 7251
rect 22979 7248 23423 7249
rect 22223 7218 23423 7248
rect 23493 7282 23565 7492
rect 23605 7497 23643 7506
rect 23605 7477 23614 7497
rect 23634 7477 23643 7497
rect 23605 7469 23643 7477
rect 23709 7501 23794 7507
rect 23819 7506 23856 7507
rect 23709 7481 23717 7501
rect 23737 7481 23794 7501
rect 23709 7473 23794 7481
rect 23818 7497 23856 7506
rect 23818 7477 23827 7497
rect 23847 7477 23856 7497
rect 23709 7472 23745 7473
rect 23818 7469 23856 7477
rect 23922 7501 24007 7507
rect 24027 7506 24064 7507
rect 23922 7481 23930 7501
rect 23950 7500 24007 7501
rect 23950 7481 23979 7500
rect 23922 7480 23979 7481
rect 24000 7480 24007 7500
rect 23922 7473 24007 7480
rect 24026 7497 24064 7506
rect 24026 7477 24035 7497
rect 24055 7477 24064 7497
rect 23922 7472 23958 7473
rect 24026 7469 24064 7477
rect 24130 7501 24274 7507
rect 24130 7481 24138 7501
rect 24158 7481 24246 7501
rect 24266 7481 24274 7501
rect 24130 7473 24274 7481
rect 24130 7472 24166 7473
rect 24238 7472 24274 7473
rect 24340 7506 24377 7507
rect 24340 7505 24378 7506
rect 24340 7497 24404 7505
rect 24340 7477 24349 7497
rect 24369 7483 24404 7497
rect 24424 7483 24427 7503
rect 24369 7478 24427 7483
rect 24369 7477 24404 7478
rect 23606 7440 23643 7469
rect 23607 7438 23643 7440
rect 23819 7438 23856 7469
rect 23607 7416 23856 7438
rect 23688 7410 23799 7416
rect 23688 7402 23729 7410
rect 23688 7382 23696 7402
rect 23715 7382 23729 7402
rect 23688 7380 23729 7382
rect 23757 7402 23799 7410
rect 23757 7382 23773 7402
rect 23792 7382 23799 7402
rect 23757 7380 23799 7382
rect 23688 7365 23799 7380
rect 23493 7243 23512 7282
rect 23557 7243 23565 7282
rect 23493 7226 23565 7243
rect 24027 7270 24064 7469
rect 24340 7465 24404 7477
rect 24027 7264 24068 7270
rect 24444 7266 24471 7617
rect 24766 7604 24861 7630
rect 24602 7582 24666 7601
rect 24602 7543 24615 7582
rect 24649 7543 24666 7582
rect 24602 7524 24666 7543
rect 24303 7264 24471 7266
rect 24027 7238 24471 7264
rect 22223 7171 22288 7218
rect 22223 7153 22246 7171
rect 22264 7153 22288 7171
rect 23136 7198 23171 7200
rect 23136 7196 23240 7198
rect 24029 7196 24068 7238
rect 24303 7237 24471 7238
rect 23136 7189 24070 7196
rect 23136 7188 23187 7189
rect 23136 7168 23139 7188
rect 23164 7169 23187 7188
rect 23219 7169 24070 7189
rect 23164 7168 24070 7169
rect 23136 7161 24070 7168
rect 23409 7160 24070 7161
rect 22223 7132 22288 7153
rect 22500 7143 22540 7146
rect 22500 7139 23403 7143
rect 22500 7119 23377 7139
rect 23397 7119 23403 7139
rect 22500 7116 23403 7119
rect 22224 7072 22289 7092
rect 22224 7054 22248 7072
rect 22266 7054 22289 7072
rect 22224 7027 22289 7054
rect 22500 7027 22540 7116
rect 22984 7114 23400 7116
rect 22984 7113 23325 7114
rect 22641 7082 22751 7096
rect 22641 7079 22684 7082
rect 22641 7074 22645 7079
rect 22223 6992 22540 7027
rect 22563 7052 22645 7074
rect 22674 7052 22684 7079
rect 22712 7055 22719 7082
rect 22748 7074 22751 7082
rect 22748 7055 22813 7074
rect 22712 7052 22813 7055
rect 22563 7050 22813 7052
rect 20924 6959 20946 6977
rect 20964 6959 20989 6977
rect 20924 6940 20989 6959
rect 20617 6915 20654 6916
rect 20040 6894 20076 6915
rect 20466 6894 20497 6915
rect 20704 6910 20712 6919
rect 20701 6894 20712 6910
rect 19873 6890 19973 6894
rect 19873 6886 19935 6890
rect 19873 6860 19880 6886
rect 19906 6864 19935 6886
rect 19961 6864 19973 6890
rect 19906 6860 19973 6864
rect 19873 6857 19973 6860
rect 20041 6857 20076 6894
rect 20138 6891 20497 6894
rect 20138 6886 20360 6891
rect 20138 6862 20151 6886
rect 20175 6867 20360 6886
rect 20384 6867 20497 6891
rect 20175 6862 20497 6867
rect 20138 6858 20497 6862
rect 20564 6886 20712 6894
rect 20564 6866 20575 6886
rect 20595 6877 20712 6886
rect 20761 6910 20768 6919
rect 22224 6916 22289 6992
rect 22563 6971 22600 7050
rect 22641 7037 22751 7050
rect 22715 6981 22746 6982
rect 22563 6951 22572 6971
rect 22592 6951 22600 6971
rect 22563 6941 22600 6951
rect 22659 6971 22746 6981
rect 22659 6951 22668 6971
rect 22688 6951 22746 6971
rect 22659 6942 22746 6951
rect 22659 6941 22696 6942
rect 20761 6877 20769 6910
rect 22224 6898 22246 6916
rect 22264 6898 22289 6916
rect 20595 6866 20769 6877
rect 20564 6859 20769 6866
rect 20564 6858 20605 6859
rect 20040 6832 20076 6857
rect 19888 6805 19925 6806
rect 19984 6805 20021 6806
rect 20040 6805 20047 6832
rect 19564 6780 19572 6800
rect 19592 6780 19601 6800
rect 19418 6769 19449 6770
rect 19413 6701 19523 6714
rect 19564 6701 19601 6780
rect 19788 6796 19926 6805
rect 19788 6776 19897 6796
rect 19917 6776 19926 6796
rect 19788 6769 19926 6776
rect 19984 6802 20047 6805
rect 20068 6805 20076 6832
rect 20095 6805 20132 6806
rect 20068 6802 20132 6805
rect 19984 6796 20132 6802
rect 19984 6776 19993 6796
rect 20013 6776 20103 6796
rect 20123 6776 20132 6796
rect 19788 6767 19884 6769
rect 19984 6766 20132 6776
rect 20191 6796 20228 6806
rect 20303 6805 20340 6806
rect 20284 6803 20340 6805
rect 20191 6776 20199 6796
rect 20219 6776 20228 6796
rect 20040 6765 20076 6766
rect 19351 6699 19601 6701
rect 19351 6696 19452 6699
rect 19351 6677 19416 6696
rect 19413 6669 19416 6677
rect 19445 6669 19452 6696
rect 19480 6672 19490 6699
rect 19519 6677 19601 6699
rect 19519 6672 19523 6677
rect 19480 6669 19523 6672
rect 19413 6655 19523 6669
rect 18839 6637 19180 6638
rect 18764 6632 19180 6637
rect 19888 6634 19925 6635
rect 20191 6634 20228 6776
rect 20253 6796 20340 6803
rect 20253 6793 20311 6796
rect 20253 6773 20258 6793
rect 20279 6776 20311 6793
rect 20331 6776 20340 6796
rect 20279 6773 20340 6776
rect 20253 6766 20340 6773
rect 20399 6796 20436 6806
rect 20399 6776 20407 6796
rect 20427 6776 20436 6796
rect 20253 6765 20284 6766
rect 20399 6697 20436 6776
rect 20466 6805 20497 6858
rect 20701 6856 20769 6859
rect 20701 6814 20713 6856
rect 20762 6814 20769 6856
rect 20516 6805 20553 6806
rect 20466 6796 20553 6805
rect 20466 6776 20524 6796
rect 20544 6776 20553 6796
rect 20466 6766 20553 6776
rect 20612 6796 20649 6806
rect 20701 6801 20769 6814
rect 20924 6878 20989 6895
rect 20924 6860 20948 6878
rect 20966 6860 20989 6878
rect 22224 6877 22289 6898
rect 22437 6896 22502 6905
rect 20612 6776 20620 6796
rect 20640 6776 20649 6796
rect 20466 6765 20497 6766
rect 20461 6697 20571 6710
rect 20612 6697 20649 6776
rect 20924 6721 20989 6860
rect 22437 6859 22447 6896
rect 22487 6888 22502 6896
rect 22715 6889 22746 6942
rect 22776 6971 22813 7050
rect 22928 6981 22959 6982
rect 22776 6951 22785 6971
rect 22805 6951 22813 6971
rect 22776 6941 22813 6951
rect 22872 6974 22959 6981
rect 22872 6971 22933 6974
rect 22872 6951 22881 6971
rect 22901 6954 22933 6971
rect 22954 6954 22959 6974
rect 22901 6951 22959 6954
rect 22872 6944 22959 6951
rect 22984 6971 23021 7113
rect 23287 7112 23324 7113
rect 24604 7053 24666 7524
rect 24766 7563 24792 7604
rect 24828 7563 24861 7604
rect 24766 7267 24861 7563
rect 24766 7223 24781 7267
rect 24841 7223 24861 7267
rect 24766 7203 24861 7223
rect 25478 7134 25521 7847
rect 25478 7114 25872 7134
rect 25892 7114 25895 7134
rect 25479 7109 25895 7114
rect 25479 7108 25820 7109
rect 25136 7077 25246 7091
rect 25136 7074 25179 7077
rect 25136 7069 25140 7074
rect 24599 7001 24674 7053
rect 25058 7047 25140 7069
rect 25169 7047 25179 7074
rect 25207 7050 25214 7077
rect 25243 7069 25246 7077
rect 25243 7050 25308 7069
rect 25207 7047 25308 7050
rect 25058 7045 25308 7047
rect 24968 7001 25014 7002
rect 23136 6981 23172 6982
rect 22984 6951 22993 6971
rect 23013 6951 23021 6971
rect 22872 6942 22928 6944
rect 22872 6941 22909 6942
rect 22984 6941 23021 6951
rect 23080 6971 23228 6981
rect 23328 6978 23424 6980
rect 23080 6951 23089 6971
rect 23109 6951 23199 6971
rect 23219 6951 23228 6971
rect 23080 6945 23228 6951
rect 23080 6942 23144 6945
rect 23080 6941 23117 6942
rect 23136 6915 23144 6942
rect 23165 6942 23228 6945
rect 23286 6971 23424 6978
rect 23286 6951 23295 6971
rect 23315 6951 23424 6971
rect 23286 6942 23424 6951
rect 24599 6966 25014 7001
rect 23165 6915 23172 6942
rect 23191 6941 23228 6942
rect 23287 6941 23324 6942
rect 23136 6890 23172 6915
rect 22607 6888 22648 6889
rect 22487 6881 22648 6888
rect 22487 6861 22617 6881
rect 22637 6861 22648 6881
rect 22487 6859 22648 6861
rect 22437 6853 22648 6859
rect 22715 6885 23074 6889
rect 22715 6880 23037 6885
rect 22715 6856 22828 6880
rect 22852 6861 23037 6880
rect 23061 6861 23074 6885
rect 22852 6856 23074 6861
rect 22715 6853 23074 6856
rect 23136 6853 23171 6890
rect 23239 6887 23339 6890
rect 23239 6883 23306 6887
rect 23239 6857 23251 6883
rect 23277 6861 23306 6883
rect 23332 6861 23339 6887
rect 23277 6857 23339 6861
rect 23239 6853 23339 6857
rect 22437 6840 22504 6853
rect 20924 6715 20946 6721
rect 20399 6695 20649 6697
rect 20399 6692 20500 6695
rect 20399 6673 20464 6692
rect 20461 6665 20464 6673
rect 20493 6665 20500 6692
rect 20528 6668 20538 6695
rect 20567 6673 20649 6695
rect 20678 6703 20946 6715
rect 20964 6703 20989 6721
rect 20678 6680 20989 6703
rect 22229 6817 22285 6837
rect 22229 6799 22248 6817
rect 22266 6799 22285 6817
rect 22229 6686 22285 6799
rect 22437 6819 22451 6840
rect 22487 6819 22504 6840
rect 22715 6832 22746 6853
rect 23136 6832 23172 6853
rect 22558 6831 22595 6832
rect 22437 6812 22504 6819
rect 22557 6822 22595 6831
rect 20678 6679 20733 6680
rect 20567 6668 20571 6673
rect 20528 6665 20571 6668
rect 20461 6651 20571 6665
rect 19887 6633 20228 6634
rect 18764 6612 18767 6632
rect 18787 6612 19180 6632
rect 19812 6632 20228 6633
rect 20678 6632 20721 6679
rect 19812 6628 20721 6632
rect 19131 6579 19176 6612
rect 19812 6608 19815 6628
rect 19835 6608 20721 6628
rect 20189 6603 20721 6608
rect 20929 6622 20988 6644
rect 20929 6604 20948 6622
rect 20966 6604 20988 6622
rect 19977 6579 20076 6581
rect 19131 6569 20076 6579
rect 19131 6543 19999 6569
rect 19132 6542 19999 6543
rect 19977 6531 19999 6542
rect 20024 6534 20043 6569
rect 20068 6534 20076 6569
rect 20024 6531 20076 6534
rect 20929 6533 20988 6604
rect 22229 6548 22284 6686
rect 22437 6660 22502 6812
rect 22557 6802 22566 6822
rect 22586 6802 22595 6822
rect 22557 6794 22595 6802
rect 22661 6826 22746 6832
rect 22771 6831 22808 6832
rect 22661 6806 22669 6826
rect 22689 6806 22746 6826
rect 22661 6798 22746 6806
rect 22770 6822 22808 6831
rect 22770 6802 22779 6822
rect 22799 6802 22808 6822
rect 22661 6797 22697 6798
rect 22770 6794 22808 6802
rect 22874 6826 22959 6832
rect 22979 6831 23016 6832
rect 22874 6806 22882 6826
rect 22902 6825 22959 6826
rect 22902 6806 22931 6825
rect 22874 6805 22931 6806
rect 22952 6805 22959 6825
rect 22874 6798 22959 6805
rect 22978 6822 23016 6831
rect 22978 6802 22987 6822
rect 23007 6802 23016 6822
rect 22874 6797 22910 6798
rect 22978 6794 23016 6802
rect 23082 6826 23226 6832
rect 23082 6806 23090 6826
rect 23110 6806 23198 6826
rect 23218 6806 23226 6826
rect 23082 6798 23226 6806
rect 23082 6797 23118 6798
rect 23190 6797 23226 6798
rect 23292 6831 23329 6832
rect 23292 6830 23330 6831
rect 23292 6822 23356 6830
rect 23292 6802 23301 6822
rect 23321 6808 23356 6822
rect 23376 6808 23379 6828
rect 23321 6803 23379 6808
rect 23321 6802 23356 6803
rect 22558 6765 22595 6794
rect 22559 6763 22595 6765
rect 22771 6763 22808 6794
rect 22559 6741 22808 6763
rect 22640 6735 22751 6741
rect 22640 6727 22681 6735
rect 22640 6707 22648 6727
rect 22667 6707 22681 6727
rect 22640 6705 22681 6707
rect 22709 6727 22751 6735
rect 22709 6707 22725 6727
rect 22744 6707 22751 6727
rect 22709 6705 22751 6707
rect 22640 6692 22751 6705
rect 22979 6695 23016 6794
rect 23292 6790 23356 6802
rect 22430 6650 22551 6660
rect 22430 6648 22499 6650
rect 22430 6607 22443 6648
rect 22480 6609 22499 6648
rect 22536 6609 22551 6650
rect 22480 6607 22551 6609
rect 22430 6589 22551 6607
rect 22222 6545 22286 6548
rect 22642 6545 22746 6551
rect 22977 6545 23018 6695
rect 23396 6687 23423 6942
rect 23485 6932 23565 6943
rect 23485 6906 23502 6932
rect 23542 6906 23565 6932
rect 23485 6879 23565 6906
rect 23485 6853 23506 6879
rect 23546 6853 23565 6879
rect 23485 6834 23565 6853
rect 23485 6808 23509 6834
rect 23549 6808 23565 6834
rect 23485 6757 23565 6808
rect 22222 6542 23018 6545
rect 23397 6556 23423 6687
rect 23397 6542 23425 6556
rect 19977 6523 20076 6531
rect 20003 6522 20075 6523
rect 19657 6496 19724 6515
rect 19657 6475 19674 6496
rect 19655 6430 19674 6475
rect 19704 6475 19724 6496
rect 19704 6430 19725 6475
rect 20194 6472 20235 6474
rect 20466 6472 20570 6474
rect 20926 6472 20990 6533
rect 19655 6222 19725 6430
rect 19787 6437 20990 6472
rect 22222 6507 23425 6542
rect 23487 6549 23557 6757
rect 24599 6682 24674 6966
rect 24968 6883 25014 6966
rect 25058 6966 25095 7045
rect 25136 7032 25246 7045
rect 25210 6976 25241 6977
rect 25058 6946 25067 6966
rect 25087 6946 25095 6966
rect 25058 6936 25095 6946
rect 25154 6966 25241 6976
rect 25154 6946 25163 6966
rect 25183 6946 25241 6966
rect 25154 6937 25241 6946
rect 25154 6936 25191 6937
rect 25210 6884 25241 6937
rect 25271 6966 25308 7045
rect 25423 6976 25454 6977
rect 25271 6946 25280 6966
rect 25300 6946 25308 6966
rect 25271 6936 25308 6946
rect 25367 6969 25454 6976
rect 25367 6966 25428 6969
rect 25367 6946 25376 6966
rect 25396 6949 25428 6966
rect 25449 6949 25454 6969
rect 25396 6946 25454 6949
rect 25367 6939 25454 6946
rect 25479 6966 25516 7108
rect 25782 7107 25819 7108
rect 25631 6976 25667 6977
rect 25479 6946 25488 6966
rect 25508 6946 25516 6966
rect 25367 6937 25423 6939
rect 25367 6936 25404 6937
rect 25479 6936 25516 6946
rect 25575 6966 25723 6976
rect 25823 6973 25919 6975
rect 25575 6946 25584 6966
rect 25604 6946 25694 6966
rect 25714 6946 25723 6966
rect 25575 6940 25723 6946
rect 25575 6937 25639 6940
rect 25575 6936 25612 6937
rect 25631 6910 25639 6937
rect 25660 6937 25723 6940
rect 25781 6966 25919 6973
rect 25781 6946 25790 6966
rect 25810 6946 25919 6966
rect 25781 6937 25919 6946
rect 25660 6910 25667 6937
rect 25686 6936 25723 6937
rect 25782 6936 25819 6937
rect 25631 6885 25667 6910
rect 25102 6883 25143 6884
rect 24968 6876 25143 6883
rect 24766 6850 24852 6869
rect 24766 6809 24781 6850
rect 24835 6809 24852 6850
rect 24968 6856 25112 6876
rect 25132 6856 25143 6876
rect 24968 6848 25143 6856
rect 25210 6880 25569 6884
rect 25210 6875 25532 6880
rect 25210 6851 25323 6875
rect 25347 6856 25532 6875
rect 25556 6856 25569 6880
rect 25347 6851 25569 6856
rect 25210 6848 25569 6851
rect 25631 6848 25666 6885
rect 25734 6882 25834 6885
rect 25734 6878 25801 6882
rect 25734 6852 25746 6878
rect 25772 6856 25801 6878
rect 25827 6856 25834 6882
rect 25772 6852 25834 6856
rect 25734 6848 25834 6852
rect 24968 6844 25014 6848
rect 25210 6827 25241 6848
rect 25631 6827 25667 6848
rect 25053 6826 25090 6827
rect 24766 6773 24852 6809
rect 25052 6817 25090 6826
rect 25052 6797 25061 6817
rect 25081 6797 25090 6817
rect 25052 6789 25090 6797
rect 25156 6821 25241 6827
rect 25266 6826 25303 6827
rect 25156 6801 25164 6821
rect 25184 6801 25241 6821
rect 25156 6793 25241 6801
rect 25265 6817 25303 6826
rect 25265 6797 25274 6817
rect 25294 6797 25303 6817
rect 25156 6792 25192 6793
rect 25265 6789 25303 6797
rect 25369 6821 25454 6827
rect 25474 6826 25511 6827
rect 25369 6801 25377 6821
rect 25397 6820 25454 6821
rect 25397 6801 25426 6820
rect 25369 6800 25426 6801
rect 25447 6800 25454 6820
rect 25369 6793 25454 6800
rect 25473 6817 25511 6826
rect 25473 6797 25482 6817
rect 25502 6797 25511 6817
rect 25369 6792 25405 6793
rect 25473 6789 25511 6797
rect 25577 6821 25721 6827
rect 25577 6801 25585 6821
rect 25605 6801 25693 6821
rect 25713 6801 25721 6821
rect 25577 6793 25721 6801
rect 25577 6792 25613 6793
rect 22222 6446 22286 6507
rect 22642 6505 22746 6507
rect 22977 6505 23018 6507
rect 23487 6504 23508 6549
rect 23488 6483 23508 6504
rect 23538 6504 23557 6549
rect 24594 6640 24674 6682
rect 23538 6483 23555 6504
rect 23488 6464 23555 6483
rect 23137 6456 23209 6457
rect 23136 6448 23235 6456
rect 19787 6423 19815 6437
rect 19789 6292 19815 6423
rect 20194 6434 20990 6437
rect 18542 6130 18624 6150
rect 18542 6107 18570 6130
rect 18596 6107 18624 6130
rect 18542 6045 18624 6107
rect 18546 6010 18624 6045
rect 19647 6171 19727 6222
rect 19647 6145 19663 6171
rect 19703 6145 19727 6171
rect 19647 6126 19727 6145
rect 19647 6100 19666 6126
rect 19706 6100 19727 6126
rect 19647 6073 19727 6100
rect 19647 6047 19670 6073
rect 19710 6047 19727 6073
rect 19647 6036 19727 6047
rect 19789 6037 19816 6292
rect 20194 6284 20235 6434
rect 20466 6428 20570 6434
rect 20926 6431 20990 6434
rect 20661 6372 20782 6390
rect 20661 6370 20732 6372
rect 20661 6329 20676 6370
rect 20713 6331 20732 6370
rect 20769 6331 20782 6372
rect 20713 6329 20782 6331
rect 20661 6319 20782 6329
rect 19856 6177 19920 6189
rect 20196 6185 20233 6284
rect 20461 6274 20572 6287
rect 20461 6272 20503 6274
rect 20461 6252 20468 6272
rect 20487 6252 20503 6272
rect 20461 6244 20503 6252
rect 20531 6272 20572 6274
rect 20531 6252 20545 6272
rect 20564 6252 20572 6272
rect 20531 6244 20572 6252
rect 20461 6238 20572 6244
rect 20404 6216 20653 6238
rect 20404 6185 20441 6216
rect 20617 6214 20653 6216
rect 20617 6185 20654 6214
rect 19856 6176 19891 6177
rect 19833 6171 19891 6176
rect 19833 6151 19836 6171
rect 19856 6157 19891 6171
rect 19911 6157 19920 6177
rect 19856 6149 19920 6157
rect 19882 6148 19920 6149
rect 19883 6147 19920 6148
rect 19986 6181 20022 6182
rect 20094 6181 20130 6182
rect 19986 6173 20130 6181
rect 19986 6153 19994 6173
rect 20014 6153 20102 6173
rect 20122 6153 20130 6173
rect 19986 6147 20130 6153
rect 20196 6177 20234 6185
rect 20302 6181 20338 6182
rect 20196 6157 20205 6177
rect 20225 6157 20234 6177
rect 20196 6148 20234 6157
rect 20253 6174 20338 6181
rect 20253 6154 20260 6174
rect 20281 6173 20338 6174
rect 20281 6154 20310 6173
rect 20253 6153 20310 6154
rect 20330 6153 20338 6173
rect 20196 6147 20233 6148
rect 20253 6147 20338 6153
rect 20404 6177 20442 6185
rect 20515 6181 20551 6182
rect 20404 6157 20413 6177
rect 20433 6157 20442 6177
rect 20404 6148 20442 6157
rect 20466 6173 20551 6181
rect 20466 6153 20523 6173
rect 20543 6153 20551 6173
rect 20404 6147 20441 6148
rect 20466 6147 20551 6153
rect 20617 6177 20655 6185
rect 20617 6157 20626 6177
rect 20646 6157 20655 6177
rect 20710 6167 20775 6319
rect 20928 6293 20983 6431
rect 22224 6375 22283 6446
rect 23136 6445 23188 6448
rect 23136 6410 23144 6445
rect 23169 6410 23188 6445
rect 23213 6437 23235 6448
rect 23213 6436 24080 6437
rect 23213 6410 24081 6436
rect 23136 6400 24081 6410
rect 23136 6398 23235 6400
rect 22224 6357 22246 6375
rect 22264 6357 22283 6375
rect 22224 6335 22283 6357
rect 22491 6371 23023 6376
rect 22491 6351 23377 6371
rect 23397 6351 23400 6371
rect 24036 6367 24081 6400
rect 22491 6347 23400 6351
rect 22491 6300 22534 6347
rect 22984 6346 23400 6347
rect 24032 6347 24425 6367
rect 24445 6347 24448 6367
rect 22984 6345 23325 6346
rect 22641 6314 22751 6328
rect 22641 6311 22684 6314
rect 22641 6306 22645 6311
rect 22479 6299 22534 6300
rect 20617 6148 20655 6157
rect 20708 6160 20775 6167
rect 20617 6147 20654 6148
rect 20040 6126 20076 6147
rect 20466 6126 20497 6147
rect 20708 6139 20725 6160
rect 20761 6139 20775 6160
rect 20927 6180 20983 6293
rect 20927 6162 20946 6180
rect 20964 6162 20983 6180
rect 20927 6142 20983 6162
rect 22223 6276 22534 6299
rect 22223 6258 22248 6276
rect 22266 6264 22534 6276
rect 22563 6284 22645 6306
rect 22674 6284 22684 6311
rect 22712 6287 22719 6314
rect 22748 6306 22751 6314
rect 22748 6287 22813 6306
rect 22712 6284 22813 6287
rect 22563 6282 22813 6284
rect 22266 6258 22288 6264
rect 20708 6126 20775 6139
rect 19873 6122 19973 6126
rect 19873 6118 19935 6122
rect 19873 6092 19880 6118
rect 19906 6096 19935 6118
rect 19961 6096 19973 6122
rect 19906 6092 19973 6096
rect 19873 6089 19973 6092
rect 20041 6089 20076 6126
rect 20138 6123 20497 6126
rect 20138 6118 20360 6123
rect 20138 6094 20151 6118
rect 20175 6099 20360 6118
rect 20384 6099 20497 6123
rect 20175 6094 20497 6099
rect 20138 6090 20497 6094
rect 20564 6120 20775 6126
rect 20564 6118 20725 6120
rect 20564 6098 20575 6118
rect 20595 6098 20725 6118
rect 20564 6091 20725 6098
rect 20564 6090 20605 6091
rect 20040 6064 20076 6089
rect 19888 6037 19925 6038
rect 19984 6037 20021 6038
rect 20040 6037 20047 6064
rect 19788 6028 19926 6037
rect 18546 5494 18608 6010
rect 19788 6008 19897 6028
rect 19917 6008 19926 6028
rect 19788 6001 19926 6008
rect 19984 6034 20047 6037
rect 20068 6037 20076 6064
rect 20095 6037 20132 6038
rect 20068 6034 20132 6037
rect 19984 6028 20132 6034
rect 19984 6008 19993 6028
rect 20013 6008 20103 6028
rect 20123 6008 20132 6028
rect 19788 5999 19884 6001
rect 19984 5998 20132 6008
rect 20191 6028 20228 6038
rect 20303 6037 20340 6038
rect 20284 6035 20340 6037
rect 20191 6008 20199 6028
rect 20219 6008 20228 6028
rect 20040 5997 20076 5998
rect 19888 5866 19925 5867
rect 20191 5866 20228 6008
rect 20253 6028 20340 6035
rect 20253 6025 20311 6028
rect 20253 6005 20258 6025
rect 20279 6008 20311 6025
rect 20331 6008 20340 6028
rect 20279 6005 20340 6008
rect 20253 5998 20340 6005
rect 20399 6028 20436 6038
rect 20399 6008 20407 6028
rect 20427 6008 20436 6028
rect 20253 5997 20284 5998
rect 20399 5929 20436 6008
rect 20466 6037 20497 6090
rect 20710 6083 20725 6091
rect 20765 6083 20775 6120
rect 22223 6119 22288 6258
rect 22563 6203 22600 6282
rect 22641 6269 22751 6282
rect 22715 6213 22746 6214
rect 22563 6183 22572 6203
rect 22592 6183 22600 6203
rect 20710 6074 20775 6083
rect 20923 6081 20988 6102
rect 22223 6101 22246 6119
rect 22264 6101 22288 6119
rect 22223 6084 22288 6101
rect 22443 6165 22511 6178
rect 22563 6173 22600 6183
rect 22659 6203 22746 6213
rect 22659 6183 22668 6203
rect 22688 6183 22746 6203
rect 22659 6174 22746 6183
rect 22659 6173 22696 6174
rect 22443 6123 22450 6165
rect 22499 6123 22511 6165
rect 22443 6120 22511 6123
rect 22715 6121 22746 6174
rect 22776 6203 22813 6282
rect 22928 6213 22959 6214
rect 22776 6183 22785 6203
rect 22805 6183 22813 6203
rect 22776 6173 22813 6183
rect 22872 6206 22959 6213
rect 22872 6203 22933 6206
rect 22872 6183 22881 6203
rect 22901 6186 22933 6203
rect 22954 6186 22959 6206
rect 22901 6183 22959 6186
rect 22872 6176 22959 6183
rect 22984 6203 23021 6345
rect 23287 6344 23324 6345
rect 24032 6342 24448 6347
rect 24032 6341 24373 6342
rect 23689 6310 23799 6324
rect 23689 6307 23732 6310
rect 23689 6302 23693 6307
rect 23611 6280 23693 6302
rect 23722 6280 23732 6307
rect 23760 6283 23767 6310
rect 23796 6302 23799 6310
rect 23796 6283 23861 6302
rect 23760 6280 23861 6283
rect 23611 6278 23861 6280
rect 23136 6213 23172 6214
rect 22984 6183 22993 6203
rect 23013 6183 23021 6203
rect 22872 6174 22928 6176
rect 22872 6173 22909 6174
rect 22984 6173 23021 6183
rect 23080 6203 23228 6213
rect 23328 6210 23424 6212
rect 23080 6183 23089 6203
rect 23109 6183 23199 6203
rect 23219 6183 23228 6203
rect 23080 6177 23228 6183
rect 23080 6174 23144 6177
rect 23080 6173 23117 6174
rect 23136 6147 23144 6174
rect 23165 6174 23228 6177
rect 23286 6203 23424 6210
rect 23286 6183 23295 6203
rect 23315 6183 23424 6203
rect 23286 6174 23424 6183
rect 23611 6199 23648 6278
rect 23689 6265 23799 6278
rect 23763 6209 23794 6210
rect 23611 6179 23620 6199
rect 23640 6179 23648 6199
rect 23165 6147 23172 6174
rect 23191 6173 23228 6174
rect 23287 6173 23324 6174
rect 23136 6122 23172 6147
rect 22607 6120 22648 6121
rect 22443 6113 22648 6120
rect 22443 6102 22617 6113
rect 20923 6063 20948 6081
rect 20966 6063 20988 6081
rect 22443 6069 22451 6102
rect 20516 6037 20553 6038
rect 20466 6028 20553 6037
rect 20466 6008 20524 6028
rect 20544 6008 20553 6028
rect 20466 5998 20553 6008
rect 20612 6028 20649 6038
rect 20612 6008 20620 6028
rect 20640 6008 20649 6028
rect 20466 5997 20497 5998
rect 20461 5929 20571 5942
rect 20612 5929 20649 6008
rect 20923 5987 20988 6063
rect 22444 6060 22451 6069
rect 22500 6093 22617 6102
rect 22637 6093 22648 6113
rect 22500 6085 22648 6093
rect 22715 6117 23074 6121
rect 22715 6112 23037 6117
rect 22715 6088 22828 6112
rect 22852 6093 23037 6112
rect 23061 6093 23074 6117
rect 22852 6088 23074 6093
rect 22715 6085 23074 6088
rect 23136 6085 23171 6122
rect 23239 6119 23339 6122
rect 23239 6115 23306 6119
rect 23239 6089 23251 6115
rect 23277 6093 23306 6115
rect 23332 6093 23339 6119
rect 23277 6089 23339 6093
rect 23239 6085 23339 6089
rect 22500 6069 22511 6085
rect 22500 6060 22508 6069
rect 22715 6064 22746 6085
rect 23136 6064 23172 6085
rect 22558 6063 22595 6064
rect 22223 6020 22288 6039
rect 22223 6002 22248 6020
rect 22266 6002 22288 6020
rect 20399 5927 20649 5929
rect 20399 5924 20500 5927
rect 20399 5905 20464 5924
rect 20461 5897 20464 5905
rect 20493 5897 20500 5924
rect 20528 5900 20538 5927
rect 20567 5905 20649 5927
rect 20672 5952 20989 5987
rect 20567 5900 20571 5905
rect 20528 5897 20571 5900
rect 20461 5883 20571 5897
rect 19887 5865 20228 5866
rect 19812 5863 20228 5865
rect 20672 5863 20712 5952
rect 20923 5925 20988 5952
rect 20923 5907 20946 5925
rect 20964 5907 20988 5925
rect 20923 5887 20988 5907
rect 19809 5860 20712 5863
rect 19809 5840 19815 5860
rect 19835 5840 20712 5860
rect 19809 5836 20712 5840
rect 20672 5833 20712 5836
rect 20924 5826 20989 5847
rect 19142 5818 19803 5819
rect 19142 5811 20076 5818
rect 19142 5810 20048 5811
rect 19142 5790 19993 5810
rect 20025 5791 20048 5810
rect 20073 5791 20076 5811
rect 20025 5790 20076 5791
rect 19142 5783 20076 5790
rect 18741 5741 18909 5742
rect 19144 5741 19183 5783
rect 19972 5781 20076 5783
rect 20041 5779 20076 5781
rect 20924 5808 20948 5826
rect 20966 5808 20989 5826
rect 20924 5761 20989 5808
rect 18741 5715 19185 5741
rect 18741 5713 18909 5715
rect 18543 5410 18612 5494
rect 18541 4931 18612 5410
rect 18741 5362 18768 5713
rect 19144 5709 19185 5715
rect 18808 5502 18872 5514
rect 19148 5510 19185 5709
rect 19647 5736 19719 5753
rect 19647 5697 19655 5736
rect 19700 5697 19719 5736
rect 19413 5599 19524 5614
rect 19413 5597 19455 5599
rect 19413 5577 19420 5597
rect 19439 5577 19455 5597
rect 19413 5569 19455 5577
rect 19483 5597 19524 5599
rect 19483 5577 19497 5597
rect 19516 5577 19524 5597
rect 19483 5569 19524 5577
rect 19413 5563 19524 5569
rect 19356 5541 19605 5563
rect 19356 5510 19393 5541
rect 19569 5539 19605 5541
rect 19569 5510 19606 5539
rect 18808 5501 18843 5502
rect 18785 5496 18843 5501
rect 18785 5476 18788 5496
rect 18808 5482 18843 5496
rect 18863 5482 18872 5502
rect 18808 5474 18872 5482
rect 18834 5473 18872 5474
rect 18835 5472 18872 5473
rect 18938 5506 18974 5507
rect 19046 5506 19082 5507
rect 18938 5498 19082 5506
rect 18938 5478 18946 5498
rect 18966 5478 19054 5498
rect 19074 5478 19082 5498
rect 18938 5472 19082 5478
rect 19148 5502 19186 5510
rect 19254 5506 19290 5507
rect 19148 5482 19157 5502
rect 19177 5482 19186 5502
rect 19148 5473 19186 5482
rect 19205 5499 19290 5506
rect 19205 5479 19212 5499
rect 19233 5498 19290 5499
rect 19233 5479 19262 5498
rect 19205 5478 19262 5479
rect 19282 5478 19290 5498
rect 19148 5472 19185 5473
rect 19205 5472 19290 5478
rect 19356 5502 19394 5510
rect 19467 5506 19503 5507
rect 19356 5482 19365 5502
rect 19385 5482 19394 5502
rect 19356 5473 19394 5482
rect 19418 5498 19503 5506
rect 19418 5478 19475 5498
rect 19495 5478 19503 5498
rect 19356 5472 19393 5473
rect 19418 5472 19503 5478
rect 19569 5502 19607 5510
rect 19569 5482 19578 5502
rect 19598 5482 19607 5502
rect 19569 5473 19607 5482
rect 19647 5487 19719 5697
rect 19789 5731 20989 5761
rect 19789 5730 20233 5731
rect 19789 5728 19957 5730
rect 19647 5473 19730 5487
rect 19569 5472 19606 5473
rect 18992 5451 19028 5472
rect 19418 5451 19449 5472
rect 19647 5451 19664 5473
rect 18825 5447 18925 5451
rect 18825 5443 18887 5447
rect 18825 5417 18832 5443
rect 18858 5421 18887 5443
rect 18913 5421 18925 5447
rect 18858 5417 18925 5421
rect 18825 5414 18925 5417
rect 18993 5414 19028 5451
rect 19090 5448 19449 5451
rect 19090 5443 19312 5448
rect 19090 5419 19103 5443
rect 19127 5424 19312 5443
rect 19336 5424 19449 5448
rect 19127 5419 19449 5424
rect 19090 5415 19449 5419
rect 19516 5443 19664 5451
rect 19516 5423 19527 5443
rect 19547 5440 19664 5443
rect 19717 5440 19730 5473
rect 19547 5423 19730 5440
rect 19516 5416 19730 5423
rect 19516 5415 19557 5416
rect 19647 5415 19730 5416
rect 18992 5389 19028 5414
rect 18840 5362 18877 5363
rect 18936 5362 18973 5363
rect 18992 5362 18999 5389
rect 18740 5353 18878 5362
rect 18740 5333 18849 5353
rect 18869 5333 18878 5353
rect 18740 5326 18878 5333
rect 18936 5359 18999 5362
rect 19020 5362 19028 5389
rect 19047 5362 19084 5363
rect 19020 5359 19084 5362
rect 18936 5353 19084 5359
rect 18936 5333 18945 5353
rect 18965 5333 19055 5353
rect 19075 5333 19084 5353
rect 18740 5324 18836 5326
rect 18936 5323 19084 5333
rect 19143 5353 19180 5363
rect 19255 5362 19292 5363
rect 19236 5360 19292 5362
rect 19143 5333 19151 5353
rect 19171 5333 19180 5353
rect 18992 5322 19028 5323
rect 18840 5191 18877 5192
rect 19143 5191 19180 5333
rect 19205 5353 19292 5360
rect 19205 5350 19263 5353
rect 19205 5330 19210 5350
rect 19231 5333 19263 5350
rect 19283 5333 19292 5353
rect 19231 5330 19292 5333
rect 19205 5323 19292 5330
rect 19351 5353 19388 5363
rect 19351 5333 19359 5353
rect 19379 5333 19388 5353
rect 19205 5322 19236 5323
rect 19351 5254 19388 5333
rect 19418 5362 19449 5415
rect 19655 5382 19669 5415
rect 19722 5382 19730 5415
rect 19655 5376 19730 5382
rect 19655 5371 19725 5376
rect 19468 5362 19505 5363
rect 19418 5353 19505 5362
rect 19418 5333 19476 5353
rect 19496 5333 19505 5353
rect 19418 5323 19505 5333
rect 19564 5353 19601 5363
rect 19789 5358 19816 5728
rect 19856 5498 19920 5510
rect 20196 5506 20233 5730
rect 20704 5711 20768 5713
rect 20700 5699 20768 5711
rect 20700 5666 20711 5699
rect 20751 5666 20768 5699
rect 20700 5656 20768 5666
rect 20461 5595 20572 5610
rect 20461 5593 20503 5595
rect 20461 5573 20468 5593
rect 20487 5573 20503 5593
rect 20461 5565 20503 5573
rect 20531 5593 20572 5595
rect 20531 5573 20545 5593
rect 20564 5573 20572 5593
rect 20531 5565 20572 5573
rect 20461 5559 20572 5565
rect 20404 5537 20653 5559
rect 20404 5506 20441 5537
rect 20617 5535 20653 5537
rect 20617 5506 20654 5535
rect 19856 5497 19891 5498
rect 19833 5492 19891 5497
rect 19833 5472 19836 5492
rect 19856 5478 19891 5492
rect 19911 5478 19920 5498
rect 19856 5470 19920 5478
rect 19882 5469 19920 5470
rect 19883 5468 19920 5469
rect 19986 5502 20022 5503
rect 20094 5502 20130 5503
rect 19986 5494 20130 5502
rect 19986 5474 19994 5494
rect 20014 5474 20102 5494
rect 20122 5474 20130 5494
rect 19986 5468 20130 5474
rect 20196 5498 20234 5506
rect 20302 5502 20338 5503
rect 20196 5478 20205 5498
rect 20225 5478 20234 5498
rect 20196 5469 20234 5478
rect 20253 5495 20338 5502
rect 20253 5475 20260 5495
rect 20281 5494 20338 5495
rect 20281 5475 20310 5494
rect 20253 5474 20310 5475
rect 20330 5474 20338 5494
rect 20196 5468 20233 5469
rect 20253 5468 20338 5474
rect 20404 5498 20442 5506
rect 20515 5502 20551 5503
rect 20404 5478 20413 5498
rect 20433 5478 20442 5498
rect 20404 5469 20442 5478
rect 20466 5494 20551 5502
rect 20466 5474 20523 5494
rect 20543 5474 20551 5494
rect 20404 5468 20441 5469
rect 20466 5468 20551 5474
rect 20617 5498 20655 5506
rect 20617 5478 20626 5498
rect 20646 5478 20655 5498
rect 20617 5469 20655 5478
rect 20704 5472 20768 5656
rect 20924 5530 20989 5731
rect 22223 5801 22288 6002
rect 22444 5876 22508 6060
rect 22557 6054 22595 6063
rect 22557 6034 22566 6054
rect 22586 6034 22595 6054
rect 22557 6026 22595 6034
rect 22661 6058 22746 6064
rect 22771 6063 22808 6064
rect 22661 6038 22669 6058
rect 22689 6038 22746 6058
rect 22661 6030 22746 6038
rect 22770 6054 22808 6063
rect 22770 6034 22779 6054
rect 22799 6034 22808 6054
rect 22661 6029 22697 6030
rect 22770 6026 22808 6034
rect 22874 6058 22959 6064
rect 22979 6063 23016 6064
rect 22874 6038 22882 6058
rect 22902 6057 22959 6058
rect 22902 6038 22931 6057
rect 22874 6037 22931 6038
rect 22952 6037 22959 6057
rect 22874 6030 22959 6037
rect 22978 6054 23016 6063
rect 22978 6034 22987 6054
rect 23007 6034 23016 6054
rect 22874 6029 22910 6030
rect 22978 6026 23016 6034
rect 23082 6058 23226 6064
rect 23082 6038 23090 6058
rect 23110 6038 23198 6058
rect 23218 6038 23226 6058
rect 23082 6030 23226 6038
rect 23082 6029 23118 6030
rect 23190 6029 23226 6030
rect 23292 6063 23329 6064
rect 23292 6062 23330 6063
rect 23292 6054 23356 6062
rect 23292 6034 23301 6054
rect 23321 6040 23356 6054
rect 23376 6040 23379 6060
rect 23321 6035 23379 6040
rect 23321 6034 23356 6035
rect 22558 5997 22595 6026
rect 22559 5995 22595 5997
rect 22771 5995 22808 6026
rect 22559 5973 22808 5995
rect 22640 5967 22751 5973
rect 22640 5959 22681 5967
rect 22640 5939 22648 5959
rect 22667 5939 22681 5959
rect 22640 5937 22681 5939
rect 22709 5959 22751 5967
rect 22709 5939 22725 5959
rect 22744 5939 22751 5959
rect 22709 5937 22751 5939
rect 22640 5922 22751 5937
rect 22444 5866 22512 5876
rect 22444 5833 22461 5866
rect 22501 5833 22512 5866
rect 22444 5821 22512 5833
rect 22444 5819 22508 5821
rect 22979 5802 23016 6026
rect 23292 6022 23356 6034
rect 23396 5804 23423 6174
rect 23611 6169 23648 6179
rect 23707 6199 23794 6209
rect 23707 6179 23716 6199
rect 23736 6179 23794 6199
rect 23707 6170 23794 6179
rect 23707 6169 23744 6170
rect 23487 6156 23557 6161
rect 23482 6150 23557 6156
rect 23482 6117 23490 6150
rect 23543 6117 23557 6150
rect 23763 6117 23794 6170
rect 23824 6199 23861 6278
rect 23976 6209 24007 6210
rect 23824 6179 23833 6199
rect 23853 6179 23861 6199
rect 23824 6169 23861 6179
rect 23920 6202 24007 6209
rect 23920 6199 23981 6202
rect 23920 6179 23929 6199
rect 23949 6182 23981 6199
rect 24002 6182 24007 6202
rect 23949 6179 24007 6182
rect 23920 6172 24007 6179
rect 24032 6199 24069 6341
rect 24335 6340 24372 6341
rect 24184 6209 24220 6210
rect 24032 6179 24041 6199
rect 24061 6179 24069 6199
rect 23920 6170 23976 6172
rect 23920 6169 23957 6170
rect 24032 6169 24069 6179
rect 24128 6199 24276 6209
rect 24376 6206 24472 6208
rect 24128 6179 24137 6199
rect 24157 6179 24247 6199
rect 24267 6179 24276 6199
rect 24128 6173 24276 6179
rect 24128 6170 24192 6173
rect 24128 6169 24165 6170
rect 24184 6143 24192 6170
rect 24213 6170 24276 6173
rect 24334 6199 24472 6206
rect 24334 6179 24343 6199
rect 24363 6179 24472 6199
rect 24334 6170 24472 6179
rect 24213 6143 24220 6170
rect 24239 6169 24276 6170
rect 24335 6169 24372 6170
rect 24184 6118 24220 6143
rect 23482 6116 23565 6117
rect 23655 6116 23696 6117
rect 23482 6109 23696 6116
rect 23482 6092 23665 6109
rect 23482 6059 23495 6092
rect 23548 6089 23665 6092
rect 23685 6089 23696 6109
rect 23548 6081 23696 6089
rect 23763 6113 24122 6117
rect 23763 6108 24085 6113
rect 23763 6084 23876 6108
rect 23900 6089 24085 6108
rect 24109 6089 24122 6113
rect 23900 6084 24122 6089
rect 23763 6081 24122 6084
rect 24184 6081 24219 6118
rect 24287 6115 24387 6118
rect 24287 6111 24354 6115
rect 24287 6085 24299 6111
rect 24325 6089 24354 6111
rect 24380 6089 24387 6115
rect 24325 6085 24387 6089
rect 24287 6081 24387 6085
rect 23548 6059 23565 6081
rect 23763 6060 23794 6081
rect 24184 6060 24220 6081
rect 23606 6059 23643 6060
rect 23482 6045 23565 6059
rect 23255 5802 23423 5804
rect 22979 5801 23423 5802
rect 22223 5771 23423 5801
rect 23493 5835 23565 6045
rect 23605 6050 23643 6059
rect 23605 6030 23614 6050
rect 23634 6030 23643 6050
rect 23605 6022 23643 6030
rect 23709 6054 23794 6060
rect 23819 6059 23856 6060
rect 23709 6034 23717 6054
rect 23737 6034 23794 6054
rect 23709 6026 23794 6034
rect 23818 6050 23856 6059
rect 23818 6030 23827 6050
rect 23847 6030 23856 6050
rect 23709 6025 23745 6026
rect 23818 6022 23856 6030
rect 23922 6054 24007 6060
rect 24027 6059 24064 6060
rect 23922 6034 23930 6054
rect 23950 6053 24007 6054
rect 23950 6034 23979 6053
rect 23922 6033 23979 6034
rect 24000 6033 24007 6053
rect 23922 6026 24007 6033
rect 24026 6050 24064 6059
rect 24026 6030 24035 6050
rect 24055 6030 24064 6050
rect 23922 6025 23958 6026
rect 24026 6022 24064 6030
rect 24130 6054 24274 6060
rect 24130 6034 24138 6054
rect 24158 6034 24246 6054
rect 24266 6034 24274 6054
rect 24130 6026 24274 6034
rect 24130 6025 24166 6026
rect 24238 6025 24274 6026
rect 24340 6059 24377 6060
rect 24340 6058 24378 6059
rect 24340 6050 24404 6058
rect 24340 6030 24349 6050
rect 24369 6036 24404 6050
rect 24424 6036 24427 6056
rect 24369 6031 24427 6036
rect 24369 6030 24404 6031
rect 23606 5993 23643 6022
rect 23607 5991 23643 5993
rect 23819 5991 23856 6022
rect 23607 5969 23856 5991
rect 23688 5963 23799 5969
rect 23688 5955 23729 5963
rect 23688 5935 23696 5955
rect 23715 5935 23729 5955
rect 23688 5933 23729 5935
rect 23757 5955 23799 5963
rect 23757 5935 23773 5955
rect 23792 5935 23799 5955
rect 23757 5933 23799 5935
rect 23688 5918 23799 5933
rect 23493 5796 23512 5835
rect 23557 5796 23565 5835
rect 23493 5779 23565 5796
rect 24027 5823 24064 6022
rect 24340 6018 24404 6030
rect 24027 5817 24068 5823
rect 24444 5819 24471 6170
rect 24594 6040 24673 6640
rect 24770 6188 24849 6773
rect 25053 6760 25090 6789
rect 25054 6758 25090 6760
rect 25266 6758 25303 6789
rect 25054 6736 25303 6758
rect 25135 6730 25246 6736
rect 25135 6722 25176 6730
rect 25135 6702 25143 6722
rect 25162 6702 25176 6722
rect 25135 6700 25176 6702
rect 25204 6722 25246 6730
rect 25204 6702 25220 6722
rect 25239 6702 25246 6722
rect 25204 6700 25246 6702
rect 25135 6685 25246 6700
rect 25474 6674 25511 6789
rect 25467 6562 25514 6674
rect 25635 6634 25665 6793
rect 25685 6792 25721 6793
rect 25787 6826 25824 6827
rect 25787 6825 25825 6826
rect 25787 6817 25851 6825
rect 25787 6797 25796 6817
rect 25816 6803 25851 6817
rect 25871 6803 25874 6823
rect 25816 6798 25874 6803
rect 25816 6797 25851 6798
rect 25787 6785 25851 6797
rect 25635 6630 25721 6634
rect 25635 6612 25650 6630
rect 25702 6612 25721 6630
rect 25635 6603 25721 6612
rect 25891 6564 25918 6937
rect 25750 6562 25918 6564
rect 25467 6536 25918 6562
rect 25467 6458 25514 6536
rect 25750 6535 25918 6536
rect 25412 6457 25514 6458
rect 25411 6449 25514 6457
rect 25411 6446 25463 6449
rect 25411 6411 25419 6446
rect 25444 6411 25463 6446
rect 25488 6411 25514 6449
rect 25411 6405 25514 6411
rect 25674 6450 25710 6454
rect 25674 6427 25682 6450
rect 25706 6427 25710 6450
rect 25674 6406 25710 6427
rect 25411 6401 25510 6405
rect 25674 6383 25682 6406
rect 25706 6383 25710 6406
rect 24303 5817 24471 5819
rect 24027 5791 24471 5817
rect 22223 5724 22288 5771
rect 22223 5706 22246 5724
rect 22264 5706 22288 5724
rect 23136 5751 23171 5753
rect 23136 5749 23240 5751
rect 24029 5749 24068 5791
rect 24303 5790 24471 5791
rect 23136 5742 24070 5749
rect 23136 5741 23187 5742
rect 23136 5721 23139 5741
rect 23164 5722 23187 5741
rect 23219 5722 24070 5742
rect 23164 5721 24070 5722
rect 23136 5714 24070 5721
rect 23409 5713 24070 5714
rect 22223 5685 22288 5706
rect 22500 5696 22540 5699
rect 22500 5692 23403 5696
rect 22500 5672 23377 5692
rect 23397 5672 23403 5692
rect 22500 5669 23403 5672
rect 22224 5625 22289 5645
rect 22224 5607 22248 5625
rect 22266 5607 22289 5625
rect 22224 5580 22289 5607
rect 22500 5580 22540 5669
rect 22984 5667 23400 5669
rect 22984 5666 23325 5667
rect 22641 5635 22751 5649
rect 22641 5632 22684 5635
rect 22641 5627 22645 5632
rect 22223 5545 22540 5580
rect 22563 5605 22645 5627
rect 22674 5605 22684 5632
rect 22712 5608 22719 5635
rect 22748 5627 22751 5635
rect 22748 5608 22813 5627
rect 22712 5605 22813 5608
rect 22563 5603 22813 5605
rect 20924 5512 20946 5530
rect 20964 5512 20989 5530
rect 20924 5493 20989 5512
rect 20617 5468 20654 5469
rect 20040 5447 20076 5468
rect 20466 5447 20497 5468
rect 20704 5463 20712 5472
rect 20701 5447 20712 5463
rect 19873 5443 19973 5447
rect 19873 5439 19935 5443
rect 19873 5413 19880 5439
rect 19906 5417 19935 5439
rect 19961 5417 19973 5443
rect 19906 5413 19973 5417
rect 19873 5410 19973 5413
rect 20041 5410 20076 5447
rect 20138 5444 20497 5447
rect 20138 5439 20360 5444
rect 20138 5415 20151 5439
rect 20175 5420 20360 5439
rect 20384 5420 20497 5444
rect 20175 5415 20497 5420
rect 20138 5411 20497 5415
rect 20564 5439 20712 5447
rect 20564 5419 20575 5439
rect 20595 5430 20712 5439
rect 20761 5463 20768 5472
rect 22224 5469 22289 5545
rect 22563 5524 22600 5603
rect 22641 5590 22751 5603
rect 22715 5534 22746 5535
rect 22563 5504 22572 5524
rect 22592 5504 22600 5524
rect 22563 5494 22600 5504
rect 22659 5524 22746 5534
rect 22659 5504 22668 5524
rect 22688 5504 22746 5524
rect 22659 5495 22746 5504
rect 22659 5494 22696 5495
rect 20761 5430 20769 5463
rect 22224 5451 22246 5469
rect 22264 5451 22289 5469
rect 20595 5419 20769 5430
rect 20564 5412 20769 5419
rect 20564 5411 20605 5412
rect 20040 5385 20076 5410
rect 19888 5358 19925 5359
rect 19984 5358 20021 5359
rect 20040 5358 20047 5385
rect 19564 5333 19572 5353
rect 19592 5333 19601 5353
rect 19418 5322 19449 5323
rect 19413 5254 19523 5267
rect 19564 5254 19601 5333
rect 19788 5349 19926 5358
rect 19788 5329 19897 5349
rect 19917 5329 19926 5349
rect 19788 5322 19926 5329
rect 19984 5355 20047 5358
rect 20068 5358 20076 5385
rect 20095 5358 20132 5359
rect 20068 5355 20132 5358
rect 19984 5349 20132 5355
rect 19984 5329 19993 5349
rect 20013 5329 20103 5349
rect 20123 5329 20132 5349
rect 19788 5320 19884 5322
rect 19984 5319 20132 5329
rect 20191 5349 20228 5359
rect 20303 5358 20340 5359
rect 20284 5356 20340 5358
rect 20191 5329 20199 5349
rect 20219 5329 20228 5349
rect 20040 5318 20076 5319
rect 19351 5252 19601 5254
rect 19351 5249 19452 5252
rect 19351 5230 19416 5249
rect 19413 5222 19416 5230
rect 19445 5222 19452 5249
rect 19480 5225 19490 5252
rect 19519 5230 19601 5252
rect 19519 5225 19523 5230
rect 19480 5222 19523 5225
rect 19413 5208 19523 5222
rect 18839 5190 19180 5191
rect 18764 5185 19180 5190
rect 19888 5187 19925 5188
rect 20191 5187 20228 5329
rect 20253 5349 20340 5356
rect 20253 5346 20311 5349
rect 20253 5326 20258 5346
rect 20279 5329 20311 5346
rect 20331 5329 20340 5349
rect 20279 5326 20340 5329
rect 20253 5319 20340 5326
rect 20399 5349 20436 5359
rect 20399 5329 20407 5349
rect 20427 5329 20436 5349
rect 20253 5318 20284 5319
rect 20399 5250 20436 5329
rect 20466 5358 20497 5411
rect 20701 5409 20769 5412
rect 20701 5367 20713 5409
rect 20762 5367 20769 5409
rect 20516 5358 20553 5359
rect 20466 5349 20553 5358
rect 20466 5329 20524 5349
rect 20544 5329 20553 5349
rect 20466 5319 20553 5329
rect 20612 5349 20649 5359
rect 20701 5354 20769 5367
rect 20924 5431 20989 5448
rect 20924 5413 20948 5431
rect 20966 5413 20989 5431
rect 22224 5430 22289 5451
rect 22437 5449 22502 5458
rect 20612 5329 20620 5349
rect 20640 5329 20649 5349
rect 20466 5318 20497 5319
rect 20461 5250 20571 5263
rect 20612 5250 20649 5329
rect 20924 5274 20989 5413
rect 22437 5412 22447 5449
rect 22487 5441 22502 5449
rect 22715 5442 22746 5495
rect 22776 5524 22813 5603
rect 22928 5534 22959 5535
rect 22776 5504 22785 5524
rect 22805 5504 22813 5524
rect 22776 5494 22813 5504
rect 22872 5527 22959 5534
rect 22872 5524 22933 5527
rect 22872 5504 22881 5524
rect 22901 5507 22933 5524
rect 22954 5507 22959 5527
rect 22901 5504 22959 5507
rect 22872 5497 22959 5504
rect 22984 5524 23021 5666
rect 23287 5665 23324 5666
rect 23136 5534 23172 5535
rect 22984 5504 22993 5524
rect 23013 5504 23021 5524
rect 22872 5495 22928 5497
rect 22872 5494 22909 5495
rect 22984 5494 23021 5504
rect 23080 5524 23228 5534
rect 23328 5531 23424 5533
rect 23080 5504 23089 5524
rect 23109 5504 23199 5524
rect 23219 5504 23228 5524
rect 23080 5498 23228 5504
rect 23080 5495 23144 5498
rect 23080 5494 23117 5495
rect 23136 5468 23144 5495
rect 23165 5495 23228 5498
rect 23286 5524 23424 5531
rect 23286 5504 23295 5524
rect 23315 5504 23424 5524
rect 23286 5495 23424 5504
rect 23165 5468 23172 5495
rect 23191 5494 23228 5495
rect 23287 5494 23324 5495
rect 23136 5443 23172 5468
rect 22607 5441 22648 5442
rect 22487 5434 22648 5441
rect 22487 5414 22617 5434
rect 22637 5414 22648 5434
rect 22487 5412 22648 5414
rect 22437 5406 22648 5412
rect 22715 5438 23074 5442
rect 22715 5433 23037 5438
rect 22715 5409 22828 5433
rect 22852 5414 23037 5433
rect 23061 5414 23074 5438
rect 22852 5409 23074 5414
rect 22715 5406 23074 5409
rect 23136 5406 23171 5443
rect 23239 5440 23339 5443
rect 23239 5436 23306 5440
rect 23239 5410 23251 5436
rect 23277 5414 23306 5436
rect 23332 5414 23339 5440
rect 23277 5410 23339 5414
rect 23239 5406 23339 5410
rect 22437 5393 22504 5406
rect 20924 5268 20946 5274
rect 20399 5248 20649 5250
rect 20399 5245 20500 5248
rect 20399 5226 20464 5245
rect 20461 5218 20464 5226
rect 20493 5218 20500 5245
rect 20528 5221 20538 5248
rect 20567 5226 20649 5248
rect 20678 5256 20946 5268
rect 20964 5256 20989 5274
rect 20678 5233 20989 5256
rect 22229 5370 22285 5390
rect 22229 5352 22248 5370
rect 22266 5352 22285 5370
rect 22229 5239 22285 5352
rect 22437 5372 22451 5393
rect 22487 5372 22504 5393
rect 22715 5385 22746 5406
rect 23136 5385 23172 5406
rect 22558 5384 22595 5385
rect 22437 5365 22504 5372
rect 22557 5375 22595 5384
rect 20678 5232 20733 5233
rect 20567 5221 20571 5226
rect 20528 5218 20571 5221
rect 20461 5204 20571 5218
rect 19887 5186 20228 5187
rect 18764 5165 18767 5185
rect 18787 5165 19180 5185
rect 19812 5185 20228 5186
rect 20678 5185 20721 5232
rect 19812 5181 20721 5185
rect 19131 5132 19176 5165
rect 19812 5161 19815 5181
rect 19835 5161 20721 5181
rect 20189 5156 20721 5161
rect 20929 5175 20988 5197
rect 20929 5157 20948 5175
rect 20966 5157 20988 5175
rect 19977 5132 20076 5134
rect 19131 5122 20076 5132
rect 19131 5096 19999 5122
rect 19132 5095 19999 5096
rect 19977 5084 19999 5095
rect 20024 5087 20043 5122
rect 20068 5087 20076 5122
rect 20024 5084 20076 5087
rect 19977 5076 20076 5084
rect 20003 5075 20075 5076
rect 20929 5027 20988 5157
rect 22229 5110 22284 5239
rect 22437 5213 22502 5365
rect 22557 5355 22566 5375
rect 22586 5355 22595 5375
rect 22557 5347 22595 5355
rect 22661 5379 22746 5385
rect 22771 5384 22808 5385
rect 22661 5359 22669 5379
rect 22689 5359 22746 5379
rect 22661 5351 22746 5359
rect 22770 5375 22808 5384
rect 22770 5355 22779 5375
rect 22799 5355 22808 5375
rect 22661 5350 22697 5351
rect 22770 5347 22808 5355
rect 22874 5379 22959 5385
rect 22979 5384 23016 5385
rect 22874 5359 22882 5379
rect 22902 5378 22959 5379
rect 22902 5359 22931 5378
rect 22874 5358 22931 5359
rect 22952 5358 22959 5378
rect 22874 5351 22959 5358
rect 22978 5375 23016 5384
rect 22978 5355 22987 5375
rect 23007 5355 23016 5375
rect 22874 5350 22910 5351
rect 22978 5347 23016 5355
rect 23082 5379 23226 5385
rect 23082 5359 23090 5379
rect 23110 5359 23198 5379
rect 23218 5359 23226 5379
rect 23082 5351 23226 5359
rect 23082 5350 23118 5351
rect 23190 5350 23226 5351
rect 23292 5384 23329 5385
rect 23292 5383 23330 5384
rect 23292 5375 23356 5383
rect 23292 5355 23301 5375
rect 23321 5361 23356 5375
rect 23376 5361 23379 5381
rect 23321 5356 23379 5361
rect 23321 5355 23356 5356
rect 22558 5318 22595 5347
rect 22559 5316 22595 5318
rect 22771 5316 22808 5347
rect 22559 5294 22808 5316
rect 22640 5288 22751 5294
rect 22640 5280 22681 5288
rect 22640 5260 22648 5280
rect 22667 5260 22681 5280
rect 22640 5258 22681 5260
rect 22709 5280 22751 5288
rect 22709 5260 22725 5280
rect 22744 5260 22751 5280
rect 22709 5258 22751 5260
rect 22640 5243 22751 5258
rect 22979 5248 23016 5347
rect 23292 5343 23356 5355
rect 22642 5234 22746 5243
rect 22430 5203 22551 5213
rect 22430 5201 22499 5203
rect 22430 5160 22443 5201
rect 22480 5162 22499 5201
rect 22536 5162 22551 5203
rect 22480 5160 22551 5162
rect 22430 5142 22551 5160
rect 22223 5098 22284 5110
rect 22977 5098 23018 5248
rect 23396 5240 23423 5495
rect 23485 5485 23565 5496
rect 23485 5459 23502 5485
rect 23542 5459 23565 5485
rect 23485 5432 23565 5459
rect 23485 5406 23506 5432
rect 23546 5406 23565 5432
rect 23485 5387 23565 5406
rect 23485 5361 23509 5387
rect 23549 5361 23565 5387
rect 23485 5310 23565 5361
rect 22223 5095 23018 5098
rect 23397 5109 23423 5240
rect 23487 5154 23557 5310
rect 23486 5138 23562 5154
rect 23397 5095 23425 5109
rect 22223 5060 23425 5095
rect 23486 5101 23501 5138
rect 23545 5101 23562 5138
rect 23486 5081 23562 5101
rect 24600 5131 24670 6040
rect 24769 5519 24850 6188
rect 25674 6083 25710 6383
rect 25598 6054 25711 6083
rect 25598 5689 25629 6054
rect 25522 5669 25915 5689
rect 25935 5669 25938 5689
rect 25522 5664 25938 5669
rect 25522 5663 25863 5664
rect 25179 5632 25289 5646
rect 25179 5629 25222 5632
rect 25179 5624 25183 5629
rect 25101 5602 25183 5624
rect 25212 5602 25222 5629
rect 25250 5605 25257 5632
rect 25286 5624 25289 5632
rect 25286 5605 25351 5624
rect 25250 5602 25351 5605
rect 25101 5600 25351 5602
rect 25101 5521 25138 5600
rect 25179 5587 25289 5600
rect 25253 5531 25284 5532
rect 24763 5439 24862 5519
rect 25101 5501 25110 5521
rect 25130 5501 25138 5521
rect 25101 5491 25138 5501
rect 25197 5521 25284 5531
rect 25197 5501 25206 5521
rect 25226 5501 25284 5521
rect 25197 5492 25284 5501
rect 25197 5491 25234 5492
rect 25253 5439 25284 5492
rect 25314 5521 25351 5600
rect 25466 5531 25497 5532
rect 25314 5501 25323 5521
rect 25343 5501 25351 5521
rect 25314 5491 25351 5501
rect 25410 5524 25497 5531
rect 25410 5521 25471 5524
rect 25410 5501 25419 5521
rect 25439 5504 25471 5521
rect 25492 5504 25497 5524
rect 25439 5501 25497 5504
rect 25410 5494 25497 5501
rect 25522 5521 25559 5663
rect 25825 5662 25862 5663
rect 25674 5531 25710 5532
rect 25522 5501 25531 5521
rect 25551 5501 25559 5521
rect 25410 5492 25466 5494
rect 25410 5491 25447 5492
rect 25522 5491 25559 5501
rect 25618 5521 25766 5531
rect 25866 5528 25962 5530
rect 25618 5501 25627 5521
rect 25647 5501 25737 5521
rect 25757 5501 25766 5521
rect 25618 5495 25766 5501
rect 25618 5492 25682 5495
rect 25618 5491 25655 5492
rect 25674 5465 25682 5492
rect 25703 5492 25766 5495
rect 25824 5521 25962 5528
rect 25824 5501 25833 5521
rect 25853 5501 25962 5521
rect 25824 5492 25962 5501
rect 25703 5465 25710 5492
rect 25729 5491 25766 5492
rect 25825 5491 25862 5492
rect 25674 5440 25710 5465
rect 24763 5438 25103 5439
rect 25145 5438 25186 5439
rect 24763 5431 25186 5438
rect 24763 5411 25155 5431
rect 25175 5411 25186 5431
rect 24763 5403 25186 5411
rect 25253 5435 25612 5439
rect 25253 5430 25575 5435
rect 25253 5406 25366 5430
rect 25390 5411 25575 5430
rect 25599 5411 25612 5435
rect 25390 5406 25612 5411
rect 25253 5403 25612 5406
rect 25674 5403 25709 5440
rect 25777 5437 25877 5440
rect 25777 5433 25844 5437
rect 25777 5407 25789 5433
rect 25815 5411 25844 5433
rect 25870 5411 25877 5437
rect 25815 5407 25877 5411
rect 25777 5403 25877 5407
rect 24763 5399 25103 5403
rect 24600 5081 24672 5131
rect 19651 4997 19727 5021
rect 19651 4931 19663 4997
rect 19717 4931 19727 4997
rect 20195 4952 20236 4954
rect 20467 4952 20571 4954
rect 20929 4952 20990 5027
rect 22223 4985 22284 5060
rect 22642 5058 22746 5060
rect 22977 5058 23018 5060
rect 23486 5015 23496 5081
rect 23550 5015 23562 5081
rect 23486 4991 23562 5015
rect 18541 4881 18613 4931
rect 18110 4609 18446 4613
rect 17336 4605 17436 4609
rect 17336 4601 17398 4605
rect 17336 4575 17343 4601
rect 17369 4579 17398 4601
rect 17424 4579 17436 4605
rect 17369 4575 17436 4579
rect 17336 4572 17436 4575
rect 17504 4572 17539 4609
rect 17601 4606 17960 4609
rect 17601 4601 17823 4606
rect 17601 4577 17614 4601
rect 17638 4582 17823 4601
rect 17847 4582 17960 4606
rect 17638 4577 17960 4582
rect 17601 4573 17960 4577
rect 18027 4601 18446 4609
rect 18027 4581 18038 4601
rect 18058 4581 18446 4601
rect 18027 4574 18446 4581
rect 18027 4573 18068 4574
rect 18110 4573 18446 4574
rect 17503 4547 17539 4572
rect 17351 4520 17388 4521
rect 17447 4520 17484 4521
rect 17503 4520 17510 4547
rect 17251 4511 17389 4520
rect 17251 4491 17360 4511
rect 17380 4491 17389 4511
rect 17251 4484 17389 4491
rect 17447 4517 17510 4520
rect 17531 4520 17539 4547
rect 17558 4520 17595 4521
rect 17531 4517 17595 4520
rect 17447 4511 17595 4517
rect 17447 4491 17456 4511
rect 17476 4491 17566 4511
rect 17586 4491 17595 4511
rect 17251 4482 17347 4484
rect 17447 4481 17595 4491
rect 17654 4511 17691 4521
rect 17766 4520 17803 4521
rect 17747 4518 17803 4520
rect 17654 4491 17662 4511
rect 17682 4491 17691 4511
rect 17503 4480 17539 4481
rect 17351 4349 17388 4350
rect 17654 4349 17691 4491
rect 17716 4511 17803 4518
rect 17716 4508 17774 4511
rect 17716 4488 17721 4508
rect 17742 4491 17774 4508
rect 17794 4491 17803 4511
rect 17742 4488 17803 4491
rect 17716 4481 17803 4488
rect 17862 4511 17899 4521
rect 17862 4491 17870 4511
rect 17890 4491 17899 4511
rect 17716 4480 17747 4481
rect 17862 4412 17899 4491
rect 17929 4520 17960 4573
rect 18354 4537 18446 4573
rect 17979 4520 18016 4521
rect 17929 4511 18016 4520
rect 17929 4491 17987 4511
rect 18007 4491 18016 4511
rect 17929 4481 18016 4491
rect 18075 4511 18112 4521
rect 18075 4491 18083 4511
rect 18103 4491 18112 4511
rect 17929 4480 17960 4481
rect 17924 4412 18034 4425
rect 18075 4412 18112 4491
rect 17862 4410 18112 4412
rect 17862 4407 17963 4410
rect 17862 4388 17927 4407
rect 17924 4380 17927 4388
rect 17956 4380 17963 4407
rect 17991 4383 18001 4410
rect 18030 4388 18112 4410
rect 18030 4383 18034 4388
rect 17991 4380 18034 4383
rect 17924 4366 18034 4380
rect 17350 4348 17691 4349
rect 17275 4343 17691 4348
rect 17275 4323 17278 4343
rect 17298 4323 17691 4343
rect 17435 4279 17540 4282
rect 17434 4256 17540 4279
rect 16554 4254 17055 4256
rect 17196 4254 17545 4256
rect 14668 4233 14705 4254
rect 14668 4196 14679 4233
rect 14696 4196 14705 4233
rect 16554 4248 17545 4254
rect 16554 4243 17506 4248
rect 16554 4222 17465 4243
rect 17485 4227 17506 4243
rect 17526 4227 17545 4248
rect 17485 4222 17545 4227
rect 16554 4197 17545 4222
rect 17030 4196 17212 4197
rect 14668 4186 14705 4196
rect 14514 4143 14908 4163
rect 14928 4143 14931 4163
rect 14515 4138 14931 4143
rect 14515 4137 14856 4138
rect 14172 4106 14282 4120
rect 14172 4103 14215 4106
rect 14172 4098 14176 4103
rect 14094 4076 14176 4098
rect 14205 4076 14215 4103
rect 14243 4079 14250 4106
rect 14279 4098 14282 4106
rect 14279 4079 14344 4098
rect 14243 4076 14344 4079
rect 14094 4074 14344 4076
rect 14094 3995 14131 4074
rect 14172 4061 14282 4074
rect 14246 4005 14277 4006
rect 14094 3975 14103 3995
rect 14123 3975 14131 3995
rect 14094 3965 14131 3975
rect 14190 3995 14277 4005
rect 14190 3975 14199 3995
rect 14219 3975 14277 3995
rect 14190 3966 14277 3975
rect 14190 3965 14227 3966
rect 14246 3913 14277 3966
rect 14307 3995 14344 4074
rect 14459 4005 14490 4006
rect 14307 3975 14316 3995
rect 14336 3975 14344 3995
rect 14307 3965 14344 3975
rect 14403 3998 14490 4005
rect 14403 3995 14464 3998
rect 14403 3975 14412 3995
rect 14432 3978 14464 3995
rect 14485 3978 14490 3998
rect 14432 3975 14490 3978
rect 14403 3968 14490 3975
rect 14515 3995 14552 4137
rect 14818 4136 14855 4137
rect 14667 4005 14703 4006
rect 14515 3975 14524 3995
rect 14544 3975 14552 3995
rect 14403 3966 14459 3968
rect 14403 3965 14440 3966
rect 14515 3965 14552 3975
rect 14611 3995 14759 4005
rect 14859 4002 14955 4004
rect 14611 3975 14620 3995
rect 14640 3975 14730 3995
rect 14750 3975 14759 3995
rect 14611 3969 14759 3975
rect 14611 3966 14675 3969
rect 14611 3965 14648 3966
rect 14667 3939 14675 3966
rect 14696 3966 14759 3969
rect 14817 3995 14955 4002
rect 14817 3975 14826 3995
rect 14846 3975 14955 3995
rect 14817 3966 14955 3975
rect 17584 3967 17615 4323
rect 14696 3939 14703 3966
rect 14722 3965 14759 3966
rect 14818 3965 14855 3966
rect 14667 3914 14703 3939
rect 14138 3912 14179 3913
rect 14058 3907 14179 3912
rect 14009 3905 14179 3907
rect 14009 3894 14148 3905
rect 14009 3871 14032 3894
rect 14058 3885 14148 3894
rect 14168 3885 14179 3905
rect 14058 3877 14179 3885
rect 14246 3909 14605 3913
rect 14246 3904 14568 3909
rect 14246 3880 14359 3904
rect 14383 3885 14568 3904
rect 14592 3885 14605 3909
rect 14383 3880 14605 3885
rect 14246 3877 14605 3880
rect 14667 3877 14702 3914
rect 14770 3911 14870 3914
rect 14770 3907 14837 3911
rect 14770 3881 14782 3907
rect 14808 3885 14837 3907
rect 14863 3885 14870 3911
rect 14808 3881 14870 3885
rect 14770 3877 14870 3881
rect 14058 3871 14066 3877
rect 14009 3863 14066 3871
rect 14246 3856 14277 3877
rect 14667 3856 14703 3877
rect 14089 3855 14126 3856
rect 14088 3846 14126 3855
rect 14088 3826 14097 3846
rect 14117 3826 14126 3846
rect 14088 3818 14126 3826
rect 14192 3850 14277 3856
rect 14302 3855 14339 3856
rect 14192 3830 14200 3850
rect 14220 3830 14277 3850
rect 14192 3822 14277 3830
rect 14301 3846 14339 3855
rect 14301 3826 14310 3846
rect 14330 3826 14339 3846
rect 14192 3821 14228 3822
rect 14301 3818 14339 3826
rect 14405 3850 14490 3856
rect 14510 3855 14547 3856
rect 14405 3830 14413 3850
rect 14433 3849 14490 3850
rect 14433 3830 14462 3849
rect 14405 3829 14462 3830
rect 14483 3829 14490 3849
rect 14405 3822 14490 3829
rect 14509 3846 14547 3855
rect 14509 3826 14518 3846
rect 14538 3826 14547 3846
rect 14405 3821 14441 3822
rect 14509 3818 14547 3826
rect 14613 3850 14757 3856
rect 14613 3830 14621 3850
rect 14641 3830 14729 3850
rect 14749 3830 14757 3850
rect 14613 3822 14757 3830
rect 14613 3821 14649 3822
rect 14721 3821 14757 3822
rect 14823 3855 14860 3856
rect 14823 3854 14861 3855
rect 14823 3846 14887 3854
rect 14823 3826 14832 3846
rect 14852 3832 14887 3846
rect 14907 3832 14910 3852
rect 14852 3827 14910 3832
rect 14852 3826 14887 3827
rect 14089 3789 14126 3818
rect 14090 3787 14126 3789
rect 14302 3787 14339 3818
rect 14090 3765 14339 3787
rect 14171 3759 14282 3765
rect 14171 3751 14212 3759
rect 14171 3731 14179 3751
rect 14198 3731 14212 3751
rect 14171 3729 14212 3731
rect 14240 3751 14282 3759
rect 14240 3731 14256 3751
rect 14275 3731 14282 3751
rect 14240 3729 14282 3731
rect 14171 3714 14282 3729
rect 14510 3703 14547 3818
rect 14823 3814 14887 3826
rect 14503 3697 14550 3703
rect 14927 3699 14954 3966
rect 17502 3938 17615 3967
rect 14786 3697 14954 3699
rect 14503 3671 14954 3697
rect 14503 3536 14550 3671
rect 14786 3670 14954 3671
rect 17503 3629 17539 3938
rect 18363 3824 18444 4537
rect 18543 3972 18613 4881
rect 19651 4911 19727 4931
rect 19651 4874 19668 4911
rect 19712 4874 19727 4911
rect 19788 4917 20990 4952
rect 19788 4903 19816 4917
rect 19651 4858 19727 4874
rect 19656 4702 19726 4858
rect 19790 4772 19816 4903
rect 20195 4914 20990 4917
rect 19648 4651 19728 4702
rect 19648 4625 19664 4651
rect 19704 4625 19728 4651
rect 19648 4606 19728 4625
rect 19648 4580 19667 4606
rect 19707 4580 19728 4606
rect 19648 4553 19728 4580
rect 19648 4527 19671 4553
rect 19711 4527 19728 4553
rect 19648 4516 19728 4527
rect 19790 4517 19817 4772
rect 20195 4764 20236 4914
rect 20929 4902 20990 4914
rect 20662 4852 20783 4870
rect 20662 4850 20733 4852
rect 20662 4809 20677 4850
rect 20714 4811 20733 4850
rect 20770 4811 20783 4852
rect 20714 4809 20783 4811
rect 20662 4799 20783 4809
rect 20467 4769 20571 4778
rect 19857 4657 19921 4669
rect 20197 4665 20234 4764
rect 20462 4754 20573 4769
rect 20462 4752 20504 4754
rect 20462 4732 20469 4752
rect 20488 4732 20504 4752
rect 20462 4724 20504 4732
rect 20532 4752 20573 4754
rect 20532 4732 20546 4752
rect 20565 4732 20573 4752
rect 20532 4724 20573 4732
rect 20462 4718 20573 4724
rect 20405 4696 20654 4718
rect 20405 4665 20442 4696
rect 20618 4694 20654 4696
rect 20618 4665 20655 4694
rect 19857 4656 19892 4657
rect 19834 4651 19892 4656
rect 19834 4631 19837 4651
rect 19857 4637 19892 4651
rect 19912 4637 19921 4657
rect 19857 4629 19921 4637
rect 19883 4628 19921 4629
rect 19884 4627 19921 4628
rect 19987 4661 20023 4662
rect 20095 4661 20131 4662
rect 19987 4653 20131 4661
rect 19987 4633 19995 4653
rect 20015 4633 20103 4653
rect 20123 4633 20131 4653
rect 19987 4627 20131 4633
rect 20197 4657 20235 4665
rect 20303 4661 20339 4662
rect 20197 4637 20206 4657
rect 20226 4637 20235 4657
rect 20197 4628 20235 4637
rect 20254 4654 20339 4661
rect 20254 4634 20261 4654
rect 20282 4653 20339 4654
rect 20282 4634 20311 4653
rect 20254 4633 20311 4634
rect 20331 4633 20339 4653
rect 20197 4627 20234 4628
rect 20254 4627 20339 4633
rect 20405 4657 20443 4665
rect 20516 4661 20552 4662
rect 20405 4637 20414 4657
rect 20434 4637 20443 4657
rect 20405 4628 20443 4637
rect 20467 4653 20552 4661
rect 20467 4633 20524 4653
rect 20544 4633 20552 4653
rect 20405 4627 20442 4628
rect 20467 4627 20552 4633
rect 20618 4657 20656 4665
rect 20618 4637 20627 4657
rect 20647 4637 20656 4657
rect 20711 4647 20776 4799
rect 20929 4773 20984 4902
rect 22225 4855 22284 4985
rect 23138 4936 23210 4937
rect 23137 4928 23236 4936
rect 23137 4925 23189 4928
rect 23137 4890 23145 4925
rect 23170 4890 23189 4925
rect 23214 4917 23236 4928
rect 23214 4916 24081 4917
rect 23214 4890 24082 4916
rect 23137 4880 24082 4890
rect 23137 4878 23236 4880
rect 22225 4837 22247 4855
rect 22265 4837 22284 4855
rect 22225 4815 22284 4837
rect 22492 4851 23024 4856
rect 22492 4831 23378 4851
rect 23398 4831 23401 4851
rect 24037 4847 24082 4880
rect 22492 4827 23401 4831
rect 22492 4780 22535 4827
rect 22985 4826 23401 4827
rect 24033 4827 24426 4847
rect 24446 4827 24449 4847
rect 22985 4825 23326 4826
rect 22642 4794 22752 4808
rect 22642 4791 22685 4794
rect 22642 4786 22646 4791
rect 22480 4779 22535 4780
rect 20618 4628 20656 4637
rect 20709 4640 20776 4647
rect 20618 4627 20655 4628
rect 20041 4606 20077 4627
rect 20467 4606 20498 4627
rect 20709 4619 20726 4640
rect 20762 4619 20776 4640
rect 20928 4660 20984 4773
rect 20928 4642 20947 4660
rect 20965 4642 20984 4660
rect 20928 4622 20984 4642
rect 22224 4756 22535 4779
rect 22224 4738 22249 4756
rect 22267 4744 22535 4756
rect 22564 4764 22646 4786
rect 22675 4764 22685 4791
rect 22713 4767 22720 4794
rect 22749 4786 22752 4794
rect 22749 4767 22814 4786
rect 22713 4764 22814 4767
rect 22564 4762 22814 4764
rect 22267 4738 22289 4744
rect 20709 4606 20776 4619
rect 19874 4602 19974 4606
rect 19874 4598 19936 4602
rect 19874 4572 19881 4598
rect 19907 4576 19936 4598
rect 19962 4576 19974 4602
rect 19907 4572 19974 4576
rect 19874 4569 19974 4572
rect 20042 4569 20077 4606
rect 20139 4603 20498 4606
rect 20139 4598 20361 4603
rect 20139 4574 20152 4598
rect 20176 4579 20361 4598
rect 20385 4579 20498 4603
rect 20176 4574 20498 4579
rect 20139 4570 20498 4574
rect 20565 4600 20776 4606
rect 20565 4598 20726 4600
rect 20565 4578 20576 4598
rect 20596 4578 20726 4598
rect 20565 4571 20726 4578
rect 20565 4570 20606 4571
rect 20041 4544 20077 4569
rect 19889 4517 19926 4518
rect 19985 4517 20022 4518
rect 20041 4517 20048 4544
rect 19789 4508 19927 4517
rect 19789 4488 19898 4508
rect 19918 4488 19927 4508
rect 19789 4481 19927 4488
rect 19985 4514 20048 4517
rect 20069 4517 20077 4544
rect 20096 4517 20133 4518
rect 20069 4514 20133 4517
rect 19985 4508 20133 4514
rect 19985 4488 19994 4508
rect 20014 4488 20104 4508
rect 20124 4488 20133 4508
rect 19789 4479 19885 4481
rect 19985 4478 20133 4488
rect 20192 4508 20229 4518
rect 20304 4517 20341 4518
rect 20285 4515 20341 4517
rect 20192 4488 20200 4508
rect 20220 4488 20229 4508
rect 20041 4477 20077 4478
rect 19889 4346 19926 4347
rect 20192 4346 20229 4488
rect 20254 4508 20341 4515
rect 20254 4505 20312 4508
rect 20254 4485 20259 4505
rect 20280 4488 20312 4505
rect 20332 4488 20341 4508
rect 20280 4485 20341 4488
rect 20254 4478 20341 4485
rect 20400 4508 20437 4518
rect 20400 4488 20408 4508
rect 20428 4488 20437 4508
rect 20254 4477 20285 4478
rect 20400 4409 20437 4488
rect 20467 4517 20498 4570
rect 20711 4563 20726 4571
rect 20766 4563 20776 4600
rect 22224 4599 22289 4738
rect 22564 4683 22601 4762
rect 22642 4749 22752 4762
rect 22716 4693 22747 4694
rect 22564 4663 22573 4683
rect 22593 4663 22601 4683
rect 20711 4554 20776 4563
rect 20924 4561 20989 4582
rect 22224 4581 22247 4599
rect 22265 4581 22289 4599
rect 22224 4564 22289 4581
rect 22444 4645 22512 4658
rect 22564 4653 22601 4663
rect 22660 4683 22747 4693
rect 22660 4663 22669 4683
rect 22689 4663 22747 4683
rect 22660 4654 22747 4663
rect 22660 4653 22697 4654
rect 22444 4603 22451 4645
rect 22500 4603 22512 4645
rect 22444 4600 22512 4603
rect 22716 4601 22747 4654
rect 22777 4683 22814 4762
rect 22929 4693 22960 4694
rect 22777 4663 22786 4683
rect 22806 4663 22814 4683
rect 22777 4653 22814 4663
rect 22873 4686 22960 4693
rect 22873 4683 22934 4686
rect 22873 4663 22882 4683
rect 22902 4666 22934 4683
rect 22955 4666 22960 4686
rect 22902 4663 22960 4666
rect 22873 4656 22960 4663
rect 22985 4683 23022 4825
rect 23288 4824 23325 4825
rect 24033 4822 24449 4827
rect 24033 4821 24374 4822
rect 23690 4790 23800 4804
rect 23690 4787 23733 4790
rect 23690 4782 23694 4787
rect 23612 4760 23694 4782
rect 23723 4760 23733 4787
rect 23761 4763 23768 4790
rect 23797 4782 23800 4790
rect 23797 4763 23862 4782
rect 23761 4760 23862 4763
rect 23612 4758 23862 4760
rect 23137 4693 23173 4694
rect 22985 4663 22994 4683
rect 23014 4663 23022 4683
rect 22873 4654 22929 4656
rect 22873 4653 22910 4654
rect 22985 4653 23022 4663
rect 23081 4683 23229 4693
rect 23329 4690 23425 4692
rect 23081 4663 23090 4683
rect 23110 4663 23200 4683
rect 23220 4663 23229 4683
rect 23081 4657 23229 4663
rect 23081 4654 23145 4657
rect 23081 4653 23118 4654
rect 23137 4627 23145 4654
rect 23166 4654 23229 4657
rect 23287 4683 23425 4690
rect 23287 4663 23296 4683
rect 23316 4663 23425 4683
rect 23287 4654 23425 4663
rect 23612 4679 23649 4758
rect 23690 4745 23800 4758
rect 23764 4689 23795 4690
rect 23612 4659 23621 4679
rect 23641 4659 23649 4679
rect 23166 4627 23173 4654
rect 23192 4653 23229 4654
rect 23288 4653 23325 4654
rect 23137 4602 23173 4627
rect 22608 4600 22649 4601
rect 22444 4593 22649 4600
rect 22444 4582 22618 4593
rect 20924 4543 20949 4561
rect 20967 4543 20989 4561
rect 22444 4549 22452 4582
rect 20517 4517 20554 4518
rect 20467 4508 20554 4517
rect 20467 4488 20525 4508
rect 20545 4488 20554 4508
rect 20467 4478 20554 4488
rect 20613 4508 20650 4518
rect 20613 4488 20621 4508
rect 20641 4488 20650 4508
rect 20467 4477 20498 4478
rect 20462 4409 20572 4422
rect 20613 4409 20650 4488
rect 20924 4467 20989 4543
rect 22445 4540 22452 4549
rect 22501 4573 22618 4582
rect 22638 4573 22649 4593
rect 22501 4565 22649 4573
rect 22716 4597 23075 4601
rect 22716 4592 23038 4597
rect 22716 4568 22829 4592
rect 22853 4573 23038 4592
rect 23062 4573 23075 4597
rect 22853 4568 23075 4573
rect 22716 4565 23075 4568
rect 23137 4565 23172 4602
rect 23240 4599 23340 4602
rect 23240 4595 23307 4599
rect 23240 4569 23252 4595
rect 23278 4573 23307 4595
rect 23333 4573 23340 4599
rect 23278 4569 23340 4573
rect 23240 4565 23340 4569
rect 22501 4549 22512 4565
rect 22501 4540 22509 4549
rect 22716 4544 22747 4565
rect 23137 4544 23173 4565
rect 22559 4543 22596 4544
rect 22224 4500 22289 4519
rect 22224 4482 22249 4500
rect 22267 4482 22289 4500
rect 20400 4407 20650 4409
rect 20400 4404 20501 4407
rect 20400 4385 20465 4404
rect 20462 4377 20465 4385
rect 20494 4377 20501 4404
rect 20529 4380 20539 4407
rect 20568 4385 20650 4407
rect 20673 4432 20990 4467
rect 20568 4380 20572 4385
rect 20529 4377 20572 4380
rect 20462 4363 20572 4377
rect 19888 4345 20229 4346
rect 19813 4343 20229 4345
rect 20673 4343 20713 4432
rect 20924 4405 20989 4432
rect 20924 4387 20947 4405
rect 20965 4387 20989 4405
rect 20924 4367 20989 4387
rect 19810 4340 20713 4343
rect 19810 4320 19816 4340
rect 19836 4320 20713 4340
rect 19810 4316 20713 4320
rect 20673 4313 20713 4316
rect 20925 4306 20990 4327
rect 19143 4298 19804 4299
rect 19143 4291 20077 4298
rect 19143 4290 20049 4291
rect 19143 4270 19994 4290
rect 20026 4271 20049 4290
rect 20074 4271 20077 4291
rect 20026 4270 20077 4271
rect 19143 4263 20077 4270
rect 18742 4221 18910 4222
rect 19145 4221 19184 4263
rect 19973 4261 20077 4263
rect 20042 4259 20077 4261
rect 20925 4288 20949 4306
rect 20967 4288 20990 4306
rect 20925 4241 20990 4288
rect 18742 4195 19186 4221
rect 18742 4193 18910 4195
rect 17503 3606 17507 3629
rect 17531 3606 17539 3629
rect 17703 3607 17802 3611
rect 17503 3585 17539 3606
rect 17503 3562 17507 3585
rect 17531 3562 17539 3585
rect 17503 3558 17539 3562
rect 17699 3601 17802 3607
rect 17699 3563 17725 3601
rect 17750 3566 17769 3601
rect 17794 3566 17802 3601
rect 17750 3563 17802 3566
rect 17699 3555 17802 3563
rect 17699 3554 17801 3555
rect 14501 3487 14560 3536
rect 14501 3459 14519 3487
rect 14547 3459 14560 3487
rect 14501 3449 14560 3459
rect 17295 3476 17463 3477
rect 17699 3476 17746 3554
rect 17295 3450 17746 3476
rect 17295 3448 17463 3450
rect 17295 3075 17322 3448
rect 17492 3400 17578 3409
rect 17492 3382 17511 3400
rect 17563 3382 17578 3400
rect 17492 3378 17578 3382
rect 17362 3215 17426 3227
rect 17362 3214 17397 3215
rect 17339 3209 17397 3214
rect 17339 3189 17342 3209
rect 17362 3195 17397 3209
rect 17417 3195 17426 3215
rect 17362 3187 17426 3195
rect 17388 3186 17426 3187
rect 17389 3185 17426 3186
rect 17492 3219 17528 3220
rect 17548 3219 17578 3378
rect 17699 3338 17746 3450
rect 17702 3223 17739 3338
rect 17967 3312 18078 3327
rect 17967 3310 18009 3312
rect 17967 3290 17974 3310
rect 17993 3290 18009 3310
rect 17967 3282 18009 3290
rect 18037 3310 18078 3312
rect 18037 3290 18051 3310
rect 18070 3290 18078 3310
rect 18037 3282 18078 3290
rect 17967 3276 18078 3282
rect 17910 3254 18159 3276
rect 17910 3223 17947 3254
rect 18123 3252 18159 3254
rect 18123 3223 18160 3252
rect 18364 3239 18443 3824
rect 18540 3372 18619 3972
rect 18742 3842 18769 4193
rect 19145 4189 19186 4195
rect 18809 3982 18873 3994
rect 19149 3990 19186 4189
rect 19648 4216 19720 4233
rect 19648 4177 19656 4216
rect 19701 4177 19720 4216
rect 19414 4079 19525 4094
rect 19414 4077 19456 4079
rect 19414 4057 19421 4077
rect 19440 4057 19456 4077
rect 19414 4049 19456 4057
rect 19484 4077 19525 4079
rect 19484 4057 19498 4077
rect 19517 4057 19525 4077
rect 19484 4049 19525 4057
rect 19414 4043 19525 4049
rect 19357 4021 19606 4043
rect 19357 3990 19394 4021
rect 19570 4019 19606 4021
rect 19570 3990 19607 4019
rect 18809 3981 18844 3982
rect 18786 3976 18844 3981
rect 18786 3956 18789 3976
rect 18809 3962 18844 3976
rect 18864 3962 18873 3982
rect 18809 3954 18873 3962
rect 18835 3953 18873 3954
rect 18836 3952 18873 3953
rect 18939 3986 18975 3987
rect 19047 3986 19083 3987
rect 18939 3978 19083 3986
rect 18939 3958 18947 3978
rect 18967 3958 19055 3978
rect 19075 3958 19083 3978
rect 18939 3952 19083 3958
rect 19149 3982 19187 3990
rect 19255 3986 19291 3987
rect 19149 3962 19158 3982
rect 19178 3962 19187 3982
rect 19149 3953 19187 3962
rect 19206 3979 19291 3986
rect 19206 3959 19213 3979
rect 19234 3978 19291 3979
rect 19234 3959 19263 3978
rect 19206 3958 19263 3959
rect 19283 3958 19291 3978
rect 19149 3952 19186 3953
rect 19206 3952 19291 3958
rect 19357 3982 19395 3990
rect 19468 3986 19504 3987
rect 19357 3962 19366 3982
rect 19386 3962 19395 3982
rect 19357 3953 19395 3962
rect 19419 3978 19504 3986
rect 19419 3958 19476 3978
rect 19496 3958 19504 3978
rect 19357 3952 19394 3953
rect 19419 3952 19504 3958
rect 19570 3982 19608 3990
rect 19570 3962 19579 3982
rect 19599 3962 19608 3982
rect 19570 3953 19608 3962
rect 19648 3967 19720 4177
rect 19790 4211 20990 4241
rect 19790 4210 20234 4211
rect 19790 4208 19958 4210
rect 19648 3953 19731 3967
rect 19570 3952 19607 3953
rect 18993 3931 19029 3952
rect 19419 3931 19450 3952
rect 19648 3931 19665 3953
rect 18826 3927 18926 3931
rect 18826 3923 18888 3927
rect 18826 3897 18833 3923
rect 18859 3901 18888 3923
rect 18914 3901 18926 3927
rect 18859 3897 18926 3901
rect 18826 3894 18926 3897
rect 18994 3894 19029 3931
rect 19091 3928 19450 3931
rect 19091 3923 19313 3928
rect 19091 3899 19104 3923
rect 19128 3904 19313 3923
rect 19337 3904 19450 3928
rect 19128 3899 19450 3904
rect 19091 3895 19450 3899
rect 19517 3923 19665 3931
rect 19517 3903 19528 3923
rect 19548 3920 19665 3923
rect 19718 3920 19731 3953
rect 19548 3903 19731 3920
rect 19517 3896 19731 3903
rect 19517 3895 19558 3896
rect 19648 3895 19731 3896
rect 18993 3869 19029 3894
rect 18841 3842 18878 3843
rect 18937 3842 18974 3843
rect 18993 3842 19000 3869
rect 18741 3833 18879 3842
rect 18741 3813 18850 3833
rect 18870 3813 18879 3833
rect 18741 3806 18879 3813
rect 18937 3839 19000 3842
rect 19021 3842 19029 3869
rect 19048 3842 19085 3843
rect 19021 3839 19085 3842
rect 18937 3833 19085 3839
rect 18937 3813 18946 3833
rect 18966 3813 19056 3833
rect 19076 3813 19085 3833
rect 18741 3804 18837 3806
rect 18937 3803 19085 3813
rect 19144 3833 19181 3843
rect 19256 3842 19293 3843
rect 19237 3840 19293 3842
rect 19144 3813 19152 3833
rect 19172 3813 19181 3833
rect 18993 3802 19029 3803
rect 18841 3671 18878 3672
rect 19144 3671 19181 3813
rect 19206 3833 19293 3840
rect 19206 3830 19264 3833
rect 19206 3810 19211 3830
rect 19232 3813 19264 3830
rect 19284 3813 19293 3833
rect 19232 3810 19293 3813
rect 19206 3803 19293 3810
rect 19352 3833 19389 3843
rect 19352 3813 19360 3833
rect 19380 3813 19389 3833
rect 19206 3802 19237 3803
rect 19352 3734 19389 3813
rect 19419 3842 19450 3895
rect 19656 3862 19670 3895
rect 19723 3862 19731 3895
rect 19656 3856 19731 3862
rect 19656 3851 19726 3856
rect 19469 3842 19506 3843
rect 19419 3833 19506 3842
rect 19419 3813 19477 3833
rect 19497 3813 19506 3833
rect 19419 3803 19506 3813
rect 19565 3833 19602 3843
rect 19790 3838 19817 4208
rect 19857 3978 19921 3990
rect 20197 3986 20234 4210
rect 20705 4191 20769 4193
rect 20701 4179 20769 4191
rect 20701 4146 20712 4179
rect 20752 4146 20769 4179
rect 20701 4136 20769 4146
rect 20462 4075 20573 4090
rect 20462 4073 20504 4075
rect 20462 4053 20469 4073
rect 20488 4053 20504 4073
rect 20462 4045 20504 4053
rect 20532 4073 20573 4075
rect 20532 4053 20546 4073
rect 20565 4053 20573 4073
rect 20532 4045 20573 4053
rect 20462 4039 20573 4045
rect 20405 4017 20654 4039
rect 20405 3986 20442 4017
rect 20618 4015 20654 4017
rect 20618 3986 20655 4015
rect 19857 3977 19892 3978
rect 19834 3972 19892 3977
rect 19834 3952 19837 3972
rect 19857 3958 19892 3972
rect 19912 3958 19921 3978
rect 19857 3950 19921 3958
rect 19883 3949 19921 3950
rect 19884 3948 19921 3949
rect 19987 3982 20023 3983
rect 20095 3982 20131 3983
rect 19987 3974 20131 3982
rect 19987 3954 19995 3974
rect 20015 3954 20103 3974
rect 20123 3954 20131 3974
rect 19987 3948 20131 3954
rect 20197 3978 20235 3986
rect 20303 3982 20339 3983
rect 20197 3958 20206 3978
rect 20226 3958 20235 3978
rect 20197 3949 20235 3958
rect 20254 3975 20339 3982
rect 20254 3955 20261 3975
rect 20282 3974 20339 3975
rect 20282 3955 20311 3974
rect 20254 3954 20311 3955
rect 20331 3954 20339 3974
rect 20197 3948 20234 3949
rect 20254 3948 20339 3954
rect 20405 3978 20443 3986
rect 20516 3982 20552 3983
rect 20405 3958 20414 3978
rect 20434 3958 20443 3978
rect 20405 3949 20443 3958
rect 20467 3974 20552 3982
rect 20467 3954 20524 3974
rect 20544 3954 20552 3974
rect 20405 3948 20442 3949
rect 20467 3948 20552 3954
rect 20618 3978 20656 3986
rect 20618 3958 20627 3978
rect 20647 3958 20656 3978
rect 20618 3949 20656 3958
rect 20705 3952 20769 4136
rect 20925 4010 20990 4211
rect 22224 4281 22289 4482
rect 22445 4356 22509 4540
rect 22558 4534 22596 4543
rect 22558 4514 22567 4534
rect 22587 4514 22596 4534
rect 22558 4506 22596 4514
rect 22662 4538 22747 4544
rect 22772 4543 22809 4544
rect 22662 4518 22670 4538
rect 22690 4518 22747 4538
rect 22662 4510 22747 4518
rect 22771 4534 22809 4543
rect 22771 4514 22780 4534
rect 22800 4514 22809 4534
rect 22662 4509 22698 4510
rect 22771 4506 22809 4514
rect 22875 4538 22960 4544
rect 22980 4543 23017 4544
rect 22875 4518 22883 4538
rect 22903 4537 22960 4538
rect 22903 4518 22932 4537
rect 22875 4517 22932 4518
rect 22953 4517 22960 4537
rect 22875 4510 22960 4517
rect 22979 4534 23017 4543
rect 22979 4514 22988 4534
rect 23008 4514 23017 4534
rect 22875 4509 22911 4510
rect 22979 4506 23017 4514
rect 23083 4538 23227 4544
rect 23083 4518 23091 4538
rect 23111 4518 23199 4538
rect 23219 4518 23227 4538
rect 23083 4510 23227 4518
rect 23083 4509 23119 4510
rect 23191 4509 23227 4510
rect 23293 4543 23330 4544
rect 23293 4542 23331 4543
rect 23293 4534 23357 4542
rect 23293 4514 23302 4534
rect 23322 4520 23357 4534
rect 23377 4520 23380 4540
rect 23322 4515 23380 4520
rect 23322 4514 23357 4515
rect 22559 4477 22596 4506
rect 22560 4475 22596 4477
rect 22772 4475 22809 4506
rect 22560 4453 22809 4475
rect 22641 4447 22752 4453
rect 22641 4439 22682 4447
rect 22641 4419 22649 4439
rect 22668 4419 22682 4439
rect 22641 4417 22682 4419
rect 22710 4439 22752 4447
rect 22710 4419 22726 4439
rect 22745 4419 22752 4439
rect 22710 4417 22752 4419
rect 22641 4402 22752 4417
rect 22445 4346 22513 4356
rect 22445 4313 22462 4346
rect 22502 4313 22513 4346
rect 22445 4301 22513 4313
rect 22445 4299 22509 4301
rect 22980 4282 23017 4506
rect 23293 4502 23357 4514
rect 23397 4284 23424 4654
rect 23612 4649 23649 4659
rect 23708 4679 23795 4689
rect 23708 4659 23717 4679
rect 23737 4659 23795 4679
rect 23708 4650 23795 4659
rect 23708 4649 23745 4650
rect 23488 4636 23558 4641
rect 23483 4630 23558 4636
rect 23483 4597 23491 4630
rect 23544 4597 23558 4630
rect 23764 4597 23795 4650
rect 23825 4679 23862 4758
rect 23977 4689 24008 4690
rect 23825 4659 23834 4679
rect 23854 4659 23862 4679
rect 23825 4649 23862 4659
rect 23921 4682 24008 4689
rect 23921 4679 23982 4682
rect 23921 4659 23930 4679
rect 23950 4662 23982 4679
rect 24003 4662 24008 4682
rect 23950 4659 24008 4662
rect 23921 4652 24008 4659
rect 24033 4679 24070 4821
rect 24336 4820 24373 4821
rect 24185 4689 24221 4690
rect 24033 4659 24042 4679
rect 24062 4659 24070 4679
rect 23921 4650 23977 4652
rect 23921 4649 23958 4650
rect 24033 4649 24070 4659
rect 24129 4679 24277 4689
rect 24377 4686 24473 4688
rect 24129 4659 24138 4679
rect 24158 4659 24248 4679
rect 24268 4659 24277 4679
rect 24129 4653 24277 4659
rect 24129 4650 24193 4653
rect 24129 4649 24166 4650
rect 24185 4623 24193 4650
rect 24214 4650 24277 4653
rect 24335 4679 24473 4686
rect 24335 4659 24344 4679
rect 24364 4659 24473 4679
rect 24335 4650 24473 4659
rect 24214 4623 24221 4650
rect 24240 4649 24277 4650
rect 24336 4649 24373 4650
rect 24185 4598 24221 4623
rect 23483 4596 23566 4597
rect 23656 4596 23697 4597
rect 23483 4589 23697 4596
rect 23483 4572 23666 4589
rect 23483 4539 23496 4572
rect 23549 4569 23666 4572
rect 23686 4569 23697 4589
rect 23549 4561 23697 4569
rect 23764 4593 24123 4597
rect 23764 4588 24086 4593
rect 23764 4564 23877 4588
rect 23901 4569 24086 4588
rect 24110 4569 24123 4593
rect 23901 4564 24123 4569
rect 23764 4561 24123 4564
rect 24185 4561 24220 4598
rect 24288 4595 24388 4598
rect 24288 4591 24355 4595
rect 24288 4565 24300 4591
rect 24326 4569 24355 4591
rect 24381 4569 24388 4595
rect 24326 4565 24388 4569
rect 24288 4561 24388 4565
rect 23549 4539 23566 4561
rect 23764 4540 23795 4561
rect 24185 4540 24221 4561
rect 23607 4539 23644 4540
rect 23483 4525 23566 4539
rect 23256 4282 23424 4284
rect 22980 4281 23424 4282
rect 22224 4251 23424 4281
rect 23494 4315 23566 4525
rect 23606 4530 23644 4539
rect 23606 4510 23615 4530
rect 23635 4510 23644 4530
rect 23606 4502 23644 4510
rect 23710 4534 23795 4540
rect 23820 4539 23857 4540
rect 23710 4514 23718 4534
rect 23738 4514 23795 4534
rect 23710 4506 23795 4514
rect 23819 4530 23857 4539
rect 23819 4510 23828 4530
rect 23848 4510 23857 4530
rect 23710 4505 23746 4506
rect 23819 4502 23857 4510
rect 23923 4534 24008 4540
rect 24028 4539 24065 4540
rect 23923 4514 23931 4534
rect 23951 4533 24008 4534
rect 23951 4514 23980 4533
rect 23923 4513 23980 4514
rect 24001 4513 24008 4533
rect 23923 4506 24008 4513
rect 24027 4530 24065 4539
rect 24027 4510 24036 4530
rect 24056 4510 24065 4530
rect 23923 4505 23959 4506
rect 24027 4502 24065 4510
rect 24131 4534 24275 4540
rect 24131 4514 24139 4534
rect 24159 4514 24247 4534
rect 24267 4514 24275 4534
rect 24131 4506 24275 4514
rect 24131 4505 24167 4506
rect 24239 4505 24275 4506
rect 24341 4539 24378 4540
rect 24341 4538 24379 4539
rect 24341 4530 24405 4538
rect 24341 4510 24350 4530
rect 24370 4516 24405 4530
rect 24425 4516 24428 4536
rect 24370 4511 24428 4516
rect 24370 4510 24405 4511
rect 23607 4473 23644 4502
rect 23608 4471 23644 4473
rect 23820 4471 23857 4502
rect 23608 4449 23857 4471
rect 23689 4443 23800 4449
rect 23689 4435 23730 4443
rect 23689 4415 23697 4435
rect 23716 4415 23730 4435
rect 23689 4413 23730 4415
rect 23758 4435 23800 4443
rect 23758 4415 23774 4435
rect 23793 4415 23800 4435
rect 23758 4413 23800 4415
rect 23689 4398 23800 4413
rect 23494 4276 23513 4315
rect 23558 4276 23566 4315
rect 23494 4259 23566 4276
rect 24028 4303 24065 4502
rect 24341 4498 24405 4510
rect 24028 4297 24069 4303
rect 24445 4299 24472 4650
rect 24601 4602 24672 5081
rect 24601 4518 24670 4602
rect 24304 4297 24472 4299
rect 24028 4271 24472 4297
rect 22224 4204 22289 4251
rect 22224 4186 22247 4204
rect 22265 4186 22289 4204
rect 23137 4231 23172 4233
rect 23137 4229 23241 4231
rect 24030 4229 24069 4271
rect 24304 4270 24472 4271
rect 23137 4222 24071 4229
rect 23137 4221 23188 4222
rect 23137 4201 23140 4221
rect 23165 4202 23188 4221
rect 23220 4202 24071 4222
rect 23165 4201 24071 4202
rect 23137 4194 24071 4201
rect 23410 4193 24071 4194
rect 22224 4165 22289 4186
rect 22501 4176 22541 4179
rect 22501 4172 23404 4176
rect 22501 4152 23378 4172
rect 23398 4152 23404 4172
rect 22501 4149 23404 4152
rect 22225 4105 22290 4125
rect 22225 4087 22249 4105
rect 22267 4087 22290 4105
rect 22225 4060 22290 4087
rect 22501 4060 22541 4149
rect 22985 4147 23401 4149
rect 22985 4146 23326 4147
rect 22642 4115 22752 4129
rect 22642 4112 22685 4115
rect 22642 4107 22646 4112
rect 22224 4025 22541 4060
rect 22564 4085 22646 4107
rect 22675 4085 22685 4112
rect 22713 4088 22720 4115
rect 22749 4107 22752 4115
rect 22749 4088 22814 4107
rect 22713 4085 22814 4088
rect 22564 4083 22814 4085
rect 20925 3992 20947 4010
rect 20965 3992 20990 4010
rect 20925 3973 20990 3992
rect 20618 3948 20655 3949
rect 20041 3927 20077 3948
rect 20467 3927 20498 3948
rect 20705 3943 20713 3952
rect 20702 3927 20713 3943
rect 19874 3923 19974 3927
rect 19874 3919 19936 3923
rect 19874 3893 19881 3919
rect 19907 3897 19936 3919
rect 19962 3897 19974 3923
rect 19907 3893 19974 3897
rect 19874 3890 19974 3893
rect 20042 3890 20077 3927
rect 20139 3924 20498 3927
rect 20139 3919 20361 3924
rect 20139 3895 20152 3919
rect 20176 3900 20361 3919
rect 20385 3900 20498 3924
rect 20176 3895 20498 3900
rect 20139 3891 20498 3895
rect 20565 3919 20713 3927
rect 20565 3899 20576 3919
rect 20596 3910 20713 3919
rect 20762 3943 20769 3952
rect 22225 3949 22290 4025
rect 22564 4004 22601 4083
rect 22642 4070 22752 4083
rect 22716 4014 22747 4015
rect 22564 3984 22573 4004
rect 22593 3984 22601 4004
rect 22564 3974 22601 3984
rect 22660 4004 22747 4014
rect 22660 3984 22669 4004
rect 22689 3984 22747 4004
rect 22660 3975 22747 3984
rect 22660 3974 22697 3975
rect 20762 3910 20770 3943
rect 22225 3931 22247 3949
rect 22265 3931 22290 3949
rect 20596 3899 20770 3910
rect 20565 3892 20770 3899
rect 20565 3891 20606 3892
rect 20041 3865 20077 3890
rect 19889 3838 19926 3839
rect 19985 3838 20022 3839
rect 20041 3838 20048 3865
rect 19565 3813 19573 3833
rect 19593 3813 19602 3833
rect 19419 3802 19450 3803
rect 19414 3734 19524 3747
rect 19565 3734 19602 3813
rect 19789 3829 19927 3838
rect 19789 3809 19898 3829
rect 19918 3809 19927 3829
rect 19789 3802 19927 3809
rect 19985 3835 20048 3838
rect 20069 3838 20077 3865
rect 20096 3838 20133 3839
rect 20069 3835 20133 3838
rect 19985 3829 20133 3835
rect 19985 3809 19994 3829
rect 20014 3809 20104 3829
rect 20124 3809 20133 3829
rect 19789 3800 19885 3802
rect 19985 3799 20133 3809
rect 20192 3829 20229 3839
rect 20304 3838 20341 3839
rect 20285 3836 20341 3838
rect 20192 3809 20200 3829
rect 20220 3809 20229 3829
rect 20041 3798 20077 3799
rect 19352 3732 19602 3734
rect 19352 3729 19453 3732
rect 19352 3710 19417 3729
rect 19414 3702 19417 3710
rect 19446 3702 19453 3729
rect 19481 3705 19491 3732
rect 19520 3710 19602 3732
rect 19520 3705 19524 3710
rect 19481 3702 19524 3705
rect 19414 3688 19524 3702
rect 18840 3670 19181 3671
rect 18765 3665 19181 3670
rect 19889 3667 19926 3668
rect 20192 3667 20229 3809
rect 20254 3829 20341 3836
rect 20254 3826 20312 3829
rect 20254 3806 20259 3826
rect 20280 3809 20312 3826
rect 20332 3809 20341 3829
rect 20280 3806 20341 3809
rect 20254 3799 20341 3806
rect 20400 3829 20437 3839
rect 20400 3809 20408 3829
rect 20428 3809 20437 3829
rect 20254 3798 20285 3799
rect 20400 3730 20437 3809
rect 20467 3838 20498 3891
rect 20702 3889 20770 3892
rect 20702 3847 20714 3889
rect 20763 3847 20770 3889
rect 20517 3838 20554 3839
rect 20467 3829 20554 3838
rect 20467 3809 20525 3829
rect 20545 3809 20554 3829
rect 20467 3799 20554 3809
rect 20613 3829 20650 3839
rect 20702 3834 20770 3847
rect 20925 3911 20990 3928
rect 20925 3893 20949 3911
rect 20967 3893 20990 3911
rect 22225 3910 22290 3931
rect 22438 3929 22503 3938
rect 20613 3809 20621 3829
rect 20641 3809 20650 3829
rect 20467 3798 20498 3799
rect 20462 3730 20572 3743
rect 20613 3730 20650 3809
rect 20925 3754 20990 3893
rect 22438 3892 22448 3929
rect 22488 3921 22503 3929
rect 22716 3922 22747 3975
rect 22777 4004 22814 4083
rect 22929 4014 22960 4015
rect 22777 3984 22786 4004
rect 22806 3984 22814 4004
rect 22777 3974 22814 3984
rect 22873 4007 22960 4014
rect 22873 4004 22934 4007
rect 22873 3984 22882 4004
rect 22902 3987 22934 4004
rect 22955 3987 22960 4007
rect 22902 3984 22960 3987
rect 22873 3977 22960 3984
rect 22985 4004 23022 4146
rect 23288 4145 23325 4146
rect 23137 4014 23173 4015
rect 22985 3984 22994 4004
rect 23014 3984 23022 4004
rect 22873 3975 22929 3977
rect 22873 3974 22910 3975
rect 22985 3974 23022 3984
rect 23081 4004 23229 4014
rect 23329 4011 23425 4013
rect 23081 3984 23090 4004
rect 23110 3984 23200 4004
rect 23220 3984 23229 4004
rect 23081 3978 23229 3984
rect 23081 3975 23145 3978
rect 23081 3974 23118 3975
rect 23137 3948 23145 3975
rect 23166 3975 23229 3978
rect 23287 4004 23425 4011
rect 24605 4006 24667 4518
rect 23287 3984 23296 4004
rect 23316 3984 23425 4004
rect 23287 3975 23425 3984
rect 23166 3948 23173 3975
rect 23192 3974 23229 3975
rect 23288 3974 23325 3975
rect 23137 3923 23173 3948
rect 22608 3921 22649 3922
rect 22488 3914 22649 3921
rect 22488 3894 22618 3914
rect 22638 3894 22649 3914
rect 22488 3892 22649 3894
rect 22438 3886 22649 3892
rect 22716 3918 23075 3922
rect 22716 3913 23038 3918
rect 22716 3889 22829 3913
rect 22853 3894 23038 3913
rect 23062 3894 23075 3918
rect 22853 3889 23075 3894
rect 22716 3886 23075 3889
rect 23137 3886 23172 3923
rect 23240 3920 23340 3923
rect 23240 3916 23307 3920
rect 23240 3890 23252 3916
rect 23278 3894 23307 3916
rect 23333 3894 23340 3920
rect 23278 3890 23340 3894
rect 23240 3886 23340 3890
rect 22438 3873 22505 3886
rect 20925 3748 20947 3754
rect 20400 3728 20650 3730
rect 20400 3725 20501 3728
rect 20400 3706 20465 3725
rect 20462 3698 20465 3706
rect 20494 3698 20501 3725
rect 20529 3701 20539 3728
rect 20568 3706 20650 3728
rect 20679 3736 20947 3748
rect 20965 3736 20990 3754
rect 20679 3713 20990 3736
rect 22230 3850 22286 3870
rect 22230 3832 22249 3850
rect 22267 3832 22286 3850
rect 22230 3719 22286 3832
rect 22438 3852 22452 3873
rect 22488 3852 22505 3873
rect 22716 3865 22747 3886
rect 23137 3865 23173 3886
rect 22559 3864 22596 3865
rect 22438 3845 22505 3852
rect 22558 3855 22596 3864
rect 20679 3712 20734 3713
rect 20568 3701 20572 3706
rect 20529 3698 20572 3701
rect 20462 3684 20572 3698
rect 19888 3666 20229 3667
rect 18765 3645 18768 3665
rect 18788 3645 19181 3665
rect 19813 3665 20229 3666
rect 20679 3665 20722 3712
rect 19813 3661 20722 3665
rect 19132 3612 19177 3645
rect 19813 3641 19816 3661
rect 19836 3641 20722 3661
rect 20190 3636 20722 3641
rect 20930 3655 20989 3677
rect 20930 3637 20949 3655
rect 20967 3637 20989 3655
rect 19978 3612 20077 3614
rect 19132 3602 20077 3612
rect 19132 3576 20000 3602
rect 19133 3575 20000 3576
rect 19978 3564 20000 3575
rect 20025 3567 20044 3602
rect 20069 3567 20077 3602
rect 20025 3564 20077 3567
rect 20930 3566 20989 3637
rect 22230 3581 22285 3719
rect 22438 3693 22503 3845
rect 22558 3835 22567 3855
rect 22587 3835 22596 3855
rect 22558 3827 22596 3835
rect 22662 3859 22747 3865
rect 22772 3864 22809 3865
rect 22662 3839 22670 3859
rect 22690 3839 22747 3859
rect 22662 3831 22747 3839
rect 22771 3855 22809 3864
rect 22771 3835 22780 3855
rect 22800 3835 22809 3855
rect 22662 3830 22698 3831
rect 22771 3827 22809 3835
rect 22875 3859 22960 3865
rect 22980 3864 23017 3865
rect 22875 3839 22883 3859
rect 22903 3858 22960 3859
rect 22903 3839 22932 3858
rect 22875 3838 22932 3839
rect 22953 3838 22960 3858
rect 22875 3831 22960 3838
rect 22979 3855 23017 3864
rect 22979 3835 22988 3855
rect 23008 3835 23017 3855
rect 22875 3830 22911 3831
rect 22979 3827 23017 3835
rect 23083 3859 23227 3865
rect 23083 3839 23091 3859
rect 23111 3839 23199 3859
rect 23219 3839 23227 3859
rect 23083 3831 23227 3839
rect 23083 3830 23119 3831
rect 23191 3830 23227 3831
rect 23293 3864 23330 3865
rect 23293 3863 23331 3864
rect 23293 3855 23357 3863
rect 23293 3835 23302 3855
rect 23322 3841 23357 3855
rect 23377 3841 23380 3861
rect 23322 3836 23380 3841
rect 23322 3835 23357 3836
rect 22559 3798 22596 3827
rect 22560 3796 22596 3798
rect 22772 3796 22809 3827
rect 22560 3774 22809 3796
rect 22641 3768 22752 3774
rect 22641 3760 22682 3768
rect 22641 3740 22649 3760
rect 22668 3740 22682 3760
rect 22641 3738 22682 3740
rect 22710 3760 22752 3768
rect 22710 3740 22726 3760
rect 22745 3740 22752 3760
rect 22710 3738 22752 3740
rect 22641 3725 22752 3738
rect 22980 3728 23017 3827
rect 23293 3823 23357 3835
rect 22431 3683 22552 3693
rect 22431 3681 22500 3683
rect 22431 3640 22444 3681
rect 22481 3642 22500 3681
rect 22537 3642 22552 3683
rect 22481 3640 22552 3642
rect 22431 3622 22552 3640
rect 22223 3578 22287 3581
rect 22643 3578 22747 3584
rect 22978 3578 23019 3728
rect 23397 3720 23424 3975
rect 23486 3965 23566 3976
rect 23486 3939 23503 3965
rect 23543 3939 23566 3965
rect 23486 3912 23566 3939
rect 24609 3967 24667 4006
rect 24609 3932 24671 3967
rect 23486 3886 23507 3912
rect 23547 3886 23566 3912
rect 23486 3867 23566 3886
rect 23486 3841 23510 3867
rect 23550 3841 23566 3867
rect 23486 3790 23566 3841
rect 24558 3905 24671 3932
rect 24558 3903 24617 3905
rect 24558 3872 24572 3903
rect 24597 3882 24617 3903
rect 24643 3882 24671 3905
rect 24597 3872 24671 3882
rect 24558 3862 24671 3872
rect 22223 3575 23019 3578
rect 23398 3589 23424 3720
rect 23398 3575 23426 3589
rect 19978 3556 20077 3564
rect 20004 3555 20076 3556
rect 19658 3529 19725 3548
rect 19658 3508 19675 3529
rect 18539 3330 18619 3372
rect 19656 3463 19675 3508
rect 19705 3508 19725 3529
rect 19705 3463 19726 3508
rect 20195 3505 20236 3507
rect 20467 3505 20571 3507
rect 20927 3505 20991 3566
rect 17600 3219 17636 3220
rect 17492 3211 17636 3219
rect 17492 3191 17500 3211
rect 17520 3191 17608 3211
rect 17628 3191 17636 3211
rect 17492 3185 17636 3191
rect 17702 3215 17740 3223
rect 17808 3219 17844 3220
rect 17702 3195 17711 3215
rect 17731 3195 17740 3215
rect 17702 3186 17740 3195
rect 17759 3212 17844 3219
rect 17759 3192 17766 3212
rect 17787 3211 17844 3212
rect 17787 3192 17816 3211
rect 17759 3191 17816 3192
rect 17836 3191 17844 3211
rect 17702 3185 17739 3186
rect 17759 3185 17844 3191
rect 17910 3215 17948 3223
rect 18021 3219 18057 3220
rect 17910 3195 17919 3215
rect 17939 3195 17948 3215
rect 17910 3186 17948 3195
rect 17972 3211 18057 3219
rect 17972 3191 18029 3211
rect 18049 3191 18057 3211
rect 17910 3185 17947 3186
rect 17972 3185 18057 3191
rect 18123 3215 18161 3223
rect 18123 3195 18132 3215
rect 18152 3195 18161 3215
rect 18123 3186 18161 3195
rect 18361 3203 18447 3239
rect 18123 3185 18160 3186
rect 17546 3164 17582 3185
rect 17972 3164 18003 3185
rect 18199 3164 18245 3168
rect 17379 3160 17479 3164
rect 17379 3156 17441 3160
rect 17379 3130 17386 3156
rect 17412 3134 17441 3156
rect 17467 3134 17479 3160
rect 17412 3130 17479 3134
rect 17379 3127 17479 3130
rect 17547 3127 17582 3164
rect 17644 3161 18003 3164
rect 17644 3156 17866 3161
rect 17644 3132 17657 3156
rect 17681 3137 17866 3156
rect 17890 3137 18003 3161
rect 17681 3132 18003 3137
rect 17644 3128 18003 3132
rect 18070 3156 18245 3164
rect 18070 3136 18081 3156
rect 18101 3136 18245 3156
rect 18361 3162 18378 3203
rect 18432 3162 18447 3203
rect 18361 3143 18447 3162
rect 18070 3129 18245 3136
rect 18070 3128 18111 3129
rect 17546 3102 17582 3127
rect 17394 3075 17431 3076
rect 17490 3075 17527 3076
rect 17546 3075 17553 3102
rect 17294 3066 17432 3075
rect 17294 3046 17403 3066
rect 17423 3046 17432 3066
rect 17294 3039 17432 3046
rect 17490 3072 17553 3075
rect 17574 3075 17582 3102
rect 17601 3075 17638 3076
rect 17574 3072 17638 3075
rect 17490 3066 17638 3072
rect 17490 3046 17499 3066
rect 17519 3046 17609 3066
rect 17629 3046 17638 3066
rect 17294 3037 17390 3039
rect 17490 3036 17638 3046
rect 17697 3066 17734 3076
rect 17809 3075 17846 3076
rect 17790 3073 17846 3075
rect 17697 3046 17705 3066
rect 17725 3046 17734 3066
rect 17546 3035 17582 3036
rect 17394 2904 17431 2905
rect 17697 2904 17734 3046
rect 17759 3066 17846 3073
rect 17759 3063 17817 3066
rect 17759 3043 17764 3063
rect 17785 3046 17817 3063
rect 17837 3046 17846 3066
rect 17785 3043 17846 3046
rect 17759 3036 17846 3043
rect 17905 3066 17942 3076
rect 17905 3046 17913 3066
rect 17933 3046 17942 3066
rect 17759 3035 17790 3036
rect 17905 2967 17942 3046
rect 17972 3075 18003 3128
rect 18022 3075 18059 3076
rect 17972 3066 18059 3075
rect 17972 3046 18030 3066
rect 18050 3046 18059 3066
rect 17972 3036 18059 3046
rect 18118 3066 18155 3076
rect 18118 3046 18126 3066
rect 18146 3046 18155 3066
rect 17972 3035 18003 3036
rect 17967 2967 18077 2980
rect 18118 2967 18155 3046
rect 18199 3046 18245 3129
rect 18539 3046 18614 3330
rect 19656 3255 19726 3463
rect 19788 3470 20991 3505
rect 22223 3540 23426 3575
rect 23488 3582 23558 3790
rect 22223 3479 22287 3540
rect 22643 3538 22747 3540
rect 22978 3538 23019 3540
rect 23488 3537 23509 3582
rect 23489 3516 23509 3537
rect 23539 3537 23558 3582
rect 23539 3516 23556 3537
rect 23489 3497 23556 3516
rect 23138 3489 23210 3490
rect 23137 3481 23236 3489
rect 19788 3456 19816 3470
rect 19790 3325 19816 3456
rect 20195 3467 20991 3470
rect 19648 3204 19728 3255
rect 19648 3178 19664 3204
rect 19704 3178 19728 3204
rect 19648 3159 19728 3178
rect 19648 3133 19667 3159
rect 19707 3133 19728 3159
rect 19648 3106 19728 3133
rect 19648 3080 19671 3106
rect 19711 3080 19728 3106
rect 19648 3069 19728 3080
rect 19790 3070 19817 3325
rect 20195 3317 20236 3467
rect 20467 3461 20571 3467
rect 20927 3464 20991 3467
rect 20662 3405 20783 3423
rect 20662 3403 20733 3405
rect 20662 3362 20677 3403
rect 20714 3364 20733 3403
rect 20770 3364 20783 3405
rect 20714 3362 20783 3364
rect 20662 3352 20783 3362
rect 19857 3210 19921 3222
rect 20197 3218 20234 3317
rect 20462 3307 20573 3320
rect 20462 3305 20504 3307
rect 20462 3285 20469 3305
rect 20488 3285 20504 3305
rect 20462 3277 20504 3285
rect 20532 3305 20573 3307
rect 20532 3285 20546 3305
rect 20565 3285 20573 3305
rect 20532 3277 20573 3285
rect 20462 3271 20573 3277
rect 20405 3249 20654 3271
rect 20405 3218 20442 3249
rect 20618 3247 20654 3249
rect 20618 3218 20655 3247
rect 19857 3209 19892 3210
rect 19834 3204 19892 3209
rect 19834 3184 19837 3204
rect 19857 3190 19892 3204
rect 19912 3190 19921 3210
rect 19857 3182 19921 3190
rect 19883 3181 19921 3182
rect 19884 3180 19921 3181
rect 19987 3214 20023 3215
rect 20095 3214 20131 3215
rect 19987 3206 20131 3214
rect 19987 3186 19995 3206
rect 20015 3186 20103 3206
rect 20123 3186 20131 3206
rect 19987 3180 20131 3186
rect 20197 3210 20235 3218
rect 20303 3214 20339 3215
rect 20197 3190 20206 3210
rect 20226 3190 20235 3210
rect 20197 3181 20235 3190
rect 20254 3207 20339 3214
rect 20254 3187 20261 3207
rect 20282 3206 20339 3207
rect 20282 3187 20311 3206
rect 20254 3186 20311 3187
rect 20331 3186 20339 3206
rect 20197 3180 20234 3181
rect 20254 3180 20339 3186
rect 20405 3210 20443 3218
rect 20516 3214 20552 3215
rect 20405 3190 20414 3210
rect 20434 3190 20443 3210
rect 20405 3181 20443 3190
rect 20467 3206 20552 3214
rect 20467 3186 20524 3206
rect 20544 3186 20552 3206
rect 20405 3180 20442 3181
rect 20467 3180 20552 3186
rect 20618 3210 20656 3218
rect 20618 3190 20627 3210
rect 20647 3190 20656 3210
rect 20711 3200 20776 3352
rect 20929 3326 20984 3464
rect 22225 3408 22284 3479
rect 23137 3478 23189 3481
rect 23137 3443 23145 3478
rect 23170 3443 23189 3478
rect 23214 3470 23236 3481
rect 23214 3469 24081 3470
rect 23214 3443 24082 3469
rect 23137 3433 24082 3443
rect 23137 3431 23236 3433
rect 22225 3390 22247 3408
rect 22265 3390 22284 3408
rect 22225 3368 22284 3390
rect 22492 3404 23024 3409
rect 22492 3384 23378 3404
rect 23398 3384 23401 3404
rect 24037 3400 24082 3433
rect 22492 3380 23401 3384
rect 22492 3333 22535 3380
rect 22985 3379 23401 3380
rect 24033 3380 24426 3400
rect 24446 3380 24449 3400
rect 22985 3378 23326 3379
rect 22642 3347 22752 3361
rect 22642 3344 22685 3347
rect 22642 3339 22646 3344
rect 22480 3332 22535 3333
rect 20618 3181 20656 3190
rect 20709 3193 20776 3200
rect 20618 3180 20655 3181
rect 20041 3159 20077 3180
rect 20467 3159 20498 3180
rect 20709 3172 20726 3193
rect 20762 3172 20776 3193
rect 20928 3213 20984 3326
rect 20928 3195 20947 3213
rect 20965 3195 20984 3213
rect 20928 3175 20984 3195
rect 22224 3309 22535 3332
rect 22224 3291 22249 3309
rect 22267 3297 22535 3309
rect 22564 3317 22646 3339
rect 22675 3317 22685 3344
rect 22713 3320 22720 3347
rect 22749 3339 22752 3347
rect 22749 3320 22814 3339
rect 22713 3317 22814 3320
rect 22564 3315 22814 3317
rect 22267 3291 22289 3297
rect 20709 3159 20776 3172
rect 19874 3155 19974 3159
rect 19874 3151 19936 3155
rect 19874 3125 19881 3151
rect 19907 3129 19936 3151
rect 19962 3129 19974 3155
rect 19907 3125 19974 3129
rect 19874 3122 19974 3125
rect 20042 3122 20077 3159
rect 20139 3156 20498 3159
rect 20139 3151 20361 3156
rect 20139 3127 20152 3151
rect 20176 3132 20361 3151
rect 20385 3132 20498 3156
rect 20176 3127 20498 3132
rect 20139 3123 20498 3127
rect 20565 3153 20776 3159
rect 20565 3151 20726 3153
rect 20565 3131 20576 3151
rect 20596 3131 20726 3151
rect 20565 3124 20726 3131
rect 20565 3123 20606 3124
rect 20041 3097 20077 3122
rect 19889 3070 19926 3071
rect 19985 3070 20022 3071
rect 20041 3070 20048 3097
rect 18199 3011 18614 3046
rect 19789 3061 19927 3070
rect 19789 3041 19898 3061
rect 19918 3041 19927 3061
rect 19789 3034 19927 3041
rect 19985 3067 20048 3070
rect 20069 3070 20077 3097
rect 20096 3070 20133 3071
rect 20069 3067 20133 3070
rect 19985 3061 20133 3067
rect 19985 3041 19994 3061
rect 20014 3041 20104 3061
rect 20124 3041 20133 3061
rect 19789 3032 19885 3034
rect 19985 3031 20133 3041
rect 20192 3061 20229 3071
rect 20304 3070 20341 3071
rect 20285 3068 20341 3070
rect 20192 3041 20200 3061
rect 20220 3041 20229 3061
rect 20041 3030 20077 3031
rect 18199 3010 18245 3011
rect 17905 2965 18155 2967
rect 17905 2962 18006 2965
rect 17905 2943 17970 2962
rect 17967 2935 17970 2943
rect 17999 2935 18006 2962
rect 18034 2938 18044 2965
rect 18073 2943 18155 2965
rect 18539 2959 18614 3011
rect 18073 2938 18077 2943
rect 18034 2935 18077 2938
rect 17967 2921 18077 2935
rect 17393 2903 17734 2904
rect 17318 2898 17734 2903
rect 17318 2878 17321 2898
rect 17341 2878 17735 2898
rect 13798 2469 16866 2494
rect 13798 2404 16661 2469
rect 16792 2404 16866 2469
rect 13798 2387 16866 2404
rect 17692 2374 17735 2878
rect 18352 2789 18447 2809
rect 18352 2745 18372 2789
rect 18432 2745 18447 2789
rect 18352 2449 18447 2745
rect 18352 2408 18385 2449
rect 18421 2408 18447 2449
rect 18547 2488 18609 2959
rect 19889 2899 19926 2900
rect 20192 2899 20229 3041
rect 20254 3061 20341 3068
rect 20254 3058 20312 3061
rect 20254 3038 20259 3058
rect 20280 3041 20312 3058
rect 20332 3041 20341 3061
rect 20280 3038 20341 3041
rect 20254 3031 20341 3038
rect 20400 3061 20437 3071
rect 20400 3041 20408 3061
rect 20428 3041 20437 3061
rect 20254 3030 20285 3031
rect 20400 2962 20437 3041
rect 20467 3070 20498 3123
rect 20711 3116 20726 3124
rect 20766 3116 20776 3153
rect 22224 3152 22289 3291
rect 22564 3236 22601 3315
rect 22642 3302 22752 3315
rect 22716 3246 22747 3247
rect 22564 3216 22573 3236
rect 22593 3216 22601 3236
rect 20711 3107 20776 3116
rect 20924 3114 20989 3135
rect 22224 3134 22247 3152
rect 22265 3134 22289 3152
rect 22224 3117 22289 3134
rect 22444 3198 22512 3211
rect 22564 3206 22601 3216
rect 22660 3236 22747 3246
rect 22660 3216 22669 3236
rect 22689 3216 22747 3236
rect 22660 3207 22747 3216
rect 22660 3206 22697 3207
rect 22444 3156 22451 3198
rect 22500 3156 22512 3198
rect 22444 3153 22512 3156
rect 22716 3154 22747 3207
rect 22777 3236 22814 3315
rect 22929 3246 22960 3247
rect 22777 3216 22786 3236
rect 22806 3216 22814 3236
rect 22777 3206 22814 3216
rect 22873 3239 22960 3246
rect 22873 3236 22934 3239
rect 22873 3216 22882 3236
rect 22902 3219 22934 3236
rect 22955 3219 22960 3239
rect 22902 3216 22960 3219
rect 22873 3209 22960 3216
rect 22985 3236 23022 3378
rect 23288 3377 23325 3378
rect 24033 3375 24449 3380
rect 24033 3374 24374 3375
rect 23690 3343 23800 3357
rect 23690 3340 23733 3343
rect 23690 3335 23694 3340
rect 23612 3313 23694 3335
rect 23723 3313 23733 3340
rect 23761 3316 23768 3343
rect 23797 3335 23800 3343
rect 23797 3316 23862 3335
rect 23761 3313 23862 3316
rect 23612 3311 23862 3313
rect 23137 3246 23173 3247
rect 22985 3216 22994 3236
rect 23014 3216 23022 3236
rect 22873 3207 22929 3209
rect 22873 3206 22910 3207
rect 22985 3206 23022 3216
rect 23081 3236 23229 3246
rect 23329 3243 23425 3245
rect 23081 3216 23090 3236
rect 23110 3216 23200 3236
rect 23220 3216 23229 3236
rect 23081 3210 23229 3216
rect 23081 3207 23145 3210
rect 23081 3206 23118 3207
rect 23137 3180 23145 3207
rect 23166 3207 23229 3210
rect 23287 3236 23425 3243
rect 23287 3216 23296 3236
rect 23316 3216 23425 3236
rect 23287 3207 23425 3216
rect 23612 3232 23649 3311
rect 23690 3298 23800 3311
rect 23764 3242 23795 3243
rect 23612 3212 23621 3232
rect 23641 3212 23649 3232
rect 23166 3180 23173 3207
rect 23192 3206 23229 3207
rect 23288 3206 23325 3207
rect 23137 3155 23173 3180
rect 22608 3153 22649 3154
rect 22444 3146 22649 3153
rect 22444 3135 22618 3146
rect 20924 3096 20949 3114
rect 20967 3096 20989 3114
rect 22444 3102 22452 3135
rect 20517 3070 20554 3071
rect 20467 3061 20554 3070
rect 20467 3041 20525 3061
rect 20545 3041 20554 3061
rect 20467 3031 20554 3041
rect 20613 3061 20650 3071
rect 20613 3041 20621 3061
rect 20641 3041 20650 3061
rect 20467 3030 20498 3031
rect 20462 2962 20572 2975
rect 20613 2962 20650 3041
rect 20924 3020 20989 3096
rect 22445 3093 22452 3102
rect 22501 3126 22618 3135
rect 22638 3126 22649 3146
rect 22501 3118 22649 3126
rect 22716 3150 23075 3154
rect 22716 3145 23038 3150
rect 22716 3121 22829 3145
rect 22853 3126 23038 3145
rect 23062 3126 23075 3150
rect 22853 3121 23075 3126
rect 22716 3118 23075 3121
rect 23137 3118 23172 3155
rect 23240 3152 23340 3155
rect 23240 3148 23307 3152
rect 23240 3122 23252 3148
rect 23278 3126 23307 3148
rect 23333 3126 23340 3152
rect 23278 3122 23340 3126
rect 23240 3118 23340 3122
rect 22501 3102 22512 3118
rect 22501 3093 22509 3102
rect 22716 3097 22747 3118
rect 23137 3097 23173 3118
rect 22559 3096 22596 3097
rect 22224 3053 22289 3072
rect 22224 3035 22249 3053
rect 22267 3035 22289 3053
rect 20400 2960 20650 2962
rect 20400 2957 20501 2960
rect 20400 2938 20465 2957
rect 20462 2930 20465 2938
rect 20494 2930 20501 2957
rect 20529 2933 20539 2960
rect 20568 2938 20650 2960
rect 20673 2985 20990 3020
rect 20568 2933 20572 2938
rect 20529 2930 20572 2933
rect 20462 2916 20572 2930
rect 19888 2898 20229 2899
rect 19813 2896 20229 2898
rect 20673 2896 20713 2985
rect 20924 2958 20989 2985
rect 20924 2940 20947 2958
rect 20965 2940 20989 2958
rect 20924 2920 20989 2940
rect 19810 2893 20713 2896
rect 19810 2873 19816 2893
rect 19836 2873 20713 2893
rect 19810 2869 20713 2873
rect 20673 2866 20713 2869
rect 20925 2859 20990 2880
rect 19143 2851 19804 2852
rect 19143 2844 20077 2851
rect 19143 2843 20049 2844
rect 19143 2823 19994 2843
rect 20026 2824 20049 2843
rect 20074 2824 20077 2844
rect 20026 2823 20077 2824
rect 19143 2816 20077 2823
rect 18742 2774 18910 2775
rect 19145 2774 19184 2816
rect 19973 2814 20077 2816
rect 20042 2812 20077 2814
rect 20925 2841 20949 2859
rect 20967 2841 20990 2859
rect 20925 2794 20990 2841
rect 18742 2748 19186 2774
rect 18742 2746 18910 2748
rect 18547 2469 18611 2488
rect 18547 2430 18564 2469
rect 18598 2430 18611 2469
rect 18547 2411 18611 2430
rect 18352 2382 18447 2408
rect 18742 2395 18769 2746
rect 19145 2742 19186 2748
rect 18809 2535 18873 2547
rect 19149 2543 19186 2742
rect 19648 2769 19720 2786
rect 19648 2730 19656 2769
rect 19701 2730 19720 2769
rect 19414 2632 19525 2647
rect 19414 2630 19456 2632
rect 19414 2610 19421 2630
rect 19440 2610 19456 2630
rect 19414 2602 19456 2610
rect 19484 2630 19525 2632
rect 19484 2610 19498 2630
rect 19517 2610 19525 2630
rect 19484 2602 19525 2610
rect 19414 2596 19525 2602
rect 19357 2574 19606 2596
rect 19357 2543 19394 2574
rect 19570 2572 19606 2574
rect 19570 2543 19607 2572
rect 18809 2534 18844 2535
rect 18786 2529 18844 2534
rect 18786 2509 18789 2529
rect 18809 2515 18844 2529
rect 18864 2515 18873 2535
rect 18809 2507 18873 2515
rect 18835 2506 18873 2507
rect 18836 2505 18873 2506
rect 18939 2539 18975 2540
rect 19047 2539 19083 2540
rect 18939 2531 19083 2539
rect 18939 2511 18947 2531
rect 18967 2511 19055 2531
rect 19075 2511 19083 2531
rect 18939 2505 19083 2511
rect 19149 2535 19187 2543
rect 19255 2539 19291 2540
rect 19149 2515 19158 2535
rect 19178 2515 19187 2535
rect 19149 2506 19187 2515
rect 19206 2532 19291 2539
rect 19206 2512 19213 2532
rect 19234 2531 19291 2532
rect 19234 2512 19263 2531
rect 19206 2511 19263 2512
rect 19283 2511 19291 2531
rect 19149 2505 19186 2506
rect 19206 2505 19291 2511
rect 19357 2535 19395 2543
rect 19468 2539 19504 2540
rect 19357 2515 19366 2535
rect 19386 2515 19395 2535
rect 19357 2506 19395 2515
rect 19419 2531 19504 2539
rect 19419 2511 19476 2531
rect 19496 2511 19504 2531
rect 19357 2505 19394 2506
rect 19419 2505 19504 2511
rect 19570 2535 19608 2543
rect 19570 2515 19579 2535
rect 19599 2515 19608 2535
rect 19570 2506 19608 2515
rect 19648 2520 19720 2730
rect 19790 2764 20990 2794
rect 19790 2763 20234 2764
rect 19790 2761 19958 2763
rect 19648 2506 19731 2520
rect 19570 2505 19607 2506
rect 18993 2484 19029 2505
rect 19419 2484 19450 2505
rect 19648 2484 19665 2506
rect 18826 2480 18926 2484
rect 18826 2476 18888 2480
rect 18826 2450 18833 2476
rect 18859 2454 18888 2476
rect 18914 2454 18926 2480
rect 18859 2450 18926 2454
rect 18826 2447 18926 2450
rect 18994 2447 19029 2484
rect 19091 2481 19450 2484
rect 19091 2476 19313 2481
rect 19091 2452 19104 2476
rect 19128 2457 19313 2476
rect 19337 2457 19450 2481
rect 19128 2452 19450 2457
rect 19091 2448 19450 2452
rect 19517 2476 19665 2484
rect 19517 2456 19528 2476
rect 19548 2473 19665 2476
rect 19718 2473 19731 2506
rect 19548 2456 19731 2473
rect 19517 2449 19731 2456
rect 19517 2448 19558 2449
rect 19648 2448 19731 2449
rect 18993 2422 19029 2447
rect 18841 2395 18878 2396
rect 18937 2395 18974 2396
rect 18993 2395 19000 2422
rect 18741 2386 18879 2395
rect 13553 2288 13710 2301
rect 13553 2284 13714 2288
rect 12433 2138 12459 2243
rect 13553 2177 13594 2284
rect 13694 2177 13714 2284
rect 13553 2148 13714 2177
rect 17690 2165 17739 2374
rect 18741 2366 18850 2386
rect 18870 2366 18879 2386
rect 18741 2359 18879 2366
rect 18937 2392 19000 2395
rect 19021 2395 19029 2422
rect 19048 2395 19085 2396
rect 19021 2392 19085 2395
rect 18937 2386 19085 2392
rect 18937 2366 18946 2386
rect 18966 2366 19056 2386
rect 19076 2366 19085 2386
rect 18741 2357 18837 2359
rect 18937 2356 19085 2366
rect 19144 2386 19181 2396
rect 19256 2395 19293 2396
rect 19237 2393 19293 2395
rect 19144 2366 19152 2386
rect 19172 2366 19181 2386
rect 18993 2355 19029 2356
rect 18841 2224 18878 2225
rect 19144 2224 19181 2366
rect 19206 2386 19293 2393
rect 19206 2383 19264 2386
rect 19206 2363 19211 2383
rect 19232 2366 19264 2383
rect 19284 2366 19293 2386
rect 19232 2363 19293 2366
rect 19206 2356 19293 2363
rect 19352 2386 19389 2396
rect 19352 2366 19360 2386
rect 19380 2366 19389 2386
rect 19206 2355 19237 2356
rect 19352 2287 19389 2366
rect 19419 2395 19450 2448
rect 19656 2415 19670 2448
rect 19723 2415 19731 2448
rect 19656 2409 19731 2415
rect 19656 2404 19726 2409
rect 19469 2395 19506 2396
rect 19419 2386 19506 2395
rect 19419 2366 19477 2386
rect 19497 2366 19506 2386
rect 19419 2356 19506 2366
rect 19565 2386 19602 2396
rect 19790 2391 19817 2761
rect 19857 2531 19921 2543
rect 20197 2539 20234 2763
rect 20705 2744 20769 2746
rect 20701 2732 20769 2744
rect 20701 2699 20712 2732
rect 20752 2699 20769 2732
rect 20701 2689 20769 2699
rect 20462 2628 20573 2643
rect 20462 2626 20504 2628
rect 20462 2606 20469 2626
rect 20488 2606 20504 2626
rect 20462 2598 20504 2606
rect 20532 2626 20573 2628
rect 20532 2606 20546 2626
rect 20565 2606 20573 2626
rect 20532 2598 20573 2606
rect 20462 2592 20573 2598
rect 20405 2570 20654 2592
rect 20405 2539 20442 2570
rect 20618 2568 20654 2570
rect 20618 2539 20655 2568
rect 19857 2530 19892 2531
rect 19834 2525 19892 2530
rect 19834 2505 19837 2525
rect 19857 2511 19892 2525
rect 19912 2511 19921 2531
rect 19857 2503 19921 2511
rect 19883 2502 19921 2503
rect 19884 2501 19921 2502
rect 19987 2535 20023 2536
rect 20095 2535 20131 2536
rect 19987 2527 20131 2535
rect 19987 2507 19995 2527
rect 20015 2507 20103 2527
rect 20123 2507 20131 2527
rect 19987 2501 20131 2507
rect 20197 2531 20235 2539
rect 20303 2535 20339 2536
rect 20197 2511 20206 2531
rect 20226 2511 20235 2531
rect 20197 2502 20235 2511
rect 20254 2528 20339 2535
rect 20254 2508 20261 2528
rect 20282 2527 20339 2528
rect 20282 2508 20311 2527
rect 20254 2507 20311 2508
rect 20331 2507 20339 2527
rect 20197 2501 20234 2502
rect 20254 2501 20339 2507
rect 20405 2531 20443 2539
rect 20516 2535 20552 2536
rect 20405 2511 20414 2531
rect 20434 2511 20443 2531
rect 20405 2502 20443 2511
rect 20467 2527 20552 2535
rect 20467 2507 20524 2527
rect 20544 2507 20552 2527
rect 20405 2501 20442 2502
rect 20467 2501 20552 2507
rect 20618 2531 20656 2539
rect 20618 2511 20627 2531
rect 20647 2511 20656 2531
rect 20618 2502 20656 2511
rect 20705 2505 20769 2689
rect 20925 2563 20990 2764
rect 22224 2834 22289 3035
rect 22445 2909 22509 3093
rect 22558 3087 22596 3096
rect 22558 3067 22567 3087
rect 22587 3067 22596 3087
rect 22558 3059 22596 3067
rect 22662 3091 22747 3097
rect 22772 3096 22809 3097
rect 22662 3071 22670 3091
rect 22690 3071 22747 3091
rect 22662 3063 22747 3071
rect 22771 3087 22809 3096
rect 22771 3067 22780 3087
rect 22800 3067 22809 3087
rect 22662 3062 22698 3063
rect 22771 3059 22809 3067
rect 22875 3091 22960 3097
rect 22980 3096 23017 3097
rect 22875 3071 22883 3091
rect 22903 3090 22960 3091
rect 22903 3071 22932 3090
rect 22875 3070 22932 3071
rect 22953 3070 22960 3090
rect 22875 3063 22960 3070
rect 22979 3087 23017 3096
rect 22979 3067 22988 3087
rect 23008 3067 23017 3087
rect 22875 3062 22911 3063
rect 22979 3059 23017 3067
rect 23083 3091 23227 3097
rect 23083 3071 23091 3091
rect 23111 3071 23199 3091
rect 23219 3071 23227 3091
rect 23083 3063 23227 3071
rect 23083 3062 23119 3063
rect 23191 3062 23227 3063
rect 23293 3096 23330 3097
rect 23293 3095 23331 3096
rect 23293 3087 23357 3095
rect 23293 3067 23302 3087
rect 23322 3073 23357 3087
rect 23377 3073 23380 3093
rect 23322 3068 23380 3073
rect 23322 3067 23357 3068
rect 22559 3030 22596 3059
rect 22560 3028 22596 3030
rect 22772 3028 22809 3059
rect 22560 3006 22809 3028
rect 22641 3000 22752 3006
rect 22641 2992 22682 3000
rect 22641 2972 22649 2992
rect 22668 2972 22682 2992
rect 22641 2970 22682 2972
rect 22710 2992 22752 3000
rect 22710 2972 22726 2992
rect 22745 2972 22752 2992
rect 22710 2970 22752 2972
rect 22641 2955 22752 2970
rect 22445 2899 22513 2909
rect 22445 2866 22462 2899
rect 22502 2866 22513 2899
rect 22445 2854 22513 2866
rect 22445 2852 22509 2854
rect 22980 2835 23017 3059
rect 23293 3055 23357 3067
rect 23397 2837 23424 3207
rect 23612 3202 23649 3212
rect 23708 3232 23795 3242
rect 23708 3212 23717 3232
rect 23737 3212 23795 3232
rect 23708 3203 23795 3212
rect 23708 3202 23745 3203
rect 23488 3189 23558 3194
rect 23483 3183 23558 3189
rect 23483 3150 23491 3183
rect 23544 3150 23558 3183
rect 23764 3150 23795 3203
rect 23825 3232 23862 3311
rect 23977 3242 24008 3243
rect 23825 3212 23834 3232
rect 23854 3212 23862 3232
rect 23825 3202 23862 3212
rect 23921 3235 24008 3242
rect 23921 3232 23982 3235
rect 23921 3212 23930 3232
rect 23950 3215 23982 3232
rect 24003 3215 24008 3235
rect 23950 3212 24008 3215
rect 23921 3205 24008 3212
rect 24033 3232 24070 3374
rect 24336 3373 24373 3374
rect 24185 3242 24221 3243
rect 24033 3212 24042 3232
rect 24062 3212 24070 3232
rect 23921 3203 23977 3205
rect 23921 3202 23958 3203
rect 24033 3202 24070 3212
rect 24129 3232 24277 3242
rect 24377 3239 24473 3241
rect 24129 3212 24138 3232
rect 24158 3212 24248 3232
rect 24268 3212 24277 3232
rect 24129 3206 24277 3212
rect 24129 3203 24193 3206
rect 24129 3202 24166 3203
rect 24185 3176 24193 3203
rect 24214 3203 24277 3206
rect 24335 3232 24473 3239
rect 24335 3212 24344 3232
rect 24364 3212 24473 3232
rect 24335 3203 24473 3212
rect 24214 3176 24221 3203
rect 24240 3202 24277 3203
rect 24336 3202 24373 3203
rect 24185 3151 24221 3176
rect 23483 3149 23566 3150
rect 23656 3149 23697 3150
rect 23483 3142 23697 3149
rect 23483 3125 23666 3142
rect 23483 3092 23496 3125
rect 23549 3122 23666 3125
rect 23686 3122 23697 3142
rect 23549 3114 23697 3122
rect 23764 3146 24123 3150
rect 23764 3141 24086 3146
rect 23764 3117 23877 3141
rect 23901 3122 24086 3141
rect 24110 3122 24123 3146
rect 23901 3117 24123 3122
rect 23764 3114 24123 3117
rect 24185 3114 24220 3151
rect 24288 3148 24388 3151
rect 24288 3144 24355 3148
rect 24288 3118 24300 3144
rect 24326 3122 24355 3144
rect 24381 3122 24388 3148
rect 24326 3118 24388 3122
rect 24288 3114 24388 3118
rect 23549 3092 23566 3114
rect 23764 3093 23795 3114
rect 24185 3093 24221 3114
rect 23607 3092 23644 3093
rect 23483 3078 23566 3092
rect 23256 2835 23424 2837
rect 22980 2834 23424 2835
rect 22224 2804 23424 2834
rect 23494 2868 23566 3078
rect 23606 3083 23644 3092
rect 23606 3063 23615 3083
rect 23635 3063 23644 3083
rect 23606 3055 23644 3063
rect 23710 3087 23795 3093
rect 23820 3092 23857 3093
rect 23710 3067 23718 3087
rect 23738 3067 23795 3087
rect 23710 3059 23795 3067
rect 23819 3083 23857 3092
rect 23819 3063 23828 3083
rect 23848 3063 23857 3083
rect 23710 3058 23746 3059
rect 23819 3055 23857 3063
rect 23923 3087 24008 3093
rect 24028 3092 24065 3093
rect 23923 3067 23931 3087
rect 23951 3086 24008 3087
rect 23951 3067 23980 3086
rect 23923 3066 23980 3067
rect 24001 3066 24008 3086
rect 23923 3059 24008 3066
rect 24027 3083 24065 3092
rect 24027 3063 24036 3083
rect 24056 3063 24065 3083
rect 23923 3058 23959 3059
rect 24027 3055 24065 3063
rect 24131 3087 24275 3093
rect 24131 3067 24139 3087
rect 24159 3067 24247 3087
rect 24267 3067 24275 3087
rect 24131 3059 24275 3067
rect 24131 3058 24167 3059
rect 24239 3058 24275 3059
rect 24341 3092 24378 3093
rect 24341 3091 24379 3092
rect 24341 3083 24405 3091
rect 24341 3063 24350 3083
rect 24370 3069 24405 3083
rect 24425 3069 24428 3089
rect 24370 3064 24428 3069
rect 24370 3063 24405 3064
rect 23607 3026 23644 3055
rect 23608 3024 23644 3026
rect 23820 3024 23857 3055
rect 23608 3002 23857 3024
rect 23689 2996 23800 3002
rect 23689 2988 23730 2996
rect 23689 2968 23697 2988
rect 23716 2968 23730 2988
rect 23689 2966 23730 2968
rect 23758 2988 23800 2996
rect 23758 2968 23774 2988
rect 23793 2968 23800 2988
rect 23758 2966 23800 2968
rect 23689 2951 23800 2966
rect 23494 2829 23513 2868
rect 23558 2829 23566 2868
rect 23494 2812 23566 2829
rect 24028 2856 24065 3055
rect 24341 3051 24405 3063
rect 24028 2850 24069 2856
rect 24445 2852 24472 3203
rect 24304 2850 24472 2852
rect 24028 2824 24472 2850
rect 22224 2757 22289 2804
rect 22224 2739 22247 2757
rect 22265 2739 22289 2757
rect 23137 2784 23172 2786
rect 23137 2782 23241 2784
rect 24030 2782 24069 2824
rect 24304 2823 24472 2824
rect 23137 2775 24071 2782
rect 23137 2774 23188 2775
rect 23137 2754 23140 2774
rect 23165 2755 23188 2774
rect 23220 2755 24071 2775
rect 23165 2754 24071 2755
rect 23137 2747 24071 2754
rect 23410 2746 24071 2747
rect 22224 2718 22289 2739
rect 22501 2729 22541 2732
rect 22501 2725 23404 2729
rect 22501 2705 23378 2725
rect 23398 2705 23404 2725
rect 22501 2702 23404 2705
rect 22225 2658 22290 2678
rect 22225 2640 22249 2658
rect 22267 2640 22290 2658
rect 22225 2613 22290 2640
rect 22501 2613 22541 2702
rect 22985 2700 23401 2702
rect 22985 2699 23326 2700
rect 22642 2668 22752 2682
rect 22642 2665 22685 2668
rect 22642 2660 22646 2665
rect 22224 2578 22541 2613
rect 22564 2638 22646 2660
rect 22675 2638 22685 2665
rect 22713 2641 22720 2668
rect 22749 2660 22752 2668
rect 22749 2641 22814 2660
rect 22713 2638 22814 2641
rect 22564 2636 22814 2638
rect 20925 2545 20947 2563
rect 20965 2545 20990 2563
rect 20925 2526 20990 2545
rect 20618 2501 20655 2502
rect 20041 2480 20077 2501
rect 20467 2480 20498 2501
rect 20705 2496 20713 2505
rect 20702 2480 20713 2496
rect 19874 2476 19974 2480
rect 19874 2472 19936 2476
rect 19874 2446 19881 2472
rect 19907 2450 19936 2472
rect 19962 2450 19974 2476
rect 19907 2446 19974 2450
rect 19874 2443 19974 2446
rect 20042 2443 20077 2480
rect 20139 2477 20498 2480
rect 20139 2472 20361 2477
rect 20139 2448 20152 2472
rect 20176 2453 20361 2472
rect 20385 2453 20498 2477
rect 20176 2448 20498 2453
rect 20139 2444 20498 2448
rect 20565 2472 20713 2480
rect 20565 2452 20576 2472
rect 20596 2463 20713 2472
rect 20762 2496 20769 2505
rect 22225 2502 22290 2578
rect 22564 2557 22601 2636
rect 22642 2623 22752 2636
rect 22716 2567 22747 2568
rect 22564 2537 22573 2557
rect 22593 2537 22601 2557
rect 22564 2527 22601 2537
rect 22660 2557 22747 2567
rect 22660 2537 22669 2557
rect 22689 2537 22747 2557
rect 22660 2528 22747 2537
rect 22660 2527 22697 2528
rect 20762 2463 20770 2496
rect 22225 2484 22247 2502
rect 22265 2484 22290 2502
rect 20596 2452 20770 2463
rect 20565 2445 20770 2452
rect 20565 2444 20606 2445
rect 20041 2418 20077 2443
rect 19889 2391 19926 2392
rect 19985 2391 20022 2392
rect 20041 2391 20048 2418
rect 19565 2366 19573 2386
rect 19593 2366 19602 2386
rect 19419 2355 19450 2356
rect 19414 2287 19524 2300
rect 19565 2287 19602 2366
rect 19789 2382 19927 2391
rect 19789 2362 19898 2382
rect 19918 2362 19927 2382
rect 19789 2355 19927 2362
rect 19985 2388 20048 2391
rect 20069 2391 20077 2418
rect 20096 2391 20133 2392
rect 20069 2388 20133 2391
rect 19985 2382 20133 2388
rect 19985 2362 19994 2382
rect 20014 2362 20104 2382
rect 20124 2362 20133 2382
rect 19789 2353 19885 2355
rect 19985 2352 20133 2362
rect 20192 2382 20229 2392
rect 20304 2391 20341 2392
rect 20285 2389 20341 2391
rect 20192 2362 20200 2382
rect 20220 2362 20229 2382
rect 20041 2351 20077 2352
rect 19352 2285 19602 2287
rect 19352 2282 19453 2285
rect 19352 2263 19417 2282
rect 19414 2255 19417 2263
rect 19446 2255 19453 2282
rect 19481 2258 19491 2285
rect 19520 2263 19602 2285
rect 19520 2258 19524 2263
rect 19481 2255 19524 2258
rect 19414 2241 19524 2255
rect 18840 2223 19181 2224
rect 18765 2218 19181 2223
rect 19889 2220 19926 2221
rect 20192 2220 20229 2362
rect 20254 2382 20341 2389
rect 20254 2379 20312 2382
rect 20254 2359 20259 2379
rect 20280 2362 20312 2379
rect 20332 2362 20341 2382
rect 20280 2359 20341 2362
rect 20254 2352 20341 2359
rect 20400 2382 20437 2392
rect 20400 2362 20408 2382
rect 20428 2362 20437 2382
rect 20254 2351 20285 2352
rect 20400 2283 20437 2362
rect 20467 2391 20498 2444
rect 20702 2442 20770 2445
rect 20702 2400 20714 2442
rect 20763 2400 20770 2442
rect 20517 2391 20554 2392
rect 20467 2382 20554 2391
rect 20467 2362 20525 2382
rect 20545 2362 20554 2382
rect 20467 2352 20554 2362
rect 20613 2382 20650 2392
rect 20702 2387 20770 2400
rect 20925 2464 20990 2481
rect 20925 2446 20949 2464
rect 20967 2446 20990 2464
rect 22225 2463 22290 2484
rect 22438 2482 22503 2491
rect 20613 2362 20621 2382
rect 20641 2362 20650 2382
rect 20467 2351 20498 2352
rect 20462 2283 20572 2296
rect 20613 2283 20650 2362
rect 20925 2307 20990 2446
rect 22438 2445 22448 2482
rect 22488 2474 22503 2482
rect 22716 2475 22747 2528
rect 22777 2557 22814 2636
rect 22929 2567 22960 2568
rect 22777 2537 22786 2557
rect 22806 2537 22814 2557
rect 22777 2527 22814 2537
rect 22873 2560 22960 2567
rect 22873 2557 22934 2560
rect 22873 2537 22882 2557
rect 22902 2540 22934 2557
rect 22955 2540 22960 2560
rect 22902 2537 22960 2540
rect 22873 2530 22960 2537
rect 22985 2557 23022 2699
rect 23288 2698 23325 2699
rect 23137 2567 23173 2568
rect 22985 2537 22994 2557
rect 23014 2537 23022 2557
rect 22873 2528 22929 2530
rect 22873 2527 22910 2528
rect 22985 2527 23022 2537
rect 23081 2557 23229 2567
rect 23329 2564 23425 2566
rect 23081 2537 23090 2557
rect 23110 2537 23200 2557
rect 23220 2537 23229 2557
rect 23081 2531 23229 2537
rect 23081 2528 23145 2531
rect 23081 2527 23118 2528
rect 23137 2501 23145 2528
rect 23166 2528 23229 2531
rect 23287 2557 23425 2564
rect 23287 2537 23296 2557
rect 23316 2537 23425 2557
rect 23287 2528 23425 2537
rect 23166 2501 23173 2528
rect 23192 2527 23229 2528
rect 23288 2527 23325 2528
rect 23137 2476 23173 2501
rect 22608 2474 22649 2475
rect 22488 2467 22649 2474
rect 22488 2447 22618 2467
rect 22638 2447 22649 2467
rect 22488 2445 22649 2447
rect 22438 2439 22649 2445
rect 22716 2471 23075 2475
rect 22716 2466 23038 2471
rect 22716 2442 22829 2466
rect 22853 2447 23038 2466
rect 23062 2447 23075 2471
rect 22853 2442 23075 2447
rect 22716 2439 23075 2442
rect 23137 2439 23172 2476
rect 23240 2473 23340 2476
rect 23240 2469 23307 2473
rect 23240 2443 23252 2469
rect 23278 2447 23307 2469
rect 23333 2447 23340 2473
rect 23278 2443 23340 2447
rect 23240 2439 23340 2443
rect 22438 2426 22505 2439
rect 22230 2403 22286 2423
rect 22230 2385 22249 2403
rect 22267 2385 22286 2403
rect 22230 2350 22286 2385
rect 20925 2301 20947 2307
rect 20400 2281 20650 2283
rect 20400 2278 20501 2281
rect 20400 2259 20465 2278
rect 20462 2251 20465 2259
rect 20494 2251 20501 2278
rect 20529 2254 20539 2281
rect 20568 2259 20650 2281
rect 20679 2289 20947 2301
rect 20965 2289 20990 2307
rect 20679 2266 20990 2289
rect 22192 2272 22286 2350
rect 22438 2405 22452 2426
rect 22488 2405 22505 2426
rect 22716 2418 22747 2439
rect 23137 2418 23173 2439
rect 22559 2417 22596 2418
rect 22438 2398 22505 2405
rect 22558 2408 22596 2417
rect 20679 2265 20734 2266
rect 20568 2254 20572 2259
rect 20529 2251 20572 2254
rect 20462 2237 20572 2251
rect 19888 2219 20229 2220
rect 18765 2198 18768 2218
rect 18788 2198 19181 2218
rect 19813 2218 20229 2219
rect 20679 2218 20722 2265
rect 19813 2214 20722 2218
rect 12433 2124 12461 2138
rect 13557 2135 13714 2148
rect 17688 2163 18505 2165
rect 18938 2163 19027 2166
rect 17688 2154 19027 2163
rect 11235 2089 12461 2124
rect 17688 2116 18950 2154
rect 18975 2119 18994 2154
rect 19019 2119 19027 2154
rect 19132 2165 19177 2198
rect 19813 2194 19816 2214
rect 19836 2194 20722 2214
rect 20190 2189 20722 2194
rect 20930 2208 20989 2230
rect 20930 2190 20949 2208
rect 20967 2190 20989 2208
rect 19978 2165 20077 2167
rect 19132 2155 20077 2165
rect 19132 2129 20000 2155
rect 19133 2128 20000 2129
rect 18975 2116 19027 2119
rect 17688 2108 19027 2116
rect 19978 2117 20000 2128
rect 20025 2120 20044 2155
rect 20069 2120 20077 2155
rect 20025 2117 20077 2120
rect 19978 2109 20077 2117
rect 20004 2108 20076 2109
rect 17688 2107 19026 2108
rect 17688 2105 18505 2107
rect 18279 2101 18505 2105
rect 527 1946 10295 2019
rect 541 1931 10295 1946
rect 11235 2013 11320 2089
rect 11678 2087 11782 2089
rect 12013 2087 12054 2089
rect 20930 2013 20989 2190
rect 22192 2131 22285 2272
rect 22438 2246 22503 2398
rect 22558 2388 22567 2408
rect 22587 2388 22596 2408
rect 22558 2380 22596 2388
rect 22662 2412 22747 2418
rect 22772 2417 22809 2418
rect 22662 2392 22670 2412
rect 22690 2392 22747 2412
rect 22662 2384 22747 2392
rect 22771 2408 22809 2417
rect 22771 2388 22780 2408
rect 22800 2388 22809 2408
rect 22662 2383 22698 2384
rect 22771 2380 22809 2388
rect 22875 2412 22960 2418
rect 22980 2417 23017 2418
rect 22875 2392 22883 2412
rect 22903 2411 22960 2412
rect 22903 2392 22932 2411
rect 22875 2391 22932 2392
rect 22953 2391 22960 2411
rect 22875 2384 22960 2391
rect 22979 2408 23017 2417
rect 22979 2388 22988 2408
rect 23008 2388 23017 2408
rect 22875 2383 22911 2384
rect 22979 2380 23017 2388
rect 23083 2412 23227 2418
rect 23083 2392 23091 2412
rect 23111 2392 23199 2412
rect 23219 2392 23227 2412
rect 23083 2384 23227 2392
rect 23083 2383 23119 2384
rect 23191 2383 23227 2384
rect 23293 2417 23330 2418
rect 23293 2416 23331 2417
rect 23293 2408 23357 2416
rect 23293 2388 23302 2408
rect 23322 2394 23357 2408
rect 23377 2394 23380 2414
rect 23322 2389 23380 2394
rect 23322 2388 23357 2389
rect 22559 2351 22596 2380
rect 22560 2349 22596 2351
rect 22772 2349 22809 2380
rect 22560 2327 22809 2349
rect 22641 2321 22752 2327
rect 22641 2313 22682 2321
rect 22641 2293 22649 2313
rect 22668 2293 22682 2313
rect 22641 2291 22682 2293
rect 22710 2313 22752 2321
rect 22710 2293 22726 2313
rect 22745 2293 22752 2313
rect 22710 2291 22752 2293
rect 22641 2276 22752 2291
rect 22980 2281 23017 2380
rect 23293 2376 23357 2388
rect 23397 2337 23424 2528
rect 22643 2267 22747 2276
rect 22431 2236 22552 2246
rect 22431 2234 22500 2236
rect 22431 2193 22444 2234
rect 22481 2195 22500 2234
rect 22537 2195 22552 2236
rect 22481 2193 22552 2195
rect 22431 2175 22552 2193
rect 22643 2131 22747 2140
rect 22978 2131 23019 2281
rect 22192 2129 23019 2131
rect 22200 2128 23019 2129
rect 23398 2247 23423 2337
rect 24558 2305 24657 3862
rect 24763 2498 24862 5399
rect 25253 5382 25284 5403
rect 25674 5382 25710 5403
rect 25096 5381 25133 5382
rect 25095 5372 25133 5381
rect 25095 5352 25104 5372
rect 25124 5352 25133 5372
rect 25095 5344 25133 5352
rect 25199 5376 25284 5382
rect 25309 5381 25346 5382
rect 25199 5356 25207 5376
rect 25227 5356 25284 5376
rect 25199 5348 25284 5356
rect 25308 5372 25346 5381
rect 25308 5352 25317 5372
rect 25337 5352 25346 5372
rect 25199 5347 25235 5348
rect 25308 5344 25346 5352
rect 25412 5376 25497 5382
rect 25517 5381 25554 5382
rect 25412 5356 25420 5376
rect 25440 5375 25497 5376
rect 25440 5356 25469 5375
rect 25412 5355 25469 5356
rect 25490 5355 25497 5375
rect 25412 5348 25497 5355
rect 25516 5372 25554 5381
rect 25516 5352 25525 5372
rect 25545 5352 25554 5372
rect 25412 5347 25448 5348
rect 25516 5344 25554 5352
rect 25620 5376 25764 5382
rect 25620 5356 25628 5376
rect 25648 5356 25736 5376
rect 25756 5356 25764 5376
rect 25620 5348 25764 5356
rect 25620 5347 25656 5348
rect 25728 5347 25764 5348
rect 25830 5381 25867 5382
rect 25830 5380 25868 5381
rect 25830 5372 25894 5380
rect 25830 5352 25839 5372
rect 25859 5358 25894 5372
rect 25914 5358 25917 5378
rect 25859 5353 25917 5358
rect 25859 5352 25894 5353
rect 25096 5315 25133 5344
rect 25097 5313 25133 5315
rect 25309 5313 25346 5344
rect 25097 5291 25346 5313
rect 25178 5285 25289 5291
rect 25178 5277 25219 5285
rect 25178 5257 25186 5277
rect 25205 5257 25219 5277
rect 25178 5255 25219 5257
rect 25247 5277 25289 5285
rect 25247 5257 25263 5277
rect 25282 5257 25289 5277
rect 25247 5255 25289 5257
rect 25178 5240 25289 5255
rect 25517 5223 25554 5344
rect 25830 5340 25894 5352
rect 25635 5223 25664 5227
rect 25934 5225 25961 5492
rect 25793 5223 25961 5225
rect 25517 5197 25961 5223
rect 25476 4929 25521 4938
rect 25476 4891 25486 4929
rect 25511 4891 25521 4929
rect 25476 4880 25521 4891
rect 25479 4872 25521 4880
rect 25479 4167 25522 4872
rect 25635 4258 25664 5197
rect 25793 5196 25961 5197
rect 26365 5047 26449 5051
rect 26917 5047 27005 7898
rect 27544 7885 27599 7897
rect 27544 7851 27562 7885
rect 27591 7851 27599 7885
rect 27544 7825 27599 7851
rect 27151 7792 27319 7793
rect 27544 7792 27561 7825
rect 27151 7791 27561 7792
rect 27590 7791 27599 7825
rect 27151 7766 27599 7791
rect 27151 7764 27319 7766
rect 27151 7497 27178 7764
rect 27544 7760 27599 7766
rect 27218 7637 27282 7649
rect 27558 7645 27595 7760
rect 27823 7734 27934 7749
rect 27823 7732 27865 7734
rect 27823 7712 27830 7732
rect 27849 7712 27865 7732
rect 27823 7704 27865 7712
rect 27893 7732 27934 7734
rect 27893 7712 27907 7732
rect 27926 7712 27934 7732
rect 27893 7704 27934 7712
rect 27823 7698 27934 7704
rect 27766 7676 28015 7698
rect 27766 7645 27803 7676
rect 27979 7674 28015 7676
rect 27979 7645 28016 7674
rect 27218 7636 27253 7637
rect 27195 7631 27253 7636
rect 27195 7611 27198 7631
rect 27218 7617 27253 7631
rect 27273 7617 27282 7637
rect 27218 7609 27282 7617
rect 27244 7608 27282 7609
rect 27245 7607 27282 7608
rect 27348 7641 27384 7642
rect 27456 7641 27492 7642
rect 27348 7633 27492 7641
rect 27348 7613 27356 7633
rect 27376 7613 27464 7633
rect 27484 7613 27492 7633
rect 27348 7607 27492 7613
rect 27558 7637 27596 7645
rect 27664 7641 27700 7642
rect 27558 7617 27567 7637
rect 27587 7617 27596 7637
rect 27558 7608 27596 7617
rect 27615 7634 27700 7641
rect 27615 7614 27622 7634
rect 27643 7633 27700 7634
rect 27643 7614 27672 7633
rect 27615 7613 27672 7614
rect 27692 7613 27700 7633
rect 27558 7607 27595 7608
rect 27615 7607 27700 7613
rect 27766 7637 27804 7645
rect 27877 7641 27913 7642
rect 27766 7617 27775 7637
rect 27795 7617 27804 7637
rect 27766 7608 27804 7617
rect 27828 7633 27913 7641
rect 27828 7613 27885 7633
rect 27905 7613 27913 7633
rect 27766 7607 27803 7608
rect 27828 7607 27913 7613
rect 27979 7637 28017 7645
rect 27979 7617 27988 7637
rect 28008 7617 28017 7637
rect 27979 7608 28017 7617
rect 27979 7607 28016 7608
rect 27402 7586 27438 7607
rect 27828 7586 27859 7607
rect 28073 7590 28144 8243
rect 28659 8177 28702 8890
rect 29319 8801 29414 8821
rect 29319 8757 29339 8801
rect 29399 8757 29414 8801
rect 29319 8461 29414 8757
rect 29319 8420 29352 8461
rect 29388 8420 29414 8461
rect 29514 8500 29576 8971
rect 30856 8911 30893 8912
rect 31159 8911 31196 9053
rect 31221 9073 31308 9080
rect 31221 9070 31279 9073
rect 31221 9050 31226 9070
rect 31247 9053 31279 9070
rect 31299 9053 31308 9073
rect 31247 9050 31308 9053
rect 31221 9043 31308 9050
rect 31367 9073 31404 9083
rect 31367 9053 31375 9073
rect 31395 9053 31404 9073
rect 31221 9042 31252 9043
rect 31367 8974 31404 9053
rect 31434 9082 31465 9135
rect 31678 9128 31693 9136
rect 31733 9128 31743 9165
rect 32934 9154 32999 9293
rect 33274 9238 33311 9317
rect 33352 9304 33462 9317
rect 33426 9248 33457 9249
rect 33274 9218 33283 9238
rect 33303 9218 33311 9238
rect 31678 9119 31743 9128
rect 31891 9126 31956 9147
rect 31891 9108 31916 9126
rect 31934 9108 31956 9126
rect 32934 9136 32957 9154
rect 32975 9136 32999 9154
rect 32934 9119 32999 9136
rect 33154 9200 33222 9213
rect 33274 9208 33311 9218
rect 33370 9238 33457 9248
rect 33370 9218 33379 9238
rect 33399 9218 33457 9238
rect 33370 9209 33457 9218
rect 33370 9208 33407 9209
rect 33154 9158 33161 9200
rect 33210 9158 33222 9200
rect 33154 9155 33222 9158
rect 33426 9156 33457 9209
rect 33487 9238 33524 9317
rect 33639 9248 33670 9249
rect 33487 9218 33496 9238
rect 33516 9218 33524 9238
rect 33487 9208 33524 9218
rect 33583 9241 33670 9248
rect 33583 9238 33644 9241
rect 33583 9218 33592 9238
rect 33612 9221 33644 9238
rect 33665 9221 33670 9241
rect 33612 9218 33670 9221
rect 33583 9211 33670 9218
rect 33695 9238 33732 9380
rect 33998 9379 34035 9380
rect 34743 9377 35159 9382
rect 34743 9376 35084 9377
rect 34400 9345 34510 9359
rect 34400 9342 34443 9345
rect 34400 9337 34404 9342
rect 34322 9315 34404 9337
rect 34433 9315 34443 9342
rect 34471 9318 34478 9345
rect 34507 9337 34510 9345
rect 34507 9318 34572 9337
rect 34471 9315 34572 9318
rect 34322 9313 34572 9315
rect 33847 9248 33883 9249
rect 33695 9218 33704 9238
rect 33724 9218 33732 9238
rect 33583 9209 33639 9211
rect 33583 9208 33620 9209
rect 33695 9208 33732 9218
rect 33791 9238 33939 9248
rect 34039 9245 34135 9247
rect 33791 9218 33800 9238
rect 33820 9218 33910 9238
rect 33930 9218 33939 9238
rect 33791 9212 33939 9218
rect 33791 9209 33855 9212
rect 33791 9208 33828 9209
rect 33847 9182 33855 9209
rect 33876 9209 33939 9212
rect 33997 9238 34135 9245
rect 33997 9218 34006 9238
rect 34026 9218 34135 9238
rect 33997 9209 34135 9218
rect 34322 9234 34359 9313
rect 34400 9300 34510 9313
rect 34474 9244 34505 9245
rect 34322 9214 34331 9234
rect 34351 9214 34359 9234
rect 33876 9182 33883 9209
rect 33902 9208 33939 9209
rect 33998 9208 34035 9209
rect 33847 9157 33883 9182
rect 33318 9155 33359 9156
rect 33154 9148 33359 9155
rect 33154 9137 33328 9148
rect 31484 9082 31521 9083
rect 31434 9073 31521 9082
rect 31434 9053 31492 9073
rect 31512 9053 31521 9073
rect 31434 9043 31521 9053
rect 31580 9073 31617 9083
rect 31580 9053 31588 9073
rect 31608 9053 31617 9073
rect 31434 9042 31465 9043
rect 31429 8974 31539 8987
rect 31580 8974 31617 9053
rect 31891 9032 31956 9108
rect 33154 9104 33162 9137
rect 33155 9095 33162 9104
rect 33211 9128 33328 9137
rect 33348 9128 33359 9148
rect 33211 9120 33359 9128
rect 33426 9152 33785 9156
rect 33426 9147 33748 9152
rect 33426 9123 33539 9147
rect 33563 9128 33748 9147
rect 33772 9128 33785 9152
rect 33563 9123 33785 9128
rect 33426 9120 33785 9123
rect 33847 9120 33882 9157
rect 33950 9154 34050 9157
rect 33950 9150 34017 9154
rect 33950 9124 33962 9150
rect 33988 9128 34017 9150
rect 34043 9128 34050 9154
rect 33988 9124 34050 9128
rect 33950 9120 34050 9124
rect 33211 9104 33222 9120
rect 33211 9095 33219 9104
rect 33426 9099 33457 9120
rect 33847 9099 33883 9120
rect 33269 9098 33306 9099
rect 32934 9055 32999 9074
rect 32934 9037 32959 9055
rect 32977 9037 32999 9055
rect 31367 8972 31617 8974
rect 31367 8969 31468 8972
rect 31367 8950 31432 8969
rect 31429 8942 31432 8950
rect 31461 8942 31468 8969
rect 31496 8945 31506 8972
rect 31535 8950 31617 8972
rect 31640 8997 31957 9032
rect 31535 8945 31539 8950
rect 31496 8942 31539 8945
rect 31429 8928 31539 8942
rect 30855 8910 31196 8911
rect 30780 8908 31196 8910
rect 31640 8908 31680 8997
rect 31891 8970 31956 8997
rect 31891 8952 31914 8970
rect 31932 8952 31956 8970
rect 31891 8932 31956 8952
rect 30777 8905 31680 8908
rect 30777 8885 30783 8905
rect 30803 8885 31680 8905
rect 30777 8881 31680 8885
rect 31640 8878 31680 8881
rect 31892 8871 31957 8892
rect 30110 8863 30771 8864
rect 30110 8856 31044 8863
rect 30110 8855 31016 8856
rect 30110 8835 30961 8855
rect 30993 8836 31016 8855
rect 31041 8836 31044 8856
rect 30993 8835 31044 8836
rect 30110 8828 31044 8835
rect 29709 8786 29877 8787
rect 30112 8786 30151 8828
rect 30940 8826 31044 8828
rect 31009 8824 31044 8826
rect 31892 8853 31916 8871
rect 31934 8853 31957 8871
rect 31892 8806 31957 8853
rect 29709 8760 30153 8786
rect 29709 8758 29877 8760
rect 29514 8481 29578 8500
rect 29514 8442 29531 8481
rect 29565 8442 29578 8481
rect 29514 8423 29578 8442
rect 29319 8394 29414 8420
rect 29709 8407 29736 8758
rect 30112 8754 30153 8760
rect 29776 8547 29840 8559
rect 30116 8555 30153 8754
rect 30615 8781 30687 8798
rect 30615 8742 30623 8781
rect 30668 8742 30687 8781
rect 30381 8644 30492 8659
rect 30381 8642 30423 8644
rect 30381 8622 30388 8642
rect 30407 8622 30423 8642
rect 30381 8614 30423 8622
rect 30451 8642 30492 8644
rect 30451 8622 30465 8642
rect 30484 8622 30492 8642
rect 30451 8614 30492 8622
rect 30381 8608 30492 8614
rect 30324 8586 30573 8608
rect 30324 8555 30361 8586
rect 30537 8584 30573 8586
rect 30537 8555 30574 8584
rect 29776 8546 29811 8547
rect 29753 8541 29811 8546
rect 29753 8521 29756 8541
rect 29776 8527 29811 8541
rect 29831 8527 29840 8547
rect 29776 8519 29840 8527
rect 29802 8518 29840 8519
rect 29803 8517 29840 8518
rect 29906 8551 29942 8552
rect 30014 8551 30050 8552
rect 29906 8543 30050 8551
rect 29906 8523 29914 8543
rect 29934 8523 30022 8543
rect 30042 8523 30050 8543
rect 29906 8517 30050 8523
rect 30116 8547 30154 8555
rect 30222 8551 30258 8552
rect 30116 8527 30125 8547
rect 30145 8527 30154 8547
rect 30116 8518 30154 8527
rect 30173 8544 30258 8551
rect 30173 8524 30180 8544
rect 30201 8543 30258 8544
rect 30201 8524 30230 8543
rect 30173 8523 30230 8524
rect 30250 8523 30258 8543
rect 30116 8517 30153 8518
rect 30173 8517 30258 8523
rect 30324 8547 30362 8555
rect 30435 8551 30471 8552
rect 30324 8527 30333 8547
rect 30353 8527 30362 8547
rect 30324 8518 30362 8527
rect 30386 8543 30471 8551
rect 30386 8523 30443 8543
rect 30463 8523 30471 8543
rect 30324 8517 30361 8518
rect 30386 8517 30471 8523
rect 30537 8547 30575 8555
rect 30537 8527 30546 8547
rect 30566 8527 30575 8547
rect 30537 8518 30575 8527
rect 30615 8532 30687 8742
rect 30757 8776 31957 8806
rect 30757 8775 31201 8776
rect 30757 8773 30925 8775
rect 30615 8518 30698 8532
rect 30537 8517 30574 8518
rect 29960 8496 29996 8517
rect 30386 8496 30417 8517
rect 30615 8496 30632 8518
rect 29793 8492 29893 8496
rect 29793 8488 29855 8492
rect 29793 8462 29800 8488
rect 29826 8466 29855 8488
rect 29881 8466 29893 8492
rect 29826 8462 29893 8466
rect 29793 8459 29893 8462
rect 29961 8459 29996 8496
rect 30058 8493 30417 8496
rect 30058 8488 30280 8493
rect 30058 8464 30071 8488
rect 30095 8469 30280 8488
rect 30304 8469 30417 8493
rect 30095 8464 30417 8469
rect 30058 8460 30417 8464
rect 30484 8488 30632 8496
rect 30484 8468 30495 8488
rect 30515 8485 30632 8488
rect 30685 8485 30698 8518
rect 30515 8468 30698 8485
rect 30484 8461 30698 8468
rect 30484 8460 30525 8461
rect 30615 8460 30698 8461
rect 29960 8434 29996 8459
rect 29808 8407 29845 8408
rect 29904 8407 29941 8408
rect 29960 8407 29967 8434
rect 29708 8398 29846 8407
rect 29708 8378 29817 8398
rect 29837 8378 29846 8398
rect 29708 8371 29846 8378
rect 29904 8404 29967 8407
rect 29988 8407 29996 8434
rect 30015 8407 30052 8408
rect 29988 8404 30052 8407
rect 29904 8398 30052 8404
rect 29904 8378 29913 8398
rect 29933 8378 30023 8398
rect 30043 8378 30052 8398
rect 29708 8369 29804 8371
rect 29904 8368 30052 8378
rect 30111 8398 30148 8408
rect 30223 8407 30260 8408
rect 30204 8405 30260 8407
rect 30111 8378 30119 8398
rect 30139 8378 30148 8398
rect 29960 8367 29996 8368
rect 29808 8236 29845 8237
rect 30111 8236 30148 8378
rect 30173 8398 30260 8405
rect 30173 8395 30231 8398
rect 30173 8375 30178 8395
rect 30199 8378 30231 8395
rect 30251 8378 30260 8398
rect 30199 8375 30260 8378
rect 30173 8368 30260 8375
rect 30319 8398 30356 8408
rect 30319 8378 30327 8398
rect 30347 8378 30356 8398
rect 30173 8367 30204 8368
rect 30319 8299 30356 8378
rect 30386 8407 30417 8460
rect 30623 8427 30637 8460
rect 30690 8427 30698 8460
rect 30623 8421 30698 8427
rect 30623 8416 30693 8421
rect 30436 8407 30473 8408
rect 30386 8398 30473 8407
rect 30386 8378 30444 8398
rect 30464 8378 30473 8398
rect 30386 8368 30473 8378
rect 30532 8398 30569 8408
rect 30757 8403 30784 8773
rect 30824 8543 30888 8555
rect 31164 8551 31201 8775
rect 31672 8756 31736 8758
rect 31668 8744 31736 8756
rect 31668 8711 31679 8744
rect 31719 8711 31736 8744
rect 31668 8701 31736 8711
rect 31429 8640 31540 8655
rect 31429 8638 31471 8640
rect 31429 8618 31436 8638
rect 31455 8618 31471 8638
rect 31429 8610 31471 8618
rect 31499 8638 31540 8640
rect 31499 8618 31513 8638
rect 31532 8618 31540 8638
rect 31499 8610 31540 8618
rect 31429 8604 31540 8610
rect 31372 8582 31621 8604
rect 31372 8551 31409 8582
rect 31585 8580 31621 8582
rect 31585 8551 31622 8580
rect 30824 8542 30859 8543
rect 30801 8537 30859 8542
rect 30801 8517 30804 8537
rect 30824 8523 30859 8537
rect 30879 8523 30888 8543
rect 30824 8515 30888 8523
rect 30850 8514 30888 8515
rect 30851 8513 30888 8514
rect 30954 8547 30990 8548
rect 31062 8547 31098 8548
rect 30954 8539 31098 8547
rect 30954 8519 30962 8539
rect 30982 8519 31070 8539
rect 31090 8519 31098 8539
rect 30954 8513 31098 8519
rect 31164 8543 31202 8551
rect 31270 8547 31306 8548
rect 31164 8523 31173 8543
rect 31193 8523 31202 8543
rect 31164 8514 31202 8523
rect 31221 8540 31306 8547
rect 31221 8520 31228 8540
rect 31249 8539 31306 8540
rect 31249 8520 31278 8539
rect 31221 8519 31278 8520
rect 31298 8519 31306 8539
rect 31164 8513 31201 8514
rect 31221 8513 31306 8519
rect 31372 8543 31410 8551
rect 31483 8547 31519 8548
rect 31372 8523 31381 8543
rect 31401 8523 31410 8543
rect 31372 8514 31410 8523
rect 31434 8539 31519 8547
rect 31434 8519 31491 8539
rect 31511 8519 31519 8539
rect 31372 8513 31409 8514
rect 31434 8513 31519 8519
rect 31585 8543 31623 8551
rect 31585 8523 31594 8543
rect 31614 8523 31623 8543
rect 31585 8514 31623 8523
rect 31672 8517 31736 8701
rect 31892 8575 31957 8776
rect 32934 8836 32999 9037
rect 33155 8911 33219 9095
rect 33268 9089 33306 9098
rect 33268 9069 33277 9089
rect 33297 9069 33306 9089
rect 33268 9061 33306 9069
rect 33372 9093 33457 9099
rect 33482 9098 33519 9099
rect 33372 9073 33380 9093
rect 33400 9073 33457 9093
rect 33372 9065 33457 9073
rect 33481 9089 33519 9098
rect 33481 9069 33490 9089
rect 33510 9069 33519 9089
rect 33372 9064 33408 9065
rect 33481 9061 33519 9069
rect 33585 9093 33670 9099
rect 33690 9098 33727 9099
rect 33585 9073 33593 9093
rect 33613 9092 33670 9093
rect 33613 9073 33642 9092
rect 33585 9072 33642 9073
rect 33663 9072 33670 9092
rect 33585 9065 33670 9072
rect 33689 9089 33727 9098
rect 33689 9069 33698 9089
rect 33718 9069 33727 9089
rect 33585 9064 33621 9065
rect 33689 9061 33727 9069
rect 33793 9093 33937 9099
rect 33793 9073 33801 9093
rect 33821 9073 33909 9093
rect 33929 9073 33937 9093
rect 33793 9065 33937 9073
rect 33793 9064 33829 9065
rect 33901 9064 33937 9065
rect 34003 9098 34040 9099
rect 34003 9097 34041 9098
rect 34003 9089 34067 9097
rect 34003 9069 34012 9089
rect 34032 9075 34067 9089
rect 34087 9075 34090 9095
rect 34032 9070 34090 9075
rect 34032 9069 34067 9070
rect 33269 9032 33306 9061
rect 33270 9030 33306 9032
rect 33482 9030 33519 9061
rect 33270 9008 33519 9030
rect 33351 9002 33462 9008
rect 33351 8994 33392 9002
rect 33351 8974 33359 8994
rect 33378 8974 33392 8994
rect 33351 8972 33392 8974
rect 33420 8994 33462 9002
rect 33420 8974 33436 8994
rect 33455 8974 33462 8994
rect 33420 8972 33462 8974
rect 33351 8957 33462 8972
rect 33155 8901 33223 8911
rect 33155 8868 33172 8901
rect 33212 8868 33223 8901
rect 33155 8856 33223 8868
rect 33155 8854 33219 8856
rect 33690 8837 33727 9061
rect 34003 9057 34067 9069
rect 34107 8839 34134 9209
rect 34322 9204 34359 9214
rect 34418 9234 34505 9244
rect 34418 9214 34427 9234
rect 34447 9214 34505 9234
rect 34418 9205 34505 9214
rect 34418 9204 34455 9205
rect 34198 9191 34268 9196
rect 34193 9185 34268 9191
rect 34193 9152 34201 9185
rect 34254 9152 34268 9185
rect 34474 9152 34505 9205
rect 34535 9234 34572 9313
rect 34687 9244 34718 9245
rect 34535 9214 34544 9234
rect 34564 9214 34572 9234
rect 34535 9204 34572 9214
rect 34631 9237 34718 9244
rect 34631 9234 34692 9237
rect 34631 9214 34640 9234
rect 34660 9217 34692 9234
rect 34713 9217 34718 9237
rect 34660 9214 34718 9217
rect 34631 9207 34718 9214
rect 34743 9234 34780 9376
rect 35046 9375 35083 9376
rect 34895 9244 34931 9245
rect 34743 9214 34752 9234
rect 34772 9214 34780 9234
rect 34631 9205 34687 9207
rect 34631 9204 34668 9205
rect 34743 9204 34780 9214
rect 34839 9234 34987 9244
rect 35087 9241 35183 9243
rect 34839 9214 34848 9234
rect 34868 9214 34958 9234
rect 34978 9214 34987 9234
rect 34839 9208 34987 9214
rect 34839 9205 34903 9208
rect 34839 9204 34876 9205
rect 34895 9178 34903 9205
rect 34924 9205 34987 9208
rect 35045 9234 35183 9241
rect 35045 9214 35054 9234
rect 35074 9214 35183 9234
rect 35045 9205 35183 9214
rect 34924 9178 34931 9205
rect 34950 9204 34987 9205
rect 35046 9204 35083 9205
rect 34895 9153 34931 9178
rect 34193 9151 34276 9152
rect 34366 9151 34407 9152
rect 34193 9144 34407 9151
rect 34193 9127 34376 9144
rect 34193 9094 34206 9127
rect 34259 9124 34376 9127
rect 34396 9124 34407 9144
rect 34259 9116 34407 9124
rect 34474 9148 34833 9152
rect 34474 9143 34796 9148
rect 34474 9119 34587 9143
rect 34611 9124 34796 9143
rect 34820 9124 34833 9148
rect 34611 9119 34833 9124
rect 34474 9116 34833 9119
rect 34895 9116 34930 9153
rect 34998 9150 35098 9153
rect 34998 9146 35065 9150
rect 34998 9120 35010 9146
rect 35036 9124 35065 9146
rect 35091 9124 35098 9150
rect 35036 9120 35098 9124
rect 34998 9116 35098 9120
rect 34259 9094 34276 9116
rect 34474 9095 34505 9116
rect 34895 9095 34931 9116
rect 34317 9094 34354 9095
rect 34193 9080 34276 9094
rect 33966 8837 34134 8839
rect 33690 8836 34134 8837
rect 32934 8806 34134 8836
rect 34204 8870 34276 9080
rect 34316 9085 34354 9094
rect 34316 9065 34325 9085
rect 34345 9065 34354 9085
rect 34316 9057 34354 9065
rect 34420 9089 34505 9095
rect 34530 9094 34567 9095
rect 34420 9069 34428 9089
rect 34448 9069 34505 9089
rect 34420 9061 34505 9069
rect 34529 9085 34567 9094
rect 34529 9065 34538 9085
rect 34558 9065 34567 9085
rect 34420 9060 34456 9061
rect 34529 9057 34567 9065
rect 34633 9089 34718 9095
rect 34738 9094 34775 9095
rect 34633 9069 34641 9089
rect 34661 9088 34718 9089
rect 34661 9069 34690 9088
rect 34633 9068 34690 9069
rect 34711 9068 34718 9088
rect 34633 9061 34718 9068
rect 34737 9085 34775 9094
rect 34737 9065 34746 9085
rect 34766 9065 34775 9085
rect 34633 9060 34669 9061
rect 34737 9057 34775 9065
rect 34841 9089 34985 9095
rect 34841 9069 34849 9089
rect 34869 9069 34957 9089
rect 34977 9069 34985 9089
rect 34841 9061 34985 9069
rect 34841 9060 34877 9061
rect 34949 9060 34985 9061
rect 35051 9094 35088 9095
rect 35051 9093 35089 9094
rect 35051 9085 35115 9093
rect 35051 9065 35060 9085
rect 35080 9071 35115 9085
rect 35135 9071 35138 9091
rect 35080 9066 35138 9071
rect 35080 9065 35115 9066
rect 34317 9028 34354 9057
rect 34318 9026 34354 9028
rect 34530 9026 34567 9057
rect 34318 9004 34567 9026
rect 34399 8998 34510 9004
rect 34399 8990 34440 8998
rect 34399 8970 34407 8990
rect 34426 8970 34440 8990
rect 34399 8968 34440 8970
rect 34468 8990 34510 8998
rect 34468 8970 34484 8990
rect 34503 8970 34510 8990
rect 34468 8968 34510 8970
rect 34399 8953 34510 8968
rect 34204 8831 34223 8870
rect 34268 8831 34276 8870
rect 34204 8814 34276 8831
rect 34738 8858 34775 9057
rect 35051 9053 35115 9065
rect 34738 8852 34779 8858
rect 35155 8854 35182 9205
rect 35014 8852 35182 8854
rect 34738 8826 35182 8852
rect 32934 8759 32999 8806
rect 32934 8741 32957 8759
rect 32975 8741 32999 8759
rect 33847 8786 33882 8788
rect 33847 8784 33951 8786
rect 34740 8784 34779 8826
rect 35014 8825 35182 8826
rect 33847 8777 34781 8784
rect 33847 8776 33898 8777
rect 33847 8756 33850 8776
rect 33875 8757 33898 8776
rect 33930 8757 34781 8777
rect 33875 8756 34781 8757
rect 33847 8749 34781 8756
rect 34120 8748 34781 8749
rect 32934 8720 32999 8741
rect 33211 8731 33251 8734
rect 33211 8727 34114 8731
rect 33211 8707 34088 8727
rect 34108 8707 34114 8727
rect 33211 8704 34114 8707
rect 32935 8660 33000 8680
rect 32935 8642 32959 8660
rect 32977 8642 33000 8660
rect 32935 8615 33000 8642
rect 33211 8615 33251 8704
rect 33695 8702 34111 8704
rect 33695 8701 34036 8702
rect 33352 8670 33462 8684
rect 33352 8667 33395 8670
rect 33352 8662 33356 8667
rect 32934 8580 33251 8615
rect 33274 8640 33356 8662
rect 33385 8640 33395 8667
rect 33423 8643 33430 8670
rect 33459 8662 33462 8670
rect 33459 8643 33524 8662
rect 33423 8640 33524 8643
rect 33274 8638 33524 8640
rect 31892 8557 31914 8575
rect 31932 8557 31957 8575
rect 31892 8538 31957 8557
rect 31585 8513 31622 8514
rect 31008 8492 31044 8513
rect 31434 8492 31465 8513
rect 31672 8508 31680 8517
rect 31669 8492 31680 8508
rect 30841 8488 30941 8492
rect 30841 8484 30903 8488
rect 30841 8458 30848 8484
rect 30874 8462 30903 8484
rect 30929 8462 30941 8488
rect 30874 8458 30941 8462
rect 30841 8455 30941 8458
rect 31009 8455 31044 8492
rect 31106 8489 31465 8492
rect 31106 8484 31328 8489
rect 31106 8460 31119 8484
rect 31143 8465 31328 8484
rect 31352 8465 31465 8489
rect 31143 8460 31465 8465
rect 31106 8456 31465 8460
rect 31532 8484 31680 8492
rect 31532 8464 31543 8484
rect 31563 8475 31680 8484
rect 31729 8508 31736 8517
rect 31729 8475 31737 8508
rect 32935 8504 33000 8580
rect 33274 8559 33311 8638
rect 33352 8625 33462 8638
rect 33426 8569 33457 8570
rect 33274 8539 33283 8559
rect 33303 8539 33311 8559
rect 33274 8529 33311 8539
rect 33370 8559 33457 8569
rect 33370 8539 33379 8559
rect 33399 8539 33457 8559
rect 33370 8530 33457 8539
rect 33370 8529 33407 8530
rect 31563 8464 31737 8475
rect 31532 8457 31737 8464
rect 31532 8456 31573 8457
rect 31008 8430 31044 8455
rect 30856 8403 30893 8404
rect 30952 8403 30989 8404
rect 31008 8403 31015 8430
rect 30532 8378 30540 8398
rect 30560 8378 30569 8398
rect 30386 8367 30417 8368
rect 30381 8299 30491 8312
rect 30532 8299 30569 8378
rect 30756 8394 30894 8403
rect 30756 8374 30865 8394
rect 30885 8374 30894 8394
rect 30756 8367 30894 8374
rect 30952 8400 31015 8403
rect 31036 8403 31044 8430
rect 31063 8403 31100 8404
rect 31036 8400 31100 8403
rect 30952 8394 31100 8400
rect 30952 8374 30961 8394
rect 30981 8374 31071 8394
rect 31091 8374 31100 8394
rect 30756 8365 30852 8367
rect 30952 8364 31100 8374
rect 31159 8394 31196 8404
rect 31271 8403 31308 8404
rect 31252 8401 31308 8403
rect 31159 8374 31167 8394
rect 31187 8374 31196 8394
rect 31008 8363 31044 8364
rect 30319 8297 30569 8299
rect 30319 8294 30420 8297
rect 30319 8275 30384 8294
rect 30381 8267 30384 8275
rect 30413 8267 30420 8294
rect 30448 8270 30458 8297
rect 30487 8275 30569 8297
rect 30487 8270 30491 8275
rect 30448 8267 30491 8270
rect 30381 8253 30491 8267
rect 29807 8235 30148 8236
rect 29732 8230 30148 8235
rect 30856 8232 30893 8233
rect 31159 8232 31196 8374
rect 31221 8394 31308 8401
rect 31221 8391 31279 8394
rect 31221 8371 31226 8391
rect 31247 8374 31279 8391
rect 31299 8374 31308 8394
rect 31247 8371 31308 8374
rect 31221 8364 31308 8371
rect 31367 8394 31404 8404
rect 31367 8374 31375 8394
rect 31395 8374 31404 8394
rect 31221 8363 31252 8364
rect 31367 8295 31404 8374
rect 31434 8403 31465 8456
rect 31669 8454 31737 8457
rect 31669 8412 31681 8454
rect 31730 8412 31737 8454
rect 31484 8403 31521 8404
rect 31434 8394 31521 8403
rect 31434 8374 31492 8394
rect 31512 8374 31521 8394
rect 31434 8364 31521 8374
rect 31580 8394 31617 8404
rect 31669 8399 31737 8412
rect 31892 8476 31957 8493
rect 31892 8458 31916 8476
rect 31934 8458 31957 8476
rect 32935 8486 32957 8504
rect 32975 8486 33000 8504
rect 32935 8465 33000 8486
rect 33148 8484 33213 8493
rect 31580 8374 31588 8394
rect 31608 8374 31617 8394
rect 31434 8363 31465 8364
rect 31429 8295 31539 8308
rect 31580 8295 31617 8374
rect 31892 8319 31957 8458
rect 33148 8447 33158 8484
rect 33198 8476 33213 8484
rect 33426 8477 33457 8530
rect 33487 8559 33524 8638
rect 33639 8569 33670 8570
rect 33487 8539 33496 8559
rect 33516 8539 33524 8559
rect 33487 8529 33524 8539
rect 33583 8562 33670 8569
rect 33583 8559 33644 8562
rect 33583 8539 33592 8559
rect 33612 8542 33644 8559
rect 33665 8542 33670 8562
rect 33612 8539 33670 8542
rect 33583 8532 33670 8539
rect 33695 8559 33732 8701
rect 33998 8700 34035 8701
rect 33847 8569 33883 8570
rect 33695 8539 33704 8559
rect 33724 8539 33732 8559
rect 33583 8530 33639 8532
rect 33583 8529 33620 8530
rect 33695 8529 33732 8539
rect 33791 8559 33939 8569
rect 34039 8566 34135 8568
rect 33791 8539 33800 8559
rect 33820 8539 33910 8559
rect 33930 8539 33939 8559
rect 33791 8533 33939 8539
rect 33791 8530 33855 8533
rect 33791 8529 33828 8530
rect 33847 8503 33855 8530
rect 33876 8530 33939 8533
rect 33997 8559 34135 8566
rect 33997 8539 34006 8559
rect 34026 8539 34135 8559
rect 33997 8530 34135 8539
rect 33876 8503 33883 8530
rect 33902 8529 33939 8530
rect 33998 8529 34035 8530
rect 33847 8478 33883 8503
rect 33318 8476 33359 8477
rect 33198 8469 33359 8476
rect 33198 8449 33328 8469
rect 33348 8449 33359 8469
rect 33198 8447 33359 8449
rect 33148 8441 33359 8447
rect 33426 8473 33785 8477
rect 33426 8468 33748 8473
rect 33426 8444 33539 8468
rect 33563 8449 33748 8468
rect 33772 8449 33785 8473
rect 33563 8444 33785 8449
rect 33426 8441 33785 8444
rect 33847 8441 33882 8478
rect 33950 8475 34050 8478
rect 33950 8471 34017 8475
rect 33950 8445 33962 8471
rect 33988 8449 34017 8471
rect 34043 8449 34050 8475
rect 33988 8445 34050 8449
rect 33950 8441 34050 8445
rect 33148 8428 33215 8441
rect 31892 8313 31914 8319
rect 31367 8293 31617 8295
rect 31367 8290 31468 8293
rect 31367 8271 31432 8290
rect 31429 8263 31432 8271
rect 31461 8263 31468 8290
rect 31496 8266 31506 8293
rect 31535 8271 31617 8293
rect 31646 8301 31914 8313
rect 31932 8301 31957 8319
rect 31646 8278 31957 8301
rect 32940 8405 32996 8425
rect 32940 8387 32959 8405
rect 32977 8387 32996 8405
rect 31646 8277 31701 8278
rect 31535 8266 31539 8271
rect 31496 8263 31539 8266
rect 31429 8249 31539 8263
rect 30855 8231 31196 8232
rect 29732 8210 29735 8230
rect 29755 8210 30148 8230
rect 30780 8230 31196 8231
rect 31646 8230 31689 8277
rect 32940 8274 32996 8387
rect 33148 8407 33162 8428
rect 33198 8407 33215 8428
rect 33426 8420 33457 8441
rect 33847 8420 33883 8441
rect 33269 8419 33306 8420
rect 33148 8400 33215 8407
rect 33268 8410 33306 8419
rect 30780 8226 31689 8230
rect 28655 8175 29366 8177
rect 29905 8175 29994 8178
rect 28655 8166 29994 8175
rect 28655 8128 29917 8166
rect 29942 8131 29961 8166
rect 29986 8131 29994 8166
rect 30099 8177 30144 8210
rect 30780 8206 30783 8226
rect 30803 8206 31689 8226
rect 31157 8201 31689 8206
rect 31897 8220 31956 8242
rect 31897 8202 31916 8220
rect 31934 8202 31956 8220
rect 30945 8177 31044 8179
rect 30099 8167 31044 8177
rect 30099 8141 30967 8167
rect 30100 8140 30967 8141
rect 29942 8128 29994 8131
rect 28655 8120 29994 8128
rect 30945 8129 30967 8140
rect 30992 8132 31011 8167
rect 31036 8132 31044 8167
rect 30992 8129 31044 8132
rect 30945 8121 31044 8129
rect 31897 8128 31956 8202
rect 32940 8167 32995 8274
rect 33148 8248 33213 8400
rect 33268 8390 33277 8410
rect 33297 8390 33306 8410
rect 33268 8382 33306 8390
rect 33372 8414 33457 8420
rect 33482 8419 33519 8420
rect 33372 8394 33380 8414
rect 33400 8394 33457 8414
rect 33372 8386 33457 8394
rect 33481 8410 33519 8419
rect 33481 8390 33490 8410
rect 33510 8390 33519 8410
rect 33372 8385 33408 8386
rect 33481 8382 33519 8390
rect 33585 8414 33670 8420
rect 33690 8419 33727 8420
rect 33585 8394 33593 8414
rect 33613 8413 33670 8414
rect 33613 8394 33642 8413
rect 33585 8393 33642 8394
rect 33663 8393 33670 8413
rect 33585 8386 33670 8393
rect 33689 8410 33727 8419
rect 33689 8390 33698 8410
rect 33718 8390 33727 8410
rect 33585 8385 33621 8386
rect 33689 8382 33727 8390
rect 33793 8414 33937 8420
rect 33793 8394 33801 8414
rect 33821 8394 33909 8414
rect 33929 8394 33937 8414
rect 33793 8386 33937 8394
rect 33793 8385 33829 8386
rect 33901 8385 33937 8386
rect 34003 8419 34040 8420
rect 34003 8418 34041 8419
rect 34003 8410 34067 8418
rect 34003 8390 34012 8410
rect 34032 8396 34067 8410
rect 34087 8396 34090 8416
rect 34032 8391 34090 8396
rect 34032 8390 34067 8391
rect 33269 8353 33306 8382
rect 33270 8351 33306 8353
rect 33482 8351 33519 8382
rect 33270 8329 33519 8351
rect 33351 8323 33462 8329
rect 33351 8315 33392 8323
rect 33351 8295 33359 8315
rect 33378 8295 33392 8315
rect 33351 8293 33392 8295
rect 33420 8315 33462 8323
rect 33420 8295 33436 8315
rect 33455 8295 33462 8315
rect 33420 8293 33462 8295
rect 33351 8278 33462 8293
rect 33690 8283 33727 8382
rect 34003 8378 34067 8390
rect 33353 8275 33457 8278
rect 33141 8238 33262 8248
rect 33141 8236 33210 8238
rect 33141 8195 33154 8236
rect 33191 8197 33210 8236
rect 33247 8197 33262 8238
rect 33191 8195 33262 8197
rect 33141 8177 33262 8195
rect 30971 8120 31043 8121
rect 28655 8119 29993 8120
rect 28655 8117 29366 8119
rect 29515 8078 29579 8082
rect 31890 8080 31956 8128
rect 32933 8133 32998 8167
rect 33353 8133 33457 8135
rect 33688 8133 33729 8283
rect 34107 8275 34134 8530
rect 34196 8520 34276 8531
rect 34196 8494 34213 8520
rect 34253 8494 34276 8520
rect 34196 8467 34276 8494
rect 34196 8441 34217 8467
rect 34257 8441 34276 8467
rect 34196 8422 34276 8441
rect 34196 8396 34220 8422
rect 34260 8396 34276 8422
rect 34196 8345 34276 8396
rect 32933 8130 33729 8133
rect 34108 8144 34134 8275
rect 34198 8145 34268 8345
rect 34108 8130 34136 8144
rect 32933 8095 34136 8130
rect 34197 8123 34269 8145
rect 29515 8069 29589 8078
rect 28030 7586 28144 7590
rect 27235 7582 27335 7586
rect 27235 7578 27297 7582
rect 27235 7552 27242 7578
rect 27268 7556 27297 7578
rect 27323 7556 27335 7582
rect 27268 7552 27335 7556
rect 27235 7549 27335 7552
rect 27403 7549 27438 7586
rect 27500 7583 27859 7586
rect 27500 7578 27722 7583
rect 27500 7554 27513 7578
rect 27537 7559 27722 7578
rect 27746 7559 27859 7583
rect 27537 7554 27859 7559
rect 27500 7550 27859 7554
rect 27926 7583 28144 7586
rect 27926 7582 28109 7583
rect 27926 7578 28052 7582
rect 27926 7558 27937 7578
rect 27957 7558 28052 7578
rect 28076 7559 28109 7582
rect 28133 7559 28144 7583
rect 28076 7558 28144 7559
rect 27926 7551 28144 7558
rect 27926 7550 27967 7551
rect 27402 7524 27438 7549
rect 27250 7497 27287 7498
rect 27346 7497 27383 7498
rect 27402 7497 27409 7524
rect 27150 7488 27288 7497
rect 27150 7468 27259 7488
rect 27279 7468 27288 7488
rect 27150 7461 27288 7468
rect 27346 7494 27409 7497
rect 27430 7497 27438 7524
rect 27457 7497 27494 7498
rect 27430 7494 27494 7497
rect 27346 7488 27494 7494
rect 27346 7468 27355 7488
rect 27375 7468 27465 7488
rect 27485 7468 27494 7488
rect 27150 7459 27246 7461
rect 27346 7458 27494 7468
rect 27553 7488 27590 7498
rect 27665 7497 27702 7498
rect 27646 7495 27702 7497
rect 27553 7468 27561 7488
rect 27581 7468 27590 7488
rect 27402 7457 27438 7458
rect 27250 7326 27287 7327
rect 27553 7326 27590 7468
rect 27615 7488 27702 7495
rect 27615 7485 27673 7488
rect 27615 7465 27620 7485
rect 27641 7468 27673 7485
rect 27693 7468 27702 7488
rect 27641 7465 27702 7468
rect 27615 7458 27702 7465
rect 27761 7488 27798 7498
rect 27761 7468 27769 7488
rect 27789 7468 27798 7488
rect 27615 7457 27646 7458
rect 27761 7389 27798 7468
rect 27828 7497 27859 7550
rect 28030 7548 28144 7551
rect 28073 7516 28144 7548
rect 29319 8027 29403 8052
rect 29319 7999 29334 8027
rect 29378 7999 29403 8027
rect 29319 7970 29403 7999
rect 29515 8021 29529 8069
rect 29566 8021 29589 8069
rect 29515 7993 29589 8021
rect 29319 7942 29331 7970
rect 29375 7942 29403 7970
rect 29319 7921 29403 7942
rect 27878 7497 27915 7498
rect 27828 7488 27915 7497
rect 27828 7468 27886 7488
rect 27906 7468 27915 7488
rect 27828 7458 27915 7468
rect 27974 7488 28011 7498
rect 27974 7468 27982 7488
rect 28002 7468 28011 7488
rect 27828 7457 27859 7458
rect 27823 7389 27933 7402
rect 27974 7389 28011 7468
rect 27761 7387 28011 7389
rect 27761 7384 27862 7387
rect 27761 7365 27826 7384
rect 27823 7357 27826 7365
rect 27855 7357 27862 7384
rect 27890 7360 27900 7387
rect 27929 7365 28011 7387
rect 27929 7360 27933 7365
rect 27890 7357 27933 7360
rect 27823 7343 27933 7357
rect 27249 7325 27590 7326
rect 27174 7322 27590 7325
rect 27174 7320 27597 7322
rect 27174 7300 27177 7320
rect 27197 7300 27597 7320
rect 26365 4959 27005 5047
rect 26365 4608 26449 4959
rect 26931 4928 26975 4934
rect 26931 4902 26939 4928
rect 26964 4902 26975 4928
rect 26931 4853 26975 4902
rect 26931 4833 27328 4853
rect 27348 4833 27351 4853
rect 26931 4828 27351 4833
rect 26931 4827 27276 4828
rect 26931 4823 26975 4827
rect 27238 4826 27275 4827
rect 26592 4796 26702 4810
rect 26592 4793 26635 4796
rect 26592 4788 26596 4793
rect 26514 4766 26596 4788
rect 26625 4766 26635 4793
rect 26663 4769 26670 4796
rect 26699 4788 26702 4796
rect 26699 4769 26764 4788
rect 26663 4766 26764 4769
rect 26514 4764 26764 4766
rect 26514 4685 26551 4764
rect 26592 4751 26702 4764
rect 26666 4695 26697 4696
rect 26514 4665 26523 4685
rect 26543 4665 26551 4685
rect 26514 4655 26551 4665
rect 26610 4685 26697 4695
rect 26610 4665 26619 4685
rect 26639 4665 26697 4685
rect 26610 4656 26697 4665
rect 26610 4655 26647 4656
rect 26365 4602 26474 4608
rect 26666 4603 26697 4656
rect 26727 4685 26764 4764
rect 26879 4695 26910 4696
rect 26727 4665 26736 4685
rect 26756 4665 26764 4685
rect 26727 4655 26764 4665
rect 26823 4688 26910 4695
rect 26823 4685 26884 4688
rect 26823 4665 26832 4685
rect 26852 4668 26884 4685
rect 26905 4668 26910 4688
rect 26852 4665 26910 4668
rect 26823 4658 26910 4665
rect 26935 4685 26972 4823
rect 27087 4695 27123 4696
rect 26935 4665 26944 4685
rect 26964 4665 26972 4685
rect 26823 4656 26879 4658
rect 26823 4655 26860 4656
rect 26935 4655 26972 4665
rect 27031 4685 27179 4695
rect 27279 4692 27375 4694
rect 27031 4665 27040 4685
rect 27060 4665 27150 4685
rect 27170 4665 27179 4685
rect 27031 4659 27179 4665
rect 27031 4656 27095 4659
rect 27031 4655 27068 4656
rect 27087 4629 27095 4656
rect 27116 4656 27179 4659
rect 27237 4685 27375 4692
rect 27237 4665 27246 4685
rect 27266 4665 27375 4685
rect 27237 4656 27375 4665
rect 27116 4629 27123 4656
rect 27142 4655 27179 4656
rect 27238 4655 27275 4656
rect 27087 4604 27123 4629
rect 26558 4602 26599 4603
rect 26365 4595 26599 4602
rect 26365 4575 26568 4595
rect 26588 4575 26599 4595
rect 26365 4567 26599 4575
rect 26666 4599 27025 4603
rect 26666 4594 26988 4599
rect 26666 4570 26779 4594
rect 26803 4575 26988 4594
rect 27012 4575 27025 4599
rect 26803 4570 27025 4575
rect 26666 4567 27025 4570
rect 27087 4567 27122 4604
rect 27190 4601 27290 4604
rect 27190 4597 27257 4601
rect 27190 4571 27202 4597
rect 27228 4575 27257 4597
rect 27283 4575 27290 4601
rect 27228 4571 27290 4575
rect 27190 4567 27290 4571
rect 26365 4549 26474 4567
rect 26666 4546 26697 4567
rect 27087 4546 27123 4567
rect 26509 4545 26546 4546
rect 26508 4536 26546 4545
rect 26508 4516 26517 4536
rect 26537 4516 26546 4536
rect 26508 4508 26546 4516
rect 26612 4540 26697 4546
rect 26722 4545 26759 4546
rect 26612 4520 26620 4540
rect 26640 4520 26697 4540
rect 26612 4512 26697 4520
rect 26721 4536 26759 4545
rect 26721 4516 26730 4536
rect 26750 4516 26759 4536
rect 26612 4511 26648 4512
rect 26721 4508 26759 4516
rect 26825 4540 26910 4546
rect 26930 4545 26967 4546
rect 26825 4520 26833 4540
rect 26853 4539 26910 4540
rect 26853 4520 26882 4539
rect 26825 4519 26882 4520
rect 26903 4519 26910 4539
rect 26825 4512 26910 4519
rect 26929 4536 26967 4545
rect 26929 4516 26938 4536
rect 26958 4516 26967 4536
rect 26825 4511 26861 4512
rect 26929 4508 26967 4516
rect 27033 4541 27177 4546
rect 27033 4540 27086 4541
rect 27033 4520 27041 4540
rect 27061 4521 27086 4540
rect 27119 4540 27177 4541
rect 27119 4521 27149 4540
rect 27061 4520 27149 4521
rect 27169 4520 27177 4540
rect 27033 4512 27177 4520
rect 27033 4511 27069 4512
rect 27141 4511 27177 4512
rect 27243 4545 27280 4546
rect 27243 4544 27281 4545
rect 27243 4536 27307 4544
rect 27243 4516 27252 4536
rect 27272 4522 27307 4536
rect 27327 4522 27330 4542
rect 27272 4517 27330 4522
rect 27272 4516 27307 4517
rect 26509 4479 26546 4508
rect 26510 4477 26546 4479
rect 26722 4477 26759 4508
rect 26510 4455 26759 4477
rect 26591 4449 26702 4455
rect 26591 4441 26632 4449
rect 26591 4421 26599 4441
rect 26618 4421 26632 4441
rect 26591 4419 26632 4421
rect 26660 4441 26702 4449
rect 26660 4421 26676 4441
rect 26695 4421 26702 4441
rect 26660 4419 26702 4421
rect 26591 4404 26702 4419
rect 26930 4387 26967 4508
rect 27243 4504 27307 4516
rect 27347 4393 27374 4656
rect 27401 4402 27437 4409
rect 27401 4393 27407 4402
rect 27325 4389 27407 4393
rect 27206 4387 27407 4389
rect 26930 4364 27407 4387
rect 27430 4364 27437 4402
rect 26930 4361 27437 4364
rect 27206 4360 27374 4361
rect 27401 4358 27437 4361
rect 27519 4260 27597 7300
rect 28653 6553 28712 6563
rect 28653 6525 28666 6553
rect 28694 6525 28712 6553
rect 28653 6476 28712 6525
rect 28259 6341 28427 6342
rect 28663 6341 28710 6476
rect 28259 6315 28710 6341
rect 28259 6313 28427 6315
rect 28259 6046 28286 6313
rect 28663 6309 28710 6315
rect 28326 6186 28390 6198
rect 28666 6194 28703 6309
rect 28931 6283 29042 6298
rect 28931 6281 28973 6283
rect 28931 6261 28938 6281
rect 28957 6261 28973 6281
rect 28931 6253 28973 6261
rect 29001 6281 29042 6283
rect 29001 6261 29015 6281
rect 29034 6261 29042 6281
rect 29001 6253 29042 6261
rect 28931 6247 29042 6253
rect 28874 6225 29123 6247
rect 28874 6194 28911 6225
rect 29087 6223 29123 6225
rect 29087 6194 29124 6223
rect 28326 6185 28361 6186
rect 28303 6180 28361 6185
rect 28303 6160 28306 6180
rect 28326 6166 28361 6180
rect 28381 6166 28390 6186
rect 28326 6158 28390 6166
rect 28352 6157 28390 6158
rect 28353 6156 28390 6157
rect 28456 6190 28492 6191
rect 28564 6190 28600 6191
rect 28456 6182 28600 6190
rect 28456 6162 28464 6182
rect 28484 6162 28572 6182
rect 28592 6162 28600 6182
rect 28456 6156 28600 6162
rect 28666 6186 28704 6194
rect 28772 6190 28808 6191
rect 28666 6166 28675 6186
rect 28695 6166 28704 6186
rect 28666 6157 28704 6166
rect 28723 6183 28808 6190
rect 28723 6163 28730 6183
rect 28751 6182 28808 6183
rect 28751 6163 28780 6182
rect 28723 6162 28780 6163
rect 28800 6162 28808 6182
rect 28666 6156 28703 6157
rect 28723 6156 28808 6162
rect 28874 6186 28912 6194
rect 28985 6190 29021 6191
rect 28874 6166 28883 6186
rect 28903 6166 28912 6186
rect 28874 6157 28912 6166
rect 28936 6182 29021 6190
rect 28936 6162 28993 6182
rect 29013 6162 29021 6182
rect 28874 6156 28911 6157
rect 28936 6156 29021 6162
rect 29087 6186 29125 6194
rect 29087 6166 29096 6186
rect 29116 6166 29125 6186
rect 29087 6157 29125 6166
rect 29087 6156 29124 6157
rect 28510 6135 28546 6156
rect 28936 6135 28967 6156
rect 29147 6141 29204 6149
rect 29147 6135 29155 6141
rect 28343 6131 28443 6135
rect 28343 6127 28405 6131
rect 28343 6101 28350 6127
rect 28376 6105 28405 6127
rect 28431 6105 28443 6131
rect 28376 6101 28443 6105
rect 28343 6098 28443 6101
rect 28511 6098 28546 6135
rect 28608 6132 28967 6135
rect 28608 6127 28830 6132
rect 28608 6103 28621 6127
rect 28645 6108 28830 6127
rect 28854 6108 28967 6132
rect 28645 6103 28967 6108
rect 28608 6099 28967 6103
rect 29034 6127 29155 6135
rect 29034 6107 29045 6127
rect 29065 6118 29155 6127
rect 29181 6118 29204 6141
rect 29065 6107 29204 6118
rect 29034 6105 29204 6107
rect 29034 6100 29155 6105
rect 29034 6099 29075 6100
rect 28510 6073 28546 6098
rect 28358 6046 28395 6047
rect 28454 6046 28491 6047
rect 28510 6046 28517 6073
rect 28258 6037 28396 6046
rect 28258 6017 28367 6037
rect 28387 6017 28396 6037
rect 28258 6010 28396 6017
rect 28454 6043 28517 6046
rect 28538 6046 28546 6073
rect 28565 6046 28602 6047
rect 28538 6043 28602 6046
rect 28454 6037 28602 6043
rect 28454 6017 28463 6037
rect 28483 6017 28573 6037
rect 28593 6017 28602 6037
rect 28258 6008 28354 6010
rect 28454 6007 28602 6017
rect 28661 6037 28698 6047
rect 28773 6046 28810 6047
rect 28754 6044 28810 6046
rect 28661 6017 28669 6037
rect 28689 6017 28698 6037
rect 28510 6006 28546 6007
rect 28358 5875 28395 5876
rect 28661 5875 28698 6017
rect 28723 6037 28810 6044
rect 28723 6034 28781 6037
rect 28723 6014 28728 6034
rect 28749 6017 28781 6034
rect 28801 6017 28810 6037
rect 28749 6014 28810 6017
rect 28723 6007 28810 6014
rect 28869 6037 28906 6047
rect 28869 6017 28877 6037
rect 28897 6017 28906 6037
rect 28723 6006 28754 6007
rect 28869 5938 28906 6017
rect 28936 6046 28967 6099
rect 28986 6046 29023 6047
rect 28936 6037 29023 6046
rect 28936 6017 28994 6037
rect 29014 6017 29023 6037
rect 28936 6007 29023 6017
rect 29082 6037 29119 6047
rect 29082 6017 29090 6037
rect 29110 6017 29119 6037
rect 28936 6006 28967 6007
rect 28931 5938 29041 5951
rect 29082 5938 29119 6017
rect 28869 5936 29119 5938
rect 28869 5933 28970 5936
rect 28869 5914 28934 5933
rect 28931 5906 28934 5914
rect 28963 5906 28970 5933
rect 28998 5909 29008 5936
rect 29037 5914 29119 5936
rect 29037 5909 29041 5914
rect 28998 5906 29041 5909
rect 28931 5892 29041 5906
rect 28357 5874 28698 5875
rect 28282 5869 28698 5874
rect 28282 5849 28285 5869
rect 28305 5849 28699 5869
rect 28508 5816 28545 5826
rect 28508 5779 28517 5816
rect 28534 5779 28545 5816
rect 28508 5758 28545 5779
rect 28217 4819 28385 4820
rect 28514 4819 28543 5758
rect 28656 5144 28699 5849
rect 28657 5136 28699 5144
rect 28657 5125 28702 5136
rect 28657 5087 28667 5125
rect 28692 5087 28702 5125
rect 28657 5078 28702 5087
rect 28217 4793 28661 4819
rect 28217 4791 28385 4793
rect 28217 4524 28244 4791
rect 28514 4789 28543 4793
rect 28284 4664 28348 4676
rect 28624 4672 28661 4793
rect 28889 4761 29000 4776
rect 28889 4759 28931 4761
rect 28889 4739 28896 4759
rect 28915 4739 28931 4759
rect 28889 4731 28931 4739
rect 28959 4759 29000 4761
rect 28959 4739 28973 4759
rect 28992 4739 29000 4759
rect 28959 4731 29000 4739
rect 28889 4725 29000 4731
rect 28832 4703 29081 4725
rect 28832 4672 28869 4703
rect 29045 4701 29081 4703
rect 29045 4672 29082 4701
rect 28284 4663 28319 4664
rect 28261 4658 28319 4663
rect 28261 4638 28264 4658
rect 28284 4644 28319 4658
rect 28339 4644 28348 4664
rect 28284 4636 28348 4644
rect 28310 4635 28348 4636
rect 28311 4634 28348 4635
rect 28414 4668 28450 4669
rect 28522 4668 28558 4669
rect 28414 4660 28558 4668
rect 28414 4640 28422 4660
rect 28442 4640 28530 4660
rect 28550 4640 28558 4660
rect 28414 4634 28558 4640
rect 28624 4664 28662 4672
rect 28730 4668 28766 4669
rect 28624 4644 28633 4664
rect 28653 4644 28662 4664
rect 28624 4635 28662 4644
rect 28681 4661 28766 4668
rect 28681 4641 28688 4661
rect 28709 4660 28766 4661
rect 28709 4641 28738 4660
rect 28681 4640 28738 4641
rect 28758 4640 28766 4660
rect 28624 4634 28661 4635
rect 28681 4634 28766 4640
rect 28832 4664 28870 4672
rect 28943 4668 28979 4669
rect 28832 4644 28841 4664
rect 28861 4644 28870 4664
rect 28832 4635 28870 4644
rect 28894 4660 28979 4668
rect 28894 4640 28951 4660
rect 28971 4640 28979 4660
rect 28832 4634 28869 4635
rect 28894 4634 28979 4640
rect 29045 4664 29083 4672
rect 29045 4644 29054 4664
rect 29074 4644 29083 4664
rect 29045 4635 29083 4644
rect 29045 4634 29082 4635
rect 28468 4613 28504 4634
rect 28894 4613 28925 4634
rect 29319 4617 29411 7921
rect 29517 6154 29589 7993
rect 30619 7943 30691 7960
rect 30619 7895 30631 7943
rect 30677 7895 30691 7943
rect 31159 7923 31200 7925
rect 31431 7923 31535 7925
rect 31890 7923 31955 8080
rect 32933 7938 32998 8095
rect 33353 8093 33457 8095
rect 33688 8093 33729 8095
rect 34197 8075 34211 8123
rect 34257 8075 34269 8123
rect 34197 8058 34269 8075
rect 35299 8025 35371 9864
rect 35477 8097 35569 11401
rect 35963 11384 35994 11405
rect 36384 11384 36420 11405
rect 35806 11383 35843 11384
rect 35805 11374 35843 11383
rect 35805 11354 35814 11374
rect 35834 11354 35843 11374
rect 35805 11346 35843 11354
rect 35909 11378 35994 11384
rect 36019 11383 36056 11384
rect 35909 11358 35917 11378
rect 35937 11358 35994 11378
rect 35909 11350 35994 11358
rect 36018 11374 36056 11383
rect 36018 11354 36027 11374
rect 36047 11354 36056 11374
rect 35909 11349 35945 11350
rect 36018 11346 36056 11354
rect 36122 11378 36207 11384
rect 36227 11383 36264 11384
rect 36122 11358 36130 11378
rect 36150 11377 36207 11378
rect 36150 11358 36179 11377
rect 36122 11357 36179 11358
rect 36200 11357 36207 11377
rect 36122 11350 36207 11357
rect 36226 11374 36264 11383
rect 36226 11354 36235 11374
rect 36255 11354 36264 11374
rect 36122 11349 36158 11350
rect 36226 11346 36264 11354
rect 36330 11378 36474 11384
rect 36330 11358 36338 11378
rect 36358 11358 36446 11378
rect 36466 11358 36474 11378
rect 36330 11350 36474 11358
rect 36330 11349 36366 11350
rect 36438 11349 36474 11350
rect 36540 11383 36577 11384
rect 36540 11382 36578 11383
rect 36540 11374 36604 11382
rect 36540 11354 36549 11374
rect 36569 11360 36604 11374
rect 36624 11360 36627 11380
rect 36569 11355 36627 11360
rect 36569 11354 36604 11355
rect 35806 11317 35843 11346
rect 35807 11315 35843 11317
rect 36019 11315 36056 11346
rect 35807 11293 36056 11315
rect 35888 11287 35999 11293
rect 35888 11279 35929 11287
rect 35888 11259 35896 11279
rect 35915 11259 35929 11279
rect 35888 11257 35929 11259
rect 35957 11279 35999 11287
rect 35957 11259 35973 11279
rect 35992 11259 35999 11279
rect 35957 11257 35999 11259
rect 35888 11242 35999 11257
rect 36227 11225 36264 11346
rect 36540 11342 36604 11354
rect 36345 11225 36374 11229
rect 36644 11227 36671 11494
rect 36503 11225 36671 11227
rect 36227 11199 36671 11225
rect 36186 10931 36231 10940
rect 36186 10893 36196 10931
rect 36221 10893 36231 10931
rect 36186 10882 36231 10893
rect 36189 10874 36231 10882
rect 36189 10169 36232 10874
rect 36345 10260 36374 11199
rect 36503 11198 36671 11199
rect 36343 10239 36380 10260
rect 36343 10202 36354 10239
rect 36371 10202 36380 10239
rect 36343 10192 36380 10202
rect 36189 10149 36583 10169
rect 36603 10149 36606 10169
rect 36190 10144 36606 10149
rect 36190 10143 36531 10144
rect 35847 10112 35957 10126
rect 35847 10109 35890 10112
rect 35847 10104 35851 10109
rect 35769 10082 35851 10104
rect 35880 10082 35890 10109
rect 35918 10085 35925 10112
rect 35954 10104 35957 10112
rect 35954 10085 36019 10104
rect 35918 10082 36019 10085
rect 35769 10080 36019 10082
rect 35769 10001 35806 10080
rect 35847 10067 35957 10080
rect 35921 10011 35952 10012
rect 35769 9981 35778 10001
rect 35798 9981 35806 10001
rect 35769 9971 35806 9981
rect 35865 10001 35952 10011
rect 35865 9981 35874 10001
rect 35894 9981 35952 10001
rect 35865 9972 35952 9981
rect 35865 9971 35902 9972
rect 35921 9919 35952 9972
rect 35982 10001 36019 10080
rect 36134 10011 36165 10012
rect 35982 9981 35991 10001
rect 36011 9981 36019 10001
rect 35982 9971 36019 9981
rect 36078 10004 36165 10011
rect 36078 10001 36139 10004
rect 36078 9981 36087 10001
rect 36107 9984 36139 10001
rect 36160 9984 36165 10004
rect 36107 9981 36165 9984
rect 36078 9974 36165 9981
rect 36190 10001 36227 10143
rect 36493 10142 36530 10143
rect 36342 10011 36378 10012
rect 36190 9981 36199 10001
rect 36219 9981 36227 10001
rect 36078 9972 36134 9974
rect 36078 9971 36115 9972
rect 36190 9971 36227 9981
rect 36286 10001 36434 10011
rect 36534 10008 36630 10010
rect 36286 9981 36295 10001
rect 36315 9981 36405 10001
rect 36425 9981 36434 10001
rect 36286 9975 36434 9981
rect 36286 9972 36350 9975
rect 36286 9971 36323 9972
rect 36342 9945 36350 9972
rect 36371 9972 36434 9975
rect 36492 10001 36630 10008
rect 36492 9981 36501 10001
rect 36521 9981 36630 10001
rect 36492 9972 36630 9981
rect 36371 9945 36378 9972
rect 36397 9971 36434 9972
rect 36493 9971 36530 9972
rect 36342 9920 36378 9945
rect 35813 9918 35854 9919
rect 35733 9913 35854 9918
rect 35684 9911 35854 9913
rect 35684 9900 35823 9911
rect 35684 9877 35707 9900
rect 35733 9891 35823 9900
rect 35843 9891 35854 9911
rect 35733 9883 35854 9891
rect 35921 9915 36280 9919
rect 35921 9910 36243 9915
rect 35921 9886 36034 9910
rect 36058 9891 36243 9910
rect 36267 9891 36280 9915
rect 36058 9886 36280 9891
rect 35921 9883 36280 9886
rect 36342 9883 36377 9920
rect 36445 9917 36545 9920
rect 36445 9913 36512 9917
rect 36445 9887 36457 9913
rect 36483 9891 36512 9913
rect 36538 9891 36545 9917
rect 36483 9887 36545 9891
rect 36445 9883 36545 9887
rect 35733 9877 35741 9883
rect 35684 9869 35741 9877
rect 35921 9862 35952 9883
rect 36342 9862 36378 9883
rect 35764 9861 35801 9862
rect 35763 9852 35801 9861
rect 35763 9832 35772 9852
rect 35792 9832 35801 9852
rect 35763 9824 35801 9832
rect 35867 9856 35952 9862
rect 35977 9861 36014 9862
rect 35867 9836 35875 9856
rect 35895 9836 35952 9856
rect 35867 9828 35952 9836
rect 35976 9852 36014 9861
rect 35976 9832 35985 9852
rect 36005 9832 36014 9852
rect 35867 9827 35903 9828
rect 35976 9824 36014 9832
rect 36080 9856 36165 9862
rect 36185 9861 36222 9862
rect 36080 9836 36088 9856
rect 36108 9855 36165 9856
rect 36108 9836 36137 9855
rect 36080 9835 36137 9836
rect 36158 9835 36165 9855
rect 36080 9828 36165 9835
rect 36184 9852 36222 9861
rect 36184 9832 36193 9852
rect 36213 9832 36222 9852
rect 36080 9827 36116 9828
rect 36184 9824 36222 9832
rect 36288 9856 36432 9862
rect 36288 9836 36296 9856
rect 36316 9836 36404 9856
rect 36424 9836 36432 9856
rect 36288 9828 36432 9836
rect 36288 9827 36324 9828
rect 36396 9827 36432 9828
rect 36498 9861 36535 9862
rect 36498 9860 36536 9861
rect 36498 9852 36562 9860
rect 36498 9832 36507 9852
rect 36527 9838 36562 9852
rect 36582 9838 36585 9858
rect 36527 9833 36585 9838
rect 36527 9832 36562 9833
rect 35764 9795 35801 9824
rect 35765 9793 35801 9795
rect 35977 9793 36014 9824
rect 35765 9771 36014 9793
rect 35846 9765 35957 9771
rect 35846 9757 35887 9765
rect 35846 9737 35854 9757
rect 35873 9737 35887 9757
rect 35846 9735 35887 9737
rect 35915 9757 35957 9765
rect 35915 9737 35931 9757
rect 35950 9737 35957 9757
rect 35915 9735 35957 9737
rect 35846 9720 35957 9735
rect 36185 9709 36222 9824
rect 36498 9820 36562 9832
rect 36178 9703 36225 9709
rect 36602 9705 36629 9972
rect 36461 9703 36629 9705
rect 36178 9677 36629 9703
rect 36178 9542 36225 9677
rect 36461 9676 36629 9677
rect 36176 9493 36235 9542
rect 36176 9465 36194 9493
rect 36222 9465 36235 9493
rect 36176 9455 36235 9465
rect 37291 8718 37369 11758
rect 37291 8698 37691 8718
rect 37711 8698 37714 8718
rect 37291 8696 37714 8698
rect 37298 8693 37714 8696
rect 37298 8692 37639 8693
rect 36955 8661 37065 8675
rect 36955 8658 36998 8661
rect 36955 8653 36959 8658
rect 36877 8631 36959 8653
rect 36988 8631 36998 8658
rect 37026 8634 37033 8661
rect 37062 8653 37065 8661
rect 37062 8634 37127 8653
rect 37026 8631 37127 8634
rect 36877 8629 37127 8631
rect 36877 8550 36914 8629
rect 36955 8616 37065 8629
rect 37029 8560 37060 8561
rect 36877 8530 36886 8550
rect 36906 8530 36914 8550
rect 36877 8520 36914 8530
rect 36973 8550 37060 8560
rect 36973 8530 36982 8550
rect 37002 8530 37060 8550
rect 36973 8521 37060 8530
rect 36973 8520 37010 8521
rect 36747 8467 36858 8470
rect 37029 8468 37060 8521
rect 37090 8550 37127 8629
rect 37242 8560 37273 8561
rect 37090 8530 37099 8550
rect 37119 8530 37127 8550
rect 37090 8520 37127 8530
rect 37186 8553 37273 8560
rect 37186 8550 37247 8553
rect 37186 8530 37195 8550
rect 37215 8533 37247 8550
rect 37268 8533 37273 8553
rect 37215 8530 37273 8533
rect 37186 8523 37273 8530
rect 37298 8550 37335 8692
rect 37601 8691 37638 8692
rect 37450 8560 37486 8561
rect 37298 8530 37307 8550
rect 37327 8530 37335 8550
rect 37186 8521 37242 8523
rect 37186 8520 37223 8521
rect 37298 8520 37335 8530
rect 37394 8550 37542 8560
rect 37642 8557 37738 8559
rect 37394 8530 37403 8550
rect 37423 8530 37513 8550
rect 37533 8530 37542 8550
rect 37394 8524 37542 8530
rect 37394 8521 37458 8524
rect 37394 8520 37431 8521
rect 37450 8494 37458 8521
rect 37479 8521 37542 8524
rect 37600 8550 37738 8557
rect 37600 8530 37609 8550
rect 37629 8530 37738 8550
rect 37600 8521 37738 8530
rect 37479 8494 37486 8521
rect 37505 8520 37542 8521
rect 37601 8520 37638 8521
rect 37450 8469 37486 8494
rect 36921 8467 36962 8468
rect 36747 8460 36962 8467
rect 36747 8459 36812 8460
rect 36747 8435 36755 8459
rect 36779 8436 36812 8459
rect 36836 8440 36931 8460
rect 36951 8440 36962 8460
rect 36836 8436 36962 8440
rect 36779 8435 36962 8436
rect 36747 8432 36962 8435
rect 37029 8464 37388 8468
rect 37029 8459 37351 8464
rect 37029 8435 37142 8459
rect 37166 8440 37351 8459
rect 37375 8440 37388 8464
rect 37166 8435 37388 8440
rect 37029 8432 37388 8435
rect 37450 8432 37485 8469
rect 37553 8466 37653 8469
rect 37553 8462 37620 8466
rect 37553 8436 37565 8462
rect 37591 8440 37620 8462
rect 37646 8440 37653 8466
rect 37591 8436 37653 8440
rect 37553 8432 37653 8436
rect 36747 8428 36858 8432
rect 37029 8411 37060 8432
rect 37450 8411 37486 8432
rect 36872 8410 36909 8411
rect 36871 8401 36909 8410
rect 36871 8381 36880 8401
rect 36900 8381 36909 8401
rect 36871 8373 36909 8381
rect 36975 8405 37060 8411
rect 37085 8410 37122 8411
rect 36975 8385 36983 8405
rect 37003 8385 37060 8405
rect 36975 8377 37060 8385
rect 37084 8401 37122 8410
rect 37084 8381 37093 8401
rect 37113 8381 37122 8401
rect 36975 8376 37011 8377
rect 37084 8373 37122 8381
rect 37188 8405 37273 8411
rect 37293 8410 37330 8411
rect 37188 8385 37196 8405
rect 37216 8404 37273 8405
rect 37216 8385 37245 8404
rect 37188 8384 37245 8385
rect 37266 8384 37273 8404
rect 37188 8377 37273 8384
rect 37292 8401 37330 8410
rect 37292 8381 37301 8401
rect 37321 8381 37330 8401
rect 37188 8376 37224 8377
rect 37292 8373 37330 8381
rect 37396 8405 37540 8411
rect 37396 8385 37404 8405
rect 37424 8404 37512 8405
rect 37424 8385 37458 8404
rect 37396 8382 37458 8385
rect 37482 8385 37512 8404
rect 37532 8385 37540 8405
rect 37482 8382 37540 8385
rect 37396 8377 37540 8382
rect 37396 8376 37432 8377
rect 37504 8376 37540 8377
rect 37606 8410 37643 8411
rect 37606 8409 37644 8410
rect 37606 8401 37670 8409
rect 37606 8381 37615 8401
rect 37635 8387 37670 8401
rect 37690 8387 37693 8407
rect 37635 8382 37693 8387
rect 37635 8381 37670 8382
rect 36872 8344 36909 8373
rect 36873 8342 36909 8344
rect 37085 8342 37122 8373
rect 36873 8320 37122 8342
rect 36954 8314 37065 8320
rect 36954 8306 36995 8314
rect 36954 8286 36962 8306
rect 36981 8286 36995 8306
rect 36954 8284 36995 8286
rect 37023 8306 37065 8314
rect 37023 8286 37039 8306
rect 37058 8286 37065 8306
rect 37023 8284 37065 8286
rect 36954 8269 37065 8284
rect 37293 8258 37330 8373
rect 37606 8369 37670 8381
rect 37289 8252 37344 8258
rect 37710 8254 37737 8521
rect 37569 8252 37737 8254
rect 37289 8227 37737 8252
rect 38050 8312 38156 13565
rect 41322 13553 41341 13579
rect 41381 13553 41402 13579
rect 41322 13526 41402 13553
rect 41322 13500 41345 13526
rect 41385 13500 41402 13526
rect 41322 13489 41402 13500
rect 41464 13490 41491 13745
rect 41869 13737 41910 13887
rect 42141 13742 42245 13887
rect 42336 13825 42457 13843
rect 42336 13823 42407 13825
rect 42336 13782 42351 13823
rect 42388 13784 42407 13823
rect 42444 13784 42457 13825
rect 42388 13782 42457 13784
rect 42336 13772 42457 13782
rect 41531 13630 41595 13642
rect 41871 13638 41908 13737
rect 42136 13727 42247 13742
rect 42136 13725 42178 13727
rect 42136 13705 42143 13725
rect 42162 13705 42178 13725
rect 42136 13697 42178 13705
rect 42206 13725 42247 13727
rect 42206 13705 42220 13725
rect 42239 13705 42247 13725
rect 42206 13697 42247 13705
rect 42136 13691 42247 13697
rect 42079 13669 42328 13691
rect 42079 13638 42116 13669
rect 42292 13667 42328 13669
rect 42292 13638 42329 13667
rect 41531 13629 41566 13630
rect 41508 13624 41566 13629
rect 41508 13604 41511 13624
rect 41531 13610 41566 13624
rect 41586 13610 41595 13630
rect 41531 13602 41595 13610
rect 41557 13601 41595 13602
rect 41558 13600 41595 13601
rect 41661 13634 41697 13635
rect 41769 13634 41805 13635
rect 41661 13626 41805 13634
rect 41661 13606 41669 13626
rect 41689 13606 41777 13626
rect 41797 13606 41805 13626
rect 41661 13600 41805 13606
rect 41871 13630 41909 13638
rect 41977 13634 42013 13635
rect 41871 13610 41880 13630
rect 41900 13610 41909 13630
rect 41871 13601 41909 13610
rect 41928 13627 42013 13634
rect 41928 13607 41935 13627
rect 41956 13626 42013 13627
rect 41956 13607 41985 13626
rect 41928 13606 41985 13607
rect 42005 13606 42013 13626
rect 41871 13600 41908 13601
rect 41928 13600 42013 13606
rect 42079 13630 42117 13638
rect 42190 13634 42226 13635
rect 42079 13610 42088 13630
rect 42108 13610 42117 13630
rect 42079 13601 42117 13610
rect 42141 13626 42226 13634
rect 42141 13606 42198 13626
rect 42218 13606 42226 13626
rect 42079 13600 42116 13601
rect 42141 13600 42226 13606
rect 42292 13630 42330 13638
rect 42292 13610 42301 13630
rect 42321 13610 42330 13630
rect 42385 13620 42450 13772
rect 42603 13746 42658 13887
rect 42292 13601 42330 13610
rect 42383 13613 42450 13620
rect 42292 13600 42329 13601
rect 41715 13579 41751 13600
rect 42141 13579 42172 13600
rect 42383 13592 42400 13613
rect 42436 13592 42450 13613
rect 42602 13633 42658 13746
rect 42602 13615 42621 13633
rect 42639 13615 42658 13633
rect 42602 13595 42658 13615
rect 42383 13579 42450 13592
rect 41548 13575 41648 13579
rect 41548 13571 41610 13575
rect 41548 13545 41555 13571
rect 41581 13549 41610 13571
rect 41636 13549 41648 13575
rect 41581 13545 41648 13549
rect 41548 13542 41648 13545
rect 41716 13542 41751 13579
rect 41813 13576 42172 13579
rect 41813 13571 42035 13576
rect 41813 13547 41826 13571
rect 41850 13552 42035 13571
rect 42059 13552 42172 13576
rect 41850 13547 42172 13552
rect 41813 13543 42172 13547
rect 42239 13573 42450 13579
rect 42239 13571 42400 13573
rect 42239 13551 42250 13571
rect 42270 13551 42400 13571
rect 42239 13544 42400 13551
rect 42239 13543 42280 13544
rect 41715 13517 41751 13542
rect 41563 13490 41600 13491
rect 41659 13490 41696 13491
rect 41715 13490 41722 13517
rect 41463 13481 41601 13490
rect 41463 13461 41572 13481
rect 41592 13461 41601 13481
rect 41463 13454 41601 13461
rect 41659 13487 41722 13490
rect 41743 13490 41751 13517
rect 41770 13490 41807 13491
rect 41743 13487 41807 13490
rect 41659 13481 41807 13487
rect 41659 13461 41668 13481
rect 41688 13461 41778 13481
rect 41798 13461 41807 13481
rect 41463 13452 41559 13454
rect 41659 13451 41807 13461
rect 41866 13481 41903 13491
rect 41978 13490 42015 13491
rect 41959 13488 42015 13490
rect 41866 13461 41874 13481
rect 41894 13461 41903 13481
rect 41715 13450 41751 13451
rect 41563 13319 41600 13320
rect 41866 13319 41903 13461
rect 41928 13481 42015 13488
rect 41928 13478 41986 13481
rect 41928 13458 41933 13478
rect 41954 13461 41986 13478
rect 42006 13461 42015 13481
rect 41954 13458 42015 13461
rect 41928 13451 42015 13458
rect 42074 13481 42111 13491
rect 42074 13461 42082 13481
rect 42102 13461 42111 13481
rect 41928 13450 41959 13451
rect 42074 13382 42111 13461
rect 42141 13490 42172 13543
rect 42385 13536 42400 13544
rect 42440 13536 42450 13573
rect 42385 13527 42450 13536
rect 42598 13534 42663 13555
rect 42598 13516 42623 13534
rect 42641 13516 42663 13534
rect 42191 13490 42228 13491
rect 42141 13481 42228 13490
rect 42141 13461 42199 13481
rect 42219 13461 42228 13481
rect 42141 13451 42228 13461
rect 42287 13481 42324 13491
rect 42287 13461 42295 13481
rect 42315 13461 42324 13481
rect 42141 13450 42172 13451
rect 42136 13382 42246 13395
rect 42287 13382 42324 13461
rect 42598 13440 42663 13516
rect 42074 13380 42324 13382
rect 42074 13377 42175 13380
rect 42074 13358 42139 13377
rect 42136 13350 42139 13358
rect 42168 13350 42175 13377
rect 42203 13353 42213 13380
rect 42242 13358 42324 13380
rect 42347 13405 42664 13440
rect 42242 13353 42246 13358
rect 42203 13350 42246 13353
rect 42136 13336 42246 13350
rect 41562 13318 41903 13319
rect 41487 13316 41903 13318
rect 42347 13316 42387 13405
rect 42598 13378 42663 13405
rect 42598 13360 42621 13378
rect 42639 13360 42663 13378
rect 42598 13340 42663 13360
rect 41484 13313 42387 13316
rect 41484 13293 41490 13313
rect 41510 13293 42387 13313
rect 41484 13289 42387 13293
rect 42347 13286 42387 13289
rect 42599 13279 42664 13300
rect 40817 13271 41478 13272
rect 40817 13264 41751 13271
rect 40817 13263 41723 13264
rect 40817 13243 41668 13263
rect 41700 13244 41723 13263
rect 41748 13244 41751 13264
rect 41700 13243 41751 13244
rect 40817 13236 41751 13243
rect 40416 13194 40584 13195
rect 40819 13194 40858 13236
rect 41647 13234 41751 13236
rect 41716 13232 41751 13234
rect 42599 13261 42623 13279
rect 42641 13261 42664 13279
rect 42599 13214 42664 13261
rect 40416 13168 40860 13194
rect 40416 13166 40584 13168
rect 40416 12815 40443 13166
rect 40819 13162 40860 13168
rect 40483 12955 40547 12967
rect 40823 12963 40860 13162
rect 41322 13189 41394 13206
rect 41322 13150 41330 13189
rect 41375 13150 41394 13189
rect 41088 13052 41199 13067
rect 41088 13050 41130 13052
rect 41088 13030 41095 13050
rect 41114 13030 41130 13050
rect 41088 13022 41130 13030
rect 41158 13050 41199 13052
rect 41158 13030 41172 13050
rect 41191 13030 41199 13050
rect 41158 13022 41199 13030
rect 41088 13016 41199 13022
rect 41031 12994 41280 13016
rect 41031 12963 41068 12994
rect 41244 12992 41280 12994
rect 41244 12963 41281 12992
rect 40483 12954 40518 12955
rect 40460 12949 40518 12954
rect 40460 12929 40463 12949
rect 40483 12935 40518 12949
rect 40538 12935 40547 12955
rect 40483 12927 40547 12935
rect 40509 12926 40547 12927
rect 40510 12925 40547 12926
rect 40613 12959 40649 12960
rect 40721 12959 40757 12960
rect 40613 12951 40757 12959
rect 40613 12931 40621 12951
rect 40641 12931 40729 12951
rect 40749 12931 40757 12951
rect 40613 12925 40757 12931
rect 40823 12955 40861 12963
rect 40929 12959 40965 12960
rect 40823 12935 40832 12955
rect 40852 12935 40861 12955
rect 40823 12926 40861 12935
rect 40880 12952 40965 12959
rect 40880 12932 40887 12952
rect 40908 12951 40965 12952
rect 40908 12932 40937 12951
rect 40880 12931 40937 12932
rect 40957 12931 40965 12951
rect 40823 12925 40860 12926
rect 40880 12925 40965 12931
rect 41031 12955 41069 12963
rect 41142 12959 41178 12960
rect 41031 12935 41040 12955
rect 41060 12935 41069 12955
rect 41031 12926 41069 12935
rect 41093 12951 41178 12959
rect 41093 12931 41150 12951
rect 41170 12931 41178 12951
rect 41031 12925 41068 12926
rect 41093 12925 41178 12931
rect 41244 12955 41282 12963
rect 41244 12935 41253 12955
rect 41273 12935 41282 12955
rect 41244 12926 41282 12935
rect 41322 12940 41394 13150
rect 41464 13184 42664 13214
rect 41464 13183 41908 13184
rect 41464 13181 41632 13183
rect 41322 12926 41405 12940
rect 41244 12925 41281 12926
rect 40667 12904 40703 12925
rect 41093 12904 41124 12925
rect 41322 12904 41339 12926
rect 40500 12900 40600 12904
rect 40500 12896 40562 12900
rect 40500 12870 40507 12896
rect 40533 12874 40562 12896
rect 40588 12874 40600 12900
rect 40533 12870 40600 12874
rect 40500 12867 40600 12870
rect 40668 12867 40703 12904
rect 40765 12901 41124 12904
rect 40765 12896 40987 12901
rect 40765 12872 40778 12896
rect 40802 12877 40987 12896
rect 41011 12877 41124 12901
rect 40802 12872 41124 12877
rect 40765 12868 41124 12872
rect 41191 12896 41339 12904
rect 41191 12876 41202 12896
rect 41222 12893 41339 12896
rect 41392 12893 41405 12926
rect 41222 12876 41405 12893
rect 41191 12869 41405 12876
rect 41191 12868 41232 12869
rect 41322 12868 41405 12869
rect 40667 12842 40703 12867
rect 40515 12815 40552 12816
rect 40611 12815 40648 12816
rect 40667 12815 40674 12842
rect 40415 12806 40553 12815
rect 40415 12786 40524 12806
rect 40544 12786 40553 12806
rect 40415 12779 40553 12786
rect 40611 12812 40674 12815
rect 40695 12815 40703 12842
rect 40722 12815 40759 12816
rect 40695 12812 40759 12815
rect 40611 12806 40759 12812
rect 40611 12786 40620 12806
rect 40640 12786 40730 12806
rect 40750 12786 40759 12806
rect 40415 12777 40511 12779
rect 40611 12776 40759 12786
rect 40818 12806 40855 12816
rect 40930 12815 40967 12816
rect 40911 12813 40967 12815
rect 40818 12786 40826 12806
rect 40846 12786 40855 12806
rect 40667 12775 40703 12776
rect 40515 12644 40552 12645
rect 40818 12644 40855 12786
rect 40880 12806 40967 12813
rect 40880 12803 40938 12806
rect 40880 12783 40885 12803
rect 40906 12786 40938 12803
rect 40958 12786 40967 12806
rect 40906 12783 40967 12786
rect 40880 12776 40967 12783
rect 41026 12806 41063 12816
rect 41026 12786 41034 12806
rect 41054 12786 41063 12806
rect 40880 12775 40911 12776
rect 41026 12707 41063 12786
rect 41093 12815 41124 12868
rect 41330 12835 41344 12868
rect 41397 12835 41405 12868
rect 41330 12829 41405 12835
rect 41330 12824 41400 12829
rect 41143 12815 41180 12816
rect 41093 12806 41180 12815
rect 41093 12786 41151 12806
rect 41171 12786 41180 12806
rect 41093 12776 41180 12786
rect 41239 12806 41276 12816
rect 41464 12811 41491 13181
rect 41531 12951 41595 12963
rect 41871 12959 41908 13183
rect 42379 13164 42443 13166
rect 42375 13152 42443 13164
rect 42375 13119 42386 13152
rect 42426 13119 42443 13152
rect 42375 13109 42443 13119
rect 42136 13048 42247 13063
rect 42136 13046 42178 13048
rect 42136 13026 42143 13046
rect 42162 13026 42178 13046
rect 42136 13018 42178 13026
rect 42206 13046 42247 13048
rect 42206 13026 42220 13046
rect 42239 13026 42247 13046
rect 42206 13018 42247 13026
rect 42136 13012 42247 13018
rect 42079 12990 42328 13012
rect 42079 12959 42116 12990
rect 42292 12988 42328 12990
rect 42292 12959 42329 12988
rect 41531 12950 41566 12951
rect 41508 12945 41566 12950
rect 41508 12925 41511 12945
rect 41531 12931 41566 12945
rect 41586 12931 41595 12951
rect 41531 12923 41595 12931
rect 41557 12922 41595 12923
rect 41558 12921 41595 12922
rect 41661 12955 41697 12956
rect 41769 12955 41805 12956
rect 41661 12947 41805 12955
rect 41661 12927 41669 12947
rect 41689 12927 41777 12947
rect 41797 12927 41805 12947
rect 41661 12921 41805 12927
rect 41871 12951 41909 12959
rect 41977 12955 42013 12956
rect 41871 12931 41880 12951
rect 41900 12931 41909 12951
rect 41871 12922 41909 12931
rect 41928 12948 42013 12955
rect 41928 12928 41935 12948
rect 41956 12947 42013 12948
rect 41956 12928 41985 12947
rect 41928 12927 41985 12928
rect 42005 12927 42013 12947
rect 41871 12921 41908 12922
rect 41928 12921 42013 12927
rect 42079 12951 42117 12959
rect 42190 12955 42226 12956
rect 42079 12931 42088 12951
rect 42108 12931 42117 12951
rect 42079 12922 42117 12931
rect 42141 12947 42226 12955
rect 42141 12927 42198 12947
rect 42218 12927 42226 12947
rect 42079 12921 42116 12922
rect 42141 12921 42226 12927
rect 42292 12951 42330 12959
rect 42292 12931 42301 12951
rect 42321 12931 42330 12951
rect 42292 12922 42330 12931
rect 42379 12925 42443 13109
rect 42599 12983 42664 13184
rect 42599 12965 42621 12983
rect 42639 12965 42664 12983
rect 42599 12946 42664 12965
rect 42292 12921 42329 12922
rect 41715 12900 41751 12921
rect 42141 12900 42172 12921
rect 42379 12916 42387 12925
rect 42376 12900 42387 12916
rect 41548 12896 41648 12900
rect 41548 12892 41610 12896
rect 41548 12866 41555 12892
rect 41581 12870 41610 12892
rect 41636 12870 41648 12896
rect 41581 12866 41648 12870
rect 41548 12863 41648 12866
rect 41716 12863 41751 12900
rect 41813 12897 42172 12900
rect 41813 12892 42035 12897
rect 41813 12868 41826 12892
rect 41850 12873 42035 12892
rect 42059 12873 42172 12897
rect 41850 12868 42172 12873
rect 41813 12864 42172 12868
rect 42239 12892 42387 12900
rect 42239 12872 42250 12892
rect 42270 12883 42387 12892
rect 42436 12916 42443 12925
rect 42436 12883 42444 12916
rect 42270 12872 42444 12883
rect 42239 12865 42444 12872
rect 42239 12864 42280 12865
rect 41715 12838 41751 12863
rect 41563 12811 41600 12812
rect 41659 12811 41696 12812
rect 41715 12811 41722 12838
rect 41239 12786 41247 12806
rect 41267 12786 41276 12806
rect 41093 12775 41124 12776
rect 41088 12707 41198 12720
rect 41239 12707 41276 12786
rect 41463 12802 41601 12811
rect 41463 12782 41572 12802
rect 41592 12782 41601 12802
rect 41463 12775 41601 12782
rect 41659 12808 41722 12811
rect 41743 12811 41751 12838
rect 41770 12811 41807 12812
rect 41743 12808 41807 12811
rect 41659 12802 41807 12808
rect 41659 12782 41668 12802
rect 41688 12782 41778 12802
rect 41798 12782 41807 12802
rect 41463 12773 41559 12775
rect 41659 12772 41807 12782
rect 41866 12802 41903 12812
rect 41978 12811 42015 12812
rect 41959 12809 42015 12811
rect 41866 12782 41874 12802
rect 41894 12782 41903 12802
rect 41715 12771 41751 12772
rect 41026 12705 41276 12707
rect 41026 12702 41127 12705
rect 41026 12683 41091 12702
rect 41088 12675 41091 12683
rect 41120 12675 41127 12702
rect 41155 12678 41165 12705
rect 41194 12683 41276 12705
rect 41194 12678 41198 12683
rect 41155 12675 41198 12678
rect 41088 12661 41198 12675
rect 40514 12643 40855 12644
rect 40439 12638 40855 12643
rect 41563 12640 41600 12641
rect 41866 12640 41903 12782
rect 41928 12802 42015 12809
rect 41928 12799 41986 12802
rect 41928 12779 41933 12799
rect 41954 12782 41986 12799
rect 42006 12782 42015 12802
rect 41954 12779 42015 12782
rect 41928 12772 42015 12779
rect 42074 12802 42111 12812
rect 42074 12782 42082 12802
rect 42102 12782 42111 12802
rect 41928 12771 41959 12772
rect 42074 12703 42111 12782
rect 42141 12811 42172 12864
rect 42376 12862 42444 12865
rect 42376 12820 42388 12862
rect 42437 12820 42444 12862
rect 42191 12811 42228 12812
rect 42141 12802 42228 12811
rect 42141 12782 42199 12802
rect 42219 12782 42228 12802
rect 42141 12772 42228 12782
rect 42287 12802 42324 12812
rect 42376 12807 42444 12820
rect 42599 12884 42664 12901
rect 42599 12866 42623 12884
rect 42641 12866 42664 12884
rect 42287 12782 42295 12802
rect 42315 12782 42324 12802
rect 42141 12771 42172 12772
rect 42136 12703 42246 12716
rect 42287 12703 42324 12782
rect 42599 12727 42664 12866
rect 42599 12721 42621 12727
rect 42074 12701 42324 12703
rect 42074 12698 42175 12701
rect 42074 12679 42139 12698
rect 42136 12671 42139 12679
rect 42168 12671 42175 12698
rect 42203 12674 42213 12701
rect 42242 12679 42324 12701
rect 42353 12709 42621 12721
rect 42639 12709 42664 12727
rect 42353 12686 42664 12709
rect 42353 12685 42408 12686
rect 42242 12674 42246 12679
rect 42203 12671 42246 12674
rect 42136 12657 42246 12671
rect 41562 12639 41903 12640
rect 40439 12618 40442 12638
rect 40462 12618 40855 12638
rect 41487 12638 41903 12639
rect 42353 12638 42396 12685
rect 41487 12634 42396 12638
rect 40806 12585 40851 12618
rect 41487 12614 41490 12634
rect 41510 12614 42396 12634
rect 41864 12609 42396 12614
rect 42604 12628 42663 12650
rect 42604 12610 42623 12628
rect 42641 12610 42663 12628
rect 41652 12585 41751 12587
rect 40806 12575 41751 12585
rect 39363 12555 39422 12565
rect 39363 12527 39376 12555
rect 39404 12527 39422 12555
rect 40806 12549 41674 12575
rect 40807 12548 41674 12549
rect 41652 12537 41674 12548
rect 41699 12540 41718 12575
rect 41743 12540 41751 12575
rect 41699 12537 41751 12540
rect 42604 12539 42663 12610
rect 41652 12529 41751 12537
rect 41678 12528 41750 12529
rect 39363 12478 39422 12527
rect 41332 12502 41399 12521
rect 41332 12481 41349 12502
rect 38969 12343 39137 12344
rect 39373 12343 39420 12478
rect 38969 12317 39420 12343
rect 38969 12315 39137 12317
rect 38969 12048 38996 12315
rect 39373 12311 39420 12317
rect 41330 12436 41349 12481
rect 41379 12481 41399 12502
rect 41379 12436 41400 12481
rect 41869 12478 41910 12480
rect 42141 12478 42245 12480
rect 42601 12478 42665 12539
rect 39036 12188 39100 12200
rect 39376 12196 39413 12311
rect 39641 12285 39752 12300
rect 39641 12283 39683 12285
rect 39641 12263 39648 12283
rect 39667 12263 39683 12283
rect 39641 12255 39683 12263
rect 39711 12283 39752 12285
rect 39711 12263 39725 12283
rect 39744 12263 39752 12283
rect 39711 12255 39752 12263
rect 39641 12249 39752 12255
rect 39584 12227 39833 12249
rect 41330 12228 41400 12436
rect 41462 12443 42665 12478
rect 41462 12429 41490 12443
rect 41464 12298 41490 12429
rect 41869 12440 42665 12443
rect 39584 12196 39621 12227
rect 39797 12225 39833 12227
rect 39797 12196 39834 12225
rect 39036 12187 39071 12188
rect 39013 12182 39071 12187
rect 39013 12162 39016 12182
rect 39036 12168 39071 12182
rect 39091 12168 39100 12188
rect 39036 12160 39100 12168
rect 39062 12159 39100 12160
rect 39063 12158 39100 12159
rect 39166 12192 39202 12193
rect 39274 12192 39310 12193
rect 39166 12184 39310 12192
rect 39166 12164 39174 12184
rect 39194 12164 39282 12184
rect 39302 12164 39310 12184
rect 39166 12158 39310 12164
rect 39376 12188 39414 12196
rect 39482 12192 39518 12193
rect 39376 12168 39385 12188
rect 39405 12168 39414 12188
rect 39376 12159 39414 12168
rect 39433 12185 39518 12192
rect 39433 12165 39440 12185
rect 39461 12184 39518 12185
rect 39461 12165 39490 12184
rect 39433 12164 39490 12165
rect 39510 12164 39518 12184
rect 39376 12158 39413 12159
rect 39433 12158 39518 12164
rect 39584 12188 39622 12196
rect 39695 12192 39731 12193
rect 39584 12168 39593 12188
rect 39613 12168 39622 12188
rect 39584 12159 39622 12168
rect 39646 12184 39731 12192
rect 39646 12164 39703 12184
rect 39723 12164 39731 12184
rect 39584 12158 39621 12159
rect 39646 12158 39731 12164
rect 39797 12188 39835 12196
rect 39797 12168 39806 12188
rect 39826 12168 39835 12188
rect 39797 12159 39835 12168
rect 41322 12177 41402 12228
rect 39797 12158 39834 12159
rect 39220 12137 39256 12158
rect 39646 12137 39677 12158
rect 39857 12143 39914 12151
rect 39857 12137 39865 12143
rect 39053 12133 39153 12137
rect 39053 12129 39115 12133
rect 39053 12103 39060 12129
rect 39086 12107 39115 12129
rect 39141 12107 39153 12133
rect 39086 12103 39153 12107
rect 39053 12100 39153 12103
rect 39221 12100 39256 12137
rect 39318 12134 39677 12137
rect 39318 12129 39540 12134
rect 39318 12105 39331 12129
rect 39355 12110 39540 12129
rect 39564 12110 39677 12134
rect 39355 12105 39677 12110
rect 39318 12101 39677 12105
rect 39744 12129 39865 12137
rect 39744 12109 39755 12129
rect 39775 12120 39865 12129
rect 39891 12120 39914 12143
rect 39775 12109 39914 12120
rect 39744 12107 39914 12109
rect 40217 12136 40289 12156
rect 40217 12113 40245 12136
rect 40271 12113 40289 12136
rect 39744 12102 39865 12107
rect 39744 12101 39785 12102
rect 39220 12075 39256 12100
rect 39068 12048 39105 12049
rect 39164 12048 39201 12049
rect 39220 12048 39227 12075
rect 38968 12039 39106 12048
rect 38968 12019 39077 12039
rect 39097 12019 39106 12039
rect 38968 12012 39106 12019
rect 39164 12045 39227 12048
rect 39248 12048 39256 12075
rect 39275 12048 39312 12049
rect 39248 12045 39312 12048
rect 39164 12039 39312 12045
rect 39164 12019 39173 12039
rect 39193 12019 39283 12039
rect 39303 12019 39312 12039
rect 38968 12010 39064 12012
rect 39164 12009 39312 12019
rect 39371 12039 39408 12049
rect 39483 12048 39520 12049
rect 39464 12046 39520 12048
rect 39371 12019 39379 12039
rect 39399 12019 39408 12039
rect 39220 12008 39256 12009
rect 39068 11877 39105 11878
rect 39371 11877 39408 12019
rect 39433 12039 39520 12046
rect 39433 12036 39491 12039
rect 39433 12016 39438 12036
rect 39459 12019 39491 12036
rect 39511 12019 39520 12039
rect 39459 12016 39520 12019
rect 39433 12009 39520 12016
rect 39579 12039 39616 12049
rect 39579 12019 39587 12039
rect 39607 12019 39616 12039
rect 39433 12008 39464 12009
rect 39579 11940 39616 12019
rect 39646 12048 39677 12101
rect 40217 12051 40289 12113
rect 41322 12151 41338 12177
rect 41378 12151 41402 12177
rect 41322 12132 41402 12151
rect 41322 12106 41341 12132
rect 41381 12106 41402 12132
rect 41322 12079 41402 12106
rect 41322 12053 41345 12079
rect 41385 12053 41402 12079
rect 39696 12048 39733 12049
rect 39646 12039 39733 12048
rect 39646 12019 39704 12039
rect 39724 12019 39733 12039
rect 39646 12009 39733 12019
rect 39792 12039 39829 12049
rect 39792 12019 39800 12039
rect 39820 12019 39829 12039
rect 39646 12008 39677 12009
rect 39641 11940 39751 11953
rect 39792 11940 39829 12019
rect 39579 11938 39829 11940
rect 39579 11935 39680 11938
rect 39579 11916 39644 11935
rect 39641 11908 39644 11916
rect 39673 11908 39680 11935
rect 39708 11911 39718 11938
rect 39747 11916 39829 11938
rect 39747 11911 39751 11916
rect 39708 11908 39751 11911
rect 39641 11894 39751 11908
rect 39067 11876 39408 11877
rect 38992 11871 39408 11876
rect 38992 11851 38995 11871
rect 39015 11851 39409 11871
rect 39218 11818 39255 11828
rect 39218 11781 39227 11818
rect 39244 11781 39255 11818
rect 39218 11760 39255 11781
rect 38927 10821 39095 10822
rect 39224 10821 39253 11760
rect 39366 11146 39409 11851
rect 40221 11500 40283 12051
rect 41322 12042 41402 12053
rect 41464 12043 41491 12298
rect 41869 12290 41910 12440
rect 42141 12434 42245 12440
rect 42601 12437 42665 12440
rect 42336 12378 42457 12396
rect 42336 12376 42407 12378
rect 42336 12335 42351 12376
rect 42388 12337 42407 12376
rect 42444 12337 42457 12378
rect 42388 12335 42457 12337
rect 42336 12325 42457 12335
rect 41531 12183 41595 12195
rect 41871 12191 41908 12290
rect 42136 12280 42247 12293
rect 42136 12278 42178 12280
rect 42136 12258 42143 12278
rect 42162 12258 42178 12278
rect 42136 12250 42178 12258
rect 42206 12278 42247 12280
rect 42206 12258 42220 12278
rect 42239 12258 42247 12278
rect 42206 12250 42247 12258
rect 42136 12244 42247 12250
rect 42079 12222 42328 12244
rect 42079 12191 42116 12222
rect 42292 12220 42328 12222
rect 42292 12191 42329 12220
rect 41531 12182 41566 12183
rect 41508 12177 41566 12182
rect 41508 12157 41511 12177
rect 41531 12163 41566 12177
rect 41586 12163 41595 12183
rect 41531 12155 41595 12163
rect 41557 12154 41595 12155
rect 41558 12153 41595 12154
rect 41661 12187 41697 12188
rect 41769 12187 41805 12188
rect 41661 12179 41805 12187
rect 41661 12159 41669 12179
rect 41689 12159 41777 12179
rect 41797 12159 41805 12179
rect 41661 12153 41805 12159
rect 41871 12183 41909 12191
rect 41977 12187 42013 12188
rect 41871 12163 41880 12183
rect 41900 12163 41909 12183
rect 41871 12154 41909 12163
rect 41928 12180 42013 12187
rect 41928 12160 41935 12180
rect 41956 12179 42013 12180
rect 41956 12160 41985 12179
rect 41928 12159 41985 12160
rect 42005 12159 42013 12179
rect 41871 12153 41908 12154
rect 41928 12153 42013 12159
rect 42079 12183 42117 12191
rect 42190 12187 42226 12188
rect 42079 12163 42088 12183
rect 42108 12163 42117 12183
rect 42079 12154 42117 12163
rect 42141 12179 42226 12187
rect 42141 12159 42198 12179
rect 42218 12159 42226 12179
rect 42079 12153 42116 12154
rect 42141 12153 42226 12159
rect 42292 12183 42330 12191
rect 42292 12163 42301 12183
rect 42321 12163 42330 12183
rect 42385 12173 42450 12325
rect 42603 12299 42658 12437
rect 42292 12154 42330 12163
rect 42383 12166 42450 12173
rect 42292 12153 42329 12154
rect 41715 12132 41751 12153
rect 42141 12132 42172 12153
rect 42383 12145 42400 12166
rect 42436 12145 42450 12166
rect 42602 12186 42658 12299
rect 42602 12168 42621 12186
rect 42639 12168 42658 12186
rect 42602 12148 42658 12168
rect 42383 12132 42450 12145
rect 41548 12128 41648 12132
rect 41548 12124 41610 12128
rect 41548 12098 41555 12124
rect 41581 12102 41610 12124
rect 41636 12102 41648 12128
rect 41581 12098 41648 12102
rect 41548 12095 41648 12098
rect 41716 12095 41751 12132
rect 41813 12129 42172 12132
rect 41813 12124 42035 12129
rect 41813 12100 41826 12124
rect 41850 12105 42035 12124
rect 42059 12105 42172 12129
rect 41850 12100 42172 12105
rect 41813 12096 42172 12100
rect 42239 12126 42450 12132
rect 42239 12124 42400 12126
rect 42239 12104 42250 12124
rect 42270 12104 42400 12124
rect 42239 12097 42400 12104
rect 42239 12096 42280 12097
rect 41715 12070 41751 12095
rect 41563 12043 41600 12044
rect 41659 12043 41696 12044
rect 41715 12043 41722 12070
rect 41463 12034 41601 12043
rect 41463 12014 41572 12034
rect 41592 12014 41601 12034
rect 41463 12007 41601 12014
rect 41659 12040 41722 12043
rect 41743 12043 41751 12070
rect 41770 12043 41807 12044
rect 41743 12040 41807 12043
rect 41659 12034 41807 12040
rect 41659 12014 41668 12034
rect 41688 12014 41778 12034
rect 41798 12014 41807 12034
rect 41463 12005 41559 12007
rect 41659 12004 41807 12014
rect 41866 12034 41903 12044
rect 41978 12043 42015 12044
rect 41959 12041 42015 12043
rect 41866 12014 41874 12034
rect 41894 12014 41903 12034
rect 41715 12003 41751 12004
rect 41563 11872 41600 11873
rect 41866 11872 41903 12014
rect 41928 12034 42015 12041
rect 41928 12031 41986 12034
rect 41928 12011 41933 12031
rect 41954 12014 41986 12031
rect 42006 12014 42015 12034
rect 41954 12011 42015 12014
rect 41928 12004 42015 12011
rect 42074 12034 42111 12044
rect 42074 12014 42082 12034
rect 42102 12014 42111 12034
rect 41928 12003 41959 12004
rect 42074 11935 42111 12014
rect 42141 12043 42172 12096
rect 42385 12089 42400 12097
rect 42440 12089 42450 12126
rect 42385 12080 42450 12089
rect 42598 12087 42663 12108
rect 42598 12069 42623 12087
rect 42641 12069 42663 12087
rect 42191 12043 42228 12044
rect 42141 12034 42228 12043
rect 42141 12014 42199 12034
rect 42219 12014 42228 12034
rect 42141 12004 42228 12014
rect 42287 12034 42324 12044
rect 42287 12014 42295 12034
rect 42315 12014 42324 12034
rect 42141 12003 42172 12004
rect 42136 11935 42246 11948
rect 42287 11935 42324 12014
rect 42598 11993 42663 12069
rect 42074 11933 42324 11935
rect 42074 11930 42175 11933
rect 42074 11911 42139 11930
rect 42136 11903 42139 11911
rect 42168 11903 42175 11930
rect 42203 11906 42213 11933
rect 42242 11911 42324 11933
rect 42347 11958 42664 11993
rect 42242 11906 42246 11911
rect 42203 11903 42246 11906
rect 42136 11889 42246 11903
rect 41562 11871 41903 11872
rect 41487 11869 41903 11871
rect 42347 11869 42387 11958
rect 42598 11931 42663 11958
rect 42598 11913 42621 11931
rect 42639 11913 42663 11931
rect 42598 11893 42663 11913
rect 41484 11866 42387 11869
rect 41484 11846 41490 11866
rect 41510 11846 42387 11866
rect 41484 11842 42387 11846
rect 42347 11839 42387 11842
rect 42599 11832 42664 11853
rect 40817 11824 41478 11825
rect 40817 11817 41751 11824
rect 40817 11816 41723 11817
rect 40817 11796 41668 11816
rect 41700 11797 41723 11816
rect 41748 11797 41751 11817
rect 41700 11796 41751 11797
rect 40817 11789 41751 11796
rect 40416 11747 40584 11748
rect 40819 11747 40858 11789
rect 41647 11787 41751 11789
rect 41716 11785 41751 11787
rect 42599 11814 42623 11832
rect 42641 11814 42664 11832
rect 42599 11767 42664 11814
rect 40416 11721 40860 11747
rect 40416 11719 40584 11721
rect 40218 11416 40287 11500
rect 39367 11138 39409 11146
rect 39367 11127 39412 11138
rect 39367 11089 39377 11127
rect 39402 11089 39412 11127
rect 39367 11080 39412 11089
rect 40216 10937 40287 11416
rect 40416 11368 40443 11719
rect 40819 11715 40860 11721
rect 40483 11508 40547 11520
rect 40823 11516 40860 11715
rect 41322 11742 41394 11759
rect 41322 11703 41330 11742
rect 41375 11703 41394 11742
rect 41088 11605 41199 11620
rect 41088 11603 41130 11605
rect 41088 11583 41095 11603
rect 41114 11583 41130 11603
rect 41088 11575 41130 11583
rect 41158 11603 41199 11605
rect 41158 11583 41172 11603
rect 41191 11583 41199 11603
rect 41158 11575 41199 11583
rect 41088 11569 41199 11575
rect 41031 11547 41280 11569
rect 41031 11516 41068 11547
rect 41244 11545 41280 11547
rect 41244 11516 41281 11545
rect 40483 11507 40518 11508
rect 40460 11502 40518 11507
rect 40460 11482 40463 11502
rect 40483 11488 40518 11502
rect 40538 11488 40547 11508
rect 40483 11480 40547 11488
rect 40509 11479 40547 11480
rect 40510 11478 40547 11479
rect 40613 11512 40649 11513
rect 40721 11512 40757 11513
rect 40613 11504 40757 11512
rect 40613 11484 40621 11504
rect 40641 11484 40729 11504
rect 40749 11484 40757 11504
rect 40613 11478 40757 11484
rect 40823 11508 40861 11516
rect 40929 11512 40965 11513
rect 40823 11488 40832 11508
rect 40852 11488 40861 11508
rect 40823 11479 40861 11488
rect 40880 11505 40965 11512
rect 40880 11485 40887 11505
rect 40908 11504 40965 11505
rect 40908 11485 40937 11504
rect 40880 11484 40937 11485
rect 40957 11484 40965 11504
rect 40823 11478 40860 11479
rect 40880 11478 40965 11484
rect 41031 11508 41069 11516
rect 41142 11512 41178 11513
rect 41031 11488 41040 11508
rect 41060 11488 41069 11508
rect 41031 11479 41069 11488
rect 41093 11504 41178 11512
rect 41093 11484 41150 11504
rect 41170 11484 41178 11504
rect 41031 11478 41068 11479
rect 41093 11478 41178 11484
rect 41244 11508 41282 11516
rect 41244 11488 41253 11508
rect 41273 11488 41282 11508
rect 41244 11479 41282 11488
rect 41322 11493 41394 11703
rect 41464 11737 42664 11767
rect 41464 11736 41908 11737
rect 41464 11734 41632 11736
rect 41322 11479 41405 11493
rect 41244 11478 41281 11479
rect 40667 11457 40703 11478
rect 41093 11457 41124 11478
rect 41322 11457 41339 11479
rect 40500 11453 40600 11457
rect 40500 11449 40562 11453
rect 40500 11423 40507 11449
rect 40533 11427 40562 11449
rect 40588 11427 40600 11453
rect 40533 11423 40600 11427
rect 40500 11420 40600 11423
rect 40668 11420 40703 11457
rect 40765 11454 41124 11457
rect 40765 11449 40987 11454
rect 40765 11425 40778 11449
rect 40802 11430 40987 11449
rect 41011 11430 41124 11454
rect 40802 11425 41124 11430
rect 40765 11421 41124 11425
rect 41191 11449 41339 11457
rect 41191 11429 41202 11449
rect 41222 11446 41339 11449
rect 41392 11446 41405 11479
rect 41222 11429 41405 11446
rect 41191 11422 41405 11429
rect 41191 11421 41232 11422
rect 41322 11421 41405 11422
rect 40667 11395 40703 11420
rect 40515 11368 40552 11369
rect 40611 11368 40648 11369
rect 40667 11368 40674 11395
rect 40415 11359 40553 11368
rect 40415 11339 40524 11359
rect 40544 11339 40553 11359
rect 40415 11332 40553 11339
rect 40611 11365 40674 11368
rect 40695 11368 40703 11395
rect 40722 11368 40759 11369
rect 40695 11365 40759 11368
rect 40611 11359 40759 11365
rect 40611 11339 40620 11359
rect 40640 11339 40730 11359
rect 40750 11339 40759 11359
rect 40415 11330 40511 11332
rect 40611 11329 40759 11339
rect 40818 11359 40855 11369
rect 40930 11368 40967 11369
rect 40911 11366 40967 11368
rect 40818 11339 40826 11359
rect 40846 11339 40855 11359
rect 40667 11328 40703 11329
rect 40515 11197 40552 11198
rect 40818 11197 40855 11339
rect 40880 11359 40967 11366
rect 40880 11356 40938 11359
rect 40880 11336 40885 11356
rect 40906 11339 40938 11356
rect 40958 11339 40967 11359
rect 40906 11336 40967 11339
rect 40880 11329 40967 11336
rect 41026 11359 41063 11369
rect 41026 11339 41034 11359
rect 41054 11339 41063 11359
rect 40880 11328 40911 11329
rect 41026 11260 41063 11339
rect 41093 11368 41124 11421
rect 41330 11388 41344 11421
rect 41397 11388 41405 11421
rect 41330 11382 41405 11388
rect 41330 11377 41400 11382
rect 41143 11368 41180 11369
rect 41093 11359 41180 11368
rect 41093 11339 41151 11359
rect 41171 11339 41180 11359
rect 41093 11329 41180 11339
rect 41239 11359 41276 11369
rect 41464 11364 41491 11734
rect 41531 11504 41595 11516
rect 41871 11512 41908 11736
rect 42379 11717 42443 11719
rect 42375 11705 42443 11717
rect 42375 11672 42386 11705
rect 42426 11672 42443 11705
rect 42375 11662 42443 11672
rect 42136 11601 42247 11616
rect 42136 11599 42178 11601
rect 42136 11579 42143 11599
rect 42162 11579 42178 11599
rect 42136 11571 42178 11579
rect 42206 11599 42247 11601
rect 42206 11579 42220 11599
rect 42239 11579 42247 11599
rect 42206 11571 42247 11579
rect 42136 11565 42247 11571
rect 42079 11543 42328 11565
rect 42079 11512 42116 11543
rect 42292 11541 42328 11543
rect 42292 11512 42329 11541
rect 41531 11503 41566 11504
rect 41508 11498 41566 11503
rect 41508 11478 41511 11498
rect 41531 11484 41566 11498
rect 41586 11484 41595 11504
rect 41531 11476 41595 11484
rect 41557 11475 41595 11476
rect 41558 11474 41595 11475
rect 41661 11508 41697 11509
rect 41769 11508 41805 11509
rect 41661 11500 41805 11508
rect 41661 11480 41669 11500
rect 41689 11480 41777 11500
rect 41797 11480 41805 11500
rect 41661 11474 41805 11480
rect 41871 11504 41909 11512
rect 41977 11508 42013 11509
rect 41871 11484 41880 11504
rect 41900 11484 41909 11504
rect 41871 11475 41909 11484
rect 41928 11501 42013 11508
rect 41928 11481 41935 11501
rect 41956 11500 42013 11501
rect 41956 11481 41985 11500
rect 41928 11480 41985 11481
rect 42005 11480 42013 11500
rect 41871 11474 41908 11475
rect 41928 11474 42013 11480
rect 42079 11504 42117 11512
rect 42190 11508 42226 11509
rect 42079 11484 42088 11504
rect 42108 11484 42117 11504
rect 42079 11475 42117 11484
rect 42141 11500 42226 11508
rect 42141 11480 42198 11500
rect 42218 11480 42226 11500
rect 42079 11474 42116 11475
rect 42141 11474 42226 11480
rect 42292 11504 42330 11512
rect 42292 11484 42301 11504
rect 42321 11484 42330 11504
rect 42292 11475 42330 11484
rect 42379 11478 42443 11662
rect 42599 11536 42664 11737
rect 42599 11518 42621 11536
rect 42639 11518 42664 11536
rect 42599 11499 42664 11518
rect 42292 11474 42329 11475
rect 41715 11453 41751 11474
rect 42141 11453 42172 11474
rect 42379 11469 42387 11478
rect 42376 11453 42387 11469
rect 41548 11449 41648 11453
rect 41548 11445 41610 11449
rect 41548 11419 41555 11445
rect 41581 11423 41610 11445
rect 41636 11423 41648 11449
rect 41581 11419 41648 11423
rect 41548 11416 41648 11419
rect 41716 11416 41751 11453
rect 41813 11450 42172 11453
rect 41813 11445 42035 11450
rect 41813 11421 41826 11445
rect 41850 11426 42035 11445
rect 42059 11426 42172 11450
rect 41850 11421 42172 11426
rect 41813 11417 42172 11421
rect 42239 11445 42387 11453
rect 42239 11425 42250 11445
rect 42270 11436 42387 11445
rect 42436 11469 42443 11478
rect 42436 11436 42444 11469
rect 42270 11425 42444 11436
rect 42239 11418 42444 11425
rect 42239 11417 42280 11418
rect 41715 11391 41751 11416
rect 41563 11364 41600 11365
rect 41659 11364 41696 11365
rect 41715 11364 41722 11391
rect 41239 11339 41247 11359
rect 41267 11339 41276 11359
rect 41093 11328 41124 11329
rect 41088 11260 41198 11273
rect 41239 11260 41276 11339
rect 41463 11355 41601 11364
rect 41463 11335 41572 11355
rect 41592 11335 41601 11355
rect 41463 11328 41601 11335
rect 41659 11361 41722 11364
rect 41743 11364 41751 11391
rect 41770 11364 41807 11365
rect 41743 11361 41807 11364
rect 41659 11355 41807 11361
rect 41659 11335 41668 11355
rect 41688 11335 41778 11355
rect 41798 11335 41807 11355
rect 41463 11326 41559 11328
rect 41659 11325 41807 11335
rect 41866 11355 41903 11365
rect 41978 11364 42015 11365
rect 41959 11362 42015 11364
rect 41866 11335 41874 11355
rect 41894 11335 41903 11355
rect 41715 11324 41751 11325
rect 41026 11258 41276 11260
rect 41026 11255 41127 11258
rect 41026 11236 41091 11255
rect 41088 11228 41091 11236
rect 41120 11228 41127 11255
rect 41155 11231 41165 11258
rect 41194 11236 41276 11258
rect 41194 11231 41198 11236
rect 41155 11228 41198 11231
rect 41088 11214 41198 11228
rect 40514 11196 40855 11197
rect 40439 11191 40855 11196
rect 41563 11193 41600 11194
rect 41866 11193 41903 11335
rect 41928 11355 42015 11362
rect 41928 11352 41986 11355
rect 41928 11332 41933 11352
rect 41954 11335 41986 11352
rect 42006 11335 42015 11355
rect 41954 11332 42015 11335
rect 41928 11325 42015 11332
rect 42074 11355 42111 11365
rect 42074 11335 42082 11355
rect 42102 11335 42111 11355
rect 41928 11324 41959 11325
rect 42074 11256 42111 11335
rect 42141 11364 42172 11417
rect 42376 11415 42444 11418
rect 42376 11373 42388 11415
rect 42437 11373 42444 11415
rect 42191 11364 42228 11365
rect 42141 11355 42228 11364
rect 42141 11335 42199 11355
rect 42219 11335 42228 11355
rect 42141 11325 42228 11335
rect 42287 11355 42324 11365
rect 42376 11360 42444 11373
rect 42599 11437 42664 11454
rect 42599 11419 42623 11437
rect 42641 11419 42664 11437
rect 42287 11335 42295 11355
rect 42315 11335 42324 11355
rect 42141 11324 42172 11325
rect 42136 11256 42246 11269
rect 42287 11256 42324 11335
rect 42599 11280 42664 11419
rect 42599 11274 42621 11280
rect 42074 11254 42324 11256
rect 42074 11251 42175 11254
rect 42074 11232 42139 11251
rect 42136 11224 42139 11232
rect 42168 11224 42175 11251
rect 42203 11227 42213 11254
rect 42242 11232 42324 11254
rect 42353 11262 42621 11274
rect 42639 11262 42664 11280
rect 42353 11239 42664 11262
rect 42353 11238 42408 11239
rect 42242 11227 42246 11232
rect 42203 11224 42246 11227
rect 42136 11210 42246 11224
rect 41562 11192 41903 11193
rect 40439 11171 40442 11191
rect 40462 11171 40855 11191
rect 41487 11191 41903 11192
rect 42353 11191 42396 11238
rect 41487 11187 42396 11191
rect 40806 11138 40851 11171
rect 41487 11167 41490 11187
rect 41510 11167 42396 11187
rect 41864 11162 42396 11167
rect 42604 11181 42663 11203
rect 42604 11163 42623 11181
rect 42641 11163 42663 11181
rect 41652 11138 41751 11140
rect 40806 11128 41751 11138
rect 40806 11102 41674 11128
rect 40807 11101 41674 11102
rect 41652 11090 41674 11101
rect 41699 11093 41718 11128
rect 41743 11093 41751 11128
rect 41699 11090 41751 11093
rect 41652 11082 41751 11090
rect 41678 11081 41750 11082
rect 42604 11033 42663 11163
rect 41326 11003 41402 11027
rect 41326 10937 41338 11003
rect 41392 10937 41402 11003
rect 41870 10958 41911 10960
rect 42142 10958 42246 10960
rect 42604 10958 42665 11033
rect 40216 10887 40288 10937
rect 38927 10795 39371 10821
rect 38927 10793 39095 10795
rect 38927 10526 38954 10793
rect 39224 10791 39253 10795
rect 38994 10666 39058 10678
rect 39334 10674 39371 10795
rect 39599 10763 39710 10778
rect 39599 10761 39641 10763
rect 39599 10741 39606 10761
rect 39625 10741 39641 10761
rect 39599 10733 39641 10741
rect 39669 10761 39710 10763
rect 39669 10741 39683 10761
rect 39702 10741 39710 10761
rect 39669 10733 39710 10741
rect 39599 10727 39710 10733
rect 39542 10705 39791 10727
rect 39542 10674 39579 10705
rect 39755 10703 39791 10705
rect 39755 10674 39792 10703
rect 38994 10665 39029 10666
rect 38971 10660 39029 10665
rect 38971 10640 38974 10660
rect 38994 10646 39029 10660
rect 39049 10646 39058 10666
rect 38994 10638 39058 10646
rect 39020 10637 39058 10638
rect 39021 10636 39058 10637
rect 39124 10670 39160 10671
rect 39232 10670 39268 10671
rect 39124 10662 39268 10670
rect 39124 10642 39132 10662
rect 39152 10642 39240 10662
rect 39260 10642 39268 10662
rect 39124 10636 39268 10642
rect 39334 10666 39372 10674
rect 39440 10670 39476 10671
rect 39334 10646 39343 10666
rect 39363 10646 39372 10666
rect 39334 10637 39372 10646
rect 39391 10663 39476 10670
rect 39391 10643 39398 10663
rect 39419 10662 39476 10663
rect 39419 10643 39448 10662
rect 39391 10642 39448 10643
rect 39468 10642 39476 10662
rect 39334 10636 39371 10637
rect 39391 10636 39476 10642
rect 39542 10666 39580 10674
rect 39653 10670 39689 10671
rect 39542 10646 39551 10666
rect 39571 10646 39580 10666
rect 39542 10637 39580 10646
rect 39604 10662 39689 10670
rect 39604 10642 39661 10662
rect 39681 10642 39689 10662
rect 39542 10636 39579 10637
rect 39604 10636 39689 10642
rect 39755 10666 39793 10674
rect 39755 10646 39764 10666
rect 39784 10646 39793 10666
rect 39755 10637 39793 10646
rect 39755 10636 39792 10637
rect 39178 10615 39214 10636
rect 39604 10615 39635 10636
rect 39785 10615 40119 10619
rect 39011 10611 39111 10615
rect 39011 10607 39073 10611
rect 39011 10581 39018 10607
rect 39044 10585 39073 10607
rect 39099 10585 39111 10611
rect 39044 10581 39111 10585
rect 39011 10578 39111 10581
rect 39179 10578 39214 10615
rect 39276 10612 39635 10615
rect 39276 10607 39498 10612
rect 39276 10583 39289 10607
rect 39313 10588 39498 10607
rect 39522 10588 39635 10612
rect 39313 10583 39635 10588
rect 39276 10579 39635 10583
rect 39702 10607 40119 10615
rect 39702 10587 39713 10607
rect 39733 10587 40119 10607
rect 39702 10580 40119 10587
rect 39702 10579 39743 10580
rect 39785 10579 40119 10580
rect 39178 10553 39214 10578
rect 39026 10526 39063 10527
rect 39122 10526 39159 10527
rect 39178 10526 39185 10553
rect 38926 10517 39064 10526
rect 38926 10497 39035 10517
rect 39055 10497 39064 10517
rect 38926 10490 39064 10497
rect 39122 10523 39185 10526
rect 39206 10526 39214 10553
rect 39233 10526 39270 10527
rect 39206 10523 39270 10526
rect 39122 10517 39270 10523
rect 39122 10497 39131 10517
rect 39151 10497 39241 10517
rect 39261 10497 39270 10517
rect 38926 10488 39022 10490
rect 39122 10487 39270 10497
rect 39329 10517 39366 10527
rect 39441 10526 39478 10527
rect 39422 10524 39478 10526
rect 39329 10497 39337 10517
rect 39357 10497 39366 10517
rect 39178 10486 39214 10487
rect 39026 10355 39063 10356
rect 39329 10355 39366 10497
rect 39391 10517 39478 10524
rect 39391 10514 39449 10517
rect 39391 10494 39396 10514
rect 39417 10497 39449 10514
rect 39469 10497 39478 10517
rect 39417 10494 39478 10497
rect 39391 10487 39478 10494
rect 39537 10517 39574 10527
rect 39537 10497 39545 10517
rect 39565 10497 39574 10517
rect 39391 10486 39422 10487
rect 39537 10418 39574 10497
rect 39604 10526 39635 10579
rect 39654 10526 39691 10527
rect 39604 10517 39691 10526
rect 39604 10497 39662 10517
rect 39682 10497 39691 10517
rect 39604 10487 39691 10497
rect 39750 10517 39787 10527
rect 39750 10497 39758 10517
rect 39778 10497 39787 10517
rect 39604 10486 39635 10487
rect 39599 10418 39709 10431
rect 39750 10418 39787 10497
rect 39537 10416 39787 10418
rect 39537 10413 39638 10416
rect 39537 10394 39602 10413
rect 39599 10386 39602 10394
rect 39631 10386 39638 10413
rect 39666 10389 39676 10416
rect 39705 10394 39787 10416
rect 39705 10389 39709 10394
rect 39666 10386 39709 10389
rect 39599 10372 39709 10386
rect 39025 10354 39366 10355
rect 38950 10349 39366 10354
rect 38950 10329 38953 10349
rect 38973 10329 39366 10349
rect 39259 9964 39290 10329
rect 39177 9935 39290 9964
rect 39178 9635 39214 9935
rect 40038 9830 40119 10579
rect 40218 9978 40288 10887
rect 41326 10917 41402 10937
rect 41326 10880 41343 10917
rect 41387 10880 41402 10917
rect 41463 10923 42665 10958
rect 41463 10909 41491 10923
rect 41326 10864 41402 10880
rect 41331 10708 41401 10864
rect 41465 10778 41491 10909
rect 41870 10920 42665 10923
rect 41323 10657 41403 10708
rect 41323 10631 41339 10657
rect 41379 10631 41403 10657
rect 41323 10612 41403 10631
rect 41323 10586 41342 10612
rect 41382 10586 41403 10612
rect 41323 10559 41403 10586
rect 41323 10533 41346 10559
rect 41386 10533 41403 10559
rect 41323 10522 41403 10533
rect 41465 10523 41492 10778
rect 41870 10770 41911 10920
rect 42604 10908 42665 10920
rect 42337 10858 42458 10876
rect 42337 10856 42408 10858
rect 42337 10815 42352 10856
rect 42389 10817 42408 10856
rect 42445 10817 42458 10858
rect 42389 10815 42458 10817
rect 42337 10805 42458 10815
rect 42142 10775 42246 10784
rect 41532 10663 41596 10675
rect 41872 10671 41909 10770
rect 42137 10760 42248 10775
rect 42137 10758 42179 10760
rect 42137 10738 42144 10758
rect 42163 10738 42179 10758
rect 42137 10730 42179 10738
rect 42207 10758 42248 10760
rect 42207 10738 42221 10758
rect 42240 10738 42248 10758
rect 42207 10730 42248 10738
rect 42137 10724 42248 10730
rect 42080 10702 42329 10724
rect 42080 10671 42117 10702
rect 42293 10700 42329 10702
rect 42293 10671 42330 10700
rect 41532 10662 41567 10663
rect 41509 10657 41567 10662
rect 41509 10637 41512 10657
rect 41532 10643 41567 10657
rect 41587 10643 41596 10663
rect 41532 10635 41596 10643
rect 41558 10634 41596 10635
rect 41559 10633 41596 10634
rect 41662 10667 41698 10668
rect 41770 10667 41806 10668
rect 41662 10659 41806 10667
rect 41662 10639 41670 10659
rect 41690 10639 41778 10659
rect 41798 10639 41806 10659
rect 41662 10633 41806 10639
rect 41872 10663 41910 10671
rect 41978 10667 42014 10668
rect 41872 10643 41881 10663
rect 41901 10643 41910 10663
rect 41872 10634 41910 10643
rect 41929 10660 42014 10667
rect 41929 10640 41936 10660
rect 41957 10659 42014 10660
rect 41957 10640 41986 10659
rect 41929 10639 41986 10640
rect 42006 10639 42014 10659
rect 41872 10633 41909 10634
rect 41929 10633 42014 10639
rect 42080 10663 42118 10671
rect 42191 10667 42227 10668
rect 42080 10643 42089 10663
rect 42109 10643 42118 10663
rect 42080 10634 42118 10643
rect 42142 10659 42227 10667
rect 42142 10639 42199 10659
rect 42219 10639 42227 10659
rect 42080 10633 42117 10634
rect 42142 10633 42227 10639
rect 42293 10663 42331 10671
rect 42293 10643 42302 10663
rect 42322 10643 42331 10663
rect 42386 10653 42451 10805
rect 42604 10779 42659 10908
rect 42293 10634 42331 10643
rect 42384 10646 42451 10653
rect 42293 10633 42330 10634
rect 41716 10612 41752 10633
rect 42142 10612 42173 10633
rect 42384 10625 42401 10646
rect 42437 10625 42451 10646
rect 42603 10666 42659 10779
rect 42603 10648 42622 10666
rect 42640 10648 42659 10666
rect 42603 10628 42659 10648
rect 42384 10612 42451 10625
rect 41549 10608 41649 10612
rect 41549 10604 41611 10608
rect 41549 10578 41556 10604
rect 41582 10582 41611 10604
rect 41637 10582 41649 10608
rect 41582 10578 41649 10582
rect 41549 10575 41649 10578
rect 41717 10575 41752 10612
rect 41814 10609 42173 10612
rect 41814 10604 42036 10609
rect 41814 10580 41827 10604
rect 41851 10585 42036 10604
rect 42060 10585 42173 10609
rect 41851 10580 42173 10585
rect 41814 10576 42173 10580
rect 42240 10606 42451 10612
rect 42240 10604 42401 10606
rect 42240 10584 42251 10604
rect 42271 10584 42401 10604
rect 42240 10577 42401 10584
rect 42240 10576 42281 10577
rect 41716 10550 41752 10575
rect 41564 10523 41601 10524
rect 41660 10523 41697 10524
rect 41716 10523 41723 10550
rect 41464 10514 41602 10523
rect 41464 10494 41573 10514
rect 41593 10494 41602 10514
rect 41464 10487 41602 10494
rect 41660 10520 41723 10523
rect 41744 10523 41752 10550
rect 41771 10523 41808 10524
rect 41744 10520 41808 10523
rect 41660 10514 41808 10520
rect 41660 10494 41669 10514
rect 41689 10494 41779 10514
rect 41799 10494 41808 10514
rect 41464 10485 41560 10487
rect 41660 10484 41808 10494
rect 41867 10514 41904 10524
rect 41979 10523 42016 10524
rect 41960 10521 42016 10523
rect 41867 10494 41875 10514
rect 41895 10494 41904 10514
rect 41716 10483 41752 10484
rect 41564 10352 41601 10353
rect 41867 10352 41904 10494
rect 41929 10514 42016 10521
rect 41929 10511 41987 10514
rect 41929 10491 41934 10511
rect 41955 10494 41987 10511
rect 42007 10494 42016 10514
rect 41955 10491 42016 10494
rect 41929 10484 42016 10491
rect 42075 10514 42112 10524
rect 42075 10494 42083 10514
rect 42103 10494 42112 10514
rect 41929 10483 41960 10484
rect 42075 10415 42112 10494
rect 42142 10523 42173 10576
rect 42386 10569 42401 10577
rect 42441 10569 42451 10606
rect 42386 10560 42451 10569
rect 42599 10567 42664 10588
rect 42599 10549 42624 10567
rect 42642 10549 42664 10567
rect 42192 10523 42229 10524
rect 42142 10514 42229 10523
rect 42142 10494 42200 10514
rect 42220 10494 42229 10514
rect 42142 10484 42229 10494
rect 42288 10514 42325 10524
rect 42288 10494 42296 10514
rect 42316 10494 42325 10514
rect 42142 10483 42173 10484
rect 42137 10415 42247 10428
rect 42288 10415 42325 10494
rect 42599 10473 42664 10549
rect 42075 10413 42325 10415
rect 42075 10410 42176 10413
rect 42075 10391 42140 10410
rect 42137 10383 42140 10391
rect 42169 10383 42176 10410
rect 42204 10386 42214 10413
rect 42243 10391 42325 10413
rect 42348 10438 42665 10473
rect 42243 10386 42247 10391
rect 42204 10383 42247 10386
rect 42137 10369 42247 10383
rect 41563 10351 41904 10352
rect 41488 10349 41904 10351
rect 42348 10349 42388 10438
rect 42599 10411 42664 10438
rect 42599 10393 42622 10411
rect 42640 10393 42664 10411
rect 42599 10373 42664 10393
rect 41485 10346 42388 10349
rect 41485 10326 41491 10346
rect 41511 10326 42388 10346
rect 41485 10322 42388 10326
rect 42348 10319 42388 10322
rect 42600 10312 42665 10333
rect 40818 10304 41479 10305
rect 40818 10297 41752 10304
rect 40818 10296 41724 10297
rect 40818 10276 41669 10296
rect 41701 10277 41724 10296
rect 41749 10277 41752 10297
rect 41701 10276 41752 10277
rect 40818 10269 41752 10276
rect 40417 10227 40585 10228
rect 40820 10227 40859 10269
rect 41648 10267 41752 10269
rect 41717 10265 41752 10267
rect 42600 10294 42624 10312
rect 42642 10294 42665 10312
rect 42600 10247 42665 10294
rect 40417 10201 40861 10227
rect 40417 10199 40585 10201
rect 39178 9612 39182 9635
rect 39206 9612 39214 9635
rect 39378 9613 39477 9617
rect 39178 9591 39214 9612
rect 39178 9568 39182 9591
rect 39206 9568 39214 9591
rect 39178 9564 39214 9568
rect 39374 9607 39477 9613
rect 39374 9569 39400 9607
rect 39425 9572 39444 9607
rect 39469 9572 39477 9607
rect 39425 9569 39477 9572
rect 39374 9561 39477 9569
rect 39374 9560 39476 9561
rect 38970 9482 39138 9483
rect 39374 9482 39421 9560
rect 38970 9456 39421 9482
rect 38970 9454 39138 9456
rect 38970 9081 38997 9454
rect 39167 9406 39253 9415
rect 39167 9388 39186 9406
rect 39238 9388 39253 9406
rect 39167 9384 39253 9388
rect 39037 9221 39101 9233
rect 39037 9220 39072 9221
rect 39014 9215 39072 9220
rect 39014 9195 39017 9215
rect 39037 9201 39072 9215
rect 39092 9201 39101 9221
rect 39037 9193 39101 9201
rect 39063 9192 39101 9193
rect 39064 9191 39101 9192
rect 39167 9225 39203 9226
rect 39223 9225 39253 9384
rect 39374 9344 39421 9456
rect 39377 9229 39414 9344
rect 39642 9318 39753 9333
rect 39642 9316 39684 9318
rect 39642 9296 39649 9316
rect 39668 9296 39684 9316
rect 39642 9288 39684 9296
rect 39712 9316 39753 9318
rect 39712 9296 39726 9316
rect 39745 9296 39753 9316
rect 39712 9288 39753 9296
rect 39642 9282 39753 9288
rect 39585 9260 39834 9282
rect 39585 9229 39622 9260
rect 39798 9258 39834 9260
rect 39798 9229 39835 9258
rect 40039 9245 40118 9830
rect 40215 9378 40294 9978
rect 40417 9848 40444 10199
rect 40820 10195 40861 10201
rect 40484 9988 40548 10000
rect 40824 9996 40861 10195
rect 41323 10222 41395 10239
rect 41323 10183 41331 10222
rect 41376 10183 41395 10222
rect 41089 10085 41200 10100
rect 41089 10083 41131 10085
rect 41089 10063 41096 10083
rect 41115 10063 41131 10083
rect 41089 10055 41131 10063
rect 41159 10083 41200 10085
rect 41159 10063 41173 10083
rect 41192 10063 41200 10083
rect 41159 10055 41200 10063
rect 41089 10049 41200 10055
rect 41032 10027 41281 10049
rect 41032 9996 41069 10027
rect 41245 10025 41281 10027
rect 41245 9996 41282 10025
rect 40484 9987 40519 9988
rect 40461 9982 40519 9987
rect 40461 9962 40464 9982
rect 40484 9968 40519 9982
rect 40539 9968 40548 9988
rect 40484 9960 40548 9968
rect 40510 9959 40548 9960
rect 40511 9958 40548 9959
rect 40614 9992 40650 9993
rect 40722 9992 40758 9993
rect 40614 9984 40758 9992
rect 40614 9964 40622 9984
rect 40642 9964 40730 9984
rect 40750 9964 40758 9984
rect 40614 9958 40758 9964
rect 40824 9988 40862 9996
rect 40930 9992 40966 9993
rect 40824 9968 40833 9988
rect 40853 9968 40862 9988
rect 40824 9959 40862 9968
rect 40881 9985 40966 9992
rect 40881 9965 40888 9985
rect 40909 9984 40966 9985
rect 40909 9965 40938 9984
rect 40881 9964 40938 9965
rect 40958 9964 40966 9984
rect 40824 9958 40861 9959
rect 40881 9958 40966 9964
rect 41032 9988 41070 9996
rect 41143 9992 41179 9993
rect 41032 9968 41041 9988
rect 41061 9968 41070 9988
rect 41032 9959 41070 9968
rect 41094 9984 41179 9992
rect 41094 9964 41151 9984
rect 41171 9964 41179 9984
rect 41032 9958 41069 9959
rect 41094 9958 41179 9964
rect 41245 9988 41283 9996
rect 41245 9968 41254 9988
rect 41274 9968 41283 9988
rect 41245 9959 41283 9968
rect 41323 9973 41395 10183
rect 41465 10217 42665 10247
rect 41465 10216 41909 10217
rect 41465 10214 41633 10216
rect 41323 9959 41406 9973
rect 41245 9958 41282 9959
rect 40668 9937 40704 9958
rect 41094 9937 41125 9958
rect 41323 9937 41340 9959
rect 40501 9933 40601 9937
rect 40501 9929 40563 9933
rect 40501 9903 40508 9929
rect 40534 9907 40563 9929
rect 40589 9907 40601 9933
rect 40534 9903 40601 9907
rect 40501 9900 40601 9903
rect 40669 9900 40704 9937
rect 40766 9934 41125 9937
rect 40766 9929 40988 9934
rect 40766 9905 40779 9929
rect 40803 9910 40988 9929
rect 41012 9910 41125 9934
rect 40803 9905 41125 9910
rect 40766 9901 41125 9905
rect 41192 9929 41340 9937
rect 41192 9909 41203 9929
rect 41223 9926 41340 9929
rect 41393 9926 41406 9959
rect 41223 9909 41406 9926
rect 41192 9902 41406 9909
rect 41192 9901 41233 9902
rect 41323 9901 41406 9902
rect 40668 9875 40704 9900
rect 40516 9848 40553 9849
rect 40612 9848 40649 9849
rect 40668 9848 40675 9875
rect 40416 9839 40554 9848
rect 40416 9819 40525 9839
rect 40545 9819 40554 9839
rect 40416 9812 40554 9819
rect 40612 9845 40675 9848
rect 40696 9848 40704 9875
rect 40723 9848 40760 9849
rect 40696 9845 40760 9848
rect 40612 9839 40760 9845
rect 40612 9819 40621 9839
rect 40641 9819 40731 9839
rect 40751 9819 40760 9839
rect 40416 9810 40512 9812
rect 40612 9809 40760 9819
rect 40819 9839 40856 9849
rect 40931 9848 40968 9849
rect 40912 9846 40968 9848
rect 40819 9819 40827 9839
rect 40847 9819 40856 9839
rect 40668 9808 40704 9809
rect 40516 9677 40553 9678
rect 40819 9677 40856 9819
rect 40881 9839 40968 9846
rect 40881 9836 40939 9839
rect 40881 9816 40886 9836
rect 40907 9819 40939 9836
rect 40959 9819 40968 9839
rect 40907 9816 40968 9819
rect 40881 9809 40968 9816
rect 41027 9839 41064 9849
rect 41027 9819 41035 9839
rect 41055 9819 41064 9839
rect 40881 9808 40912 9809
rect 41027 9740 41064 9819
rect 41094 9848 41125 9901
rect 41331 9868 41345 9901
rect 41398 9868 41406 9901
rect 41331 9862 41406 9868
rect 41331 9857 41401 9862
rect 41144 9848 41181 9849
rect 41094 9839 41181 9848
rect 41094 9819 41152 9839
rect 41172 9819 41181 9839
rect 41094 9809 41181 9819
rect 41240 9839 41277 9849
rect 41465 9844 41492 10214
rect 41532 9984 41596 9996
rect 41872 9992 41909 10216
rect 42380 10197 42444 10199
rect 42376 10185 42444 10197
rect 42376 10152 42387 10185
rect 42427 10152 42444 10185
rect 42376 10142 42444 10152
rect 42137 10081 42248 10096
rect 42137 10079 42179 10081
rect 42137 10059 42144 10079
rect 42163 10059 42179 10079
rect 42137 10051 42179 10059
rect 42207 10079 42248 10081
rect 42207 10059 42221 10079
rect 42240 10059 42248 10079
rect 42207 10051 42248 10059
rect 42137 10045 42248 10051
rect 42080 10023 42329 10045
rect 42080 9992 42117 10023
rect 42293 10021 42329 10023
rect 42293 9992 42330 10021
rect 41532 9983 41567 9984
rect 41509 9978 41567 9983
rect 41509 9958 41512 9978
rect 41532 9964 41567 9978
rect 41587 9964 41596 9984
rect 41532 9956 41596 9964
rect 41558 9955 41596 9956
rect 41559 9954 41596 9955
rect 41662 9988 41698 9989
rect 41770 9988 41806 9989
rect 41662 9980 41806 9988
rect 41662 9960 41670 9980
rect 41690 9960 41778 9980
rect 41798 9960 41806 9980
rect 41662 9954 41806 9960
rect 41872 9984 41910 9992
rect 41978 9988 42014 9989
rect 41872 9964 41881 9984
rect 41901 9964 41910 9984
rect 41872 9955 41910 9964
rect 41929 9981 42014 9988
rect 41929 9961 41936 9981
rect 41957 9980 42014 9981
rect 41957 9961 41986 9980
rect 41929 9960 41986 9961
rect 42006 9960 42014 9980
rect 41872 9954 41909 9955
rect 41929 9954 42014 9960
rect 42080 9984 42118 9992
rect 42191 9988 42227 9989
rect 42080 9964 42089 9984
rect 42109 9964 42118 9984
rect 42080 9955 42118 9964
rect 42142 9980 42227 9988
rect 42142 9960 42199 9980
rect 42219 9960 42227 9980
rect 42080 9954 42117 9955
rect 42142 9954 42227 9960
rect 42293 9984 42331 9992
rect 42293 9964 42302 9984
rect 42322 9964 42331 9984
rect 42293 9955 42331 9964
rect 42380 9958 42444 10142
rect 42600 10016 42665 10217
rect 42600 9998 42622 10016
rect 42640 9998 42665 10016
rect 42600 9979 42665 9998
rect 42293 9954 42330 9955
rect 41716 9933 41752 9954
rect 42142 9933 42173 9954
rect 42380 9949 42388 9958
rect 42377 9933 42388 9949
rect 41549 9929 41649 9933
rect 41549 9925 41611 9929
rect 41549 9899 41556 9925
rect 41582 9903 41611 9925
rect 41637 9903 41649 9929
rect 41582 9899 41649 9903
rect 41549 9896 41649 9899
rect 41717 9896 41752 9933
rect 41814 9930 42173 9933
rect 41814 9925 42036 9930
rect 41814 9901 41827 9925
rect 41851 9906 42036 9925
rect 42060 9906 42173 9930
rect 41851 9901 42173 9906
rect 41814 9897 42173 9901
rect 42240 9925 42388 9933
rect 42240 9905 42251 9925
rect 42271 9916 42388 9925
rect 42437 9949 42444 9958
rect 42437 9916 42445 9949
rect 42271 9905 42445 9916
rect 42240 9898 42445 9905
rect 42240 9897 42281 9898
rect 41716 9871 41752 9896
rect 41564 9844 41601 9845
rect 41660 9844 41697 9845
rect 41716 9844 41723 9871
rect 41240 9819 41248 9839
rect 41268 9819 41277 9839
rect 41094 9808 41125 9809
rect 41089 9740 41199 9753
rect 41240 9740 41277 9819
rect 41464 9835 41602 9844
rect 41464 9815 41573 9835
rect 41593 9815 41602 9835
rect 41464 9808 41602 9815
rect 41660 9841 41723 9844
rect 41744 9844 41752 9871
rect 41771 9844 41808 9845
rect 41744 9841 41808 9844
rect 41660 9835 41808 9841
rect 41660 9815 41669 9835
rect 41689 9815 41779 9835
rect 41799 9815 41808 9835
rect 41464 9806 41560 9808
rect 41660 9805 41808 9815
rect 41867 9835 41904 9845
rect 41979 9844 42016 9845
rect 41960 9842 42016 9844
rect 41867 9815 41875 9835
rect 41895 9815 41904 9835
rect 41716 9804 41752 9805
rect 41027 9738 41277 9740
rect 41027 9735 41128 9738
rect 41027 9716 41092 9735
rect 41089 9708 41092 9716
rect 41121 9708 41128 9735
rect 41156 9711 41166 9738
rect 41195 9716 41277 9738
rect 41195 9711 41199 9716
rect 41156 9708 41199 9711
rect 41089 9694 41199 9708
rect 40515 9676 40856 9677
rect 40440 9671 40856 9676
rect 41564 9673 41601 9674
rect 41867 9673 41904 9815
rect 41929 9835 42016 9842
rect 41929 9832 41987 9835
rect 41929 9812 41934 9832
rect 41955 9815 41987 9832
rect 42007 9815 42016 9835
rect 41955 9812 42016 9815
rect 41929 9805 42016 9812
rect 42075 9835 42112 9845
rect 42075 9815 42083 9835
rect 42103 9815 42112 9835
rect 41929 9804 41960 9805
rect 42075 9736 42112 9815
rect 42142 9844 42173 9897
rect 42377 9895 42445 9898
rect 42377 9853 42389 9895
rect 42438 9853 42445 9895
rect 42192 9844 42229 9845
rect 42142 9835 42229 9844
rect 42142 9815 42200 9835
rect 42220 9815 42229 9835
rect 42142 9805 42229 9815
rect 42288 9835 42325 9845
rect 42377 9840 42445 9853
rect 42600 9917 42665 9934
rect 42600 9899 42624 9917
rect 42642 9899 42665 9917
rect 42288 9815 42296 9835
rect 42316 9815 42325 9835
rect 42142 9804 42173 9805
rect 42137 9736 42247 9749
rect 42288 9736 42325 9815
rect 42600 9760 42665 9899
rect 42600 9754 42622 9760
rect 42075 9734 42325 9736
rect 42075 9731 42176 9734
rect 42075 9712 42140 9731
rect 42137 9704 42140 9712
rect 42169 9704 42176 9731
rect 42204 9707 42214 9734
rect 42243 9712 42325 9734
rect 42354 9742 42622 9754
rect 42640 9742 42665 9760
rect 42354 9719 42665 9742
rect 42354 9718 42409 9719
rect 42243 9707 42247 9712
rect 42204 9704 42247 9707
rect 42137 9690 42247 9704
rect 41563 9672 41904 9673
rect 40440 9651 40443 9671
rect 40463 9651 40856 9671
rect 41488 9671 41904 9672
rect 42354 9671 42397 9718
rect 41488 9667 42397 9671
rect 40807 9618 40852 9651
rect 41488 9647 41491 9667
rect 41511 9647 42397 9667
rect 41865 9642 42397 9647
rect 42605 9661 42664 9683
rect 42605 9643 42624 9661
rect 42642 9643 42664 9661
rect 41653 9618 41752 9620
rect 40807 9608 41752 9618
rect 40807 9582 41675 9608
rect 40808 9581 41675 9582
rect 41653 9570 41675 9581
rect 41700 9573 41719 9608
rect 41744 9573 41752 9608
rect 41700 9570 41752 9573
rect 42605 9572 42664 9643
rect 41653 9562 41752 9570
rect 41679 9561 41751 9562
rect 41333 9535 41400 9554
rect 41333 9514 41350 9535
rect 40214 9336 40294 9378
rect 41331 9469 41350 9514
rect 41380 9514 41400 9535
rect 41380 9469 41401 9514
rect 41870 9511 41911 9513
rect 42142 9511 42246 9513
rect 42602 9511 42666 9572
rect 39275 9225 39311 9226
rect 39167 9217 39311 9225
rect 39167 9197 39175 9217
rect 39195 9197 39283 9217
rect 39303 9197 39311 9217
rect 39167 9191 39311 9197
rect 39377 9221 39415 9229
rect 39483 9225 39519 9226
rect 39377 9201 39386 9221
rect 39406 9201 39415 9221
rect 39377 9192 39415 9201
rect 39434 9218 39519 9225
rect 39434 9198 39441 9218
rect 39462 9217 39519 9218
rect 39462 9198 39491 9217
rect 39434 9197 39491 9198
rect 39511 9197 39519 9217
rect 39377 9191 39414 9192
rect 39434 9191 39519 9197
rect 39585 9221 39623 9229
rect 39696 9225 39732 9226
rect 39585 9201 39594 9221
rect 39614 9201 39623 9221
rect 39585 9192 39623 9201
rect 39647 9217 39732 9225
rect 39647 9197 39704 9217
rect 39724 9197 39732 9217
rect 39585 9191 39622 9192
rect 39647 9191 39732 9197
rect 39798 9221 39836 9229
rect 39798 9201 39807 9221
rect 39827 9201 39836 9221
rect 39798 9192 39836 9201
rect 40036 9209 40122 9245
rect 39798 9191 39835 9192
rect 39221 9170 39257 9191
rect 39647 9170 39678 9191
rect 39874 9170 39920 9174
rect 39054 9166 39154 9170
rect 39054 9162 39116 9166
rect 39054 9136 39061 9162
rect 39087 9140 39116 9162
rect 39142 9140 39154 9166
rect 39087 9136 39154 9140
rect 39054 9133 39154 9136
rect 39222 9133 39257 9170
rect 39319 9167 39678 9170
rect 39319 9162 39541 9167
rect 39319 9138 39332 9162
rect 39356 9143 39541 9162
rect 39565 9143 39678 9167
rect 39356 9138 39678 9143
rect 39319 9134 39678 9138
rect 39745 9162 39920 9170
rect 39745 9142 39756 9162
rect 39776 9142 39920 9162
rect 40036 9168 40053 9209
rect 40107 9168 40122 9209
rect 40036 9149 40122 9168
rect 39745 9135 39920 9142
rect 39745 9134 39786 9135
rect 39221 9108 39257 9133
rect 39069 9081 39106 9082
rect 39165 9081 39202 9082
rect 39221 9081 39228 9108
rect 38969 9072 39107 9081
rect 38969 9052 39078 9072
rect 39098 9052 39107 9072
rect 38969 9045 39107 9052
rect 39165 9078 39228 9081
rect 39249 9081 39257 9108
rect 39276 9081 39313 9082
rect 39249 9078 39313 9081
rect 39165 9072 39313 9078
rect 39165 9052 39174 9072
rect 39194 9052 39284 9072
rect 39304 9052 39313 9072
rect 38969 9043 39065 9045
rect 39165 9042 39313 9052
rect 39372 9072 39409 9082
rect 39484 9081 39521 9082
rect 39465 9079 39521 9081
rect 39372 9052 39380 9072
rect 39400 9052 39409 9072
rect 39221 9041 39257 9042
rect 39069 8910 39106 8911
rect 39372 8910 39409 9052
rect 39434 9072 39521 9079
rect 39434 9069 39492 9072
rect 39434 9049 39439 9069
rect 39460 9052 39492 9069
rect 39512 9052 39521 9072
rect 39460 9049 39521 9052
rect 39434 9042 39521 9049
rect 39580 9072 39617 9082
rect 39580 9052 39588 9072
rect 39608 9052 39617 9072
rect 39434 9041 39465 9042
rect 39580 8973 39617 9052
rect 39647 9081 39678 9134
rect 39697 9081 39734 9082
rect 39647 9072 39734 9081
rect 39647 9052 39705 9072
rect 39725 9052 39734 9072
rect 39647 9042 39734 9052
rect 39793 9072 39830 9082
rect 39793 9052 39801 9072
rect 39821 9052 39830 9072
rect 39647 9041 39678 9042
rect 39642 8973 39752 8986
rect 39793 8973 39830 9052
rect 39874 9052 39920 9135
rect 40214 9052 40289 9336
rect 41331 9261 41401 9469
rect 41463 9476 42666 9511
rect 41463 9462 41491 9476
rect 41465 9331 41491 9462
rect 41870 9473 42666 9476
rect 41323 9210 41403 9261
rect 41323 9184 41339 9210
rect 41379 9184 41403 9210
rect 41323 9165 41403 9184
rect 41323 9139 41342 9165
rect 41382 9139 41403 9165
rect 41323 9112 41403 9139
rect 41323 9086 41346 9112
rect 41386 9086 41403 9112
rect 41323 9075 41403 9086
rect 41465 9076 41492 9331
rect 41870 9323 41911 9473
rect 42142 9467 42246 9473
rect 42602 9470 42666 9473
rect 42337 9411 42458 9429
rect 42337 9409 42408 9411
rect 42337 9368 42352 9409
rect 42389 9370 42408 9409
rect 42445 9370 42458 9411
rect 42389 9368 42458 9370
rect 42337 9358 42458 9368
rect 41532 9216 41596 9228
rect 41872 9224 41909 9323
rect 42137 9313 42248 9326
rect 42137 9311 42179 9313
rect 42137 9291 42144 9311
rect 42163 9291 42179 9311
rect 42137 9283 42179 9291
rect 42207 9311 42248 9313
rect 42207 9291 42221 9311
rect 42240 9291 42248 9311
rect 42207 9283 42248 9291
rect 42137 9277 42248 9283
rect 42080 9255 42329 9277
rect 42080 9224 42117 9255
rect 42293 9253 42329 9255
rect 42293 9224 42330 9253
rect 41532 9215 41567 9216
rect 41509 9210 41567 9215
rect 41509 9190 41512 9210
rect 41532 9196 41567 9210
rect 41587 9196 41596 9216
rect 41532 9188 41596 9196
rect 41558 9187 41596 9188
rect 41559 9186 41596 9187
rect 41662 9220 41698 9221
rect 41770 9220 41806 9221
rect 41662 9212 41806 9220
rect 41662 9192 41670 9212
rect 41690 9192 41778 9212
rect 41798 9192 41806 9212
rect 41662 9186 41806 9192
rect 41872 9216 41910 9224
rect 41978 9220 42014 9221
rect 41872 9196 41881 9216
rect 41901 9196 41910 9216
rect 41872 9187 41910 9196
rect 41929 9213 42014 9220
rect 41929 9193 41936 9213
rect 41957 9212 42014 9213
rect 41957 9193 41986 9212
rect 41929 9192 41986 9193
rect 42006 9192 42014 9212
rect 41872 9186 41909 9187
rect 41929 9186 42014 9192
rect 42080 9216 42118 9224
rect 42191 9220 42227 9221
rect 42080 9196 42089 9216
rect 42109 9196 42118 9216
rect 42080 9187 42118 9196
rect 42142 9212 42227 9220
rect 42142 9192 42199 9212
rect 42219 9192 42227 9212
rect 42080 9186 42117 9187
rect 42142 9186 42227 9192
rect 42293 9216 42331 9224
rect 42293 9196 42302 9216
rect 42322 9196 42331 9216
rect 42386 9206 42451 9358
rect 42604 9332 42659 9470
rect 42293 9187 42331 9196
rect 42384 9199 42451 9206
rect 42293 9186 42330 9187
rect 41716 9165 41752 9186
rect 42142 9165 42173 9186
rect 42384 9178 42401 9199
rect 42437 9178 42451 9199
rect 42603 9219 42659 9332
rect 42603 9201 42622 9219
rect 42640 9201 42659 9219
rect 42603 9181 42659 9201
rect 42384 9165 42451 9178
rect 41549 9161 41649 9165
rect 41549 9157 41611 9161
rect 41549 9131 41556 9157
rect 41582 9135 41611 9157
rect 41637 9135 41649 9161
rect 41582 9131 41649 9135
rect 41549 9128 41649 9131
rect 41717 9128 41752 9165
rect 41814 9162 42173 9165
rect 41814 9157 42036 9162
rect 41814 9133 41827 9157
rect 41851 9138 42036 9157
rect 42060 9138 42173 9162
rect 41851 9133 42173 9138
rect 41814 9129 42173 9133
rect 42240 9159 42451 9165
rect 42240 9157 42401 9159
rect 42240 9137 42251 9157
rect 42271 9137 42401 9157
rect 42240 9130 42401 9137
rect 42240 9129 42281 9130
rect 41716 9103 41752 9128
rect 41564 9076 41601 9077
rect 41660 9076 41697 9077
rect 41716 9076 41723 9103
rect 39874 9017 40289 9052
rect 41464 9067 41602 9076
rect 41464 9047 41573 9067
rect 41593 9047 41602 9067
rect 41464 9040 41602 9047
rect 41660 9073 41723 9076
rect 41744 9076 41752 9103
rect 41771 9076 41808 9077
rect 41744 9073 41808 9076
rect 41660 9067 41808 9073
rect 41660 9047 41669 9067
rect 41689 9047 41779 9067
rect 41799 9047 41808 9067
rect 41464 9038 41560 9040
rect 41660 9037 41808 9047
rect 41867 9067 41904 9077
rect 41979 9076 42016 9077
rect 41960 9074 42016 9076
rect 41867 9047 41875 9067
rect 41895 9047 41904 9067
rect 41716 9036 41752 9037
rect 39874 9016 39920 9017
rect 39580 8971 39830 8973
rect 39580 8968 39681 8971
rect 39580 8949 39645 8968
rect 39642 8941 39645 8949
rect 39674 8941 39681 8968
rect 39709 8944 39719 8971
rect 39748 8949 39830 8971
rect 40214 8965 40289 9017
rect 39748 8944 39752 8949
rect 39709 8941 39752 8944
rect 39642 8927 39752 8941
rect 39068 8909 39409 8910
rect 38993 8904 39409 8909
rect 38993 8884 38996 8904
rect 39016 8884 39410 8904
rect 38050 8237 38856 8312
rect 37289 8193 37298 8227
rect 37327 8226 37737 8227
rect 37327 8193 37344 8226
rect 37569 8225 37737 8226
rect 37289 8167 37344 8193
rect 37289 8133 37297 8167
rect 37326 8133 37344 8167
rect 37289 8121 37344 8133
rect 35485 8076 35569 8097
rect 35485 8048 35513 8076
rect 35557 8048 35569 8076
rect 35299 7997 35373 8025
rect 35299 7949 35322 7997
rect 35359 7949 35373 7997
rect 35485 8019 35569 8048
rect 35485 7991 35510 8019
rect 35554 7991 35569 8019
rect 35485 7966 35569 7991
rect 37625 7980 37713 7984
rect 35299 7940 35373 7949
rect 30619 7873 30691 7895
rect 30752 7888 31955 7923
rect 30752 7874 30780 7888
rect 30620 7673 30690 7873
rect 30754 7743 30780 7874
rect 31159 7885 31955 7888
rect 30612 7622 30692 7673
rect 30612 7596 30628 7622
rect 30668 7596 30692 7622
rect 30612 7577 30692 7596
rect 30612 7551 30631 7577
rect 30671 7551 30692 7577
rect 30612 7524 30692 7551
rect 30612 7498 30635 7524
rect 30675 7498 30692 7524
rect 30612 7487 30692 7498
rect 30754 7488 30781 7743
rect 31159 7735 31200 7885
rect 31431 7883 31535 7885
rect 31890 7851 31955 7885
rect 32932 7890 32998 7938
rect 35309 7936 35373 7940
rect 37625 7963 37889 7980
rect 37625 7909 37805 7963
rect 37868 7909 37889 7963
rect 35522 7899 36233 7901
rect 34895 7898 36233 7899
rect 33845 7897 33917 7898
rect 31626 7823 31747 7841
rect 31626 7821 31697 7823
rect 31626 7780 31641 7821
rect 31678 7782 31697 7821
rect 31734 7782 31747 7823
rect 31678 7780 31747 7782
rect 31626 7770 31747 7780
rect 31431 7740 31535 7743
rect 30821 7628 30885 7640
rect 31161 7636 31198 7735
rect 31426 7725 31537 7740
rect 31426 7723 31468 7725
rect 31426 7703 31433 7723
rect 31452 7703 31468 7723
rect 31426 7695 31468 7703
rect 31496 7723 31537 7725
rect 31496 7703 31510 7723
rect 31529 7703 31537 7723
rect 31496 7695 31537 7703
rect 31426 7689 31537 7695
rect 31369 7667 31618 7689
rect 31369 7636 31406 7667
rect 31582 7665 31618 7667
rect 31582 7636 31619 7665
rect 30821 7627 30856 7628
rect 30798 7622 30856 7627
rect 30798 7602 30801 7622
rect 30821 7608 30856 7622
rect 30876 7608 30885 7628
rect 30821 7600 30885 7608
rect 30847 7599 30885 7600
rect 30848 7598 30885 7599
rect 30951 7632 30987 7633
rect 31059 7632 31095 7633
rect 30951 7624 31095 7632
rect 30951 7604 30959 7624
rect 30979 7604 31067 7624
rect 31087 7604 31095 7624
rect 30951 7598 31095 7604
rect 31161 7628 31199 7636
rect 31267 7632 31303 7633
rect 31161 7608 31170 7628
rect 31190 7608 31199 7628
rect 31161 7599 31199 7608
rect 31218 7625 31303 7632
rect 31218 7605 31225 7625
rect 31246 7624 31303 7625
rect 31246 7605 31275 7624
rect 31218 7604 31275 7605
rect 31295 7604 31303 7624
rect 31161 7598 31198 7599
rect 31218 7598 31303 7604
rect 31369 7628 31407 7636
rect 31480 7632 31516 7633
rect 31369 7608 31378 7628
rect 31398 7608 31407 7628
rect 31369 7599 31407 7608
rect 31431 7624 31516 7632
rect 31431 7604 31488 7624
rect 31508 7604 31516 7624
rect 31369 7598 31406 7599
rect 31431 7598 31516 7604
rect 31582 7628 31620 7636
rect 31582 7608 31591 7628
rect 31611 7608 31620 7628
rect 31675 7618 31740 7770
rect 31893 7744 31948 7851
rect 32932 7816 32991 7890
rect 33844 7889 33943 7897
rect 33844 7886 33896 7889
rect 33844 7851 33852 7886
rect 33877 7851 33896 7886
rect 33921 7878 33943 7889
rect 34894 7890 36233 7898
rect 34894 7887 34946 7890
rect 33921 7877 34788 7878
rect 33921 7851 34789 7877
rect 33844 7841 34789 7851
rect 33844 7839 33943 7841
rect 32932 7798 32954 7816
rect 32972 7798 32991 7816
rect 32932 7776 32991 7798
rect 33199 7812 33731 7817
rect 33199 7792 34085 7812
rect 34105 7792 34108 7812
rect 34744 7808 34789 7841
rect 34894 7852 34902 7887
rect 34927 7852 34946 7887
rect 34971 7852 36233 7890
rect 34894 7843 36233 7852
rect 34894 7840 34983 7843
rect 35522 7841 36233 7843
rect 37625 7892 37889 7909
rect 33199 7788 34108 7792
rect 31582 7599 31620 7608
rect 31673 7611 31740 7618
rect 31582 7598 31619 7599
rect 31005 7577 31041 7598
rect 31431 7577 31462 7598
rect 31673 7590 31690 7611
rect 31726 7590 31740 7611
rect 31892 7631 31948 7744
rect 33199 7741 33242 7788
rect 33692 7787 34108 7788
rect 34740 7788 35133 7808
rect 35153 7788 35156 7808
rect 33692 7786 34033 7787
rect 33349 7755 33459 7769
rect 33349 7752 33392 7755
rect 33349 7747 33353 7752
rect 33187 7740 33242 7741
rect 31892 7613 31911 7631
rect 31929 7613 31948 7631
rect 31892 7593 31948 7613
rect 32931 7717 33242 7740
rect 32931 7699 32956 7717
rect 32974 7705 33242 7717
rect 33271 7725 33353 7747
rect 33382 7725 33392 7752
rect 33420 7728 33427 7755
rect 33456 7747 33459 7755
rect 33456 7728 33521 7747
rect 33420 7725 33521 7728
rect 33271 7723 33521 7725
rect 32974 7699 32996 7705
rect 31673 7577 31740 7590
rect 30838 7573 30938 7577
rect 30838 7569 30900 7573
rect 30838 7543 30845 7569
rect 30871 7547 30900 7569
rect 30926 7547 30938 7573
rect 30871 7543 30938 7547
rect 30838 7540 30938 7543
rect 31006 7540 31041 7577
rect 31103 7574 31462 7577
rect 31103 7569 31325 7574
rect 31103 7545 31116 7569
rect 31140 7550 31325 7569
rect 31349 7550 31462 7574
rect 31140 7545 31462 7550
rect 31103 7541 31462 7545
rect 31529 7571 31740 7577
rect 31529 7569 31690 7571
rect 31529 7549 31540 7569
rect 31560 7549 31690 7569
rect 31529 7542 31690 7549
rect 31529 7541 31570 7542
rect 31005 7515 31041 7540
rect 30853 7488 30890 7489
rect 30949 7488 30986 7489
rect 31005 7488 31012 7515
rect 30753 7479 30891 7488
rect 30753 7459 30862 7479
rect 30882 7459 30891 7479
rect 30753 7452 30891 7459
rect 30949 7485 31012 7488
rect 31033 7488 31041 7515
rect 31060 7488 31097 7489
rect 31033 7485 31097 7488
rect 30949 7479 31097 7485
rect 30949 7459 30958 7479
rect 30978 7459 31068 7479
rect 31088 7459 31097 7479
rect 30753 7450 30849 7452
rect 30949 7449 31097 7459
rect 31156 7479 31193 7489
rect 31268 7488 31305 7489
rect 31249 7486 31305 7488
rect 31156 7459 31164 7479
rect 31184 7459 31193 7479
rect 31005 7448 31041 7449
rect 30853 7317 30890 7318
rect 31156 7317 31193 7459
rect 31218 7479 31305 7486
rect 31218 7476 31276 7479
rect 31218 7456 31223 7476
rect 31244 7459 31276 7476
rect 31296 7459 31305 7479
rect 31244 7456 31305 7459
rect 31218 7449 31305 7456
rect 31364 7479 31401 7489
rect 31364 7459 31372 7479
rect 31392 7459 31401 7479
rect 31218 7448 31249 7449
rect 31364 7380 31401 7459
rect 31431 7488 31462 7541
rect 31675 7534 31690 7542
rect 31730 7534 31740 7571
rect 32931 7560 32996 7699
rect 33271 7644 33308 7723
rect 33349 7710 33459 7723
rect 33423 7654 33454 7655
rect 33271 7624 33280 7644
rect 33300 7624 33308 7644
rect 31675 7525 31740 7534
rect 31888 7532 31953 7553
rect 31888 7514 31913 7532
rect 31931 7514 31953 7532
rect 32931 7542 32954 7560
rect 32972 7542 32996 7560
rect 32931 7525 32996 7542
rect 33151 7606 33219 7619
rect 33271 7614 33308 7624
rect 33367 7644 33454 7654
rect 33367 7624 33376 7644
rect 33396 7624 33454 7644
rect 33367 7615 33454 7624
rect 33367 7614 33404 7615
rect 33151 7564 33158 7606
rect 33207 7564 33219 7606
rect 33151 7561 33219 7564
rect 33423 7562 33454 7615
rect 33484 7644 33521 7723
rect 33636 7654 33667 7655
rect 33484 7624 33493 7644
rect 33513 7624 33521 7644
rect 33484 7614 33521 7624
rect 33580 7647 33667 7654
rect 33580 7644 33641 7647
rect 33580 7624 33589 7644
rect 33609 7627 33641 7644
rect 33662 7627 33667 7647
rect 33609 7624 33667 7627
rect 33580 7617 33667 7624
rect 33692 7644 33729 7786
rect 33995 7785 34032 7786
rect 34740 7783 35156 7788
rect 34740 7782 35081 7783
rect 34397 7751 34507 7765
rect 34397 7748 34440 7751
rect 34397 7743 34401 7748
rect 34319 7721 34401 7743
rect 34430 7721 34440 7748
rect 34468 7724 34475 7751
rect 34504 7743 34507 7751
rect 34504 7724 34569 7743
rect 34468 7721 34569 7724
rect 34319 7719 34569 7721
rect 33844 7654 33880 7655
rect 33692 7624 33701 7644
rect 33721 7624 33729 7644
rect 33580 7615 33636 7617
rect 33580 7614 33617 7615
rect 33692 7614 33729 7624
rect 33788 7644 33936 7654
rect 34036 7651 34132 7653
rect 33788 7624 33797 7644
rect 33817 7624 33907 7644
rect 33927 7624 33936 7644
rect 33788 7618 33936 7624
rect 33788 7615 33852 7618
rect 33788 7614 33825 7615
rect 33844 7588 33852 7615
rect 33873 7615 33936 7618
rect 33994 7644 34132 7651
rect 33994 7624 34003 7644
rect 34023 7624 34132 7644
rect 33994 7615 34132 7624
rect 34319 7640 34356 7719
rect 34397 7706 34507 7719
rect 34471 7650 34502 7651
rect 34319 7620 34328 7640
rect 34348 7620 34356 7640
rect 33873 7588 33880 7615
rect 33899 7614 33936 7615
rect 33995 7614 34032 7615
rect 33844 7563 33880 7588
rect 33315 7561 33356 7562
rect 33151 7554 33356 7561
rect 33151 7543 33325 7554
rect 31481 7488 31518 7489
rect 31431 7479 31518 7488
rect 31431 7459 31489 7479
rect 31509 7459 31518 7479
rect 31431 7449 31518 7459
rect 31577 7479 31614 7489
rect 31577 7459 31585 7479
rect 31605 7459 31614 7479
rect 31431 7448 31462 7449
rect 31426 7380 31536 7393
rect 31577 7380 31614 7459
rect 31888 7438 31953 7514
rect 33151 7510 33159 7543
rect 33152 7501 33159 7510
rect 33208 7534 33325 7543
rect 33345 7534 33356 7554
rect 33208 7526 33356 7534
rect 33423 7558 33782 7562
rect 33423 7553 33745 7558
rect 33423 7529 33536 7553
rect 33560 7534 33745 7553
rect 33769 7534 33782 7558
rect 33560 7529 33782 7534
rect 33423 7526 33782 7529
rect 33844 7526 33879 7563
rect 33947 7560 34047 7563
rect 33947 7556 34014 7560
rect 33947 7530 33959 7556
rect 33985 7534 34014 7556
rect 34040 7534 34047 7560
rect 33985 7530 34047 7534
rect 33947 7526 34047 7530
rect 33208 7510 33219 7526
rect 33208 7501 33216 7510
rect 33423 7505 33454 7526
rect 33844 7505 33880 7526
rect 33266 7504 33303 7505
rect 32931 7461 32996 7480
rect 32931 7443 32956 7461
rect 32974 7443 32996 7461
rect 31364 7378 31614 7380
rect 31364 7375 31465 7378
rect 31364 7356 31429 7375
rect 31426 7348 31429 7356
rect 31458 7348 31465 7375
rect 31493 7351 31503 7378
rect 31532 7356 31614 7378
rect 31637 7403 31954 7438
rect 31532 7351 31536 7356
rect 31493 7348 31536 7351
rect 31426 7334 31536 7348
rect 30852 7316 31193 7317
rect 30777 7314 31193 7316
rect 31637 7314 31677 7403
rect 31888 7376 31953 7403
rect 31888 7358 31911 7376
rect 31929 7358 31953 7376
rect 31888 7338 31953 7358
rect 30774 7311 31677 7314
rect 30774 7291 30780 7311
rect 30800 7291 31677 7311
rect 30774 7287 31677 7291
rect 31637 7284 31677 7287
rect 31889 7277 31954 7298
rect 30107 7269 30768 7270
rect 30107 7262 31041 7269
rect 30107 7261 31013 7262
rect 30107 7241 30958 7261
rect 30990 7242 31013 7261
rect 31038 7242 31041 7262
rect 30990 7241 31041 7242
rect 30107 7234 31041 7241
rect 29706 7192 29874 7193
rect 30109 7192 30148 7234
rect 30937 7232 31041 7234
rect 31006 7230 31041 7232
rect 31889 7259 31913 7277
rect 31931 7259 31954 7277
rect 31889 7212 31954 7259
rect 29706 7166 30150 7192
rect 29706 7164 29874 7166
rect 29706 6813 29733 7164
rect 30109 7160 30150 7166
rect 29773 6953 29837 6965
rect 30113 6961 30150 7160
rect 30612 7187 30684 7204
rect 30612 7148 30620 7187
rect 30665 7148 30684 7187
rect 30378 7050 30489 7065
rect 30378 7048 30420 7050
rect 30378 7028 30385 7048
rect 30404 7028 30420 7048
rect 30378 7020 30420 7028
rect 30448 7048 30489 7050
rect 30448 7028 30462 7048
rect 30481 7028 30489 7048
rect 30448 7020 30489 7028
rect 30378 7014 30489 7020
rect 30321 6992 30570 7014
rect 30321 6961 30358 6992
rect 30534 6990 30570 6992
rect 30534 6961 30571 6990
rect 29773 6952 29808 6953
rect 29750 6947 29808 6952
rect 29750 6927 29753 6947
rect 29773 6933 29808 6947
rect 29828 6933 29837 6953
rect 29773 6925 29837 6933
rect 29799 6924 29837 6925
rect 29800 6923 29837 6924
rect 29903 6957 29939 6958
rect 30011 6957 30047 6958
rect 29903 6949 30047 6957
rect 29903 6929 29911 6949
rect 29931 6929 30019 6949
rect 30039 6929 30047 6949
rect 29903 6923 30047 6929
rect 30113 6953 30151 6961
rect 30219 6957 30255 6958
rect 30113 6933 30122 6953
rect 30142 6933 30151 6953
rect 30113 6924 30151 6933
rect 30170 6950 30255 6957
rect 30170 6930 30177 6950
rect 30198 6949 30255 6950
rect 30198 6930 30227 6949
rect 30170 6929 30227 6930
rect 30247 6929 30255 6949
rect 30113 6923 30150 6924
rect 30170 6923 30255 6929
rect 30321 6953 30359 6961
rect 30432 6957 30468 6958
rect 30321 6933 30330 6953
rect 30350 6933 30359 6953
rect 30321 6924 30359 6933
rect 30383 6949 30468 6957
rect 30383 6929 30440 6949
rect 30460 6929 30468 6949
rect 30321 6923 30358 6924
rect 30383 6923 30468 6929
rect 30534 6953 30572 6961
rect 30534 6933 30543 6953
rect 30563 6933 30572 6953
rect 30534 6924 30572 6933
rect 30612 6938 30684 7148
rect 30754 7182 31954 7212
rect 30754 7181 31198 7182
rect 30754 7179 30922 7181
rect 30612 6924 30695 6938
rect 30534 6923 30571 6924
rect 29957 6902 29993 6923
rect 30383 6902 30414 6923
rect 30612 6902 30629 6924
rect 29790 6898 29890 6902
rect 29790 6894 29852 6898
rect 29790 6868 29797 6894
rect 29823 6872 29852 6894
rect 29878 6872 29890 6898
rect 29823 6868 29890 6872
rect 29790 6865 29890 6868
rect 29958 6865 29993 6902
rect 30055 6899 30414 6902
rect 30055 6894 30277 6899
rect 30055 6870 30068 6894
rect 30092 6875 30277 6894
rect 30301 6875 30414 6899
rect 30092 6870 30414 6875
rect 30055 6866 30414 6870
rect 30481 6894 30629 6902
rect 30481 6874 30492 6894
rect 30512 6891 30629 6894
rect 30682 6891 30695 6924
rect 30512 6874 30695 6891
rect 30481 6867 30695 6874
rect 30481 6866 30522 6867
rect 30612 6866 30695 6867
rect 29957 6840 29993 6865
rect 29805 6813 29842 6814
rect 29901 6813 29938 6814
rect 29957 6813 29964 6840
rect 29705 6804 29843 6813
rect 29705 6784 29814 6804
rect 29834 6784 29843 6804
rect 29705 6777 29843 6784
rect 29901 6810 29964 6813
rect 29985 6813 29993 6840
rect 30012 6813 30049 6814
rect 29985 6810 30049 6813
rect 29901 6804 30049 6810
rect 29901 6784 29910 6804
rect 29930 6784 30020 6804
rect 30040 6784 30049 6804
rect 29705 6775 29801 6777
rect 29901 6774 30049 6784
rect 30108 6804 30145 6814
rect 30220 6813 30257 6814
rect 30201 6811 30257 6813
rect 30108 6784 30116 6804
rect 30136 6784 30145 6804
rect 29957 6773 29993 6774
rect 29805 6642 29842 6643
rect 30108 6642 30145 6784
rect 30170 6804 30257 6811
rect 30170 6801 30228 6804
rect 30170 6781 30175 6801
rect 30196 6784 30228 6801
rect 30248 6784 30257 6804
rect 30196 6781 30257 6784
rect 30170 6774 30257 6781
rect 30316 6804 30353 6814
rect 30316 6784 30324 6804
rect 30344 6784 30353 6804
rect 30170 6773 30201 6774
rect 30316 6705 30353 6784
rect 30383 6813 30414 6866
rect 30620 6833 30634 6866
rect 30687 6833 30695 6866
rect 30620 6827 30695 6833
rect 30620 6822 30690 6827
rect 30433 6813 30470 6814
rect 30383 6804 30470 6813
rect 30383 6784 30441 6804
rect 30461 6784 30470 6804
rect 30383 6774 30470 6784
rect 30529 6804 30566 6814
rect 30754 6809 30781 7179
rect 30821 6949 30885 6961
rect 31161 6957 31198 7181
rect 31669 7162 31733 7164
rect 31665 7150 31733 7162
rect 31665 7117 31676 7150
rect 31716 7117 31733 7150
rect 31665 7107 31733 7117
rect 31426 7046 31537 7061
rect 31426 7044 31468 7046
rect 31426 7024 31433 7044
rect 31452 7024 31468 7044
rect 31426 7016 31468 7024
rect 31496 7044 31537 7046
rect 31496 7024 31510 7044
rect 31529 7024 31537 7044
rect 31496 7016 31537 7024
rect 31426 7010 31537 7016
rect 31369 6988 31618 7010
rect 31369 6957 31406 6988
rect 31582 6986 31618 6988
rect 31582 6957 31619 6986
rect 30821 6948 30856 6949
rect 30798 6943 30856 6948
rect 30798 6923 30801 6943
rect 30821 6929 30856 6943
rect 30876 6929 30885 6949
rect 30821 6921 30885 6929
rect 30847 6920 30885 6921
rect 30848 6919 30885 6920
rect 30951 6953 30987 6954
rect 31059 6953 31095 6954
rect 30951 6945 31095 6953
rect 30951 6925 30959 6945
rect 30979 6925 31067 6945
rect 31087 6925 31095 6945
rect 30951 6919 31095 6925
rect 31161 6949 31199 6957
rect 31267 6953 31303 6954
rect 31161 6929 31170 6949
rect 31190 6929 31199 6949
rect 31161 6920 31199 6929
rect 31218 6946 31303 6953
rect 31218 6926 31225 6946
rect 31246 6945 31303 6946
rect 31246 6926 31275 6945
rect 31218 6925 31275 6926
rect 31295 6925 31303 6945
rect 31161 6919 31198 6920
rect 31218 6919 31303 6925
rect 31369 6949 31407 6957
rect 31480 6953 31516 6954
rect 31369 6929 31378 6949
rect 31398 6929 31407 6949
rect 31369 6920 31407 6929
rect 31431 6945 31516 6953
rect 31431 6925 31488 6945
rect 31508 6925 31516 6945
rect 31369 6919 31406 6920
rect 31431 6919 31516 6925
rect 31582 6949 31620 6957
rect 31582 6929 31591 6949
rect 31611 6929 31620 6949
rect 31582 6920 31620 6929
rect 31669 6923 31733 7107
rect 31889 6981 31954 7182
rect 32931 7242 32996 7443
rect 33152 7317 33216 7501
rect 33265 7495 33303 7504
rect 33265 7475 33274 7495
rect 33294 7475 33303 7495
rect 33265 7467 33303 7475
rect 33369 7499 33454 7505
rect 33479 7504 33516 7505
rect 33369 7479 33377 7499
rect 33397 7479 33454 7499
rect 33369 7471 33454 7479
rect 33478 7495 33516 7504
rect 33478 7475 33487 7495
rect 33507 7475 33516 7495
rect 33369 7470 33405 7471
rect 33478 7467 33516 7475
rect 33582 7499 33667 7505
rect 33687 7504 33724 7505
rect 33582 7479 33590 7499
rect 33610 7498 33667 7499
rect 33610 7479 33639 7498
rect 33582 7478 33639 7479
rect 33660 7478 33667 7498
rect 33582 7471 33667 7478
rect 33686 7495 33724 7504
rect 33686 7475 33695 7495
rect 33715 7475 33724 7495
rect 33582 7470 33618 7471
rect 33686 7467 33724 7475
rect 33790 7499 33934 7505
rect 33790 7479 33798 7499
rect 33818 7479 33906 7499
rect 33926 7479 33934 7499
rect 33790 7471 33934 7479
rect 33790 7470 33826 7471
rect 33898 7470 33934 7471
rect 34000 7504 34037 7505
rect 34000 7503 34038 7504
rect 34000 7495 34064 7503
rect 34000 7475 34009 7495
rect 34029 7481 34064 7495
rect 34084 7481 34087 7501
rect 34029 7476 34087 7481
rect 34029 7475 34064 7476
rect 33266 7438 33303 7467
rect 33267 7436 33303 7438
rect 33479 7436 33516 7467
rect 33267 7414 33516 7436
rect 33348 7408 33459 7414
rect 33348 7400 33389 7408
rect 33348 7380 33356 7400
rect 33375 7380 33389 7400
rect 33348 7378 33389 7380
rect 33417 7400 33459 7408
rect 33417 7380 33433 7400
rect 33452 7380 33459 7400
rect 33417 7378 33459 7380
rect 33348 7363 33459 7378
rect 33152 7307 33220 7317
rect 33152 7274 33169 7307
rect 33209 7274 33220 7307
rect 33152 7262 33220 7274
rect 33152 7260 33216 7262
rect 33687 7243 33724 7467
rect 34000 7463 34064 7475
rect 34104 7245 34131 7615
rect 34319 7610 34356 7620
rect 34415 7640 34502 7650
rect 34415 7620 34424 7640
rect 34444 7620 34502 7640
rect 34415 7611 34502 7620
rect 34415 7610 34452 7611
rect 34195 7597 34265 7602
rect 34190 7591 34265 7597
rect 34190 7558 34198 7591
rect 34251 7558 34265 7591
rect 34471 7558 34502 7611
rect 34532 7640 34569 7719
rect 34684 7650 34715 7651
rect 34532 7620 34541 7640
rect 34561 7620 34569 7640
rect 34532 7610 34569 7620
rect 34628 7643 34715 7650
rect 34628 7640 34689 7643
rect 34628 7620 34637 7640
rect 34657 7623 34689 7640
rect 34710 7623 34715 7643
rect 34657 7620 34715 7623
rect 34628 7613 34715 7620
rect 34740 7640 34777 7782
rect 35043 7781 35080 7782
rect 34892 7650 34928 7651
rect 34740 7620 34749 7640
rect 34769 7620 34777 7640
rect 34628 7611 34684 7613
rect 34628 7610 34665 7611
rect 34740 7610 34777 7620
rect 34836 7640 34984 7650
rect 35084 7647 35180 7649
rect 34836 7620 34845 7640
rect 34865 7620 34955 7640
rect 34975 7620 34984 7640
rect 34836 7614 34984 7620
rect 34836 7611 34900 7614
rect 34836 7610 34873 7611
rect 34892 7584 34900 7611
rect 34921 7611 34984 7614
rect 35042 7640 35180 7647
rect 35042 7620 35051 7640
rect 35071 7620 35180 7640
rect 35042 7611 35180 7620
rect 34921 7584 34928 7611
rect 34947 7610 34984 7611
rect 35043 7610 35080 7611
rect 34892 7559 34928 7584
rect 34190 7557 34273 7558
rect 34363 7557 34404 7558
rect 34190 7550 34404 7557
rect 34190 7533 34373 7550
rect 34190 7500 34203 7533
rect 34256 7530 34373 7533
rect 34393 7530 34404 7550
rect 34256 7522 34404 7530
rect 34471 7554 34830 7558
rect 34471 7549 34793 7554
rect 34471 7525 34584 7549
rect 34608 7530 34793 7549
rect 34817 7530 34830 7554
rect 34608 7525 34830 7530
rect 34471 7522 34830 7525
rect 34892 7522 34927 7559
rect 34995 7556 35095 7559
rect 34995 7552 35062 7556
rect 34995 7526 35007 7552
rect 35033 7530 35062 7552
rect 35088 7530 35095 7556
rect 35033 7526 35095 7530
rect 34995 7522 35095 7526
rect 34256 7500 34273 7522
rect 34471 7501 34502 7522
rect 34892 7501 34928 7522
rect 34314 7500 34351 7501
rect 34190 7486 34273 7500
rect 33963 7243 34131 7245
rect 33687 7242 34131 7243
rect 32931 7212 34131 7242
rect 34201 7276 34273 7486
rect 34313 7491 34351 7500
rect 34313 7471 34322 7491
rect 34342 7471 34351 7491
rect 34313 7463 34351 7471
rect 34417 7495 34502 7501
rect 34527 7500 34564 7501
rect 34417 7475 34425 7495
rect 34445 7475 34502 7495
rect 34417 7467 34502 7475
rect 34526 7491 34564 7500
rect 34526 7471 34535 7491
rect 34555 7471 34564 7491
rect 34417 7466 34453 7467
rect 34526 7463 34564 7471
rect 34630 7495 34715 7501
rect 34735 7500 34772 7501
rect 34630 7475 34638 7495
rect 34658 7494 34715 7495
rect 34658 7475 34687 7494
rect 34630 7474 34687 7475
rect 34708 7474 34715 7494
rect 34630 7467 34715 7474
rect 34734 7491 34772 7500
rect 34734 7471 34743 7491
rect 34763 7471 34772 7491
rect 34630 7466 34666 7467
rect 34734 7463 34772 7471
rect 34838 7495 34982 7501
rect 34838 7475 34846 7495
rect 34866 7475 34954 7495
rect 34974 7475 34982 7495
rect 34838 7467 34982 7475
rect 34838 7466 34874 7467
rect 34946 7466 34982 7467
rect 35048 7500 35085 7501
rect 35048 7499 35086 7500
rect 35048 7491 35112 7499
rect 35048 7471 35057 7491
rect 35077 7477 35112 7491
rect 35132 7477 35135 7497
rect 35077 7472 35135 7477
rect 35077 7471 35112 7472
rect 34314 7434 34351 7463
rect 34315 7432 34351 7434
rect 34527 7432 34564 7463
rect 34315 7410 34564 7432
rect 34396 7404 34507 7410
rect 34396 7396 34437 7404
rect 34396 7376 34404 7396
rect 34423 7376 34437 7396
rect 34396 7374 34437 7376
rect 34465 7396 34507 7404
rect 34465 7376 34481 7396
rect 34500 7376 34507 7396
rect 34465 7374 34507 7376
rect 34396 7359 34507 7374
rect 34201 7237 34220 7276
rect 34265 7237 34273 7276
rect 34201 7220 34273 7237
rect 34735 7264 34772 7463
rect 35048 7459 35112 7471
rect 34735 7258 34776 7264
rect 35152 7260 35179 7611
rect 35474 7598 35569 7624
rect 35310 7576 35374 7595
rect 35310 7537 35323 7576
rect 35357 7537 35374 7576
rect 35310 7518 35374 7537
rect 35011 7258 35179 7260
rect 34735 7232 35179 7258
rect 32931 7165 32996 7212
rect 32931 7147 32954 7165
rect 32972 7147 32996 7165
rect 33844 7192 33879 7194
rect 33844 7190 33948 7192
rect 34737 7190 34776 7232
rect 35011 7231 35179 7232
rect 33844 7183 34778 7190
rect 33844 7182 33895 7183
rect 33844 7162 33847 7182
rect 33872 7163 33895 7182
rect 33927 7163 34778 7183
rect 33872 7162 34778 7163
rect 33844 7155 34778 7162
rect 34117 7154 34778 7155
rect 32931 7126 32996 7147
rect 33208 7137 33248 7140
rect 33208 7133 34111 7137
rect 33208 7113 34085 7133
rect 34105 7113 34111 7133
rect 33208 7110 34111 7113
rect 32932 7066 32997 7086
rect 32932 7048 32956 7066
rect 32974 7048 32997 7066
rect 32932 7021 32997 7048
rect 33208 7021 33248 7110
rect 33692 7108 34108 7110
rect 33692 7107 34033 7108
rect 33349 7076 33459 7090
rect 33349 7073 33392 7076
rect 33349 7068 33353 7073
rect 32931 6986 33248 7021
rect 33271 7046 33353 7068
rect 33382 7046 33392 7073
rect 33420 7049 33427 7076
rect 33456 7068 33459 7076
rect 33456 7049 33521 7068
rect 33420 7046 33521 7049
rect 33271 7044 33521 7046
rect 31889 6963 31911 6981
rect 31929 6963 31954 6981
rect 31889 6944 31954 6963
rect 31582 6919 31619 6920
rect 31005 6898 31041 6919
rect 31431 6898 31462 6919
rect 31669 6914 31677 6923
rect 31666 6898 31677 6914
rect 30838 6894 30938 6898
rect 30838 6890 30900 6894
rect 30838 6864 30845 6890
rect 30871 6868 30900 6890
rect 30926 6868 30938 6894
rect 30871 6864 30938 6868
rect 30838 6861 30938 6864
rect 31006 6861 31041 6898
rect 31103 6895 31462 6898
rect 31103 6890 31325 6895
rect 31103 6866 31116 6890
rect 31140 6871 31325 6890
rect 31349 6871 31462 6895
rect 31140 6866 31462 6871
rect 31103 6862 31462 6866
rect 31529 6890 31677 6898
rect 31529 6870 31540 6890
rect 31560 6881 31677 6890
rect 31726 6914 31733 6923
rect 31726 6881 31734 6914
rect 32932 6910 32997 6986
rect 33271 6965 33308 7044
rect 33349 7031 33459 7044
rect 33423 6975 33454 6976
rect 33271 6945 33280 6965
rect 33300 6945 33308 6965
rect 33271 6935 33308 6945
rect 33367 6965 33454 6975
rect 33367 6945 33376 6965
rect 33396 6945 33454 6965
rect 33367 6936 33454 6945
rect 33367 6935 33404 6936
rect 31560 6870 31734 6881
rect 31529 6863 31734 6870
rect 31529 6862 31570 6863
rect 31005 6836 31041 6861
rect 30853 6809 30890 6810
rect 30949 6809 30986 6810
rect 31005 6809 31012 6836
rect 30529 6784 30537 6804
rect 30557 6784 30566 6804
rect 30383 6773 30414 6774
rect 30378 6705 30488 6718
rect 30529 6705 30566 6784
rect 30753 6800 30891 6809
rect 30753 6780 30862 6800
rect 30882 6780 30891 6800
rect 30753 6773 30891 6780
rect 30949 6806 31012 6809
rect 31033 6809 31041 6836
rect 31060 6809 31097 6810
rect 31033 6806 31097 6809
rect 30949 6800 31097 6806
rect 30949 6780 30958 6800
rect 30978 6780 31068 6800
rect 31088 6780 31097 6800
rect 30753 6771 30849 6773
rect 30949 6770 31097 6780
rect 31156 6800 31193 6810
rect 31268 6809 31305 6810
rect 31249 6807 31305 6809
rect 31156 6780 31164 6800
rect 31184 6780 31193 6800
rect 31005 6769 31041 6770
rect 30316 6703 30566 6705
rect 30316 6700 30417 6703
rect 30316 6681 30381 6700
rect 30378 6673 30381 6681
rect 30410 6673 30417 6700
rect 30445 6676 30455 6703
rect 30484 6681 30566 6703
rect 30484 6676 30488 6681
rect 30445 6673 30488 6676
rect 30378 6659 30488 6673
rect 29804 6641 30145 6642
rect 29729 6636 30145 6641
rect 30853 6638 30890 6639
rect 31156 6638 31193 6780
rect 31218 6800 31305 6807
rect 31218 6797 31276 6800
rect 31218 6777 31223 6797
rect 31244 6780 31276 6797
rect 31296 6780 31305 6800
rect 31244 6777 31305 6780
rect 31218 6770 31305 6777
rect 31364 6800 31401 6810
rect 31364 6780 31372 6800
rect 31392 6780 31401 6800
rect 31218 6769 31249 6770
rect 31364 6701 31401 6780
rect 31431 6809 31462 6862
rect 31666 6860 31734 6863
rect 31666 6818 31678 6860
rect 31727 6818 31734 6860
rect 31481 6809 31518 6810
rect 31431 6800 31518 6809
rect 31431 6780 31489 6800
rect 31509 6780 31518 6800
rect 31431 6770 31518 6780
rect 31577 6800 31614 6810
rect 31666 6805 31734 6818
rect 31889 6882 31954 6899
rect 31889 6864 31913 6882
rect 31931 6864 31954 6882
rect 32932 6892 32954 6910
rect 32972 6892 32997 6910
rect 32932 6871 32997 6892
rect 33145 6890 33210 6899
rect 31577 6780 31585 6800
rect 31605 6780 31614 6800
rect 31431 6769 31462 6770
rect 31426 6701 31536 6714
rect 31577 6701 31614 6780
rect 31889 6725 31954 6864
rect 33145 6853 33155 6890
rect 33195 6882 33210 6890
rect 33423 6883 33454 6936
rect 33484 6965 33521 7044
rect 33636 6975 33667 6976
rect 33484 6945 33493 6965
rect 33513 6945 33521 6965
rect 33484 6935 33521 6945
rect 33580 6968 33667 6975
rect 33580 6965 33641 6968
rect 33580 6945 33589 6965
rect 33609 6948 33641 6965
rect 33662 6948 33667 6968
rect 33609 6945 33667 6948
rect 33580 6938 33667 6945
rect 33692 6965 33729 7107
rect 33995 7106 34032 7107
rect 35312 7047 35374 7518
rect 35474 7557 35500 7598
rect 35536 7557 35569 7598
rect 35474 7261 35569 7557
rect 35474 7217 35489 7261
rect 35549 7217 35569 7261
rect 35474 7197 35569 7217
rect 36186 7128 36229 7841
rect 36186 7108 36580 7128
rect 36600 7108 36603 7128
rect 36187 7103 36603 7108
rect 36187 7102 36528 7103
rect 35844 7071 35954 7085
rect 35844 7068 35887 7071
rect 35844 7063 35848 7068
rect 35307 6995 35382 7047
rect 35766 7041 35848 7063
rect 35877 7041 35887 7068
rect 35915 7044 35922 7071
rect 35951 7063 35954 7071
rect 35951 7044 36016 7063
rect 35915 7041 36016 7044
rect 35766 7039 36016 7041
rect 35676 6995 35722 6996
rect 33844 6975 33880 6976
rect 33692 6945 33701 6965
rect 33721 6945 33729 6965
rect 33580 6936 33636 6938
rect 33580 6935 33617 6936
rect 33692 6935 33729 6945
rect 33788 6965 33936 6975
rect 34036 6972 34132 6974
rect 33788 6945 33797 6965
rect 33817 6945 33907 6965
rect 33927 6945 33936 6965
rect 33788 6939 33936 6945
rect 33788 6936 33852 6939
rect 33788 6935 33825 6936
rect 33844 6909 33852 6936
rect 33873 6936 33936 6939
rect 33994 6965 34132 6972
rect 33994 6945 34003 6965
rect 34023 6945 34132 6965
rect 33994 6936 34132 6945
rect 35307 6960 35722 6995
rect 33873 6909 33880 6936
rect 33899 6935 33936 6936
rect 33995 6935 34032 6936
rect 33844 6884 33880 6909
rect 33315 6882 33356 6883
rect 33195 6875 33356 6882
rect 33195 6855 33325 6875
rect 33345 6855 33356 6875
rect 33195 6853 33356 6855
rect 33145 6847 33356 6853
rect 33423 6879 33782 6883
rect 33423 6874 33745 6879
rect 33423 6850 33536 6874
rect 33560 6855 33745 6874
rect 33769 6855 33782 6879
rect 33560 6850 33782 6855
rect 33423 6847 33782 6850
rect 33844 6847 33879 6884
rect 33947 6881 34047 6884
rect 33947 6877 34014 6881
rect 33947 6851 33959 6877
rect 33985 6855 34014 6877
rect 34040 6855 34047 6881
rect 33985 6851 34047 6855
rect 33947 6847 34047 6851
rect 33145 6834 33212 6847
rect 31889 6719 31911 6725
rect 31364 6699 31614 6701
rect 31364 6696 31465 6699
rect 31364 6677 31429 6696
rect 31426 6669 31429 6677
rect 31458 6669 31465 6696
rect 31493 6672 31503 6699
rect 31532 6677 31614 6699
rect 31643 6707 31911 6719
rect 31929 6707 31954 6725
rect 31643 6684 31954 6707
rect 32937 6811 32993 6831
rect 32937 6793 32956 6811
rect 32974 6793 32993 6811
rect 31643 6683 31698 6684
rect 31532 6672 31536 6677
rect 31493 6669 31536 6672
rect 31426 6655 31536 6669
rect 30852 6637 31193 6638
rect 29729 6616 29732 6636
rect 29752 6616 30145 6636
rect 30777 6636 31193 6637
rect 31643 6636 31686 6683
rect 32937 6680 32993 6793
rect 33145 6813 33159 6834
rect 33195 6813 33212 6834
rect 33423 6826 33454 6847
rect 33844 6826 33880 6847
rect 33266 6825 33303 6826
rect 33145 6806 33212 6813
rect 33265 6816 33303 6825
rect 30777 6632 31686 6636
rect 30096 6583 30141 6616
rect 30777 6612 30780 6632
rect 30800 6612 31686 6632
rect 31154 6607 31686 6612
rect 31894 6626 31953 6648
rect 31894 6608 31913 6626
rect 31931 6608 31953 6626
rect 30942 6583 31041 6585
rect 30096 6573 31041 6583
rect 30096 6547 30964 6573
rect 30097 6546 30964 6547
rect 30942 6535 30964 6546
rect 30989 6538 31008 6573
rect 31033 6538 31041 6573
rect 30989 6535 31041 6538
rect 31894 6537 31953 6608
rect 32937 6542 32992 6680
rect 33145 6654 33210 6806
rect 33265 6796 33274 6816
rect 33294 6796 33303 6816
rect 33265 6788 33303 6796
rect 33369 6820 33454 6826
rect 33479 6825 33516 6826
rect 33369 6800 33377 6820
rect 33397 6800 33454 6820
rect 33369 6792 33454 6800
rect 33478 6816 33516 6825
rect 33478 6796 33487 6816
rect 33507 6796 33516 6816
rect 33369 6791 33405 6792
rect 33478 6788 33516 6796
rect 33582 6820 33667 6826
rect 33687 6825 33724 6826
rect 33582 6800 33590 6820
rect 33610 6819 33667 6820
rect 33610 6800 33639 6819
rect 33582 6799 33639 6800
rect 33660 6799 33667 6819
rect 33582 6792 33667 6799
rect 33686 6816 33724 6825
rect 33686 6796 33695 6816
rect 33715 6796 33724 6816
rect 33582 6791 33618 6792
rect 33686 6788 33724 6796
rect 33790 6820 33934 6826
rect 33790 6800 33798 6820
rect 33818 6800 33906 6820
rect 33926 6800 33934 6820
rect 33790 6792 33934 6800
rect 33790 6791 33826 6792
rect 33898 6791 33934 6792
rect 34000 6825 34037 6826
rect 34000 6824 34038 6825
rect 34000 6816 34064 6824
rect 34000 6796 34009 6816
rect 34029 6802 34064 6816
rect 34084 6802 34087 6822
rect 34029 6797 34087 6802
rect 34029 6796 34064 6797
rect 33266 6759 33303 6788
rect 33267 6757 33303 6759
rect 33479 6757 33516 6788
rect 33267 6735 33516 6757
rect 33348 6729 33459 6735
rect 33348 6721 33389 6729
rect 33348 6701 33356 6721
rect 33375 6701 33389 6721
rect 33348 6699 33389 6701
rect 33417 6721 33459 6729
rect 33417 6701 33433 6721
rect 33452 6701 33459 6721
rect 33417 6699 33459 6701
rect 33348 6686 33459 6699
rect 33687 6689 33724 6788
rect 34000 6784 34064 6796
rect 33138 6644 33259 6654
rect 33138 6642 33207 6644
rect 33138 6601 33151 6642
rect 33188 6603 33207 6642
rect 33244 6603 33259 6644
rect 33188 6601 33259 6603
rect 33138 6583 33259 6601
rect 32930 6539 32994 6542
rect 33350 6539 33454 6545
rect 33685 6539 33726 6689
rect 34104 6681 34131 6936
rect 34193 6926 34273 6937
rect 34193 6900 34210 6926
rect 34250 6900 34273 6926
rect 34193 6873 34273 6900
rect 34193 6847 34214 6873
rect 34254 6847 34273 6873
rect 34193 6828 34273 6847
rect 34193 6802 34217 6828
rect 34257 6802 34273 6828
rect 34193 6751 34273 6802
rect 30942 6527 31041 6535
rect 30968 6526 31040 6527
rect 30622 6500 30689 6519
rect 30622 6479 30639 6500
rect 30620 6434 30639 6479
rect 30669 6479 30689 6500
rect 30669 6434 30690 6479
rect 31159 6476 31200 6478
rect 31431 6476 31535 6478
rect 31891 6476 31955 6537
rect 30620 6226 30690 6434
rect 30752 6441 31955 6476
rect 30752 6427 30780 6441
rect 30754 6296 30780 6427
rect 31159 6438 31955 6441
rect 32930 6536 33726 6539
rect 34105 6550 34131 6681
rect 34105 6536 34133 6550
rect 32930 6501 34133 6536
rect 34195 6543 34265 6751
rect 35307 6676 35382 6960
rect 35676 6877 35722 6960
rect 35766 6960 35803 7039
rect 35844 7026 35954 7039
rect 35918 6970 35949 6971
rect 35766 6940 35775 6960
rect 35795 6940 35803 6960
rect 35766 6930 35803 6940
rect 35862 6960 35949 6970
rect 35862 6940 35871 6960
rect 35891 6940 35949 6960
rect 35862 6931 35949 6940
rect 35862 6930 35899 6931
rect 35918 6878 35949 6931
rect 35979 6960 36016 7039
rect 36131 6970 36162 6971
rect 35979 6940 35988 6960
rect 36008 6940 36016 6960
rect 35979 6930 36016 6940
rect 36075 6963 36162 6970
rect 36075 6960 36136 6963
rect 36075 6940 36084 6960
rect 36104 6943 36136 6960
rect 36157 6943 36162 6963
rect 36104 6940 36162 6943
rect 36075 6933 36162 6940
rect 36187 6960 36224 7102
rect 36490 7101 36527 7102
rect 36339 6970 36375 6971
rect 36187 6940 36196 6960
rect 36216 6940 36224 6960
rect 36075 6931 36131 6933
rect 36075 6930 36112 6931
rect 36187 6930 36224 6940
rect 36283 6960 36431 6970
rect 36531 6967 36627 6969
rect 36283 6940 36292 6960
rect 36312 6940 36402 6960
rect 36422 6940 36431 6960
rect 36283 6934 36431 6940
rect 36283 6931 36347 6934
rect 36283 6930 36320 6931
rect 36339 6904 36347 6931
rect 36368 6931 36431 6934
rect 36489 6960 36627 6967
rect 36489 6940 36498 6960
rect 36518 6940 36627 6960
rect 36489 6931 36627 6940
rect 36368 6904 36375 6931
rect 36394 6930 36431 6931
rect 36490 6930 36527 6931
rect 36339 6879 36375 6904
rect 35810 6877 35851 6878
rect 35676 6870 35851 6877
rect 35474 6844 35560 6863
rect 35474 6803 35489 6844
rect 35543 6803 35560 6844
rect 35676 6850 35820 6870
rect 35840 6850 35851 6870
rect 35676 6842 35851 6850
rect 35918 6874 36277 6878
rect 35918 6869 36240 6874
rect 35918 6845 36031 6869
rect 36055 6850 36240 6869
rect 36264 6850 36277 6874
rect 36055 6845 36277 6850
rect 35918 6842 36277 6845
rect 36339 6842 36374 6879
rect 36442 6876 36542 6879
rect 36442 6872 36509 6876
rect 36442 6846 36454 6872
rect 36480 6850 36509 6872
rect 36535 6850 36542 6876
rect 36480 6846 36542 6850
rect 36442 6842 36542 6846
rect 35676 6838 35722 6842
rect 35918 6821 35949 6842
rect 36339 6821 36375 6842
rect 35761 6820 35798 6821
rect 35474 6767 35560 6803
rect 35760 6811 35798 6820
rect 35760 6791 35769 6811
rect 35789 6791 35798 6811
rect 35760 6783 35798 6791
rect 35864 6815 35949 6821
rect 35974 6820 36011 6821
rect 35864 6795 35872 6815
rect 35892 6795 35949 6815
rect 35864 6787 35949 6795
rect 35973 6811 36011 6820
rect 35973 6791 35982 6811
rect 36002 6791 36011 6811
rect 35864 6786 35900 6787
rect 35973 6783 36011 6791
rect 36077 6815 36162 6821
rect 36182 6820 36219 6821
rect 36077 6795 36085 6815
rect 36105 6814 36162 6815
rect 36105 6795 36134 6814
rect 36077 6794 36134 6795
rect 36155 6794 36162 6814
rect 36077 6787 36162 6794
rect 36181 6811 36219 6820
rect 36181 6791 36190 6811
rect 36210 6791 36219 6811
rect 36077 6786 36113 6787
rect 36181 6783 36219 6791
rect 36285 6815 36429 6821
rect 36285 6795 36293 6815
rect 36313 6795 36401 6815
rect 36421 6795 36429 6815
rect 36285 6787 36429 6795
rect 36285 6786 36321 6787
rect 32930 6440 32994 6501
rect 33350 6499 33454 6501
rect 33685 6499 33726 6501
rect 34195 6498 34216 6543
rect 34196 6477 34216 6498
rect 34246 6498 34265 6543
rect 35302 6634 35382 6676
rect 34246 6477 34263 6498
rect 34196 6458 34263 6477
rect 33845 6450 33917 6451
rect 33844 6442 33943 6450
rect 29507 6134 29589 6154
rect 29507 6111 29535 6134
rect 29561 6111 29589 6134
rect 29507 6049 29589 6111
rect 29511 6014 29589 6049
rect 30612 6175 30692 6226
rect 30612 6149 30628 6175
rect 30668 6149 30692 6175
rect 30612 6130 30692 6149
rect 30612 6104 30631 6130
rect 30671 6104 30692 6130
rect 30612 6077 30692 6104
rect 30612 6051 30635 6077
rect 30675 6051 30692 6077
rect 30612 6040 30692 6051
rect 30754 6041 30781 6296
rect 31159 6288 31200 6438
rect 31431 6432 31535 6438
rect 31891 6435 31955 6438
rect 31626 6376 31747 6394
rect 31626 6374 31697 6376
rect 31626 6333 31641 6374
rect 31678 6335 31697 6374
rect 31734 6335 31747 6376
rect 31678 6333 31747 6335
rect 31626 6323 31747 6333
rect 30821 6181 30885 6193
rect 31161 6189 31198 6288
rect 31426 6278 31537 6291
rect 31426 6276 31468 6278
rect 31426 6256 31433 6276
rect 31452 6256 31468 6276
rect 31426 6248 31468 6256
rect 31496 6276 31537 6278
rect 31496 6256 31510 6276
rect 31529 6256 31537 6276
rect 31496 6248 31537 6256
rect 31426 6242 31537 6248
rect 31369 6220 31618 6242
rect 31369 6189 31406 6220
rect 31582 6218 31618 6220
rect 31582 6189 31619 6218
rect 30821 6180 30856 6181
rect 30798 6175 30856 6180
rect 30798 6155 30801 6175
rect 30821 6161 30856 6175
rect 30876 6161 30885 6181
rect 30821 6153 30885 6161
rect 30847 6152 30885 6153
rect 30848 6151 30885 6152
rect 30951 6185 30987 6186
rect 31059 6185 31095 6186
rect 30951 6177 31095 6185
rect 30951 6157 30959 6177
rect 30979 6157 31067 6177
rect 31087 6157 31095 6177
rect 30951 6151 31095 6157
rect 31161 6181 31199 6189
rect 31267 6185 31303 6186
rect 31161 6161 31170 6181
rect 31190 6161 31199 6181
rect 31161 6152 31199 6161
rect 31218 6178 31303 6185
rect 31218 6158 31225 6178
rect 31246 6177 31303 6178
rect 31246 6158 31275 6177
rect 31218 6157 31275 6158
rect 31295 6157 31303 6177
rect 31161 6151 31198 6152
rect 31218 6151 31303 6157
rect 31369 6181 31407 6189
rect 31480 6185 31516 6186
rect 31369 6161 31378 6181
rect 31398 6161 31407 6181
rect 31369 6152 31407 6161
rect 31431 6177 31516 6185
rect 31431 6157 31488 6177
rect 31508 6157 31516 6177
rect 31369 6151 31406 6152
rect 31431 6151 31516 6157
rect 31582 6181 31620 6189
rect 31582 6161 31591 6181
rect 31611 6161 31620 6181
rect 31675 6171 31740 6323
rect 31893 6297 31948 6435
rect 32932 6369 32991 6440
rect 33844 6439 33896 6442
rect 33844 6404 33852 6439
rect 33877 6404 33896 6439
rect 33921 6431 33943 6442
rect 33921 6430 34788 6431
rect 33921 6404 34789 6430
rect 33844 6394 34789 6404
rect 33844 6392 33943 6394
rect 32932 6351 32954 6369
rect 32972 6351 32991 6369
rect 32932 6329 32991 6351
rect 33199 6365 33731 6370
rect 33199 6345 34085 6365
rect 34105 6345 34108 6365
rect 34744 6361 34789 6394
rect 33199 6341 34108 6345
rect 31582 6152 31620 6161
rect 31673 6164 31740 6171
rect 31582 6151 31619 6152
rect 31005 6130 31041 6151
rect 31431 6130 31462 6151
rect 31673 6143 31690 6164
rect 31726 6143 31740 6164
rect 31892 6184 31948 6297
rect 33199 6294 33242 6341
rect 33692 6340 34108 6341
rect 34740 6341 35133 6361
rect 35153 6341 35156 6361
rect 33692 6339 34033 6340
rect 33349 6308 33459 6322
rect 33349 6305 33392 6308
rect 33349 6300 33353 6305
rect 33187 6293 33242 6294
rect 31892 6166 31911 6184
rect 31929 6166 31948 6184
rect 31892 6146 31948 6166
rect 32931 6270 33242 6293
rect 32931 6252 32956 6270
rect 32974 6258 33242 6270
rect 33271 6278 33353 6300
rect 33382 6278 33392 6305
rect 33420 6281 33427 6308
rect 33456 6300 33459 6308
rect 33456 6281 33521 6300
rect 33420 6278 33521 6281
rect 33271 6276 33521 6278
rect 32974 6252 32996 6258
rect 31673 6130 31740 6143
rect 30838 6126 30938 6130
rect 30838 6122 30900 6126
rect 30838 6096 30845 6122
rect 30871 6100 30900 6122
rect 30926 6100 30938 6126
rect 30871 6096 30938 6100
rect 30838 6093 30938 6096
rect 31006 6093 31041 6130
rect 31103 6127 31462 6130
rect 31103 6122 31325 6127
rect 31103 6098 31116 6122
rect 31140 6103 31325 6122
rect 31349 6103 31462 6127
rect 31140 6098 31462 6103
rect 31103 6094 31462 6098
rect 31529 6124 31740 6130
rect 31529 6122 31690 6124
rect 31529 6102 31540 6122
rect 31560 6102 31690 6122
rect 31529 6095 31690 6102
rect 31529 6094 31570 6095
rect 31005 6068 31041 6093
rect 30853 6041 30890 6042
rect 30949 6041 30986 6042
rect 31005 6041 31012 6068
rect 30753 6032 30891 6041
rect 29511 5498 29573 6014
rect 30753 6012 30862 6032
rect 30882 6012 30891 6032
rect 30753 6005 30891 6012
rect 30949 6038 31012 6041
rect 31033 6041 31041 6068
rect 31060 6041 31097 6042
rect 31033 6038 31097 6041
rect 30949 6032 31097 6038
rect 30949 6012 30958 6032
rect 30978 6012 31068 6032
rect 31088 6012 31097 6032
rect 30753 6003 30849 6005
rect 30949 6002 31097 6012
rect 31156 6032 31193 6042
rect 31268 6041 31305 6042
rect 31249 6039 31305 6041
rect 31156 6012 31164 6032
rect 31184 6012 31193 6032
rect 31005 6001 31041 6002
rect 30853 5870 30890 5871
rect 31156 5870 31193 6012
rect 31218 6032 31305 6039
rect 31218 6029 31276 6032
rect 31218 6009 31223 6029
rect 31244 6012 31276 6029
rect 31296 6012 31305 6032
rect 31244 6009 31305 6012
rect 31218 6002 31305 6009
rect 31364 6032 31401 6042
rect 31364 6012 31372 6032
rect 31392 6012 31401 6032
rect 31218 6001 31249 6002
rect 31364 5933 31401 6012
rect 31431 6041 31462 6094
rect 31675 6087 31690 6095
rect 31730 6087 31740 6124
rect 32931 6113 32996 6252
rect 33271 6197 33308 6276
rect 33349 6263 33459 6276
rect 33423 6207 33454 6208
rect 33271 6177 33280 6197
rect 33300 6177 33308 6197
rect 31675 6078 31740 6087
rect 31888 6085 31953 6106
rect 31888 6067 31913 6085
rect 31931 6067 31953 6085
rect 32931 6095 32954 6113
rect 32972 6095 32996 6113
rect 32931 6078 32996 6095
rect 33151 6159 33219 6172
rect 33271 6167 33308 6177
rect 33367 6197 33454 6207
rect 33367 6177 33376 6197
rect 33396 6177 33454 6197
rect 33367 6168 33454 6177
rect 33367 6167 33404 6168
rect 33151 6117 33158 6159
rect 33207 6117 33219 6159
rect 33151 6114 33219 6117
rect 33423 6115 33454 6168
rect 33484 6197 33521 6276
rect 33636 6207 33667 6208
rect 33484 6177 33493 6197
rect 33513 6177 33521 6197
rect 33484 6167 33521 6177
rect 33580 6200 33667 6207
rect 33580 6197 33641 6200
rect 33580 6177 33589 6197
rect 33609 6180 33641 6197
rect 33662 6180 33667 6200
rect 33609 6177 33667 6180
rect 33580 6170 33667 6177
rect 33692 6197 33729 6339
rect 33995 6338 34032 6339
rect 34740 6336 35156 6341
rect 34740 6335 35081 6336
rect 34397 6304 34507 6318
rect 34397 6301 34440 6304
rect 34397 6296 34401 6301
rect 34319 6274 34401 6296
rect 34430 6274 34440 6301
rect 34468 6277 34475 6304
rect 34504 6296 34507 6304
rect 34504 6277 34569 6296
rect 34468 6274 34569 6277
rect 34319 6272 34569 6274
rect 33844 6207 33880 6208
rect 33692 6177 33701 6197
rect 33721 6177 33729 6197
rect 33580 6168 33636 6170
rect 33580 6167 33617 6168
rect 33692 6167 33729 6177
rect 33788 6197 33936 6207
rect 34036 6204 34132 6206
rect 33788 6177 33797 6197
rect 33817 6177 33907 6197
rect 33927 6177 33936 6197
rect 33788 6171 33936 6177
rect 33788 6168 33852 6171
rect 33788 6167 33825 6168
rect 33844 6141 33852 6168
rect 33873 6168 33936 6171
rect 33994 6197 34132 6204
rect 33994 6177 34003 6197
rect 34023 6177 34132 6197
rect 33994 6168 34132 6177
rect 34319 6193 34356 6272
rect 34397 6259 34507 6272
rect 34471 6203 34502 6204
rect 34319 6173 34328 6193
rect 34348 6173 34356 6193
rect 33873 6141 33880 6168
rect 33899 6167 33936 6168
rect 33995 6167 34032 6168
rect 33844 6116 33880 6141
rect 33315 6114 33356 6115
rect 33151 6107 33356 6114
rect 33151 6096 33325 6107
rect 31481 6041 31518 6042
rect 31431 6032 31518 6041
rect 31431 6012 31489 6032
rect 31509 6012 31518 6032
rect 31431 6002 31518 6012
rect 31577 6032 31614 6042
rect 31577 6012 31585 6032
rect 31605 6012 31614 6032
rect 31431 6001 31462 6002
rect 31426 5933 31536 5946
rect 31577 5933 31614 6012
rect 31888 5991 31953 6067
rect 33151 6063 33159 6096
rect 33152 6054 33159 6063
rect 33208 6087 33325 6096
rect 33345 6087 33356 6107
rect 33208 6079 33356 6087
rect 33423 6111 33782 6115
rect 33423 6106 33745 6111
rect 33423 6082 33536 6106
rect 33560 6087 33745 6106
rect 33769 6087 33782 6111
rect 33560 6082 33782 6087
rect 33423 6079 33782 6082
rect 33844 6079 33879 6116
rect 33947 6113 34047 6116
rect 33947 6109 34014 6113
rect 33947 6083 33959 6109
rect 33985 6087 34014 6109
rect 34040 6087 34047 6113
rect 33985 6083 34047 6087
rect 33947 6079 34047 6083
rect 33208 6063 33219 6079
rect 33208 6054 33216 6063
rect 33423 6058 33454 6079
rect 33844 6058 33880 6079
rect 33266 6057 33303 6058
rect 32931 6014 32996 6033
rect 32931 5996 32956 6014
rect 32974 5996 32996 6014
rect 31364 5931 31614 5933
rect 31364 5928 31465 5931
rect 31364 5909 31429 5928
rect 31426 5901 31429 5909
rect 31458 5901 31465 5928
rect 31493 5904 31503 5931
rect 31532 5909 31614 5931
rect 31637 5956 31954 5991
rect 31532 5904 31536 5909
rect 31493 5901 31536 5904
rect 31426 5887 31536 5901
rect 30852 5869 31193 5870
rect 30777 5867 31193 5869
rect 31637 5867 31677 5956
rect 31888 5929 31953 5956
rect 31888 5911 31911 5929
rect 31929 5911 31953 5929
rect 31888 5891 31953 5911
rect 30774 5864 31677 5867
rect 30774 5844 30780 5864
rect 30800 5844 31677 5864
rect 30774 5840 31677 5844
rect 31637 5837 31677 5840
rect 31889 5830 31954 5851
rect 30107 5822 30768 5823
rect 30107 5815 31041 5822
rect 30107 5814 31013 5815
rect 30107 5794 30958 5814
rect 30990 5795 31013 5814
rect 31038 5795 31041 5815
rect 30990 5794 31041 5795
rect 30107 5787 31041 5794
rect 29706 5745 29874 5746
rect 30109 5745 30148 5787
rect 30937 5785 31041 5787
rect 31006 5783 31041 5785
rect 31889 5812 31913 5830
rect 31931 5812 31954 5830
rect 31889 5765 31954 5812
rect 29706 5719 30150 5745
rect 29706 5717 29874 5719
rect 29508 5414 29577 5498
rect 29506 4935 29577 5414
rect 29706 5366 29733 5717
rect 30109 5713 30150 5719
rect 29773 5506 29837 5518
rect 30113 5514 30150 5713
rect 30612 5740 30684 5757
rect 30612 5701 30620 5740
rect 30665 5701 30684 5740
rect 30378 5603 30489 5618
rect 30378 5601 30420 5603
rect 30378 5581 30385 5601
rect 30404 5581 30420 5601
rect 30378 5573 30420 5581
rect 30448 5601 30489 5603
rect 30448 5581 30462 5601
rect 30481 5581 30489 5601
rect 30448 5573 30489 5581
rect 30378 5567 30489 5573
rect 30321 5545 30570 5567
rect 30321 5514 30358 5545
rect 30534 5543 30570 5545
rect 30534 5514 30571 5543
rect 29773 5505 29808 5506
rect 29750 5500 29808 5505
rect 29750 5480 29753 5500
rect 29773 5486 29808 5500
rect 29828 5486 29837 5506
rect 29773 5478 29837 5486
rect 29799 5477 29837 5478
rect 29800 5476 29837 5477
rect 29903 5510 29939 5511
rect 30011 5510 30047 5511
rect 29903 5502 30047 5510
rect 29903 5482 29911 5502
rect 29931 5482 30019 5502
rect 30039 5482 30047 5502
rect 29903 5476 30047 5482
rect 30113 5506 30151 5514
rect 30219 5510 30255 5511
rect 30113 5486 30122 5506
rect 30142 5486 30151 5506
rect 30113 5477 30151 5486
rect 30170 5503 30255 5510
rect 30170 5483 30177 5503
rect 30198 5502 30255 5503
rect 30198 5483 30227 5502
rect 30170 5482 30227 5483
rect 30247 5482 30255 5502
rect 30113 5476 30150 5477
rect 30170 5476 30255 5482
rect 30321 5506 30359 5514
rect 30432 5510 30468 5511
rect 30321 5486 30330 5506
rect 30350 5486 30359 5506
rect 30321 5477 30359 5486
rect 30383 5502 30468 5510
rect 30383 5482 30440 5502
rect 30460 5482 30468 5502
rect 30321 5476 30358 5477
rect 30383 5476 30468 5482
rect 30534 5506 30572 5514
rect 30534 5486 30543 5506
rect 30563 5486 30572 5506
rect 30534 5477 30572 5486
rect 30612 5491 30684 5701
rect 30754 5735 31954 5765
rect 30754 5734 31198 5735
rect 30754 5732 30922 5734
rect 30612 5477 30695 5491
rect 30534 5476 30571 5477
rect 29957 5455 29993 5476
rect 30383 5455 30414 5476
rect 30612 5455 30629 5477
rect 29790 5451 29890 5455
rect 29790 5447 29852 5451
rect 29790 5421 29797 5447
rect 29823 5425 29852 5447
rect 29878 5425 29890 5451
rect 29823 5421 29890 5425
rect 29790 5418 29890 5421
rect 29958 5418 29993 5455
rect 30055 5452 30414 5455
rect 30055 5447 30277 5452
rect 30055 5423 30068 5447
rect 30092 5428 30277 5447
rect 30301 5428 30414 5452
rect 30092 5423 30414 5428
rect 30055 5419 30414 5423
rect 30481 5447 30629 5455
rect 30481 5427 30492 5447
rect 30512 5444 30629 5447
rect 30682 5444 30695 5477
rect 30512 5427 30695 5444
rect 30481 5420 30695 5427
rect 30481 5419 30522 5420
rect 30612 5419 30695 5420
rect 29957 5393 29993 5418
rect 29805 5366 29842 5367
rect 29901 5366 29938 5367
rect 29957 5366 29964 5393
rect 29705 5357 29843 5366
rect 29705 5337 29814 5357
rect 29834 5337 29843 5357
rect 29705 5330 29843 5337
rect 29901 5363 29964 5366
rect 29985 5366 29993 5393
rect 30012 5366 30049 5367
rect 29985 5363 30049 5366
rect 29901 5357 30049 5363
rect 29901 5337 29910 5357
rect 29930 5337 30020 5357
rect 30040 5337 30049 5357
rect 29705 5328 29801 5330
rect 29901 5327 30049 5337
rect 30108 5357 30145 5367
rect 30220 5366 30257 5367
rect 30201 5364 30257 5366
rect 30108 5337 30116 5357
rect 30136 5337 30145 5357
rect 29957 5326 29993 5327
rect 29805 5195 29842 5196
rect 30108 5195 30145 5337
rect 30170 5357 30257 5364
rect 30170 5354 30228 5357
rect 30170 5334 30175 5354
rect 30196 5337 30228 5354
rect 30248 5337 30257 5357
rect 30196 5334 30257 5337
rect 30170 5327 30257 5334
rect 30316 5357 30353 5367
rect 30316 5337 30324 5357
rect 30344 5337 30353 5357
rect 30170 5326 30201 5327
rect 30316 5258 30353 5337
rect 30383 5366 30414 5419
rect 30620 5386 30634 5419
rect 30687 5386 30695 5419
rect 30620 5380 30695 5386
rect 30620 5375 30690 5380
rect 30433 5366 30470 5367
rect 30383 5357 30470 5366
rect 30383 5337 30441 5357
rect 30461 5337 30470 5357
rect 30383 5327 30470 5337
rect 30529 5357 30566 5367
rect 30754 5362 30781 5732
rect 30821 5502 30885 5514
rect 31161 5510 31198 5734
rect 31669 5715 31733 5717
rect 31665 5703 31733 5715
rect 31665 5670 31676 5703
rect 31716 5670 31733 5703
rect 31665 5660 31733 5670
rect 31426 5599 31537 5614
rect 31426 5597 31468 5599
rect 31426 5577 31433 5597
rect 31452 5577 31468 5597
rect 31426 5569 31468 5577
rect 31496 5597 31537 5599
rect 31496 5577 31510 5597
rect 31529 5577 31537 5597
rect 31496 5569 31537 5577
rect 31426 5563 31537 5569
rect 31369 5541 31618 5563
rect 31369 5510 31406 5541
rect 31582 5539 31618 5541
rect 31582 5510 31619 5539
rect 30821 5501 30856 5502
rect 30798 5496 30856 5501
rect 30798 5476 30801 5496
rect 30821 5482 30856 5496
rect 30876 5482 30885 5502
rect 30821 5474 30885 5482
rect 30847 5473 30885 5474
rect 30848 5472 30885 5473
rect 30951 5506 30987 5507
rect 31059 5506 31095 5507
rect 30951 5498 31095 5506
rect 30951 5478 30959 5498
rect 30979 5478 31067 5498
rect 31087 5478 31095 5498
rect 30951 5472 31095 5478
rect 31161 5502 31199 5510
rect 31267 5506 31303 5507
rect 31161 5482 31170 5502
rect 31190 5482 31199 5502
rect 31161 5473 31199 5482
rect 31218 5499 31303 5506
rect 31218 5479 31225 5499
rect 31246 5498 31303 5499
rect 31246 5479 31275 5498
rect 31218 5478 31275 5479
rect 31295 5478 31303 5498
rect 31161 5472 31198 5473
rect 31218 5472 31303 5478
rect 31369 5502 31407 5510
rect 31480 5506 31516 5507
rect 31369 5482 31378 5502
rect 31398 5482 31407 5502
rect 31369 5473 31407 5482
rect 31431 5498 31516 5506
rect 31431 5478 31488 5498
rect 31508 5478 31516 5498
rect 31369 5472 31406 5473
rect 31431 5472 31516 5478
rect 31582 5502 31620 5510
rect 31582 5482 31591 5502
rect 31611 5482 31620 5502
rect 31582 5473 31620 5482
rect 31669 5476 31733 5660
rect 31889 5534 31954 5735
rect 32931 5795 32996 5996
rect 33152 5870 33216 6054
rect 33265 6048 33303 6057
rect 33265 6028 33274 6048
rect 33294 6028 33303 6048
rect 33265 6020 33303 6028
rect 33369 6052 33454 6058
rect 33479 6057 33516 6058
rect 33369 6032 33377 6052
rect 33397 6032 33454 6052
rect 33369 6024 33454 6032
rect 33478 6048 33516 6057
rect 33478 6028 33487 6048
rect 33507 6028 33516 6048
rect 33369 6023 33405 6024
rect 33478 6020 33516 6028
rect 33582 6052 33667 6058
rect 33687 6057 33724 6058
rect 33582 6032 33590 6052
rect 33610 6051 33667 6052
rect 33610 6032 33639 6051
rect 33582 6031 33639 6032
rect 33660 6031 33667 6051
rect 33582 6024 33667 6031
rect 33686 6048 33724 6057
rect 33686 6028 33695 6048
rect 33715 6028 33724 6048
rect 33582 6023 33618 6024
rect 33686 6020 33724 6028
rect 33790 6052 33934 6058
rect 33790 6032 33798 6052
rect 33818 6032 33906 6052
rect 33926 6032 33934 6052
rect 33790 6024 33934 6032
rect 33790 6023 33826 6024
rect 33898 6023 33934 6024
rect 34000 6057 34037 6058
rect 34000 6056 34038 6057
rect 34000 6048 34064 6056
rect 34000 6028 34009 6048
rect 34029 6034 34064 6048
rect 34084 6034 34087 6054
rect 34029 6029 34087 6034
rect 34029 6028 34064 6029
rect 33266 5991 33303 6020
rect 33267 5989 33303 5991
rect 33479 5989 33516 6020
rect 33267 5967 33516 5989
rect 33348 5961 33459 5967
rect 33348 5953 33389 5961
rect 33348 5933 33356 5953
rect 33375 5933 33389 5953
rect 33348 5931 33389 5933
rect 33417 5953 33459 5961
rect 33417 5933 33433 5953
rect 33452 5933 33459 5953
rect 33417 5931 33459 5933
rect 33348 5916 33459 5931
rect 33152 5860 33220 5870
rect 33152 5827 33169 5860
rect 33209 5827 33220 5860
rect 33152 5815 33220 5827
rect 33152 5813 33216 5815
rect 33687 5796 33724 6020
rect 34000 6016 34064 6028
rect 34104 5798 34131 6168
rect 34319 6163 34356 6173
rect 34415 6193 34502 6203
rect 34415 6173 34424 6193
rect 34444 6173 34502 6193
rect 34415 6164 34502 6173
rect 34415 6163 34452 6164
rect 34195 6150 34265 6155
rect 34190 6144 34265 6150
rect 34190 6111 34198 6144
rect 34251 6111 34265 6144
rect 34471 6111 34502 6164
rect 34532 6193 34569 6272
rect 34684 6203 34715 6204
rect 34532 6173 34541 6193
rect 34561 6173 34569 6193
rect 34532 6163 34569 6173
rect 34628 6196 34715 6203
rect 34628 6193 34689 6196
rect 34628 6173 34637 6193
rect 34657 6176 34689 6193
rect 34710 6176 34715 6196
rect 34657 6173 34715 6176
rect 34628 6166 34715 6173
rect 34740 6193 34777 6335
rect 35043 6334 35080 6335
rect 34892 6203 34928 6204
rect 34740 6173 34749 6193
rect 34769 6173 34777 6193
rect 34628 6164 34684 6166
rect 34628 6163 34665 6164
rect 34740 6163 34777 6173
rect 34836 6193 34984 6203
rect 35084 6200 35180 6202
rect 34836 6173 34845 6193
rect 34865 6173 34955 6193
rect 34975 6173 34984 6193
rect 34836 6167 34984 6173
rect 34836 6164 34900 6167
rect 34836 6163 34873 6164
rect 34892 6137 34900 6164
rect 34921 6164 34984 6167
rect 35042 6193 35180 6200
rect 35042 6173 35051 6193
rect 35071 6173 35180 6193
rect 35042 6164 35180 6173
rect 34921 6137 34928 6164
rect 34947 6163 34984 6164
rect 35043 6163 35080 6164
rect 34892 6112 34928 6137
rect 34190 6110 34273 6111
rect 34363 6110 34404 6111
rect 34190 6103 34404 6110
rect 34190 6086 34373 6103
rect 34190 6053 34203 6086
rect 34256 6083 34373 6086
rect 34393 6083 34404 6103
rect 34256 6075 34404 6083
rect 34471 6107 34830 6111
rect 34471 6102 34793 6107
rect 34471 6078 34584 6102
rect 34608 6083 34793 6102
rect 34817 6083 34830 6107
rect 34608 6078 34830 6083
rect 34471 6075 34830 6078
rect 34892 6075 34927 6112
rect 34995 6109 35095 6112
rect 34995 6105 35062 6109
rect 34995 6079 35007 6105
rect 35033 6083 35062 6105
rect 35088 6083 35095 6109
rect 35033 6079 35095 6083
rect 34995 6075 35095 6079
rect 34256 6053 34273 6075
rect 34471 6054 34502 6075
rect 34892 6054 34928 6075
rect 34314 6053 34351 6054
rect 34190 6039 34273 6053
rect 33963 5796 34131 5798
rect 33687 5795 34131 5796
rect 32931 5765 34131 5795
rect 34201 5829 34273 6039
rect 34313 6044 34351 6053
rect 34313 6024 34322 6044
rect 34342 6024 34351 6044
rect 34313 6016 34351 6024
rect 34417 6048 34502 6054
rect 34527 6053 34564 6054
rect 34417 6028 34425 6048
rect 34445 6028 34502 6048
rect 34417 6020 34502 6028
rect 34526 6044 34564 6053
rect 34526 6024 34535 6044
rect 34555 6024 34564 6044
rect 34417 6019 34453 6020
rect 34526 6016 34564 6024
rect 34630 6048 34715 6054
rect 34735 6053 34772 6054
rect 34630 6028 34638 6048
rect 34658 6047 34715 6048
rect 34658 6028 34687 6047
rect 34630 6027 34687 6028
rect 34708 6027 34715 6047
rect 34630 6020 34715 6027
rect 34734 6044 34772 6053
rect 34734 6024 34743 6044
rect 34763 6024 34772 6044
rect 34630 6019 34666 6020
rect 34734 6016 34772 6024
rect 34838 6048 34982 6054
rect 34838 6028 34846 6048
rect 34866 6028 34954 6048
rect 34974 6028 34982 6048
rect 34838 6020 34982 6028
rect 34838 6019 34874 6020
rect 34946 6019 34982 6020
rect 35048 6053 35085 6054
rect 35048 6052 35086 6053
rect 35048 6044 35112 6052
rect 35048 6024 35057 6044
rect 35077 6030 35112 6044
rect 35132 6030 35135 6050
rect 35077 6025 35135 6030
rect 35077 6024 35112 6025
rect 34314 5987 34351 6016
rect 34315 5985 34351 5987
rect 34527 5985 34564 6016
rect 34315 5963 34564 5985
rect 34396 5957 34507 5963
rect 34396 5949 34437 5957
rect 34396 5929 34404 5949
rect 34423 5929 34437 5949
rect 34396 5927 34437 5929
rect 34465 5949 34507 5957
rect 34465 5929 34481 5949
rect 34500 5929 34507 5949
rect 34465 5927 34507 5929
rect 34396 5912 34507 5927
rect 34201 5790 34220 5829
rect 34265 5790 34273 5829
rect 34201 5773 34273 5790
rect 34735 5817 34772 6016
rect 35048 6012 35112 6024
rect 34735 5811 34776 5817
rect 35152 5813 35179 6164
rect 35302 6034 35381 6634
rect 35478 6182 35557 6767
rect 35761 6754 35798 6783
rect 35762 6752 35798 6754
rect 35974 6752 36011 6783
rect 35762 6730 36011 6752
rect 35843 6724 35954 6730
rect 35843 6716 35884 6724
rect 35843 6696 35851 6716
rect 35870 6696 35884 6716
rect 35843 6694 35884 6696
rect 35912 6716 35954 6724
rect 35912 6696 35928 6716
rect 35947 6696 35954 6716
rect 35912 6694 35954 6696
rect 35843 6679 35954 6694
rect 36182 6668 36219 6783
rect 36175 6556 36222 6668
rect 36343 6628 36373 6787
rect 36393 6786 36429 6787
rect 36495 6820 36532 6821
rect 36495 6819 36533 6820
rect 36495 6811 36559 6819
rect 36495 6791 36504 6811
rect 36524 6797 36559 6811
rect 36579 6797 36582 6817
rect 36524 6792 36582 6797
rect 36524 6791 36559 6792
rect 36495 6779 36559 6791
rect 36343 6624 36429 6628
rect 36343 6606 36358 6624
rect 36410 6606 36429 6624
rect 36343 6597 36429 6606
rect 36599 6558 36626 6931
rect 36458 6556 36626 6558
rect 36175 6530 36626 6556
rect 36175 6452 36222 6530
rect 36458 6529 36626 6530
rect 36120 6451 36222 6452
rect 36119 6443 36222 6451
rect 36119 6440 36171 6443
rect 36119 6405 36127 6440
rect 36152 6405 36171 6440
rect 36196 6405 36222 6443
rect 36119 6399 36222 6405
rect 36382 6444 36418 6448
rect 36382 6421 36390 6444
rect 36414 6421 36418 6444
rect 36382 6400 36418 6421
rect 36119 6395 36218 6399
rect 36382 6377 36390 6400
rect 36414 6377 36418 6400
rect 35011 5811 35179 5813
rect 34735 5785 35179 5811
rect 32931 5718 32996 5765
rect 32931 5700 32954 5718
rect 32972 5700 32996 5718
rect 33844 5745 33879 5747
rect 33844 5743 33948 5745
rect 34737 5743 34776 5785
rect 35011 5784 35179 5785
rect 33844 5736 34778 5743
rect 33844 5735 33895 5736
rect 33844 5715 33847 5735
rect 33872 5716 33895 5735
rect 33927 5716 34778 5736
rect 33872 5715 34778 5716
rect 33844 5708 34778 5715
rect 34117 5707 34778 5708
rect 32931 5679 32996 5700
rect 33208 5690 33248 5693
rect 33208 5686 34111 5690
rect 33208 5666 34085 5686
rect 34105 5666 34111 5686
rect 33208 5663 34111 5666
rect 32932 5619 32997 5639
rect 32932 5601 32956 5619
rect 32974 5601 32997 5619
rect 32932 5574 32997 5601
rect 33208 5574 33248 5663
rect 33692 5661 34108 5663
rect 33692 5660 34033 5661
rect 33349 5629 33459 5643
rect 33349 5626 33392 5629
rect 33349 5621 33353 5626
rect 32931 5539 33248 5574
rect 33271 5599 33353 5621
rect 33382 5599 33392 5626
rect 33420 5602 33427 5629
rect 33456 5621 33459 5629
rect 33456 5602 33521 5621
rect 33420 5599 33521 5602
rect 33271 5597 33521 5599
rect 31889 5516 31911 5534
rect 31929 5516 31954 5534
rect 31889 5497 31954 5516
rect 31582 5472 31619 5473
rect 31005 5451 31041 5472
rect 31431 5451 31462 5472
rect 31669 5467 31677 5476
rect 31666 5451 31677 5467
rect 30838 5447 30938 5451
rect 30838 5443 30900 5447
rect 30838 5417 30845 5443
rect 30871 5421 30900 5443
rect 30926 5421 30938 5447
rect 30871 5417 30938 5421
rect 30838 5414 30938 5417
rect 31006 5414 31041 5451
rect 31103 5448 31462 5451
rect 31103 5443 31325 5448
rect 31103 5419 31116 5443
rect 31140 5424 31325 5443
rect 31349 5424 31462 5448
rect 31140 5419 31462 5424
rect 31103 5415 31462 5419
rect 31529 5443 31677 5451
rect 31529 5423 31540 5443
rect 31560 5434 31677 5443
rect 31726 5467 31733 5476
rect 31726 5434 31734 5467
rect 32932 5463 32997 5539
rect 33271 5518 33308 5597
rect 33349 5584 33459 5597
rect 33423 5528 33454 5529
rect 33271 5498 33280 5518
rect 33300 5498 33308 5518
rect 33271 5488 33308 5498
rect 33367 5518 33454 5528
rect 33367 5498 33376 5518
rect 33396 5498 33454 5518
rect 33367 5489 33454 5498
rect 33367 5488 33404 5489
rect 31560 5423 31734 5434
rect 31529 5416 31734 5423
rect 31529 5415 31570 5416
rect 31005 5389 31041 5414
rect 30853 5362 30890 5363
rect 30949 5362 30986 5363
rect 31005 5362 31012 5389
rect 30529 5337 30537 5357
rect 30557 5337 30566 5357
rect 30383 5326 30414 5327
rect 30378 5258 30488 5271
rect 30529 5258 30566 5337
rect 30753 5353 30891 5362
rect 30753 5333 30862 5353
rect 30882 5333 30891 5353
rect 30753 5326 30891 5333
rect 30949 5359 31012 5362
rect 31033 5362 31041 5389
rect 31060 5362 31097 5363
rect 31033 5359 31097 5362
rect 30949 5353 31097 5359
rect 30949 5333 30958 5353
rect 30978 5333 31068 5353
rect 31088 5333 31097 5353
rect 30753 5324 30849 5326
rect 30949 5323 31097 5333
rect 31156 5353 31193 5363
rect 31268 5362 31305 5363
rect 31249 5360 31305 5362
rect 31156 5333 31164 5353
rect 31184 5333 31193 5353
rect 31005 5322 31041 5323
rect 30316 5256 30566 5258
rect 30316 5253 30417 5256
rect 30316 5234 30381 5253
rect 30378 5226 30381 5234
rect 30410 5226 30417 5253
rect 30445 5229 30455 5256
rect 30484 5234 30566 5256
rect 30484 5229 30488 5234
rect 30445 5226 30488 5229
rect 30378 5212 30488 5226
rect 29804 5194 30145 5195
rect 29729 5189 30145 5194
rect 30853 5191 30890 5192
rect 31156 5191 31193 5333
rect 31218 5353 31305 5360
rect 31218 5350 31276 5353
rect 31218 5330 31223 5350
rect 31244 5333 31276 5350
rect 31296 5333 31305 5353
rect 31244 5330 31305 5333
rect 31218 5323 31305 5330
rect 31364 5353 31401 5363
rect 31364 5333 31372 5353
rect 31392 5333 31401 5353
rect 31218 5322 31249 5323
rect 31364 5254 31401 5333
rect 31431 5362 31462 5415
rect 31666 5413 31734 5416
rect 31666 5371 31678 5413
rect 31727 5371 31734 5413
rect 31481 5362 31518 5363
rect 31431 5353 31518 5362
rect 31431 5333 31489 5353
rect 31509 5333 31518 5353
rect 31431 5323 31518 5333
rect 31577 5353 31614 5363
rect 31666 5358 31734 5371
rect 31889 5435 31954 5452
rect 31889 5417 31913 5435
rect 31931 5417 31954 5435
rect 32932 5445 32954 5463
rect 32972 5445 32997 5463
rect 32932 5424 32997 5445
rect 33145 5443 33210 5452
rect 31577 5333 31585 5353
rect 31605 5333 31614 5353
rect 31431 5322 31462 5323
rect 31426 5254 31536 5267
rect 31577 5254 31614 5333
rect 31889 5278 31954 5417
rect 33145 5406 33155 5443
rect 33195 5435 33210 5443
rect 33423 5436 33454 5489
rect 33484 5518 33521 5597
rect 33636 5528 33667 5529
rect 33484 5498 33493 5518
rect 33513 5498 33521 5518
rect 33484 5488 33521 5498
rect 33580 5521 33667 5528
rect 33580 5518 33641 5521
rect 33580 5498 33589 5518
rect 33609 5501 33641 5518
rect 33662 5501 33667 5521
rect 33609 5498 33667 5501
rect 33580 5491 33667 5498
rect 33692 5518 33729 5660
rect 33995 5659 34032 5660
rect 33844 5528 33880 5529
rect 33692 5498 33701 5518
rect 33721 5498 33729 5518
rect 33580 5489 33636 5491
rect 33580 5488 33617 5489
rect 33692 5488 33729 5498
rect 33788 5518 33936 5528
rect 34036 5525 34132 5527
rect 33788 5498 33797 5518
rect 33817 5498 33907 5518
rect 33927 5498 33936 5518
rect 33788 5492 33936 5498
rect 33788 5489 33852 5492
rect 33788 5488 33825 5489
rect 33844 5462 33852 5489
rect 33873 5489 33936 5492
rect 33994 5518 34132 5525
rect 33994 5498 34003 5518
rect 34023 5498 34132 5518
rect 33994 5489 34132 5498
rect 33873 5462 33880 5489
rect 33899 5488 33936 5489
rect 33995 5488 34032 5489
rect 33844 5437 33880 5462
rect 33315 5435 33356 5436
rect 33195 5428 33356 5435
rect 33195 5408 33325 5428
rect 33345 5408 33356 5428
rect 33195 5406 33356 5408
rect 33145 5400 33356 5406
rect 33423 5432 33782 5436
rect 33423 5427 33745 5432
rect 33423 5403 33536 5427
rect 33560 5408 33745 5427
rect 33769 5408 33782 5432
rect 33560 5403 33782 5408
rect 33423 5400 33782 5403
rect 33844 5400 33879 5437
rect 33947 5434 34047 5437
rect 33947 5430 34014 5434
rect 33947 5404 33959 5430
rect 33985 5408 34014 5430
rect 34040 5408 34047 5434
rect 33985 5404 34047 5408
rect 33947 5400 34047 5404
rect 33145 5387 33212 5400
rect 31889 5272 31911 5278
rect 31364 5252 31614 5254
rect 31364 5249 31465 5252
rect 31364 5230 31429 5249
rect 31426 5222 31429 5230
rect 31458 5222 31465 5249
rect 31493 5225 31503 5252
rect 31532 5230 31614 5252
rect 31643 5260 31911 5272
rect 31929 5260 31954 5278
rect 31643 5237 31954 5260
rect 32937 5364 32993 5384
rect 32937 5346 32956 5364
rect 32974 5346 32993 5364
rect 31643 5236 31698 5237
rect 31532 5225 31536 5230
rect 31493 5222 31536 5225
rect 31426 5208 31536 5222
rect 30852 5190 31193 5191
rect 29729 5169 29732 5189
rect 29752 5169 30145 5189
rect 30777 5189 31193 5190
rect 31643 5189 31686 5236
rect 32937 5233 32993 5346
rect 33145 5366 33159 5387
rect 33195 5366 33212 5387
rect 33423 5379 33454 5400
rect 33844 5379 33880 5400
rect 33266 5378 33303 5379
rect 33145 5359 33212 5366
rect 33265 5369 33303 5378
rect 30777 5185 31686 5189
rect 30096 5136 30141 5169
rect 30777 5165 30780 5185
rect 30800 5165 31686 5185
rect 31154 5160 31686 5165
rect 31894 5179 31953 5201
rect 31894 5161 31913 5179
rect 31931 5161 31953 5179
rect 30942 5136 31041 5138
rect 30096 5126 31041 5136
rect 30096 5100 30964 5126
rect 30097 5099 30964 5100
rect 30942 5088 30964 5099
rect 30989 5091 31008 5126
rect 31033 5091 31041 5126
rect 30989 5088 31041 5091
rect 30942 5080 31041 5088
rect 30968 5079 31040 5080
rect 31894 5031 31953 5161
rect 32937 5104 32992 5233
rect 33145 5207 33210 5359
rect 33265 5349 33274 5369
rect 33294 5349 33303 5369
rect 33265 5341 33303 5349
rect 33369 5373 33454 5379
rect 33479 5378 33516 5379
rect 33369 5353 33377 5373
rect 33397 5353 33454 5373
rect 33369 5345 33454 5353
rect 33478 5369 33516 5378
rect 33478 5349 33487 5369
rect 33507 5349 33516 5369
rect 33369 5344 33405 5345
rect 33478 5341 33516 5349
rect 33582 5373 33667 5379
rect 33687 5378 33724 5379
rect 33582 5353 33590 5373
rect 33610 5372 33667 5373
rect 33610 5353 33639 5372
rect 33582 5352 33639 5353
rect 33660 5352 33667 5372
rect 33582 5345 33667 5352
rect 33686 5369 33724 5378
rect 33686 5349 33695 5369
rect 33715 5349 33724 5369
rect 33582 5344 33618 5345
rect 33686 5341 33724 5349
rect 33790 5373 33934 5379
rect 33790 5353 33798 5373
rect 33818 5353 33906 5373
rect 33926 5353 33934 5373
rect 33790 5345 33934 5353
rect 33790 5344 33826 5345
rect 33898 5344 33934 5345
rect 34000 5378 34037 5379
rect 34000 5377 34038 5378
rect 34000 5369 34064 5377
rect 34000 5349 34009 5369
rect 34029 5355 34064 5369
rect 34084 5355 34087 5375
rect 34029 5350 34087 5355
rect 34029 5349 34064 5350
rect 33266 5312 33303 5341
rect 33267 5310 33303 5312
rect 33479 5310 33516 5341
rect 33267 5288 33516 5310
rect 33348 5282 33459 5288
rect 33348 5274 33389 5282
rect 33348 5254 33356 5274
rect 33375 5254 33389 5274
rect 33348 5252 33389 5254
rect 33417 5274 33459 5282
rect 33417 5254 33433 5274
rect 33452 5254 33459 5274
rect 33417 5252 33459 5254
rect 33348 5237 33459 5252
rect 33687 5242 33724 5341
rect 34000 5337 34064 5349
rect 33350 5228 33454 5237
rect 33138 5197 33259 5207
rect 33138 5195 33207 5197
rect 33138 5154 33151 5195
rect 33188 5156 33207 5195
rect 33244 5156 33259 5197
rect 33188 5154 33259 5156
rect 33138 5136 33259 5154
rect 32931 5092 32992 5104
rect 33685 5092 33726 5242
rect 34104 5234 34131 5489
rect 34193 5479 34273 5490
rect 34193 5453 34210 5479
rect 34250 5453 34273 5479
rect 34193 5426 34273 5453
rect 34193 5400 34214 5426
rect 34254 5400 34273 5426
rect 34193 5381 34273 5400
rect 34193 5355 34217 5381
rect 34257 5355 34273 5381
rect 34193 5304 34273 5355
rect 32931 5089 33726 5092
rect 34105 5103 34131 5234
rect 34195 5148 34265 5304
rect 34194 5132 34270 5148
rect 34105 5089 34133 5103
rect 32931 5054 34133 5089
rect 34194 5095 34209 5132
rect 34253 5095 34270 5132
rect 34194 5075 34270 5095
rect 35308 5125 35378 6034
rect 35477 5513 35558 6182
rect 36382 6077 36418 6377
rect 36306 6048 36419 6077
rect 36306 5683 36337 6048
rect 36230 5663 36623 5683
rect 36643 5663 36646 5683
rect 36230 5658 36646 5663
rect 36230 5657 36571 5658
rect 35887 5626 35997 5640
rect 35887 5623 35930 5626
rect 35887 5618 35891 5623
rect 35809 5596 35891 5618
rect 35920 5596 35930 5623
rect 35958 5599 35965 5626
rect 35994 5618 35997 5626
rect 35994 5599 36059 5618
rect 35958 5596 36059 5599
rect 35809 5594 36059 5596
rect 35809 5515 35846 5594
rect 35887 5581 35997 5594
rect 35961 5525 35992 5526
rect 35471 5433 35570 5513
rect 35809 5495 35818 5515
rect 35838 5495 35846 5515
rect 35809 5485 35846 5495
rect 35905 5515 35992 5525
rect 35905 5495 35914 5515
rect 35934 5495 35992 5515
rect 35905 5486 35992 5495
rect 35905 5485 35942 5486
rect 35961 5433 35992 5486
rect 36022 5515 36059 5594
rect 36174 5525 36205 5526
rect 36022 5495 36031 5515
rect 36051 5495 36059 5515
rect 36022 5485 36059 5495
rect 36118 5518 36205 5525
rect 36118 5515 36179 5518
rect 36118 5495 36127 5515
rect 36147 5498 36179 5515
rect 36200 5498 36205 5518
rect 36147 5495 36205 5498
rect 36118 5488 36205 5495
rect 36230 5515 36267 5657
rect 36533 5656 36570 5657
rect 36382 5525 36418 5526
rect 36230 5495 36239 5515
rect 36259 5495 36267 5515
rect 36118 5486 36174 5488
rect 36118 5485 36155 5486
rect 36230 5485 36267 5495
rect 36326 5515 36474 5525
rect 36574 5522 36670 5524
rect 36326 5495 36335 5515
rect 36355 5495 36445 5515
rect 36465 5495 36474 5515
rect 36326 5489 36474 5495
rect 36326 5486 36390 5489
rect 36326 5485 36363 5486
rect 36382 5459 36390 5486
rect 36411 5486 36474 5489
rect 36532 5515 36670 5522
rect 36532 5495 36541 5515
rect 36561 5495 36670 5515
rect 36532 5486 36670 5495
rect 36411 5459 36418 5486
rect 36437 5485 36474 5486
rect 36533 5485 36570 5486
rect 36382 5434 36418 5459
rect 35471 5432 35811 5433
rect 35853 5432 35894 5433
rect 35471 5425 35894 5432
rect 35471 5405 35863 5425
rect 35883 5405 35894 5425
rect 35471 5397 35894 5405
rect 35961 5429 36320 5433
rect 35961 5424 36283 5429
rect 35961 5400 36074 5424
rect 36098 5405 36283 5424
rect 36307 5405 36320 5429
rect 36098 5400 36320 5405
rect 35961 5397 36320 5400
rect 36382 5397 36417 5434
rect 36485 5431 36585 5434
rect 36485 5427 36552 5431
rect 36485 5401 36497 5427
rect 36523 5405 36552 5427
rect 36578 5405 36585 5431
rect 36523 5401 36585 5405
rect 36485 5397 36585 5401
rect 35471 5393 35811 5397
rect 35308 5075 35380 5125
rect 30616 5001 30692 5025
rect 30616 4935 30628 5001
rect 30682 4935 30692 5001
rect 31160 4956 31201 4958
rect 31432 4956 31536 4958
rect 31894 4956 31955 5031
rect 32931 4979 32992 5054
rect 33350 5052 33454 5054
rect 33685 5052 33726 5054
rect 34194 5009 34204 5075
rect 34258 5009 34270 5075
rect 34194 4985 34270 5009
rect 29506 4885 29578 4935
rect 29075 4613 29411 4617
rect 28301 4609 28401 4613
rect 28301 4605 28363 4609
rect 28301 4579 28308 4605
rect 28334 4583 28363 4605
rect 28389 4583 28401 4609
rect 28334 4579 28401 4583
rect 28301 4576 28401 4579
rect 28469 4576 28504 4613
rect 28566 4610 28925 4613
rect 28566 4605 28788 4610
rect 28566 4581 28579 4605
rect 28603 4586 28788 4605
rect 28812 4586 28925 4610
rect 28603 4581 28925 4586
rect 28566 4577 28925 4581
rect 28992 4605 29411 4613
rect 28992 4585 29003 4605
rect 29023 4585 29411 4605
rect 28992 4578 29411 4585
rect 28992 4577 29033 4578
rect 29075 4577 29411 4578
rect 28468 4551 28504 4576
rect 28316 4524 28353 4525
rect 28412 4524 28449 4525
rect 28468 4524 28475 4551
rect 28216 4515 28354 4524
rect 28216 4495 28325 4515
rect 28345 4495 28354 4515
rect 28216 4488 28354 4495
rect 28412 4521 28475 4524
rect 28496 4524 28504 4551
rect 28523 4524 28560 4525
rect 28496 4521 28560 4524
rect 28412 4515 28560 4521
rect 28412 4495 28421 4515
rect 28441 4495 28531 4515
rect 28551 4495 28560 4515
rect 28216 4486 28312 4488
rect 28412 4485 28560 4495
rect 28619 4515 28656 4525
rect 28731 4524 28768 4525
rect 28712 4522 28768 4524
rect 28619 4495 28627 4515
rect 28647 4495 28656 4515
rect 28468 4484 28504 4485
rect 28316 4353 28353 4354
rect 28619 4353 28656 4495
rect 28681 4515 28768 4522
rect 28681 4512 28739 4515
rect 28681 4492 28686 4512
rect 28707 4495 28739 4512
rect 28759 4495 28768 4515
rect 28707 4492 28768 4495
rect 28681 4485 28768 4492
rect 28827 4515 28864 4525
rect 28827 4495 28835 4515
rect 28855 4495 28864 4515
rect 28681 4484 28712 4485
rect 28827 4416 28864 4495
rect 28894 4524 28925 4577
rect 29319 4541 29411 4577
rect 28944 4524 28981 4525
rect 28894 4515 28981 4524
rect 28894 4495 28952 4515
rect 28972 4495 28981 4515
rect 28894 4485 28981 4495
rect 29040 4515 29077 4525
rect 29040 4495 29048 4515
rect 29068 4495 29077 4515
rect 28894 4484 28925 4485
rect 28889 4416 28999 4429
rect 29040 4416 29077 4495
rect 28827 4414 29077 4416
rect 28827 4411 28928 4414
rect 28827 4392 28892 4411
rect 28889 4384 28892 4392
rect 28921 4384 28928 4411
rect 28956 4387 28966 4414
rect 28995 4392 29077 4414
rect 28995 4387 28999 4392
rect 28956 4384 28999 4387
rect 28889 4370 28999 4384
rect 28315 4352 28656 4353
rect 28240 4347 28656 4352
rect 28240 4327 28243 4347
rect 28263 4327 28656 4347
rect 28400 4283 28505 4286
rect 28399 4260 28505 4283
rect 27519 4258 28020 4260
rect 28161 4258 28510 4260
rect 25633 4237 25670 4258
rect 25633 4200 25644 4237
rect 25661 4200 25670 4237
rect 27519 4252 28510 4258
rect 27519 4247 28471 4252
rect 27519 4226 28430 4247
rect 28450 4231 28471 4247
rect 28491 4231 28510 4252
rect 28450 4226 28510 4231
rect 27519 4201 28510 4226
rect 27995 4200 28177 4201
rect 25633 4190 25670 4200
rect 25479 4147 25873 4167
rect 25893 4147 25896 4167
rect 25480 4142 25896 4147
rect 25480 4141 25821 4142
rect 25137 4110 25247 4124
rect 25137 4107 25180 4110
rect 25137 4102 25141 4107
rect 25059 4080 25141 4102
rect 25170 4080 25180 4107
rect 25208 4083 25215 4110
rect 25244 4102 25247 4110
rect 25244 4083 25309 4102
rect 25208 4080 25309 4083
rect 25059 4078 25309 4080
rect 25059 3999 25096 4078
rect 25137 4065 25247 4078
rect 25211 4009 25242 4010
rect 25059 3979 25068 3999
rect 25088 3979 25096 3999
rect 25059 3969 25096 3979
rect 25155 3999 25242 4009
rect 25155 3979 25164 3999
rect 25184 3979 25242 3999
rect 25155 3970 25242 3979
rect 25155 3969 25192 3970
rect 25211 3917 25242 3970
rect 25272 3999 25309 4078
rect 25424 4009 25455 4010
rect 25272 3979 25281 3999
rect 25301 3979 25309 3999
rect 25272 3969 25309 3979
rect 25368 4002 25455 4009
rect 25368 3999 25429 4002
rect 25368 3979 25377 3999
rect 25397 3982 25429 3999
rect 25450 3982 25455 4002
rect 25397 3979 25455 3982
rect 25368 3972 25455 3979
rect 25480 3999 25517 4141
rect 25783 4140 25820 4141
rect 25632 4009 25668 4010
rect 25480 3979 25489 3999
rect 25509 3979 25517 3999
rect 25368 3970 25424 3972
rect 25368 3969 25405 3970
rect 25480 3969 25517 3979
rect 25576 3999 25724 4009
rect 25824 4006 25920 4008
rect 25576 3979 25585 3999
rect 25605 3979 25695 3999
rect 25715 3979 25724 3999
rect 25576 3973 25724 3979
rect 25576 3970 25640 3973
rect 25576 3969 25613 3970
rect 25632 3943 25640 3970
rect 25661 3970 25724 3973
rect 25782 3999 25920 4006
rect 25782 3979 25791 3999
rect 25811 3979 25920 3999
rect 25782 3970 25920 3979
rect 28549 3971 28580 4327
rect 25661 3943 25668 3970
rect 25687 3969 25724 3970
rect 25783 3969 25820 3970
rect 25632 3918 25668 3943
rect 25103 3916 25144 3917
rect 25023 3911 25144 3916
rect 24974 3909 25144 3911
rect 24974 3898 25113 3909
rect 24974 3875 24997 3898
rect 25023 3889 25113 3898
rect 25133 3889 25144 3909
rect 25023 3881 25144 3889
rect 25211 3913 25570 3917
rect 25211 3908 25533 3913
rect 25211 3884 25324 3908
rect 25348 3889 25533 3908
rect 25557 3889 25570 3913
rect 25348 3884 25570 3889
rect 25211 3881 25570 3884
rect 25632 3881 25667 3918
rect 25735 3915 25835 3918
rect 25735 3911 25802 3915
rect 25735 3885 25747 3911
rect 25773 3889 25802 3911
rect 25828 3889 25835 3915
rect 25773 3885 25835 3889
rect 25735 3881 25835 3885
rect 25023 3875 25031 3881
rect 24974 3867 25031 3875
rect 25211 3860 25242 3881
rect 25632 3860 25668 3881
rect 25054 3859 25091 3860
rect 25053 3850 25091 3859
rect 25053 3830 25062 3850
rect 25082 3830 25091 3850
rect 25053 3822 25091 3830
rect 25157 3854 25242 3860
rect 25267 3859 25304 3860
rect 25157 3834 25165 3854
rect 25185 3834 25242 3854
rect 25157 3826 25242 3834
rect 25266 3850 25304 3859
rect 25266 3830 25275 3850
rect 25295 3830 25304 3850
rect 25157 3825 25193 3826
rect 25266 3822 25304 3830
rect 25370 3854 25455 3860
rect 25475 3859 25512 3860
rect 25370 3834 25378 3854
rect 25398 3853 25455 3854
rect 25398 3834 25427 3853
rect 25370 3833 25427 3834
rect 25448 3833 25455 3853
rect 25370 3826 25455 3833
rect 25474 3850 25512 3859
rect 25474 3830 25483 3850
rect 25503 3830 25512 3850
rect 25370 3825 25406 3826
rect 25474 3822 25512 3830
rect 25578 3854 25722 3860
rect 25578 3834 25586 3854
rect 25606 3834 25694 3854
rect 25714 3834 25722 3854
rect 25578 3826 25722 3834
rect 25578 3825 25614 3826
rect 25686 3825 25722 3826
rect 25788 3859 25825 3860
rect 25788 3858 25826 3859
rect 25788 3850 25852 3858
rect 25788 3830 25797 3850
rect 25817 3836 25852 3850
rect 25872 3836 25875 3856
rect 25817 3831 25875 3836
rect 25817 3830 25852 3831
rect 25054 3793 25091 3822
rect 25055 3791 25091 3793
rect 25267 3791 25304 3822
rect 25055 3769 25304 3791
rect 25136 3763 25247 3769
rect 25136 3755 25177 3763
rect 25136 3735 25144 3755
rect 25163 3735 25177 3755
rect 25136 3733 25177 3735
rect 25205 3755 25247 3763
rect 25205 3735 25221 3755
rect 25240 3735 25247 3755
rect 25205 3733 25247 3735
rect 25136 3718 25247 3733
rect 25475 3707 25512 3822
rect 25788 3818 25852 3830
rect 25468 3701 25515 3707
rect 25892 3703 25919 3970
rect 28467 3942 28580 3971
rect 25751 3701 25919 3703
rect 25468 3675 25919 3701
rect 25468 3540 25515 3675
rect 25751 3674 25919 3675
rect 28468 3633 28504 3942
rect 29328 3828 29409 4541
rect 29508 3976 29578 4885
rect 30616 4915 30692 4935
rect 30616 4878 30633 4915
rect 30677 4878 30692 4915
rect 30753 4921 31955 4956
rect 30753 4907 30781 4921
rect 30616 4862 30692 4878
rect 30621 4706 30691 4862
rect 30755 4776 30781 4907
rect 31160 4918 31955 4921
rect 30613 4655 30693 4706
rect 30613 4629 30629 4655
rect 30669 4629 30693 4655
rect 30613 4610 30693 4629
rect 30613 4584 30632 4610
rect 30672 4584 30693 4610
rect 30613 4557 30693 4584
rect 30613 4531 30636 4557
rect 30676 4531 30693 4557
rect 30613 4520 30693 4531
rect 30755 4521 30782 4776
rect 31160 4768 31201 4918
rect 31894 4906 31955 4918
rect 31627 4856 31748 4874
rect 31627 4854 31698 4856
rect 31627 4813 31642 4854
rect 31679 4815 31698 4854
rect 31735 4815 31748 4856
rect 31679 4813 31748 4815
rect 31627 4803 31748 4813
rect 31432 4773 31536 4782
rect 30822 4661 30886 4673
rect 31162 4669 31199 4768
rect 31427 4758 31538 4773
rect 31427 4756 31469 4758
rect 31427 4736 31434 4756
rect 31453 4736 31469 4756
rect 31427 4728 31469 4736
rect 31497 4756 31538 4758
rect 31497 4736 31511 4756
rect 31530 4736 31538 4756
rect 31497 4728 31538 4736
rect 31427 4722 31538 4728
rect 31370 4700 31619 4722
rect 31370 4669 31407 4700
rect 31583 4698 31619 4700
rect 31583 4669 31620 4698
rect 30822 4660 30857 4661
rect 30799 4655 30857 4660
rect 30799 4635 30802 4655
rect 30822 4641 30857 4655
rect 30877 4641 30886 4661
rect 30822 4633 30886 4641
rect 30848 4632 30886 4633
rect 30849 4631 30886 4632
rect 30952 4665 30988 4666
rect 31060 4665 31096 4666
rect 30952 4657 31096 4665
rect 30952 4637 30960 4657
rect 30980 4637 31068 4657
rect 31088 4637 31096 4657
rect 30952 4631 31096 4637
rect 31162 4661 31200 4669
rect 31268 4665 31304 4666
rect 31162 4641 31171 4661
rect 31191 4641 31200 4661
rect 31162 4632 31200 4641
rect 31219 4658 31304 4665
rect 31219 4638 31226 4658
rect 31247 4657 31304 4658
rect 31247 4638 31276 4657
rect 31219 4637 31276 4638
rect 31296 4637 31304 4657
rect 31162 4631 31199 4632
rect 31219 4631 31304 4637
rect 31370 4661 31408 4669
rect 31481 4665 31517 4666
rect 31370 4641 31379 4661
rect 31399 4641 31408 4661
rect 31370 4632 31408 4641
rect 31432 4657 31517 4665
rect 31432 4637 31489 4657
rect 31509 4637 31517 4657
rect 31370 4631 31407 4632
rect 31432 4631 31517 4637
rect 31583 4661 31621 4669
rect 31583 4641 31592 4661
rect 31612 4641 31621 4661
rect 31676 4651 31741 4803
rect 31894 4777 31949 4906
rect 32933 4849 32992 4979
rect 33846 4930 33918 4931
rect 33845 4922 33944 4930
rect 33845 4919 33897 4922
rect 33845 4884 33853 4919
rect 33878 4884 33897 4919
rect 33922 4911 33944 4922
rect 33922 4910 34789 4911
rect 33922 4884 34790 4910
rect 33845 4874 34790 4884
rect 33845 4872 33944 4874
rect 32933 4831 32955 4849
rect 32973 4831 32992 4849
rect 32933 4809 32992 4831
rect 33200 4845 33732 4850
rect 33200 4825 34086 4845
rect 34106 4825 34109 4845
rect 34745 4841 34790 4874
rect 33200 4821 34109 4825
rect 31583 4632 31621 4641
rect 31674 4644 31741 4651
rect 31583 4631 31620 4632
rect 31006 4610 31042 4631
rect 31432 4610 31463 4631
rect 31674 4623 31691 4644
rect 31727 4623 31741 4644
rect 31893 4664 31949 4777
rect 33200 4774 33243 4821
rect 33693 4820 34109 4821
rect 34741 4821 35134 4841
rect 35154 4821 35157 4841
rect 33693 4819 34034 4820
rect 33350 4788 33460 4802
rect 33350 4785 33393 4788
rect 33350 4780 33354 4785
rect 33188 4773 33243 4774
rect 31893 4646 31912 4664
rect 31930 4646 31949 4664
rect 31893 4626 31949 4646
rect 32932 4750 33243 4773
rect 32932 4732 32957 4750
rect 32975 4738 33243 4750
rect 33272 4758 33354 4780
rect 33383 4758 33393 4785
rect 33421 4761 33428 4788
rect 33457 4780 33460 4788
rect 33457 4761 33522 4780
rect 33421 4758 33522 4761
rect 33272 4756 33522 4758
rect 32975 4732 32997 4738
rect 31674 4610 31741 4623
rect 30839 4606 30939 4610
rect 30839 4602 30901 4606
rect 30839 4576 30846 4602
rect 30872 4580 30901 4602
rect 30927 4580 30939 4606
rect 30872 4576 30939 4580
rect 30839 4573 30939 4576
rect 31007 4573 31042 4610
rect 31104 4607 31463 4610
rect 31104 4602 31326 4607
rect 31104 4578 31117 4602
rect 31141 4583 31326 4602
rect 31350 4583 31463 4607
rect 31141 4578 31463 4583
rect 31104 4574 31463 4578
rect 31530 4604 31741 4610
rect 31530 4602 31691 4604
rect 31530 4582 31541 4602
rect 31561 4582 31691 4602
rect 31530 4575 31691 4582
rect 31530 4574 31571 4575
rect 31006 4548 31042 4573
rect 30854 4521 30891 4522
rect 30950 4521 30987 4522
rect 31006 4521 31013 4548
rect 30754 4512 30892 4521
rect 30754 4492 30863 4512
rect 30883 4492 30892 4512
rect 30754 4485 30892 4492
rect 30950 4518 31013 4521
rect 31034 4521 31042 4548
rect 31061 4521 31098 4522
rect 31034 4518 31098 4521
rect 30950 4512 31098 4518
rect 30950 4492 30959 4512
rect 30979 4492 31069 4512
rect 31089 4492 31098 4512
rect 30754 4483 30850 4485
rect 30950 4482 31098 4492
rect 31157 4512 31194 4522
rect 31269 4521 31306 4522
rect 31250 4519 31306 4521
rect 31157 4492 31165 4512
rect 31185 4492 31194 4512
rect 31006 4481 31042 4482
rect 30854 4350 30891 4351
rect 31157 4350 31194 4492
rect 31219 4512 31306 4519
rect 31219 4509 31277 4512
rect 31219 4489 31224 4509
rect 31245 4492 31277 4509
rect 31297 4492 31306 4512
rect 31245 4489 31306 4492
rect 31219 4482 31306 4489
rect 31365 4512 31402 4522
rect 31365 4492 31373 4512
rect 31393 4492 31402 4512
rect 31219 4481 31250 4482
rect 31365 4413 31402 4492
rect 31432 4521 31463 4574
rect 31676 4567 31691 4575
rect 31731 4567 31741 4604
rect 32932 4593 32997 4732
rect 33272 4677 33309 4756
rect 33350 4743 33460 4756
rect 33424 4687 33455 4688
rect 33272 4657 33281 4677
rect 33301 4657 33309 4677
rect 31676 4558 31741 4567
rect 31889 4565 31954 4586
rect 31889 4547 31914 4565
rect 31932 4547 31954 4565
rect 32932 4575 32955 4593
rect 32973 4575 32997 4593
rect 32932 4558 32997 4575
rect 33152 4639 33220 4652
rect 33272 4647 33309 4657
rect 33368 4677 33455 4687
rect 33368 4657 33377 4677
rect 33397 4657 33455 4677
rect 33368 4648 33455 4657
rect 33368 4647 33405 4648
rect 33152 4597 33159 4639
rect 33208 4597 33220 4639
rect 33152 4594 33220 4597
rect 33424 4595 33455 4648
rect 33485 4677 33522 4756
rect 33637 4687 33668 4688
rect 33485 4657 33494 4677
rect 33514 4657 33522 4677
rect 33485 4647 33522 4657
rect 33581 4680 33668 4687
rect 33581 4677 33642 4680
rect 33581 4657 33590 4677
rect 33610 4660 33642 4677
rect 33663 4660 33668 4680
rect 33610 4657 33668 4660
rect 33581 4650 33668 4657
rect 33693 4677 33730 4819
rect 33996 4818 34033 4819
rect 34741 4816 35157 4821
rect 34741 4815 35082 4816
rect 34398 4784 34508 4798
rect 34398 4781 34441 4784
rect 34398 4776 34402 4781
rect 34320 4754 34402 4776
rect 34431 4754 34441 4781
rect 34469 4757 34476 4784
rect 34505 4776 34508 4784
rect 34505 4757 34570 4776
rect 34469 4754 34570 4757
rect 34320 4752 34570 4754
rect 33845 4687 33881 4688
rect 33693 4657 33702 4677
rect 33722 4657 33730 4677
rect 33581 4648 33637 4650
rect 33581 4647 33618 4648
rect 33693 4647 33730 4657
rect 33789 4677 33937 4687
rect 34037 4684 34133 4686
rect 33789 4657 33798 4677
rect 33818 4657 33908 4677
rect 33928 4657 33937 4677
rect 33789 4651 33937 4657
rect 33789 4648 33853 4651
rect 33789 4647 33826 4648
rect 33845 4621 33853 4648
rect 33874 4648 33937 4651
rect 33995 4677 34133 4684
rect 33995 4657 34004 4677
rect 34024 4657 34133 4677
rect 33995 4648 34133 4657
rect 34320 4673 34357 4752
rect 34398 4739 34508 4752
rect 34472 4683 34503 4684
rect 34320 4653 34329 4673
rect 34349 4653 34357 4673
rect 33874 4621 33881 4648
rect 33900 4647 33937 4648
rect 33996 4647 34033 4648
rect 33845 4596 33881 4621
rect 33316 4594 33357 4595
rect 33152 4587 33357 4594
rect 33152 4576 33326 4587
rect 31482 4521 31519 4522
rect 31432 4512 31519 4521
rect 31432 4492 31490 4512
rect 31510 4492 31519 4512
rect 31432 4482 31519 4492
rect 31578 4512 31615 4522
rect 31578 4492 31586 4512
rect 31606 4492 31615 4512
rect 31432 4481 31463 4482
rect 31427 4413 31537 4426
rect 31578 4413 31615 4492
rect 31889 4471 31954 4547
rect 33152 4543 33160 4576
rect 33153 4534 33160 4543
rect 33209 4567 33326 4576
rect 33346 4567 33357 4587
rect 33209 4559 33357 4567
rect 33424 4591 33783 4595
rect 33424 4586 33746 4591
rect 33424 4562 33537 4586
rect 33561 4567 33746 4586
rect 33770 4567 33783 4591
rect 33561 4562 33783 4567
rect 33424 4559 33783 4562
rect 33845 4559 33880 4596
rect 33948 4593 34048 4596
rect 33948 4589 34015 4593
rect 33948 4563 33960 4589
rect 33986 4567 34015 4589
rect 34041 4567 34048 4593
rect 33986 4563 34048 4567
rect 33948 4559 34048 4563
rect 33209 4543 33220 4559
rect 33209 4534 33217 4543
rect 33424 4538 33455 4559
rect 33845 4538 33881 4559
rect 33267 4537 33304 4538
rect 32932 4494 32997 4513
rect 32932 4476 32957 4494
rect 32975 4476 32997 4494
rect 31365 4411 31615 4413
rect 31365 4408 31466 4411
rect 31365 4389 31430 4408
rect 31427 4381 31430 4389
rect 31459 4381 31466 4408
rect 31494 4384 31504 4411
rect 31533 4389 31615 4411
rect 31638 4436 31955 4471
rect 31533 4384 31537 4389
rect 31494 4381 31537 4384
rect 31427 4367 31537 4381
rect 30853 4349 31194 4350
rect 30778 4347 31194 4349
rect 31638 4347 31678 4436
rect 31889 4409 31954 4436
rect 31889 4391 31912 4409
rect 31930 4391 31954 4409
rect 31889 4371 31954 4391
rect 30775 4344 31678 4347
rect 30775 4324 30781 4344
rect 30801 4324 31678 4344
rect 30775 4320 31678 4324
rect 31638 4317 31678 4320
rect 31890 4310 31955 4331
rect 30108 4302 30769 4303
rect 30108 4295 31042 4302
rect 30108 4294 31014 4295
rect 30108 4274 30959 4294
rect 30991 4275 31014 4294
rect 31039 4275 31042 4295
rect 30991 4274 31042 4275
rect 30108 4267 31042 4274
rect 29707 4225 29875 4226
rect 30110 4225 30149 4267
rect 30938 4265 31042 4267
rect 31007 4263 31042 4265
rect 31890 4292 31914 4310
rect 31932 4292 31955 4310
rect 31890 4245 31955 4292
rect 29707 4199 30151 4225
rect 29707 4197 29875 4199
rect 28468 3610 28472 3633
rect 28496 3610 28504 3633
rect 28668 3611 28767 3615
rect 28468 3589 28504 3610
rect 28468 3566 28472 3589
rect 28496 3566 28504 3589
rect 28468 3562 28504 3566
rect 28664 3605 28767 3611
rect 28664 3567 28690 3605
rect 28715 3570 28734 3605
rect 28759 3570 28767 3605
rect 28715 3567 28767 3570
rect 28664 3559 28767 3567
rect 28664 3558 28766 3559
rect 25466 3491 25525 3540
rect 25466 3463 25484 3491
rect 25512 3463 25525 3491
rect 25466 3453 25525 3463
rect 28260 3480 28428 3481
rect 28664 3480 28711 3558
rect 28260 3454 28711 3480
rect 28260 3452 28428 3454
rect 28260 3079 28287 3452
rect 28457 3404 28543 3413
rect 28457 3386 28476 3404
rect 28528 3386 28543 3404
rect 28457 3382 28543 3386
rect 28327 3219 28391 3231
rect 28327 3218 28362 3219
rect 28304 3213 28362 3218
rect 28304 3193 28307 3213
rect 28327 3199 28362 3213
rect 28382 3199 28391 3219
rect 28327 3191 28391 3199
rect 28353 3190 28391 3191
rect 28354 3189 28391 3190
rect 28457 3223 28493 3224
rect 28513 3223 28543 3382
rect 28664 3342 28711 3454
rect 28667 3227 28704 3342
rect 28932 3316 29043 3331
rect 28932 3314 28974 3316
rect 28932 3294 28939 3314
rect 28958 3294 28974 3314
rect 28932 3286 28974 3294
rect 29002 3314 29043 3316
rect 29002 3294 29016 3314
rect 29035 3294 29043 3314
rect 29002 3286 29043 3294
rect 28932 3280 29043 3286
rect 28875 3258 29124 3280
rect 28875 3227 28912 3258
rect 29088 3256 29124 3258
rect 29088 3227 29125 3256
rect 29329 3243 29408 3828
rect 29505 3376 29584 3976
rect 29707 3846 29734 4197
rect 30110 4193 30151 4199
rect 29774 3986 29838 3998
rect 30114 3994 30151 4193
rect 30613 4220 30685 4237
rect 30613 4181 30621 4220
rect 30666 4181 30685 4220
rect 30379 4083 30490 4098
rect 30379 4081 30421 4083
rect 30379 4061 30386 4081
rect 30405 4061 30421 4081
rect 30379 4053 30421 4061
rect 30449 4081 30490 4083
rect 30449 4061 30463 4081
rect 30482 4061 30490 4081
rect 30449 4053 30490 4061
rect 30379 4047 30490 4053
rect 30322 4025 30571 4047
rect 30322 3994 30359 4025
rect 30535 4023 30571 4025
rect 30535 3994 30572 4023
rect 29774 3985 29809 3986
rect 29751 3980 29809 3985
rect 29751 3960 29754 3980
rect 29774 3966 29809 3980
rect 29829 3966 29838 3986
rect 29774 3958 29838 3966
rect 29800 3957 29838 3958
rect 29801 3956 29838 3957
rect 29904 3990 29940 3991
rect 30012 3990 30048 3991
rect 29904 3982 30048 3990
rect 29904 3962 29912 3982
rect 29932 3962 30020 3982
rect 30040 3962 30048 3982
rect 29904 3956 30048 3962
rect 30114 3986 30152 3994
rect 30220 3990 30256 3991
rect 30114 3966 30123 3986
rect 30143 3966 30152 3986
rect 30114 3957 30152 3966
rect 30171 3983 30256 3990
rect 30171 3963 30178 3983
rect 30199 3982 30256 3983
rect 30199 3963 30228 3982
rect 30171 3962 30228 3963
rect 30248 3962 30256 3982
rect 30114 3956 30151 3957
rect 30171 3956 30256 3962
rect 30322 3986 30360 3994
rect 30433 3990 30469 3991
rect 30322 3966 30331 3986
rect 30351 3966 30360 3986
rect 30322 3957 30360 3966
rect 30384 3982 30469 3990
rect 30384 3962 30441 3982
rect 30461 3962 30469 3982
rect 30322 3956 30359 3957
rect 30384 3956 30469 3962
rect 30535 3986 30573 3994
rect 30535 3966 30544 3986
rect 30564 3966 30573 3986
rect 30535 3957 30573 3966
rect 30613 3971 30685 4181
rect 30755 4215 31955 4245
rect 30755 4214 31199 4215
rect 30755 4212 30923 4214
rect 30613 3957 30696 3971
rect 30535 3956 30572 3957
rect 29958 3935 29994 3956
rect 30384 3935 30415 3956
rect 30613 3935 30630 3957
rect 29791 3931 29891 3935
rect 29791 3927 29853 3931
rect 29791 3901 29798 3927
rect 29824 3905 29853 3927
rect 29879 3905 29891 3931
rect 29824 3901 29891 3905
rect 29791 3898 29891 3901
rect 29959 3898 29994 3935
rect 30056 3932 30415 3935
rect 30056 3927 30278 3932
rect 30056 3903 30069 3927
rect 30093 3908 30278 3927
rect 30302 3908 30415 3932
rect 30093 3903 30415 3908
rect 30056 3899 30415 3903
rect 30482 3927 30630 3935
rect 30482 3907 30493 3927
rect 30513 3924 30630 3927
rect 30683 3924 30696 3957
rect 30513 3907 30696 3924
rect 30482 3900 30696 3907
rect 30482 3899 30523 3900
rect 30613 3899 30696 3900
rect 29958 3873 29994 3898
rect 29806 3846 29843 3847
rect 29902 3846 29939 3847
rect 29958 3846 29965 3873
rect 29706 3837 29844 3846
rect 29706 3817 29815 3837
rect 29835 3817 29844 3837
rect 29706 3810 29844 3817
rect 29902 3843 29965 3846
rect 29986 3846 29994 3873
rect 30013 3846 30050 3847
rect 29986 3843 30050 3846
rect 29902 3837 30050 3843
rect 29902 3817 29911 3837
rect 29931 3817 30021 3837
rect 30041 3817 30050 3837
rect 29706 3808 29802 3810
rect 29902 3807 30050 3817
rect 30109 3837 30146 3847
rect 30221 3846 30258 3847
rect 30202 3844 30258 3846
rect 30109 3817 30117 3837
rect 30137 3817 30146 3837
rect 29958 3806 29994 3807
rect 29806 3675 29843 3676
rect 30109 3675 30146 3817
rect 30171 3837 30258 3844
rect 30171 3834 30229 3837
rect 30171 3814 30176 3834
rect 30197 3817 30229 3834
rect 30249 3817 30258 3837
rect 30197 3814 30258 3817
rect 30171 3807 30258 3814
rect 30317 3837 30354 3847
rect 30317 3817 30325 3837
rect 30345 3817 30354 3837
rect 30171 3806 30202 3807
rect 30317 3738 30354 3817
rect 30384 3846 30415 3899
rect 30621 3866 30635 3899
rect 30688 3866 30696 3899
rect 30621 3860 30696 3866
rect 30621 3855 30691 3860
rect 30434 3846 30471 3847
rect 30384 3837 30471 3846
rect 30384 3817 30442 3837
rect 30462 3817 30471 3837
rect 30384 3807 30471 3817
rect 30530 3837 30567 3847
rect 30755 3842 30782 4212
rect 30822 3982 30886 3994
rect 31162 3990 31199 4214
rect 31670 4195 31734 4197
rect 31666 4183 31734 4195
rect 31666 4150 31677 4183
rect 31717 4150 31734 4183
rect 31666 4140 31734 4150
rect 31427 4079 31538 4094
rect 31427 4077 31469 4079
rect 31427 4057 31434 4077
rect 31453 4057 31469 4077
rect 31427 4049 31469 4057
rect 31497 4077 31538 4079
rect 31497 4057 31511 4077
rect 31530 4057 31538 4077
rect 31497 4049 31538 4057
rect 31427 4043 31538 4049
rect 31370 4021 31619 4043
rect 31370 3990 31407 4021
rect 31583 4019 31619 4021
rect 31583 3990 31620 4019
rect 30822 3981 30857 3982
rect 30799 3976 30857 3981
rect 30799 3956 30802 3976
rect 30822 3962 30857 3976
rect 30877 3962 30886 3982
rect 30822 3954 30886 3962
rect 30848 3953 30886 3954
rect 30849 3952 30886 3953
rect 30952 3986 30988 3987
rect 31060 3986 31096 3987
rect 30952 3978 31096 3986
rect 30952 3958 30960 3978
rect 30980 3958 31068 3978
rect 31088 3958 31096 3978
rect 30952 3952 31096 3958
rect 31162 3982 31200 3990
rect 31268 3986 31304 3987
rect 31162 3962 31171 3982
rect 31191 3962 31200 3982
rect 31162 3953 31200 3962
rect 31219 3979 31304 3986
rect 31219 3959 31226 3979
rect 31247 3978 31304 3979
rect 31247 3959 31276 3978
rect 31219 3958 31276 3959
rect 31296 3958 31304 3978
rect 31162 3952 31199 3953
rect 31219 3952 31304 3958
rect 31370 3982 31408 3990
rect 31481 3986 31517 3987
rect 31370 3962 31379 3982
rect 31399 3962 31408 3982
rect 31370 3953 31408 3962
rect 31432 3978 31517 3986
rect 31432 3958 31489 3978
rect 31509 3958 31517 3978
rect 31370 3952 31407 3953
rect 31432 3952 31517 3958
rect 31583 3982 31621 3990
rect 31583 3962 31592 3982
rect 31612 3962 31621 3982
rect 31583 3953 31621 3962
rect 31670 3956 31734 4140
rect 31890 4014 31955 4215
rect 32932 4275 32997 4476
rect 33153 4350 33217 4534
rect 33266 4528 33304 4537
rect 33266 4508 33275 4528
rect 33295 4508 33304 4528
rect 33266 4500 33304 4508
rect 33370 4532 33455 4538
rect 33480 4537 33517 4538
rect 33370 4512 33378 4532
rect 33398 4512 33455 4532
rect 33370 4504 33455 4512
rect 33479 4528 33517 4537
rect 33479 4508 33488 4528
rect 33508 4508 33517 4528
rect 33370 4503 33406 4504
rect 33479 4500 33517 4508
rect 33583 4532 33668 4538
rect 33688 4537 33725 4538
rect 33583 4512 33591 4532
rect 33611 4531 33668 4532
rect 33611 4512 33640 4531
rect 33583 4511 33640 4512
rect 33661 4511 33668 4531
rect 33583 4504 33668 4511
rect 33687 4528 33725 4537
rect 33687 4508 33696 4528
rect 33716 4508 33725 4528
rect 33583 4503 33619 4504
rect 33687 4500 33725 4508
rect 33791 4532 33935 4538
rect 33791 4512 33799 4532
rect 33819 4512 33907 4532
rect 33927 4512 33935 4532
rect 33791 4504 33935 4512
rect 33791 4503 33827 4504
rect 33899 4503 33935 4504
rect 34001 4537 34038 4538
rect 34001 4536 34039 4537
rect 34001 4528 34065 4536
rect 34001 4508 34010 4528
rect 34030 4514 34065 4528
rect 34085 4514 34088 4534
rect 34030 4509 34088 4514
rect 34030 4508 34065 4509
rect 33267 4471 33304 4500
rect 33268 4469 33304 4471
rect 33480 4469 33517 4500
rect 33268 4447 33517 4469
rect 33349 4441 33460 4447
rect 33349 4433 33390 4441
rect 33349 4413 33357 4433
rect 33376 4413 33390 4433
rect 33349 4411 33390 4413
rect 33418 4433 33460 4441
rect 33418 4413 33434 4433
rect 33453 4413 33460 4433
rect 33418 4411 33460 4413
rect 33349 4396 33460 4411
rect 33153 4340 33221 4350
rect 33153 4307 33170 4340
rect 33210 4307 33221 4340
rect 33153 4295 33221 4307
rect 33153 4293 33217 4295
rect 33688 4276 33725 4500
rect 34001 4496 34065 4508
rect 34105 4278 34132 4648
rect 34320 4643 34357 4653
rect 34416 4673 34503 4683
rect 34416 4653 34425 4673
rect 34445 4653 34503 4673
rect 34416 4644 34503 4653
rect 34416 4643 34453 4644
rect 34196 4630 34266 4635
rect 34191 4624 34266 4630
rect 34191 4591 34199 4624
rect 34252 4591 34266 4624
rect 34472 4591 34503 4644
rect 34533 4673 34570 4752
rect 34685 4683 34716 4684
rect 34533 4653 34542 4673
rect 34562 4653 34570 4673
rect 34533 4643 34570 4653
rect 34629 4676 34716 4683
rect 34629 4673 34690 4676
rect 34629 4653 34638 4673
rect 34658 4656 34690 4673
rect 34711 4656 34716 4676
rect 34658 4653 34716 4656
rect 34629 4646 34716 4653
rect 34741 4673 34778 4815
rect 35044 4814 35081 4815
rect 34893 4683 34929 4684
rect 34741 4653 34750 4673
rect 34770 4653 34778 4673
rect 34629 4644 34685 4646
rect 34629 4643 34666 4644
rect 34741 4643 34778 4653
rect 34837 4673 34985 4683
rect 35085 4680 35181 4682
rect 34837 4653 34846 4673
rect 34866 4653 34956 4673
rect 34976 4653 34985 4673
rect 34837 4647 34985 4653
rect 34837 4644 34901 4647
rect 34837 4643 34874 4644
rect 34893 4617 34901 4644
rect 34922 4644 34985 4647
rect 35043 4673 35181 4680
rect 35043 4653 35052 4673
rect 35072 4653 35181 4673
rect 35043 4644 35181 4653
rect 34922 4617 34929 4644
rect 34948 4643 34985 4644
rect 35044 4643 35081 4644
rect 34893 4592 34929 4617
rect 34191 4590 34274 4591
rect 34364 4590 34405 4591
rect 34191 4583 34405 4590
rect 34191 4566 34374 4583
rect 34191 4533 34204 4566
rect 34257 4563 34374 4566
rect 34394 4563 34405 4583
rect 34257 4555 34405 4563
rect 34472 4587 34831 4591
rect 34472 4582 34794 4587
rect 34472 4558 34585 4582
rect 34609 4563 34794 4582
rect 34818 4563 34831 4587
rect 34609 4558 34831 4563
rect 34472 4555 34831 4558
rect 34893 4555 34928 4592
rect 34996 4589 35096 4592
rect 34996 4585 35063 4589
rect 34996 4559 35008 4585
rect 35034 4563 35063 4585
rect 35089 4563 35096 4589
rect 35034 4559 35096 4563
rect 34996 4555 35096 4559
rect 34257 4533 34274 4555
rect 34472 4534 34503 4555
rect 34893 4534 34929 4555
rect 34315 4533 34352 4534
rect 34191 4519 34274 4533
rect 33964 4276 34132 4278
rect 33688 4275 34132 4276
rect 32932 4245 34132 4275
rect 34202 4309 34274 4519
rect 34314 4524 34352 4533
rect 34314 4504 34323 4524
rect 34343 4504 34352 4524
rect 34314 4496 34352 4504
rect 34418 4528 34503 4534
rect 34528 4533 34565 4534
rect 34418 4508 34426 4528
rect 34446 4508 34503 4528
rect 34418 4500 34503 4508
rect 34527 4524 34565 4533
rect 34527 4504 34536 4524
rect 34556 4504 34565 4524
rect 34418 4499 34454 4500
rect 34527 4496 34565 4504
rect 34631 4528 34716 4534
rect 34736 4533 34773 4534
rect 34631 4508 34639 4528
rect 34659 4527 34716 4528
rect 34659 4508 34688 4527
rect 34631 4507 34688 4508
rect 34709 4507 34716 4527
rect 34631 4500 34716 4507
rect 34735 4524 34773 4533
rect 34735 4504 34744 4524
rect 34764 4504 34773 4524
rect 34631 4499 34667 4500
rect 34735 4496 34773 4504
rect 34839 4528 34983 4534
rect 34839 4508 34847 4528
rect 34867 4508 34955 4528
rect 34975 4508 34983 4528
rect 34839 4500 34983 4508
rect 34839 4499 34875 4500
rect 34947 4499 34983 4500
rect 35049 4533 35086 4534
rect 35049 4532 35087 4533
rect 35049 4524 35113 4532
rect 35049 4504 35058 4524
rect 35078 4510 35113 4524
rect 35133 4510 35136 4530
rect 35078 4505 35136 4510
rect 35078 4504 35113 4505
rect 34315 4467 34352 4496
rect 34316 4465 34352 4467
rect 34528 4465 34565 4496
rect 34316 4443 34565 4465
rect 34397 4437 34508 4443
rect 34397 4429 34438 4437
rect 34397 4409 34405 4429
rect 34424 4409 34438 4429
rect 34397 4407 34438 4409
rect 34466 4429 34508 4437
rect 34466 4409 34482 4429
rect 34501 4409 34508 4429
rect 34466 4407 34508 4409
rect 34397 4392 34508 4407
rect 34202 4270 34221 4309
rect 34266 4270 34274 4309
rect 34202 4253 34274 4270
rect 34736 4297 34773 4496
rect 35049 4492 35113 4504
rect 34736 4291 34777 4297
rect 35153 4293 35180 4644
rect 35309 4596 35380 5075
rect 35309 4512 35378 4596
rect 35012 4291 35180 4293
rect 34736 4265 35180 4291
rect 32932 4198 32997 4245
rect 32932 4180 32955 4198
rect 32973 4180 32997 4198
rect 33845 4225 33880 4227
rect 33845 4223 33949 4225
rect 34738 4223 34777 4265
rect 35012 4264 35180 4265
rect 33845 4216 34779 4223
rect 33845 4215 33896 4216
rect 33845 4195 33848 4215
rect 33873 4196 33896 4215
rect 33928 4196 34779 4216
rect 33873 4195 34779 4196
rect 33845 4188 34779 4195
rect 34118 4187 34779 4188
rect 32932 4159 32997 4180
rect 33209 4170 33249 4173
rect 33209 4166 34112 4170
rect 33209 4146 34086 4166
rect 34106 4146 34112 4166
rect 33209 4143 34112 4146
rect 32933 4099 32998 4119
rect 32933 4081 32957 4099
rect 32975 4081 32998 4099
rect 32933 4054 32998 4081
rect 33209 4054 33249 4143
rect 33693 4141 34109 4143
rect 33693 4140 34034 4141
rect 33350 4109 33460 4123
rect 33350 4106 33393 4109
rect 33350 4101 33354 4106
rect 32932 4019 33249 4054
rect 33272 4079 33354 4101
rect 33383 4079 33393 4106
rect 33421 4082 33428 4109
rect 33457 4101 33460 4109
rect 33457 4082 33522 4101
rect 33421 4079 33522 4082
rect 33272 4077 33522 4079
rect 31890 3996 31912 4014
rect 31930 3996 31955 4014
rect 31890 3977 31955 3996
rect 31583 3952 31620 3953
rect 31006 3931 31042 3952
rect 31432 3931 31463 3952
rect 31670 3947 31678 3956
rect 31667 3931 31678 3947
rect 30839 3927 30939 3931
rect 30839 3923 30901 3927
rect 30839 3897 30846 3923
rect 30872 3901 30901 3923
rect 30927 3901 30939 3927
rect 30872 3897 30939 3901
rect 30839 3894 30939 3897
rect 31007 3894 31042 3931
rect 31104 3928 31463 3931
rect 31104 3923 31326 3928
rect 31104 3899 31117 3923
rect 31141 3904 31326 3923
rect 31350 3904 31463 3928
rect 31141 3899 31463 3904
rect 31104 3895 31463 3899
rect 31530 3923 31678 3931
rect 31530 3903 31541 3923
rect 31561 3914 31678 3923
rect 31727 3947 31734 3956
rect 31727 3914 31735 3947
rect 32933 3943 32998 4019
rect 33272 3998 33309 4077
rect 33350 4064 33460 4077
rect 33424 4008 33455 4009
rect 33272 3978 33281 3998
rect 33301 3978 33309 3998
rect 33272 3968 33309 3978
rect 33368 3998 33455 4008
rect 33368 3978 33377 3998
rect 33397 3978 33455 3998
rect 33368 3969 33455 3978
rect 33368 3968 33405 3969
rect 31561 3903 31735 3914
rect 31530 3896 31735 3903
rect 31530 3895 31571 3896
rect 31006 3869 31042 3894
rect 30854 3842 30891 3843
rect 30950 3842 30987 3843
rect 31006 3842 31013 3869
rect 30530 3817 30538 3837
rect 30558 3817 30567 3837
rect 30384 3806 30415 3807
rect 30379 3738 30489 3751
rect 30530 3738 30567 3817
rect 30754 3833 30892 3842
rect 30754 3813 30863 3833
rect 30883 3813 30892 3833
rect 30754 3806 30892 3813
rect 30950 3839 31013 3842
rect 31034 3842 31042 3869
rect 31061 3842 31098 3843
rect 31034 3839 31098 3842
rect 30950 3833 31098 3839
rect 30950 3813 30959 3833
rect 30979 3813 31069 3833
rect 31089 3813 31098 3833
rect 30754 3804 30850 3806
rect 30950 3803 31098 3813
rect 31157 3833 31194 3843
rect 31269 3842 31306 3843
rect 31250 3840 31306 3842
rect 31157 3813 31165 3833
rect 31185 3813 31194 3833
rect 31006 3802 31042 3803
rect 30317 3736 30567 3738
rect 30317 3733 30418 3736
rect 30317 3714 30382 3733
rect 30379 3706 30382 3714
rect 30411 3706 30418 3733
rect 30446 3709 30456 3736
rect 30485 3714 30567 3736
rect 30485 3709 30489 3714
rect 30446 3706 30489 3709
rect 30379 3692 30489 3706
rect 29805 3674 30146 3675
rect 29730 3669 30146 3674
rect 30854 3671 30891 3672
rect 31157 3671 31194 3813
rect 31219 3833 31306 3840
rect 31219 3830 31277 3833
rect 31219 3810 31224 3830
rect 31245 3813 31277 3830
rect 31297 3813 31306 3833
rect 31245 3810 31306 3813
rect 31219 3803 31306 3810
rect 31365 3833 31402 3843
rect 31365 3813 31373 3833
rect 31393 3813 31402 3833
rect 31219 3802 31250 3803
rect 31365 3734 31402 3813
rect 31432 3842 31463 3895
rect 31667 3893 31735 3896
rect 31667 3851 31679 3893
rect 31728 3851 31735 3893
rect 31482 3842 31519 3843
rect 31432 3833 31519 3842
rect 31432 3813 31490 3833
rect 31510 3813 31519 3833
rect 31432 3803 31519 3813
rect 31578 3833 31615 3843
rect 31667 3838 31735 3851
rect 31890 3915 31955 3932
rect 31890 3897 31914 3915
rect 31932 3897 31955 3915
rect 32933 3925 32955 3943
rect 32973 3925 32998 3943
rect 32933 3904 32998 3925
rect 33146 3923 33211 3932
rect 31578 3813 31586 3833
rect 31606 3813 31615 3833
rect 31432 3802 31463 3803
rect 31427 3734 31537 3747
rect 31578 3734 31615 3813
rect 31890 3758 31955 3897
rect 33146 3886 33156 3923
rect 33196 3915 33211 3923
rect 33424 3916 33455 3969
rect 33485 3998 33522 4077
rect 33637 4008 33668 4009
rect 33485 3978 33494 3998
rect 33514 3978 33522 3998
rect 33485 3968 33522 3978
rect 33581 4001 33668 4008
rect 33581 3998 33642 4001
rect 33581 3978 33590 3998
rect 33610 3981 33642 3998
rect 33663 3981 33668 4001
rect 33610 3978 33668 3981
rect 33581 3971 33668 3978
rect 33693 3998 33730 4140
rect 33996 4139 34033 4140
rect 33845 4008 33881 4009
rect 33693 3978 33702 3998
rect 33722 3978 33730 3998
rect 33581 3969 33637 3971
rect 33581 3968 33618 3969
rect 33693 3968 33730 3978
rect 33789 3998 33937 4008
rect 34037 4005 34133 4007
rect 33789 3978 33798 3998
rect 33818 3978 33908 3998
rect 33928 3978 33937 3998
rect 33789 3972 33937 3978
rect 33789 3969 33853 3972
rect 33789 3968 33826 3969
rect 33845 3942 33853 3969
rect 33874 3969 33937 3972
rect 33995 3998 34133 4005
rect 35313 4000 35375 4512
rect 33995 3978 34004 3998
rect 34024 3978 34133 3998
rect 33995 3969 34133 3978
rect 33874 3942 33881 3969
rect 33900 3968 33937 3969
rect 33996 3968 34033 3969
rect 33845 3917 33881 3942
rect 33316 3915 33357 3916
rect 33196 3908 33357 3915
rect 33196 3888 33326 3908
rect 33346 3888 33357 3908
rect 33196 3886 33357 3888
rect 33146 3880 33357 3886
rect 33424 3912 33783 3916
rect 33424 3907 33746 3912
rect 33424 3883 33537 3907
rect 33561 3888 33746 3907
rect 33770 3888 33783 3912
rect 33561 3883 33783 3888
rect 33424 3880 33783 3883
rect 33845 3880 33880 3917
rect 33948 3914 34048 3917
rect 33948 3910 34015 3914
rect 33948 3884 33960 3910
rect 33986 3888 34015 3910
rect 34041 3888 34048 3914
rect 33986 3884 34048 3888
rect 33948 3880 34048 3884
rect 33146 3867 33213 3880
rect 31890 3752 31912 3758
rect 31365 3732 31615 3734
rect 31365 3729 31466 3732
rect 31365 3710 31430 3729
rect 31427 3702 31430 3710
rect 31459 3702 31466 3729
rect 31494 3705 31504 3732
rect 31533 3710 31615 3732
rect 31644 3740 31912 3752
rect 31930 3740 31955 3758
rect 31644 3717 31955 3740
rect 32938 3844 32994 3864
rect 32938 3826 32957 3844
rect 32975 3826 32994 3844
rect 31644 3716 31699 3717
rect 31533 3705 31537 3710
rect 31494 3702 31537 3705
rect 31427 3688 31537 3702
rect 30853 3670 31194 3671
rect 29730 3649 29733 3669
rect 29753 3649 30146 3669
rect 30778 3669 31194 3670
rect 31644 3669 31687 3716
rect 32938 3713 32994 3826
rect 33146 3846 33160 3867
rect 33196 3846 33213 3867
rect 33424 3859 33455 3880
rect 33845 3859 33881 3880
rect 33267 3858 33304 3859
rect 33146 3839 33213 3846
rect 33266 3849 33304 3858
rect 30778 3665 31687 3669
rect 30097 3616 30142 3649
rect 30778 3645 30781 3665
rect 30801 3645 31687 3665
rect 31155 3640 31687 3645
rect 31895 3659 31954 3681
rect 31895 3641 31914 3659
rect 31932 3641 31954 3659
rect 30943 3616 31042 3618
rect 30097 3606 31042 3616
rect 30097 3580 30965 3606
rect 30098 3579 30965 3580
rect 30943 3568 30965 3579
rect 30990 3571 31009 3606
rect 31034 3571 31042 3606
rect 30990 3568 31042 3571
rect 31895 3570 31954 3641
rect 32938 3575 32993 3713
rect 33146 3687 33211 3839
rect 33266 3829 33275 3849
rect 33295 3829 33304 3849
rect 33266 3821 33304 3829
rect 33370 3853 33455 3859
rect 33480 3858 33517 3859
rect 33370 3833 33378 3853
rect 33398 3833 33455 3853
rect 33370 3825 33455 3833
rect 33479 3849 33517 3858
rect 33479 3829 33488 3849
rect 33508 3829 33517 3849
rect 33370 3824 33406 3825
rect 33479 3821 33517 3829
rect 33583 3853 33668 3859
rect 33688 3858 33725 3859
rect 33583 3833 33591 3853
rect 33611 3852 33668 3853
rect 33611 3833 33640 3852
rect 33583 3832 33640 3833
rect 33661 3832 33668 3852
rect 33583 3825 33668 3832
rect 33687 3849 33725 3858
rect 33687 3829 33696 3849
rect 33716 3829 33725 3849
rect 33583 3824 33619 3825
rect 33687 3821 33725 3829
rect 33791 3853 33935 3859
rect 33791 3833 33799 3853
rect 33819 3833 33907 3853
rect 33927 3833 33935 3853
rect 33791 3825 33935 3833
rect 33791 3824 33827 3825
rect 33899 3824 33935 3825
rect 34001 3858 34038 3859
rect 34001 3857 34039 3858
rect 34001 3849 34065 3857
rect 34001 3829 34010 3849
rect 34030 3835 34065 3849
rect 34085 3835 34088 3855
rect 34030 3830 34088 3835
rect 34030 3829 34065 3830
rect 33267 3792 33304 3821
rect 33268 3790 33304 3792
rect 33480 3790 33517 3821
rect 33268 3768 33517 3790
rect 33349 3762 33460 3768
rect 33349 3754 33390 3762
rect 33349 3734 33357 3754
rect 33376 3734 33390 3754
rect 33349 3732 33390 3734
rect 33418 3754 33460 3762
rect 33418 3734 33434 3754
rect 33453 3734 33460 3754
rect 33418 3732 33460 3734
rect 33349 3719 33460 3732
rect 33688 3722 33725 3821
rect 34001 3817 34065 3829
rect 33139 3677 33260 3687
rect 33139 3675 33208 3677
rect 33139 3634 33152 3675
rect 33189 3636 33208 3675
rect 33245 3636 33260 3677
rect 33189 3634 33260 3636
rect 33139 3616 33260 3634
rect 32931 3572 32995 3575
rect 33351 3572 33455 3578
rect 33686 3572 33727 3722
rect 34105 3714 34132 3969
rect 34194 3959 34274 3970
rect 34194 3933 34211 3959
rect 34251 3933 34274 3959
rect 34194 3906 34274 3933
rect 35317 3961 35375 4000
rect 35317 3926 35379 3961
rect 34194 3880 34215 3906
rect 34255 3880 34274 3906
rect 34194 3861 34274 3880
rect 34194 3835 34218 3861
rect 34258 3835 34274 3861
rect 34194 3784 34274 3835
rect 35266 3899 35379 3926
rect 35266 3897 35325 3899
rect 35266 3866 35280 3897
rect 35305 3876 35325 3897
rect 35351 3876 35379 3899
rect 35305 3866 35379 3876
rect 35266 3856 35379 3866
rect 30943 3560 31042 3568
rect 30969 3559 31041 3560
rect 30623 3533 30690 3552
rect 30623 3512 30640 3533
rect 29504 3334 29584 3376
rect 30621 3467 30640 3512
rect 30670 3512 30690 3533
rect 30670 3467 30691 3512
rect 31160 3509 31201 3511
rect 31432 3509 31536 3511
rect 31892 3509 31956 3570
rect 28565 3223 28601 3224
rect 28457 3215 28601 3223
rect 28457 3195 28465 3215
rect 28485 3195 28573 3215
rect 28593 3195 28601 3215
rect 28457 3189 28601 3195
rect 28667 3219 28705 3227
rect 28773 3223 28809 3224
rect 28667 3199 28676 3219
rect 28696 3199 28705 3219
rect 28667 3190 28705 3199
rect 28724 3216 28809 3223
rect 28724 3196 28731 3216
rect 28752 3215 28809 3216
rect 28752 3196 28781 3215
rect 28724 3195 28781 3196
rect 28801 3195 28809 3215
rect 28667 3189 28704 3190
rect 28724 3189 28809 3195
rect 28875 3219 28913 3227
rect 28986 3223 29022 3224
rect 28875 3199 28884 3219
rect 28904 3199 28913 3219
rect 28875 3190 28913 3199
rect 28937 3215 29022 3223
rect 28937 3195 28994 3215
rect 29014 3195 29022 3215
rect 28875 3189 28912 3190
rect 28937 3189 29022 3195
rect 29088 3219 29126 3227
rect 29088 3199 29097 3219
rect 29117 3199 29126 3219
rect 29088 3190 29126 3199
rect 29326 3207 29412 3243
rect 29088 3189 29125 3190
rect 28511 3168 28547 3189
rect 28937 3168 28968 3189
rect 29164 3168 29210 3172
rect 28344 3164 28444 3168
rect 28344 3160 28406 3164
rect 28344 3134 28351 3160
rect 28377 3138 28406 3160
rect 28432 3138 28444 3164
rect 28377 3134 28444 3138
rect 28344 3131 28444 3134
rect 28512 3131 28547 3168
rect 28609 3165 28968 3168
rect 28609 3160 28831 3165
rect 28609 3136 28622 3160
rect 28646 3141 28831 3160
rect 28855 3141 28968 3165
rect 28646 3136 28968 3141
rect 28609 3132 28968 3136
rect 29035 3160 29210 3168
rect 29035 3140 29046 3160
rect 29066 3140 29210 3160
rect 29326 3166 29343 3207
rect 29397 3166 29412 3207
rect 29326 3147 29412 3166
rect 29035 3133 29210 3140
rect 29035 3132 29076 3133
rect 28511 3106 28547 3131
rect 28359 3079 28396 3080
rect 28455 3079 28492 3080
rect 28511 3079 28518 3106
rect 28259 3070 28397 3079
rect 28259 3050 28368 3070
rect 28388 3050 28397 3070
rect 28259 3043 28397 3050
rect 28455 3076 28518 3079
rect 28539 3079 28547 3106
rect 28566 3079 28603 3080
rect 28539 3076 28603 3079
rect 28455 3070 28603 3076
rect 28455 3050 28464 3070
rect 28484 3050 28574 3070
rect 28594 3050 28603 3070
rect 28259 3041 28355 3043
rect 28455 3040 28603 3050
rect 28662 3070 28699 3080
rect 28774 3079 28811 3080
rect 28755 3077 28811 3079
rect 28662 3050 28670 3070
rect 28690 3050 28699 3070
rect 28511 3039 28547 3040
rect 28359 2908 28396 2909
rect 28662 2908 28699 3050
rect 28724 3070 28811 3077
rect 28724 3067 28782 3070
rect 28724 3047 28729 3067
rect 28750 3050 28782 3067
rect 28802 3050 28811 3070
rect 28750 3047 28811 3050
rect 28724 3040 28811 3047
rect 28870 3070 28907 3080
rect 28870 3050 28878 3070
rect 28898 3050 28907 3070
rect 28724 3039 28755 3040
rect 28870 2971 28907 3050
rect 28937 3079 28968 3132
rect 28987 3079 29024 3080
rect 28937 3070 29024 3079
rect 28937 3050 28995 3070
rect 29015 3050 29024 3070
rect 28937 3040 29024 3050
rect 29083 3070 29120 3080
rect 29083 3050 29091 3070
rect 29111 3050 29120 3070
rect 28937 3039 28968 3040
rect 28932 2971 29042 2984
rect 29083 2971 29120 3050
rect 29164 3050 29210 3133
rect 29504 3050 29579 3334
rect 30621 3259 30691 3467
rect 30753 3474 31956 3509
rect 30753 3460 30781 3474
rect 30755 3329 30781 3460
rect 31160 3471 31956 3474
rect 32931 3569 33727 3572
rect 34106 3583 34132 3714
rect 34106 3569 34134 3583
rect 32931 3534 34134 3569
rect 34196 3576 34266 3784
rect 32931 3473 32995 3534
rect 33351 3532 33455 3534
rect 33686 3532 33727 3534
rect 34196 3531 34217 3576
rect 34197 3510 34217 3531
rect 34247 3531 34266 3576
rect 34247 3510 34264 3531
rect 34197 3491 34264 3510
rect 33846 3483 33918 3484
rect 33845 3475 33944 3483
rect 30613 3208 30693 3259
rect 30613 3182 30629 3208
rect 30669 3182 30693 3208
rect 30613 3163 30693 3182
rect 30613 3137 30632 3163
rect 30672 3137 30693 3163
rect 30613 3110 30693 3137
rect 30613 3084 30636 3110
rect 30676 3084 30693 3110
rect 30613 3073 30693 3084
rect 30755 3074 30782 3329
rect 31160 3321 31201 3471
rect 31432 3465 31536 3471
rect 31892 3468 31956 3471
rect 31627 3409 31748 3427
rect 31627 3407 31698 3409
rect 31627 3366 31642 3407
rect 31679 3368 31698 3407
rect 31735 3368 31748 3409
rect 31679 3366 31748 3368
rect 31627 3356 31748 3366
rect 30822 3214 30886 3226
rect 31162 3222 31199 3321
rect 31427 3311 31538 3324
rect 31427 3309 31469 3311
rect 31427 3289 31434 3309
rect 31453 3289 31469 3309
rect 31427 3281 31469 3289
rect 31497 3309 31538 3311
rect 31497 3289 31511 3309
rect 31530 3289 31538 3309
rect 31497 3281 31538 3289
rect 31427 3275 31538 3281
rect 31370 3253 31619 3275
rect 31370 3222 31407 3253
rect 31583 3251 31619 3253
rect 31583 3222 31620 3251
rect 30822 3213 30857 3214
rect 30799 3208 30857 3213
rect 30799 3188 30802 3208
rect 30822 3194 30857 3208
rect 30877 3194 30886 3214
rect 30822 3186 30886 3194
rect 30848 3185 30886 3186
rect 30849 3184 30886 3185
rect 30952 3218 30988 3219
rect 31060 3218 31096 3219
rect 30952 3210 31096 3218
rect 30952 3190 30960 3210
rect 30980 3190 31068 3210
rect 31088 3190 31096 3210
rect 30952 3184 31096 3190
rect 31162 3214 31200 3222
rect 31268 3218 31304 3219
rect 31162 3194 31171 3214
rect 31191 3194 31200 3214
rect 31162 3185 31200 3194
rect 31219 3211 31304 3218
rect 31219 3191 31226 3211
rect 31247 3210 31304 3211
rect 31247 3191 31276 3210
rect 31219 3190 31276 3191
rect 31296 3190 31304 3210
rect 31162 3184 31199 3185
rect 31219 3184 31304 3190
rect 31370 3214 31408 3222
rect 31481 3218 31517 3219
rect 31370 3194 31379 3214
rect 31399 3194 31408 3214
rect 31370 3185 31408 3194
rect 31432 3210 31517 3218
rect 31432 3190 31489 3210
rect 31509 3190 31517 3210
rect 31370 3184 31407 3185
rect 31432 3184 31517 3190
rect 31583 3214 31621 3222
rect 31583 3194 31592 3214
rect 31612 3194 31621 3214
rect 31676 3204 31741 3356
rect 31894 3330 31949 3468
rect 32933 3402 32992 3473
rect 33845 3472 33897 3475
rect 33845 3437 33853 3472
rect 33878 3437 33897 3472
rect 33922 3464 33944 3475
rect 33922 3463 34789 3464
rect 33922 3437 34790 3463
rect 33845 3427 34790 3437
rect 33845 3425 33944 3427
rect 32933 3384 32955 3402
rect 32973 3384 32992 3402
rect 32933 3362 32992 3384
rect 33200 3398 33732 3403
rect 33200 3378 34086 3398
rect 34106 3378 34109 3398
rect 34745 3394 34790 3427
rect 33200 3374 34109 3378
rect 31583 3185 31621 3194
rect 31674 3197 31741 3204
rect 31583 3184 31620 3185
rect 31006 3163 31042 3184
rect 31432 3163 31463 3184
rect 31674 3176 31691 3197
rect 31727 3176 31741 3197
rect 31893 3217 31949 3330
rect 33200 3327 33243 3374
rect 33693 3373 34109 3374
rect 34741 3374 35134 3394
rect 35154 3374 35157 3394
rect 33693 3372 34034 3373
rect 33350 3341 33460 3355
rect 33350 3338 33393 3341
rect 33350 3333 33354 3338
rect 33188 3326 33243 3327
rect 31893 3199 31912 3217
rect 31930 3199 31949 3217
rect 31893 3179 31949 3199
rect 32932 3303 33243 3326
rect 32932 3285 32957 3303
rect 32975 3291 33243 3303
rect 33272 3311 33354 3333
rect 33383 3311 33393 3338
rect 33421 3314 33428 3341
rect 33457 3333 33460 3341
rect 33457 3314 33522 3333
rect 33421 3311 33522 3314
rect 33272 3309 33522 3311
rect 32975 3285 32997 3291
rect 31674 3163 31741 3176
rect 30839 3159 30939 3163
rect 30839 3155 30901 3159
rect 30839 3129 30846 3155
rect 30872 3133 30901 3155
rect 30927 3133 30939 3159
rect 30872 3129 30939 3133
rect 30839 3126 30939 3129
rect 31007 3126 31042 3163
rect 31104 3160 31463 3163
rect 31104 3155 31326 3160
rect 31104 3131 31117 3155
rect 31141 3136 31326 3155
rect 31350 3136 31463 3160
rect 31141 3131 31463 3136
rect 31104 3127 31463 3131
rect 31530 3157 31741 3163
rect 31530 3155 31691 3157
rect 31530 3135 31541 3155
rect 31561 3135 31691 3155
rect 31530 3128 31691 3135
rect 31530 3127 31571 3128
rect 31006 3101 31042 3126
rect 30854 3074 30891 3075
rect 30950 3074 30987 3075
rect 31006 3074 31013 3101
rect 29164 3015 29579 3050
rect 30754 3065 30892 3074
rect 30754 3045 30863 3065
rect 30883 3045 30892 3065
rect 30754 3038 30892 3045
rect 30950 3071 31013 3074
rect 31034 3074 31042 3101
rect 31061 3074 31098 3075
rect 31034 3071 31098 3074
rect 30950 3065 31098 3071
rect 30950 3045 30959 3065
rect 30979 3045 31069 3065
rect 31089 3045 31098 3065
rect 30754 3036 30850 3038
rect 30950 3035 31098 3045
rect 31157 3065 31194 3075
rect 31269 3074 31306 3075
rect 31250 3072 31306 3074
rect 31157 3045 31165 3065
rect 31185 3045 31194 3065
rect 31006 3034 31042 3035
rect 29164 3014 29210 3015
rect 28870 2969 29120 2971
rect 28870 2966 28971 2969
rect 28870 2947 28935 2966
rect 28932 2939 28935 2947
rect 28964 2939 28971 2966
rect 28999 2942 29009 2969
rect 29038 2947 29120 2969
rect 29504 2963 29579 3015
rect 29038 2942 29042 2947
rect 28999 2939 29042 2942
rect 28932 2925 29042 2939
rect 28358 2907 28699 2908
rect 28283 2902 28699 2907
rect 28283 2882 28286 2902
rect 28306 2882 28700 2902
rect 24763 2473 27831 2498
rect 24763 2408 27626 2473
rect 27757 2408 27831 2473
rect 24763 2391 27831 2408
rect 28657 2378 28700 2882
rect 29317 2793 29412 2813
rect 29317 2749 29337 2793
rect 29397 2749 29412 2793
rect 29317 2453 29412 2749
rect 29317 2412 29350 2453
rect 29386 2412 29412 2453
rect 29512 2492 29574 2963
rect 30854 2903 30891 2904
rect 31157 2903 31194 3045
rect 31219 3065 31306 3072
rect 31219 3062 31277 3065
rect 31219 3042 31224 3062
rect 31245 3045 31277 3062
rect 31297 3045 31306 3065
rect 31245 3042 31306 3045
rect 31219 3035 31306 3042
rect 31365 3065 31402 3075
rect 31365 3045 31373 3065
rect 31393 3045 31402 3065
rect 31219 3034 31250 3035
rect 31365 2966 31402 3045
rect 31432 3074 31463 3127
rect 31676 3120 31691 3128
rect 31731 3120 31741 3157
rect 32932 3146 32997 3285
rect 33272 3230 33309 3309
rect 33350 3296 33460 3309
rect 33424 3240 33455 3241
rect 33272 3210 33281 3230
rect 33301 3210 33309 3230
rect 31676 3111 31741 3120
rect 31889 3118 31954 3139
rect 31889 3100 31914 3118
rect 31932 3100 31954 3118
rect 32932 3128 32955 3146
rect 32973 3128 32997 3146
rect 32932 3111 32997 3128
rect 33152 3192 33220 3205
rect 33272 3200 33309 3210
rect 33368 3230 33455 3240
rect 33368 3210 33377 3230
rect 33397 3210 33455 3230
rect 33368 3201 33455 3210
rect 33368 3200 33405 3201
rect 33152 3150 33159 3192
rect 33208 3150 33220 3192
rect 33152 3147 33220 3150
rect 33424 3148 33455 3201
rect 33485 3230 33522 3309
rect 33637 3240 33668 3241
rect 33485 3210 33494 3230
rect 33514 3210 33522 3230
rect 33485 3200 33522 3210
rect 33581 3233 33668 3240
rect 33581 3230 33642 3233
rect 33581 3210 33590 3230
rect 33610 3213 33642 3230
rect 33663 3213 33668 3233
rect 33610 3210 33668 3213
rect 33581 3203 33668 3210
rect 33693 3230 33730 3372
rect 33996 3371 34033 3372
rect 34741 3369 35157 3374
rect 34741 3368 35082 3369
rect 34398 3337 34508 3351
rect 34398 3334 34441 3337
rect 34398 3329 34402 3334
rect 34320 3307 34402 3329
rect 34431 3307 34441 3334
rect 34469 3310 34476 3337
rect 34505 3329 34508 3337
rect 34505 3310 34570 3329
rect 34469 3307 34570 3310
rect 34320 3305 34570 3307
rect 33845 3240 33881 3241
rect 33693 3210 33702 3230
rect 33722 3210 33730 3230
rect 33581 3201 33637 3203
rect 33581 3200 33618 3201
rect 33693 3200 33730 3210
rect 33789 3230 33937 3240
rect 34037 3237 34133 3239
rect 33789 3210 33798 3230
rect 33818 3210 33908 3230
rect 33928 3210 33937 3230
rect 33789 3204 33937 3210
rect 33789 3201 33853 3204
rect 33789 3200 33826 3201
rect 33845 3174 33853 3201
rect 33874 3201 33937 3204
rect 33995 3230 34133 3237
rect 33995 3210 34004 3230
rect 34024 3210 34133 3230
rect 33995 3201 34133 3210
rect 34320 3226 34357 3305
rect 34398 3292 34508 3305
rect 34472 3236 34503 3237
rect 34320 3206 34329 3226
rect 34349 3206 34357 3226
rect 33874 3174 33881 3201
rect 33900 3200 33937 3201
rect 33996 3200 34033 3201
rect 33845 3149 33881 3174
rect 33316 3147 33357 3148
rect 33152 3140 33357 3147
rect 33152 3129 33326 3140
rect 31482 3074 31519 3075
rect 31432 3065 31519 3074
rect 31432 3045 31490 3065
rect 31510 3045 31519 3065
rect 31432 3035 31519 3045
rect 31578 3065 31615 3075
rect 31578 3045 31586 3065
rect 31606 3045 31615 3065
rect 31432 3034 31463 3035
rect 31427 2966 31537 2979
rect 31578 2966 31615 3045
rect 31889 3024 31954 3100
rect 33152 3096 33160 3129
rect 33153 3087 33160 3096
rect 33209 3120 33326 3129
rect 33346 3120 33357 3140
rect 33209 3112 33357 3120
rect 33424 3144 33783 3148
rect 33424 3139 33746 3144
rect 33424 3115 33537 3139
rect 33561 3120 33746 3139
rect 33770 3120 33783 3144
rect 33561 3115 33783 3120
rect 33424 3112 33783 3115
rect 33845 3112 33880 3149
rect 33948 3146 34048 3149
rect 33948 3142 34015 3146
rect 33948 3116 33960 3142
rect 33986 3120 34015 3142
rect 34041 3120 34048 3146
rect 33986 3116 34048 3120
rect 33948 3112 34048 3116
rect 33209 3096 33220 3112
rect 33209 3087 33217 3096
rect 33424 3091 33455 3112
rect 33845 3091 33881 3112
rect 33267 3090 33304 3091
rect 32932 3047 32997 3066
rect 32932 3029 32957 3047
rect 32975 3029 32997 3047
rect 31365 2964 31615 2966
rect 31365 2961 31466 2964
rect 31365 2942 31430 2961
rect 31427 2934 31430 2942
rect 31459 2934 31466 2961
rect 31494 2937 31504 2964
rect 31533 2942 31615 2964
rect 31638 2989 31955 3024
rect 31533 2937 31537 2942
rect 31494 2934 31537 2937
rect 31427 2920 31537 2934
rect 30853 2902 31194 2903
rect 30778 2900 31194 2902
rect 31638 2900 31678 2989
rect 31889 2962 31954 2989
rect 31889 2944 31912 2962
rect 31930 2944 31954 2962
rect 31889 2924 31954 2944
rect 30775 2897 31678 2900
rect 30775 2877 30781 2897
rect 30801 2877 31678 2897
rect 30775 2873 31678 2877
rect 31638 2870 31678 2873
rect 31890 2863 31955 2884
rect 30108 2855 30769 2856
rect 30108 2848 31042 2855
rect 30108 2847 31014 2848
rect 30108 2827 30959 2847
rect 30991 2828 31014 2847
rect 31039 2828 31042 2848
rect 30991 2827 31042 2828
rect 30108 2820 31042 2827
rect 29707 2778 29875 2779
rect 30110 2778 30149 2820
rect 30938 2818 31042 2820
rect 31007 2816 31042 2818
rect 31890 2845 31914 2863
rect 31932 2845 31955 2863
rect 31890 2798 31955 2845
rect 29707 2752 30151 2778
rect 29707 2750 29875 2752
rect 29512 2473 29576 2492
rect 29512 2434 29529 2473
rect 29563 2434 29576 2473
rect 29512 2415 29576 2434
rect 29317 2386 29412 2412
rect 29707 2399 29734 2750
rect 30110 2746 30151 2752
rect 29774 2539 29838 2551
rect 30114 2547 30151 2746
rect 30613 2773 30685 2790
rect 30613 2734 30621 2773
rect 30666 2734 30685 2773
rect 30379 2636 30490 2651
rect 30379 2634 30421 2636
rect 30379 2614 30386 2634
rect 30405 2614 30421 2634
rect 30379 2606 30421 2614
rect 30449 2634 30490 2636
rect 30449 2614 30463 2634
rect 30482 2614 30490 2634
rect 30449 2606 30490 2614
rect 30379 2600 30490 2606
rect 30322 2578 30571 2600
rect 30322 2547 30359 2578
rect 30535 2576 30571 2578
rect 30535 2547 30572 2576
rect 29774 2538 29809 2539
rect 29751 2533 29809 2538
rect 29751 2513 29754 2533
rect 29774 2519 29809 2533
rect 29829 2519 29838 2539
rect 29774 2511 29838 2519
rect 29800 2510 29838 2511
rect 29801 2509 29838 2510
rect 29904 2543 29940 2544
rect 30012 2543 30048 2544
rect 29904 2535 30048 2543
rect 29904 2515 29912 2535
rect 29932 2515 30020 2535
rect 30040 2515 30048 2535
rect 29904 2509 30048 2515
rect 30114 2539 30152 2547
rect 30220 2543 30256 2544
rect 30114 2519 30123 2539
rect 30143 2519 30152 2539
rect 30114 2510 30152 2519
rect 30171 2536 30256 2543
rect 30171 2516 30178 2536
rect 30199 2535 30256 2536
rect 30199 2516 30228 2535
rect 30171 2515 30228 2516
rect 30248 2515 30256 2535
rect 30114 2509 30151 2510
rect 30171 2509 30256 2515
rect 30322 2539 30360 2547
rect 30433 2543 30469 2544
rect 30322 2519 30331 2539
rect 30351 2519 30360 2539
rect 30322 2510 30360 2519
rect 30384 2535 30469 2543
rect 30384 2515 30441 2535
rect 30461 2515 30469 2535
rect 30322 2509 30359 2510
rect 30384 2509 30469 2515
rect 30535 2539 30573 2547
rect 30535 2519 30544 2539
rect 30564 2519 30573 2539
rect 30535 2510 30573 2519
rect 30613 2524 30685 2734
rect 30755 2768 31955 2798
rect 30755 2767 31199 2768
rect 30755 2765 30923 2767
rect 30613 2510 30696 2524
rect 30535 2509 30572 2510
rect 29958 2488 29994 2509
rect 30384 2488 30415 2509
rect 30613 2488 30630 2510
rect 29791 2484 29891 2488
rect 29791 2480 29853 2484
rect 29791 2454 29798 2480
rect 29824 2458 29853 2480
rect 29879 2458 29891 2484
rect 29824 2454 29891 2458
rect 29791 2451 29891 2454
rect 29959 2451 29994 2488
rect 30056 2485 30415 2488
rect 30056 2480 30278 2485
rect 30056 2456 30069 2480
rect 30093 2461 30278 2480
rect 30302 2461 30415 2485
rect 30093 2456 30415 2461
rect 30056 2452 30415 2456
rect 30482 2480 30630 2488
rect 30482 2460 30493 2480
rect 30513 2477 30630 2480
rect 30683 2477 30696 2510
rect 30513 2460 30696 2477
rect 30482 2453 30696 2460
rect 30482 2452 30523 2453
rect 30613 2452 30696 2453
rect 29958 2426 29994 2451
rect 29806 2399 29843 2400
rect 29902 2399 29939 2400
rect 29958 2399 29965 2426
rect 29706 2390 29844 2399
rect 24518 2292 24675 2305
rect 24518 2288 24679 2292
rect 23398 2142 23424 2247
rect 24518 2181 24559 2288
rect 24659 2181 24679 2288
rect 24518 2152 24679 2181
rect 28655 2169 28704 2378
rect 29706 2370 29815 2390
rect 29835 2370 29844 2390
rect 29706 2363 29844 2370
rect 29902 2396 29965 2399
rect 29986 2399 29994 2426
rect 30013 2399 30050 2400
rect 29986 2396 30050 2399
rect 29902 2390 30050 2396
rect 29902 2370 29911 2390
rect 29931 2370 30021 2390
rect 30041 2370 30050 2390
rect 29706 2361 29802 2363
rect 29902 2360 30050 2370
rect 30109 2390 30146 2400
rect 30221 2399 30258 2400
rect 30202 2397 30258 2399
rect 30109 2370 30117 2390
rect 30137 2370 30146 2390
rect 29958 2359 29994 2360
rect 29806 2228 29843 2229
rect 30109 2228 30146 2370
rect 30171 2390 30258 2397
rect 30171 2387 30229 2390
rect 30171 2367 30176 2387
rect 30197 2370 30229 2387
rect 30249 2370 30258 2390
rect 30197 2367 30258 2370
rect 30171 2360 30258 2367
rect 30317 2390 30354 2400
rect 30317 2370 30325 2390
rect 30345 2370 30354 2390
rect 30171 2359 30202 2360
rect 30317 2291 30354 2370
rect 30384 2399 30415 2452
rect 30621 2419 30635 2452
rect 30688 2419 30696 2452
rect 30621 2413 30696 2419
rect 30621 2408 30691 2413
rect 30434 2399 30471 2400
rect 30384 2390 30471 2399
rect 30384 2370 30442 2390
rect 30462 2370 30471 2390
rect 30384 2360 30471 2370
rect 30530 2390 30567 2400
rect 30755 2395 30782 2765
rect 30822 2535 30886 2547
rect 31162 2543 31199 2767
rect 31670 2748 31734 2750
rect 31666 2736 31734 2748
rect 31666 2703 31677 2736
rect 31717 2703 31734 2736
rect 31666 2693 31734 2703
rect 31427 2632 31538 2647
rect 31427 2630 31469 2632
rect 31427 2610 31434 2630
rect 31453 2610 31469 2630
rect 31427 2602 31469 2610
rect 31497 2630 31538 2632
rect 31497 2610 31511 2630
rect 31530 2610 31538 2630
rect 31497 2602 31538 2610
rect 31427 2596 31538 2602
rect 31370 2574 31619 2596
rect 31370 2543 31407 2574
rect 31583 2572 31619 2574
rect 31583 2543 31620 2572
rect 30822 2534 30857 2535
rect 30799 2529 30857 2534
rect 30799 2509 30802 2529
rect 30822 2515 30857 2529
rect 30877 2515 30886 2535
rect 30822 2507 30886 2515
rect 30848 2506 30886 2507
rect 30849 2505 30886 2506
rect 30952 2539 30988 2540
rect 31060 2539 31096 2540
rect 30952 2531 31096 2539
rect 30952 2511 30960 2531
rect 30980 2511 31068 2531
rect 31088 2511 31096 2531
rect 30952 2505 31096 2511
rect 31162 2535 31200 2543
rect 31268 2539 31304 2540
rect 31162 2515 31171 2535
rect 31191 2515 31200 2535
rect 31162 2506 31200 2515
rect 31219 2532 31304 2539
rect 31219 2512 31226 2532
rect 31247 2531 31304 2532
rect 31247 2512 31276 2531
rect 31219 2511 31276 2512
rect 31296 2511 31304 2531
rect 31162 2505 31199 2506
rect 31219 2505 31304 2511
rect 31370 2535 31408 2543
rect 31481 2539 31517 2540
rect 31370 2515 31379 2535
rect 31399 2515 31408 2535
rect 31370 2506 31408 2515
rect 31432 2531 31517 2539
rect 31432 2511 31489 2531
rect 31509 2511 31517 2531
rect 31370 2505 31407 2506
rect 31432 2505 31517 2511
rect 31583 2535 31621 2543
rect 31583 2515 31592 2535
rect 31612 2515 31621 2535
rect 31583 2506 31621 2515
rect 31670 2509 31734 2693
rect 31890 2567 31955 2768
rect 32932 2828 32997 3029
rect 33153 2903 33217 3087
rect 33266 3081 33304 3090
rect 33266 3061 33275 3081
rect 33295 3061 33304 3081
rect 33266 3053 33304 3061
rect 33370 3085 33455 3091
rect 33480 3090 33517 3091
rect 33370 3065 33378 3085
rect 33398 3065 33455 3085
rect 33370 3057 33455 3065
rect 33479 3081 33517 3090
rect 33479 3061 33488 3081
rect 33508 3061 33517 3081
rect 33370 3056 33406 3057
rect 33479 3053 33517 3061
rect 33583 3085 33668 3091
rect 33688 3090 33725 3091
rect 33583 3065 33591 3085
rect 33611 3084 33668 3085
rect 33611 3065 33640 3084
rect 33583 3064 33640 3065
rect 33661 3064 33668 3084
rect 33583 3057 33668 3064
rect 33687 3081 33725 3090
rect 33687 3061 33696 3081
rect 33716 3061 33725 3081
rect 33583 3056 33619 3057
rect 33687 3053 33725 3061
rect 33791 3085 33935 3091
rect 33791 3065 33799 3085
rect 33819 3065 33907 3085
rect 33927 3065 33935 3085
rect 33791 3057 33935 3065
rect 33791 3056 33827 3057
rect 33899 3056 33935 3057
rect 34001 3090 34038 3091
rect 34001 3089 34039 3090
rect 34001 3081 34065 3089
rect 34001 3061 34010 3081
rect 34030 3067 34065 3081
rect 34085 3067 34088 3087
rect 34030 3062 34088 3067
rect 34030 3061 34065 3062
rect 33267 3024 33304 3053
rect 33268 3022 33304 3024
rect 33480 3022 33517 3053
rect 33268 3000 33517 3022
rect 33349 2994 33460 3000
rect 33349 2986 33390 2994
rect 33349 2966 33357 2986
rect 33376 2966 33390 2986
rect 33349 2964 33390 2966
rect 33418 2986 33460 2994
rect 33418 2966 33434 2986
rect 33453 2966 33460 2986
rect 33418 2964 33460 2966
rect 33349 2949 33460 2964
rect 33153 2893 33221 2903
rect 33153 2860 33170 2893
rect 33210 2860 33221 2893
rect 33153 2848 33221 2860
rect 33153 2846 33217 2848
rect 33688 2829 33725 3053
rect 34001 3049 34065 3061
rect 34105 2831 34132 3201
rect 34320 3196 34357 3206
rect 34416 3226 34503 3236
rect 34416 3206 34425 3226
rect 34445 3206 34503 3226
rect 34416 3197 34503 3206
rect 34416 3196 34453 3197
rect 34196 3183 34266 3188
rect 34191 3177 34266 3183
rect 34191 3144 34199 3177
rect 34252 3144 34266 3177
rect 34472 3144 34503 3197
rect 34533 3226 34570 3305
rect 34685 3236 34716 3237
rect 34533 3206 34542 3226
rect 34562 3206 34570 3226
rect 34533 3196 34570 3206
rect 34629 3229 34716 3236
rect 34629 3226 34690 3229
rect 34629 3206 34638 3226
rect 34658 3209 34690 3226
rect 34711 3209 34716 3229
rect 34658 3206 34716 3209
rect 34629 3199 34716 3206
rect 34741 3226 34778 3368
rect 35044 3367 35081 3368
rect 34893 3236 34929 3237
rect 34741 3206 34750 3226
rect 34770 3206 34778 3226
rect 34629 3197 34685 3199
rect 34629 3196 34666 3197
rect 34741 3196 34778 3206
rect 34837 3226 34985 3236
rect 35085 3233 35181 3235
rect 34837 3206 34846 3226
rect 34866 3206 34956 3226
rect 34976 3206 34985 3226
rect 34837 3200 34985 3206
rect 34837 3197 34901 3200
rect 34837 3196 34874 3197
rect 34893 3170 34901 3197
rect 34922 3197 34985 3200
rect 35043 3226 35181 3233
rect 35043 3206 35052 3226
rect 35072 3206 35181 3226
rect 35043 3197 35181 3206
rect 34922 3170 34929 3197
rect 34948 3196 34985 3197
rect 35044 3196 35081 3197
rect 34893 3145 34929 3170
rect 34191 3143 34274 3144
rect 34364 3143 34405 3144
rect 34191 3136 34405 3143
rect 34191 3119 34374 3136
rect 34191 3086 34204 3119
rect 34257 3116 34374 3119
rect 34394 3116 34405 3136
rect 34257 3108 34405 3116
rect 34472 3140 34831 3144
rect 34472 3135 34794 3140
rect 34472 3111 34585 3135
rect 34609 3116 34794 3135
rect 34818 3116 34831 3140
rect 34609 3111 34831 3116
rect 34472 3108 34831 3111
rect 34893 3108 34928 3145
rect 34996 3142 35096 3145
rect 34996 3138 35063 3142
rect 34996 3112 35008 3138
rect 35034 3116 35063 3138
rect 35089 3116 35096 3142
rect 35034 3112 35096 3116
rect 34996 3108 35096 3112
rect 34257 3086 34274 3108
rect 34472 3087 34503 3108
rect 34893 3087 34929 3108
rect 34315 3086 34352 3087
rect 34191 3072 34274 3086
rect 33964 2829 34132 2831
rect 33688 2828 34132 2829
rect 32932 2798 34132 2828
rect 34202 2862 34274 3072
rect 34314 3077 34352 3086
rect 34314 3057 34323 3077
rect 34343 3057 34352 3077
rect 34314 3049 34352 3057
rect 34418 3081 34503 3087
rect 34528 3086 34565 3087
rect 34418 3061 34426 3081
rect 34446 3061 34503 3081
rect 34418 3053 34503 3061
rect 34527 3077 34565 3086
rect 34527 3057 34536 3077
rect 34556 3057 34565 3077
rect 34418 3052 34454 3053
rect 34527 3049 34565 3057
rect 34631 3081 34716 3087
rect 34736 3086 34773 3087
rect 34631 3061 34639 3081
rect 34659 3080 34716 3081
rect 34659 3061 34688 3080
rect 34631 3060 34688 3061
rect 34709 3060 34716 3080
rect 34631 3053 34716 3060
rect 34735 3077 34773 3086
rect 34735 3057 34744 3077
rect 34764 3057 34773 3077
rect 34631 3052 34667 3053
rect 34735 3049 34773 3057
rect 34839 3081 34983 3087
rect 34839 3061 34847 3081
rect 34867 3061 34955 3081
rect 34975 3061 34983 3081
rect 34839 3053 34983 3061
rect 34839 3052 34875 3053
rect 34947 3052 34983 3053
rect 35049 3086 35086 3087
rect 35049 3085 35087 3086
rect 35049 3077 35113 3085
rect 35049 3057 35058 3077
rect 35078 3063 35113 3077
rect 35133 3063 35136 3083
rect 35078 3058 35136 3063
rect 35078 3057 35113 3058
rect 34315 3020 34352 3049
rect 34316 3018 34352 3020
rect 34528 3018 34565 3049
rect 34316 2996 34565 3018
rect 34397 2990 34508 2996
rect 34397 2982 34438 2990
rect 34397 2962 34405 2982
rect 34424 2962 34438 2982
rect 34397 2960 34438 2962
rect 34466 2982 34508 2990
rect 34466 2962 34482 2982
rect 34501 2962 34508 2982
rect 34466 2960 34508 2962
rect 34397 2945 34508 2960
rect 34202 2823 34221 2862
rect 34266 2823 34274 2862
rect 34202 2806 34274 2823
rect 34736 2850 34773 3049
rect 35049 3045 35113 3057
rect 34736 2844 34777 2850
rect 35153 2846 35180 3197
rect 35012 2844 35180 2846
rect 34736 2818 35180 2844
rect 32932 2751 32997 2798
rect 32932 2733 32955 2751
rect 32973 2733 32997 2751
rect 33845 2778 33880 2780
rect 33845 2776 33949 2778
rect 34738 2776 34777 2818
rect 35012 2817 35180 2818
rect 33845 2769 34779 2776
rect 33845 2768 33896 2769
rect 33845 2748 33848 2768
rect 33873 2749 33896 2768
rect 33928 2749 34779 2769
rect 33873 2748 34779 2749
rect 33845 2741 34779 2748
rect 34118 2740 34779 2741
rect 32932 2712 32997 2733
rect 33209 2723 33249 2726
rect 33209 2719 34112 2723
rect 33209 2699 34086 2719
rect 34106 2699 34112 2719
rect 33209 2696 34112 2699
rect 32933 2652 32998 2672
rect 32933 2634 32957 2652
rect 32975 2634 32998 2652
rect 32933 2607 32998 2634
rect 33209 2607 33249 2696
rect 33693 2694 34109 2696
rect 33693 2693 34034 2694
rect 33350 2662 33460 2676
rect 33350 2659 33393 2662
rect 33350 2654 33354 2659
rect 32932 2572 33249 2607
rect 33272 2632 33354 2654
rect 33383 2632 33393 2659
rect 33421 2635 33428 2662
rect 33457 2654 33460 2662
rect 33457 2635 33522 2654
rect 33421 2632 33522 2635
rect 33272 2630 33522 2632
rect 31890 2549 31912 2567
rect 31930 2549 31955 2567
rect 31890 2530 31955 2549
rect 31583 2505 31620 2506
rect 31006 2484 31042 2505
rect 31432 2484 31463 2505
rect 31670 2500 31678 2509
rect 31667 2484 31678 2500
rect 30839 2480 30939 2484
rect 30839 2476 30901 2480
rect 30839 2450 30846 2476
rect 30872 2454 30901 2476
rect 30927 2454 30939 2480
rect 30872 2450 30939 2454
rect 30839 2447 30939 2450
rect 31007 2447 31042 2484
rect 31104 2481 31463 2484
rect 31104 2476 31326 2481
rect 31104 2452 31117 2476
rect 31141 2457 31326 2476
rect 31350 2457 31463 2481
rect 31141 2452 31463 2457
rect 31104 2448 31463 2452
rect 31530 2476 31678 2484
rect 31530 2456 31541 2476
rect 31561 2467 31678 2476
rect 31727 2500 31734 2509
rect 31727 2467 31735 2500
rect 32933 2496 32998 2572
rect 33272 2551 33309 2630
rect 33350 2617 33460 2630
rect 33424 2561 33455 2562
rect 33272 2531 33281 2551
rect 33301 2531 33309 2551
rect 33272 2521 33309 2531
rect 33368 2551 33455 2561
rect 33368 2531 33377 2551
rect 33397 2531 33455 2551
rect 33368 2522 33455 2531
rect 33368 2521 33405 2522
rect 31561 2456 31735 2467
rect 31530 2449 31735 2456
rect 31530 2448 31571 2449
rect 31006 2422 31042 2447
rect 30854 2395 30891 2396
rect 30950 2395 30987 2396
rect 31006 2395 31013 2422
rect 30530 2370 30538 2390
rect 30558 2370 30567 2390
rect 30384 2359 30415 2360
rect 30379 2291 30489 2304
rect 30530 2291 30567 2370
rect 30754 2386 30892 2395
rect 30754 2366 30863 2386
rect 30883 2366 30892 2386
rect 30754 2359 30892 2366
rect 30950 2392 31013 2395
rect 31034 2395 31042 2422
rect 31061 2395 31098 2396
rect 31034 2392 31098 2395
rect 30950 2386 31098 2392
rect 30950 2366 30959 2386
rect 30979 2366 31069 2386
rect 31089 2366 31098 2386
rect 30754 2357 30850 2359
rect 30950 2356 31098 2366
rect 31157 2386 31194 2396
rect 31269 2395 31306 2396
rect 31250 2393 31306 2395
rect 31157 2366 31165 2386
rect 31185 2366 31194 2386
rect 31006 2355 31042 2356
rect 30317 2289 30567 2291
rect 30317 2286 30418 2289
rect 30317 2267 30382 2286
rect 30379 2259 30382 2267
rect 30411 2259 30418 2286
rect 30446 2262 30456 2289
rect 30485 2267 30567 2289
rect 30485 2262 30489 2267
rect 30446 2259 30489 2262
rect 30379 2245 30489 2259
rect 29805 2227 30146 2228
rect 29730 2222 30146 2227
rect 30854 2224 30891 2225
rect 31157 2224 31194 2366
rect 31219 2386 31306 2393
rect 31219 2383 31277 2386
rect 31219 2363 31224 2383
rect 31245 2366 31277 2383
rect 31297 2366 31306 2386
rect 31245 2363 31306 2366
rect 31219 2356 31306 2363
rect 31365 2386 31402 2396
rect 31365 2366 31373 2386
rect 31393 2366 31402 2386
rect 31219 2355 31250 2356
rect 31365 2287 31402 2366
rect 31432 2395 31463 2448
rect 31667 2446 31735 2449
rect 31667 2404 31679 2446
rect 31728 2404 31735 2446
rect 31482 2395 31519 2396
rect 31432 2386 31519 2395
rect 31432 2366 31490 2386
rect 31510 2366 31519 2386
rect 31432 2356 31519 2366
rect 31578 2386 31615 2396
rect 31667 2391 31735 2404
rect 31890 2468 31955 2485
rect 31890 2450 31914 2468
rect 31932 2450 31955 2468
rect 32933 2478 32955 2496
rect 32973 2478 32998 2496
rect 32933 2457 32998 2478
rect 33146 2476 33211 2485
rect 31578 2366 31586 2386
rect 31606 2366 31615 2386
rect 31432 2355 31463 2356
rect 31427 2287 31537 2300
rect 31578 2287 31615 2366
rect 31890 2311 31955 2450
rect 33146 2439 33156 2476
rect 33196 2468 33211 2476
rect 33424 2469 33455 2522
rect 33485 2551 33522 2630
rect 33637 2561 33668 2562
rect 33485 2531 33494 2551
rect 33514 2531 33522 2551
rect 33485 2521 33522 2531
rect 33581 2554 33668 2561
rect 33581 2551 33642 2554
rect 33581 2531 33590 2551
rect 33610 2534 33642 2551
rect 33663 2534 33668 2554
rect 33610 2531 33668 2534
rect 33581 2524 33668 2531
rect 33693 2551 33730 2693
rect 33996 2692 34033 2693
rect 33845 2561 33881 2562
rect 33693 2531 33702 2551
rect 33722 2531 33730 2551
rect 33581 2522 33637 2524
rect 33581 2521 33618 2522
rect 33693 2521 33730 2531
rect 33789 2551 33937 2561
rect 34037 2558 34133 2560
rect 33789 2531 33798 2551
rect 33818 2531 33908 2551
rect 33928 2531 33937 2551
rect 33789 2525 33937 2531
rect 33789 2522 33853 2525
rect 33789 2521 33826 2522
rect 33845 2495 33853 2522
rect 33874 2522 33937 2525
rect 33995 2551 34133 2558
rect 33995 2531 34004 2551
rect 34024 2531 34133 2551
rect 33995 2522 34133 2531
rect 33874 2495 33881 2522
rect 33900 2521 33937 2522
rect 33996 2521 34033 2522
rect 33845 2470 33881 2495
rect 33316 2468 33357 2469
rect 33196 2461 33357 2468
rect 33196 2441 33326 2461
rect 33346 2441 33357 2461
rect 33196 2439 33357 2441
rect 33146 2433 33357 2439
rect 33424 2465 33783 2469
rect 33424 2460 33746 2465
rect 33424 2436 33537 2460
rect 33561 2441 33746 2460
rect 33770 2441 33783 2465
rect 33561 2436 33783 2441
rect 33424 2433 33783 2436
rect 33845 2433 33880 2470
rect 33948 2467 34048 2470
rect 33948 2463 34015 2467
rect 33948 2437 33960 2463
rect 33986 2441 34015 2463
rect 34041 2441 34048 2467
rect 33986 2437 34048 2441
rect 33948 2433 34048 2437
rect 33146 2420 33213 2433
rect 32938 2397 32994 2417
rect 32938 2379 32957 2397
rect 32975 2379 32994 2397
rect 32938 2344 32994 2379
rect 31890 2305 31912 2311
rect 31365 2285 31615 2287
rect 31365 2282 31466 2285
rect 31365 2263 31430 2282
rect 31427 2255 31430 2263
rect 31459 2255 31466 2282
rect 31494 2258 31504 2285
rect 31533 2263 31615 2285
rect 31644 2293 31912 2305
rect 31930 2293 31955 2311
rect 31644 2270 31955 2293
rect 31644 2269 31699 2270
rect 31533 2258 31537 2263
rect 31494 2255 31537 2258
rect 31427 2241 31537 2255
rect 30853 2223 31194 2224
rect 29730 2202 29733 2222
rect 29753 2202 30146 2222
rect 30778 2222 31194 2223
rect 31644 2222 31687 2269
rect 32900 2266 32994 2344
rect 33146 2399 33160 2420
rect 33196 2399 33213 2420
rect 33424 2412 33455 2433
rect 33845 2412 33881 2433
rect 33267 2411 33304 2412
rect 33146 2392 33213 2399
rect 33266 2402 33304 2411
rect 30778 2218 31687 2222
rect 23398 2128 23426 2142
rect 24522 2139 24679 2152
rect 28653 2167 29470 2169
rect 29903 2167 29992 2170
rect 28653 2158 29992 2167
rect 22200 2093 23426 2128
rect 28653 2120 29915 2158
rect 29940 2123 29959 2158
rect 29984 2123 29992 2158
rect 30097 2169 30142 2202
rect 30778 2198 30781 2218
rect 30801 2198 31687 2218
rect 31155 2193 31687 2198
rect 31895 2212 31954 2234
rect 31895 2194 31914 2212
rect 31932 2194 31954 2212
rect 30943 2169 31042 2171
rect 30097 2159 31042 2169
rect 30097 2133 30965 2159
rect 30098 2132 30965 2133
rect 29940 2120 29992 2123
rect 28653 2112 29992 2120
rect 30943 2121 30965 2132
rect 30990 2124 31009 2159
rect 31034 2124 31042 2159
rect 30990 2121 31042 2124
rect 30943 2113 31042 2121
rect 30969 2112 31041 2113
rect 28653 2111 29991 2112
rect 28653 2109 29470 2111
rect 29244 2105 29470 2109
rect 22200 2017 22285 2093
rect 22643 2091 22747 2093
rect 22978 2091 23019 2093
rect 31895 2017 31954 2194
rect 32900 2125 32993 2266
rect 33146 2240 33211 2392
rect 33266 2382 33275 2402
rect 33295 2382 33304 2402
rect 33266 2374 33304 2382
rect 33370 2406 33455 2412
rect 33480 2411 33517 2412
rect 33370 2386 33378 2406
rect 33398 2386 33455 2406
rect 33370 2378 33455 2386
rect 33479 2402 33517 2411
rect 33479 2382 33488 2402
rect 33508 2382 33517 2402
rect 33370 2377 33406 2378
rect 33479 2374 33517 2382
rect 33583 2406 33668 2412
rect 33688 2411 33725 2412
rect 33583 2386 33591 2406
rect 33611 2405 33668 2406
rect 33611 2386 33640 2405
rect 33583 2385 33640 2386
rect 33661 2385 33668 2405
rect 33583 2378 33668 2385
rect 33687 2402 33725 2411
rect 33687 2382 33696 2402
rect 33716 2382 33725 2402
rect 33583 2377 33619 2378
rect 33687 2374 33725 2382
rect 33791 2406 33935 2412
rect 33791 2386 33799 2406
rect 33819 2386 33907 2406
rect 33927 2386 33935 2406
rect 33791 2378 33935 2386
rect 33791 2377 33827 2378
rect 33899 2377 33935 2378
rect 34001 2411 34038 2412
rect 34001 2410 34039 2411
rect 34001 2402 34065 2410
rect 34001 2382 34010 2402
rect 34030 2388 34065 2402
rect 34085 2388 34088 2408
rect 34030 2383 34088 2388
rect 34030 2382 34065 2383
rect 33267 2345 33304 2374
rect 33268 2343 33304 2345
rect 33480 2343 33517 2374
rect 33268 2321 33517 2343
rect 33349 2315 33460 2321
rect 33349 2307 33390 2315
rect 33349 2287 33357 2307
rect 33376 2287 33390 2307
rect 33349 2285 33390 2287
rect 33418 2307 33460 2315
rect 33418 2287 33434 2307
rect 33453 2287 33460 2307
rect 33418 2285 33460 2287
rect 33349 2270 33460 2285
rect 33688 2275 33725 2374
rect 34001 2370 34065 2382
rect 34105 2331 34132 2522
rect 33351 2261 33455 2270
rect 33139 2230 33260 2240
rect 33139 2228 33208 2230
rect 33139 2187 33152 2228
rect 33189 2189 33208 2228
rect 33245 2189 33260 2230
rect 33189 2187 33260 2189
rect 33139 2169 33260 2187
rect 33351 2125 33455 2134
rect 33686 2125 33727 2275
rect 32900 2123 33727 2125
rect 32908 2122 33727 2123
rect 34106 2241 34131 2331
rect 35266 2299 35365 3856
rect 35471 2492 35570 5393
rect 35961 5376 35992 5397
rect 36382 5376 36418 5397
rect 35804 5375 35841 5376
rect 35803 5366 35841 5375
rect 35803 5346 35812 5366
rect 35832 5346 35841 5366
rect 35803 5338 35841 5346
rect 35907 5370 35992 5376
rect 36017 5375 36054 5376
rect 35907 5350 35915 5370
rect 35935 5350 35992 5370
rect 35907 5342 35992 5350
rect 36016 5366 36054 5375
rect 36016 5346 36025 5366
rect 36045 5346 36054 5366
rect 35907 5341 35943 5342
rect 36016 5338 36054 5346
rect 36120 5370 36205 5376
rect 36225 5375 36262 5376
rect 36120 5350 36128 5370
rect 36148 5369 36205 5370
rect 36148 5350 36177 5369
rect 36120 5349 36177 5350
rect 36198 5349 36205 5369
rect 36120 5342 36205 5349
rect 36224 5366 36262 5375
rect 36224 5346 36233 5366
rect 36253 5346 36262 5366
rect 36120 5341 36156 5342
rect 36224 5338 36262 5346
rect 36328 5370 36472 5376
rect 36328 5350 36336 5370
rect 36356 5350 36444 5370
rect 36464 5350 36472 5370
rect 36328 5342 36472 5350
rect 36328 5341 36364 5342
rect 36436 5341 36472 5342
rect 36538 5375 36575 5376
rect 36538 5374 36576 5375
rect 36538 5366 36602 5374
rect 36538 5346 36547 5366
rect 36567 5352 36602 5366
rect 36622 5352 36625 5372
rect 36567 5347 36625 5352
rect 36567 5346 36602 5347
rect 35804 5309 35841 5338
rect 35805 5307 35841 5309
rect 36017 5307 36054 5338
rect 35805 5285 36054 5307
rect 35886 5279 35997 5285
rect 35886 5271 35927 5279
rect 35886 5251 35894 5271
rect 35913 5251 35927 5271
rect 35886 5249 35927 5251
rect 35955 5271 35997 5279
rect 35955 5251 35971 5271
rect 35990 5251 35997 5271
rect 35955 5249 35997 5251
rect 35886 5234 35997 5249
rect 36225 5217 36262 5338
rect 36538 5334 36602 5346
rect 36343 5217 36372 5221
rect 36642 5219 36669 5486
rect 36501 5217 36669 5219
rect 36225 5191 36669 5217
rect 36184 4923 36229 4932
rect 36184 4885 36194 4923
rect 36219 4885 36229 4923
rect 36184 4874 36229 4885
rect 36187 4866 36229 4874
rect 36187 4161 36230 4866
rect 36343 4252 36372 5191
rect 36501 5190 36669 5191
rect 37073 5041 37157 5045
rect 37625 5041 37713 7892
rect 38252 7879 38307 7891
rect 38252 7845 38270 7879
rect 38299 7845 38307 7879
rect 38252 7819 38307 7845
rect 37859 7786 38027 7787
rect 38252 7786 38269 7819
rect 37859 7785 38269 7786
rect 38298 7785 38307 7819
rect 37859 7760 38307 7785
rect 37859 7758 38027 7760
rect 37859 7491 37886 7758
rect 38252 7754 38307 7760
rect 37926 7631 37990 7643
rect 38266 7639 38303 7754
rect 38531 7728 38642 7743
rect 38531 7726 38573 7728
rect 38531 7706 38538 7726
rect 38557 7706 38573 7726
rect 38531 7698 38573 7706
rect 38601 7726 38642 7728
rect 38601 7706 38615 7726
rect 38634 7706 38642 7726
rect 38601 7698 38642 7706
rect 38531 7692 38642 7698
rect 38474 7670 38723 7692
rect 38474 7639 38511 7670
rect 38687 7668 38723 7670
rect 38687 7639 38724 7668
rect 37926 7630 37961 7631
rect 37903 7625 37961 7630
rect 37903 7605 37906 7625
rect 37926 7611 37961 7625
rect 37981 7611 37990 7631
rect 37926 7603 37990 7611
rect 37952 7602 37990 7603
rect 37953 7601 37990 7602
rect 38056 7635 38092 7636
rect 38164 7635 38200 7636
rect 38056 7627 38200 7635
rect 38056 7607 38064 7627
rect 38084 7607 38172 7627
rect 38192 7607 38200 7627
rect 38056 7601 38200 7607
rect 38266 7631 38304 7639
rect 38372 7635 38408 7636
rect 38266 7611 38275 7631
rect 38295 7611 38304 7631
rect 38266 7602 38304 7611
rect 38323 7628 38408 7635
rect 38323 7608 38330 7628
rect 38351 7627 38408 7628
rect 38351 7608 38380 7627
rect 38323 7607 38380 7608
rect 38400 7607 38408 7627
rect 38266 7601 38303 7602
rect 38323 7601 38408 7607
rect 38474 7631 38512 7639
rect 38585 7635 38621 7636
rect 38474 7611 38483 7631
rect 38503 7611 38512 7631
rect 38474 7602 38512 7611
rect 38536 7627 38621 7635
rect 38536 7607 38593 7627
rect 38613 7607 38621 7627
rect 38474 7601 38511 7602
rect 38536 7601 38621 7607
rect 38687 7631 38725 7639
rect 38687 7611 38696 7631
rect 38716 7611 38725 7631
rect 38687 7602 38725 7611
rect 38687 7601 38724 7602
rect 38110 7580 38146 7601
rect 38536 7580 38567 7601
rect 38781 7584 38852 8237
rect 39367 8171 39410 8884
rect 40027 8795 40122 8815
rect 40027 8751 40047 8795
rect 40107 8751 40122 8795
rect 40027 8455 40122 8751
rect 40027 8414 40060 8455
rect 40096 8414 40122 8455
rect 40222 8494 40284 8965
rect 41564 8905 41601 8906
rect 41867 8905 41904 9047
rect 41929 9067 42016 9074
rect 41929 9064 41987 9067
rect 41929 9044 41934 9064
rect 41955 9047 41987 9064
rect 42007 9047 42016 9067
rect 41955 9044 42016 9047
rect 41929 9037 42016 9044
rect 42075 9067 42112 9077
rect 42075 9047 42083 9067
rect 42103 9047 42112 9067
rect 41929 9036 41960 9037
rect 42075 8968 42112 9047
rect 42142 9076 42173 9129
rect 42386 9122 42401 9130
rect 42441 9122 42451 9159
rect 42386 9113 42451 9122
rect 42599 9120 42664 9141
rect 42599 9102 42624 9120
rect 42642 9102 42664 9120
rect 42192 9076 42229 9077
rect 42142 9067 42229 9076
rect 42142 9047 42200 9067
rect 42220 9047 42229 9067
rect 42142 9037 42229 9047
rect 42288 9067 42325 9077
rect 42288 9047 42296 9067
rect 42316 9047 42325 9067
rect 42142 9036 42173 9037
rect 42137 8968 42247 8981
rect 42288 8968 42325 9047
rect 42599 9026 42664 9102
rect 42075 8966 42325 8968
rect 42075 8963 42176 8966
rect 42075 8944 42140 8963
rect 42137 8936 42140 8944
rect 42169 8936 42176 8963
rect 42204 8939 42214 8966
rect 42243 8944 42325 8966
rect 42348 8991 42665 9026
rect 42243 8939 42247 8944
rect 42204 8936 42247 8939
rect 42137 8922 42247 8936
rect 41563 8904 41904 8905
rect 41488 8902 41904 8904
rect 42348 8902 42388 8991
rect 42599 8964 42664 8991
rect 42599 8946 42622 8964
rect 42640 8946 42664 8964
rect 42599 8926 42664 8946
rect 41485 8899 42388 8902
rect 41485 8879 41491 8899
rect 41511 8879 42388 8899
rect 41485 8875 42388 8879
rect 42348 8872 42388 8875
rect 42600 8865 42665 8886
rect 40818 8857 41479 8858
rect 40818 8850 41752 8857
rect 40818 8849 41724 8850
rect 40818 8829 41669 8849
rect 41701 8830 41724 8849
rect 41749 8830 41752 8850
rect 41701 8829 41752 8830
rect 40818 8822 41752 8829
rect 40417 8780 40585 8781
rect 40820 8780 40859 8822
rect 41648 8820 41752 8822
rect 41717 8818 41752 8820
rect 42600 8847 42624 8865
rect 42642 8847 42665 8865
rect 42600 8800 42665 8847
rect 40417 8754 40861 8780
rect 40417 8752 40585 8754
rect 40222 8475 40286 8494
rect 40222 8436 40239 8475
rect 40273 8436 40286 8475
rect 40222 8417 40286 8436
rect 40027 8388 40122 8414
rect 40417 8401 40444 8752
rect 40820 8748 40861 8754
rect 40484 8541 40548 8553
rect 40824 8549 40861 8748
rect 41323 8775 41395 8792
rect 41323 8736 41331 8775
rect 41376 8736 41395 8775
rect 41089 8638 41200 8653
rect 41089 8636 41131 8638
rect 41089 8616 41096 8636
rect 41115 8616 41131 8636
rect 41089 8608 41131 8616
rect 41159 8636 41200 8638
rect 41159 8616 41173 8636
rect 41192 8616 41200 8636
rect 41159 8608 41200 8616
rect 41089 8602 41200 8608
rect 41032 8580 41281 8602
rect 41032 8549 41069 8580
rect 41245 8578 41281 8580
rect 41245 8549 41282 8578
rect 40484 8540 40519 8541
rect 40461 8535 40519 8540
rect 40461 8515 40464 8535
rect 40484 8521 40519 8535
rect 40539 8521 40548 8541
rect 40484 8513 40548 8521
rect 40510 8512 40548 8513
rect 40511 8511 40548 8512
rect 40614 8545 40650 8546
rect 40722 8545 40758 8546
rect 40614 8537 40758 8545
rect 40614 8517 40622 8537
rect 40642 8517 40730 8537
rect 40750 8517 40758 8537
rect 40614 8511 40758 8517
rect 40824 8541 40862 8549
rect 40930 8545 40966 8546
rect 40824 8521 40833 8541
rect 40853 8521 40862 8541
rect 40824 8512 40862 8521
rect 40881 8538 40966 8545
rect 40881 8518 40888 8538
rect 40909 8537 40966 8538
rect 40909 8518 40938 8537
rect 40881 8517 40938 8518
rect 40958 8517 40966 8537
rect 40824 8511 40861 8512
rect 40881 8511 40966 8517
rect 41032 8541 41070 8549
rect 41143 8545 41179 8546
rect 41032 8521 41041 8541
rect 41061 8521 41070 8541
rect 41032 8512 41070 8521
rect 41094 8537 41179 8545
rect 41094 8517 41151 8537
rect 41171 8517 41179 8537
rect 41032 8511 41069 8512
rect 41094 8511 41179 8517
rect 41245 8541 41283 8549
rect 41245 8521 41254 8541
rect 41274 8521 41283 8541
rect 41245 8512 41283 8521
rect 41323 8526 41395 8736
rect 41465 8770 42665 8800
rect 41465 8769 41909 8770
rect 41465 8767 41633 8769
rect 41323 8512 41406 8526
rect 41245 8511 41282 8512
rect 40668 8490 40704 8511
rect 41094 8490 41125 8511
rect 41323 8490 41340 8512
rect 40501 8486 40601 8490
rect 40501 8482 40563 8486
rect 40501 8456 40508 8482
rect 40534 8460 40563 8482
rect 40589 8460 40601 8486
rect 40534 8456 40601 8460
rect 40501 8453 40601 8456
rect 40669 8453 40704 8490
rect 40766 8487 41125 8490
rect 40766 8482 40988 8487
rect 40766 8458 40779 8482
rect 40803 8463 40988 8482
rect 41012 8463 41125 8487
rect 40803 8458 41125 8463
rect 40766 8454 41125 8458
rect 41192 8482 41340 8490
rect 41192 8462 41203 8482
rect 41223 8479 41340 8482
rect 41393 8479 41406 8512
rect 41223 8462 41406 8479
rect 41192 8455 41406 8462
rect 41192 8454 41233 8455
rect 41323 8454 41406 8455
rect 40668 8428 40704 8453
rect 40516 8401 40553 8402
rect 40612 8401 40649 8402
rect 40668 8401 40675 8428
rect 40416 8392 40554 8401
rect 40416 8372 40525 8392
rect 40545 8372 40554 8392
rect 40416 8365 40554 8372
rect 40612 8398 40675 8401
rect 40696 8401 40704 8428
rect 40723 8401 40760 8402
rect 40696 8398 40760 8401
rect 40612 8392 40760 8398
rect 40612 8372 40621 8392
rect 40641 8372 40731 8392
rect 40751 8372 40760 8392
rect 40416 8363 40512 8365
rect 40612 8362 40760 8372
rect 40819 8392 40856 8402
rect 40931 8401 40968 8402
rect 40912 8399 40968 8401
rect 40819 8372 40827 8392
rect 40847 8372 40856 8392
rect 40668 8361 40704 8362
rect 40516 8230 40553 8231
rect 40819 8230 40856 8372
rect 40881 8392 40968 8399
rect 40881 8389 40939 8392
rect 40881 8369 40886 8389
rect 40907 8372 40939 8389
rect 40959 8372 40968 8392
rect 40907 8369 40968 8372
rect 40881 8362 40968 8369
rect 41027 8392 41064 8402
rect 41027 8372 41035 8392
rect 41055 8372 41064 8392
rect 40881 8361 40912 8362
rect 41027 8293 41064 8372
rect 41094 8401 41125 8454
rect 41331 8421 41345 8454
rect 41398 8421 41406 8454
rect 41331 8415 41406 8421
rect 41331 8410 41401 8415
rect 41144 8401 41181 8402
rect 41094 8392 41181 8401
rect 41094 8372 41152 8392
rect 41172 8372 41181 8392
rect 41094 8362 41181 8372
rect 41240 8392 41277 8402
rect 41465 8397 41492 8767
rect 41532 8537 41596 8549
rect 41872 8545 41909 8769
rect 42380 8750 42444 8752
rect 42376 8738 42444 8750
rect 42376 8705 42387 8738
rect 42427 8705 42444 8738
rect 42376 8695 42444 8705
rect 42137 8634 42248 8649
rect 42137 8632 42179 8634
rect 42137 8612 42144 8632
rect 42163 8612 42179 8632
rect 42137 8604 42179 8612
rect 42207 8632 42248 8634
rect 42207 8612 42221 8632
rect 42240 8612 42248 8632
rect 42207 8604 42248 8612
rect 42137 8598 42248 8604
rect 42080 8576 42329 8598
rect 42080 8545 42117 8576
rect 42293 8574 42329 8576
rect 42293 8545 42330 8574
rect 41532 8536 41567 8537
rect 41509 8531 41567 8536
rect 41509 8511 41512 8531
rect 41532 8517 41567 8531
rect 41587 8517 41596 8537
rect 41532 8509 41596 8517
rect 41558 8508 41596 8509
rect 41559 8507 41596 8508
rect 41662 8541 41698 8542
rect 41770 8541 41806 8542
rect 41662 8533 41806 8541
rect 41662 8513 41670 8533
rect 41690 8513 41778 8533
rect 41798 8513 41806 8533
rect 41662 8507 41806 8513
rect 41872 8537 41910 8545
rect 41978 8541 42014 8542
rect 41872 8517 41881 8537
rect 41901 8517 41910 8537
rect 41872 8508 41910 8517
rect 41929 8534 42014 8541
rect 41929 8514 41936 8534
rect 41957 8533 42014 8534
rect 41957 8514 41986 8533
rect 41929 8513 41986 8514
rect 42006 8513 42014 8533
rect 41872 8507 41909 8508
rect 41929 8507 42014 8513
rect 42080 8537 42118 8545
rect 42191 8541 42227 8542
rect 42080 8517 42089 8537
rect 42109 8517 42118 8537
rect 42080 8508 42118 8517
rect 42142 8533 42227 8541
rect 42142 8513 42199 8533
rect 42219 8513 42227 8533
rect 42080 8507 42117 8508
rect 42142 8507 42227 8513
rect 42293 8537 42331 8545
rect 42293 8517 42302 8537
rect 42322 8517 42331 8537
rect 42293 8508 42331 8517
rect 42380 8511 42444 8695
rect 42600 8569 42665 8770
rect 42600 8551 42622 8569
rect 42640 8551 42665 8569
rect 42600 8532 42665 8551
rect 42293 8507 42330 8508
rect 41716 8486 41752 8507
rect 42142 8486 42173 8507
rect 42380 8502 42388 8511
rect 42377 8486 42388 8502
rect 41549 8482 41649 8486
rect 41549 8478 41611 8482
rect 41549 8452 41556 8478
rect 41582 8456 41611 8478
rect 41637 8456 41649 8482
rect 41582 8452 41649 8456
rect 41549 8449 41649 8452
rect 41717 8449 41752 8486
rect 41814 8483 42173 8486
rect 41814 8478 42036 8483
rect 41814 8454 41827 8478
rect 41851 8459 42036 8478
rect 42060 8459 42173 8483
rect 41851 8454 42173 8459
rect 41814 8450 42173 8454
rect 42240 8478 42388 8486
rect 42240 8458 42251 8478
rect 42271 8469 42388 8478
rect 42437 8502 42444 8511
rect 42437 8469 42445 8502
rect 42271 8458 42445 8469
rect 42240 8451 42445 8458
rect 42240 8450 42281 8451
rect 41716 8424 41752 8449
rect 41564 8397 41601 8398
rect 41660 8397 41697 8398
rect 41716 8397 41723 8424
rect 41240 8372 41248 8392
rect 41268 8372 41277 8392
rect 41094 8361 41125 8362
rect 41089 8293 41199 8306
rect 41240 8293 41277 8372
rect 41464 8388 41602 8397
rect 41464 8368 41573 8388
rect 41593 8368 41602 8388
rect 41464 8361 41602 8368
rect 41660 8394 41723 8397
rect 41744 8397 41752 8424
rect 41771 8397 41808 8398
rect 41744 8394 41808 8397
rect 41660 8388 41808 8394
rect 41660 8368 41669 8388
rect 41689 8368 41779 8388
rect 41799 8368 41808 8388
rect 41464 8359 41560 8361
rect 41660 8358 41808 8368
rect 41867 8388 41904 8398
rect 41979 8397 42016 8398
rect 41960 8395 42016 8397
rect 41867 8368 41875 8388
rect 41895 8368 41904 8388
rect 41716 8357 41752 8358
rect 41027 8291 41277 8293
rect 41027 8288 41128 8291
rect 41027 8269 41092 8288
rect 41089 8261 41092 8269
rect 41121 8261 41128 8288
rect 41156 8264 41166 8291
rect 41195 8269 41277 8291
rect 41195 8264 41199 8269
rect 41156 8261 41199 8264
rect 41089 8247 41199 8261
rect 40515 8229 40856 8230
rect 40440 8224 40856 8229
rect 41564 8226 41601 8227
rect 41867 8226 41904 8368
rect 41929 8388 42016 8395
rect 41929 8385 41987 8388
rect 41929 8365 41934 8385
rect 41955 8368 41987 8385
rect 42007 8368 42016 8388
rect 41955 8365 42016 8368
rect 41929 8358 42016 8365
rect 42075 8388 42112 8398
rect 42075 8368 42083 8388
rect 42103 8368 42112 8388
rect 41929 8357 41960 8358
rect 42075 8289 42112 8368
rect 42142 8397 42173 8450
rect 42377 8448 42445 8451
rect 42377 8406 42389 8448
rect 42438 8406 42445 8448
rect 42192 8397 42229 8398
rect 42142 8388 42229 8397
rect 42142 8368 42200 8388
rect 42220 8368 42229 8388
rect 42142 8358 42229 8368
rect 42288 8388 42325 8398
rect 42377 8393 42445 8406
rect 42600 8470 42665 8487
rect 42600 8452 42624 8470
rect 42642 8452 42665 8470
rect 42288 8368 42296 8388
rect 42316 8368 42325 8388
rect 42142 8357 42173 8358
rect 42137 8289 42247 8302
rect 42288 8289 42325 8368
rect 42600 8313 42665 8452
rect 42600 8307 42622 8313
rect 42075 8287 42325 8289
rect 42075 8284 42176 8287
rect 42075 8265 42140 8284
rect 42137 8257 42140 8265
rect 42169 8257 42176 8284
rect 42204 8260 42214 8287
rect 42243 8265 42325 8287
rect 42354 8295 42622 8307
rect 42640 8295 42665 8313
rect 42354 8272 42665 8295
rect 42354 8271 42409 8272
rect 42243 8260 42247 8265
rect 42204 8257 42247 8260
rect 42137 8243 42247 8257
rect 41563 8225 41904 8226
rect 40440 8204 40443 8224
rect 40463 8204 40856 8224
rect 41488 8224 41904 8225
rect 42354 8224 42397 8271
rect 41488 8220 42397 8224
rect 39363 8169 40074 8171
rect 40613 8169 40702 8172
rect 39363 8160 40702 8169
rect 39363 8122 40625 8160
rect 40650 8125 40669 8160
rect 40694 8125 40702 8160
rect 40807 8171 40852 8204
rect 41488 8200 41491 8220
rect 41511 8200 42397 8220
rect 41865 8195 42397 8200
rect 42605 8214 42664 8236
rect 42605 8196 42624 8214
rect 42642 8196 42664 8214
rect 41653 8171 41752 8173
rect 40807 8161 41752 8171
rect 40807 8135 41675 8161
rect 40808 8134 41675 8135
rect 40650 8122 40702 8125
rect 39363 8114 40702 8122
rect 41653 8123 41675 8134
rect 41700 8126 41719 8161
rect 41744 8126 41752 8161
rect 41700 8123 41752 8126
rect 41653 8115 41752 8123
rect 42605 8122 42664 8196
rect 41679 8114 41751 8115
rect 39363 8113 40701 8114
rect 39363 8111 40074 8113
rect 40223 8072 40287 8076
rect 42598 8074 42664 8122
rect 40223 8063 40297 8072
rect 38738 7580 38852 7584
rect 37943 7576 38043 7580
rect 37943 7572 38005 7576
rect 37943 7546 37950 7572
rect 37976 7550 38005 7572
rect 38031 7550 38043 7576
rect 37976 7546 38043 7550
rect 37943 7543 38043 7546
rect 38111 7543 38146 7580
rect 38208 7577 38567 7580
rect 38208 7572 38430 7577
rect 38208 7548 38221 7572
rect 38245 7553 38430 7572
rect 38454 7553 38567 7577
rect 38245 7548 38567 7553
rect 38208 7544 38567 7548
rect 38634 7577 38852 7580
rect 38634 7576 38817 7577
rect 38634 7572 38760 7576
rect 38634 7552 38645 7572
rect 38665 7552 38760 7572
rect 38784 7553 38817 7576
rect 38841 7553 38852 7577
rect 38784 7552 38852 7553
rect 38634 7545 38852 7552
rect 38634 7544 38675 7545
rect 38110 7518 38146 7543
rect 37958 7491 37995 7492
rect 38054 7491 38091 7492
rect 38110 7491 38117 7518
rect 37858 7482 37996 7491
rect 37858 7462 37967 7482
rect 37987 7462 37996 7482
rect 37858 7455 37996 7462
rect 38054 7488 38117 7491
rect 38138 7491 38146 7518
rect 38165 7491 38202 7492
rect 38138 7488 38202 7491
rect 38054 7482 38202 7488
rect 38054 7462 38063 7482
rect 38083 7462 38173 7482
rect 38193 7462 38202 7482
rect 37858 7453 37954 7455
rect 38054 7452 38202 7462
rect 38261 7482 38298 7492
rect 38373 7491 38410 7492
rect 38354 7489 38410 7491
rect 38261 7462 38269 7482
rect 38289 7462 38298 7482
rect 38110 7451 38146 7452
rect 37958 7320 37995 7321
rect 38261 7320 38298 7462
rect 38323 7482 38410 7489
rect 38323 7479 38381 7482
rect 38323 7459 38328 7479
rect 38349 7462 38381 7479
rect 38401 7462 38410 7482
rect 38349 7459 38410 7462
rect 38323 7452 38410 7459
rect 38469 7482 38506 7492
rect 38469 7462 38477 7482
rect 38497 7462 38506 7482
rect 38323 7451 38354 7452
rect 38469 7383 38506 7462
rect 38536 7491 38567 7544
rect 38738 7542 38852 7545
rect 38781 7510 38852 7542
rect 40027 8021 40111 8046
rect 40027 7993 40042 8021
rect 40086 7993 40111 8021
rect 40027 7964 40111 7993
rect 40223 8015 40237 8063
rect 40274 8015 40297 8063
rect 40223 7987 40297 8015
rect 40027 7936 40039 7964
rect 40083 7936 40111 7964
rect 40027 7915 40111 7936
rect 38586 7491 38623 7492
rect 38536 7482 38623 7491
rect 38536 7462 38594 7482
rect 38614 7462 38623 7482
rect 38536 7452 38623 7462
rect 38682 7482 38719 7492
rect 38682 7462 38690 7482
rect 38710 7462 38719 7482
rect 38536 7451 38567 7452
rect 38531 7383 38641 7396
rect 38682 7383 38719 7462
rect 38469 7381 38719 7383
rect 38469 7378 38570 7381
rect 38469 7359 38534 7378
rect 38531 7351 38534 7359
rect 38563 7351 38570 7378
rect 38598 7354 38608 7381
rect 38637 7359 38719 7381
rect 38637 7354 38641 7359
rect 38598 7351 38641 7354
rect 38531 7337 38641 7351
rect 37957 7319 38298 7320
rect 37882 7316 38298 7319
rect 37882 7314 38305 7316
rect 37882 7294 37885 7314
rect 37905 7294 38305 7314
rect 37073 4953 37713 5041
rect 37073 4602 37157 4953
rect 37639 4922 37683 4928
rect 37639 4896 37647 4922
rect 37672 4896 37683 4922
rect 37639 4847 37683 4896
rect 37639 4827 38036 4847
rect 38056 4827 38059 4847
rect 37639 4822 38059 4827
rect 37639 4821 37984 4822
rect 37639 4817 37683 4821
rect 37946 4820 37983 4821
rect 37300 4790 37410 4804
rect 37300 4787 37343 4790
rect 37300 4782 37304 4787
rect 37222 4760 37304 4782
rect 37333 4760 37343 4787
rect 37371 4763 37378 4790
rect 37407 4782 37410 4790
rect 37407 4763 37472 4782
rect 37371 4760 37472 4763
rect 37222 4758 37472 4760
rect 37222 4679 37259 4758
rect 37300 4745 37410 4758
rect 37374 4689 37405 4690
rect 37222 4659 37231 4679
rect 37251 4659 37259 4679
rect 37222 4649 37259 4659
rect 37318 4679 37405 4689
rect 37318 4659 37327 4679
rect 37347 4659 37405 4679
rect 37318 4650 37405 4659
rect 37318 4649 37355 4650
rect 37073 4596 37182 4602
rect 37374 4597 37405 4650
rect 37435 4679 37472 4758
rect 37587 4689 37618 4690
rect 37435 4659 37444 4679
rect 37464 4659 37472 4679
rect 37435 4649 37472 4659
rect 37531 4682 37618 4689
rect 37531 4679 37592 4682
rect 37531 4659 37540 4679
rect 37560 4662 37592 4679
rect 37613 4662 37618 4682
rect 37560 4659 37618 4662
rect 37531 4652 37618 4659
rect 37643 4679 37680 4817
rect 37795 4689 37831 4690
rect 37643 4659 37652 4679
rect 37672 4659 37680 4679
rect 37531 4650 37587 4652
rect 37531 4649 37568 4650
rect 37643 4649 37680 4659
rect 37739 4679 37887 4689
rect 37987 4686 38083 4688
rect 37739 4659 37748 4679
rect 37768 4659 37858 4679
rect 37878 4659 37887 4679
rect 37739 4653 37887 4659
rect 37739 4650 37803 4653
rect 37739 4649 37776 4650
rect 37795 4623 37803 4650
rect 37824 4650 37887 4653
rect 37945 4679 38083 4686
rect 37945 4659 37954 4679
rect 37974 4659 38083 4679
rect 37945 4650 38083 4659
rect 37824 4623 37831 4650
rect 37850 4649 37887 4650
rect 37946 4649 37983 4650
rect 37795 4598 37831 4623
rect 37266 4596 37307 4597
rect 37073 4589 37307 4596
rect 37073 4569 37276 4589
rect 37296 4569 37307 4589
rect 37073 4561 37307 4569
rect 37374 4593 37733 4597
rect 37374 4588 37696 4593
rect 37374 4564 37487 4588
rect 37511 4569 37696 4588
rect 37720 4569 37733 4593
rect 37511 4564 37733 4569
rect 37374 4561 37733 4564
rect 37795 4561 37830 4598
rect 37898 4595 37998 4598
rect 37898 4591 37965 4595
rect 37898 4565 37910 4591
rect 37936 4569 37965 4591
rect 37991 4569 37998 4595
rect 37936 4565 37998 4569
rect 37898 4561 37998 4565
rect 37073 4543 37182 4561
rect 37374 4540 37405 4561
rect 37795 4540 37831 4561
rect 37217 4539 37254 4540
rect 37216 4530 37254 4539
rect 37216 4510 37225 4530
rect 37245 4510 37254 4530
rect 37216 4502 37254 4510
rect 37320 4534 37405 4540
rect 37430 4539 37467 4540
rect 37320 4514 37328 4534
rect 37348 4514 37405 4534
rect 37320 4506 37405 4514
rect 37429 4530 37467 4539
rect 37429 4510 37438 4530
rect 37458 4510 37467 4530
rect 37320 4505 37356 4506
rect 37429 4502 37467 4510
rect 37533 4534 37618 4540
rect 37638 4539 37675 4540
rect 37533 4514 37541 4534
rect 37561 4533 37618 4534
rect 37561 4514 37590 4533
rect 37533 4513 37590 4514
rect 37611 4513 37618 4533
rect 37533 4506 37618 4513
rect 37637 4530 37675 4539
rect 37637 4510 37646 4530
rect 37666 4510 37675 4530
rect 37533 4505 37569 4506
rect 37637 4502 37675 4510
rect 37741 4535 37885 4540
rect 37741 4534 37794 4535
rect 37741 4514 37749 4534
rect 37769 4515 37794 4534
rect 37827 4534 37885 4535
rect 37827 4515 37857 4534
rect 37769 4514 37857 4515
rect 37877 4514 37885 4534
rect 37741 4506 37885 4514
rect 37741 4505 37777 4506
rect 37849 4505 37885 4506
rect 37951 4539 37988 4540
rect 37951 4538 37989 4539
rect 37951 4530 38015 4538
rect 37951 4510 37960 4530
rect 37980 4516 38015 4530
rect 38035 4516 38038 4536
rect 37980 4511 38038 4516
rect 37980 4510 38015 4511
rect 37217 4473 37254 4502
rect 37218 4471 37254 4473
rect 37430 4471 37467 4502
rect 37218 4449 37467 4471
rect 37299 4443 37410 4449
rect 37299 4435 37340 4443
rect 37299 4415 37307 4435
rect 37326 4415 37340 4435
rect 37299 4413 37340 4415
rect 37368 4435 37410 4443
rect 37368 4415 37384 4435
rect 37403 4415 37410 4435
rect 37368 4413 37410 4415
rect 37299 4398 37410 4413
rect 37638 4381 37675 4502
rect 37951 4498 38015 4510
rect 38055 4387 38082 4650
rect 38109 4396 38145 4403
rect 38109 4387 38115 4396
rect 38033 4383 38115 4387
rect 37914 4381 38115 4383
rect 37638 4358 38115 4381
rect 38138 4358 38145 4396
rect 37638 4355 38145 4358
rect 37914 4354 38082 4355
rect 38109 4352 38145 4355
rect 38227 4254 38305 7294
rect 39361 6547 39420 6557
rect 39361 6519 39374 6547
rect 39402 6519 39420 6547
rect 39361 6470 39420 6519
rect 38967 6335 39135 6336
rect 39371 6335 39418 6470
rect 38967 6309 39418 6335
rect 38967 6307 39135 6309
rect 38967 6040 38994 6307
rect 39371 6303 39418 6309
rect 39034 6180 39098 6192
rect 39374 6188 39411 6303
rect 39639 6277 39750 6292
rect 39639 6275 39681 6277
rect 39639 6255 39646 6275
rect 39665 6255 39681 6275
rect 39639 6247 39681 6255
rect 39709 6275 39750 6277
rect 39709 6255 39723 6275
rect 39742 6255 39750 6275
rect 39709 6247 39750 6255
rect 39639 6241 39750 6247
rect 39582 6219 39831 6241
rect 39582 6188 39619 6219
rect 39795 6217 39831 6219
rect 39795 6188 39832 6217
rect 39034 6179 39069 6180
rect 39011 6174 39069 6179
rect 39011 6154 39014 6174
rect 39034 6160 39069 6174
rect 39089 6160 39098 6180
rect 39034 6152 39098 6160
rect 39060 6151 39098 6152
rect 39061 6150 39098 6151
rect 39164 6184 39200 6185
rect 39272 6184 39308 6185
rect 39164 6176 39308 6184
rect 39164 6156 39172 6176
rect 39192 6156 39280 6176
rect 39300 6156 39308 6176
rect 39164 6150 39308 6156
rect 39374 6180 39412 6188
rect 39480 6184 39516 6185
rect 39374 6160 39383 6180
rect 39403 6160 39412 6180
rect 39374 6151 39412 6160
rect 39431 6177 39516 6184
rect 39431 6157 39438 6177
rect 39459 6176 39516 6177
rect 39459 6157 39488 6176
rect 39431 6156 39488 6157
rect 39508 6156 39516 6176
rect 39374 6150 39411 6151
rect 39431 6150 39516 6156
rect 39582 6180 39620 6188
rect 39693 6184 39729 6185
rect 39582 6160 39591 6180
rect 39611 6160 39620 6180
rect 39582 6151 39620 6160
rect 39644 6176 39729 6184
rect 39644 6156 39701 6176
rect 39721 6156 39729 6176
rect 39582 6150 39619 6151
rect 39644 6150 39729 6156
rect 39795 6180 39833 6188
rect 39795 6160 39804 6180
rect 39824 6160 39833 6180
rect 39795 6151 39833 6160
rect 39795 6150 39832 6151
rect 39218 6129 39254 6150
rect 39644 6129 39675 6150
rect 39855 6135 39912 6143
rect 39855 6129 39863 6135
rect 39051 6125 39151 6129
rect 39051 6121 39113 6125
rect 39051 6095 39058 6121
rect 39084 6099 39113 6121
rect 39139 6099 39151 6125
rect 39084 6095 39151 6099
rect 39051 6092 39151 6095
rect 39219 6092 39254 6129
rect 39316 6126 39675 6129
rect 39316 6121 39538 6126
rect 39316 6097 39329 6121
rect 39353 6102 39538 6121
rect 39562 6102 39675 6126
rect 39353 6097 39675 6102
rect 39316 6093 39675 6097
rect 39742 6121 39863 6129
rect 39742 6101 39753 6121
rect 39773 6112 39863 6121
rect 39889 6112 39912 6135
rect 39773 6101 39912 6112
rect 39742 6099 39912 6101
rect 39742 6094 39863 6099
rect 39742 6093 39783 6094
rect 39218 6067 39254 6092
rect 39066 6040 39103 6041
rect 39162 6040 39199 6041
rect 39218 6040 39225 6067
rect 38966 6031 39104 6040
rect 38966 6011 39075 6031
rect 39095 6011 39104 6031
rect 38966 6004 39104 6011
rect 39162 6037 39225 6040
rect 39246 6040 39254 6067
rect 39273 6040 39310 6041
rect 39246 6037 39310 6040
rect 39162 6031 39310 6037
rect 39162 6011 39171 6031
rect 39191 6011 39281 6031
rect 39301 6011 39310 6031
rect 38966 6002 39062 6004
rect 39162 6001 39310 6011
rect 39369 6031 39406 6041
rect 39481 6040 39518 6041
rect 39462 6038 39518 6040
rect 39369 6011 39377 6031
rect 39397 6011 39406 6031
rect 39218 6000 39254 6001
rect 39066 5869 39103 5870
rect 39369 5869 39406 6011
rect 39431 6031 39518 6038
rect 39431 6028 39489 6031
rect 39431 6008 39436 6028
rect 39457 6011 39489 6028
rect 39509 6011 39518 6031
rect 39457 6008 39518 6011
rect 39431 6001 39518 6008
rect 39577 6031 39614 6041
rect 39577 6011 39585 6031
rect 39605 6011 39614 6031
rect 39431 6000 39462 6001
rect 39577 5932 39614 6011
rect 39644 6040 39675 6093
rect 39694 6040 39731 6041
rect 39644 6031 39731 6040
rect 39644 6011 39702 6031
rect 39722 6011 39731 6031
rect 39644 6001 39731 6011
rect 39790 6031 39827 6041
rect 39790 6011 39798 6031
rect 39818 6011 39827 6031
rect 39644 6000 39675 6001
rect 39639 5932 39749 5945
rect 39790 5932 39827 6011
rect 39577 5930 39827 5932
rect 39577 5927 39678 5930
rect 39577 5908 39642 5927
rect 39639 5900 39642 5908
rect 39671 5900 39678 5927
rect 39706 5903 39716 5930
rect 39745 5908 39827 5930
rect 39745 5903 39749 5908
rect 39706 5900 39749 5903
rect 39639 5886 39749 5900
rect 39065 5868 39406 5869
rect 38990 5863 39406 5868
rect 38990 5843 38993 5863
rect 39013 5843 39407 5863
rect 39216 5810 39253 5820
rect 39216 5773 39225 5810
rect 39242 5773 39253 5810
rect 39216 5752 39253 5773
rect 38925 4813 39093 4814
rect 39222 4813 39251 5752
rect 39364 5138 39407 5843
rect 39365 5130 39407 5138
rect 39365 5119 39410 5130
rect 39365 5081 39375 5119
rect 39400 5081 39410 5119
rect 39365 5072 39410 5081
rect 38925 4787 39369 4813
rect 38925 4785 39093 4787
rect 38925 4518 38952 4785
rect 39222 4783 39251 4787
rect 38992 4658 39056 4670
rect 39332 4666 39369 4787
rect 39597 4755 39708 4770
rect 39597 4753 39639 4755
rect 39597 4733 39604 4753
rect 39623 4733 39639 4753
rect 39597 4725 39639 4733
rect 39667 4753 39708 4755
rect 39667 4733 39681 4753
rect 39700 4733 39708 4753
rect 39667 4725 39708 4733
rect 39597 4719 39708 4725
rect 39540 4697 39789 4719
rect 39540 4666 39577 4697
rect 39753 4695 39789 4697
rect 39753 4666 39790 4695
rect 38992 4657 39027 4658
rect 38969 4652 39027 4657
rect 38969 4632 38972 4652
rect 38992 4638 39027 4652
rect 39047 4638 39056 4658
rect 38992 4630 39056 4638
rect 39018 4629 39056 4630
rect 39019 4628 39056 4629
rect 39122 4662 39158 4663
rect 39230 4662 39266 4663
rect 39122 4654 39266 4662
rect 39122 4634 39130 4654
rect 39150 4634 39238 4654
rect 39258 4634 39266 4654
rect 39122 4628 39266 4634
rect 39332 4658 39370 4666
rect 39438 4662 39474 4663
rect 39332 4638 39341 4658
rect 39361 4638 39370 4658
rect 39332 4629 39370 4638
rect 39389 4655 39474 4662
rect 39389 4635 39396 4655
rect 39417 4654 39474 4655
rect 39417 4635 39446 4654
rect 39389 4634 39446 4635
rect 39466 4634 39474 4654
rect 39332 4628 39369 4629
rect 39389 4628 39474 4634
rect 39540 4658 39578 4666
rect 39651 4662 39687 4663
rect 39540 4638 39549 4658
rect 39569 4638 39578 4658
rect 39540 4629 39578 4638
rect 39602 4654 39687 4662
rect 39602 4634 39659 4654
rect 39679 4634 39687 4654
rect 39540 4628 39577 4629
rect 39602 4628 39687 4634
rect 39753 4658 39791 4666
rect 39753 4638 39762 4658
rect 39782 4638 39791 4658
rect 39753 4629 39791 4638
rect 39753 4628 39790 4629
rect 39176 4607 39212 4628
rect 39602 4607 39633 4628
rect 40027 4611 40119 7915
rect 40225 6148 40297 7987
rect 41327 7937 41399 7954
rect 41327 7889 41339 7937
rect 41385 7889 41399 7937
rect 41867 7917 41908 7919
rect 42139 7917 42243 7919
rect 42598 7917 42663 8074
rect 41327 7867 41399 7889
rect 41460 7882 42663 7917
rect 41460 7868 41488 7882
rect 41328 7667 41398 7867
rect 41462 7737 41488 7868
rect 41867 7879 42663 7882
rect 41320 7616 41400 7667
rect 41320 7590 41336 7616
rect 41376 7590 41400 7616
rect 41320 7571 41400 7590
rect 41320 7545 41339 7571
rect 41379 7545 41400 7571
rect 41320 7518 41400 7545
rect 41320 7492 41343 7518
rect 41383 7492 41400 7518
rect 41320 7481 41400 7492
rect 41462 7482 41489 7737
rect 41867 7729 41908 7879
rect 42139 7877 42243 7879
rect 42598 7845 42663 7879
rect 42334 7817 42455 7835
rect 42334 7815 42405 7817
rect 42334 7774 42349 7815
rect 42386 7776 42405 7815
rect 42442 7776 42455 7817
rect 42386 7774 42455 7776
rect 42334 7764 42455 7774
rect 42139 7734 42243 7737
rect 41529 7622 41593 7634
rect 41869 7630 41906 7729
rect 42134 7719 42245 7734
rect 42134 7717 42176 7719
rect 42134 7697 42141 7717
rect 42160 7697 42176 7717
rect 42134 7689 42176 7697
rect 42204 7717 42245 7719
rect 42204 7697 42218 7717
rect 42237 7697 42245 7717
rect 42204 7689 42245 7697
rect 42134 7683 42245 7689
rect 42077 7661 42326 7683
rect 42077 7630 42114 7661
rect 42290 7659 42326 7661
rect 42290 7630 42327 7659
rect 41529 7621 41564 7622
rect 41506 7616 41564 7621
rect 41506 7596 41509 7616
rect 41529 7602 41564 7616
rect 41584 7602 41593 7622
rect 41529 7594 41593 7602
rect 41555 7593 41593 7594
rect 41556 7592 41593 7593
rect 41659 7626 41695 7627
rect 41767 7626 41803 7627
rect 41659 7618 41803 7626
rect 41659 7598 41667 7618
rect 41687 7598 41775 7618
rect 41795 7598 41803 7618
rect 41659 7592 41803 7598
rect 41869 7622 41907 7630
rect 41975 7626 42011 7627
rect 41869 7602 41878 7622
rect 41898 7602 41907 7622
rect 41869 7593 41907 7602
rect 41926 7619 42011 7626
rect 41926 7599 41933 7619
rect 41954 7618 42011 7619
rect 41954 7599 41983 7618
rect 41926 7598 41983 7599
rect 42003 7598 42011 7618
rect 41869 7592 41906 7593
rect 41926 7592 42011 7598
rect 42077 7622 42115 7630
rect 42188 7626 42224 7627
rect 42077 7602 42086 7622
rect 42106 7602 42115 7622
rect 42077 7593 42115 7602
rect 42139 7618 42224 7626
rect 42139 7598 42196 7618
rect 42216 7598 42224 7618
rect 42077 7592 42114 7593
rect 42139 7592 42224 7598
rect 42290 7622 42328 7630
rect 42290 7602 42299 7622
rect 42319 7602 42328 7622
rect 42383 7612 42448 7764
rect 42601 7738 42656 7845
rect 42290 7593 42328 7602
rect 42381 7605 42448 7612
rect 42290 7592 42327 7593
rect 41713 7571 41749 7592
rect 42139 7571 42170 7592
rect 42381 7584 42398 7605
rect 42434 7584 42448 7605
rect 42600 7625 42656 7738
rect 42600 7607 42619 7625
rect 42637 7607 42656 7625
rect 42600 7587 42656 7607
rect 42381 7571 42448 7584
rect 41546 7567 41646 7571
rect 41546 7563 41608 7567
rect 41546 7537 41553 7563
rect 41579 7541 41608 7563
rect 41634 7541 41646 7567
rect 41579 7537 41646 7541
rect 41546 7534 41646 7537
rect 41714 7534 41749 7571
rect 41811 7568 42170 7571
rect 41811 7563 42033 7568
rect 41811 7539 41824 7563
rect 41848 7544 42033 7563
rect 42057 7544 42170 7568
rect 41848 7539 42170 7544
rect 41811 7535 42170 7539
rect 42237 7565 42448 7571
rect 42237 7563 42398 7565
rect 42237 7543 42248 7563
rect 42268 7543 42398 7563
rect 42237 7536 42398 7543
rect 42237 7535 42278 7536
rect 41713 7509 41749 7534
rect 41561 7482 41598 7483
rect 41657 7482 41694 7483
rect 41713 7482 41720 7509
rect 41461 7473 41599 7482
rect 41461 7453 41570 7473
rect 41590 7453 41599 7473
rect 41461 7446 41599 7453
rect 41657 7479 41720 7482
rect 41741 7482 41749 7509
rect 41768 7482 41805 7483
rect 41741 7479 41805 7482
rect 41657 7473 41805 7479
rect 41657 7453 41666 7473
rect 41686 7453 41776 7473
rect 41796 7453 41805 7473
rect 41461 7444 41557 7446
rect 41657 7443 41805 7453
rect 41864 7473 41901 7483
rect 41976 7482 42013 7483
rect 41957 7480 42013 7482
rect 41864 7453 41872 7473
rect 41892 7453 41901 7473
rect 41713 7442 41749 7443
rect 41561 7311 41598 7312
rect 41864 7311 41901 7453
rect 41926 7473 42013 7480
rect 41926 7470 41984 7473
rect 41926 7450 41931 7470
rect 41952 7453 41984 7470
rect 42004 7453 42013 7473
rect 41952 7450 42013 7453
rect 41926 7443 42013 7450
rect 42072 7473 42109 7483
rect 42072 7453 42080 7473
rect 42100 7453 42109 7473
rect 41926 7442 41957 7443
rect 42072 7374 42109 7453
rect 42139 7482 42170 7535
rect 42383 7528 42398 7536
rect 42438 7528 42448 7565
rect 42383 7519 42448 7528
rect 42596 7526 42661 7547
rect 42596 7508 42621 7526
rect 42639 7508 42661 7526
rect 42189 7482 42226 7483
rect 42139 7473 42226 7482
rect 42139 7453 42197 7473
rect 42217 7453 42226 7473
rect 42139 7443 42226 7453
rect 42285 7473 42322 7483
rect 42285 7453 42293 7473
rect 42313 7453 42322 7473
rect 42139 7442 42170 7443
rect 42134 7374 42244 7387
rect 42285 7374 42322 7453
rect 42596 7432 42661 7508
rect 42072 7372 42322 7374
rect 42072 7369 42173 7372
rect 42072 7350 42137 7369
rect 42134 7342 42137 7350
rect 42166 7342 42173 7369
rect 42201 7345 42211 7372
rect 42240 7350 42322 7372
rect 42345 7397 42662 7432
rect 42240 7345 42244 7350
rect 42201 7342 42244 7345
rect 42134 7328 42244 7342
rect 41560 7310 41901 7311
rect 41485 7308 41901 7310
rect 42345 7308 42385 7397
rect 42596 7370 42661 7397
rect 42596 7352 42619 7370
rect 42637 7352 42661 7370
rect 42596 7332 42661 7352
rect 41482 7305 42385 7308
rect 41482 7285 41488 7305
rect 41508 7285 42385 7305
rect 41482 7281 42385 7285
rect 42345 7278 42385 7281
rect 42597 7271 42662 7292
rect 40815 7263 41476 7264
rect 40815 7256 41749 7263
rect 40815 7255 41721 7256
rect 40815 7235 41666 7255
rect 41698 7236 41721 7255
rect 41746 7236 41749 7256
rect 41698 7235 41749 7236
rect 40815 7228 41749 7235
rect 40414 7186 40582 7187
rect 40817 7186 40856 7228
rect 41645 7226 41749 7228
rect 41714 7224 41749 7226
rect 42597 7253 42621 7271
rect 42639 7253 42662 7271
rect 42597 7206 42662 7253
rect 40414 7160 40858 7186
rect 40414 7158 40582 7160
rect 40414 6807 40441 7158
rect 40817 7154 40858 7160
rect 40481 6947 40545 6959
rect 40821 6955 40858 7154
rect 41320 7181 41392 7198
rect 41320 7142 41328 7181
rect 41373 7142 41392 7181
rect 41086 7044 41197 7059
rect 41086 7042 41128 7044
rect 41086 7022 41093 7042
rect 41112 7022 41128 7042
rect 41086 7014 41128 7022
rect 41156 7042 41197 7044
rect 41156 7022 41170 7042
rect 41189 7022 41197 7042
rect 41156 7014 41197 7022
rect 41086 7008 41197 7014
rect 41029 6986 41278 7008
rect 41029 6955 41066 6986
rect 41242 6984 41278 6986
rect 41242 6955 41279 6984
rect 40481 6946 40516 6947
rect 40458 6941 40516 6946
rect 40458 6921 40461 6941
rect 40481 6927 40516 6941
rect 40536 6927 40545 6947
rect 40481 6919 40545 6927
rect 40507 6918 40545 6919
rect 40508 6917 40545 6918
rect 40611 6951 40647 6952
rect 40719 6951 40755 6952
rect 40611 6943 40755 6951
rect 40611 6923 40619 6943
rect 40639 6923 40727 6943
rect 40747 6923 40755 6943
rect 40611 6917 40755 6923
rect 40821 6947 40859 6955
rect 40927 6951 40963 6952
rect 40821 6927 40830 6947
rect 40850 6927 40859 6947
rect 40821 6918 40859 6927
rect 40878 6944 40963 6951
rect 40878 6924 40885 6944
rect 40906 6943 40963 6944
rect 40906 6924 40935 6943
rect 40878 6923 40935 6924
rect 40955 6923 40963 6943
rect 40821 6917 40858 6918
rect 40878 6917 40963 6923
rect 41029 6947 41067 6955
rect 41140 6951 41176 6952
rect 41029 6927 41038 6947
rect 41058 6927 41067 6947
rect 41029 6918 41067 6927
rect 41091 6943 41176 6951
rect 41091 6923 41148 6943
rect 41168 6923 41176 6943
rect 41029 6917 41066 6918
rect 41091 6917 41176 6923
rect 41242 6947 41280 6955
rect 41242 6927 41251 6947
rect 41271 6927 41280 6947
rect 41242 6918 41280 6927
rect 41320 6932 41392 7142
rect 41462 7176 42662 7206
rect 41462 7175 41906 7176
rect 41462 7173 41630 7175
rect 41320 6918 41403 6932
rect 41242 6917 41279 6918
rect 40665 6896 40701 6917
rect 41091 6896 41122 6917
rect 41320 6896 41337 6918
rect 40498 6892 40598 6896
rect 40498 6888 40560 6892
rect 40498 6862 40505 6888
rect 40531 6866 40560 6888
rect 40586 6866 40598 6892
rect 40531 6862 40598 6866
rect 40498 6859 40598 6862
rect 40666 6859 40701 6896
rect 40763 6893 41122 6896
rect 40763 6888 40985 6893
rect 40763 6864 40776 6888
rect 40800 6869 40985 6888
rect 41009 6869 41122 6893
rect 40800 6864 41122 6869
rect 40763 6860 41122 6864
rect 41189 6888 41337 6896
rect 41189 6868 41200 6888
rect 41220 6885 41337 6888
rect 41390 6885 41403 6918
rect 41220 6868 41403 6885
rect 41189 6861 41403 6868
rect 41189 6860 41230 6861
rect 41320 6860 41403 6861
rect 40665 6834 40701 6859
rect 40513 6807 40550 6808
rect 40609 6807 40646 6808
rect 40665 6807 40672 6834
rect 40413 6798 40551 6807
rect 40413 6778 40522 6798
rect 40542 6778 40551 6798
rect 40413 6771 40551 6778
rect 40609 6804 40672 6807
rect 40693 6807 40701 6834
rect 40720 6807 40757 6808
rect 40693 6804 40757 6807
rect 40609 6798 40757 6804
rect 40609 6778 40618 6798
rect 40638 6778 40728 6798
rect 40748 6778 40757 6798
rect 40413 6769 40509 6771
rect 40609 6768 40757 6778
rect 40816 6798 40853 6808
rect 40928 6807 40965 6808
rect 40909 6805 40965 6807
rect 40816 6778 40824 6798
rect 40844 6778 40853 6798
rect 40665 6767 40701 6768
rect 40513 6636 40550 6637
rect 40816 6636 40853 6778
rect 40878 6798 40965 6805
rect 40878 6795 40936 6798
rect 40878 6775 40883 6795
rect 40904 6778 40936 6795
rect 40956 6778 40965 6798
rect 40904 6775 40965 6778
rect 40878 6768 40965 6775
rect 41024 6798 41061 6808
rect 41024 6778 41032 6798
rect 41052 6778 41061 6798
rect 40878 6767 40909 6768
rect 41024 6699 41061 6778
rect 41091 6807 41122 6860
rect 41328 6827 41342 6860
rect 41395 6827 41403 6860
rect 41328 6821 41403 6827
rect 41328 6816 41398 6821
rect 41141 6807 41178 6808
rect 41091 6798 41178 6807
rect 41091 6778 41149 6798
rect 41169 6778 41178 6798
rect 41091 6768 41178 6778
rect 41237 6798 41274 6808
rect 41462 6803 41489 7173
rect 41529 6943 41593 6955
rect 41869 6951 41906 7175
rect 42377 7156 42441 7158
rect 42373 7144 42441 7156
rect 42373 7111 42384 7144
rect 42424 7111 42441 7144
rect 42373 7101 42441 7111
rect 42134 7040 42245 7055
rect 42134 7038 42176 7040
rect 42134 7018 42141 7038
rect 42160 7018 42176 7038
rect 42134 7010 42176 7018
rect 42204 7038 42245 7040
rect 42204 7018 42218 7038
rect 42237 7018 42245 7038
rect 42204 7010 42245 7018
rect 42134 7004 42245 7010
rect 42077 6982 42326 7004
rect 42077 6951 42114 6982
rect 42290 6980 42326 6982
rect 42290 6951 42327 6980
rect 41529 6942 41564 6943
rect 41506 6937 41564 6942
rect 41506 6917 41509 6937
rect 41529 6923 41564 6937
rect 41584 6923 41593 6943
rect 41529 6915 41593 6923
rect 41555 6914 41593 6915
rect 41556 6913 41593 6914
rect 41659 6947 41695 6948
rect 41767 6947 41803 6948
rect 41659 6939 41803 6947
rect 41659 6919 41667 6939
rect 41687 6919 41775 6939
rect 41795 6919 41803 6939
rect 41659 6913 41803 6919
rect 41869 6943 41907 6951
rect 41975 6947 42011 6948
rect 41869 6923 41878 6943
rect 41898 6923 41907 6943
rect 41869 6914 41907 6923
rect 41926 6940 42011 6947
rect 41926 6920 41933 6940
rect 41954 6939 42011 6940
rect 41954 6920 41983 6939
rect 41926 6919 41983 6920
rect 42003 6919 42011 6939
rect 41869 6913 41906 6914
rect 41926 6913 42011 6919
rect 42077 6943 42115 6951
rect 42188 6947 42224 6948
rect 42077 6923 42086 6943
rect 42106 6923 42115 6943
rect 42077 6914 42115 6923
rect 42139 6939 42224 6947
rect 42139 6919 42196 6939
rect 42216 6919 42224 6939
rect 42077 6913 42114 6914
rect 42139 6913 42224 6919
rect 42290 6943 42328 6951
rect 42290 6923 42299 6943
rect 42319 6923 42328 6943
rect 42290 6914 42328 6923
rect 42377 6917 42441 7101
rect 42597 6975 42662 7176
rect 42597 6957 42619 6975
rect 42637 6957 42662 6975
rect 42597 6938 42662 6957
rect 42290 6913 42327 6914
rect 41713 6892 41749 6913
rect 42139 6892 42170 6913
rect 42377 6908 42385 6917
rect 42374 6892 42385 6908
rect 41546 6888 41646 6892
rect 41546 6884 41608 6888
rect 41546 6858 41553 6884
rect 41579 6862 41608 6884
rect 41634 6862 41646 6888
rect 41579 6858 41646 6862
rect 41546 6855 41646 6858
rect 41714 6855 41749 6892
rect 41811 6889 42170 6892
rect 41811 6884 42033 6889
rect 41811 6860 41824 6884
rect 41848 6865 42033 6884
rect 42057 6865 42170 6889
rect 41848 6860 42170 6865
rect 41811 6856 42170 6860
rect 42237 6884 42385 6892
rect 42237 6864 42248 6884
rect 42268 6875 42385 6884
rect 42434 6908 42441 6917
rect 42434 6875 42442 6908
rect 42268 6864 42442 6875
rect 42237 6857 42442 6864
rect 42237 6856 42278 6857
rect 41713 6830 41749 6855
rect 41561 6803 41598 6804
rect 41657 6803 41694 6804
rect 41713 6803 41720 6830
rect 41237 6778 41245 6798
rect 41265 6778 41274 6798
rect 41091 6767 41122 6768
rect 41086 6699 41196 6712
rect 41237 6699 41274 6778
rect 41461 6794 41599 6803
rect 41461 6774 41570 6794
rect 41590 6774 41599 6794
rect 41461 6767 41599 6774
rect 41657 6800 41720 6803
rect 41741 6803 41749 6830
rect 41768 6803 41805 6804
rect 41741 6800 41805 6803
rect 41657 6794 41805 6800
rect 41657 6774 41666 6794
rect 41686 6774 41776 6794
rect 41796 6774 41805 6794
rect 41461 6765 41557 6767
rect 41657 6764 41805 6774
rect 41864 6794 41901 6804
rect 41976 6803 42013 6804
rect 41957 6801 42013 6803
rect 41864 6774 41872 6794
rect 41892 6774 41901 6794
rect 41713 6763 41749 6764
rect 41024 6697 41274 6699
rect 41024 6694 41125 6697
rect 41024 6675 41089 6694
rect 41086 6667 41089 6675
rect 41118 6667 41125 6694
rect 41153 6670 41163 6697
rect 41192 6675 41274 6697
rect 41192 6670 41196 6675
rect 41153 6667 41196 6670
rect 41086 6653 41196 6667
rect 40512 6635 40853 6636
rect 40437 6630 40853 6635
rect 41561 6632 41598 6633
rect 41864 6632 41901 6774
rect 41926 6794 42013 6801
rect 41926 6791 41984 6794
rect 41926 6771 41931 6791
rect 41952 6774 41984 6791
rect 42004 6774 42013 6794
rect 41952 6771 42013 6774
rect 41926 6764 42013 6771
rect 42072 6794 42109 6804
rect 42072 6774 42080 6794
rect 42100 6774 42109 6794
rect 41926 6763 41957 6764
rect 42072 6695 42109 6774
rect 42139 6803 42170 6856
rect 42374 6854 42442 6857
rect 42374 6812 42386 6854
rect 42435 6812 42442 6854
rect 42189 6803 42226 6804
rect 42139 6794 42226 6803
rect 42139 6774 42197 6794
rect 42217 6774 42226 6794
rect 42139 6764 42226 6774
rect 42285 6794 42322 6804
rect 42374 6799 42442 6812
rect 42597 6876 42662 6893
rect 42597 6858 42621 6876
rect 42639 6858 42662 6876
rect 42285 6774 42293 6794
rect 42313 6774 42322 6794
rect 42139 6763 42170 6764
rect 42134 6695 42244 6708
rect 42285 6695 42322 6774
rect 42597 6719 42662 6858
rect 42597 6713 42619 6719
rect 42072 6693 42322 6695
rect 42072 6690 42173 6693
rect 42072 6671 42137 6690
rect 42134 6663 42137 6671
rect 42166 6663 42173 6690
rect 42201 6666 42211 6693
rect 42240 6671 42322 6693
rect 42351 6701 42619 6713
rect 42637 6701 42662 6719
rect 42351 6678 42662 6701
rect 42351 6677 42406 6678
rect 42240 6666 42244 6671
rect 42201 6663 42244 6666
rect 42134 6649 42244 6663
rect 41560 6631 41901 6632
rect 40437 6610 40440 6630
rect 40460 6610 40853 6630
rect 41485 6630 41901 6631
rect 42351 6630 42394 6677
rect 41485 6626 42394 6630
rect 40804 6577 40849 6610
rect 41485 6606 41488 6626
rect 41508 6606 42394 6626
rect 41862 6601 42394 6606
rect 42602 6620 42661 6642
rect 42602 6602 42621 6620
rect 42639 6602 42661 6620
rect 41650 6577 41749 6579
rect 40804 6567 41749 6577
rect 40804 6541 41672 6567
rect 40805 6540 41672 6541
rect 41650 6529 41672 6540
rect 41697 6532 41716 6567
rect 41741 6532 41749 6567
rect 41697 6529 41749 6532
rect 42602 6531 42661 6602
rect 41650 6521 41749 6529
rect 41676 6520 41748 6521
rect 41330 6494 41397 6513
rect 41330 6473 41347 6494
rect 41328 6428 41347 6473
rect 41377 6473 41397 6494
rect 41377 6428 41398 6473
rect 41867 6470 41908 6472
rect 42139 6470 42243 6472
rect 42599 6470 42663 6531
rect 41328 6220 41398 6428
rect 41460 6435 42663 6470
rect 41460 6421 41488 6435
rect 41462 6290 41488 6421
rect 41867 6432 42663 6435
rect 40215 6128 40297 6148
rect 40215 6105 40243 6128
rect 40269 6105 40297 6128
rect 40215 6043 40297 6105
rect 40219 6008 40297 6043
rect 41320 6169 41400 6220
rect 41320 6143 41336 6169
rect 41376 6143 41400 6169
rect 41320 6124 41400 6143
rect 41320 6098 41339 6124
rect 41379 6098 41400 6124
rect 41320 6071 41400 6098
rect 41320 6045 41343 6071
rect 41383 6045 41400 6071
rect 41320 6034 41400 6045
rect 41462 6035 41489 6290
rect 41867 6282 41908 6432
rect 42139 6426 42243 6432
rect 42599 6429 42663 6432
rect 42334 6370 42455 6388
rect 42334 6368 42405 6370
rect 42334 6327 42349 6368
rect 42386 6329 42405 6368
rect 42442 6329 42455 6370
rect 42386 6327 42455 6329
rect 42334 6317 42455 6327
rect 41529 6175 41593 6187
rect 41869 6183 41906 6282
rect 42134 6272 42245 6285
rect 42134 6270 42176 6272
rect 42134 6250 42141 6270
rect 42160 6250 42176 6270
rect 42134 6242 42176 6250
rect 42204 6270 42245 6272
rect 42204 6250 42218 6270
rect 42237 6250 42245 6270
rect 42204 6242 42245 6250
rect 42134 6236 42245 6242
rect 42077 6214 42326 6236
rect 42077 6183 42114 6214
rect 42290 6212 42326 6214
rect 42290 6183 42327 6212
rect 41529 6174 41564 6175
rect 41506 6169 41564 6174
rect 41506 6149 41509 6169
rect 41529 6155 41564 6169
rect 41584 6155 41593 6175
rect 41529 6147 41593 6155
rect 41555 6146 41593 6147
rect 41556 6145 41593 6146
rect 41659 6179 41695 6180
rect 41767 6179 41803 6180
rect 41659 6171 41803 6179
rect 41659 6151 41667 6171
rect 41687 6151 41775 6171
rect 41795 6151 41803 6171
rect 41659 6145 41803 6151
rect 41869 6175 41907 6183
rect 41975 6179 42011 6180
rect 41869 6155 41878 6175
rect 41898 6155 41907 6175
rect 41869 6146 41907 6155
rect 41926 6172 42011 6179
rect 41926 6152 41933 6172
rect 41954 6171 42011 6172
rect 41954 6152 41983 6171
rect 41926 6151 41983 6152
rect 42003 6151 42011 6171
rect 41869 6145 41906 6146
rect 41926 6145 42011 6151
rect 42077 6175 42115 6183
rect 42188 6179 42224 6180
rect 42077 6155 42086 6175
rect 42106 6155 42115 6175
rect 42077 6146 42115 6155
rect 42139 6171 42224 6179
rect 42139 6151 42196 6171
rect 42216 6151 42224 6171
rect 42077 6145 42114 6146
rect 42139 6145 42224 6151
rect 42290 6175 42328 6183
rect 42290 6155 42299 6175
rect 42319 6155 42328 6175
rect 42383 6165 42448 6317
rect 42601 6291 42656 6429
rect 42290 6146 42328 6155
rect 42381 6158 42448 6165
rect 42290 6145 42327 6146
rect 41713 6124 41749 6145
rect 42139 6124 42170 6145
rect 42381 6137 42398 6158
rect 42434 6137 42448 6158
rect 42600 6178 42656 6291
rect 42600 6160 42619 6178
rect 42637 6160 42656 6178
rect 42600 6140 42656 6160
rect 42381 6124 42448 6137
rect 41546 6120 41646 6124
rect 41546 6116 41608 6120
rect 41546 6090 41553 6116
rect 41579 6094 41608 6116
rect 41634 6094 41646 6120
rect 41579 6090 41646 6094
rect 41546 6087 41646 6090
rect 41714 6087 41749 6124
rect 41811 6121 42170 6124
rect 41811 6116 42033 6121
rect 41811 6092 41824 6116
rect 41848 6097 42033 6116
rect 42057 6097 42170 6121
rect 41848 6092 42170 6097
rect 41811 6088 42170 6092
rect 42237 6118 42448 6124
rect 42237 6116 42398 6118
rect 42237 6096 42248 6116
rect 42268 6096 42398 6116
rect 42237 6089 42398 6096
rect 42237 6088 42278 6089
rect 41713 6062 41749 6087
rect 41561 6035 41598 6036
rect 41657 6035 41694 6036
rect 41713 6035 41720 6062
rect 41461 6026 41599 6035
rect 40219 5492 40281 6008
rect 41461 6006 41570 6026
rect 41590 6006 41599 6026
rect 41461 5999 41599 6006
rect 41657 6032 41720 6035
rect 41741 6035 41749 6062
rect 41768 6035 41805 6036
rect 41741 6032 41805 6035
rect 41657 6026 41805 6032
rect 41657 6006 41666 6026
rect 41686 6006 41776 6026
rect 41796 6006 41805 6026
rect 41461 5997 41557 5999
rect 41657 5996 41805 6006
rect 41864 6026 41901 6036
rect 41976 6035 42013 6036
rect 41957 6033 42013 6035
rect 41864 6006 41872 6026
rect 41892 6006 41901 6026
rect 41713 5995 41749 5996
rect 41561 5864 41598 5865
rect 41864 5864 41901 6006
rect 41926 6026 42013 6033
rect 41926 6023 41984 6026
rect 41926 6003 41931 6023
rect 41952 6006 41984 6023
rect 42004 6006 42013 6026
rect 41952 6003 42013 6006
rect 41926 5996 42013 6003
rect 42072 6026 42109 6036
rect 42072 6006 42080 6026
rect 42100 6006 42109 6026
rect 41926 5995 41957 5996
rect 42072 5927 42109 6006
rect 42139 6035 42170 6088
rect 42383 6081 42398 6089
rect 42438 6081 42448 6118
rect 42383 6072 42448 6081
rect 42596 6079 42661 6100
rect 42596 6061 42621 6079
rect 42639 6061 42661 6079
rect 42189 6035 42226 6036
rect 42139 6026 42226 6035
rect 42139 6006 42197 6026
rect 42217 6006 42226 6026
rect 42139 5996 42226 6006
rect 42285 6026 42322 6036
rect 42285 6006 42293 6026
rect 42313 6006 42322 6026
rect 42139 5995 42170 5996
rect 42134 5927 42244 5940
rect 42285 5927 42322 6006
rect 42596 5985 42661 6061
rect 42072 5925 42322 5927
rect 42072 5922 42173 5925
rect 42072 5903 42137 5922
rect 42134 5895 42137 5903
rect 42166 5895 42173 5922
rect 42201 5898 42211 5925
rect 42240 5903 42322 5925
rect 42345 5950 42662 5985
rect 42240 5898 42244 5903
rect 42201 5895 42244 5898
rect 42134 5881 42244 5895
rect 41560 5863 41901 5864
rect 41485 5861 41901 5863
rect 42345 5861 42385 5950
rect 42596 5923 42661 5950
rect 42596 5905 42619 5923
rect 42637 5905 42661 5923
rect 42596 5885 42661 5905
rect 41482 5858 42385 5861
rect 41482 5838 41488 5858
rect 41508 5838 42385 5858
rect 41482 5834 42385 5838
rect 42345 5831 42385 5834
rect 42597 5824 42662 5845
rect 40815 5816 41476 5817
rect 40815 5809 41749 5816
rect 40815 5808 41721 5809
rect 40815 5788 41666 5808
rect 41698 5789 41721 5808
rect 41746 5789 41749 5809
rect 41698 5788 41749 5789
rect 40815 5781 41749 5788
rect 40414 5739 40582 5740
rect 40817 5739 40856 5781
rect 41645 5779 41749 5781
rect 41714 5777 41749 5779
rect 42597 5806 42621 5824
rect 42639 5806 42662 5824
rect 42597 5759 42662 5806
rect 40414 5713 40858 5739
rect 40414 5711 40582 5713
rect 40216 5408 40285 5492
rect 40214 4929 40285 5408
rect 40414 5360 40441 5711
rect 40817 5707 40858 5713
rect 40481 5500 40545 5512
rect 40821 5508 40858 5707
rect 41320 5734 41392 5751
rect 41320 5695 41328 5734
rect 41373 5695 41392 5734
rect 41086 5597 41197 5612
rect 41086 5595 41128 5597
rect 41086 5575 41093 5595
rect 41112 5575 41128 5595
rect 41086 5567 41128 5575
rect 41156 5595 41197 5597
rect 41156 5575 41170 5595
rect 41189 5575 41197 5595
rect 41156 5567 41197 5575
rect 41086 5561 41197 5567
rect 41029 5539 41278 5561
rect 41029 5508 41066 5539
rect 41242 5537 41278 5539
rect 41242 5508 41279 5537
rect 40481 5499 40516 5500
rect 40458 5494 40516 5499
rect 40458 5474 40461 5494
rect 40481 5480 40516 5494
rect 40536 5480 40545 5500
rect 40481 5472 40545 5480
rect 40507 5471 40545 5472
rect 40508 5470 40545 5471
rect 40611 5504 40647 5505
rect 40719 5504 40755 5505
rect 40611 5496 40755 5504
rect 40611 5476 40619 5496
rect 40639 5476 40727 5496
rect 40747 5476 40755 5496
rect 40611 5470 40755 5476
rect 40821 5500 40859 5508
rect 40927 5504 40963 5505
rect 40821 5480 40830 5500
rect 40850 5480 40859 5500
rect 40821 5471 40859 5480
rect 40878 5497 40963 5504
rect 40878 5477 40885 5497
rect 40906 5496 40963 5497
rect 40906 5477 40935 5496
rect 40878 5476 40935 5477
rect 40955 5476 40963 5496
rect 40821 5470 40858 5471
rect 40878 5470 40963 5476
rect 41029 5500 41067 5508
rect 41140 5504 41176 5505
rect 41029 5480 41038 5500
rect 41058 5480 41067 5500
rect 41029 5471 41067 5480
rect 41091 5496 41176 5504
rect 41091 5476 41148 5496
rect 41168 5476 41176 5496
rect 41029 5470 41066 5471
rect 41091 5470 41176 5476
rect 41242 5500 41280 5508
rect 41242 5480 41251 5500
rect 41271 5480 41280 5500
rect 41242 5471 41280 5480
rect 41320 5485 41392 5695
rect 41462 5729 42662 5759
rect 41462 5728 41906 5729
rect 41462 5726 41630 5728
rect 41320 5471 41403 5485
rect 41242 5470 41279 5471
rect 40665 5449 40701 5470
rect 41091 5449 41122 5470
rect 41320 5449 41337 5471
rect 40498 5445 40598 5449
rect 40498 5441 40560 5445
rect 40498 5415 40505 5441
rect 40531 5419 40560 5441
rect 40586 5419 40598 5445
rect 40531 5415 40598 5419
rect 40498 5412 40598 5415
rect 40666 5412 40701 5449
rect 40763 5446 41122 5449
rect 40763 5441 40985 5446
rect 40763 5417 40776 5441
rect 40800 5422 40985 5441
rect 41009 5422 41122 5446
rect 40800 5417 41122 5422
rect 40763 5413 41122 5417
rect 41189 5441 41337 5449
rect 41189 5421 41200 5441
rect 41220 5438 41337 5441
rect 41390 5438 41403 5471
rect 41220 5421 41403 5438
rect 41189 5414 41403 5421
rect 41189 5413 41230 5414
rect 41320 5413 41403 5414
rect 40665 5387 40701 5412
rect 40513 5360 40550 5361
rect 40609 5360 40646 5361
rect 40665 5360 40672 5387
rect 40413 5351 40551 5360
rect 40413 5331 40522 5351
rect 40542 5331 40551 5351
rect 40413 5324 40551 5331
rect 40609 5357 40672 5360
rect 40693 5360 40701 5387
rect 40720 5360 40757 5361
rect 40693 5357 40757 5360
rect 40609 5351 40757 5357
rect 40609 5331 40618 5351
rect 40638 5331 40728 5351
rect 40748 5331 40757 5351
rect 40413 5322 40509 5324
rect 40609 5321 40757 5331
rect 40816 5351 40853 5361
rect 40928 5360 40965 5361
rect 40909 5358 40965 5360
rect 40816 5331 40824 5351
rect 40844 5331 40853 5351
rect 40665 5320 40701 5321
rect 40513 5189 40550 5190
rect 40816 5189 40853 5331
rect 40878 5351 40965 5358
rect 40878 5348 40936 5351
rect 40878 5328 40883 5348
rect 40904 5331 40936 5348
rect 40956 5331 40965 5351
rect 40904 5328 40965 5331
rect 40878 5321 40965 5328
rect 41024 5351 41061 5361
rect 41024 5331 41032 5351
rect 41052 5331 41061 5351
rect 40878 5320 40909 5321
rect 41024 5252 41061 5331
rect 41091 5360 41122 5413
rect 41328 5380 41342 5413
rect 41395 5380 41403 5413
rect 41328 5374 41403 5380
rect 41328 5369 41398 5374
rect 41141 5360 41178 5361
rect 41091 5351 41178 5360
rect 41091 5331 41149 5351
rect 41169 5331 41178 5351
rect 41091 5321 41178 5331
rect 41237 5351 41274 5361
rect 41462 5356 41489 5726
rect 41529 5496 41593 5508
rect 41869 5504 41906 5728
rect 42377 5709 42441 5711
rect 42373 5697 42441 5709
rect 42373 5664 42384 5697
rect 42424 5664 42441 5697
rect 42373 5654 42441 5664
rect 42134 5593 42245 5608
rect 42134 5591 42176 5593
rect 42134 5571 42141 5591
rect 42160 5571 42176 5591
rect 42134 5563 42176 5571
rect 42204 5591 42245 5593
rect 42204 5571 42218 5591
rect 42237 5571 42245 5591
rect 42204 5563 42245 5571
rect 42134 5557 42245 5563
rect 42077 5535 42326 5557
rect 42077 5504 42114 5535
rect 42290 5533 42326 5535
rect 42290 5504 42327 5533
rect 41529 5495 41564 5496
rect 41506 5490 41564 5495
rect 41506 5470 41509 5490
rect 41529 5476 41564 5490
rect 41584 5476 41593 5496
rect 41529 5468 41593 5476
rect 41555 5467 41593 5468
rect 41556 5466 41593 5467
rect 41659 5500 41695 5501
rect 41767 5500 41803 5501
rect 41659 5492 41803 5500
rect 41659 5472 41667 5492
rect 41687 5472 41775 5492
rect 41795 5472 41803 5492
rect 41659 5466 41803 5472
rect 41869 5496 41907 5504
rect 41975 5500 42011 5501
rect 41869 5476 41878 5496
rect 41898 5476 41907 5496
rect 41869 5467 41907 5476
rect 41926 5493 42011 5500
rect 41926 5473 41933 5493
rect 41954 5492 42011 5493
rect 41954 5473 41983 5492
rect 41926 5472 41983 5473
rect 42003 5472 42011 5492
rect 41869 5466 41906 5467
rect 41926 5466 42011 5472
rect 42077 5496 42115 5504
rect 42188 5500 42224 5501
rect 42077 5476 42086 5496
rect 42106 5476 42115 5496
rect 42077 5467 42115 5476
rect 42139 5492 42224 5500
rect 42139 5472 42196 5492
rect 42216 5472 42224 5492
rect 42077 5466 42114 5467
rect 42139 5466 42224 5472
rect 42290 5496 42328 5504
rect 42290 5476 42299 5496
rect 42319 5476 42328 5496
rect 42290 5467 42328 5476
rect 42377 5470 42441 5654
rect 42597 5528 42662 5729
rect 42597 5510 42619 5528
rect 42637 5510 42662 5528
rect 42597 5491 42662 5510
rect 42290 5466 42327 5467
rect 41713 5445 41749 5466
rect 42139 5445 42170 5466
rect 42377 5461 42385 5470
rect 42374 5445 42385 5461
rect 41546 5441 41646 5445
rect 41546 5437 41608 5441
rect 41546 5411 41553 5437
rect 41579 5415 41608 5437
rect 41634 5415 41646 5441
rect 41579 5411 41646 5415
rect 41546 5408 41646 5411
rect 41714 5408 41749 5445
rect 41811 5442 42170 5445
rect 41811 5437 42033 5442
rect 41811 5413 41824 5437
rect 41848 5418 42033 5437
rect 42057 5418 42170 5442
rect 41848 5413 42170 5418
rect 41811 5409 42170 5413
rect 42237 5437 42385 5445
rect 42237 5417 42248 5437
rect 42268 5428 42385 5437
rect 42434 5461 42441 5470
rect 42434 5428 42442 5461
rect 42268 5417 42442 5428
rect 42237 5410 42442 5417
rect 42237 5409 42278 5410
rect 41713 5383 41749 5408
rect 41561 5356 41598 5357
rect 41657 5356 41694 5357
rect 41713 5356 41720 5383
rect 41237 5331 41245 5351
rect 41265 5331 41274 5351
rect 41091 5320 41122 5321
rect 41086 5252 41196 5265
rect 41237 5252 41274 5331
rect 41461 5347 41599 5356
rect 41461 5327 41570 5347
rect 41590 5327 41599 5347
rect 41461 5320 41599 5327
rect 41657 5353 41720 5356
rect 41741 5356 41749 5383
rect 41768 5356 41805 5357
rect 41741 5353 41805 5356
rect 41657 5347 41805 5353
rect 41657 5327 41666 5347
rect 41686 5327 41776 5347
rect 41796 5327 41805 5347
rect 41461 5318 41557 5320
rect 41657 5317 41805 5327
rect 41864 5347 41901 5357
rect 41976 5356 42013 5357
rect 41957 5354 42013 5356
rect 41864 5327 41872 5347
rect 41892 5327 41901 5347
rect 41713 5316 41749 5317
rect 41024 5250 41274 5252
rect 41024 5247 41125 5250
rect 41024 5228 41089 5247
rect 41086 5220 41089 5228
rect 41118 5220 41125 5247
rect 41153 5223 41163 5250
rect 41192 5228 41274 5250
rect 41192 5223 41196 5228
rect 41153 5220 41196 5223
rect 41086 5206 41196 5220
rect 40512 5188 40853 5189
rect 40437 5183 40853 5188
rect 41561 5185 41598 5186
rect 41864 5185 41901 5327
rect 41926 5347 42013 5354
rect 41926 5344 41984 5347
rect 41926 5324 41931 5344
rect 41952 5327 41984 5344
rect 42004 5327 42013 5347
rect 41952 5324 42013 5327
rect 41926 5317 42013 5324
rect 42072 5347 42109 5357
rect 42072 5327 42080 5347
rect 42100 5327 42109 5347
rect 41926 5316 41957 5317
rect 42072 5248 42109 5327
rect 42139 5356 42170 5409
rect 42374 5407 42442 5410
rect 42374 5365 42386 5407
rect 42435 5365 42442 5407
rect 42189 5356 42226 5357
rect 42139 5347 42226 5356
rect 42139 5327 42197 5347
rect 42217 5327 42226 5347
rect 42139 5317 42226 5327
rect 42285 5347 42322 5357
rect 42374 5352 42442 5365
rect 42597 5429 42662 5446
rect 42597 5411 42621 5429
rect 42639 5411 42662 5429
rect 42285 5327 42293 5347
rect 42313 5327 42322 5347
rect 42139 5316 42170 5317
rect 42134 5248 42244 5261
rect 42285 5248 42322 5327
rect 42597 5272 42662 5411
rect 42597 5266 42619 5272
rect 42072 5246 42322 5248
rect 42072 5243 42173 5246
rect 42072 5224 42137 5243
rect 42134 5216 42137 5224
rect 42166 5216 42173 5243
rect 42201 5219 42211 5246
rect 42240 5224 42322 5246
rect 42351 5254 42619 5266
rect 42637 5254 42662 5272
rect 42351 5231 42662 5254
rect 42351 5230 42406 5231
rect 42240 5219 42244 5224
rect 42201 5216 42244 5219
rect 42134 5202 42244 5216
rect 41560 5184 41901 5185
rect 40437 5163 40440 5183
rect 40460 5163 40853 5183
rect 41485 5183 41901 5184
rect 42351 5183 42394 5230
rect 41485 5179 42394 5183
rect 40804 5130 40849 5163
rect 41485 5159 41488 5179
rect 41508 5159 42394 5179
rect 41862 5154 42394 5159
rect 42602 5173 42661 5195
rect 42602 5155 42621 5173
rect 42639 5155 42661 5173
rect 41650 5130 41749 5132
rect 40804 5120 41749 5130
rect 40804 5094 41672 5120
rect 40805 5093 41672 5094
rect 41650 5082 41672 5093
rect 41697 5085 41716 5120
rect 41741 5085 41749 5120
rect 41697 5082 41749 5085
rect 41650 5074 41749 5082
rect 41676 5073 41748 5074
rect 42602 5025 42661 5155
rect 41324 4995 41400 5019
rect 41324 4929 41336 4995
rect 41390 4929 41400 4995
rect 41868 4950 41909 4952
rect 42140 4950 42244 4952
rect 42602 4950 42663 5025
rect 40214 4879 40286 4929
rect 39783 4607 40119 4611
rect 39009 4603 39109 4607
rect 39009 4599 39071 4603
rect 39009 4573 39016 4599
rect 39042 4577 39071 4599
rect 39097 4577 39109 4603
rect 39042 4573 39109 4577
rect 39009 4570 39109 4573
rect 39177 4570 39212 4607
rect 39274 4604 39633 4607
rect 39274 4599 39496 4604
rect 39274 4575 39287 4599
rect 39311 4580 39496 4599
rect 39520 4580 39633 4604
rect 39311 4575 39633 4580
rect 39274 4571 39633 4575
rect 39700 4599 40119 4607
rect 39700 4579 39711 4599
rect 39731 4579 40119 4599
rect 39700 4572 40119 4579
rect 39700 4571 39741 4572
rect 39783 4571 40119 4572
rect 39176 4545 39212 4570
rect 39024 4518 39061 4519
rect 39120 4518 39157 4519
rect 39176 4518 39183 4545
rect 38924 4509 39062 4518
rect 38924 4489 39033 4509
rect 39053 4489 39062 4509
rect 38924 4482 39062 4489
rect 39120 4515 39183 4518
rect 39204 4518 39212 4545
rect 39231 4518 39268 4519
rect 39204 4515 39268 4518
rect 39120 4509 39268 4515
rect 39120 4489 39129 4509
rect 39149 4489 39239 4509
rect 39259 4489 39268 4509
rect 38924 4480 39020 4482
rect 39120 4479 39268 4489
rect 39327 4509 39364 4519
rect 39439 4518 39476 4519
rect 39420 4516 39476 4518
rect 39327 4489 39335 4509
rect 39355 4489 39364 4509
rect 39176 4478 39212 4479
rect 39024 4347 39061 4348
rect 39327 4347 39364 4489
rect 39389 4509 39476 4516
rect 39389 4506 39447 4509
rect 39389 4486 39394 4506
rect 39415 4489 39447 4506
rect 39467 4489 39476 4509
rect 39415 4486 39476 4489
rect 39389 4479 39476 4486
rect 39535 4509 39572 4519
rect 39535 4489 39543 4509
rect 39563 4489 39572 4509
rect 39389 4478 39420 4479
rect 39535 4410 39572 4489
rect 39602 4518 39633 4571
rect 40027 4535 40119 4571
rect 39652 4518 39689 4519
rect 39602 4509 39689 4518
rect 39602 4489 39660 4509
rect 39680 4489 39689 4509
rect 39602 4479 39689 4489
rect 39748 4509 39785 4519
rect 39748 4489 39756 4509
rect 39776 4489 39785 4509
rect 39602 4478 39633 4479
rect 39597 4410 39707 4423
rect 39748 4410 39785 4489
rect 39535 4408 39785 4410
rect 39535 4405 39636 4408
rect 39535 4386 39600 4405
rect 39597 4378 39600 4386
rect 39629 4378 39636 4405
rect 39664 4381 39674 4408
rect 39703 4386 39785 4408
rect 39703 4381 39707 4386
rect 39664 4378 39707 4381
rect 39597 4364 39707 4378
rect 39023 4346 39364 4347
rect 38948 4341 39364 4346
rect 38948 4321 38951 4341
rect 38971 4321 39364 4341
rect 39108 4277 39213 4280
rect 39107 4254 39213 4277
rect 38227 4252 38728 4254
rect 38869 4252 39218 4254
rect 36341 4231 36378 4252
rect 36341 4194 36352 4231
rect 36369 4194 36378 4231
rect 38227 4246 39218 4252
rect 38227 4241 39179 4246
rect 38227 4220 39138 4241
rect 39158 4225 39179 4241
rect 39199 4225 39218 4246
rect 39158 4220 39218 4225
rect 38227 4195 39218 4220
rect 38703 4194 38885 4195
rect 36341 4184 36378 4194
rect 36187 4141 36581 4161
rect 36601 4141 36604 4161
rect 36188 4136 36604 4141
rect 36188 4135 36529 4136
rect 35845 4104 35955 4118
rect 35845 4101 35888 4104
rect 35845 4096 35849 4101
rect 35767 4074 35849 4096
rect 35878 4074 35888 4101
rect 35916 4077 35923 4104
rect 35952 4096 35955 4104
rect 35952 4077 36017 4096
rect 35916 4074 36017 4077
rect 35767 4072 36017 4074
rect 35767 3993 35804 4072
rect 35845 4059 35955 4072
rect 35919 4003 35950 4004
rect 35767 3973 35776 3993
rect 35796 3973 35804 3993
rect 35767 3963 35804 3973
rect 35863 3993 35950 4003
rect 35863 3973 35872 3993
rect 35892 3973 35950 3993
rect 35863 3964 35950 3973
rect 35863 3963 35900 3964
rect 35919 3911 35950 3964
rect 35980 3993 36017 4072
rect 36132 4003 36163 4004
rect 35980 3973 35989 3993
rect 36009 3973 36017 3993
rect 35980 3963 36017 3973
rect 36076 3996 36163 4003
rect 36076 3993 36137 3996
rect 36076 3973 36085 3993
rect 36105 3976 36137 3993
rect 36158 3976 36163 3996
rect 36105 3973 36163 3976
rect 36076 3966 36163 3973
rect 36188 3993 36225 4135
rect 36491 4134 36528 4135
rect 36340 4003 36376 4004
rect 36188 3973 36197 3993
rect 36217 3973 36225 3993
rect 36076 3964 36132 3966
rect 36076 3963 36113 3964
rect 36188 3963 36225 3973
rect 36284 3993 36432 4003
rect 36532 4000 36628 4002
rect 36284 3973 36293 3993
rect 36313 3973 36403 3993
rect 36423 3973 36432 3993
rect 36284 3967 36432 3973
rect 36284 3964 36348 3967
rect 36284 3963 36321 3964
rect 36340 3937 36348 3964
rect 36369 3964 36432 3967
rect 36490 3993 36628 4000
rect 36490 3973 36499 3993
rect 36519 3973 36628 3993
rect 36490 3964 36628 3973
rect 39257 3965 39288 4321
rect 36369 3937 36376 3964
rect 36395 3963 36432 3964
rect 36491 3963 36528 3964
rect 36340 3912 36376 3937
rect 35811 3910 35852 3911
rect 35731 3905 35852 3910
rect 35682 3903 35852 3905
rect 35682 3892 35821 3903
rect 35682 3869 35705 3892
rect 35731 3883 35821 3892
rect 35841 3883 35852 3903
rect 35731 3875 35852 3883
rect 35919 3907 36278 3911
rect 35919 3902 36241 3907
rect 35919 3878 36032 3902
rect 36056 3883 36241 3902
rect 36265 3883 36278 3907
rect 36056 3878 36278 3883
rect 35919 3875 36278 3878
rect 36340 3875 36375 3912
rect 36443 3909 36543 3912
rect 36443 3905 36510 3909
rect 36443 3879 36455 3905
rect 36481 3883 36510 3905
rect 36536 3883 36543 3909
rect 36481 3879 36543 3883
rect 36443 3875 36543 3879
rect 35731 3869 35739 3875
rect 35682 3861 35739 3869
rect 35919 3854 35950 3875
rect 36340 3854 36376 3875
rect 35762 3853 35799 3854
rect 35761 3844 35799 3853
rect 35761 3824 35770 3844
rect 35790 3824 35799 3844
rect 35761 3816 35799 3824
rect 35865 3848 35950 3854
rect 35975 3853 36012 3854
rect 35865 3828 35873 3848
rect 35893 3828 35950 3848
rect 35865 3820 35950 3828
rect 35974 3844 36012 3853
rect 35974 3824 35983 3844
rect 36003 3824 36012 3844
rect 35865 3819 35901 3820
rect 35974 3816 36012 3824
rect 36078 3848 36163 3854
rect 36183 3853 36220 3854
rect 36078 3828 36086 3848
rect 36106 3847 36163 3848
rect 36106 3828 36135 3847
rect 36078 3827 36135 3828
rect 36156 3827 36163 3847
rect 36078 3820 36163 3827
rect 36182 3844 36220 3853
rect 36182 3824 36191 3844
rect 36211 3824 36220 3844
rect 36078 3819 36114 3820
rect 36182 3816 36220 3824
rect 36286 3848 36430 3854
rect 36286 3828 36294 3848
rect 36314 3828 36402 3848
rect 36422 3828 36430 3848
rect 36286 3820 36430 3828
rect 36286 3819 36322 3820
rect 36394 3819 36430 3820
rect 36496 3853 36533 3854
rect 36496 3852 36534 3853
rect 36496 3844 36560 3852
rect 36496 3824 36505 3844
rect 36525 3830 36560 3844
rect 36580 3830 36583 3850
rect 36525 3825 36583 3830
rect 36525 3824 36560 3825
rect 35762 3787 35799 3816
rect 35763 3785 35799 3787
rect 35975 3785 36012 3816
rect 35763 3763 36012 3785
rect 35844 3757 35955 3763
rect 35844 3749 35885 3757
rect 35844 3729 35852 3749
rect 35871 3729 35885 3749
rect 35844 3727 35885 3729
rect 35913 3749 35955 3757
rect 35913 3729 35929 3749
rect 35948 3729 35955 3749
rect 35913 3727 35955 3729
rect 35844 3712 35955 3727
rect 36183 3701 36220 3816
rect 36496 3812 36560 3824
rect 36176 3695 36223 3701
rect 36600 3697 36627 3964
rect 39175 3936 39288 3965
rect 36459 3695 36627 3697
rect 36176 3669 36627 3695
rect 36176 3534 36223 3669
rect 36459 3668 36627 3669
rect 39176 3627 39212 3936
rect 40036 3822 40117 4535
rect 40216 3970 40286 4879
rect 41324 4909 41400 4929
rect 41324 4872 41341 4909
rect 41385 4872 41400 4909
rect 41461 4915 42663 4950
rect 41461 4901 41489 4915
rect 41324 4856 41400 4872
rect 41329 4700 41399 4856
rect 41463 4770 41489 4901
rect 41868 4912 42663 4915
rect 41321 4649 41401 4700
rect 41321 4623 41337 4649
rect 41377 4623 41401 4649
rect 41321 4604 41401 4623
rect 41321 4578 41340 4604
rect 41380 4578 41401 4604
rect 41321 4551 41401 4578
rect 41321 4525 41344 4551
rect 41384 4525 41401 4551
rect 41321 4514 41401 4525
rect 41463 4515 41490 4770
rect 41868 4762 41909 4912
rect 42602 4900 42663 4912
rect 42335 4850 42456 4868
rect 42335 4848 42406 4850
rect 42335 4807 42350 4848
rect 42387 4809 42406 4848
rect 42443 4809 42456 4850
rect 42387 4807 42456 4809
rect 42335 4797 42456 4807
rect 42140 4767 42244 4776
rect 41530 4655 41594 4667
rect 41870 4663 41907 4762
rect 42135 4752 42246 4767
rect 42135 4750 42177 4752
rect 42135 4730 42142 4750
rect 42161 4730 42177 4750
rect 42135 4722 42177 4730
rect 42205 4750 42246 4752
rect 42205 4730 42219 4750
rect 42238 4730 42246 4750
rect 42205 4722 42246 4730
rect 42135 4716 42246 4722
rect 42078 4694 42327 4716
rect 42078 4663 42115 4694
rect 42291 4692 42327 4694
rect 42291 4663 42328 4692
rect 41530 4654 41565 4655
rect 41507 4649 41565 4654
rect 41507 4629 41510 4649
rect 41530 4635 41565 4649
rect 41585 4635 41594 4655
rect 41530 4627 41594 4635
rect 41556 4626 41594 4627
rect 41557 4625 41594 4626
rect 41660 4659 41696 4660
rect 41768 4659 41804 4660
rect 41660 4651 41804 4659
rect 41660 4631 41668 4651
rect 41688 4631 41776 4651
rect 41796 4631 41804 4651
rect 41660 4625 41804 4631
rect 41870 4655 41908 4663
rect 41976 4659 42012 4660
rect 41870 4635 41879 4655
rect 41899 4635 41908 4655
rect 41870 4626 41908 4635
rect 41927 4652 42012 4659
rect 41927 4632 41934 4652
rect 41955 4651 42012 4652
rect 41955 4632 41984 4651
rect 41927 4631 41984 4632
rect 42004 4631 42012 4651
rect 41870 4625 41907 4626
rect 41927 4625 42012 4631
rect 42078 4655 42116 4663
rect 42189 4659 42225 4660
rect 42078 4635 42087 4655
rect 42107 4635 42116 4655
rect 42078 4626 42116 4635
rect 42140 4651 42225 4659
rect 42140 4631 42197 4651
rect 42217 4631 42225 4651
rect 42078 4625 42115 4626
rect 42140 4625 42225 4631
rect 42291 4655 42329 4663
rect 42291 4635 42300 4655
rect 42320 4635 42329 4655
rect 42384 4645 42449 4797
rect 42602 4771 42657 4900
rect 42291 4626 42329 4635
rect 42382 4638 42449 4645
rect 42291 4625 42328 4626
rect 41714 4604 41750 4625
rect 42140 4604 42171 4625
rect 42382 4617 42399 4638
rect 42435 4617 42449 4638
rect 42601 4658 42657 4771
rect 42601 4640 42620 4658
rect 42638 4640 42657 4658
rect 42601 4620 42657 4640
rect 42382 4604 42449 4617
rect 41547 4600 41647 4604
rect 41547 4596 41609 4600
rect 41547 4570 41554 4596
rect 41580 4574 41609 4596
rect 41635 4574 41647 4600
rect 41580 4570 41647 4574
rect 41547 4567 41647 4570
rect 41715 4567 41750 4604
rect 41812 4601 42171 4604
rect 41812 4596 42034 4601
rect 41812 4572 41825 4596
rect 41849 4577 42034 4596
rect 42058 4577 42171 4601
rect 41849 4572 42171 4577
rect 41812 4568 42171 4572
rect 42238 4598 42449 4604
rect 42238 4596 42399 4598
rect 42238 4576 42249 4596
rect 42269 4576 42399 4596
rect 42238 4569 42399 4576
rect 42238 4568 42279 4569
rect 41714 4542 41750 4567
rect 41562 4515 41599 4516
rect 41658 4515 41695 4516
rect 41714 4515 41721 4542
rect 41462 4506 41600 4515
rect 41462 4486 41571 4506
rect 41591 4486 41600 4506
rect 41462 4479 41600 4486
rect 41658 4512 41721 4515
rect 41742 4515 41750 4542
rect 41769 4515 41806 4516
rect 41742 4512 41806 4515
rect 41658 4506 41806 4512
rect 41658 4486 41667 4506
rect 41687 4486 41777 4506
rect 41797 4486 41806 4506
rect 41462 4477 41558 4479
rect 41658 4476 41806 4486
rect 41865 4506 41902 4516
rect 41977 4515 42014 4516
rect 41958 4513 42014 4515
rect 41865 4486 41873 4506
rect 41893 4486 41902 4506
rect 41714 4475 41750 4476
rect 41562 4344 41599 4345
rect 41865 4344 41902 4486
rect 41927 4506 42014 4513
rect 41927 4503 41985 4506
rect 41927 4483 41932 4503
rect 41953 4486 41985 4503
rect 42005 4486 42014 4506
rect 41953 4483 42014 4486
rect 41927 4476 42014 4483
rect 42073 4506 42110 4516
rect 42073 4486 42081 4506
rect 42101 4486 42110 4506
rect 41927 4475 41958 4476
rect 42073 4407 42110 4486
rect 42140 4515 42171 4568
rect 42384 4561 42399 4569
rect 42439 4561 42449 4598
rect 42384 4552 42449 4561
rect 42597 4559 42662 4580
rect 42597 4541 42622 4559
rect 42640 4541 42662 4559
rect 42190 4515 42227 4516
rect 42140 4506 42227 4515
rect 42140 4486 42198 4506
rect 42218 4486 42227 4506
rect 42140 4476 42227 4486
rect 42286 4506 42323 4516
rect 42286 4486 42294 4506
rect 42314 4486 42323 4506
rect 42140 4475 42171 4476
rect 42135 4407 42245 4420
rect 42286 4407 42323 4486
rect 42597 4465 42662 4541
rect 42073 4405 42323 4407
rect 42073 4402 42174 4405
rect 42073 4383 42138 4402
rect 42135 4375 42138 4383
rect 42167 4375 42174 4402
rect 42202 4378 42212 4405
rect 42241 4383 42323 4405
rect 42346 4430 42663 4465
rect 42241 4378 42245 4383
rect 42202 4375 42245 4378
rect 42135 4361 42245 4375
rect 41561 4343 41902 4344
rect 41486 4341 41902 4343
rect 42346 4341 42386 4430
rect 42597 4403 42662 4430
rect 42597 4385 42620 4403
rect 42638 4385 42662 4403
rect 42597 4365 42662 4385
rect 41483 4338 42386 4341
rect 41483 4318 41489 4338
rect 41509 4318 42386 4338
rect 41483 4314 42386 4318
rect 42346 4311 42386 4314
rect 42598 4304 42663 4325
rect 40816 4296 41477 4297
rect 40816 4289 41750 4296
rect 40816 4288 41722 4289
rect 40816 4268 41667 4288
rect 41699 4269 41722 4288
rect 41747 4269 41750 4289
rect 41699 4268 41750 4269
rect 40816 4261 41750 4268
rect 40415 4219 40583 4220
rect 40818 4219 40857 4261
rect 41646 4259 41750 4261
rect 41715 4257 41750 4259
rect 42598 4286 42622 4304
rect 42640 4286 42663 4304
rect 42598 4239 42663 4286
rect 40415 4193 40859 4219
rect 40415 4191 40583 4193
rect 39176 3604 39180 3627
rect 39204 3604 39212 3627
rect 39376 3605 39475 3609
rect 39176 3583 39212 3604
rect 39176 3560 39180 3583
rect 39204 3560 39212 3583
rect 39176 3556 39212 3560
rect 39372 3599 39475 3605
rect 39372 3561 39398 3599
rect 39423 3564 39442 3599
rect 39467 3564 39475 3599
rect 39423 3561 39475 3564
rect 39372 3553 39475 3561
rect 39372 3552 39474 3553
rect 36174 3485 36233 3534
rect 36174 3457 36192 3485
rect 36220 3457 36233 3485
rect 36174 3447 36233 3457
rect 38968 3474 39136 3475
rect 39372 3474 39419 3552
rect 38968 3448 39419 3474
rect 38968 3446 39136 3448
rect 38968 3073 38995 3446
rect 39165 3398 39251 3407
rect 39165 3380 39184 3398
rect 39236 3380 39251 3398
rect 39165 3376 39251 3380
rect 39035 3213 39099 3225
rect 39035 3212 39070 3213
rect 39012 3207 39070 3212
rect 39012 3187 39015 3207
rect 39035 3193 39070 3207
rect 39090 3193 39099 3213
rect 39035 3185 39099 3193
rect 39061 3184 39099 3185
rect 39062 3183 39099 3184
rect 39165 3217 39201 3218
rect 39221 3217 39251 3376
rect 39372 3336 39419 3448
rect 39375 3221 39412 3336
rect 39640 3310 39751 3325
rect 39640 3308 39682 3310
rect 39640 3288 39647 3308
rect 39666 3288 39682 3308
rect 39640 3280 39682 3288
rect 39710 3308 39751 3310
rect 39710 3288 39724 3308
rect 39743 3288 39751 3308
rect 39710 3280 39751 3288
rect 39640 3274 39751 3280
rect 39583 3252 39832 3274
rect 39583 3221 39620 3252
rect 39796 3250 39832 3252
rect 39796 3221 39833 3250
rect 40037 3237 40116 3822
rect 40213 3370 40292 3970
rect 40415 3840 40442 4191
rect 40818 4187 40859 4193
rect 40482 3980 40546 3992
rect 40822 3988 40859 4187
rect 41321 4214 41393 4231
rect 41321 4175 41329 4214
rect 41374 4175 41393 4214
rect 41087 4077 41198 4092
rect 41087 4075 41129 4077
rect 41087 4055 41094 4075
rect 41113 4055 41129 4075
rect 41087 4047 41129 4055
rect 41157 4075 41198 4077
rect 41157 4055 41171 4075
rect 41190 4055 41198 4075
rect 41157 4047 41198 4055
rect 41087 4041 41198 4047
rect 41030 4019 41279 4041
rect 41030 3988 41067 4019
rect 41243 4017 41279 4019
rect 41243 3988 41280 4017
rect 40482 3979 40517 3980
rect 40459 3974 40517 3979
rect 40459 3954 40462 3974
rect 40482 3960 40517 3974
rect 40537 3960 40546 3980
rect 40482 3952 40546 3960
rect 40508 3951 40546 3952
rect 40509 3950 40546 3951
rect 40612 3984 40648 3985
rect 40720 3984 40756 3985
rect 40612 3976 40756 3984
rect 40612 3956 40620 3976
rect 40640 3956 40728 3976
rect 40748 3956 40756 3976
rect 40612 3950 40756 3956
rect 40822 3980 40860 3988
rect 40928 3984 40964 3985
rect 40822 3960 40831 3980
rect 40851 3960 40860 3980
rect 40822 3951 40860 3960
rect 40879 3977 40964 3984
rect 40879 3957 40886 3977
rect 40907 3976 40964 3977
rect 40907 3957 40936 3976
rect 40879 3956 40936 3957
rect 40956 3956 40964 3976
rect 40822 3950 40859 3951
rect 40879 3950 40964 3956
rect 41030 3980 41068 3988
rect 41141 3984 41177 3985
rect 41030 3960 41039 3980
rect 41059 3960 41068 3980
rect 41030 3951 41068 3960
rect 41092 3976 41177 3984
rect 41092 3956 41149 3976
rect 41169 3956 41177 3976
rect 41030 3950 41067 3951
rect 41092 3950 41177 3956
rect 41243 3980 41281 3988
rect 41243 3960 41252 3980
rect 41272 3960 41281 3980
rect 41243 3951 41281 3960
rect 41321 3965 41393 4175
rect 41463 4209 42663 4239
rect 41463 4208 41907 4209
rect 41463 4206 41631 4208
rect 41321 3951 41404 3965
rect 41243 3950 41280 3951
rect 40666 3929 40702 3950
rect 41092 3929 41123 3950
rect 41321 3929 41338 3951
rect 40499 3925 40599 3929
rect 40499 3921 40561 3925
rect 40499 3895 40506 3921
rect 40532 3899 40561 3921
rect 40587 3899 40599 3925
rect 40532 3895 40599 3899
rect 40499 3892 40599 3895
rect 40667 3892 40702 3929
rect 40764 3926 41123 3929
rect 40764 3921 40986 3926
rect 40764 3897 40777 3921
rect 40801 3902 40986 3921
rect 41010 3902 41123 3926
rect 40801 3897 41123 3902
rect 40764 3893 41123 3897
rect 41190 3921 41338 3929
rect 41190 3901 41201 3921
rect 41221 3918 41338 3921
rect 41391 3918 41404 3951
rect 41221 3901 41404 3918
rect 41190 3894 41404 3901
rect 41190 3893 41231 3894
rect 41321 3893 41404 3894
rect 40666 3867 40702 3892
rect 40514 3840 40551 3841
rect 40610 3840 40647 3841
rect 40666 3840 40673 3867
rect 40414 3831 40552 3840
rect 40414 3811 40523 3831
rect 40543 3811 40552 3831
rect 40414 3804 40552 3811
rect 40610 3837 40673 3840
rect 40694 3840 40702 3867
rect 40721 3840 40758 3841
rect 40694 3837 40758 3840
rect 40610 3831 40758 3837
rect 40610 3811 40619 3831
rect 40639 3811 40729 3831
rect 40749 3811 40758 3831
rect 40414 3802 40510 3804
rect 40610 3801 40758 3811
rect 40817 3831 40854 3841
rect 40929 3840 40966 3841
rect 40910 3838 40966 3840
rect 40817 3811 40825 3831
rect 40845 3811 40854 3831
rect 40666 3800 40702 3801
rect 40514 3669 40551 3670
rect 40817 3669 40854 3811
rect 40879 3831 40966 3838
rect 40879 3828 40937 3831
rect 40879 3808 40884 3828
rect 40905 3811 40937 3828
rect 40957 3811 40966 3831
rect 40905 3808 40966 3811
rect 40879 3801 40966 3808
rect 41025 3831 41062 3841
rect 41025 3811 41033 3831
rect 41053 3811 41062 3831
rect 40879 3800 40910 3801
rect 41025 3732 41062 3811
rect 41092 3840 41123 3893
rect 41329 3860 41343 3893
rect 41396 3860 41404 3893
rect 41329 3854 41404 3860
rect 41329 3849 41399 3854
rect 41142 3840 41179 3841
rect 41092 3831 41179 3840
rect 41092 3811 41150 3831
rect 41170 3811 41179 3831
rect 41092 3801 41179 3811
rect 41238 3831 41275 3841
rect 41463 3836 41490 4206
rect 41530 3976 41594 3988
rect 41870 3984 41907 4208
rect 42378 4189 42442 4191
rect 42374 4177 42442 4189
rect 42374 4144 42385 4177
rect 42425 4144 42442 4177
rect 42374 4134 42442 4144
rect 42135 4073 42246 4088
rect 42135 4071 42177 4073
rect 42135 4051 42142 4071
rect 42161 4051 42177 4071
rect 42135 4043 42177 4051
rect 42205 4071 42246 4073
rect 42205 4051 42219 4071
rect 42238 4051 42246 4071
rect 42205 4043 42246 4051
rect 42135 4037 42246 4043
rect 42078 4015 42327 4037
rect 42078 3984 42115 4015
rect 42291 4013 42327 4015
rect 42291 3984 42328 4013
rect 41530 3975 41565 3976
rect 41507 3970 41565 3975
rect 41507 3950 41510 3970
rect 41530 3956 41565 3970
rect 41585 3956 41594 3976
rect 41530 3948 41594 3956
rect 41556 3947 41594 3948
rect 41557 3946 41594 3947
rect 41660 3980 41696 3981
rect 41768 3980 41804 3981
rect 41660 3972 41804 3980
rect 41660 3952 41668 3972
rect 41688 3952 41776 3972
rect 41796 3952 41804 3972
rect 41660 3946 41804 3952
rect 41870 3976 41908 3984
rect 41976 3980 42012 3981
rect 41870 3956 41879 3976
rect 41899 3956 41908 3976
rect 41870 3947 41908 3956
rect 41927 3973 42012 3980
rect 41927 3953 41934 3973
rect 41955 3972 42012 3973
rect 41955 3953 41984 3972
rect 41927 3952 41984 3953
rect 42004 3952 42012 3972
rect 41870 3946 41907 3947
rect 41927 3946 42012 3952
rect 42078 3976 42116 3984
rect 42189 3980 42225 3981
rect 42078 3956 42087 3976
rect 42107 3956 42116 3976
rect 42078 3947 42116 3956
rect 42140 3972 42225 3980
rect 42140 3952 42197 3972
rect 42217 3952 42225 3972
rect 42078 3946 42115 3947
rect 42140 3946 42225 3952
rect 42291 3976 42329 3984
rect 42291 3956 42300 3976
rect 42320 3956 42329 3976
rect 42291 3947 42329 3956
rect 42378 3950 42442 4134
rect 42598 4008 42663 4209
rect 42598 3990 42620 4008
rect 42638 3990 42663 4008
rect 42598 3971 42663 3990
rect 42291 3946 42328 3947
rect 41714 3925 41750 3946
rect 42140 3925 42171 3946
rect 42378 3941 42386 3950
rect 42375 3925 42386 3941
rect 41547 3921 41647 3925
rect 41547 3917 41609 3921
rect 41547 3891 41554 3917
rect 41580 3895 41609 3917
rect 41635 3895 41647 3921
rect 41580 3891 41647 3895
rect 41547 3888 41647 3891
rect 41715 3888 41750 3925
rect 41812 3922 42171 3925
rect 41812 3917 42034 3922
rect 41812 3893 41825 3917
rect 41849 3898 42034 3917
rect 42058 3898 42171 3922
rect 41849 3893 42171 3898
rect 41812 3889 42171 3893
rect 42238 3917 42386 3925
rect 42238 3897 42249 3917
rect 42269 3908 42386 3917
rect 42435 3941 42442 3950
rect 42435 3908 42443 3941
rect 42269 3897 42443 3908
rect 42238 3890 42443 3897
rect 42238 3889 42279 3890
rect 41714 3863 41750 3888
rect 41562 3836 41599 3837
rect 41658 3836 41695 3837
rect 41714 3836 41721 3863
rect 41238 3811 41246 3831
rect 41266 3811 41275 3831
rect 41092 3800 41123 3801
rect 41087 3732 41197 3745
rect 41238 3732 41275 3811
rect 41462 3827 41600 3836
rect 41462 3807 41571 3827
rect 41591 3807 41600 3827
rect 41462 3800 41600 3807
rect 41658 3833 41721 3836
rect 41742 3836 41750 3863
rect 41769 3836 41806 3837
rect 41742 3833 41806 3836
rect 41658 3827 41806 3833
rect 41658 3807 41667 3827
rect 41687 3807 41777 3827
rect 41797 3807 41806 3827
rect 41462 3798 41558 3800
rect 41658 3797 41806 3807
rect 41865 3827 41902 3837
rect 41977 3836 42014 3837
rect 41958 3834 42014 3836
rect 41865 3807 41873 3827
rect 41893 3807 41902 3827
rect 41714 3796 41750 3797
rect 41025 3730 41275 3732
rect 41025 3727 41126 3730
rect 41025 3708 41090 3727
rect 41087 3700 41090 3708
rect 41119 3700 41126 3727
rect 41154 3703 41164 3730
rect 41193 3708 41275 3730
rect 41193 3703 41197 3708
rect 41154 3700 41197 3703
rect 41087 3686 41197 3700
rect 40513 3668 40854 3669
rect 40438 3663 40854 3668
rect 41562 3665 41599 3666
rect 41865 3665 41902 3807
rect 41927 3827 42014 3834
rect 41927 3824 41985 3827
rect 41927 3804 41932 3824
rect 41953 3807 41985 3824
rect 42005 3807 42014 3827
rect 41953 3804 42014 3807
rect 41927 3797 42014 3804
rect 42073 3827 42110 3837
rect 42073 3807 42081 3827
rect 42101 3807 42110 3827
rect 41927 3796 41958 3797
rect 42073 3728 42110 3807
rect 42140 3836 42171 3889
rect 42375 3887 42443 3890
rect 42375 3845 42387 3887
rect 42436 3845 42443 3887
rect 42190 3836 42227 3837
rect 42140 3827 42227 3836
rect 42140 3807 42198 3827
rect 42218 3807 42227 3827
rect 42140 3797 42227 3807
rect 42286 3827 42323 3837
rect 42375 3832 42443 3845
rect 42598 3909 42663 3926
rect 42598 3891 42622 3909
rect 42640 3891 42663 3909
rect 42286 3807 42294 3827
rect 42314 3807 42323 3827
rect 42140 3796 42171 3797
rect 42135 3728 42245 3741
rect 42286 3728 42323 3807
rect 42598 3752 42663 3891
rect 42598 3746 42620 3752
rect 42073 3726 42323 3728
rect 42073 3723 42174 3726
rect 42073 3704 42138 3723
rect 42135 3696 42138 3704
rect 42167 3696 42174 3723
rect 42202 3699 42212 3726
rect 42241 3704 42323 3726
rect 42352 3734 42620 3746
rect 42638 3734 42663 3752
rect 42352 3711 42663 3734
rect 42352 3710 42407 3711
rect 42241 3699 42245 3704
rect 42202 3696 42245 3699
rect 42135 3682 42245 3696
rect 41561 3664 41902 3665
rect 40438 3643 40441 3663
rect 40461 3643 40854 3663
rect 41486 3663 41902 3664
rect 42352 3663 42395 3710
rect 41486 3659 42395 3663
rect 40805 3610 40850 3643
rect 41486 3639 41489 3659
rect 41509 3639 42395 3659
rect 41863 3634 42395 3639
rect 42603 3653 42662 3675
rect 42603 3635 42622 3653
rect 42640 3635 42662 3653
rect 41651 3610 41750 3612
rect 40805 3600 41750 3610
rect 40805 3574 41673 3600
rect 40806 3573 41673 3574
rect 41651 3562 41673 3573
rect 41698 3565 41717 3600
rect 41742 3565 41750 3600
rect 41698 3562 41750 3565
rect 42603 3564 42662 3635
rect 41651 3554 41750 3562
rect 41677 3553 41749 3554
rect 41331 3527 41398 3546
rect 41331 3506 41348 3527
rect 40212 3328 40292 3370
rect 41329 3461 41348 3506
rect 41378 3506 41398 3527
rect 41378 3461 41399 3506
rect 41868 3503 41909 3505
rect 42140 3503 42244 3505
rect 42600 3503 42664 3564
rect 39273 3217 39309 3218
rect 39165 3209 39309 3217
rect 39165 3189 39173 3209
rect 39193 3189 39281 3209
rect 39301 3189 39309 3209
rect 39165 3183 39309 3189
rect 39375 3213 39413 3221
rect 39481 3217 39517 3218
rect 39375 3193 39384 3213
rect 39404 3193 39413 3213
rect 39375 3184 39413 3193
rect 39432 3210 39517 3217
rect 39432 3190 39439 3210
rect 39460 3209 39517 3210
rect 39460 3190 39489 3209
rect 39432 3189 39489 3190
rect 39509 3189 39517 3209
rect 39375 3183 39412 3184
rect 39432 3183 39517 3189
rect 39583 3213 39621 3221
rect 39694 3217 39730 3218
rect 39583 3193 39592 3213
rect 39612 3193 39621 3213
rect 39583 3184 39621 3193
rect 39645 3209 39730 3217
rect 39645 3189 39702 3209
rect 39722 3189 39730 3209
rect 39583 3183 39620 3184
rect 39645 3183 39730 3189
rect 39796 3213 39834 3221
rect 39796 3193 39805 3213
rect 39825 3193 39834 3213
rect 39796 3184 39834 3193
rect 40034 3201 40120 3237
rect 39796 3183 39833 3184
rect 39219 3162 39255 3183
rect 39645 3162 39676 3183
rect 39872 3162 39918 3166
rect 39052 3158 39152 3162
rect 39052 3154 39114 3158
rect 39052 3128 39059 3154
rect 39085 3132 39114 3154
rect 39140 3132 39152 3158
rect 39085 3128 39152 3132
rect 39052 3125 39152 3128
rect 39220 3125 39255 3162
rect 39317 3159 39676 3162
rect 39317 3154 39539 3159
rect 39317 3130 39330 3154
rect 39354 3135 39539 3154
rect 39563 3135 39676 3159
rect 39354 3130 39676 3135
rect 39317 3126 39676 3130
rect 39743 3154 39918 3162
rect 39743 3134 39754 3154
rect 39774 3134 39918 3154
rect 40034 3160 40051 3201
rect 40105 3160 40120 3201
rect 40034 3141 40120 3160
rect 39743 3127 39918 3134
rect 39743 3126 39784 3127
rect 39219 3100 39255 3125
rect 39067 3073 39104 3074
rect 39163 3073 39200 3074
rect 39219 3073 39226 3100
rect 38967 3064 39105 3073
rect 38967 3044 39076 3064
rect 39096 3044 39105 3064
rect 38967 3037 39105 3044
rect 39163 3070 39226 3073
rect 39247 3073 39255 3100
rect 39274 3073 39311 3074
rect 39247 3070 39311 3073
rect 39163 3064 39311 3070
rect 39163 3044 39172 3064
rect 39192 3044 39282 3064
rect 39302 3044 39311 3064
rect 38967 3035 39063 3037
rect 39163 3034 39311 3044
rect 39370 3064 39407 3074
rect 39482 3073 39519 3074
rect 39463 3071 39519 3073
rect 39370 3044 39378 3064
rect 39398 3044 39407 3064
rect 39219 3033 39255 3034
rect 39067 2902 39104 2903
rect 39370 2902 39407 3044
rect 39432 3064 39519 3071
rect 39432 3061 39490 3064
rect 39432 3041 39437 3061
rect 39458 3044 39490 3061
rect 39510 3044 39519 3064
rect 39458 3041 39519 3044
rect 39432 3034 39519 3041
rect 39578 3064 39615 3074
rect 39578 3044 39586 3064
rect 39606 3044 39615 3064
rect 39432 3033 39463 3034
rect 39578 2965 39615 3044
rect 39645 3073 39676 3126
rect 39695 3073 39732 3074
rect 39645 3064 39732 3073
rect 39645 3044 39703 3064
rect 39723 3044 39732 3064
rect 39645 3034 39732 3044
rect 39791 3064 39828 3074
rect 39791 3044 39799 3064
rect 39819 3044 39828 3064
rect 39645 3033 39676 3034
rect 39640 2965 39750 2978
rect 39791 2965 39828 3044
rect 39872 3044 39918 3127
rect 40212 3044 40287 3328
rect 41329 3253 41399 3461
rect 41461 3468 42664 3503
rect 41461 3454 41489 3468
rect 41463 3323 41489 3454
rect 41868 3465 42664 3468
rect 41321 3202 41401 3253
rect 41321 3176 41337 3202
rect 41377 3176 41401 3202
rect 41321 3157 41401 3176
rect 41321 3131 41340 3157
rect 41380 3131 41401 3157
rect 41321 3104 41401 3131
rect 41321 3078 41344 3104
rect 41384 3078 41401 3104
rect 41321 3067 41401 3078
rect 41463 3068 41490 3323
rect 41868 3315 41909 3465
rect 42140 3459 42244 3465
rect 42600 3462 42664 3465
rect 42335 3403 42456 3421
rect 42335 3401 42406 3403
rect 42335 3360 42350 3401
rect 42387 3362 42406 3401
rect 42443 3362 42456 3403
rect 42387 3360 42456 3362
rect 42335 3350 42456 3360
rect 41530 3208 41594 3220
rect 41870 3216 41907 3315
rect 42135 3305 42246 3318
rect 42135 3303 42177 3305
rect 42135 3283 42142 3303
rect 42161 3283 42177 3303
rect 42135 3275 42177 3283
rect 42205 3303 42246 3305
rect 42205 3283 42219 3303
rect 42238 3283 42246 3303
rect 42205 3275 42246 3283
rect 42135 3269 42246 3275
rect 42078 3247 42327 3269
rect 42078 3216 42115 3247
rect 42291 3245 42327 3247
rect 42291 3216 42328 3245
rect 41530 3207 41565 3208
rect 41507 3202 41565 3207
rect 41507 3182 41510 3202
rect 41530 3188 41565 3202
rect 41585 3188 41594 3208
rect 41530 3180 41594 3188
rect 41556 3179 41594 3180
rect 41557 3178 41594 3179
rect 41660 3212 41696 3213
rect 41768 3212 41804 3213
rect 41660 3204 41804 3212
rect 41660 3184 41668 3204
rect 41688 3184 41776 3204
rect 41796 3184 41804 3204
rect 41660 3178 41804 3184
rect 41870 3208 41908 3216
rect 41976 3212 42012 3213
rect 41870 3188 41879 3208
rect 41899 3188 41908 3208
rect 41870 3179 41908 3188
rect 41927 3205 42012 3212
rect 41927 3185 41934 3205
rect 41955 3204 42012 3205
rect 41955 3185 41984 3204
rect 41927 3184 41984 3185
rect 42004 3184 42012 3204
rect 41870 3178 41907 3179
rect 41927 3178 42012 3184
rect 42078 3208 42116 3216
rect 42189 3212 42225 3213
rect 42078 3188 42087 3208
rect 42107 3188 42116 3208
rect 42078 3179 42116 3188
rect 42140 3204 42225 3212
rect 42140 3184 42197 3204
rect 42217 3184 42225 3204
rect 42078 3178 42115 3179
rect 42140 3178 42225 3184
rect 42291 3208 42329 3216
rect 42291 3188 42300 3208
rect 42320 3188 42329 3208
rect 42384 3198 42449 3350
rect 42602 3324 42657 3462
rect 42291 3179 42329 3188
rect 42382 3191 42449 3198
rect 42291 3178 42328 3179
rect 41714 3157 41750 3178
rect 42140 3157 42171 3178
rect 42382 3170 42399 3191
rect 42435 3170 42449 3191
rect 42601 3211 42657 3324
rect 42601 3193 42620 3211
rect 42638 3193 42657 3211
rect 42601 3173 42657 3193
rect 42382 3157 42449 3170
rect 41547 3153 41647 3157
rect 41547 3149 41609 3153
rect 41547 3123 41554 3149
rect 41580 3127 41609 3149
rect 41635 3127 41647 3153
rect 41580 3123 41647 3127
rect 41547 3120 41647 3123
rect 41715 3120 41750 3157
rect 41812 3154 42171 3157
rect 41812 3149 42034 3154
rect 41812 3125 41825 3149
rect 41849 3130 42034 3149
rect 42058 3130 42171 3154
rect 41849 3125 42171 3130
rect 41812 3121 42171 3125
rect 42238 3151 42449 3157
rect 42238 3149 42399 3151
rect 42238 3129 42249 3149
rect 42269 3129 42399 3149
rect 42238 3122 42399 3129
rect 42238 3121 42279 3122
rect 41714 3095 41750 3120
rect 41562 3068 41599 3069
rect 41658 3068 41695 3069
rect 41714 3068 41721 3095
rect 39872 3009 40287 3044
rect 41462 3059 41600 3068
rect 41462 3039 41571 3059
rect 41591 3039 41600 3059
rect 41462 3032 41600 3039
rect 41658 3065 41721 3068
rect 41742 3068 41750 3095
rect 41769 3068 41806 3069
rect 41742 3065 41806 3068
rect 41658 3059 41806 3065
rect 41658 3039 41667 3059
rect 41687 3039 41777 3059
rect 41797 3039 41806 3059
rect 41462 3030 41558 3032
rect 41658 3029 41806 3039
rect 41865 3059 41902 3069
rect 41977 3068 42014 3069
rect 41958 3066 42014 3068
rect 41865 3039 41873 3059
rect 41893 3039 41902 3059
rect 41714 3028 41750 3029
rect 39872 3008 39918 3009
rect 39578 2963 39828 2965
rect 39578 2960 39679 2963
rect 39578 2941 39643 2960
rect 39640 2933 39643 2941
rect 39672 2933 39679 2960
rect 39707 2936 39717 2963
rect 39746 2941 39828 2963
rect 40212 2957 40287 3009
rect 39746 2936 39750 2941
rect 39707 2933 39750 2936
rect 39640 2919 39750 2933
rect 39066 2901 39407 2902
rect 38991 2896 39407 2901
rect 38991 2876 38994 2896
rect 39014 2876 39408 2896
rect 35471 2467 38539 2492
rect 35471 2402 38334 2467
rect 38465 2402 38539 2467
rect 35471 2385 38539 2402
rect 39365 2372 39408 2876
rect 40025 2787 40120 2807
rect 40025 2743 40045 2787
rect 40105 2743 40120 2787
rect 40025 2447 40120 2743
rect 40025 2406 40058 2447
rect 40094 2406 40120 2447
rect 40220 2486 40282 2957
rect 41562 2897 41599 2898
rect 41865 2897 41902 3039
rect 41927 3059 42014 3066
rect 41927 3056 41985 3059
rect 41927 3036 41932 3056
rect 41953 3039 41985 3056
rect 42005 3039 42014 3059
rect 41953 3036 42014 3039
rect 41927 3029 42014 3036
rect 42073 3059 42110 3069
rect 42073 3039 42081 3059
rect 42101 3039 42110 3059
rect 41927 3028 41958 3029
rect 42073 2960 42110 3039
rect 42140 3068 42171 3121
rect 42384 3114 42399 3122
rect 42439 3114 42449 3151
rect 42384 3105 42449 3114
rect 42597 3112 42662 3133
rect 42597 3094 42622 3112
rect 42640 3094 42662 3112
rect 42190 3068 42227 3069
rect 42140 3059 42227 3068
rect 42140 3039 42198 3059
rect 42218 3039 42227 3059
rect 42140 3029 42227 3039
rect 42286 3059 42323 3069
rect 42286 3039 42294 3059
rect 42314 3039 42323 3059
rect 42140 3028 42171 3029
rect 42135 2960 42245 2973
rect 42286 2960 42323 3039
rect 42597 3018 42662 3094
rect 42073 2958 42323 2960
rect 42073 2955 42174 2958
rect 42073 2936 42138 2955
rect 42135 2928 42138 2936
rect 42167 2928 42174 2955
rect 42202 2931 42212 2958
rect 42241 2936 42323 2958
rect 42346 2983 42663 3018
rect 42241 2931 42245 2936
rect 42202 2928 42245 2931
rect 42135 2914 42245 2928
rect 41561 2896 41902 2897
rect 41486 2894 41902 2896
rect 42346 2894 42386 2983
rect 42597 2956 42662 2983
rect 42597 2938 42620 2956
rect 42638 2938 42662 2956
rect 42597 2918 42662 2938
rect 41483 2891 42386 2894
rect 41483 2871 41489 2891
rect 41509 2871 42386 2891
rect 41483 2867 42386 2871
rect 42346 2864 42386 2867
rect 42598 2857 42663 2878
rect 40816 2849 41477 2850
rect 40816 2842 41750 2849
rect 40816 2841 41722 2842
rect 40816 2821 41667 2841
rect 41699 2822 41722 2841
rect 41747 2822 41750 2842
rect 41699 2821 41750 2822
rect 40816 2814 41750 2821
rect 40415 2772 40583 2773
rect 40818 2772 40857 2814
rect 41646 2812 41750 2814
rect 41715 2810 41750 2812
rect 42598 2839 42622 2857
rect 42640 2839 42663 2857
rect 42598 2792 42663 2839
rect 40415 2746 40859 2772
rect 40415 2744 40583 2746
rect 40220 2467 40284 2486
rect 40220 2428 40237 2467
rect 40271 2428 40284 2467
rect 40220 2409 40284 2428
rect 40025 2380 40120 2406
rect 40415 2393 40442 2744
rect 40818 2740 40859 2746
rect 40482 2533 40546 2545
rect 40822 2541 40859 2740
rect 41321 2767 41393 2784
rect 41321 2728 41329 2767
rect 41374 2728 41393 2767
rect 41087 2630 41198 2645
rect 41087 2628 41129 2630
rect 41087 2608 41094 2628
rect 41113 2608 41129 2628
rect 41087 2600 41129 2608
rect 41157 2628 41198 2630
rect 41157 2608 41171 2628
rect 41190 2608 41198 2628
rect 41157 2600 41198 2608
rect 41087 2594 41198 2600
rect 41030 2572 41279 2594
rect 41030 2541 41067 2572
rect 41243 2570 41279 2572
rect 41243 2541 41280 2570
rect 40482 2532 40517 2533
rect 40459 2527 40517 2532
rect 40459 2507 40462 2527
rect 40482 2513 40517 2527
rect 40537 2513 40546 2533
rect 40482 2505 40546 2513
rect 40508 2504 40546 2505
rect 40509 2503 40546 2504
rect 40612 2537 40648 2538
rect 40720 2537 40756 2538
rect 40612 2529 40756 2537
rect 40612 2509 40620 2529
rect 40640 2509 40728 2529
rect 40748 2509 40756 2529
rect 40612 2503 40756 2509
rect 40822 2533 40860 2541
rect 40928 2537 40964 2538
rect 40822 2513 40831 2533
rect 40851 2513 40860 2533
rect 40822 2504 40860 2513
rect 40879 2530 40964 2537
rect 40879 2510 40886 2530
rect 40907 2529 40964 2530
rect 40907 2510 40936 2529
rect 40879 2509 40936 2510
rect 40956 2509 40964 2529
rect 40822 2503 40859 2504
rect 40879 2503 40964 2509
rect 41030 2533 41068 2541
rect 41141 2537 41177 2538
rect 41030 2513 41039 2533
rect 41059 2513 41068 2533
rect 41030 2504 41068 2513
rect 41092 2529 41177 2537
rect 41092 2509 41149 2529
rect 41169 2509 41177 2529
rect 41030 2503 41067 2504
rect 41092 2503 41177 2509
rect 41243 2533 41281 2541
rect 41243 2513 41252 2533
rect 41272 2513 41281 2533
rect 41243 2504 41281 2513
rect 41321 2518 41393 2728
rect 41463 2762 42663 2792
rect 41463 2761 41907 2762
rect 41463 2759 41631 2761
rect 41321 2504 41404 2518
rect 41243 2503 41280 2504
rect 40666 2482 40702 2503
rect 41092 2482 41123 2503
rect 41321 2482 41338 2504
rect 40499 2478 40599 2482
rect 40499 2474 40561 2478
rect 40499 2448 40506 2474
rect 40532 2452 40561 2474
rect 40587 2452 40599 2478
rect 40532 2448 40599 2452
rect 40499 2445 40599 2448
rect 40667 2445 40702 2482
rect 40764 2479 41123 2482
rect 40764 2474 40986 2479
rect 40764 2450 40777 2474
rect 40801 2455 40986 2474
rect 41010 2455 41123 2479
rect 40801 2450 41123 2455
rect 40764 2446 41123 2450
rect 41190 2474 41338 2482
rect 41190 2454 41201 2474
rect 41221 2471 41338 2474
rect 41391 2471 41404 2504
rect 41221 2454 41404 2471
rect 41190 2447 41404 2454
rect 41190 2446 41231 2447
rect 41321 2446 41404 2447
rect 40666 2420 40702 2445
rect 40514 2393 40551 2394
rect 40610 2393 40647 2394
rect 40666 2393 40673 2420
rect 40414 2384 40552 2393
rect 35226 2286 35383 2299
rect 35226 2282 35387 2286
rect 34106 2136 34132 2241
rect 35226 2175 35267 2282
rect 35367 2175 35387 2282
rect 35226 2146 35387 2175
rect 39363 2163 39412 2372
rect 40414 2364 40523 2384
rect 40543 2364 40552 2384
rect 40414 2357 40552 2364
rect 40610 2390 40673 2393
rect 40694 2393 40702 2420
rect 40721 2393 40758 2394
rect 40694 2390 40758 2393
rect 40610 2384 40758 2390
rect 40610 2364 40619 2384
rect 40639 2364 40729 2384
rect 40749 2364 40758 2384
rect 40414 2355 40510 2357
rect 40610 2354 40758 2364
rect 40817 2384 40854 2394
rect 40929 2393 40966 2394
rect 40910 2391 40966 2393
rect 40817 2364 40825 2384
rect 40845 2364 40854 2384
rect 40666 2353 40702 2354
rect 40514 2222 40551 2223
rect 40817 2222 40854 2364
rect 40879 2384 40966 2391
rect 40879 2381 40937 2384
rect 40879 2361 40884 2381
rect 40905 2364 40937 2381
rect 40957 2364 40966 2384
rect 40905 2361 40966 2364
rect 40879 2354 40966 2361
rect 41025 2384 41062 2394
rect 41025 2364 41033 2384
rect 41053 2364 41062 2384
rect 40879 2353 40910 2354
rect 41025 2285 41062 2364
rect 41092 2393 41123 2446
rect 41329 2413 41343 2446
rect 41396 2413 41404 2446
rect 41329 2407 41404 2413
rect 41329 2402 41399 2407
rect 41142 2393 41179 2394
rect 41092 2384 41179 2393
rect 41092 2364 41150 2384
rect 41170 2364 41179 2384
rect 41092 2354 41179 2364
rect 41238 2384 41275 2394
rect 41463 2389 41490 2759
rect 41530 2529 41594 2541
rect 41870 2537 41907 2761
rect 42378 2742 42442 2744
rect 42374 2730 42442 2742
rect 42374 2697 42385 2730
rect 42425 2697 42442 2730
rect 42374 2687 42442 2697
rect 42135 2626 42246 2641
rect 42135 2624 42177 2626
rect 42135 2604 42142 2624
rect 42161 2604 42177 2624
rect 42135 2596 42177 2604
rect 42205 2624 42246 2626
rect 42205 2604 42219 2624
rect 42238 2604 42246 2624
rect 42205 2596 42246 2604
rect 42135 2590 42246 2596
rect 42078 2568 42327 2590
rect 42078 2537 42115 2568
rect 42291 2566 42327 2568
rect 42291 2537 42328 2566
rect 41530 2528 41565 2529
rect 41507 2523 41565 2528
rect 41507 2503 41510 2523
rect 41530 2509 41565 2523
rect 41585 2509 41594 2529
rect 41530 2501 41594 2509
rect 41556 2500 41594 2501
rect 41557 2499 41594 2500
rect 41660 2533 41696 2534
rect 41768 2533 41804 2534
rect 41660 2525 41804 2533
rect 41660 2505 41668 2525
rect 41688 2505 41776 2525
rect 41796 2505 41804 2525
rect 41660 2499 41804 2505
rect 41870 2529 41908 2537
rect 41976 2533 42012 2534
rect 41870 2509 41879 2529
rect 41899 2509 41908 2529
rect 41870 2500 41908 2509
rect 41927 2526 42012 2533
rect 41927 2506 41934 2526
rect 41955 2525 42012 2526
rect 41955 2506 41984 2525
rect 41927 2505 41984 2506
rect 42004 2505 42012 2525
rect 41870 2499 41907 2500
rect 41927 2499 42012 2505
rect 42078 2529 42116 2537
rect 42189 2533 42225 2534
rect 42078 2509 42087 2529
rect 42107 2509 42116 2529
rect 42078 2500 42116 2509
rect 42140 2525 42225 2533
rect 42140 2505 42197 2525
rect 42217 2505 42225 2525
rect 42078 2499 42115 2500
rect 42140 2499 42225 2505
rect 42291 2529 42329 2537
rect 42291 2509 42300 2529
rect 42320 2509 42329 2529
rect 42291 2500 42329 2509
rect 42378 2503 42442 2687
rect 42598 2561 42663 2762
rect 42598 2543 42620 2561
rect 42638 2543 42663 2561
rect 42598 2524 42663 2543
rect 42291 2499 42328 2500
rect 41714 2478 41750 2499
rect 42140 2478 42171 2499
rect 42378 2494 42386 2503
rect 42375 2478 42386 2494
rect 41547 2474 41647 2478
rect 41547 2470 41609 2474
rect 41547 2444 41554 2470
rect 41580 2448 41609 2470
rect 41635 2448 41647 2474
rect 41580 2444 41647 2448
rect 41547 2441 41647 2444
rect 41715 2441 41750 2478
rect 41812 2475 42171 2478
rect 41812 2470 42034 2475
rect 41812 2446 41825 2470
rect 41849 2451 42034 2470
rect 42058 2451 42171 2475
rect 41849 2446 42171 2451
rect 41812 2442 42171 2446
rect 42238 2470 42386 2478
rect 42238 2450 42249 2470
rect 42269 2461 42386 2470
rect 42435 2494 42442 2503
rect 42435 2461 42443 2494
rect 42269 2450 42443 2461
rect 42238 2443 42443 2450
rect 42238 2442 42279 2443
rect 41714 2416 41750 2441
rect 41562 2389 41599 2390
rect 41658 2389 41695 2390
rect 41714 2389 41721 2416
rect 41238 2364 41246 2384
rect 41266 2364 41275 2384
rect 41092 2353 41123 2354
rect 41087 2285 41197 2298
rect 41238 2285 41275 2364
rect 41462 2380 41600 2389
rect 41462 2360 41571 2380
rect 41591 2360 41600 2380
rect 41462 2353 41600 2360
rect 41658 2386 41721 2389
rect 41742 2389 41750 2416
rect 41769 2389 41806 2390
rect 41742 2386 41806 2389
rect 41658 2380 41806 2386
rect 41658 2360 41667 2380
rect 41687 2360 41777 2380
rect 41797 2360 41806 2380
rect 41462 2351 41558 2353
rect 41658 2350 41806 2360
rect 41865 2380 41902 2390
rect 41977 2389 42014 2390
rect 41958 2387 42014 2389
rect 41865 2360 41873 2380
rect 41893 2360 41902 2380
rect 41714 2349 41750 2350
rect 41025 2283 41275 2285
rect 41025 2280 41126 2283
rect 41025 2261 41090 2280
rect 41087 2253 41090 2261
rect 41119 2253 41126 2280
rect 41154 2256 41164 2283
rect 41193 2261 41275 2283
rect 41193 2256 41197 2261
rect 41154 2253 41197 2256
rect 41087 2239 41197 2253
rect 40513 2221 40854 2222
rect 40438 2216 40854 2221
rect 41562 2218 41599 2219
rect 41865 2218 41902 2360
rect 41927 2380 42014 2387
rect 41927 2377 41985 2380
rect 41927 2357 41932 2377
rect 41953 2360 41985 2377
rect 42005 2360 42014 2380
rect 41953 2357 42014 2360
rect 41927 2350 42014 2357
rect 42073 2380 42110 2390
rect 42073 2360 42081 2380
rect 42101 2360 42110 2380
rect 41927 2349 41958 2350
rect 42073 2281 42110 2360
rect 42140 2389 42171 2442
rect 42375 2440 42443 2443
rect 42375 2398 42387 2440
rect 42436 2398 42443 2440
rect 42190 2389 42227 2390
rect 42140 2380 42227 2389
rect 42140 2360 42198 2380
rect 42218 2360 42227 2380
rect 42140 2350 42227 2360
rect 42286 2380 42323 2390
rect 42375 2385 42443 2398
rect 42598 2462 42663 2479
rect 42598 2444 42622 2462
rect 42640 2444 42663 2462
rect 42286 2360 42294 2380
rect 42314 2360 42323 2380
rect 42140 2349 42171 2350
rect 42135 2281 42245 2294
rect 42286 2281 42323 2360
rect 42598 2305 42663 2444
rect 42598 2299 42620 2305
rect 42073 2279 42323 2281
rect 42073 2276 42174 2279
rect 42073 2257 42138 2276
rect 42135 2249 42138 2257
rect 42167 2249 42174 2276
rect 42202 2252 42212 2279
rect 42241 2257 42323 2279
rect 42352 2287 42620 2299
rect 42638 2287 42663 2305
rect 42352 2264 42663 2287
rect 42352 2263 42407 2264
rect 42241 2252 42245 2257
rect 42202 2249 42245 2252
rect 42135 2235 42245 2249
rect 41561 2217 41902 2218
rect 40438 2196 40441 2216
rect 40461 2196 40854 2216
rect 41486 2216 41902 2217
rect 42352 2216 42395 2263
rect 41486 2212 42395 2216
rect 34106 2122 34134 2136
rect 35230 2133 35387 2146
rect 39361 2161 40178 2163
rect 40611 2161 40700 2164
rect 39361 2152 40700 2161
rect 32908 2087 34134 2122
rect 39361 2114 40623 2152
rect 40648 2117 40667 2152
rect 40692 2117 40700 2152
rect 40805 2163 40850 2196
rect 41486 2192 41489 2212
rect 41509 2192 42395 2212
rect 41863 2187 42395 2192
rect 42603 2206 42662 2228
rect 42603 2188 42622 2206
rect 42640 2188 42662 2206
rect 41651 2163 41750 2165
rect 40805 2153 41750 2163
rect 40805 2127 41673 2153
rect 40806 2126 41673 2127
rect 40648 2114 40700 2117
rect 39361 2106 40700 2114
rect 41651 2115 41673 2126
rect 41698 2118 41717 2153
rect 41742 2118 41750 2153
rect 41698 2115 41750 2118
rect 41651 2107 41750 2115
rect 41677 2106 41749 2107
rect 39361 2105 40699 2106
rect 39361 2103 40178 2105
rect 39952 2099 40178 2103
rect 11235 1940 21003 2013
rect 22200 1944 31968 2017
rect 7610 1926 7764 1931
rect 11249 1925 21003 1940
rect 22214 1929 31968 1944
rect 32908 2011 32993 2087
rect 33351 2085 33455 2087
rect 33686 2085 33727 2087
rect 42603 2011 42662 2188
rect 32908 1938 42676 2011
rect 18318 1920 18472 1925
rect 29283 1924 29437 1929
rect 32922 1923 42676 1938
rect 39991 1918 40145 1923
rect 10191 786 11078 788
rect 10191 775 11085 786
rect 10191 729 10213 775
rect 10289 729 11085 775
rect 31864 784 32751 786
rect 31864 773 32758 784
rect 10191 716 11085 729
rect 11019 568 11085 716
rect 16276 743 16386 757
rect 16276 741 22349 743
rect 16276 718 22538 741
rect 11660 699 11725 705
rect 11660 651 11675 699
rect 11716 651 11725 699
rect 11660 631 11725 651
rect 16276 662 22334 718
rect 22413 708 22538 718
rect 31864 727 31886 773
rect 31962 727 32758 773
rect 31864 714 32758 727
rect 22413 662 22464 708
rect 16276 657 22464 662
rect 22510 657 22538 708
rect 16276 639 22538 657
rect 16276 634 22349 639
rect 11019 548 11416 568
rect 11436 548 11439 568
rect 11019 543 11439 548
rect 11019 542 11364 543
rect 11019 530 11085 542
rect 11326 541 11363 542
rect 10680 511 10790 525
rect 10680 508 10723 511
rect 10680 503 10684 508
rect 10602 481 10684 503
rect 10713 481 10723 508
rect 10751 484 10758 511
rect 10787 503 10790 511
rect 10787 484 10852 503
rect 10751 481 10852 484
rect 10602 479 10852 481
rect 10602 400 10639 479
rect 10680 466 10790 479
rect 10754 410 10785 411
rect 10602 380 10611 400
rect 10631 380 10639 400
rect 10602 370 10639 380
rect 10698 400 10785 410
rect 10698 380 10707 400
rect 10727 380 10785 400
rect 10698 371 10785 380
rect 10698 370 10735 371
rect 10163 333 10292 340
rect 10163 274 10187 333
rect 10218 274 10249 333
rect 10280 318 10292 333
rect 10754 318 10785 371
rect 10815 400 10852 479
rect 10967 410 10998 411
rect 10815 380 10824 400
rect 10844 380 10852 400
rect 10815 370 10852 380
rect 10911 403 10998 410
rect 10911 400 10972 403
rect 10911 380 10920 400
rect 10940 383 10972 400
rect 10993 383 10998 403
rect 10940 380 10998 383
rect 10911 373 10998 380
rect 11023 400 11060 530
rect 11175 410 11211 411
rect 11023 380 11032 400
rect 11052 380 11060 400
rect 10911 371 10967 373
rect 10911 370 10948 371
rect 11023 370 11060 380
rect 11119 400 11267 410
rect 11367 407 11463 409
rect 11119 380 11128 400
rect 11148 380 11238 400
rect 11258 380 11267 400
rect 11119 374 11267 380
rect 11119 371 11183 374
rect 11119 370 11156 371
rect 11175 344 11183 371
rect 11204 371 11267 374
rect 11325 400 11463 407
rect 11325 380 11334 400
rect 11354 380 11463 400
rect 11325 371 11463 380
rect 11204 344 11211 371
rect 11230 370 11267 371
rect 11326 370 11363 371
rect 11175 319 11211 344
rect 10280 317 10577 318
rect 10646 317 10687 318
rect 10280 310 10687 317
rect 10280 290 10656 310
rect 10676 290 10687 310
rect 10280 282 10687 290
rect 10754 314 11113 318
rect 10754 309 11076 314
rect 10754 285 10867 309
rect 10891 290 11076 309
rect 11100 290 11113 314
rect 10891 285 11113 290
rect 10754 282 11113 285
rect 11175 282 11210 319
rect 11278 316 11378 319
rect 11278 312 11345 316
rect 11278 286 11290 312
rect 11316 290 11345 312
rect 11371 290 11378 316
rect 11316 286 11378 290
rect 11278 282 11378 286
rect 10280 274 10577 282
rect 10163 261 10292 274
rect 10754 261 10785 282
rect 11175 261 11211 282
rect 10164 151 10270 261
rect 10597 260 10634 261
rect 10596 251 10634 260
rect 10596 231 10605 251
rect 10625 231 10634 251
rect 10596 223 10634 231
rect 10700 255 10785 261
rect 10810 260 10847 261
rect 10700 235 10708 255
rect 10728 235 10785 255
rect 10700 227 10785 235
rect 10809 251 10847 260
rect 10809 231 10818 251
rect 10838 231 10847 251
rect 10700 226 10736 227
rect 10809 223 10847 231
rect 10913 255 10998 261
rect 11018 260 11055 261
rect 10913 235 10921 255
rect 10941 254 10998 255
rect 10941 235 10970 254
rect 10913 234 10970 235
rect 10991 234 10998 254
rect 10913 227 10998 234
rect 11017 251 11055 260
rect 11017 231 11026 251
rect 11046 231 11055 251
rect 10913 226 10949 227
rect 11017 223 11055 231
rect 11121 255 11265 261
rect 11121 235 11129 255
rect 11149 235 11184 255
rect 11121 232 11184 235
rect 11204 235 11237 255
rect 11257 235 11265 255
rect 11204 232 11265 235
rect 11121 227 11265 232
rect 11121 226 11157 227
rect 11229 226 11265 227
rect 11331 260 11368 261
rect 11331 259 11369 260
rect 11331 251 11395 259
rect 11331 231 11340 251
rect 11360 237 11395 251
rect 11415 237 11418 257
rect 11360 232 11418 237
rect 11360 231 11395 232
rect 10597 194 10634 223
rect 10598 192 10634 194
rect 10810 192 10847 223
rect 10598 170 10847 192
rect 10160 49 10270 151
rect 10679 164 10790 170
rect 10679 156 10720 164
rect 10679 136 10687 156
rect 10706 136 10720 156
rect 10679 134 10720 136
rect 10748 156 10790 164
rect 10748 136 10764 156
rect 10783 136 10790 156
rect 10748 134 10790 136
rect 10679 119 10790 134
rect 11018 102 11055 223
rect 11331 219 11395 231
rect 11435 109 11462 371
rect 11660 109 11708 631
rect 16276 568 16386 634
rect 20148 572 20217 582
rect 11413 104 11708 109
rect 11294 102 11708 104
rect 11018 76 11708 102
rect 11294 75 11708 76
rect 11413 74 11708 75
rect 11660 69 11708 74
rect 11812 450 16394 568
rect 20148 547 20162 572
rect 20203 565 20217 572
rect 32692 566 32758 714
rect 33333 697 33398 703
rect 33333 649 33348 697
rect 33389 649 33398 697
rect 33333 629 33398 649
rect 20203 555 21751 565
rect 20203 547 22053 555
rect 20148 538 22053 547
rect 21660 535 22053 538
rect 22073 535 22076 555
rect 21660 530 22076 535
rect 32692 546 33089 566
rect 33109 546 33112 566
rect 32692 541 33112 546
rect 32692 540 33037 541
rect 21660 529 22001 530
rect 21317 498 21427 512
rect 21317 495 21360 498
rect 21317 490 21321 495
rect 21239 468 21321 490
rect 21350 468 21360 495
rect 21388 471 21395 498
rect 21424 490 21427 498
rect 21424 471 21489 490
rect 21388 468 21489 471
rect 21239 466 21489 468
rect 10160 -136 10266 49
rect 10160 -137 11505 -136
rect 11812 -137 11940 450
rect 21239 387 21276 466
rect 21317 453 21427 466
rect 21391 397 21422 398
rect 21239 367 21248 387
rect 21268 367 21276 387
rect 21239 357 21276 367
rect 21335 387 21422 397
rect 21335 367 21344 387
rect 21364 367 21422 387
rect 21335 358 21422 367
rect 21335 357 21372 358
rect 20512 319 20816 337
rect 20512 266 20556 319
rect 20753 312 20816 319
rect 20753 306 21185 312
rect 20753 304 21218 306
rect 21391 305 21422 358
rect 21452 387 21489 466
rect 21604 397 21635 398
rect 21452 367 21461 387
rect 21481 367 21489 387
rect 21452 357 21489 367
rect 21548 390 21635 397
rect 21548 387 21609 390
rect 21548 367 21557 387
rect 21577 370 21609 387
rect 21630 370 21635 390
rect 21577 367 21635 370
rect 21548 360 21635 367
rect 21660 387 21697 529
rect 21963 528 22000 529
rect 32692 528 32758 540
rect 32999 539 33036 540
rect 32353 509 32463 523
rect 32353 506 32396 509
rect 32353 501 32357 506
rect 32275 479 32357 501
rect 32386 479 32396 506
rect 32424 482 32431 509
rect 32460 501 32463 509
rect 32460 482 32525 501
rect 32424 479 32525 482
rect 32275 477 32525 479
rect 32275 398 32312 477
rect 32353 464 32463 477
rect 32427 408 32458 409
rect 21812 397 21848 398
rect 21660 367 21669 387
rect 21689 367 21697 387
rect 21548 358 21604 360
rect 21548 357 21585 358
rect 21660 357 21697 367
rect 21756 387 21904 397
rect 22004 394 22100 396
rect 21756 367 21765 387
rect 21785 367 21875 387
rect 21895 367 21904 387
rect 21756 361 21904 367
rect 21756 358 21820 361
rect 21756 357 21793 358
rect 21812 331 21820 358
rect 21841 358 21904 361
rect 21962 387 22100 394
rect 21962 367 21971 387
rect 21991 367 22100 387
rect 32275 378 32284 398
rect 32304 378 32312 398
rect 32275 368 32312 378
rect 32371 398 32458 408
rect 32371 378 32380 398
rect 32400 378 32458 398
rect 32371 369 32458 378
rect 32371 368 32408 369
rect 21962 358 22100 367
rect 21841 331 21848 358
rect 21867 357 21904 358
rect 21963 357 22000 358
rect 21812 306 21848 331
rect 21283 304 21324 305
rect 20753 297 21324 304
rect 20753 277 21293 297
rect 21313 277 21324 297
rect 20753 269 21324 277
rect 21391 301 21750 305
rect 21391 296 21713 301
rect 21391 272 21504 296
rect 21528 277 21713 296
rect 21737 277 21750 301
rect 21528 272 21750 277
rect 21391 269 21750 272
rect 21812 269 21847 306
rect 21915 303 22015 306
rect 21915 299 21982 303
rect 21915 273 21927 299
rect 21953 277 21982 299
rect 22008 277 22015 303
rect 21953 273 22015 277
rect 21915 269 22015 273
rect 20753 267 21185 269
rect 20753 266 20816 267
rect 20512 246 20816 266
rect 21391 248 21422 269
rect 21812 248 21848 269
rect 21234 247 21271 248
rect 21233 238 21271 247
rect 21233 218 21242 238
rect 21262 218 21271 238
rect 21233 210 21271 218
rect 21337 242 21422 248
rect 21447 247 21484 248
rect 21337 222 21345 242
rect 21365 222 21422 242
rect 21337 214 21422 222
rect 21446 238 21484 247
rect 21446 218 21455 238
rect 21475 218 21484 238
rect 21337 213 21373 214
rect 21446 210 21484 218
rect 21550 242 21635 248
rect 21655 247 21692 248
rect 21550 222 21558 242
rect 21578 241 21635 242
rect 21578 222 21607 241
rect 21550 221 21607 222
rect 21628 221 21635 241
rect 21550 214 21635 221
rect 21654 238 21692 247
rect 21654 218 21663 238
rect 21683 218 21692 238
rect 21550 213 21586 214
rect 21654 210 21692 218
rect 21758 243 21902 248
rect 21758 242 21823 243
rect 21758 222 21766 242
rect 21786 222 21823 242
rect 21758 221 21823 222
rect 21841 242 21902 243
rect 21841 222 21874 242
rect 21894 222 21902 242
rect 21841 221 21902 222
rect 21758 214 21902 221
rect 21758 213 21794 214
rect 21866 213 21902 214
rect 21968 247 22005 248
rect 21968 246 22006 247
rect 21968 238 22032 246
rect 21968 218 21977 238
rect 21997 224 22032 238
rect 22052 224 22055 244
rect 21997 219 22055 224
rect 21997 218 22032 219
rect 21234 181 21271 210
rect 21235 179 21271 181
rect 21447 179 21484 210
rect 21235 157 21484 179
rect 21316 151 21427 157
rect 21316 143 21357 151
rect 21316 123 21324 143
rect 21343 123 21357 143
rect 21316 121 21357 123
rect 21385 143 21427 151
rect 21385 123 21401 143
rect 21420 123 21427 143
rect 21385 121 21427 123
rect 21316 106 21427 121
rect 21655 89 21692 210
rect 21968 206 22032 218
rect 22072 95 22099 358
rect 31836 331 31965 338
rect 31836 272 31860 331
rect 31891 272 31922 331
rect 31953 316 31965 331
rect 32427 316 32458 369
rect 32488 398 32525 477
rect 32640 408 32671 409
rect 32488 378 32497 398
rect 32517 378 32525 398
rect 32488 368 32525 378
rect 32584 401 32671 408
rect 32584 398 32645 401
rect 32584 378 32593 398
rect 32613 381 32645 398
rect 32666 381 32671 401
rect 32613 378 32671 381
rect 32584 371 32671 378
rect 32696 398 32733 528
rect 32848 408 32884 409
rect 32696 378 32705 398
rect 32725 378 32733 398
rect 32584 369 32640 371
rect 32584 368 32621 369
rect 32696 368 32733 378
rect 32792 398 32940 408
rect 33040 405 33136 407
rect 32792 378 32801 398
rect 32821 378 32911 398
rect 32931 378 32940 398
rect 32792 372 32940 378
rect 32792 369 32856 372
rect 32792 368 32829 369
rect 32848 342 32856 369
rect 32877 369 32940 372
rect 32998 398 33136 405
rect 32998 378 33007 398
rect 33027 378 33136 398
rect 32998 369 33136 378
rect 32877 342 32884 369
rect 32903 368 32940 369
rect 32999 368 33036 369
rect 32848 317 32884 342
rect 31953 315 32250 316
rect 32319 315 32360 316
rect 31953 308 32360 315
rect 31953 288 32329 308
rect 32349 288 32360 308
rect 31953 280 32360 288
rect 32427 312 32786 316
rect 32427 307 32749 312
rect 32427 283 32540 307
rect 32564 288 32749 307
rect 32773 288 32786 312
rect 32564 283 32786 288
rect 32427 280 32786 283
rect 32848 280 32883 317
rect 32951 314 33051 317
rect 32951 310 33018 314
rect 32951 284 32963 310
rect 32989 288 33018 310
rect 33044 288 33051 314
rect 32989 284 33051 288
rect 32951 280 33051 284
rect 31953 272 32250 280
rect 31836 259 31965 272
rect 32427 259 32458 280
rect 32848 259 32884 280
rect 32270 258 32307 259
rect 32269 249 32307 258
rect 32269 229 32278 249
rect 32298 229 32307 249
rect 32269 221 32307 229
rect 32373 253 32458 259
rect 32483 258 32520 259
rect 32373 233 32381 253
rect 32401 233 32458 253
rect 32373 225 32458 233
rect 32482 249 32520 258
rect 32482 229 32491 249
rect 32511 229 32520 249
rect 32373 224 32409 225
rect 32482 221 32520 229
rect 32586 253 32671 259
rect 32691 258 32728 259
rect 32586 233 32594 253
rect 32614 252 32671 253
rect 32614 233 32643 252
rect 32586 232 32643 233
rect 32664 232 32671 252
rect 32586 225 32671 232
rect 32690 249 32728 258
rect 32690 229 32699 249
rect 32719 229 32728 249
rect 32586 224 32622 225
rect 32690 221 32728 229
rect 32794 253 32938 259
rect 32794 233 32802 253
rect 32822 233 32857 253
rect 32794 230 32857 233
rect 32877 233 32910 253
rect 32930 233 32938 253
rect 32877 230 32938 233
rect 32794 225 32938 230
rect 32794 224 32830 225
rect 32902 224 32938 225
rect 33004 258 33041 259
rect 33004 257 33042 258
rect 33004 249 33068 257
rect 33004 229 33013 249
rect 33033 235 33068 249
rect 33088 235 33091 255
rect 33033 230 33091 235
rect 33033 229 33068 230
rect 32270 192 32307 221
rect 32271 190 32307 192
rect 32483 190 32520 221
rect 32271 168 32520 190
rect 32352 162 32463 168
rect 32352 154 32393 162
rect 32352 134 32360 154
rect 32379 134 32393 154
rect 32352 132 32393 134
rect 32421 154 32463 162
rect 32421 134 32437 154
rect 32456 134 32463 154
rect 32421 132 32463 134
rect 32352 117 32463 132
rect 32691 100 32728 221
rect 33004 217 33068 229
rect 33108 107 33135 369
rect 33333 107 33381 629
rect 33086 102 33381 107
rect 32967 100 33381 102
rect 22059 91 22117 95
rect 21931 89 22117 91
rect 21655 71 22117 89
rect 32691 74 33381 100
rect 32967 73 33381 74
rect 33086 72 33381 73
rect 21655 63 22076 71
rect 21931 62 22076 63
rect 22059 13 22076 62
rect 22105 13 22117 71
rect 33333 67 33381 72
rect 22059 -9 22117 13
rect 10160 -224 11940 -137
rect 11349 -227 11940 -224
<< viali >>
rect 2943 14408 2980 14456
rect 1473 13867 1498 13902
rect 1517 13867 1542 13905
rect 1706 13808 1726 13828
rect 2523 13868 2548 13903
rect 2567 13868 2592 13906
rect 2754 13804 2774 13824
rect 974 13741 1003 13768
rect 1048 13744 1077 13771
rect 779 13580 828 13622
rect 1262 13643 1283 13663
rect 2022 13737 2051 13764
rect 2096 13740 2125 13767
rect 1473 13604 1494 13634
rect 780 13517 829 13559
rect 1635 13550 1661 13576
rect 1260 13494 1281 13514
rect 1685 13497 1705 13517
rect 977 13396 996 13416
rect 1054 13396 1073 13416
rect 790 13290 830 13323
rect 1819 13574 1872 13607
rect 2310 13639 2331 13659
rect 2521 13600 2542 13630
rect 1824 13516 1877 13549
rect 2683 13546 2709 13572
rect 2308 13490 2329 13510
rect 2733 13493 2753 13513
rect 2025 13392 2044 13412
rect 2102 13392 2121 13412
rect 1841 13253 1886 13292
rect 2944 13553 2978 13592
rect 1468 13178 1493 13198
rect 1516 13179 1548 13199
rect 1706 13129 1726 13149
rect 974 13062 1003 13089
rect 1048 13065 1077 13092
rect 776 12869 816 12906
rect 1262 12964 1283 12984
rect 3121 13573 3157 13614
rect 3110 13233 3170 13277
rect 4916 13680 5002 13747
rect 8957 13606 8997 13632
rect 8960 13561 9000 13587
rect 4201 13124 4221 13144
rect 3469 13057 3498 13084
rect 3543 13060 3572 13087
rect 1473 12925 1494 12955
rect 1635 12871 1661 12897
rect 780 12829 816 12850
rect 1260 12815 1281 12835
rect 1685 12818 1705 12838
rect 977 12717 996 12737
rect 1054 12717 1073 12737
rect 772 12617 809 12658
rect 828 12619 865 12660
rect 1831 12916 1871 12942
rect 1835 12863 1875 12889
rect 1838 12818 1878 12844
rect 3757 12959 3778 12979
rect 3968 12920 3989 12950
rect 3110 12819 3164 12860
rect 4130 12866 4156 12892
rect 3755 12810 3776 12830
rect 1837 12493 1867 12559
rect 1473 12420 1498 12455
rect 1517 12420 1542 12458
rect 1706 12361 1726 12381
rect 2754 12357 2774 12377
rect 974 12294 1003 12321
rect 1048 12297 1077 12324
rect 779 12133 828 12175
rect 1262 12196 1283 12216
rect 2022 12290 2051 12317
rect 2096 12293 2125 12320
rect 1473 12157 1494 12187
rect 780 12070 829 12112
rect 1635 12103 1661 12129
rect 1260 12047 1281 12067
rect 1685 12050 1705 12070
rect 977 11949 996 11969
rect 1054 11949 1073 11969
rect 790 11843 830 11876
rect 1819 12127 1872 12160
rect 2310 12192 2331 12212
rect 2521 12153 2542 12183
rect 1824 12069 1877 12102
rect 2683 12099 2709 12125
rect 2308 12043 2329 12063
rect 2733 12046 2753 12066
rect 2025 11945 2044 11965
rect 2102 11945 2121 11965
rect 1841 11806 1886 11845
rect 3472 12712 3491 12732
rect 3549 12712 3568 12732
rect 4180 12813 4200 12833
rect 3979 12622 4031 12640
rect 3748 12421 3773 12456
rect 3792 12421 3817 12459
rect 4011 12437 4035 12460
rect 4011 12393 4035 12416
rect 1468 11731 1493 11751
rect 1516 11732 1548 11752
rect 1706 11682 1726 11702
rect 974 11615 1003 11642
rect 1048 11618 1077 11645
rect 776 11422 816 11459
rect 1262 11517 1283 11537
rect 1473 11478 1494 11508
rect 1635 11424 1661 11450
rect 780 11382 816 11403
rect 1260 11368 1281 11388
rect 1685 11371 1705 11391
rect 977 11270 996 11290
rect 1054 11270 1073 11290
rect 772 11170 809 11211
rect 828 11172 865 11213
rect 1831 11469 1871 11495
rect 1835 11416 1875 11442
rect 1838 11371 1878 11397
rect 1830 11111 1874 11148
rect 4016 11774 4036 11795
rect 4057 11779 4077 11800
rect 4244 11679 4264 11699
rect 3512 11612 3541 11639
rect 3586 11615 3615 11642
rect 3800 11514 3821 11534
rect 4011 11475 4032 11505
rect 4173 11421 4199 11447
rect 1825 11025 1879 11091
rect 1474 10900 1499 10935
rect 1518 10900 1543 10938
rect 1707 10841 1727 10861
rect 2755 10837 2775 10857
rect 975 10774 1004 10801
rect 1049 10777 1078 10804
rect 780 10613 829 10655
rect 1263 10676 1284 10696
rect 2023 10770 2052 10797
rect 2097 10773 2126 10800
rect 1474 10637 1495 10667
rect 781 10550 830 10592
rect 1636 10583 1662 10609
rect 1261 10527 1282 10547
rect 1686 10530 1706 10550
rect 978 10429 997 10449
rect 1055 10429 1074 10449
rect 791 10323 831 10356
rect 1820 10607 1873 10640
rect 2311 10672 2332 10692
rect 2522 10633 2543 10663
rect 1825 10549 1878 10582
rect 2684 10579 2710 10605
rect 2309 10523 2330 10543
rect 2734 10526 2754 10546
rect 2026 10425 2045 10445
rect 2103 10425 2122 10445
rect 1842 10286 1887 10325
rect 1469 10211 1494 10231
rect 1517 10212 1549 10232
rect 1707 10162 1727 10182
rect 975 10095 1004 10122
rect 1049 10098 1078 10125
rect 777 9902 817 9939
rect 1263 9997 1284 10017
rect 1474 9958 1495 9988
rect 1636 9904 1662 9930
rect 781 9862 817 9883
rect 1261 9848 1282 9868
rect 1686 9851 1706 9871
rect 978 9750 997 9770
rect 1055 9750 1074 9770
rect 773 9650 810 9691
rect 829 9652 866 9693
rect 1832 9949 1872 9975
rect 1836 9896 1876 9922
rect 1839 9851 1879 9877
rect 2946 9892 2972 9915
rect 1838 9526 1868 9592
rect 1474 9453 1499 9488
rect 1518 9453 1543 9491
rect 1707 9394 1727 9414
rect 2755 9390 2775 9410
rect 975 9327 1004 9354
rect 1049 9330 1078 9357
rect 780 9166 829 9208
rect 1263 9229 1284 9249
rect 2023 9323 2052 9350
rect 2097 9326 2126 9353
rect 1474 9190 1495 9220
rect 781 9103 830 9145
rect 1636 9136 1662 9162
rect 1261 9080 1282 9100
rect 1686 9083 1706 9103
rect 978 8982 997 9002
rect 1055 8982 1074 9002
rect 791 8876 831 8909
rect 1820 9160 1873 9193
rect 2311 9225 2332 9245
rect 2522 9186 2543 9216
rect 1825 9102 1878 9135
rect 2684 9132 2710 9158
rect 2309 9076 2330 9096
rect 2734 9079 2754 9099
rect 2026 8978 2045 8998
rect 2103 8978 2122 8998
rect 1842 8839 1887 8878
rect 1469 8764 1494 8784
rect 1517 8765 1549 8785
rect 1707 8715 1727 8735
rect 975 8648 1004 8675
rect 1049 8651 1078 8678
rect 777 8455 817 8492
rect 1263 8550 1284 8570
rect 1474 8511 1495 8541
rect 1636 8457 1662 8483
rect 781 8415 817 8436
rect 1261 8401 1282 8421
rect 1686 8404 1706 8424
rect 978 8303 997 8323
rect 1055 8303 1074 8323
rect 773 8203 810 8244
rect 829 8205 866 8246
rect 1832 8502 1872 8528
rect 1836 8449 1876 8475
rect 1839 8404 1879 8430
rect 1830 8083 1876 8131
rect 3798 11365 3819 11385
rect 4223 11368 4243 11388
rect 3515 11267 3534 11287
rect 3592 11267 3611 11287
rect 3815 10901 3840 10939
rect 3973 10210 3990 10247
rect 4202 10157 4222 10177
rect 3470 10090 3499 10117
rect 3544 10093 3573 10120
rect 3758 9992 3779 10012
rect 3969 9953 3990 9983
rect 3326 9885 3352 9908
rect 4131 9899 4157 9925
rect 3756 9843 3777 9863
rect 4181 9846 4201 9866
rect 3473 9745 3492 9765
rect 3550 9745 3569 9765
rect 3813 9473 3841 9501
rect 5310 8706 5330 8726
rect 4578 8639 4607 8666
rect 4652 8642 4681 8669
rect 4866 8541 4887 8561
rect 5077 8502 5098 8532
rect 4374 8443 4398 8467
rect 4431 8444 4455 8468
rect 5239 8448 5265 8474
rect 4864 8392 4885 8412
rect 5077 8390 5101 8412
rect 5289 8395 5309 8415
rect 4581 8294 4600 8314
rect 4658 8294 4677 8314
rect 8964 13508 9004 13534
rect 9970 13790 10007 13831
rect 10026 13792 10063 13833
rect 9762 13713 9781 13733
rect 9839 13713 9858 13733
rect 9130 13612 9150 13632
rect 9554 13615 9575 13635
rect 12181 13861 12206 13896
rect 12225 13861 12250 13899
rect 12414 13802 12434 13822
rect 13231 13862 13256 13897
rect 13275 13862 13300 13900
rect 10019 13600 10055 13621
rect 13462 13798 13482 13818
rect 11682 13735 11711 13762
rect 11756 13738 11785 13765
rect 9174 13553 9200 13579
rect 9341 13495 9362 13525
rect 9552 13466 9573 13486
rect 10019 13544 10059 13581
rect 11487 13574 11536 13616
rect 11970 13637 11991 13657
rect 12730 13731 12759 13758
rect 12804 13734 12833 13761
rect 12181 13598 12202 13628
rect 11488 13511 11537 13553
rect 12343 13544 12369 13570
rect 9758 13358 9787 13385
rect 9832 13361 9861 13388
rect 9109 13301 9129 13321
rect 9287 13251 9319 13271
rect 9342 13252 9367 13272
rect 8949 13158 8994 13197
rect 8714 13038 8733 13058
rect 8791 13038 8810 13058
rect 8082 12937 8102 12957
rect 8506 12940 8527 12960
rect 8126 12878 8152 12904
rect 8958 12901 9011 12934
rect 8293 12820 8314 12850
rect 8504 12791 8525 12811
rect 8963 12843 9016 12876
rect 10005 13127 10045 13160
rect 9762 13034 9781 13054
rect 9839 13034 9858 13054
rect 9130 12933 9150 12953
rect 9554 12936 9575 12956
rect 11968 13488 11989 13508
rect 12393 13491 12413 13511
rect 11685 13390 11704 13410
rect 11762 13390 11781 13410
rect 11498 13284 11538 13317
rect 12527 13568 12580 13601
rect 13018 13633 13039 13653
rect 13229 13594 13250 13624
rect 12532 13510 12585 13543
rect 13391 13540 13417 13566
rect 13016 13484 13037 13504
rect 13441 13487 13461 13507
rect 12733 13386 12752 13406
rect 12810 13386 12829 13406
rect 12549 13247 12594 13286
rect 13652 13547 13686 13586
rect 12176 13172 12201 13192
rect 12224 13173 12256 13193
rect 12414 13123 12434 13143
rect 11682 13056 11711 13083
rect 11756 13059 11785 13086
rect 9174 12874 9200 12900
rect 10006 12891 10055 12933
rect 9341 12816 9362 12846
rect 8710 12683 8739 12710
rect 8784 12686 8813 12713
rect 9552 12787 9573 12807
rect 10007 12828 10056 12870
rect 11484 12863 11524 12900
rect 11970 12958 11991 12978
rect 13829 13567 13865 13608
rect 13818 13227 13878 13271
rect 15130 13669 15168 13766
rect 15190 13675 15228 13772
rect 19665 13600 19705 13626
rect 14909 13118 14929 13138
rect 14177 13051 14206 13078
rect 14251 13054 14280 13081
rect 12181 12919 12202 12949
rect 12343 12865 12369 12891
rect 9758 12679 9787 12706
rect 9832 12682 9861 12709
rect 8061 12626 8081 12646
rect 11488 12823 11524 12844
rect 9109 12622 9129 12642
rect 6995 12535 7023 12563
rect 9293 12545 9318 12583
rect 9337 12548 9362 12583
rect 11968 12809 11989 12829
rect 12393 12812 12413 12832
rect 11685 12711 11704 12731
rect 11762 12711 11781 12731
rect 11480 12611 11517 12652
rect 11536 12613 11573 12654
rect 12539 12910 12579 12936
rect 12543 12857 12583 12883
rect 12546 12812 12586 12838
rect 8968 12444 8998 12510
rect 7267 12271 7286 12291
rect 7344 12271 7363 12291
rect 14465 12953 14486 12973
rect 14676 12914 14697 12944
rect 13818 12813 13872 12854
rect 14838 12860 14864 12886
rect 14463 12804 14484 12824
rect 12545 12487 12575 12553
rect 6635 12170 6655 12190
rect 7059 12173 7080 12193
rect 6679 12111 6705 12137
rect 7484 12128 7510 12151
rect 7864 12121 7890 12144
rect 6846 12053 6867 12083
rect 7057 12024 7078 12044
rect 8957 12159 8997 12185
rect 8960 12114 9000 12140
rect 8964 12061 9004 12087
rect 7263 11916 7292 11943
rect 7337 11919 7366 11946
rect 6614 11859 6634 11879
rect 6846 11789 6863 11826
rect 9970 12343 10007 12384
rect 10026 12345 10063 12386
rect 9762 12266 9781 12286
rect 9839 12266 9858 12286
rect 9130 12165 9150 12185
rect 9554 12168 9575 12188
rect 12181 12414 12206 12449
rect 12225 12414 12250 12452
rect 12414 12355 12434 12375
rect 10019 12153 10055 12174
rect 13462 12351 13482 12371
rect 11682 12288 11711 12315
rect 11756 12291 11785 12318
rect 9174 12106 9200 12132
rect 9341 12048 9362 12078
rect 9552 12019 9573 12039
rect 10019 12097 10059 12134
rect 11487 12127 11536 12169
rect 11970 12190 11991 12210
rect 12730 12284 12759 12311
rect 12804 12287 12833 12314
rect 12181 12151 12202 12181
rect 11488 12064 11537 12106
rect 12343 12097 12369 12123
rect 9758 11911 9787 11938
rect 9832 11914 9861 11941
rect 9109 11854 9129 11874
rect 9287 11804 9319 11824
rect 9342 11805 9367 11825
rect 6996 11097 7021 11135
rect 8949 11711 8994 11750
rect 8714 11591 8733 11611
rect 8791 11591 8810 11611
rect 8082 11490 8102 11510
rect 8506 11493 8527 11513
rect 8126 11431 8152 11457
rect 8958 11454 9011 11487
rect 8293 11373 8314 11403
rect 8504 11344 8525 11364
rect 8963 11396 9016 11429
rect 10005 11680 10045 11713
rect 9762 11587 9781 11607
rect 9839 11587 9858 11607
rect 9130 11486 9150 11506
rect 9554 11489 9575 11509
rect 11968 12041 11989 12061
rect 12393 12044 12413 12064
rect 11685 11943 11704 11963
rect 11762 11943 11781 11963
rect 11498 11837 11538 11870
rect 12527 12121 12580 12154
rect 13018 12186 13039 12206
rect 13229 12147 13250 12177
rect 12532 12063 12585 12096
rect 13391 12093 13417 12119
rect 13016 12037 13037 12057
rect 13441 12040 13461 12060
rect 12733 11939 12752 11959
rect 12810 11939 12829 11959
rect 12549 11800 12594 11839
rect 14180 12706 14199 12726
rect 14257 12706 14276 12726
rect 14888 12807 14908 12827
rect 14687 12616 14739 12634
rect 14456 12415 14481 12450
rect 14500 12415 14525 12453
rect 14719 12431 14743 12454
rect 14719 12387 14743 12410
rect 12176 11725 12201 11745
rect 12224 11726 12256 11746
rect 12414 11676 12434 11696
rect 11682 11609 11711 11636
rect 11756 11612 11785 11639
rect 9174 11427 9200 11453
rect 10006 11444 10055 11486
rect 9341 11369 9362 11399
rect 8710 11236 8739 11263
rect 8784 11239 8813 11266
rect 9552 11340 9573 11360
rect 10007 11381 10056 11423
rect 11484 11416 11524 11453
rect 11970 11511 11991 11531
rect 12181 11472 12202 11502
rect 12343 11418 12369 11444
rect 9758 11232 9787 11259
rect 9832 11235 9861 11262
rect 8061 11179 8081 11199
rect 11488 11376 11524 11397
rect 9109 11175 9129 11195
rect 9293 11098 9318 11136
rect 9337 11101 9362 11136
rect 11968 11362 11989 11382
rect 12393 11365 12413 11385
rect 11685 11264 11704 11284
rect 11762 11264 11781 11284
rect 11480 11164 11517 11205
rect 11536 11166 11573 11207
rect 12539 11463 12579 11489
rect 12543 11410 12583 11436
rect 12546 11365 12586 11391
rect 12538 11105 12582 11142
rect 14724 11768 14744 11789
rect 14765 11773 14785 11794
rect 14952 11673 14972 11693
rect 14220 11606 14249 11633
rect 14294 11609 14323 11636
rect 14508 11508 14529 11528
rect 14719 11469 14740 11499
rect 14881 11415 14907 11441
rect 8957 10945 9011 11011
rect 12533 11019 12587 11085
rect 7225 10749 7244 10769
rect 7302 10749 7321 10769
rect 6593 10648 6613 10668
rect 7017 10651 7038 10671
rect 6637 10589 6663 10615
rect 6804 10531 6825 10561
rect 7015 10502 7036 10522
rect 7221 10394 7250 10421
rect 7295 10397 7324 10424
rect 6572 10337 6592 10357
rect 8962 10888 9006 10925
rect 8958 10639 8998 10665
rect 8961 10594 9001 10620
rect 8965 10541 9005 10567
rect 9971 10823 10008 10864
rect 10027 10825 10064 10866
rect 9763 10746 9782 10766
rect 9840 10746 9859 10766
rect 9131 10645 9151 10665
rect 9555 10648 9576 10668
rect 12182 10894 12207 10929
rect 12226 10894 12251 10932
rect 12415 10835 12435 10855
rect 10020 10633 10056 10654
rect 13463 10831 13483 10851
rect 11683 10768 11712 10795
rect 11757 10771 11786 10798
rect 9175 10586 9201 10612
rect 9342 10528 9363 10558
rect 9553 10499 9574 10519
rect 10020 10577 10060 10614
rect 11488 10607 11537 10649
rect 11971 10670 11992 10690
rect 12731 10764 12760 10791
rect 12805 10767 12834 10794
rect 12182 10631 12203 10661
rect 11489 10544 11538 10586
rect 12344 10577 12370 10603
rect 9759 10391 9788 10418
rect 9833 10394 9862 10421
rect 9110 10334 9130 10354
rect 9288 10284 9320 10304
rect 9343 10285 9368 10305
rect 6801 9620 6825 9643
rect 6801 9576 6825 9599
rect 7019 9577 7044 9615
rect 7063 9580 7088 9615
rect 6805 9396 6857 9414
rect 6636 9203 6656 9223
rect 7268 9304 7287 9324
rect 7345 9304 7364 9324
rect 8950 10191 8995 10230
rect 8715 10071 8734 10091
rect 8792 10071 8811 10091
rect 8083 9970 8103 9990
rect 8507 9973 8528 9993
rect 8127 9911 8153 9937
rect 8959 9934 9012 9967
rect 8294 9853 8315 9883
rect 8505 9824 8526 9844
rect 8964 9876 9017 9909
rect 10006 10160 10046 10193
rect 9763 10067 9782 10087
rect 9840 10067 9859 10087
rect 9131 9966 9151 9986
rect 9555 9969 9576 9989
rect 11969 10521 11990 10541
rect 12394 10524 12414 10544
rect 11686 10423 11705 10443
rect 11763 10423 11782 10443
rect 11499 10317 11539 10350
rect 12528 10601 12581 10634
rect 13019 10666 13040 10686
rect 13230 10627 13251 10657
rect 12533 10543 12586 10576
rect 13392 10573 13418 10599
rect 13017 10517 13038 10537
rect 13442 10520 13462 10540
rect 12734 10419 12753 10439
rect 12811 10419 12830 10439
rect 12550 10280 12595 10319
rect 12177 10205 12202 10225
rect 12225 10206 12257 10226
rect 12415 10156 12435 10176
rect 11683 10089 11712 10116
rect 11757 10092 11786 10119
rect 9175 9907 9201 9933
rect 10007 9924 10056 9966
rect 9342 9849 9363 9879
rect 8711 9716 8740 9743
rect 8785 9719 8814 9746
rect 9553 9820 9574 9840
rect 10008 9861 10057 9903
rect 11485 9896 11525 9933
rect 11971 9991 11992 10011
rect 12182 9952 12203 9982
rect 12344 9898 12370 9924
rect 9759 9712 9788 9739
rect 9833 9715 9862 9742
rect 8062 9659 8082 9679
rect 11489 9856 11525 9877
rect 9110 9655 9130 9675
rect 9294 9578 9319 9616
rect 9338 9581 9363 9616
rect 11969 9842 11990 9862
rect 12394 9845 12414 9865
rect 11686 9744 11705 9764
rect 11763 9744 11782 9764
rect 11481 9644 11518 9685
rect 11537 9646 11574 9687
rect 12540 9943 12580 9969
rect 12544 9890 12584 9916
rect 12547 9845 12587 9871
rect 13654 9886 13680 9909
rect 8969 9477 8999 9543
rect 7060 9206 7081 9226
rect 6680 9144 6706 9170
rect 7672 9176 7726 9217
rect 6847 9086 6868 9116
rect 7058 9057 7079 9077
rect 12546 9520 12576 9586
rect 8958 9192 8998 9218
rect 8961 9147 9001 9173
rect 8965 9094 9005 9120
rect 9971 9376 10008 9417
rect 10027 9378 10064 9419
rect 9763 9299 9782 9319
rect 9840 9299 9859 9319
rect 9131 9198 9151 9218
rect 9555 9201 9576 9221
rect 12182 9447 12207 9482
rect 12226 9447 12251 9485
rect 12415 9388 12435 9408
rect 10020 9186 10056 9207
rect 13463 9384 13483 9404
rect 11683 9321 11712 9348
rect 11757 9324 11786 9351
rect 9175 9139 9201 9165
rect 9342 9081 9363 9111
rect 7264 8949 7293 8976
rect 7338 8952 7367 8979
rect 6615 8892 6635 8912
rect 4917 8201 4946 8235
rect 4916 8141 4945 8175
rect 3132 8056 3176 8084
rect 2941 7957 2978 8005
rect 3129 7999 3173 8027
rect 5424 7917 5487 7971
rect 1471 7859 1496 7894
rect 1515 7859 1540 7897
rect 1704 7800 1724 7820
rect 2521 7860 2546 7895
rect 2565 7860 2590 7898
rect 2752 7796 2772 7816
rect 972 7733 1001 7760
rect 1046 7736 1075 7763
rect 777 7572 826 7614
rect 1260 7635 1281 7655
rect 2020 7729 2049 7756
rect 2094 7732 2123 7759
rect 1471 7596 1492 7626
rect 778 7509 827 7551
rect 1633 7542 1659 7568
rect 1258 7486 1279 7506
rect 1683 7489 1703 7509
rect 975 7388 994 7408
rect 1052 7388 1071 7408
rect 788 7282 828 7315
rect 1817 7566 1870 7599
rect 2308 7631 2329 7651
rect 2519 7592 2540 7622
rect 1822 7508 1875 7541
rect 2681 7538 2707 7564
rect 2306 7482 2327 7502
rect 2731 7485 2751 7505
rect 2023 7384 2042 7404
rect 2100 7384 2119 7404
rect 1839 7245 1884 7284
rect 2942 7545 2976 7584
rect 1466 7170 1491 7190
rect 1514 7171 1546 7191
rect 1704 7121 1724 7141
rect 972 7054 1001 7081
rect 1046 7057 1075 7084
rect 774 6861 814 6898
rect 1260 6956 1281 6976
rect 3119 7565 3155 7606
rect 3108 7225 3168 7269
rect 4199 7116 4219 7136
rect 3467 7049 3496 7076
rect 3541 7052 3570 7079
rect 1471 6917 1492 6947
rect 1633 6863 1659 6889
rect 778 6821 814 6842
rect 1258 6807 1279 6827
rect 1683 6810 1703 6830
rect 975 6709 994 6729
rect 1052 6709 1071 6729
rect 770 6609 807 6650
rect 826 6611 863 6652
rect 1829 6908 1869 6934
rect 1833 6855 1873 6881
rect 1836 6810 1876 6836
rect 3755 6951 3776 6971
rect 3966 6912 3987 6942
rect 3108 6811 3162 6852
rect 4128 6858 4154 6884
rect 3753 6802 3774 6822
rect 1835 6485 1865 6551
rect 1471 6412 1496 6447
rect 1515 6412 1540 6450
rect 1704 6353 1724 6373
rect 2752 6349 2772 6369
rect 972 6286 1001 6313
rect 1046 6289 1075 6316
rect 777 6125 826 6167
rect 1260 6188 1281 6208
rect 2020 6282 2049 6309
rect 2094 6285 2123 6312
rect 1471 6149 1492 6179
rect 778 6062 827 6104
rect 1633 6095 1659 6121
rect 1258 6039 1279 6059
rect 1683 6042 1703 6062
rect 975 5941 994 5961
rect 1052 5941 1071 5961
rect 788 5835 828 5868
rect 1817 6119 1870 6152
rect 2308 6184 2329 6204
rect 2519 6145 2540 6175
rect 1822 6061 1875 6094
rect 2681 6091 2707 6117
rect 2306 6035 2327 6055
rect 2731 6038 2751 6058
rect 2023 5937 2042 5957
rect 2100 5937 2119 5957
rect 1839 5798 1884 5837
rect 3470 6704 3489 6724
rect 3547 6704 3566 6724
rect 4178 6805 4198 6825
rect 3977 6614 4029 6632
rect 3746 6413 3771 6448
rect 3790 6413 3815 6451
rect 4009 6429 4033 6452
rect 4009 6385 4033 6408
rect 1466 5723 1491 5743
rect 1514 5724 1546 5744
rect 1704 5674 1724 5694
rect 972 5607 1001 5634
rect 1046 5610 1075 5637
rect 774 5414 814 5451
rect 1260 5509 1281 5529
rect 1471 5470 1492 5500
rect 1633 5416 1659 5442
rect 778 5374 814 5395
rect 1258 5360 1279 5380
rect 1683 5363 1703 5383
rect 975 5262 994 5282
rect 1052 5262 1071 5282
rect 770 5162 807 5203
rect 826 5164 863 5205
rect 1829 5461 1869 5487
rect 1833 5408 1873 5434
rect 1836 5363 1876 5389
rect 1828 5103 1872 5140
rect 4242 5671 4262 5691
rect 3510 5604 3539 5631
rect 3584 5607 3613 5634
rect 3798 5506 3819 5526
rect 4009 5467 4030 5497
rect 4171 5413 4197 5439
rect 1823 5017 1877 5083
rect 1472 4892 1497 4927
rect 1516 4892 1541 4930
rect 1705 4833 1725 4853
rect 2753 4829 2773 4849
rect 973 4766 1002 4793
rect 1047 4769 1076 4796
rect 778 4605 827 4647
rect 1261 4668 1282 4688
rect 2021 4762 2050 4789
rect 2095 4765 2124 4792
rect 1472 4629 1493 4659
rect 779 4542 828 4584
rect 1634 4575 1660 4601
rect 1259 4519 1280 4539
rect 1684 4522 1704 4542
rect 976 4421 995 4441
rect 1053 4421 1072 4441
rect 789 4315 829 4348
rect 1818 4599 1871 4632
rect 2309 4664 2330 4684
rect 2520 4625 2541 4655
rect 1823 4541 1876 4574
rect 2682 4571 2708 4597
rect 2307 4515 2328 4535
rect 2732 4518 2752 4538
rect 2024 4417 2043 4437
rect 2101 4417 2120 4437
rect 1840 4278 1885 4317
rect 1467 4203 1492 4223
rect 1515 4204 1547 4224
rect 1705 4154 1725 4174
rect 973 4087 1002 4114
rect 1047 4090 1076 4117
rect 775 3894 815 3931
rect 1261 3989 1282 4009
rect 1472 3950 1493 3980
rect 1634 3896 1660 3922
rect 779 3854 815 3875
rect 1259 3840 1280 3860
rect 1684 3843 1704 3863
rect 976 3742 995 3762
rect 1053 3742 1072 3762
rect 771 3642 808 3683
rect 827 3644 864 3685
rect 1830 3941 1870 3967
rect 1834 3888 1874 3914
rect 1837 3843 1877 3869
rect 2899 3874 2924 3905
rect 2944 3884 2970 3907
rect 1836 3518 1866 3584
rect 1472 3445 1497 3480
rect 1516 3445 1541 3483
rect 1705 3386 1725 3406
rect 2753 3382 2773 3402
rect 973 3319 1002 3346
rect 1047 3322 1076 3349
rect 778 3158 827 3200
rect 1261 3221 1282 3241
rect 2021 3315 2050 3342
rect 2095 3318 2124 3345
rect 1472 3182 1493 3212
rect 779 3095 828 3137
rect 1634 3128 1660 3154
rect 1259 3072 1280 3092
rect 1684 3075 1704 3095
rect 976 2974 995 2994
rect 1053 2974 1072 2994
rect 789 2868 829 2901
rect 1818 3152 1871 3185
rect 2309 3217 2330 3237
rect 2520 3178 2541 3208
rect 1823 3094 1876 3127
rect 2682 3124 2708 3150
rect 2307 3068 2328 3088
rect 2732 3071 2752 3091
rect 2024 2970 2043 2990
rect 2101 2970 2120 2990
rect 1840 2831 1885 2870
rect 1467 2756 1492 2776
rect 1515 2757 1547 2777
rect 1705 2707 1725 2727
rect 973 2640 1002 2667
rect 1047 2643 1076 2670
rect 775 2447 815 2484
rect 1261 2542 1282 2562
rect 1472 2503 1493 2533
rect 1634 2449 1660 2475
rect 779 2407 815 2428
rect 1259 2393 1280 2413
rect 1684 2396 1704 2416
rect 976 2295 995 2315
rect 1053 2295 1072 2315
rect 771 2195 808 2236
rect 827 2197 864 2238
rect 3796 5357 3817 5377
rect 4221 5360 4241 5380
rect 3513 5259 3532 5279
rect 3590 5259 3609 5279
rect 3813 4893 3838 4931
rect 5889 7853 5918 7887
rect 5888 7793 5917 7827
rect 6157 7714 6176 7734
rect 6234 7714 6253 7734
rect 5525 7613 5545 7633
rect 5949 7616 5970 7636
rect 7666 8759 7726 8803
rect 7679 8422 7715 8463
rect 9553 9052 9574 9072
rect 10020 9130 10060 9167
rect 11488 9160 11537 9202
rect 11971 9223 11992 9243
rect 12731 9317 12760 9344
rect 12805 9320 12834 9347
rect 12182 9184 12203 9214
rect 11489 9097 11538 9139
rect 12344 9130 12370 9156
rect 9759 8944 9788 8971
rect 9833 8947 9862 8974
rect 9110 8887 9130 8907
rect 9288 8837 9320 8857
rect 9343 8838 9368 8858
rect 7858 8444 7892 8483
rect 8950 8744 8995 8783
rect 8715 8624 8734 8644
rect 8792 8624 8811 8644
rect 8083 8523 8103 8543
rect 8507 8526 8528 8546
rect 8127 8464 8153 8490
rect 8959 8487 9012 8520
rect 8294 8406 8315 8436
rect 8505 8377 8526 8397
rect 8964 8429 9017 8462
rect 10006 8713 10046 8746
rect 9763 8620 9782 8640
rect 9840 8620 9859 8640
rect 9131 8519 9151 8539
rect 9555 8522 9576 8542
rect 11969 9074 11990 9094
rect 12394 9077 12414 9097
rect 11686 8976 11705 8996
rect 11763 8976 11782 8996
rect 11499 8870 11539 8903
rect 12528 9154 12581 9187
rect 13019 9219 13040 9239
rect 13230 9180 13251 9210
rect 12533 9096 12586 9129
rect 13392 9126 13418 9152
rect 13017 9070 13038 9090
rect 13442 9073 13462 9093
rect 12734 8972 12753 8992
rect 12811 8972 12830 8992
rect 12550 8833 12595 8872
rect 12177 8758 12202 8778
rect 12225 8759 12257 8779
rect 12415 8709 12435 8729
rect 11683 8642 11712 8669
rect 11757 8645 11786 8672
rect 9175 8460 9201 8486
rect 10007 8477 10056 8519
rect 9342 8402 9363 8432
rect 8711 8269 8740 8296
rect 8785 8272 8814 8299
rect 9553 8373 9574 8393
rect 10008 8414 10057 8456
rect 11485 8449 11525 8486
rect 11971 8544 11992 8564
rect 12182 8505 12203 8535
rect 12344 8451 12370 8477
rect 9759 8265 9788 8292
rect 9833 8268 9862 8295
rect 8062 8212 8082 8232
rect 11489 8409 11525 8430
rect 8244 8130 8269 8168
rect 8288 8133 8313 8168
rect 9110 8208 9130 8228
rect 9294 8131 9319 8169
rect 9338 8134 9363 8169
rect 11969 8395 11990 8415
rect 12394 8398 12414 8418
rect 11686 8297 11705 8317
rect 11763 8297 11782 8317
rect 11481 8197 11518 8238
rect 11537 8199 11574 8240
rect 12540 8496 12580 8522
rect 12544 8443 12584 8469
rect 12547 8398 12587 8424
rect 5569 7554 5595 7580
rect 6379 7560 6403 7584
rect 6436 7561 6460 7585
rect 5736 7496 5757 7526
rect 5947 7467 5968 7487
rect 7661 8001 7705 8029
rect 7856 8023 7893 8071
rect 7658 7944 7702 7972
rect 6153 7359 6182 7386
rect 6227 7362 6256 7389
rect 5504 7302 5524 7322
rect 5266 4904 5291 4930
rect 5655 4835 5675 4855
rect 4923 4768 4952 4795
rect 4997 4771 5026 4798
rect 5211 4670 5232 4690
rect 5422 4631 5443 4661
rect 5584 4577 5610 4603
rect 5209 4521 5230 4541
rect 5413 4523 5446 4543
rect 5634 4524 5654 4544
rect 4926 4423 4945 4443
rect 5003 4423 5022 4443
rect 5734 4366 5757 4404
rect 6993 6527 7021 6555
rect 7265 6263 7284 6283
rect 7342 6263 7361 6283
rect 6633 6162 6653 6182
rect 7057 6165 7078 6185
rect 6677 6103 6703 6129
rect 7482 6120 7508 6143
rect 6844 6045 6865 6075
rect 7055 6016 7076 6036
rect 7261 5908 7290 5935
rect 7335 5911 7364 5938
rect 6612 5851 6632 5871
rect 6844 5781 6861 5818
rect 6994 5089 7019 5127
rect 7223 4741 7242 4761
rect 7300 4741 7319 4761
rect 6591 4640 6611 4660
rect 7015 4643 7036 4663
rect 8958 7897 9004 7945
rect 12538 8077 12584 8125
rect 14506 11359 14527 11379
rect 14931 11362 14951 11382
rect 14223 11261 14242 11281
rect 14300 11261 14319 11281
rect 14523 10895 14548 10933
rect 14681 10204 14698 10241
rect 14910 10151 14930 10171
rect 14178 10084 14207 10111
rect 14252 10087 14281 10114
rect 14466 9986 14487 10006
rect 14677 9947 14698 9977
rect 14034 9879 14060 9902
rect 14839 9893 14865 9919
rect 14464 9837 14485 9857
rect 14889 9840 14909 9860
rect 14181 9739 14200 9759
rect 14258 9739 14277 9759
rect 14521 9467 14549 9495
rect 16018 8700 16038 8720
rect 15286 8633 15315 8660
rect 15360 8636 15389 8663
rect 15574 8535 15595 8555
rect 15785 8496 15806 8526
rect 15082 8437 15106 8461
rect 15139 8438 15163 8462
rect 15947 8442 15973 8468
rect 15572 8386 15593 8406
rect 15785 8384 15809 8406
rect 15997 8389 16017 8409
rect 15289 8288 15308 8308
rect 15366 8288 15385 8308
rect 19668 13555 19708 13581
rect 19672 13502 19712 13528
rect 23146 13865 23171 13900
rect 23190 13865 23215 13903
rect 20678 13784 20715 13825
rect 20734 13786 20771 13827
rect 20470 13707 20489 13727
rect 20547 13707 20566 13727
rect 19838 13606 19858 13626
rect 20262 13609 20283 13629
rect 23379 13806 23399 13826
rect 24196 13866 24221 13901
rect 24240 13866 24265 13904
rect 24427 13802 24447 13822
rect 20727 13594 20763 13615
rect 22647 13739 22676 13766
rect 22721 13742 22750 13769
rect 19882 13547 19908 13573
rect 20049 13489 20070 13519
rect 20260 13460 20281 13480
rect 20727 13538 20767 13575
rect 22452 13578 22501 13620
rect 22935 13641 22956 13661
rect 23695 13735 23724 13762
rect 23769 13738 23798 13765
rect 23146 13602 23167 13632
rect 22453 13515 22502 13557
rect 23308 13548 23334 13574
rect 20466 13352 20495 13379
rect 20540 13355 20569 13382
rect 19817 13295 19837 13315
rect 19995 13245 20027 13265
rect 20050 13246 20075 13266
rect 19657 13152 19702 13191
rect 19422 13032 19441 13052
rect 19499 13032 19518 13052
rect 18790 12931 18810 12951
rect 19214 12934 19235 12954
rect 18834 12872 18860 12898
rect 19666 12895 19719 12928
rect 19001 12814 19022 12844
rect 19212 12785 19233 12805
rect 19671 12837 19724 12870
rect 20713 13121 20753 13154
rect 20470 13028 20489 13048
rect 20547 13028 20566 13048
rect 19838 12927 19858 12947
rect 20262 12930 20283 12950
rect 22933 13492 22954 13512
rect 23358 13495 23378 13515
rect 22650 13394 22669 13414
rect 22727 13394 22746 13414
rect 22463 13288 22503 13321
rect 23492 13572 23545 13605
rect 23983 13637 24004 13657
rect 24194 13598 24215 13628
rect 23497 13514 23550 13547
rect 24356 13544 24382 13570
rect 23981 13488 24002 13508
rect 24406 13491 24426 13511
rect 23698 13390 23717 13410
rect 23775 13390 23794 13410
rect 23514 13251 23559 13290
rect 24617 13551 24651 13590
rect 23141 13176 23166 13196
rect 23189 13177 23221 13197
rect 23379 13127 23399 13147
rect 22647 13060 22676 13087
rect 22721 13063 22750 13090
rect 19882 12868 19908 12894
rect 20714 12885 20763 12927
rect 20049 12810 20070 12840
rect 19418 12677 19447 12704
rect 19492 12680 19521 12707
rect 20260 12781 20281 12801
rect 20715 12822 20764 12864
rect 22449 12867 22489 12904
rect 22935 12962 22956 12982
rect 24794 13571 24830 13612
rect 24783 13231 24843 13275
rect 26589 13678 26675 13745
rect 30630 13604 30670 13630
rect 30633 13559 30673 13585
rect 25874 13122 25894 13142
rect 25142 13055 25171 13082
rect 25216 13058 25245 13085
rect 23146 12923 23167 12953
rect 23308 12869 23334 12895
rect 20466 12673 20495 12700
rect 20540 12676 20569 12703
rect 22453 12827 22489 12848
rect 18769 12620 18789 12640
rect 19817 12616 19837 12636
rect 17703 12529 17731 12557
rect 20001 12539 20026 12577
rect 20045 12542 20070 12577
rect 22933 12813 22954 12833
rect 23358 12816 23378 12836
rect 22650 12715 22669 12735
rect 22727 12715 22746 12735
rect 22445 12615 22482 12656
rect 22501 12617 22538 12658
rect 23504 12914 23544 12940
rect 23508 12861 23548 12887
rect 23511 12816 23551 12842
rect 19676 12438 19706 12504
rect 17975 12265 17994 12285
rect 18052 12265 18071 12285
rect 25430 12957 25451 12977
rect 25641 12918 25662 12948
rect 24783 12817 24837 12858
rect 25803 12864 25829 12890
rect 25428 12808 25449 12828
rect 23510 12491 23540 12557
rect 17343 12164 17363 12184
rect 17767 12167 17788 12187
rect 17387 12105 17413 12131
rect 18192 12122 18218 12145
rect 18572 12115 18598 12138
rect 17554 12047 17575 12077
rect 17765 12018 17786 12038
rect 19665 12153 19705 12179
rect 19668 12108 19708 12134
rect 19672 12055 19712 12081
rect 17971 11910 18000 11937
rect 18045 11913 18074 11940
rect 17322 11853 17342 11873
rect 17554 11783 17571 11820
rect 20678 12337 20715 12378
rect 20734 12339 20771 12380
rect 20470 12260 20489 12280
rect 20547 12260 20566 12280
rect 19838 12159 19858 12179
rect 20262 12162 20283 12182
rect 23146 12418 23171 12453
rect 23190 12418 23215 12456
rect 23379 12359 23399 12379
rect 24427 12355 24447 12375
rect 20727 12147 20763 12168
rect 22647 12292 22676 12319
rect 22721 12295 22750 12322
rect 19882 12100 19908 12126
rect 20049 12042 20070 12072
rect 20260 12013 20281 12033
rect 20727 12091 20767 12128
rect 22452 12131 22501 12173
rect 22935 12194 22956 12214
rect 23695 12288 23724 12315
rect 23769 12291 23798 12318
rect 23146 12155 23167 12185
rect 22453 12068 22502 12110
rect 23308 12101 23334 12127
rect 20466 11905 20495 11932
rect 20540 11908 20569 11935
rect 19817 11848 19837 11868
rect 19995 11798 20027 11818
rect 20050 11799 20075 11819
rect 17704 11091 17729 11129
rect 19657 11705 19702 11744
rect 19422 11585 19441 11605
rect 19499 11585 19518 11605
rect 18790 11484 18810 11504
rect 19214 11487 19235 11507
rect 18834 11425 18860 11451
rect 19666 11448 19719 11481
rect 19001 11367 19022 11397
rect 19212 11338 19233 11358
rect 19671 11390 19724 11423
rect 20713 11674 20753 11707
rect 20470 11581 20489 11601
rect 20547 11581 20566 11601
rect 19838 11480 19858 11500
rect 20262 11483 20283 11503
rect 22933 12045 22954 12065
rect 23358 12048 23378 12068
rect 22650 11947 22669 11967
rect 22727 11947 22746 11967
rect 22463 11841 22503 11874
rect 23492 12125 23545 12158
rect 23983 12190 24004 12210
rect 24194 12151 24215 12181
rect 23497 12067 23550 12100
rect 24356 12097 24382 12123
rect 23981 12041 24002 12061
rect 24406 12044 24426 12064
rect 23698 11943 23717 11963
rect 23775 11943 23794 11963
rect 23514 11804 23559 11843
rect 25145 12710 25164 12730
rect 25222 12710 25241 12730
rect 25853 12811 25873 12831
rect 25652 12620 25704 12638
rect 25421 12419 25446 12454
rect 25465 12419 25490 12457
rect 25684 12435 25708 12458
rect 25684 12391 25708 12414
rect 23141 11729 23166 11749
rect 23189 11730 23221 11750
rect 23379 11680 23399 11700
rect 22647 11613 22676 11640
rect 22721 11616 22750 11643
rect 19882 11421 19908 11447
rect 20714 11438 20763 11480
rect 20049 11363 20070 11393
rect 19418 11230 19447 11257
rect 19492 11233 19521 11260
rect 20260 11334 20281 11354
rect 20715 11375 20764 11417
rect 22449 11420 22489 11457
rect 22935 11515 22956 11535
rect 23146 11476 23167 11506
rect 23308 11422 23334 11448
rect 20466 11226 20495 11253
rect 20540 11229 20569 11256
rect 22453 11380 22489 11401
rect 18769 11173 18789 11193
rect 19817 11169 19837 11189
rect 20001 11092 20026 11130
rect 20045 11095 20070 11130
rect 22933 11366 22954 11386
rect 23358 11369 23378 11389
rect 22650 11268 22669 11288
rect 22727 11268 22746 11288
rect 22445 11168 22482 11209
rect 22501 11170 22538 11211
rect 23504 11467 23544 11493
rect 23508 11414 23548 11440
rect 23511 11369 23551 11395
rect 23503 11109 23547 11146
rect 25689 11772 25709 11793
rect 25730 11777 25750 11798
rect 25917 11677 25937 11697
rect 25185 11610 25214 11637
rect 25259 11613 25288 11640
rect 25473 11512 25494 11532
rect 25684 11473 25705 11503
rect 25846 11419 25872 11445
rect 19665 10939 19719 11005
rect 23498 11023 23552 11089
rect 17933 10743 17952 10763
rect 18010 10743 18029 10763
rect 17301 10642 17321 10662
rect 17725 10645 17746 10665
rect 17345 10583 17371 10609
rect 17512 10525 17533 10555
rect 17723 10496 17744 10516
rect 17929 10388 17958 10415
rect 18003 10391 18032 10418
rect 17280 10331 17300 10351
rect 19670 10882 19714 10919
rect 19666 10633 19706 10659
rect 19669 10588 19709 10614
rect 19673 10535 19713 10561
rect 20679 10817 20716 10858
rect 20735 10819 20772 10860
rect 20471 10740 20490 10760
rect 20548 10740 20567 10760
rect 19839 10639 19859 10659
rect 20263 10642 20284 10662
rect 23147 10898 23172 10933
rect 23191 10898 23216 10936
rect 23380 10839 23400 10859
rect 24428 10835 24448 10855
rect 20728 10627 20764 10648
rect 22648 10772 22677 10799
rect 22722 10775 22751 10802
rect 19883 10580 19909 10606
rect 20050 10522 20071 10552
rect 20261 10493 20282 10513
rect 20728 10571 20768 10608
rect 22453 10611 22502 10653
rect 22936 10674 22957 10694
rect 23696 10768 23725 10795
rect 23770 10771 23799 10798
rect 23147 10635 23168 10665
rect 22454 10548 22503 10590
rect 23309 10581 23335 10607
rect 20467 10385 20496 10412
rect 20541 10388 20570 10415
rect 19818 10328 19838 10348
rect 19996 10278 20028 10298
rect 20051 10279 20076 10299
rect 17509 9614 17533 9637
rect 17509 9570 17533 9593
rect 17727 9571 17752 9609
rect 17771 9574 17796 9609
rect 17513 9390 17565 9408
rect 17344 9197 17364 9217
rect 17976 9298 17995 9318
rect 18053 9298 18072 9318
rect 19658 10185 19703 10224
rect 19423 10065 19442 10085
rect 19500 10065 19519 10085
rect 18791 9964 18811 9984
rect 19215 9967 19236 9987
rect 18835 9905 18861 9931
rect 19667 9928 19720 9961
rect 19002 9847 19023 9877
rect 19213 9818 19234 9838
rect 19672 9870 19725 9903
rect 20714 10154 20754 10187
rect 20471 10061 20490 10081
rect 20548 10061 20567 10081
rect 19839 9960 19859 9980
rect 20263 9963 20284 9983
rect 22934 10525 22955 10545
rect 23359 10528 23379 10548
rect 22651 10427 22670 10447
rect 22728 10427 22747 10447
rect 22464 10321 22504 10354
rect 23493 10605 23546 10638
rect 23984 10670 24005 10690
rect 24195 10631 24216 10661
rect 23498 10547 23551 10580
rect 24357 10577 24383 10603
rect 23982 10521 24003 10541
rect 24407 10524 24427 10544
rect 23699 10423 23718 10443
rect 23776 10423 23795 10443
rect 23515 10284 23560 10323
rect 23142 10209 23167 10229
rect 23190 10210 23222 10230
rect 23380 10160 23400 10180
rect 22648 10093 22677 10120
rect 22722 10096 22751 10123
rect 19883 9901 19909 9927
rect 20715 9918 20764 9960
rect 20050 9843 20071 9873
rect 19419 9710 19448 9737
rect 19493 9713 19522 9740
rect 20261 9814 20282 9834
rect 20716 9855 20765 9897
rect 22450 9900 22490 9937
rect 22936 9995 22957 10015
rect 23147 9956 23168 9986
rect 23309 9902 23335 9928
rect 20467 9706 20496 9733
rect 20541 9709 20570 9736
rect 22454 9860 22490 9881
rect 18770 9653 18790 9673
rect 19818 9649 19838 9669
rect 20002 9572 20027 9610
rect 20046 9575 20071 9610
rect 22934 9846 22955 9866
rect 23359 9849 23379 9869
rect 22651 9748 22670 9768
rect 22728 9748 22747 9768
rect 22446 9648 22483 9689
rect 22502 9650 22539 9691
rect 23505 9947 23545 9973
rect 23509 9894 23549 9920
rect 23512 9849 23552 9875
rect 24619 9890 24645 9913
rect 19677 9471 19707 9537
rect 17768 9200 17789 9220
rect 17388 9138 17414 9164
rect 18380 9170 18434 9211
rect 17555 9080 17576 9110
rect 17766 9051 17787 9071
rect 23511 9524 23541 9590
rect 19666 9186 19706 9212
rect 19669 9141 19709 9167
rect 19673 9088 19713 9114
rect 20679 9370 20716 9411
rect 20735 9372 20772 9413
rect 20471 9293 20490 9313
rect 20548 9293 20567 9313
rect 19839 9192 19859 9212
rect 20263 9195 20284 9215
rect 23147 9451 23172 9486
rect 23191 9451 23216 9489
rect 23380 9392 23400 9412
rect 24428 9388 24448 9408
rect 20728 9180 20764 9201
rect 22648 9325 22677 9352
rect 22722 9328 22751 9355
rect 19883 9133 19909 9159
rect 20050 9075 20071 9105
rect 17972 8943 18001 8970
rect 18046 8946 18075 8973
rect 17323 8886 17343 8906
rect 15625 8195 15654 8229
rect 15624 8135 15653 8169
rect 13840 8050 13884 8078
rect 13649 7951 13686 7999
rect 13837 7993 13881 8021
rect 8955 7598 8995 7624
rect 8958 7553 8998 7579
rect 8962 7500 9002 7526
rect 16132 7911 16195 7965
rect 9968 7782 10005 7823
rect 10024 7784 10061 7825
rect 9760 7705 9779 7725
rect 9837 7705 9856 7725
rect 9128 7604 9148 7624
rect 9552 7607 9573 7627
rect 12179 7853 12204 7888
rect 12223 7853 12248 7891
rect 12412 7794 12432 7814
rect 13229 7854 13254 7889
rect 13273 7854 13298 7892
rect 10017 7592 10053 7613
rect 13460 7790 13480 7810
rect 11680 7727 11709 7754
rect 11754 7730 11783 7757
rect 9172 7545 9198 7571
rect 9339 7487 9360 7517
rect 9550 7458 9571 7478
rect 10017 7536 10057 7573
rect 11485 7566 11534 7608
rect 11968 7629 11989 7649
rect 12728 7723 12757 7750
rect 12802 7726 12831 7753
rect 12179 7590 12200 7620
rect 11486 7503 11535 7545
rect 12341 7536 12367 7562
rect 9756 7350 9785 7377
rect 9830 7353 9859 7380
rect 9107 7293 9127 7313
rect 9285 7243 9317 7263
rect 9340 7244 9365 7264
rect 8947 7150 8992 7189
rect 8712 7030 8731 7050
rect 8789 7030 8808 7050
rect 8080 6929 8100 6949
rect 8504 6932 8525 6952
rect 8124 6870 8150 6896
rect 8956 6893 9009 6926
rect 8291 6812 8312 6842
rect 8502 6783 8523 6803
rect 8961 6835 9014 6868
rect 10003 7119 10043 7152
rect 9760 7026 9779 7046
rect 9837 7026 9856 7046
rect 9128 6925 9148 6945
rect 9552 6928 9573 6948
rect 11966 7480 11987 7500
rect 12391 7483 12411 7503
rect 11683 7382 11702 7402
rect 11760 7382 11779 7402
rect 11496 7276 11536 7309
rect 12525 7560 12578 7593
rect 13016 7625 13037 7645
rect 13227 7586 13248 7616
rect 12530 7502 12583 7535
rect 13389 7532 13415 7558
rect 13014 7476 13035 7496
rect 13439 7479 13459 7499
rect 12731 7378 12750 7398
rect 12808 7378 12827 7398
rect 12547 7239 12592 7278
rect 13650 7539 13684 7578
rect 12174 7164 12199 7184
rect 12222 7165 12254 7185
rect 12412 7115 12432 7135
rect 11680 7048 11709 7075
rect 11754 7051 11783 7078
rect 9172 6866 9198 6892
rect 10004 6883 10053 6925
rect 9339 6808 9360 6838
rect 8708 6675 8737 6702
rect 8782 6678 8811 6705
rect 9550 6779 9571 6799
rect 10005 6820 10054 6862
rect 11482 6855 11522 6892
rect 11968 6950 11989 6970
rect 13827 7559 13863 7600
rect 13816 7219 13876 7263
rect 14907 7110 14927 7130
rect 14175 7043 14204 7070
rect 14249 7046 14278 7073
rect 12179 6911 12200 6941
rect 12341 6857 12367 6883
rect 9756 6671 9785 6698
rect 9830 6674 9859 6701
rect 8059 6618 8079 6638
rect 11486 6815 11522 6836
rect 9107 6614 9127 6634
rect 9291 6537 9316 6575
rect 9335 6540 9360 6575
rect 11966 6801 11987 6821
rect 12391 6804 12411 6824
rect 11683 6703 11702 6723
rect 11760 6703 11779 6723
rect 11478 6603 11515 6644
rect 11534 6605 11571 6646
rect 12537 6902 12577 6928
rect 12541 6849 12581 6875
rect 12544 6804 12584 6830
rect 8966 6436 8996 6502
rect 14463 6945 14484 6965
rect 14674 6906 14695 6936
rect 13816 6805 13870 6846
rect 14836 6852 14862 6878
rect 14461 6796 14482 6816
rect 12543 6479 12573 6545
rect 7862 6113 7888 6136
rect 8955 6151 8995 6177
rect 8958 6106 8998 6132
rect 8962 6053 9002 6079
rect 9968 6335 10005 6376
rect 10024 6337 10061 6378
rect 9760 6258 9779 6278
rect 9837 6258 9856 6278
rect 9128 6157 9148 6177
rect 9552 6160 9573 6180
rect 12179 6406 12204 6441
rect 12223 6406 12248 6444
rect 12412 6347 12432 6367
rect 10017 6145 10053 6166
rect 13460 6343 13480 6363
rect 11680 6280 11709 6307
rect 11754 6283 11783 6310
rect 9172 6098 9198 6124
rect 9339 6040 9360 6070
rect 9550 6011 9571 6031
rect 10017 6089 10057 6126
rect 11485 6119 11534 6161
rect 11968 6182 11989 6202
rect 12728 6276 12757 6303
rect 12802 6279 12831 6306
rect 12179 6143 12200 6173
rect 11486 6056 11535 6098
rect 12341 6089 12367 6115
rect 9756 5903 9785 5930
rect 9830 5906 9859 5933
rect 9107 5846 9127 5866
rect 9285 5796 9317 5816
rect 9340 5797 9365 5817
rect 8947 5703 8992 5742
rect 8712 5583 8731 5603
rect 8789 5583 8808 5603
rect 8080 5482 8100 5502
rect 8504 5485 8525 5505
rect 8124 5423 8150 5449
rect 8956 5446 9009 5479
rect 8291 5365 8312 5395
rect 8502 5336 8523 5356
rect 8961 5388 9014 5421
rect 10003 5672 10043 5705
rect 9760 5579 9779 5599
rect 9837 5579 9856 5599
rect 9128 5478 9148 5498
rect 9552 5481 9573 5501
rect 11966 6033 11987 6053
rect 12391 6036 12411 6056
rect 11683 5935 11702 5955
rect 11760 5935 11779 5955
rect 11496 5829 11536 5862
rect 12525 6113 12578 6146
rect 13016 6178 13037 6198
rect 13227 6139 13248 6169
rect 12530 6055 12583 6088
rect 13389 6085 13415 6111
rect 13014 6029 13035 6049
rect 13439 6032 13459 6052
rect 12731 5931 12750 5951
rect 12808 5931 12827 5951
rect 12547 5792 12592 5831
rect 14178 6698 14197 6718
rect 14255 6698 14274 6718
rect 14886 6799 14906 6819
rect 14685 6608 14737 6626
rect 14454 6407 14479 6442
rect 14498 6407 14523 6445
rect 14717 6423 14741 6446
rect 14717 6379 14741 6402
rect 12174 5717 12199 5737
rect 12222 5718 12254 5738
rect 12412 5668 12432 5688
rect 11680 5601 11709 5628
rect 11754 5604 11783 5631
rect 9172 5419 9198 5445
rect 10004 5436 10053 5478
rect 9339 5361 9360 5391
rect 8708 5228 8737 5255
rect 8782 5231 8811 5258
rect 9550 5332 9571 5352
rect 10005 5373 10054 5415
rect 11482 5408 11522 5445
rect 11968 5503 11989 5523
rect 12179 5464 12200 5494
rect 12341 5410 12367 5436
rect 9756 5224 9785 5251
rect 9830 5227 9859 5254
rect 8059 5171 8079 5191
rect 11486 5368 11522 5389
rect 9107 5167 9127 5187
rect 9291 5090 9316 5128
rect 9335 5093 9360 5128
rect 11966 5354 11987 5374
rect 12391 5357 12411 5377
rect 11683 5256 11702 5276
rect 11760 5256 11779 5276
rect 11478 5156 11515 5197
rect 11534 5158 11571 5199
rect 12537 5455 12577 5481
rect 12541 5402 12581 5428
rect 12544 5357 12584 5383
rect 12536 5097 12580 5134
rect 14950 5665 14970 5685
rect 14218 5598 14247 5625
rect 14292 5601 14321 5628
rect 14506 5500 14527 5520
rect 14717 5461 14738 5491
rect 14879 5407 14905 5433
rect 8955 4937 9009 5003
rect 12531 5011 12585 5077
rect 6635 4581 6661 4607
rect 6802 4523 6823 4553
rect 7013 4494 7034 4514
rect 7219 4386 7248 4413
rect 7293 4389 7322 4416
rect 6570 4329 6590 4349
rect 3971 4202 3988 4239
rect 6757 4228 6777 4249
rect 6798 4233 6818 4254
rect 4200 4149 4220 4169
rect 3468 4082 3497 4109
rect 3542 4085 3571 4112
rect 3756 3984 3777 4004
rect 3967 3945 3988 3975
rect 3324 3877 3350 3900
rect 4129 3891 4155 3917
rect 3754 3835 3775 3855
rect 4179 3838 4199 3858
rect 3471 3737 3490 3757
rect 3548 3737 3567 3757
rect 8960 4880 9004 4917
rect 8956 4631 8996 4657
rect 8959 4586 8999 4612
rect 8963 4533 9003 4559
rect 9969 4815 10006 4856
rect 10025 4817 10062 4858
rect 9761 4738 9780 4758
rect 9838 4738 9857 4758
rect 9129 4637 9149 4657
rect 9553 4640 9574 4660
rect 12180 4886 12205 4921
rect 12224 4886 12249 4924
rect 12413 4827 12433 4847
rect 10018 4625 10054 4646
rect 13461 4823 13481 4843
rect 11681 4760 11710 4787
rect 11755 4763 11784 4790
rect 9173 4578 9199 4604
rect 9340 4520 9361 4550
rect 9551 4491 9572 4511
rect 10018 4569 10058 4606
rect 11486 4599 11535 4641
rect 11969 4662 11990 4682
rect 12729 4756 12758 4783
rect 12803 4759 12832 4786
rect 12180 4623 12201 4653
rect 11487 4536 11536 4578
rect 12342 4569 12368 4595
rect 9757 4383 9786 4410
rect 9831 4386 9860 4413
rect 9108 4326 9128 4346
rect 9286 4276 9318 4296
rect 9341 4277 9366 4297
rect 6799 3612 6823 3635
rect 6799 3568 6823 3591
rect 7017 3569 7042 3607
rect 7061 3572 7086 3607
rect 3811 3465 3839 3493
rect 6803 3388 6855 3406
rect 6634 3195 6654 3215
rect 7266 3296 7285 3316
rect 7343 3296 7362 3316
rect 8948 4183 8993 4222
rect 8713 4063 8732 4083
rect 8790 4063 8809 4083
rect 8081 3962 8101 3982
rect 8505 3965 8526 3985
rect 8125 3903 8151 3929
rect 8957 3926 9010 3959
rect 8292 3845 8313 3875
rect 8503 3816 8524 3836
rect 8962 3868 9015 3901
rect 10004 4152 10044 4185
rect 9761 4059 9780 4079
rect 9838 4059 9857 4079
rect 9129 3958 9149 3978
rect 9553 3961 9574 3981
rect 11967 4513 11988 4533
rect 12392 4516 12412 4536
rect 11684 4415 11703 4435
rect 11761 4415 11780 4435
rect 11497 4309 11537 4342
rect 12526 4593 12579 4626
rect 13017 4658 13038 4678
rect 13228 4619 13249 4649
rect 12531 4535 12584 4568
rect 13390 4565 13416 4591
rect 13015 4509 13036 4529
rect 13440 4512 13460 4532
rect 12732 4411 12751 4431
rect 12809 4411 12828 4431
rect 12548 4272 12593 4311
rect 12175 4197 12200 4217
rect 12223 4198 12255 4218
rect 12413 4148 12433 4168
rect 11681 4081 11710 4108
rect 11755 4084 11784 4111
rect 9173 3899 9199 3925
rect 10005 3916 10054 3958
rect 9340 3841 9361 3871
rect 8709 3708 8738 3735
rect 8783 3711 8812 3738
rect 9551 3812 9572 3832
rect 10006 3853 10055 3895
rect 11483 3888 11523 3925
rect 11969 3983 11990 4003
rect 12180 3944 12201 3974
rect 12342 3890 12368 3916
rect 9757 3704 9786 3731
rect 9831 3707 9860 3734
rect 8060 3651 8080 3671
rect 11487 3848 11523 3869
rect 9108 3647 9128 3667
rect 9292 3570 9317 3608
rect 9336 3573 9361 3608
rect 11967 3834 11988 3854
rect 12392 3837 12412 3857
rect 11684 3736 11703 3756
rect 11761 3736 11780 3756
rect 11479 3636 11516 3677
rect 11535 3638 11572 3679
rect 12538 3935 12578 3961
rect 12542 3882 12582 3908
rect 12545 3837 12585 3863
rect 13607 3868 13632 3899
rect 13652 3878 13678 3901
rect 8967 3469 8997 3535
rect 7058 3198 7079 3218
rect 6678 3136 6704 3162
rect 7670 3168 7724 3209
rect 6845 3078 6866 3108
rect 7056 3049 7077 3069
rect 12544 3512 12574 3578
rect 8956 3184 8996 3210
rect 8959 3139 8999 3165
rect 8963 3086 9003 3112
rect 9969 3368 10006 3409
rect 10025 3370 10062 3411
rect 9761 3291 9780 3311
rect 9838 3291 9857 3311
rect 9129 3190 9149 3210
rect 9553 3193 9574 3213
rect 12180 3439 12205 3474
rect 12224 3439 12249 3477
rect 12413 3380 12433 3400
rect 10018 3178 10054 3199
rect 13461 3376 13481 3396
rect 11681 3313 11710 3340
rect 11755 3316 11784 3343
rect 9173 3131 9199 3157
rect 9340 3073 9361 3103
rect 7262 2941 7291 2968
rect 7336 2944 7365 2971
rect 6613 2884 6633 2904
rect 5953 2410 6084 2475
rect 7664 2751 7724 2795
rect 7677 2414 7713 2455
rect 9551 3044 9572 3064
rect 10018 3122 10058 3159
rect 11486 3152 11535 3194
rect 11969 3215 11990 3235
rect 12729 3309 12758 3336
rect 12803 3312 12832 3339
rect 12180 3176 12201 3206
rect 11487 3089 11536 3131
rect 12342 3122 12368 3148
rect 9757 2936 9786 2963
rect 9831 2939 9860 2966
rect 9108 2879 9128 2899
rect 9286 2829 9318 2849
rect 9341 2830 9366 2850
rect 7856 2436 7890 2475
rect 8948 2736 8993 2775
rect 8713 2616 8732 2636
rect 8790 2616 8809 2636
rect 8081 2515 8101 2535
rect 8505 2518 8526 2538
rect 8125 2456 8151 2482
rect 8957 2479 9010 2512
rect 2886 2183 2986 2290
rect 8292 2398 8313 2428
rect 8503 2369 8524 2389
rect 8962 2421 9015 2454
rect 10004 2705 10044 2738
rect 9761 2612 9780 2632
rect 9838 2612 9857 2632
rect 9129 2511 9149 2531
rect 9553 2514 9574 2534
rect 11967 3066 11988 3086
rect 12392 3069 12412 3089
rect 11684 2968 11703 2988
rect 11761 2968 11780 2988
rect 11497 2862 11537 2895
rect 12526 3146 12579 3179
rect 13017 3211 13038 3231
rect 13228 3172 13249 3202
rect 12531 3088 12584 3121
rect 13390 3118 13416 3144
rect 13015 3062 13036 3082
rect 13440 3065 13460 3085
rect 12732 2964 12751 2984
rect 12809 2964 12828 2984
rect 12548 2825 12593 2864
rect 12175 2750 12200 2770
rect 12223 2751 12255 2771
rect 12413 2701 12433 2721
rect 11681 2634 11710 2661
rect 11755 2637 11784 2664
rect 9173 2452 9199 2478
rect 10005 2469 10054 2511
rect 9340 2394 9361 2424
rect 8709 2261 8738 2288
rect 8783 2264 8812 2291
rect 9551 2365 9572 2385
rect 10006 2406 10055 2448
rect 11483 2441 11523 2478
rect 11969 2536 11990 2556
rect 12180 2497 12201 2527
rect 12342 2443 12368 2469
rect 9757 2257 9786 2284
rect 9831 2260 9860 2287
rect 8060 2204 8080 2224
rect 11487 2401 11523 2422
rect 8242 2122 8267 2160
rect 8286 2125 8311 2160
rect 9108 2200 9128 2220
rect 9292 2123 9317 2161
rect 9336 2126 9361 2161
rect 11967 2387 11988 2407
rect 12392 2390 12412 2410
rect 11684 2289 11703 2309
rect 11761 2289 11780 2309
rect 11479 2189 11516 2230
rect 11535 2191 11572 2232
rect 14504 5351 14525 5371
rect 14929 5354 14949 5374
rect 14221 5253 14240 5273
rect 14298 5253 14317 5273
rect 14521 4887 14546 4925
rect 16597 7847 16626 7881
rect 16596 7787 16625 7821
rect 16865 7708 16884 7728
rect 16942 7708 16961 7728
rect 16233 7607 16253 7627
rect 16657 7610 16678 7630
rect 18374 8753 18434 8797
rect 18387 8416 18423 8457
rect 20261 9046 20282 9066
rect 20728 9124 20768 9161
rect 22453 9164 22502 9206
rect 22936 9227 22957 9247
rect 23696 9321 23725 9348
rect 23770 9324 23799 9351
rect 23147 9188 23168 9218
rect 22454 9101 22503 9143
rect 23309 9134 23335 9160
rect 20467 8938 20496 8965
rect 20541 8941 20570 8968
rect 19818 8881 19838 8901
rect 19996 8831 20028 8851
rect 20051 8832 20076 8852
rect 18566 8438 18600 8477
rect 19658 8738 19703 8777
rect 19423 8618 19442 8638
rect 19500 8618 19519 8638
rect 18791 8517 18811 8537
rect 19215 8520 19236 8540
rect 18835 8458 18861 8484
rect 19667 8481 19720 8514
rect 19002 8400 19023 8430
rect 19213 8371 19234 8391
rect 19672 8423 19725 8456
rect 20714 8707 20754 8740
rect 20471 8614 20490 8634
rect 20548 8614 20567 8634
rect 19839 8513 19859 8533
rect 20263 8516 20284 8536
rect 22934 9078 22955 9098
rect 23359 9081 23379 9101
rect 22651 8980 22670 9000
rect 22728 8980 22747 9000
rect 22464 8874 22504 8907
rect 23493 9158 23546 9191
rect 23984 9223 24005 9243
rect 24195 9184 24216 9214
rect 23498 9100 23551 9133
rect 24357 9130 24383 9156
rect 23982 9074 24003 9094
rect 24407 9077 24427 9097
rect 23699 8976 23718 8996
rect 23776 8976 23795 8996
rect 23515 8837 23560 8876
rect 23142 8762 23167 8782
rect 23190 8763 23222 8783
rect 23380 8713 23400 8733
rect 22648 8646 22677 8673
rect 22722 8649 22751 8676
rect 19883 8454 19909 8480
rect 20715 8471 20764 8513
rect 20050 8396 20071 8426
rect 19419 8263 19448 8290
rect 19493 8266 19522 8293
rect 20261 8367 20282 8387
rect 20716 8408 20765 8450
rect 22450 8453 22490 8490
rect 22936 8548 22957 8568
rect 23147 8509 23168 8539
rect 23309 8455 23335 8481
rect 20467 8259 20496 8286
rect 20541 8262 20570 8289
rect 22454 8413 22490 8434
rect 18770 8206 18790 8226
rect 18952 8124 18977 8162
rect 18996 8127 19021 8162
rect 19818 8202 19838 8222
rect 20002 8125 20027 8163
rect 20046 8128 20071 8163
rect 22934 8399 22955 8419
rect 23359 8402 23379 8422
rect 22651 8301 22670 8321
rect 22728 8301 22747 8321
rect 22446 8201 22483 8242
rect 22502 8203 22539 8244
rect 23505 8500 23545 8526
rect 23509 8447 23549 8473
rect 23512 8402 23552 8428
rect 16277 7548 16303 7574
rect 17087 7554 17111 7578
rect 17144 7555 17168 7579
rect 16444 7490 16465 7520
rect 16655 7461 16676 7481
rect 18369 7995 18413 8023
rect 18564 8017 18601 8065
rect 18366 7938 18410 7966
rect 16861 7353 16890 7380
rect 16935 7356 16964 7383
rect 16212 7296 16232 7316
rect 15974 4898 15999 4924
rect 16363 4829 16383 4849
rect 15631 4762 15660 4789
rect 15705 4765 15734 4792
rect 15919 4664 15940 4684
rect 16130 4625 16151 4655
rect 16292 4571 16318 4597
rect 15917 4515 15938 4535
rect 16121 4517 16154 4537
rect 16342 4518 16362 4538
rect 15634 4417 15653 4437
rect 15711 4417 15730 4437
rect 16442 4360 16465 4398
rect 17701 6521 17729 6549
rect 17973 6257 17992 6277
rect 18050 6257 18069 6277
rect 17341 6156 17361 6176
rect 17765 6159 17786 6179
rect 17385 6097 17411 6123
rect 18190 6114 18216 6137
rect 17552 6039 17573 6069
rect 17763 6010 17784 6030
rect 17969 5902 17998 5929
rect 18043 5905 18072 5932
rect 17320 5845 17340 5865
rect 17552 5775 17569 5812
rect 17702 5083 17727 5121
rect 17931 4735 17950 4755
rect 18008 4735 18027 4755
rect 17299 4634 17319 4654
rect 17723 4637 17744 4657
rect 19666 7891 19712 7939
rect 23503 8081 23549 8129
rect 25471 11363 25492 11383
rect 25896 11366 25916 11386
rect 25188 11265 25207 11285
rect 25265 11265 25284 11285
rect 25488 10899 25513 10937
rect 25646 10208 25663 10245
rect 25875 10155 25895 10175
rect 25143 10088 25172 10115
rect 25217 10091 25246 10118
rect 25431 9990 25452 10010
rect 25642 9951 25663 9981
rect 24999 9883 25025 9906
rect 25804 9897 25830 9923
rect 25429 9841 25450 9861
rect 25854 9844 25874 9864
rect 25146 9743 25165 9763
rect 25223 9743 25242 9763
rect 25486 9471 25514 9499
rect 26983 8704 27003 8724
rect 26251 8637 26280 8664
rect 26325 8640 26354 8667
rect 26539 8539 26560 8559
rect 26750 8500 26771 8530
rect 26047 8441 26071 8465
rect 26104 8442 26128 8466
rect 26912 8446 26938 8472
rect 26537 8390 26558 8410
rect 26750 8388 26774 8410
rect 26962 8393 26982 8413
rect 26254 8292 26273 8312
rect 26331 8292 26350 8312
rect 30637 13506 30677 13532
rect 31643 13788 31680 13829
rect 31699 13790 31736 13831
rect 31435 13711 31454 13731
rect 31512 13711 31531 13731
rect 30803 13610 30823 13630
rect 31227 13613 31248 13633
rect 33854 13859 33879 13894
rect 33898 13859 33923 13897
rect 34087 13800 34107 13820
rect 34904 13860 34929 13895
rect 34948 13860 34973 13898
rect 31692 13598 31728 13619
rect 35135 13796 35155 13816
rect 33355 13733 33384 13760
rect 33429 13736 33458 13763
rect 30847 13551 30873 13577
rect 31014 13493 31035 13523
rect 31225 13464 31246 13484
rect 31692 13542 31732 13579
rect 33160 13572 33209 13614
rect 33643 13635 33664 13655
rect 34403 13729 34432 13756
rect 34477 13732 34506 13759
rect 33854 13596 33875 13626
rect 33161 13509 33210 13551
rect 34016 13542 34042 13568
rect 31431 13356 31460 13383
rect 31505 13359 31534 13386
rect 30782 13299 30802 13319
rect 30960 13249 30992 13269
rect 31015 13250 31040 13270
rect 30622 13156 30667 13195
rect 30387 13036 30406 13056
rect 30464 13036 30483 13056
rect 29755 12935 29775 12955
rect 30179 12938 30200 12958
rect 29799 12876 29825 12902
rect 30631 12899 30684 12932
rect 29966 12818 29987 12848
rect 30177 12789 30198 12809
rect 30636 12841 30689 12874
rect 31678 13125 31718 13158
rect 31435 13032 31454 13052
rect 31512 13032 31531 13052
rect 30803 12931 30823 12951
rect 31227 12934 31248 12954
rect 33641 13486 33662 13506
rect 34066 13489 34086 13509
rect 33358 13388 33377 13408
rect 33435 13388 33454 13408
rect 33171 13282 33211 13315
rect 34200 13566 34253 13599
rect 34691 13631 34712 13651
rect 34902 13592 34923 13622
rect 34205 13508 34258 13541
rect 35064 13538 35090 13564
rect 34689 13482 34710 13502
rect 35114 13485 35134 13505
rect 34406 13384 34425 13404
rect 34483 13384 34502 13404
rect 34222 13245 34267 13284
rect 35325 13545 35359 13584
rect 33849 13170 33874 13190
rect 33897 13171 33929 13191
rect 34087 13121 34107 13141
rect 33355 13054 33384 13081
rect 33429 13057 33458 13084
rect 30847 12872 30873 12898
rect 31679 12889 31728 12931
rect 31014 12814 31035 12844
rect 30383 12681 30412 12708
rect 30457 12684 30486 12711
rect 31225 12785 31246 12805
rect 31680 12826 31729 12868
rect 33157 12861 33197 12898
rect 33643 12956 33664 12976
rect 35502 13565 35538 13606
rect 35491 13225 35551 13269
rect 36803 13667 36841 13764
rect 36863 13673 36901 13770
rect 41338 13598 41378 13624
rect 36582 13116 36602 13136
rect 35850 13049 35879 13076
rect 35924 13052 35953 13079
rect 33854 12917 33875 12947
rect 34016 12863 34042 12889
rect 31431 12677 31460 12704
rect 31505 12680 31534 12707
rect 29734 12624 29754 12644
rect 33161 12821 33197 12842
rect 30782 12620 30802 12640
rect 28668 12533 28696 12561
rect 30966 12543 30991 12581
rect 31010 12546 31035 12581
rect 33641 12807 33662 12827
rect 34066 12810 34086 12830
rect 33358 12709 33377 12729
rect 33435 12709 33454 12729
rect 33153 12609 33190 12650
rect 33209 12611 33246 12652
rect 34212 12908 34252 12934
rect 34216 12855 34256 12881
rect 34219 12810 34259 12836
rect 30641 12442 30671 12508
rect 28940 12269 28959 12289
rect 29017 12269 29036 12289
rect 36138 12951 36159 12971
rect 36349 12912 36370 12942
rect 35491 12811 35545 12852
rect 36511 12858 36537 12884
rect 36136 12802 36157 12822
rect 34218 12485 34248 12551
rect 28308 12168 28328 12188
rect 28732 12171 28753 12191
rect 28352 12109 28378 12135
rect 29157 12126 29183 12149
rect 29537 12119 29563 12142
rect 28519 12051 28540 12081
rect 28730 12022 28751 12042
rect 30630 12157 30670 12183
rect 30633 12112 30673 12138
rect 30637 12059 30677 12085
rect 28936 11914 28965 11941
rect 29010 11917 29039 11944
rect 28287 11857 28307 11877
rect 28519 11787 28536 11824
rect 31643 12341 31680 12382
rect 31699 12343 31736 12384
rect 31435 12264 31454 12284
rect 31512 12264 31531 12284
rect 30803 12163 30823 12183
rect 31227 12166 31248 12186
rect 33854 12412 33879 12447
rect 33898 12412 33923 12450
rect 34087 12353 34107 12373
rect 31692 12151 31728 12172
rect 35135 12349 35155 12369
rect 33355 12286 33384 12313
rect 33429 12289 33458 12316
rect 30847 12104 30873 12130
rect 31014 12046 31035 12076
rect 31225 12017 31246 12037
rect 31692 12095 31732 12132
rect 33160 12125 33209 12167
rect 33643 12188 33664 12208
rect 34403 12282 34432 12309
rect 34477 12285 34506 12312
rect 33854 12149 33875 12179
rect 33161 12062 33210 12104
rect 34016 12095 34042 12121
rect 31431 11909 31460 11936
rect 31505 11912 31534 11939
rect 30782 11852 30802 11872
rect 30960 11802 30992 11822
rect 31015 11803 31040 11823
rect 28669 11095 28694 11133
rect 30622 11709 30667 11748
rect 30387 11589 30406 11609
rect 30464 11589 30483 11609
rect 29755 11488 29775 11508
rect 30179 11491 30200 11511
rect 29799 11429 29825 11455
rect 30631 11452 30684 11485
rect 29966 11371 29987 11401
rect 30177 11342 30198 11362
rect 30636 11394 30689 11427
rect 31678 11678 31718 11711
rect 31435 11585 31454 11605
rect 31512 11585 31531 11605
rect 30803 11484 30823 11504
rect 31227 11487 31248 11507
rect 33641 12039 33662 12059
rect 34066 12042 34086 12062
rect 33358 11941 33377 11961
rect 33435 11941 33454 11961
rect 33171 11835 33211 11868
rect 34200 12119 34253 12152
rect 34691 12184 34712 12204
rect 34902 12145 34923 12175
rect 34205 12061 34258 12094
rect 35064 12091 35090 12117
rect 34689 12035 34710 12055
rect 35114 12038 35134 12058
rect 34406 11937 34425 11957
rect 34483 11937 34502 11957
rect 34222 11798 34267 11837
rect 35853 12704 35872 12724
rect 35930 12704 35949 12724
rect 36561 12805 36581 12825
rect 36360 12614 36412 12632
rect 36129 12413 36154 12448
rect 36173 12413 36198 12451
rect 36392 12429 36416 12452
rect 36392 12385 36416 12408
rect 33849 11723 33874 11743
rect 33897 11724 33929 11744
rect 34087 11674 34107 11694
rect 33355 11607 33384 11634
rect 33429 11610 33458 11637
rect 30847 11425 30873 11451
rect 31679 11442 31728 11484
rect 31014 11367 31035 11397
rect 30383 11234 30412 11261
rect 30457 11237 30486 11264
rect 31225 11338 31246 11358
rect 31680 11379 31729 11421
rect 33157 11414 33197 11451
rect 33643 11509 33664 11529
rect 33854 11470 33875 11500
rect 34016 11416 34042 11442
rect 31431 11230 31460 11257
rect 31505 11233 31534 11260
rect 29734 11177 29754 11197
rect 33161 11374 33197 11395
rect 30782 11173 30802 11193
rect 30966 11096 30991 11134
rect 31010 11099 31035 11134
rect 33641 11360 33662 11380
rect 34066 11363 34086 11383
rect 33358 11262 33377 11282
rect 33435 11262 33454 11282
rect 33153 11162 33190 11203
rect 33209 11164 33246 11205
rect 34212 11461 34252 11487
rect 34216 11408 34256 11434
rect 34219 11363 34259 11389
rect 34211 11103 34255 11140
rect 36397 11766 36417 11787
rect 36438 11771 36458 11792
rect 36625 11671 36645 11691
rect 35893 11604 35922 11631
rect 35967 11607 35996 11634
rect 36181 11506 36202 11526
rect 36392 11467 36413 11497
rect 36554 11413 36580 11439
rect 30630 10943 30684 11009
rect 34206 11017 34260 11083
rect 28898 10747 28917 10767
rect 28975 10747 28994 10767
rect 28266 10646 28286 10666
rect 28690 10649 28711 10669
rect 28310 10587 28336 10613
rect 28477 10529 28498 10559
rect 28688 10500 28709 10520
rect 28894 10392 28923 10419
rect 28968 10395 28997 10422
rect 28245 10335 28265 10355
rect 30635 10886 30679 10923
rect 30631 10637 30671 10663
rect 30634 10592 30674 10618
rect 30638 10539 30678 10565
rect 31644 10821 31681 10862
rect 31700 10823 31737 10864
rect 31436 10744 31455 10764
rect 31513 10744 31532 10764
rect 30804 10643 30824 10663
rect 31228 10646 31249 10666
rect 33855 10892 33880 10927
rect 33899 10892 33924 10930
rect 34088 10833 34108 10853
rect 31693 10631 31729 10652
rect 35136 10829 35156 10849
rect 33356 10766 33385 10793
rect 33430 10769 33459 10796
rect 30848 10584 30874 10610
rect 31015 10526 31036 10556
rect 31226 10497 31247 10517
rect 31693 10575 31733 10612
rect 33161 10605 33210 10647
rect 33644 10668 33665 10688
rect 34404 10762 34433 10789
rect 34478 10765 34507 10792
rect 33855 10629 33876 10659
rect 33162 10542 33211 10584
rect 34017 10575 34043 10601
rect 31432 10389 31461 10416
rect 31506 10392 31535 10419
rect 30783 10332 30803 10352
rect 30961 10282 30993 10302
rect 31016 10283 31041 10303
rect 28474 9618 28498 9641
rect 28474 9574 28498 9597
rect 28692 9575 28717 9613
rect 28736 9578 28761 9613
rect 28478 9394 28530 9412
rect 28309 9201 28329 9221
rect 28941 9302 28960 9322
rect 29018 9302 29037 9322
rect 30623 10189 30668 10228
rect 30388 10069 30407 10089
rect 30465 10069 30484 10089
rect 29756 9968 29776 9988
rect 30180 9971 30201 9991
rect 29800 9909 29826 9935
rect 30632 9932 30685 9965
rect 29967 9851 29988 9881
rect 30178 9822 30199 9842
rect 30637 9874 30690 9907
rect 31679 10158 31719 10191
rect 31436 10065 31455 10085
rect 31513 10065 31532 10085
rect 30804 9964 30824 9984
rect 31228 9967 31249 9987
rect 33642 10519 33663 10539
rect 34067 10522 34087 10542
rect 33359 10421 33378 10441
rect 33436 10421 33455 10441
rect 33172 10315 33212 10348
rect 34201 10599 34254 10632
rect 34692 10664 34713 10684
rect 34903 10625 34924 10655
rect 34206 10541 34259 10574
rect 35065 10571 35091 10597
rect 34690 10515 34711 10535
rect 35115 10518 35135 10538
rect 34407 10417 34426 10437
rect 34484 10417 34503 10437
rect 34223 10278 34268 10317
rect 33850 10203 33875 10223
rect 33898 10204 33930 10224
rect 34088 10154 34108 10174
rect 33356 10087 33385 10114
rect 33430 10090 33459 10117
rect 30848 9905 30874 9931
rect 31680 9922 31729 9964
rect 31015 9847 31036 9877
rect 30384 9714 30413 9741
rect 30458 9717 30487 9744
rect 31226 9818 31247 9838
rect 31681 9859 31730 9901
rect 33158 9894 33198 9931
rect 33644 9989 33665 10009
rect 33855 9950 33876 9980
rect 34017 9896 34043 9922
rect 31432 9710 31461 9737
rect 31506 9713 31535 9740
rect 29735 9657 29755 9677
rect 33162 9854 33198 9875
rect 30783 9653 30803 9673
rect 30967 9576 30992 9614
rect 31011 9579 31036 9614
rect 33642 9840 33663 9860
rect 34067 9843 34087 9863
rect 33359 9742 33378 9762
rect 33436 9742 33455 9762
rect 33154 9642 33191 9683
rect 33210 9644 33247 9685
rect 34213 9941 34253 9967
rect 34217 9888 34257 9914
rect 34220 9843 34260 9869
rect 35327 9884 35353 9907
rect 30642 9475 30672 9541
rect 28733 9204 28754 9224
rect 28353 9142 28379 9168
rect 29345 9174 29399 9215
rect 28520 9084 28541 9114
rect 28731 9055 28752 9075
rect 34219 9518 34249 9584
rect 30631 9190 30671 9216
rect 30634 9145 30674 9171
rect 30638 9092 30678 9118
rect 31644 9374 31681 9415
rect 31700 9376 31737 9417
rect 31436 9297 31455 9317
rect 31513 9297 31532 9317
rect 30804 9196 30824 9216
rect 31228 9199 31249 9219
rect 33855 9445 33880 9480
rect 33899 9445 33924 9483
rect 34088 9386 34108 9406
rect 31693 9184 31729 9205
rect 35136 9382 35156 9402
rect 33356 9319 33385 9346
rect 33430 9322 33459 9349
rect 30848 9137 30874 9163
rect 31015 9079 31036 9109
rect 28937 8947 28966 8974
rect 29011 8950 29040 8977
rect 28288 8890 28308 8910
rect 26590 8199 26619 8233
rect 26589 8139 26618 8173
rect 24805 8054 24849 8082
rect 24614 7955 24651 8003
rect 24802 7997 24846 8025
rect 19663 7592 19703 7618
rect 19666 7547 19706 7573
rect 19670 7494 19710 7520
rect 27097 7915 27160 7969
rect 20676 7776 20713 7817
rect 20732 7778 20769 7819
rect 20468 7699 20487 7719
rect 20545 7699 20564 7719
rect 19836 7598 19856 7618
rect 20260 7601 20281 7621
rect 23144 7857 23169 7892
rect 23188 7857 23213 7895
rect 23377 7798 23397 7818
rect 24194 7858 24219 7893
rect 24238 7858 24263 7896
rect 24425 7794 24445 7814
rect 20725 7586 20761 7607
rect 22645 7731 22674 7758
rect 22719 7734 22748 7761
rect 19880 7539 19906 7565
rect 20047 7481 20068 7511
rect 20258 7452 20279 7472
rect 20725 7530 20765 7567
rect 22450 7570 22499 7612
rect 22933 7633 22954 7653
rect 23693 7727 23722 7754
rect 23767 7730 23796 7757
rect 23144 7594 23165 7624
rect 22451 7507 22500 7549
rect 23306 7540 23332 7566
rect 20464 7344 20493 7371
rect 20538 7347 20567 7374
rect 19815 7287 19835 7307
rect 19993 7237 20025 7257
rect 20048 7238 20073 7258
rect 19655 7144 19700 7183
rect 19420 7024 19439 7044
rect 19497 7024 19516 7044
rect 18788 6923 18808 6943
rect 19212 6926 19233 6946
rect 18832 6864 18858 6890
rect 19664 6887 19717 6920
rect 18999 6806 19020 6836
rect 19210 6777 19231 6797
rect 19669 6829 19722 6862
rect 20711 7113 20751 7146
rect 20468 7020 20487 7040
rect 20545 7020 20564 7040
rect 19836 6919 19856 6939
rect 20260 6922 20281 6942
rect 22931 7484 22952 7504
rect 23356 7487 23376 7507
rect 22648 7386 22667 7406
rect 22725 7386 22744 7406
rect 22461 7280 22501 7313
rect 23490 7564 23543 7597
rect 23981 7629 24002 7649
rect 24192 7590 24213 7620
rect 23495 7506 23548 7539
rect 24354 7536 24380 7562
rect 23979 7480 24000 7500
rect 24404 7483 24424 7503
rect 23696 7382 23715 7402
rect 23773 7382 23792 7402
rect 23512 7243 23557 7282
rect 24615 7543 24649 7582
rect 23139 7168 23164 7188
rect 23187 7169 23219 7189
rect 23377 7119 23397 7139
rect 22645 7052 22674 7079
rect 22719 7055 22748 7082
rect 19880 6860 19906 6886
rect 20712 6877 20761 6919
rect 20047 6802 20068 6832
rect 19416 6669 19445 6696
rect 19490 6672 19519 6699
rect 20258 6773 20279 6793
rect 20713 6814 20762 6856
rect 22447 6859 22487 6896
rect 22933 6954 22954 6974
rect 24792 7563 24828 7604
rect 24781 7223 24841 7267
rect 25872 7114 25892 7134
rect 25140 7047 25169 7074
rect 25214 7050 25243 7077
rect 23144 6915 23165 6945
rect 23306 6861 23332 6887
rect 20464 6665 20493 6692
rect 20538 6668 20567 6695
rect 22451 6819 22487 6840
rect 18767 6612 18787 6632
rect 19815 6608 19835 6628
rect 19999 6531 20024 6569
rect 20043 6534 20068 6569
rect 22931 6805 22952 6825
rect 23356 6808 23376 6828
rect 22648 6707 22667 6727
rect 22725 6707 22744 6727
rect 22443 6607 22480 6648
rect 22499 6609 22536 6650
rect 23502 6906 23542 6932
rect 23506 6853 23546 6879
rect 23509 6808 23549 6834
rect 19674 6430 19704 6496
rect 25428 6949 25449 6969
rect 25639 6910 25660 6940
rect 24781 6809 24835 6850
rect 25801 6856 25827 6882
rect 25426 6800 25447 6820
rect 23508 6483 23538 6549
rect 18570 6107 18596 6130
rect 19663 6145 19703 6171
rect 19666 6100 19706 6126
rect 19670 6047 19710 6073
rect 20676 6329 20713 6370
rect 20732 6331 20769 6372
rect 20468 6252 20487 6272
rect 20545 6252 20564 6272
rect 19836 6151 19856 6171
rect 20260 6154 20281 6174
rect 23144 6410 23169 6445
rect 23188 6410 23213 6448
rect 23377 6351 23397 6371
rect 24425 6347 24445 6367
rect 20725 6139 20761 6160
rect 22645 6284 22674 6311
rect 22719 6287 22748 6314
rect 19880 6092 19906 6118
rect 20047 6034 20068 6064
rect 20258 6005 20279 6025
rect 20725 6083 20765 6120
rect 22450 6123 22499 6165
rect 22933 6186 22954 6206
rect 23693 6280 23722 6307
rect 23767 6283 23796 6310
rect 23144 6147 23165 6177
rect 22451 6060 22500 6102
rect 23306 6093 23332 6119
rect 20464 5897 20493 5924
rect 20538 5900 20567 5927
rect 19815 5840 19835 5860
rect 19993 5790 20025 5810
rect 20048 5791 20073 5811
rect 19655 5697 19700 5736
rect 19420 5577 19439 5597
rect 19497 5577 19516 5597
rect 18788 5476 18808 5496
rect 19212 5479 19233 5499
rect 18832 5417 18858 5443
rect 19664 5440 19717 5473
rect 18999 5359 19020 5389
rect 19210 5330 19231 5350
rect 19669 5382 19722 5415
rect 20711 5666 20751 5699
rect 20468 5573 20487 5593
rect 20545 5573 20564 5593
rect 19836 5472 19856 5492
rect 20260 5475 20281 5495
rect 22931 6037 22952 6057
rect 23356 6040 23376 6060
rect 22648 5939 22667 5959
rect 22725 5939 22744 5959
rect 22461 5833 22501 5866
rect 23490 6117 23543 6150
rect 23981 6182 24002 6202
rect 24192 6143 24213 6173
rect 23495 6059 23548 6092
rect 24354 6089 24380 6115
rect 23979 6033 24000 6053
rect 24404 6036 24424 6056
rect 23696 5935 23715 5955
rect 23773 5935 23792 5955
rect 23512 5796 23557 5835
rect 25143 6702 25162 6722
rect 25220 6702 25239 6722
rect 25851 6803 25871 6823
rect 25650 6612 25702 6630
rect 25419 6411 25444 6446
rect 25463 6411 25488 6449
rect 25682 6427 25706 6450
rect 25682 6383 25706 6406
rect 23139 5721 23164 5741
rect 23187 5722 23219 5742
rect 23377 5672 23397 5692
rect 22645 5605 22674 5632
rect 22719 5608 22748 5635
rect 19880 5413 19906 5439
rect 20712 5430 20761 5472
rect 20047 5355 20068 5385
rect 19416 5222 19445 5249
rect 19490 5225 19519 5252
rect 20258 5326 20279 5346
rect 20713 5367 20762 5409
rect 22447 5412 22487 5449
rect 22933 5507 22954 5527
rect 23144 5468 23165 5498
rect 23306 5414 23332 5440
rect 20464 5218 20493 5245
rect 20538 5221 20567 5248
rect 22451 5372 22487 5393
rect 18767 5165 18787 5185
rect 19815 5161 19835 5181
rect 19999 5084 20024 5122
rect 20043 5087 20068 5122
rect 22931 5358 22952 5378
rect 23356 5361 23376 5381
rect 22648 5260 22667 5280
rect 22725 5260 22744 5280
rect 22443 5160 22480 5201
rect 22499 5162 22536 5203
rect 23502 5459 23542 5485
rect 23506 5406 23546 5432
rect 23509 5361 23549 5387
rect 23501 5101 23545 5138
rect 25915 5669 25935 5689
rect 25183 5602 25212 5629
rect 25257 5605 25286 5632
rect 25471 5504 25492 5524
rect 25682 5465 25703 5495
rect 25844 5411 25870 5437
rect 19663 4931 19717 4997
rect 23496 5015 23550 5081
rect 17343 4575 17369 4601
rect 17510 4517 17531 4547
rect 17721 4488 17742 4508
rect 17927 4380 17956 4407
rect 18001 4383 18030 4410
rect 17278 4323 17298 4343
rect 14679 4196 14696 4233
rect 17465 4222 17485 4243
rect 17506 4227 17526 4248
rect 14908 4143 14928 4163
rect 14176 4076 14205 4103
rect 14250 4079 14279 4106
rect 14464 3978 14485 3998
rect 14675 3939 14696 3969
rect 14032 3871 14058 3894
rect 14837 3885 14863 3911
rect 14462 3829 14483 3849
rect 14887 3832 14907 3852
rect 14179 3731 14198 3751
rect 14256 3731 14275 3751
rect 19668 4874 19712 4911
rect 19664 4625 19704 4651
rect 19667 4580 19707 4606
rect 19671 4527 19711 4553
rect 20677 4809 20714 4850
rect 20733 4811 20770 4852
rect 20469 4732 20488 4752
rect 20546 4732 20565 4752
rect 19837 4631 19857 4651
rect 20261 4634 20282 4654
rect 23145 4890 23170 4925
rect 23189 4890 23214 4928
rect 23378 4831 23398 4851
rect 24426 4827 24446 4847
rect 20726 4619 20762 4640
rect 22646 4764 22675 4791
rect 22720 4767 22749 4794
rect 19881 4572 19907 4598
rect 20048 4514 20069 4544
rect 20259 4485 20280 4505
rect 20726 4563 20766 4600
rect 22451 4603 22500 4645
rect 22934 4666 22955 4686
rect 23694 4760 23723 4787
rect 23768 4763 23797 4790
rect 23145 4627 23166 4657
rect 22452 4540 22501 4582
rect 23307 4573 23333 4599
rect 20465 4377 20494 4404
rect 20539 4380 20568 4407
rect 19816 4320 19836 4340
rect 19994 4270 20026 4290
rect 20049 4271 20074 4291
rect 17507 3606 17531 3629
rect 17507 3562 17531 3585
rect 17725 3563 17750 3601
rect 17769 3566 17794 3601
rect 14519 3459 14547 3487
rect 17511 3382 17563 3400
rect 17342 3189 17362 3209
rect 17974 3290 17993 3310
rect 18051 3290 18070 3310
rect 19656 4177 19701 4216
rect 19421 4057 19440 4077
rect 19498 4057 19517 4077
rect 18789 3956 18809 3976
rect 19213 3959 19234 3979
rect 18833 3897 18859 3923
rect 19665 3920 19718 3953
rect 19000 3839 19021 3869
rect 19211 3810 19232 3830
rect 19670 3862 19723 3895
rect 20712 4146 20752 4179
rect 20469 4053 20488 4073
rect 20546 4053 20565 4073
rect 19837 3952 19857 3972
rect 20261 3955 20282 3975
rect 22932 4517 22953 4537
rect 23357 4520 23377 4540
rect 22649 4419 22668 4439
rect 22726 4419 22745 4439
rect 22462 4313 22502 4346
rect 23491 4597 23544 4630
rect 23982 4662 24003 4682
rect 24193 4623 24214 4653
rect 23496 4539 23549 4572
rect 24355 4569 24381 4595
rect 23980 4513 24001 4533
rect 24405 4516 24425 4536
rect 23697 4415 23716 4435
rect 23774 4415 23793 4435
rect 23513 4276 23558 4315
rect 23140 4201 23165 4221
rect 23188 4202 23220 4222
rect 23378 4152 23398 4172
rect 22646 4085 22675 4112
rect 22720 4088 22749 4115
rect 19881 3893 19907 3919
rect 20713 3910 20762 3952
rect 20048 3835 20069 3865
rect 19417 3702 19446 3729
rect 19491 3705 19520 3732
rect 20259 3806 20280 3826
rect 20714 3847 20763 3889
rect 22448 3892 22488 3929
rect 22934 3987 22955 4007
rect 23145 3948 23166 3978
rect 23307 3894 23333 3920
rect 20465 3698 20494 3725
rect 20539 3701 20568 3728
rect 22452 3852 22488 3873
rect 18768 3645 18788 3665
rect 19816 3641 19836 3661
rect 20000 3564 20025 3602
rect 20044 3567 20069 3602
rect 22932 3838 22953 3858
rect 23357 3841 23377 3861
rect 22649 3740 22668 3760
rect 22726 3740 22745 3760
rect 22444 3640 22481 3681
rect 22500 3642 22537 3683
rect 23503 3939 23543 3965
rect 23507 3886 23547 3912
rect 23510 3841 23550 3867
rect 24572 3872 24597 3903
rect 24617 3882 24643 3905
rect 19675 3463 19705 3529
rect 17766 3192 17787 3212
rect 17386 3130 17412 3156
rect 18378 3162 18432 3203
rect 17553 3072 17574 3102
rect 17764 3043 17785 3063
rect 23509 3516 23539 3582
rect 19664 3178 19704 3204
rect 19667 3133 19707 3159
rect 19671 3080 19711 3106
rect 20677 3362 20714 3403
rect 20733 3364 20770 3405
rect 20469 3285 20488 3305
rect 20546 3285 20565 3305
rect 19837 3184 19857 3204
rect 20261 3187 20282 3207
rect 23145 3443 23170 3478
rect 23189 3443 23214 3481
rect 23378 3384 23398 3404
rect 24426 3380 24446 3400
rect 20726 3172 20762 3193
rect 22646 3317 22675 3344
rect 22720 3320 22749 3347
rect 19881 3125 19907 3151
rect 20048 3067 20069 3097
rect 17970 2935 17999 2962
rect 18044 2938 18073 2965
rect 17321 2878 17341 2898
rect 16661 2404 16792 2469
rect 18372 2745 18432 2789
rect 18385 2408 18421 2449
rect 20259 3038 20280 3058
rect 20726 3116 20766 3153
rect 22451 3156 22500 3198
rect 22934 3219 22955 3239
rect 23694 3313 23723 3340
rect 23768 3316 23797 3343
rect 23145 3180 23166 3210
rect 22452 3093 22501 3135
rect 23307 3126 23333 3152
rect 20465 2930 20494 2957
rect 20539 2933 20568 2960
rect 19816 2873 19836 2893
rect 19994 2823 20026 2843
rect 20049 2824 20074 2844
rect 18564 2430 18598 2469
rect 19656 2730 19701 2769
rect 19421 2610 19440 2630
rect 19498 2610 19517 2630
rect 18789 2509 18809 2529
rect 19213 2512 19234 2532
rect 18833 2450 18859 2476
rect 19665 2473 19718 2506
rect 13594 2177 13694 2284
rect 19000 2392 19021 2422
rect 19211 2363 19232 2383
rect 19670 2415 19723 2448
rect 20712 2699 20752 2732
rect 20469 2606 20488 2626
rect 20546 2606 20565 2626
rect 19837 2505 19857 2525
rect 20261 2508 20282 2528
rect 22932 3070 22953 3090
rect 23357 3073 23377 3093
rect 22649 2972 22668 2992
rect 22726 2972 22745 2992
rect 22462 2866 22502 2899
rect 23491 3150 23544 3183
rect 23982 3215 24003 3235
rect 24193 3176 24214 3206
rect 23496 3092 23549 3125
rect 24355 3122 24381 3148
rect 23980 3066 24001 3086
rect 24405 3069 24425 3089
rect 23697 2968 23716 2988
rect 23774 2968 23793 2988
rect 23513 2829 23558 2868
rect 23140 2754 23165 2774
rect 23188 2755 23220 2775
rect 23378 2705 23398 2725
rect 22646 2638 22675 2665
rect 22720 2641 22749 2668
rect 19881 2446 19907 2472
rect 20713 2463 20762 2505
rect 20048 2388 20069 2418
rect 19417 2255 19446 2282
rect 19491 2258 19520 2285
rect 20259 2359 20280 2379
rect 20714 2400 20763 2442
rect 22448 2445 22488 2482
rect 22934 2540 22955 2560
rect 23145 2501 23166 2531
rect 23307 2447 23333 2473
rect 20465 2251 20494 2278
rect 20539 2254 20568 2281
rect 22452 2405 22488 2426
rect 18768 2198 18788 2218
rect 18950 2116 18975 2154
rect 18994 2119 19019 2154
rect 19816 2194 19836 2214
rect 20000 2117 20025 2155
rect 20044 2120 20069 2155
rect 22932 2391 22953 2411
rect 23357 2394 23377 2414
rect 22649 2293 22668 2313
rect 22726 2293 22745 2313
rect 22444 2193 22481 2234
rect 22500 2195 22537 2236
rect 25469 5355 25490 5375
rect 25894 5358 25914 5378
rect 25186 5257 25205 5277
rect 25263 5257 25282 5277
rect 25486 4891 25511 4929
rect 27562 7851 27591 7885
rect 27561 7791 27590 7825
rect 27830 7712 27849 7732
rect 27907 7712 27926 7732
rect 27198 7611 27218 7631
rect 27622 7614 27643 7634
rect 29339 8757 29399 8801
rect 29352 8420 29388 8461
rect 31226 9050 31247 9070
rect 31693 9128 31733 9165
rect 33161 9158 33210 9200
rect 33644 9221 33665 9241
rect 34404 9315 34433 9342
rect 34478 9318 34507 9345
rect 33855 9182 33876 9212
rect 33162 9095 33211 9137
rect 34017 9128 34043 9154
rect 31432 8942 31461 8969
rect 31506 8945 31535 8972
rect 30783 8885 30803 8905
rect 30961 8835 30993 8855
rect 31016 8836 31041 8856
rect 29531 8442 29565 8481
rect 30623 8742 30668 8781
rect 30388 8622 30407 8642
rect 30465 8622 30484 8642
rect 29756 8521 29776 8541
rect 30180 8524 30201 8544
rect 29800 8462 29826 8488
rect 30632 8485 30685 8518
rect 29967 8404 29988 8434
rect 30178 8375 30199 8395
rect 30637 8427 30690 8460
rect 31679 8711 31719 8744
rect 31436 8618 31455 8638
rect 31513 8618 31532 8638
rect 30804 8517 30824 8537
rect 31228 8520 31249 8540
rect 33642 9072 33663 9092
rect 34067 9075 34087 9095
rect 33359 8974 33378 8994
rect 33436 8974 33455 8994
rect 33172 8868 33212 8901
rect 34201 9152 34254 9185
rect 34692 9217 34713 9237
rect 34903 9178 34924 9208
rect 34206 9094 34259 9127
rect 35065 9124 35091 9150
rect 34690 9068 34711 9088
rect 35115 9071 35135 9091
rect 34407 8970 34426 8990
rect 34484 8970 34503 8990
rect 34223 8831 34268 8870
rect 33850 8756 33875 8776
rect 33898 8757 33930 8777
rect 34088 8707 34108 8727
rect 33356 8640 33385 8667
rect 33430 8643 33459 8670
rect 30848 8458 30874 8484
rect 31680 8475 31729 8517
rect 31015 8400 31036 8430
rect 30384 8267 30413 8294
rect 30458 8270 30487 8297
rect 31226 8371 31247 8391
rect 31681 8412 31730 8454
rect 33158 8447 33198 8484
rect 33644 8542 33665 8562
rect 33855 8503 33876 8533
rect 34017 8449 34043 8475
rect 31432 8263 31461 8290
rect 31506 8266 31535 8293
rect 29735 8210 29755 8230
rect 33162 8407 33198 8428
rect 29917 8128 29942 8166
rect 29961 8131 29986 8166
rect 30783 8206 30803 8226
rect 30967 8129 30992 8167
rect 31011 8132 31036 8167
rect 33642 8393 33663 8413
rect 34067 8396 34087 8416
rect 33359 8295 33378 8315
rect 33436 8295 33455 8315
rect 33154 8195 33191 8236
rect 33210 8197 33247 8238
rect 34213 8494 34253 8520
rect 34217 8441 34257 8467
rect 34220 8396 34260 8422
rect 27242 7552 27268 7578
rect 28052 7558 28076 7582
rect 28109 7559 28133 7583
rect 27409 7494 27430 7524
rect 27620 7465 27641 7485
rect 29334 7999 29378 8027
rect 29529 8021 29566 8069
rect 29331 7942 29375 7970
rect 27826 7357 27855 7384
rect 27900 7360 27929 7387
rect 27177 7300 27197 7320
rect 26939 4902 26964 4928
rect 27328 4833 27348 4853
rect 26596 4766 26625 4793
rect 26670 4769 26699 4796
rect 26884 4668 26905 4688
rect 27095 4629 27116 4659
rect 27257 4575 27283 4601
rect 26882 4519 26903 4539
rect 27086 4521 27119 4541
rect 27307 4522 27327 4542
rect 26599 4421 26618 4441
rect 26676 4421 26695 4441
rect 27407 4364 27430 4402
rect 28666 6525 28694 6553
rect 28938 6261 28957 6281
rect 29015 6261 29034 6281
rect 28306 6160 28326 6180
rect 28730 6163 28751 6183
rect 28350 6101 28376 6127
rect 29155 6118 29181 6141
rect 28517 6043 28538 6073
rect 28728 6014 28749 6034
rect 28934 5906 28963 5933
rect 29008 5909 29037 5936
rect 28285 5849 28305 5869
rect 28517 5779 28534 5816
rect 28667 5087 28692 5125
rect 28896 4739 28915 4759
rect 28973 4739 28992 4759
rect 28264 4638 28284 4658
rect 28688 4641 28709 4661
rect 30631 7895 30677 7943
rect 34211 8075 34257 8123
rect 36179 11357 36200 11377
rect 36604 11360 36624 11380
rect 35896 11259 35915 11279
rect 35973 11259 35992 11279
rect 36196 10893 36221 10931
rect 36354 10202 36371 10239
rect 36583 10149 36603 10169
rect 35851 10082 35880 10109
rect 35925 10085 35954 10112
rect 36139 9984 36160 10004
rect 36350 9945 36371 9975
rect 35707 9877 35733 9900
rect 36512 9891 36538 9917
rect 36137 9835 36158 9855
rect 36562 9838 36582 9858
rect 35854 9737 35873 9757
rect 35931 9737 35950 9757
rect 36194 9465 36222 9493
rect 37691 8698 37711 8718
rect 36959 8631 36988 8658
rect 37033 8634 37062 8661
rect 37247 8533 37268 8553
rect 37458 8494 37479 8524
rect 36755 8435 36779 8459
rect 36812 8436 36836 8460
rect 37620 8440 37646 8466
rect 37245 8384 37266 8404
rect 37458 8382 37482 8404
rect 37670 8387 37690 8407
rect 36962 8286 36981 8306
rect 37039 8286 37058 8306
rect 41341 13553 41381 13579
rect 41345 13500 41385 13526
rect 42351 13782 42388 13823
rect 42407 13784 42444 13825
rect 42143 13705 42162 13725
rect 42220 13705 42239 13725
rect 41511 13604 41531 13624
rect 41935 13607 41956 13627
rect 42400 13592 42436 13613
rect 41555 13545 41581 13571
rect 41722 13487 41743 13517
rect 41933 13458 41954 13478
rect 42400 13536 42440 13573
rect 42139 13350 42168 13377
rect 42213 13353 42242 13380
rect 41490 13293 41510 13313
rect 41668 13243 41700 13263
rect 41723 13244 41748 13264
rect 41330 13150 41375 13189
rect 41095 13030 41114 13050
rect 41172 13030 41191 13050
rect 40463 12929 40483 12949
rect 40887 12932 40908 12952
rect 40507 12870 40533 12896
rect 41339 12893 41392 12926
rect 40674 12812 40695 12842
rect 40885 12783 40906 12803
rect 41344 12835 41397 12868
rect 42386 13119 42426 13152
rect 42143 13026 42162 13046
rect 42220 13026 42239 13046
rect 41511 12925 41531 12945
rect 41935 12928 41956 12948
rect 41555 12866 41581 12892
rect 42387 12883 42436 12925
rect 41722 12808 41743 12838
rect 41091 12675 41120 12702
rect 41165 12678 41194 12705
rect 41933 12779 41954 12799
rect 42388 12820 42437 12862
rect 42139 12671 42168 12698
rect 42213 12674 42242 12701
rect 40442 12618 40462 12638
rect 41490 12614 41510 12634
rect 39376 12527 39404 12555
rect 41674 12537 41699 12575
rect 41718 12540 41743 12575
rect 41349 12436 41379 12502
rect 39648 12263 39667 12283
rect 39725 12263 39744 12283
rect 39016 12162 39036 12182
rect 39440 12165 39461 12185
rect 39060 12103 39086 12129
rect 39865 12120 39891 12143
rect 40245 12113 40271 12136
rect 39227 12045 39248 12075
rect 39438 12016 39459 12036
rect 41338 12151 41378 12177
rect 41341 12106 41381 12132
rect 41345 12053 41385 12079
rect 39644 11908 39673 11935
rect 39718 11911 39747 11938
rect 38995 11851 39015 11871
rect 39227 11781 39244 11818
rect 42351 12335 42388 12376
rect 42407 12337 42444 12378
rect 42143 12258 42162 12278
rect 42220 12258 42239 12278
rect 41511 12157 41531 12177
rect 41935 12160 41956 12180
rect 42400 12145 42436 12166
rect 41555 12098 41581 12124
rect 41722 12040 41743 12070
rect 41933 12011 41954 12031
rect 42400 12089 42440 12126
rect 42139 11903 42168 11930
rect 42213 11906 42242 11933
rect 41490 11846 41510 11866
rect 41668 11796 41700 11816
rect 41723 11797 41748 11817
rect 39377 11089 39402 11127
rect 41330 11703 41375 11742
rect 41095 11583 41114 11603
rect 41172 11583 41191 11603
rect 40463 11482 40483 11502
rect 40887 11485 40908 11505
rect 40507 11423 40533 11449
rect 41339 11446 41392 11479
rect 40674 11365 40695 11395
rect 40885 11336 40906 11356
rect 41344 11388 41397 11421
rect 42386 11672 42426 11705
rect 42143 11579 42162 11599
rect 42220 11579 42239 11599
rect 41511 11478 41531 11498
rect 41935 11481 41956 11501
rect 41555 11419 41581 11445
rect 42387 11436 42436 11478
rect 41722 11361 41743 11391
rect 41091 11228 41120 11255
rect 41165 11231 41194 11258
rect 41933 11332 41954 11352
rect 42388 11373 42437 11415
rect 42139 11224 42168 11251
rect 42213 11227 42242 11254
rect 40442 11171 40462 11191
rect 41490 11167 41510 11187
rect 41674 11090 41699 11128
rect 41718 11093 41743 11128
rect 41338 10937 41392 11003
rect 39606 10741 39625 10761
rect 39683 10741 39702 10761
rect 38974 10640 38994 10660
rect 39398 10643 39419 10663
rect 39018 10581 39044 10607
rect 39185 10523 39206 10553
rect 39396 10494 39417 10514
rect 39602 10386 39631 10413
rect 39676 10389 39705 10416
rect 38953 10329 38973 10349
rect 41343 10880 41387 10917
rect 41339 10631 41379 10657
rect 41342 10586 41382 10612
rect 41346 10533 41386 10559
rect 42352 10815 42389 10856
rect 42408 10817 42445 10858
rect 42144 10738 42163 10758
rect 42221 10738 42240 10758
rect 41512 10637 41532 10657
rect 41936 10640 41957 10660
rect 42401 10625 42437 10646
rect 41556 10578 41582 10604
rect 41723 10520 41744 10550
rect 41934 10491 41955 10511
rect 42401 10569 42441 10606
rect 42140 10383 42169 10410
rect 42214 10386 42243 10413
rect 41491 10326 41511 10346
rect 41669 10276 41701 10296
rect 41724 10277 41749 10297
rect 39182 9612 39206 9635
rect 39182 9568 39206 9591
rect 39400 9569 39425 9607
rect 39444 9572 39469 9607
rect 39186 9388 39238 9406
rect 39017 9195 39037 9215
rect 39649 9296 39668 9316
rect 39726 9296 39745 9316
rect 41331 10183 41376 10222
rect 41096 10063 41115 10083
rect 41173 10063 41192 10083
rect 40464 9962 40484 9982
rect 40888 9965 40909 9985
rect 40508 9903 40534 9929
rect 41340 9926 41393 9959
rect 40675 9845 40696 9875
rect 40886 9816 40907 9836
rect 41345 9868 41398 9901
rect 42387 10152 42427 10185
rect 42144 10059 42163 10079
rect 42221 10059 42240 10079
rect 41512 9958 41532 9978
rect 41936 9961 41957 9981
rect 41556 9899 41582 9925
rect 42388 9916 42437 9958
rect 41723 9841 41744 9871
rect 41092 9708 41121 9735
rect 41166 9711 41195 9738
rect 41934 9812 41955 9832
rect 42389 9853 42438 9895
rect 42140 9704 42169 9731
rect 42214 9707 42243 9734
rect 40443 9651 40463 9671
rect 41491 9647 41511 9667
rect 41675 9570 41700 9608
rect 41719 9573 41744 9608
rect 41350 9469 41380 9535
rect 39441 9198 39462 9218
rect 39061 9136 39087 9162
rect 40053 9168 40107 9209
rect 39228 9078 39249 9108
rect 39439 9049 39460 9069
rect 41339 9184 41379 9210
rect 41342 9139 41382 9165
rect 41346 9086 41386 9112
rect 42352 9368 42389 9409
rect 42408 9370 42445 9411
rect 42144 9291 42163 9311
rect 42221 9291 42240 9311
rect 41512 9190 41532 9210
rect 41936 9193 41957 9213
rect 42401 9178 42437 9199
rect 41556 9131 41582 9157
rect 41723 9073 41744 9103
rect 39645 8941 39674 8968
rect 39719 8944 39748 8971
rect 38996 8884 39016 8904
rect 37298 8193 37327 8227
rect 37297 8133 37326 8167
rect 35513 8048 35557 8076
rect 35322 7949 35359 7997
rect 35510 7991 35554 8019
rect 30628 7596 30668 7622
rect 30631 7551 30671 7577
rect 30635 7498 30675 7524
rect 37805 7909 37868 7963
rect 31641 7780 31678 7821
rect 31697 7782 31734 7823
rect 31433 7703 31452 7723
rect 31510 7703 31529 7723
rect 30801 7602 30821 7622
rect 31225 7605 31246 7625
rect 33852 7851 33877 7886
rect 33896 7851 33921 7889
rect 34085 7792 34105 7812
rect 34902 7852 34927 7887
rect 34946 7852 34971 7890
rect 31690 7590 31726 7611
rect 35133 7788 35153 7808
rect 33353 7725 33382 7752
rect 33427 7728 33456 7755
rect 30845 7543 30871 7569
rect 31012 7485 31033 7515
rect 31223 7456 31244 7476
rect 31690 7534 31730 7571
rect 33158 7564 33207 7606
rect 33641 7627 33662 7647
rect 34401 7721 34430 7748
rect 34475 7724 34504 7751
rect 33852 7588 33873 7618
rect 33159 7501 33208 7543
rect 34014 7534 34040 7560
rect 31429 7348 31458 7375
rect 31503 7351 31532 7378
rect 30780 7291 30800 7311
rect 30958 7241 30990 7261
rect 31013 7242 31038 7262
rect 30620 7148 30665 7187
rect 30385 7028 30404 7048
rect 30462 7028 30481 7048
rect 29753 6927 29773 6947
rect 30177 6930 30198 6950
rect 29797 6868 29823 6894
rect 30629 6891 30682 6924
rect 29964 6810 29985 6840
rect 30175 6781 30196 6801
rect 30634 6833 30687 6866
rect 31676 7117 31716 7150
rect 31433 7024 31452 7044
rect 31510 7024 31529 7044
rect 30801 6923 30821 6943
rect 31225 6926 31246 6946
rect 33639 7478 33660 7498
rect 34064 7481 34084 7501
rect 33356 7380 33375 7400
rect 33433 7380 33452 7400
rect 33169 7274 33209 7307
rect 34198 7558 34251 7591
rect 34689 7623 34710 7643
rect 34900 7584 34921 7614
rect 34203 7500 34256 7533
rect 35062 7530 35088 7556
rect 34687 7474 34708 7494
rect 35112 7477 35132 7497
rect 34404 7376 34423 7396
rect 34481 7376 34500 7396
rect 34220 7237 34265 7276
rect 35323 7537 35357 7576
rect 33847 7162 33872 7182
rect 33895 7163 33927 7183
rect 34085 7113 34105 7133
rect 33353 7046 33382 7073
rect 33427 7049 33456 7076
rect 30845 6864 30871 6890
rect 31677 6881 31726 6923
rect 31012 6806 31033 6836
rect 30381 6673 30410 6700
rect 30455 6676 30484 6703
rect 31223 6777 31244 6797
rect 31678 6818 31727 6860
rect 33155 6853 33195 6890
rect 33641 6948 33662 6968
rect 35500 7557 35536 7598
rect 35489 7217 35549 7261
rect 36580 7108 36600 7128
rect 35848 7041 35877 7068
rect 35922 7044 35951 7071
rect 33852 6909 33873 6939
rect 34014 6855 34040 6881
rect 31429 6669 31458 6696
rect 31503 6672 31532 6699
rect 29732 6616 29752 6636
rect 33159 6813 33195 6834
rect 30780 6612 30800 6632
rect 30964 6535 30989 6573
rect 31008 6538 31033 6573
rect 33639 6799 33660 6819
rect 34064 6802 34084 6822
rect 33356 6701 33375 6721
rect 33433 6701 33452 6721
rect 33151 6601 33188 6642
rect 33207 6603 33244 6644
rect 34210 6900 34250 6926
rect 34214 6847 34254 6873
rect 34217 6802 34257 6828
rect 30639 6434 30669 6500
rect 36136 6943 36157 6963
rect 36347 6904 36368 6934
rect 35489 6803 35543 6844
rect 36509 6850 36535 6876
rect 36134 6794 36155 6814
rect 34216 6477 34246 6543
rect 29535 6111 29561 6134
rect 30628 6149 30668 6175
rect 30631 6104 30671 6130
rect 30635 6051 30675 6077
rect 31641 6333 31678 6374
rect 31697 6335 31734 6376
rect 31433 6256 31452 6276
rect 31510 6256 31529 6276
rect 30801 6155 30821 6175
rect 31225 6158 31246 6178
rect 33852 6404 33877 6439
rect 33896 6404 33921 6442
rect 34085 6345 34105 6365
rect 31690 6143 31726 6164
rect 35133 6341 35153 6361
rect 33353 6278 33382 6305
rect 33427 6281 33456 6308
rect 30845 6096 30871 6122
rect 31012 6038 31033 6068
rect 31223 6009 31244 6029
rect 31690 6087 31730 6124
rect 33158 6117 33207 6159
rect 33641 6180 33662 6200
rect 34401 6274 34430 6301
rect 34475 6277 34504 6304
rect 33852 6141 33873 6171
rect 33159 6054 33208 6096
rect 34014 6087 34040 6113
rect 31429 5901 31458 5928
rect 31503 5904 31532 5931
rect 30780 5844 30800 5864
rect 30958 5794 30990 5814
rect 31013 5795 31038 5815
rect 30620 5701 30665 5740
rect 30385 5581 30404 5601
rect 30462 5581 30481 5601
rect 29753 5480 29773 5500
rect 30177 5483 30198 5503
rect 29797 5421 29823 5447
rect 30629 5444 30682 5477
rect 29964 5363 29985 5393
rect 30175 5334 30196 5354
rect 30634 5386 30687 5419
rect 31676 5670 31716 5703
rect 31433 5577 31452 5597
rect 31510 5577 31529 5597
rect 30801 5476 30821 5496
rect 31225 5479 31246 5499
rect 33639 6031 33660 6051
rect 34064 6034 34084 6054
rect 33356 5933 33375 5953
rect 33433 5933 33452 5953
rect 33169 5827 33209 5860
rect 34198 6111 34251 6144
rect 34689 6176 34710 6196
rect 34900 6137 34921 6167
rect 34203 6053 34256 6086
rect 35062 6083 35088 6109
rect 34687 6027 34708 6047
rect 35112 6030 35132 6050
rect 34404 5929 34423 5949
rect 34481 5929 34500 5949
rect 34220 5790 34265 5829
rect 35851 6696 35870 6716
rect 35928 6696 35947 6716
rect 36559 6797 36579 6817
rect 36358 6606 36410 6624
rect 36127 6405 36152 6440
rect 36171 6405 36196 6443
rect 36390 6421 36414 6444
rect 36390 6377 36414 6400
rect 33847 5715 33872 5735
rect 33895 5716 33927 5736
rect 34085 5666 34105 5686
rect 33353 5599 33382 5626
rect 33427 5602 33456 5629
rect 30845 5417 30871 5443
rect 31677 5434 31726 5476
rect 31012 5359 31033 5389
rect 30381 5226 30410 5253
rect 30455 5229 30484 5256
rect 31223 5330 31244 5350
rect 31678 5371 31727 5413
rect 33155 5406 33195 5443
rect 33641 5501 33662 5521
rect 33852 5462 33873 5492
rect 34014 5408 34040 5434
rect 31429 5222 31458 5249
rect 31503 5225 31532 5252
rect 29732 5169 29752 5189
rect 33159 5366 33195 5387
rect 30780 5165 30800 5185
rect 30964 5088 30989 5126
rect 31008 5091 31033 5126
rect 33639 5352 33660 5372
rect 34064 5355 34084 5375
rect 33356 5254 33375 5274
rect 33433 5254 33452 5274
rect 33151 5154 33188 5195
rect 33207 5156 33244 5197
rect 34210 5453 34250 5479
rect 34214 5400 34254 5426
rect 34217 5355 34257 5381
rect 34209 5095 34253 5132
rect 36623 5663 36643 5683
rect 35891 5596 35920 5623
rect 35965 5599 35994 5626
rect 36179 5498 36200 5518
rect 36390 5459 36411 5489
rect 36552 5405 36578 5431
rect 30628 4935 30682 5001
rect 34204 5009 34258 5075
rect 28308 4579 28334 4605
rect 28475 4521 28496 4551
rect 28686 4492 28707 4512
rect 28892 4384 28921 4411
rect 28966 4387 28995 4414
rect 28243 4327 28263 4347
rect 25644 4200 25661 4237
rect 28430 4226 28450 4247
rect 28471 4231 28491 4252
rect 25873 4147 25893 4167
rect 25141 4080 25170 4107
rect 25215 4083 25244 4110
rect 25429 3982 25450 4002
rect 25640 3943 25661 3973
rect 24997 3875 25023 3898
rect 25802 3889 25828 3915
rect 25427 3833 25448 3853
rect 25852 3836 25872 3856
rect 25144 3735 25163 3755
rect 25221 3735 25240 3755
rect 30633 4878 30677 4915
rect 30629 4629 30669 4655
rect 30632 4584 30672 4610
rect 30636 4531 30676 4557
rect 31642 4813 31679 4854
rect 31698 4815 31735 4856
rect 31434 4736 31453 4756
rect 31511 4736 31530 4756
rect 30802 4635 30822 4655
rect 31226 4638 31247 4658
rect 33853 4884 33878 4919
rect 33897 4884 33922 4922
rect 34086 4825 34106 4845
rect 31691 4623 31727 4644
rect 35134 4821 35154 4841
rect 33354 4758 33383 4785
rect 33428 4761 33457 4788
rect 30846 4576 30872 4602
rect 31013 4518 31034 4548
rect 31224 4489 31245 4509
rect 31691 4567 31731 4604
rect 33159 4597 33208 4639
rect 33642 4660 33663 4680
rect 34402 4754 34431 4781
rect 34476 4757 34505 4784
rect 33853 4621 33874 4651
rect 33160 4534 33209 4576
rect 34015 4567 34041 4593
rect 31430 4381 31459 4408
rect 31504 4384 31533 4411
rect 30781 4324 30801 4344
rect 30959 4274 30991 4294
rect 31014 4275 31039 4295
rect 28472 3610 28496 3633
rect 28472 3566 28496 3589
rect 28690 3567 28715 3605
rect 28734 3570 28759 3605
rect 25484 3463 25512 3491
rect 28476 3386 28528 3404
rect 28307 3193 28327 3213
rect 28939 3294 28958 3314
rect 29016 3294 29035 3314
rect 30621 4181 30666 4220
rect 30386 4061 30405 4081
rect 30463 4061 30482 4081
rect 29754 3960 29774 3980
rect 30178 3963 30199 3983
rect 29798 3901 29824 3927
rect 30630 3924 30683 3957
rect 29965 3843 29986 3873
rect 30176 3814 30197 3834
rect 30635 3866 30688 3899
rect 31677 4150 31717 4183
rect 31434 4057 31453 4077
rect 31511 4057 31530 4077
rect 30802 3956 30822 3976
rect 31226 3959 31247 3979
rect 33640 4511 33661 4531
rect 34065 4514 34085 4534
rect 33357 4413 33376 4433
rect 33434 4413 33453 4433
rect 33170 4307 33210 4340
rect 34199 4591 34252 4624
rect 34690 4656 34711 4676
rect 34901 4617 34922 4647
rect 34204 4533 34257 4566
rect 35063 4563 35089 4589
rect 34688 4507 34709 4527
rect 35113 4510 35133 4530
rect 34405 4409 34424 4429
rect 34482 4409 34501 4429
rect 34221 4270 34266 4309
rect 33848 4195 33873 4215
rect 33896 4196 33928 4216
rect 34086 4146 34106 4166
rect 33354 4079 33383 4106
rect 33428 4082 33457 4109
rect 30846 3897 30872 3923
rect 31678 3914 31727 3956
rect 31013 3839 31034 3869
rect 30382 3706 30411 3733
rect 30456 3709 30485 3736
rect 31224 3810 31245 3830
rect 31679 3851 31728 3893
rect 33156 3886 33196 3923
rect 33642 3981 33663 4001
rect 33853 3942 33874 3972
rect 34015 3888 34041 3914
rect 31430 3702 31459 3729
rect 31504 3705 31533 3732
rect 29733 3649 29753 3669
rect 33160 3846 33196 3867
rect 30781 3645 30801 3665
rect 30965 3568 30990 3606
rect 31009 3571 31034 3606
rect 33640 3832 33661 3852
rect 34065 3835 34085 3855
rect 33357 3734 33376 3754
rect 33434 3734 33453 3754
rect 33152 3634 33189 3675
rect 33208 3636 33245 3677
rect 34211 3933 34251 3959
rect 34215 3880 34255 3906
rect 34218 3835 34258 3861
rect 35280 3866 35305 3897
rect 35325 3876 35351 3899
rect 30640 3467 30670 3533
rect 28731 3196 28752 3216
rect 28351 3134 28377 3160
rect 29343 3166 29397 3207
rect 28518 3076 28539 3106
rect 28729 3047 28750 3067
rect 34217 3510 34247 3576
rect 30629 3182 30669 3208
rect 30632 3137 30672 3163
rect 30636 3084 30676 3110
rect 31642 3366 31679 3407
rect 31698 3368 31735 3409
rect 31434 3289 31453 3309
rect 31511 3289 31530 3309
rect 30802 3188 30822 3208
rect 31226 3191 31247 3211
rect 33853 3437 33878 3472
rect 33897 3437 33922 3475
rect 34086 3378 34106 3398
rect 31691 3176 31727 3197
rect 35134 3374 35154 3394
rect 33354 3311 33383 3338
rect 33428 3314 33457 3341
rect 30846 3129 30872 3155
rect 31013 3071 31034 3101
rect 28935 2939 28964 2966
rect 29009 2942 29038 2969
rect 28286 2882 28306 2902
rect 27626 2408 27757 2473
rect 29337 2749 29397 2793
rect 29350 2412 29386 2453
rect 31224 3042 31245 3062
rect 31691 3120 31731 3157
rect 33159 3150 33208 3192
rect 33642 3213 33663 3233
rect 34402 3307 34431 3334
rect 34476 3310 34505 3337
rect 33853 3174 33874 3204
rect 33160 3087 33209 3129
rect 34015 3120 34041 3146
rect 31430 2934 31459 2961
rect 31504 2937 31533 2964
rect 30781 2877 30801 2897
rect 30959 2827 30991 2847
rect 31014 2828 31039 2848
rect 29529 2434 29563 2473
rect 30621 2734 30666 2773
rect 30386 2614 30405 2634
rect 30463 2614 30482 2634
rect 29754 2513 29774 2533
rect 30178 2516 30199 2536
rect 29798 2454 29824 2480
rect 30630 2477 30683 2510
rect 24559 2181 24659 2288
rect 29965 2396 29986 2426
rect 30176 2367 30197 2387
rect 30635 2419 30688 2452
rect 31677 2703 31717 2736
rect 31434 2610 31453 2630
rect 31511 2610 31530 2630
rect 30802 2509 30822 2529
rect 31226 2512 31247 2532
rect 33640 3064 33661 3084
rect 34065 3067 34085 3087
rect 33357 2966 33376 2986
rect 33434 2966 33453 2986
rect 33170 2860 33210 2893
rect 34199 3144 34252 3177
rect 34690 3209 34711 3229
rect 34901 3170 34922 3200
rect 34204 3086 34257 3119
rect 35063 3116 35089 3142
rect 34688 3060 34709 3080
rect 35113 3063 35133 3083
rect 34405 2962 34424 2982
rect 34482 2962 34501 2982
rect 34221 2823 34266 2862
rect 33848 2748 33873 2768
rect 33896 2749 33928 2769
rect 34086 2699 34106 2719
rect 33354 2632 33383 2659
rect 33428 2635 33457 2662
rect 30846 2450 30872 2476
rect 31678 2467 31727 2509
rect 31013 2392 31034 2422
rect 30382 2259 30411 2286
rect 30456 2262 30485 2289
rect 31224 2363 31245 2383
rect 31679 2404 31728 2446
rect 33156 2439 33196 2476
rect 33642 2534 33663 2554
rect 33853 2495 33874 2525
rect 34015 2441 34041 2467
rect 31430 2255 31459 2282
rect 31504 2258 31533 2285
rect 29733 2202 29753 2222
rect 33160 2399 33196 2420
rect 29915 2120 29940 2158
rect 29959 2123 29984 2158
rect 30781 2198 30801 2218
rect 30965 2121 30990 2159
rect 31009 2124 31034 2159
rect 33640 2385 33661 2405
rect 34065 2388 34085 2408
rect 33357 2287 33376 2307
rect 33434 2287 33453 2307
rect 33152 2187 33189 2228
rect 33208 2189 33245 2230
rect 36177 5349 36198 5369
rect 36602 5352 36622 5372
rect 35894 5251 35913 5271
rect 35971 5251 35990 5271
rect 36194 4885 36219 4923
rect 38270 7845 38299 7879
rect 38269 7785 38298 7819
rect 38538 7706 38557 7726
rect 38615 7706 38634 7726
rect 37906 7605 37926 7625
rect 38330 7608 38351 7628
rect 40047 8751 40107 8795
rect 40060 8414 40096 8455
rect 41934 9044 41955 9064
rect 42401 9122 42441 9159
rect 42140 8936 42169 8963
rect 42214 8939 42243 8966
rect 41491 8879 41511 8899
rect 41669 8829 41701 8849
rect 41724 8830 41749 8850
rect 40239 8436 40273 8475
rect 41331 8736 41376 8775
rect 41096 8616 41115 8636
rect 41173 8616 41192 8636
rect 40464 8515 40484 8535
rect 40888 8518 40909 8538
rect 40508 8456 40534 8482
rect 41340 8479 41393 8512
rect 40675 8398 40696 8428
rect 40886 8369 40907 8389
rect 41345 8421 41398 8454
rect 42387 8705 42427 8738
rect 42144 8612 42163 8632
rect 42221 8612 42240 8632
rect 41512 8511 41532 8531
rect 41936 8514 41957 8534
rect 41556 8452 41582 8478
rect 42388 8469 42437 8511
rect 41723 8394 41744 8424
rect 41092 8261 41121 8288
rect 41166 8264 41195 8291
rect 41934 8365 41955 8385
rect 42389 8406 42438 8448
rect 42140 8257 42169 8284
rect 42214 8260 42243 8287
rect 40443 8204 40463 8224
rect 40625 8122 40650 8160
rect 40669 8125 40694 8160
rect 41491 8200 41511 8220
rect 41675 8123 41700 8161
rect 41719 8126 41744 8161
rect 37950 7546 37976 7572
rect 38760 7552 38784 7576
rect 38817 7553 38841 7577
rect 38117 7488 38138 7518
rect 38328 7459 38349 7479
rect 40042 7993 40086 8021
rect 40237 8015 40274 8063
rect 40039 7936 40083 7964
rect 38534 7351 38563 7378
rect 38608 7354 38637 7381
rect 37885 7294 37905 7314
rect 37647 4896 37672 4922
rect 38036 4827 38056 4847
rect 37304 4760 37333 4787
rect 37378 4763 37407 4790
rect 37592 4662 37613 4682
rect 37803 4623 37824 4653
rect 37965 4569 37991 4595
rect 37590 4513 37611 4533
rect 37794 4515 37827 4535
rect 38015 4516 38035 4536
rect 37307 4415 37326 4435
rect 37384 4415 37403 4435
rect 38115 4358 38138 4396
rect 39374 6519 39402 6547
rect 39646 6255 39665 6275
rect 39723 6255 39742 6275
rect 39014 6154 39034 6174
rect 39438 6157 39459 6177
rect 39058 6095 39084 6121
rect 39863 6112 39889 6135
rect 39225 6037 39246 6067
rect 39436 6008 39457 6028
rect 39642 5900 39671 5927
rect 39716 5903 39745 5930
rect 38993 5843 39013 5863
rect 39225 5773 39242 5810
rect 39375 5081 39400 5119
rect 39604 4733 39623 4753
rect 39681 4733 39700 4753
rect 38972 4632 38992 4652
rect 39396 4635 39417 4655
rect 41339 7889 41385 7937
rect 41336 7590 41376 7616
rect 41339 7545 41379 7571
rect 41343 7492 41383 7518
rect 42349 7774 42386 7815
rect 42405 7776 42442 7817
rect 42141 7697 42160 7717
rect 42218 7697 42237 7717
rect 41509 7596 41529 7616
rect 41933 7599 41954 7619
rect 42398 7584 42434 7605
rect 41553 7537 41579 7563
rect 41720 7479 41741 7509
rect 41931 7450 41952 7470
rect 42398 7528 42438 7565
rect 42137 7342 42166 7369
rect 42211 7345 42240 7372
rect 41488 7285 41508 7305
rect 41666 7235 41698 7255
rect 41721 7236 41746 7256
rect 41328 7142 41373 7181
rect 41093 7022 41112 7042
rect 41170 7022 41189 7042
rect 40461 6921 40481 6941
rect 40885 6924 40906 6944
rect 40505 6862 40531 6888
rect 41337 6885 41390 6918
rect 40672 6804 40693 6834
rect 40883 6775 40904 6795
rect 41342 6827 41395 6860
rect 42384 7111 42424 7144
rect 42141 7018 42160 7038
rect 42218 7018 42237 7038
rect 41509 6917 41529 6937
rect 41933 6920 41954 6940
rect 41553 6858 41579 6884
rect 42385 6875 42434 6917
rect 41720 6800 41741 6830
rect 41089 6667 41118 6694
rect 41163 6670 41192 6697
rect 41931 6771 41952 6791
rect 42386 6812 42435 6854
rect 42137 6663 42166 6690
rect 42211 6666 42240 6693
rect 40440 6610 40460 6630
rect 41488 6606 41508 6626
rect 41672 6529 41697 6567
rect 41716 6532 41741 6567
rect 41347 6428 41377 6494
rect 40243 6105 40269 6128
rect 41336 6143 41376 6169
rect 41339 6098 41379 6124
rect 41343 6045 41383 6071
rect 42349 6327 42386 6368
rect 42405 6329 42442 6370
rect 42141 6250 42160 6270
rect 42218 6250 42237 6270
rect 41509 6149 41529 6169
rect 41933 6152 41954 6172
rect 42398 6137 42434 6158
rect 41553 6090 41579 6116
rect 41720 6032 41741 6062
rect 41931 6003 41952 6023
rect 42398 6081 42438 6118
rect 42137 5895 42166 5922
rect 42211 5898 42240 5925
rect 41488 5838 41508 5858
rect 41666 5788 41698 5808
rect 41721 5789 41746 5809
rect 41328 5695 41373 5734
rect 41093 5575 41112 5595
rect 41170 5575 41189 5595
rect 40461 5474 40481 5494
rect 40885 5477 40906 5497
rect 40505 5415 40531 5441
rect 41337 5438 41390 5471
rect 40672 5357 40693 5387
rect 40883 5328 40904 5348
rect 41342 5380 41395 5413
rect 42384 5664 42424 5697
rect 42141 5571 42160 5591
rect 42218 5571 42237 5591
rect 41509 5470 41529 5490
rect 41933 5473 41954 5493
rect 41553 5411 41579 5437
rect 42385 5428 42434 5470
rect 41720 5353 41741 5383
rect 41089 5220 41118 5247
rect 41163 5223 41192 5250
rect 41931 5324 41952 5344
rect 42386 5365 42435 5407
rect 42137 5216 42166 5243
rect 42211 5219 42240 5246
rect 40440 5163 40460 5183
rect 41488 5159 41508 5179
rect 41672 5082 41697 5120
rect 41716 5085 41741 5120
rect 41336 4929 41390 4995
rect 39016 4573 39042 4599
rect 39183 4515 39204 4545
rect 39394 4486 39415 4506
rect 39600 4378 39629 4405
rect 39674 4381 39703 4408
rect 38951 4321 38971 4341
rect 36352 4194 36369 4231
rect 39138 4220 39158 4241
rect 39179 4225 39199 4246
rect 36581 4141 36601 4161
rect 35849 4074 35878 4101
rect 35923 4077 35952 4104
rect 36137 3976 36158 3996
rect 36348 3937 36369 3967
rect 35705 3869 35731 3892
rect 36510 3883 36536 3909
rect 36135 3827 36156 3847
rect 36560 3830 36580 3850
rect 35852 3729 35871 3749
rect 35929 3729 35948 3749
rect 41341 4872 41385 4909
rect 41337 4623 41377 4649
rect 41340 4578 41380 4604
rect 41344 4525 41384 4551
rect 42350 4807 42387 4848
rect 42406 4809 42443 4850
rect 42142 4730 42161 4750
rect 42219 4730 42238 4750
rect 41510 4629 41530 4649
rect 41934 4632 41955 4652
rect 42399 4617 42435 4638
rect 41554 4570 41580 4596
rect 41721 4512 41742 4542
rect 41932 4483 41953 4503
rect 42399 4561 42439 4598
rect 42138 4375 42167 4402
rect 42212 4378 42241 4405
rect 41489 4318 41509 4338
rect 41667 4268 41699 4288
rect 41722 4269 41747 4289
rect 39180 3604 39204 3627
rect 39180 3560 39204 3583
rect 39398 3561 39423 3599
rect 39442 3564 39467 3599
rect 36192 3457 36220 3485
rect 39184 3380 39236 3398
rect 39015 3187 39035 3207
rect 39647 3288 39666 3308
rect 39724 3288 39743 3308
rect 41329 4175 41374 4214
rect 41094 4055 41113 4075
rect 41171 4055 41190 4075
rect 40462 3954 40482 3974
rect 40886 3957 40907 3977
rect 40506 3895 40532 3921
rect 41338 3918 41391 3951
rect 40673 3837 40694 3867
rect 40884 3808 40905 3828
rect 41343 3860 41396 3893
rect 42385 4144 42425 4177
rect 42142 4051 42161 4071
rect 42219 4051 42238 4071
rect 41510 3950 41530 3970
rect 41934 3953 41955 3973
rect 41554 3891 41580 3917
rect 42386 3908 42435 3950
rect 41721 3833 41742 3863
rect 41090 3700 41119 3727
rect 41164 3703 41193 3730
rect 41932 3804 41953 3824
rect 42387 3845 42436 3887
rect 42138 3696 42167 3723
rect 42212 3699 42241 3726
rect 40441 3643 40461 3663
rect 41489 3639 41509 3659
rect 41673 3562 41698 3600
rect 41717 3565 41742 3600
rect 41348 3461 41378 3527
rect 39439 3190 39460 3210
rect 39059 3128 39085 3154
rect 40051 3160 40105 3201
rect 39226 3070 39247 3100
rect 39437 3041 39458 3061
rect 41337 3176 41377 3202
rect 41340 3131 41380 3157
rect 41344 3078 41384 3104
rect 42350 3360 42387 3401
rect 42406 3362 42443 3403
rect 42142 3283 42161 3303
rect 42219 3283 42238 3303
rect 41510 3182 41530 3202
rect 41934 3185 41955 3205
rect 42399 3170 42435 3191
rect 41554 3123 41580 3149
rect 41721 3065 41742 3095
rect 39643 2933 39672 2960
rect 39717 2936 39746 2963
rect 38994 2876 39014 2896
rect 38334 2402 38465 2467
rect 40045 2743 40105 2787
rect 40058 2406 40094 2447
rect 41932 3036 41953 3056
rect 42399 3114 42439 3151
rect 42138 2928 42167 2955
rect 42212 2931 42241 2958
rect 41489 2871 41509 2891
rect 41667 2821 41699 2841
rect 41722 2822 41747 2842
rect 40237 2428 40271 2467
rect 41329 2728 41374 2767
rect 41094 2608 41113 2628
rect 41171 2608 41190 2628
rect 40462 2507 40482 2527
rect 40886 2510 40907 2530
rect 40506 2448 40532 2474
rect 41338 2471 41391 2504
rect 35267 2175 35367 2282
rect 40673 2390 40694 2420
rect 40884 2361 40905 2381
rect 41343 2413 41396 2446
rect 42385 2697 42425 2730
rect 42142 2604 42161 2624
rect 42219 2604 42238 2624
rect 41510 2503 41530 2523
rect 41934 2506 41955 2526
rect 41554 2444 41580 2470
rect 42386 2461 42435 2503
rect 41721 2386 41742 2416
rect 41090 2253 41119 2280
rect 41164 2256 41193 2283
rect 41932 2357 41953 2377
rect 42387 2398 42436 2440
rect 42138 2249 42167 2276
rect 42212 2252 42241 2279
rect 40441 2196 40461 2216
rect 40623 2114 40648 2152
rect 40667 2117 40692 2152
rect 41489 2192 41509 2212
rect 41673 2115 41698 2153
rect 41717 2118 41742 2153
rect 10213 729 10289 775
rect 11675 651 11716 699
rect 22334 662 22413 718
rect 31886 727 31962 773
rect 22464 657 22510 708
rect 11416 548 11436 568
rect 10684 481 10713 508
rect 10758 484 10787 511
rect 10187 274 10218 333
rect 10249 274 10280 333
rect 10972 383 10993 403
rect 11183 344 11204 374
rect 11345 290 11371 316
rect 10970 234 10991 254
rect 11184 232 11204 255
rect 11395 237 11415 257
rect 10687 136 10706 156
rect 10764 136 10783 156
rect 20162 547 20203 572
rect 33348 649 33389 697
rect 22053 535 22073 555
rect 33089 546 33109 566
rect 21321 468 21350 495
rect 21395 471 21424 498
rect 20556 266 20753 319
rect 21609 370 21630 390
rect 32357 479 32386 506
rect 32431 482 32460 509
rect 21820 331 21841 361
rect 21982 277 22008 303
rect 21607 221 21628 241
rect 21823 221 21841 243
rect 22032 224 22052 244
rect 21324 123 21343 143
rect 21401 123 21420 143
rect 31860 272 31891 331
rect 31922 272 31953 331
rect 32645 381 32666 401
rect 32856 342 32877 372
rect 33018 288 33044 314
rect 32643 232 32664 252
rect 32857 230 32877 253
rect 33068 235 33088 255
rect 32360 134 32379 154
rect 32437 134 32456 154
rect 22076 13 22105 71
<< metal1 >>
rect 2930 14456 2995 14491
rect 2930 14452 2943 14456
rect 2931 14408 2943 14452
rect 2980 14452 2995 14456
rect 2980 14408 2993 14452
rect 291 13434 398 14224
rect 770 13622 842 14215
rect 1466 13913 1538 13914
rect 1465 13905 1564 13913
rect 1465 13902 1517 13905
rect 1465 13867 1473 13902
rect 1498 13867 1517 13902
rect 1542 13867 1564 13905
rect 1465 13855 1564 13867
rect 1466 13836 1534 13855
rect 1467 13833 1500 13836
rect 1702 13833 1734 13834
rect 877 13772 1080 13785
rect 877 13739 901 13772
rect 937 13771 1080 13772
rect 937 13768 1048 13771
rect 937 13741 974 13768
rect 1003 13744 1048 13768
rect 1077 13744 1080 13771
rect 1003 13741 1080 13744
rect 937 13739 1080 13741
rect 877 13726 1080 13739
rect 877 13725 978 13726
rect 770 13580 779 13622
rect 828 13580 842 13622
rect 770 13559 842 13580
rect 770 13517 780 13559
rect 829 13517 842 13559
rect 770 13499 842 13517
rect 1255 13663 1287 13670
rect 1255 13643 1262 13663
rect 1283 13643 1287 13663
rect 1255 13578 1287 13643
rect 1467 13634 1498 13833
rect 1699 13828 1734 13833
rect 1699 13808 1706 13828
rect 1726 13808 1734 13828
rect 1699 13800 1734 13808
rect 1467 13604 1473 13634
rect 1494 13604 1498 13634
rect 1467 13596 1498 13604
rect 1625 13578 1665 13579
rect 1255 13576 1667 13578
rect 1255 13550 1635 13576
rect 1661 13550 1667 13576
rect 1255 13542 1667 13550
rect 1255 13514 1287 13542
rect 1700 13522 1734 13800
rect 1816 13613 1886 14216
rect 2516 13914 2588 13915
rect 2515 13906 2604 13914
rect 2515 13903 2567 13906
rect 2515 13868 2523 13903
rect 2548 13868 2567 13903
rect 2592 13868 2604 13906
rect 2515 13856 2604 13868
rect 2515 13855 2584 13856
rect 2515 13837 2551 13855
rect 1925 13768 2128 13781
rect 1925 13735 1949 13768
rect 1985 13767 2128 13768
rect 1985 13764 2096 13767
rect 1985 13737 2022 13764
rect 2051 13740 2096 13764
rect 2125 13740 2128 13767
rect 2051 13737 2128 13740
rect 1985 13735 2128 13737
rect 1925 13722 2128 13735
rect 1925 13721 2026 13722
rect 1255 13494 1260 13514
rect 1281 13494 1287 13514
rect 1255 13487 1287 13494
rect 1678 13517 1734 13522
rect 1678 13497 1685 13517
rect 1705 13497 1734 13517
rect 1811 13607 1886 13613
rect 1811 13574 1819 13607
rect 1872 13574 1886 13607
rect 1811 13549 1886 13574
rect 1811 13516 1824 13549
rect 1877 13516 1886 13549
rect 1811 13507 1886 13516
rect 2303 13659 2335 13666
rect 2303 13639 2310 13659
rect 2331 13639 2335 13659
rect 2303 13574 2335 13639
rect 2515 13630 2546 13837
rect 2750 13829 2782 13830
rect 2747 13824 2782 13829
rect 2747 13804 2754 13824
rect 2774 13804 2782 13824
rect 2747 13796 2782 13804
rect 2515 13600 2521 13630
rect 2542 13600 2546 13630
rect 2515 13592 2546 13600
rect 2673 13574 2713 13575
rect 2303 13572 2715 13574
rect 2303 13546 2683 13572
rect 2709 13546 2715 13572
rect 2303 13538 2715 13546
rect 2303 13510 2335 13538
rect 2748 13518 2782 13796
rect 2931 13611 2993 14408
rect 3100 14079 3182 14486
rect 4367 14180 4416 14526
rect 5404 14519 5506 14535
rect 5404 14294 5512 14519
rect 5404 14236 5424 14294
rect 5502 14236 5512 14294
rect 16126 14291 16234 14311
rect 16126 14285 16143 14291
rect 4345 14169 4444 14180
rect 4345 14114 4361 14169
rect 4427 14114 4444 14169
rect 4345 14100 4444 14114
rect 3085 14058 3206 14079
rect 3085 13985 3099 14058
rect 3169 13985 3206 14058
rect 3085 13969 3206 13985
rect 3100 13614 3182 13969
rect 4367 13763 4416 14100
rect 4884 13775 5022 13779
rect 4864 13763 5022 13775
rect 4357 13747 5022 13763
rect 4357 13680 4916 13747
rect 5002 13680 5022 13747
rect 4357 13664 5022 13680
rect 2931 13592 2995 13611
rect 2931 13553 2944 13592
rect 2978 13553 2995 13592
rect 2931 13534 2995 13553
rect 3100 13573 3121 13614
rect 3157 13573 3182 13614
rect 3100 13544 3182 13573
rect 1811 13502 1869 13507
rect 1678 13490 1734 13497
rect 2303 13490 2308 13510
rect 2329 13490 2335 13510
rect 1678 13489 1713 13490
rect 2303 13483 2335 13490
rect 2726 13513 2782 13518
rect 2726 13493 2733 13513
rect 2753 13493 2782 13513
rect 2726 13486 2782 13493
rect 2726 13485 2761 13486
rect 969 13434 1080 13438
rect 2752 13434 3865 13435
rect 291 13416 3865 13434
rect 291 13396 977 13416
rect 996 13396 1054 13416
rect 1073 13412 3865 13416
rect 1073 13396 2025 13412
rect 291 13392 2025 13396
rect 2044 13392 2102 13412
rect 2121 13392 3865 13412
rect 291 13378 3865 13392
rect 291 12755 398 13378
rect 2017 13375 2128 13378
rect 777 13329 841 13333
rect 773 13323 841 13329
rect 773 13290 790 13323
rect 830 13290 841 13323
rect 773 13278 841 13290
rect 1824 13292 1889 13314
rect 773 13276 830 13278
rect 777 12915 828 13276
rect 1824 13253 1841 13292
rect 1886 13253 1889 13292
rect 1465 13208 1500 13210
rect 1465 13199 1569 13208
rect 1465 13198 1516 13199
rect 1465 13178 1468 13198
rect 1493 13179 1516 13198
rect 1548 13179 1569 13199
rect 1493 13178 1569 13179
rect 1465 13171 1569 13178
rect 1465 13159 1500 13171
rect 877 13093 1080 13106
rect 877 13060 901 13093
rect 937 13092 1080 13093
rect 937 13089 1048 13092
rect 937 13062 974 13089
rect 1003 13065 1048 13089
rect 1077 13065 1080 13092
rect 1003 13062 1080 13065
rect 937 13060 1080 13062
rect 877 13047 1080 13060
rect 877 13046 978 13047
rect 1255 12984 1287 12991
rect 1255 12964 1262 12984
rect 1283 12964 1287 12984
rect 766 12906 831 12915
rect 766 12869 776 12906
rect 816 12872 831 12906
rect 1255 12899 1287 12964
rect 1467 12955 1498 13159
rect 1702 13154 1734 13155
rect 1699 13149 1734 13154
rect 1699 13129 1706 13149
rect 1726 13129 1734 13149
rect 1699 13121 1734 13129
rect 1467 12925 1473 12955
rect 1494 12925 1498 12955
rect 1467 12917 1498 12925
rect 1625 12899 1665 12900
rect 1255 12897 1667 12899
rect 816 12869 833 12872
rect 766 12850 833 12869
rect 766 12829 780 12850
rect 816 12829 833 12850
rect 766 12822 833 12829
rect 1255 12871 1635 12897
rect 1661 12871 1667 12897
rect 1255 12863 1667 12871
rect 1255 12835 1287 12863
rect 1700 12843 1734 13121
rect 1824 12953 1889 13253
rect 3095 13277 3188 13292
rect 3095 13233 3110 13277
rect 3170 13233 3188 13277
rect 1255 12815 1260 12835
rect 1281 12815 1287 12835
rect 1255 12808 1287 12815
rect 1678 12838 1734 12843
rect 1678 12818 1685 12838
rect 1705 12818 1734 12838
rect 1678 12811 1734 12818
rect 1814 12942 1894 12953
rect 1814 12916 1831 12942
rect 1871 12916 1894 12942
rect 1814 12889 1894 12916
rect 1814 12863 1835 12889
rect 1875 12863 1894 12889
rect 1814 12844 1894 12863
rect 1814 12818 1838 12844
rect 1878 12818 1894 12844
rect 1678 12810 1713 12811
rect 1814 12806 1894 12818
rect 3095 12860 3188 13233
rect 3372 13088 3575 13101
rect 3372 13055 3396 13088
rect 3432 13087 3575 13088
rect 3432 13084 3543 13087
rect 3432 13057 3469 13084
rect 3498 13060 3543 13084
rect 3572 13060 3575 13087
rect 3498 13057 3575 13060
rect 3432 13055 3575 13057
rect 3372 13042 3575 13055
rect 3372 13041 3473 13042
rect 3095 12819 3110 12860
rect 3164 12819 3188 12860
rect 3095 12812 3188 12819
rect 3750 12979 3782 12986
rect 3750 12959 3757 12979
rect 3778 12959 3782 12979
rect 3750 12894 3782 12959
rect 3962 12950 3993 13151
rect 4197 13149 4229 13150
rect 4194 13144 4229 13149
rect 4194 13124 4201 13144
rect 4221 13124 4229 13144
rect 4194 13116 4229 13124
rect 3962 12920 3968 12950
rect 3989 12920 3993 12950
rect 3962 12912 3993 12920
rect 4120 12894 4160 12895
rect 3750 12892 4162 12894
rect 3750 12866 4130 12892
rect 4156 12866 4162 12892
rect 3750 12858 4162 12866
rect 3750 12830 3782 12858
rect 4195 12838 4229 13116
rect 3750 12810 3755 12830
rect 3776 12810 3782 12830
rect 3750 12803 3782 12810
rect 4173 12833 4229 12838
rect 4173 12813 4180 12833
rect 4200 12813 4229 12833
rect 4173 12806 4229 12813
rect 4173 12805 4208 12806
rect 969 12755 1080 12759
rect 2711 12755 4260 12758
rect 289 12737 4260 12755
rect 289 12717 977 12737
rect 996 12717 1054 12737
rect 1073 12732 4260 12737
rect 1073 12717 3472 12732
rect 289 12712 3472 12717
rect 3491 12712 3549 12732
rect 3568 12712 4260 12732
rect 289 12702 4260 12712
rect 289 12699 914 12702
rect 1101 12699 4260 12702
rect 291 12471 398 12699
rect 2711 12698 4260 12699
rect 3464 12695 3575 12698
rect 759 12660 880 12670
rect 759 12658 828 12660
rect 759 12617 772 12658
rect 809 12619 828 12658
rect 865 12619 880 12660
rect 809 12617 880 12619
rect 759 12599 880 12617
rect 3964 12640 4050 12644
rect 3964 12622 3979 12640
rect 4031 12622 4050 12640
rect 3964 12613 4050 12622
rect 765 12497 844 12599
rect 1817 12559 1884 12578
rect 1817 12539 1837 12559
rect 291 12416 399 12471
rect 766 12416 844 12497
rect 1816 12493 1837 12539
rect 1867 12539 1884 12559
rect 1867 12509 1886 12539
rect 1867 12493 1887 12509
rect 1816 12477 1887 12493
rect 1466 12466 1538 12467
rect 1465 12458 1564 12466
rect 1465 12455 1517 12458
rect 1465 12420 1473 12455
rect 1498 12420 1517 12455
rect 1542 12420 1564 12458
rect 291 11987 398 12416
rect 770 12175 842 12416
rect 1465 12408 1564 12420
rect 1466 12389 1534 12408
rect 1467 12386 1500 12389
rect 1702 12386 1734 12387
rect 877 12325 1080 12338
rect 877 12292 901 12325
rect 937 12324 1080 12325
rect 937 12321 1048 12324
rect 937 12294 974 12321
rect 1003 12297 1048 12321
rect 1077 12297 1080 12324
rect 1003 12294 1080 12297
rect 937 12292 1080 12294
rect 877 12279 1080 12292
rect 877 12278 978 12279
rect 770 12133 779 12175
rect 828 12133 842 12175
rect 770 12112 842 12133
rect 770 12070 780 12112
rect 829 12070 842 12112
rect 770 12052 842 12070
rect 1255 12216 1287 12223
rect 1255 12196 1262 12216
rect 1283 12196 1287 12216
rect 1255 12131 1287 12196
rect 1467 12187 1498 12386
rect 1699 12381 1734 12386
rect 1699 12361 1706 12381
rect 1726 12361 1734 12381
rect 1699 12353 1734 12361
rect 1467 12157 1473 12187
rect 1494 12157 1498 12187
rect 1467 12149 1498 12157
rect 1625 12131 1665 12132
rect 1255 12129 1667 12131
rect 1255 12103 1635 12129
rect 1661 12103 1667 12129
rect 1255 12095 1667 12103
rect 1255 12067 1287 12095
rect 1700 12075 1734 12353
rect 1816 12166 1886 12477
rect 3741 12467 3813 12468
rect 3740 12464 3829 12467
rect 2512 12462 3829 12464
rect 2509 12459 3829 12462
rect 2509 12456 3792 12459
rect 2509 12421 3748 12456
rect 3773 12421 3792 12456
rect 3817 12421 3829 12459
rect 2509 12411 3829 12421
rect 4005 12460 4041 12613
rect 4005 12437 4011 12460
rect 4035 12437 4041 12460
rect 4005 12416 4041 12437
rect 2509 12409 3794 12411
rect 2509 12399 2606 12409
rect 2515 12390 2551 12399
rect 4005 12393 4011 12416
rect 4035 12393 4041 12416
rect 1925 12321 2128 12334
rect 1925 12288 1949 12321
rect 1985 12320 2128 12321
rect 1985 12317 2096 12320
rect 1985 12290 2022 12317
rect 2051 12293 2096 12317
rect 2125 12293 2128 12320
rect 2051 12290 2128 12293
rect 1985 12288 2128 12290
rect 1925 12275 2128 12288
rect 1925 12274 2026 12275
rect 1255 12047 1260 12067
rect 1281 12047 1287 12067
rect 1255 12040 1287 12047
rect 1678 12070 1734 12075
rect 1678 12050 1685 12070
rect 1705 12050 1734 12070
rect 1811 12160 1886 12166
rect 1811 12127 1819 12160
rect 1872 12127 1886 12160
rect 1811 12102 1886 12127
rect 1811 12069 1824 12102
rect 1877 12069 1886 12102
rect 1811 12060 1886 12069
rect 2303 12212 2335 12219
rect 2303 12192 2310 12212
rect 2331 12192 2335 12212
rect 2303 12127 2335 12192
rect 2515 12183 2546 12390
rect 2750 12382 2782 12383
rect 4005 12382 4041 12393
rect 2747 12377 2782 12382
rect 2747 12357 2754 12377
rect 2774 12357 2782 12377
rect 2747 12349 2782 12357
rect 2515 12153 2521 12183
rect 2542 12153 2546 12183
rect 2515 12145 2546 12153
rect 2673 12127 2713 12128
rect 2303 12125 2715 12127
rect 2303 12099 2683 12125
rect 2709 12099 2715 12125
rect 2303 12091 2715 12099
rect 2303 12063 2335 12091
rect 2748 12071 2782 12349
rect 1811 12055 1869 12060
rect 1678 12043 1734 12050
rect 2303 12043 2308 12063
rect 2329 12043 2335 12063
rect 1678 12042 1713 12043
rect 2303 12036 2335 12043
rect 2726 12066 2782 12071
rect 2726 12046 2733 12066
rect 2753 12046 2782 12066
rect 2726 12039 2782 12046
rect 2726 12038 2761 12039
rect 969 11987 1080 11991
rect 2844 11987 4085 11988
rect 291 11969 4085 11987
rect 291 11949 977 11969
rect 996 11949 1054 11969
rect 1073 11965 4085 11969
rect 1073 11949 2025 11965
rect 291 11945 2025 11949
rect 2044 11945 2102 11965
rect 2121 11945 4085 11965
rect 291 11931 4085 11945
rect 291 11308 398 11931
rect 2017 11928 2128 11931
rect 777 11882 841 11886
rect 773 11876 841 11882
rect 773 11843 790 11876
rect 830 11843 841 11876
rect 773 11831 841 11843
rect 1824 11845 1889 11867
rect 773 11829 830 11831
rect 777 11468 828 11829
rect 1824 11806 1841 11845
rect 1886 11806 1889 11845
rect 1465 11761 1500 11763
rect 1465 11752 1569 11761
rect 1465 11751 1516 11752
rect 1465 11731 1468 11751
rect 1493 11732 1516 11751
rect 1548 11732 1569 11752
rect 1493 11731 1569 11732
rect 1465 11724 1569 11731
rect 1465 11712 1500 11724
rect 877 11646 1080 11659
rect 877 11613 901 11646
rect 937 11645 1080 11646
rect 937 11642 1048 11645
rect 937 11615 974 11642
rect 1003 11618 1048 11642
rect 1077 11618 1080 11645
rect 1003 11615 1080 11618
rect 937 11613 1080 11615
rect 877 11600 1080 11613
rect 877 11599 978 11600
rect 1255 11537 1287 11544
rect 1255 11517 1262 11537
rect 1283 11517 1287 11537
rect 766 11459 831 11468
rect 766 11422 776 11459
rect 816 11425 831 11459
rect 1255 11452 1287 11517
rect 1467 11508 1498 11712
rect 1702 11707 1734 11708
rect 1699 11702 1734 11707
rect 1699 11682 1706 11702
rect 1726 11682 1734 11702
rect 1699 11674 1734 11682
rect 1467 11478 1473 11508
rect 1494 11478 1498 11508
rect 1467 11470 1498 11478
rect 1625 11452 1665 11453
rect 1255 11450 1667 11452
rect 816 11422 833 11425
rect 766 11403 833 11422
rect 766 11382 780 11403
rect 816 11382 833 11403
rect 766 11375 833 11382
rect 1255 11424 1635 11450
rect 1661 11424 1667 11450
rect 1255 11416 1667 11424
rect 1255 11388 1287 11416
rect 1700 11396 1734 11674
rect 1824 11506 1889 11806
rect 4003 11800 4108 11809
rect 4003 11795 4057 11800
rect 4003 11774 4016 11795
rect 4036 11779 4057 11795
rect 4077 11779 4108 11800
rect 4036 11774 4108 11779
rect 4003 11743 4108 11774
rect 4006 11726 4041 11743
rect 4005 11708 4041 11726
rect 3415 11643 3618 11656
rect 3415 11610 3439 11643
rect 3475 11642 3618 11643
rect 3475 11639 3586 11642
rect 3475 11612 3512 11639
rect 3541 11615 3586 11639
rect 3615 11615 3618 11642
rect 3541 11612 3618 11615
rect 3475 11610 3618 11612
rect 3415 11597 3618 11610
rect 3415 11596 3516 11597
rect 3793 11534 3825 11541
rect 3793 11514 3800 11534
rect 3821 11514 3825 11534
rect 1255 11368 1260 11388
rect 1281 11368 1287 11388
rect 1255 11361 1287 11368
rect 1678 11391 1734 11396
rect 1678 11371 1685 11391
rect 1705 11371 1734 11391
rect 1678 11364 1734 11371
rect 1814 11495 1894 11506
rect 1814 11469 1831 11495
rect 1871 11469 1894 11495
rect 1814 11442 1894 11469
rect 1814 11416 1835 11442
rect 1875 11416 1894 11442
rect 1814 11397 1894 11416
rect 1814 11371 1838 11397
rect 1878 11371 1894 11397
rect 1678 11363 1713 11364
rect 1814 11359 1894 11371
rect 3793 11449 3825 11514
rect 4005 11505 4036 11708
rect 4240 11704 4272 11705
rect 4237 11699 4272 11704
rect 4237 11679 4244 11699
rect 4264 11679 4272 11699
rect 4237 11671 4272 11679
rect 4005 11475 4011 11505
rect 4032 11475 4036 11505
rect 4005 11467 4036 11475
rect 4163 11449 4203 11450
rect 3793 11447 4205 11449
rect 3793 11421 4173 11447
rect 4199 11421 4205 11447
rect 3793 11413 4205 11421
rect 3793 11385 3825 11413
rect 4238 11393 4272 11671
rect 3793 11365 3798 11385
rect 3819 11365 3825 11385
rect 3793 11358 3825 11365
rect 4216 11388 4272 11393
rect 4216 11368 4223 11388
rect 4243 11368 4272 11388
rect 4216 11361 4272 11368
rect 4216 11360 4251 11361
rect 969 11308 1080 11312
rect 2724 11308 2931 11309
rect 3507 11308 3618 11309
rect 289 11290 4309 11308
rect 289 11270 977 11290
rect 996 11270 1054 11290
rect 1073 11287 4309 11290
rect 1073 11270 3515 11287
rect 289 11267 3515 11270
rect 3534 11267 3592 11287
rect 3611 11267 4309 11287
rect 289 11252 4309 11267
rect 291 11064 398 11252
rect 2886 11250 4309 11252
rect 759 11213 880 11223
rect 759 11211 828 11213
rect 759 11170 772 11211
rect 809 11172 828 11211
rect 865 11172 880 11213
rect 809 11170 880 11172
rect 759 11152 880 11170
rect 291 11060 399 11064
rect 765 11060 842 11152
rect 1815 11148 1891 11164
rect 1815 11125 1830 11148
rect 292 10467 399 11060
rect 767 11009 842 11060
rect 1808 11111 1830 11125
rect 1874 11111 1891 11148
rect 1808 11091 1891 11111
rect 1808 11025 1825 11091
rect 1879 11025 1891 11091
rect 767 10966 843 11009
rect 771 10655 843 10966
rect 1808 11001 1891 11025
rect 1808 10981 1884 11001
rect 1808 10962 1887 10981
rect 1467 10946 1539 10947
rect 1466 10938 1565 10946
rect 1466 10935 1518 10938
rect 1466 10900 1474 10935
rect 1499 10900 1518 10935
rect 1543 10900 1565 10938
rect 1466 10888 1565 10900
rect 1467 10869 1535 10888
rect 1468 10866 1501 10869
rect 1703 10866 1735 10867
rect 878 10805 1081 10818
rect 878 10772 902 10805
rect 938 10804 1081 10805
rect 938 10801 1049 10804
rect 938 10774 975 10801
rect 1004 10777 1049 10801
rect 1078 10777 1081 10804
rect 1004 10774 1081 10777
rect 938 10772 1081 10774
rect 878 10759 1081 10772
rect 878 10758 979 10759
rect 771 10613 780 10655
rect 829 10613 843 10655
rect 771 10592 843 10613
rect 771 10550 781 10592
rect 830 10550 843 10592
rect 771 10532 843 10550
rect 1256 10696 1288 10703
rect 1256 10676 1263 10696
rect 1284 10676 1288 10696
rect 1256 10611 1288 10676
rect 1468 10667 1499 10866
rect 1700 10861 1735 10866
rect 1700 10841 1707 10861
rect 1727 10841 1735 10861
rect 1700 10833 1735 10841
rect 1468 10637 1474 10667
rect 1495 10637 1499 10667
rect 1468 10629 1499 10637
rect 1626 10611 1666 10612
rect 1256 10609 1668 10611
rect 1256 10583 1636 10609
rect 1662 10583 1668 10609
rect 1256 10575 1668 10583
rect 1256 10547 1288 10575
rect 1701 10555 1735 10833
rect 1817 10646 1887 10962
rect 3805 10947 3836 10948
rect 3805 10939 3850 10947
rect 2885 10916 3049 10923
rect 3805 10916 3815 10939
rect 2511 10901 3815 10916
rect 3840 10901 3850 10939
rect 2511 10883 3850 10901
rect 2516 10870 2552 10883
rect 2885 10880 3049 10883
rect 1926 10801 2129 10814
rect 1926 10768 1950 10801
rect 1986 10800 2129 10801
rect 1986 10797 2097 10800
rect 1986 10770 2023 10797
rect 2052 10773 2097 10797
rect 2126 10773 2129 10800
rect 2052 10770 2129 10773
rect 1986 10768 2129 10770
rect 1926 10755 2129 10768
rect 1926 10754 2027 10755
rect 1256 10527 1261 10547
rect 1282 10527 1288 10547
rect 1256 10520 1288 10527
rect 1679 10550 1735 10555
rect 1679 10530 1686 10550
rect 1706 10530 1735 10550
rect 1812 10640 1887 10646
rect 1812 10607 1820 10640
rect 1873 10607 1887 10640
rect 1812 10582 1887 10607
rect 1812 10549 1825 10582
rect 1878 10549 1887 10582
rect 1812 10540 1887 10549
rect 2304 10692 2336 10699
rect 2304 10672 2311 10692
rect 2332 10672 2336 10692
rect 2304 10607 2336 10672
rect 2516 10663 2547 10870
rect 2751 10862 2783 10863
rect 2748 10857 2783 10862
rect 2748 10837 2755 10857
rect 2775 10837 2783 10857
rect 2748 10829 2783 10837
rect 2516 10633 2522 10663
rect 2543 10633 2547 10663
rect 2516 10625 2547 10633
rect 2674 10607 2714 10608
rect 2304 10605 2716 10607
rect 2304 10579 2684 10605
rect 2710 10579 2716 10605
rect 2304 10571 2716 10579
rect 2304 10543 2336 10571
rect 2749 10551 2783 10829
rect 1812 10535 1870 10540
rect 1679 10523 1735 10530
rect 2304 10523 2309 10543
rect 2330 10523 2336 10543
rect 1679 10522 1714 10523
rect 2304 10516 2336 10523
rect 2727 10546 2783 10551
rect 2727 10526 2734 10546
rect 2754 10526 2783 10546
rect 2727 10519 2783 10526
rect 2727 10518 2762 10519
rect 970 10467 1081 10471
rect 2753 10467 4053 10468
rect 292 10449 4053 10467
rect 292 10429 978 10449
rect 997 10429 1055 10449
rect 1074 10445 4053 10449
rect 1074 10429 2026 10445
rect 292 10425 2026 10429
rect 2045 10425 2103 10445
rect 2122 10425 4053 10445
rect 292 10411 4053 10425
rect 292 9788 399 10411
rect 2018 10408 2129 10411
rect 778 10362 842 10366
rect 774 10356 842 10362
rect 774 10323 791 10356
rect 831 10323 842 10356
rect 774 10311 842 10323
rect 1825 10325 1890 10347
rect 774 10309 831 10311
rect 778 9948 829 10309
rect 1825 10286 1842 10325
rect 1887 10286 1890 10325
rect 1466 10241 1501 10243
rect 1466 10232 1570 10241
rect 1466 10231 1517 10232
rect 1466 10211 1469 10231
rect 1494 10212 1517 10231
rect 1549 10212 1570 10232
rect 1494 10211 1570 10212
rect 1466 10204 1570 10211
rect 1466 10192 1501 10204
rect 878 10126 1081 10139
rect 878 10093 902 10126
rect 938 10125 1081 10126
rect 938 10122 1049 10125
rect 938 10095 975 10122
rect 1004 10098 1049 10122
rect 1078 10098 1081 10125
rect 1004 10095 1081 10098
rect 938 10093 1081 10095
rect 878 10080 1081 10093
rect 878 10079 979 10080
rect 1256 10017 1288 10024
rect 1256 9997 1263 10017
rect 1284 9997 1288 10017
rect 767 9939 832 9948
rect 767 9902 777 9939
rect 817 9905 832 9939
rect 1256 9932 1288 9997
rect 1468 9988 1499 10192
rect 1703 10187 1735 10188
rect 1700 10182 1735 10187
rect 1700 10162 1707 10182
rect 1727 10162 1735 10182
rect 1700 10154 1735 10162
rect 1468 9958 1474 9988
rect 1495 9958 1499 9988
rect 1468 9950 1499 9958
rect 1626 9932 1666 9933
rect 1256 9930 1668 9932
rect 817 9902 834 9905
rect 767 9883 834 9902
rect 767 9862 781 9883
rect 817 9862 834 9883
rect 767 9855 834 9862
rect 1256 9904 1636 9930
rect 1662 9904 1668 9930
rect 1256 9896 1668 9904
rect 1256 9868 1288 9896
rect 1701 9876 1735 10154
rect 1825 9986 1890 10286
rect 3962 10247 3999 10268
rect 3962 10210 3973 10247
rect 3990 10223 3999 10247
rect 3990 10210 4000 10223
rect 3962 10200 4000 10210
rect 3963 10196 4000 10200
rect 3963 10190 3996 10196
rect 3373 10121 3576 10134
rect 3373 10088 3397 10121
rect 3433 10120 3576 10121
rect 3433 10117 3544 10120
rect 3433 10090 3470 10117
rect 3499 10093 3544 10117
rect 3573 10093 3576 10120
rect 3499 10090 3576 10093
rect 3433 10088 3576 10090
rect 3373 10075 3576 10088
rect 3373 10074 3474 10075
rect 3751 10012 3783 10019
rect 3751 9992 3758 10012
rect 3779 9992 3783 10012
rect 1256 9848 1261 9868
rect 1282 9848 1288 9868
rect 1256 9841 1288 9848
rect 1679 9871 1735 9876
rect 1679 9851 1686 9871
rect 1706 9851 1735 9871
rect 1679 9844 1735 9851
rect 1815 9975 1895 9986
rect 1815 9949 1832 9975
rect 1872 9949 1895 9975
rect 1815 9922 1895 9949
rect 1815 9896 1836 9922
rect 1876 9896 1895 9922
rect 3751 9927 3783 9992
rect 3963 9983 3994 10190
rect 4198 10182 4230 10183
rect 4195 10177 4230 10182
rect 4195 10157 4202 10177
rect 4222 10157 4230 10177
rect 4195 10149 4230 10157
rect 3963 9953 3969 9983
rect 3990 9953 3994 9983
rect 3963 9945 3994 9953
rect 4121 9927 4161 9928
rect 3751 9925 4163 9927
rect 1815 9877 1895 9896
rect 1815 9851 1839 9877
rect 1879 9851 1895 9877
rect 2928 9915 3365 9921
rect 2928 9892 2946 9915
rect 2972 9908 3365 9915
rect 2972 9892 3326 9908
rect 2928 9885 3326 9892
rect 3352 9885 3365 9908
rect 2928 9872 3365 9885
rect 3751 9899 4131 9925
rect 4157 9899 4163 9925
rect 3751 9891 4163 9899
rect 1679 9843 1714 9844
rect 1815 9839 1895 9851
rect 3751 9863 3783 9891
rect 4196 9871 4230 10149
rect 3751 9843 3756 9863
rect 3777 9843 3783 9863
rect 3751 9836 3783 9843
rect 4174 9866 4230 9871
rect 4174 9846 4181 9866
rect 4201 9846 4230 9866
rect 4174 9839 4230 9846
rect 4174 9838 4209 9839
rect 970 9788 1081 9792
rect 2712 9788 4262 9791
rect 290 9770 4262 9788
rect 290 9750 978 9770
rect 997 9750 1055 9770
rect 1074 9765 4262 9770
rect 1074 9750 3473 9765
rect 290 9745 3473 9750
rect 3492 9745 3550 9765
rect 3569 9745 4262 9765
rect 290 9735 4262 9745
rect 290 9732 915 9735
rect 1102 9732 4262 9735
rect 292 9504 399 9732
rect 2712 9731 4262 9732
rect 3465 9728 3576 9731
rect 760 9693 881 9703
rect 760 9691 829 9693
rect 760 9650 773 9691
rect 810 9652 829 9691
rect 866 9652 881 9693
rect 810 9650 881 9652
rect 760 9632 881 9650
rect 766 9530 845 9632
rect 1818 9592 1885 9611
rect 1818 9572 1838 9592
rect 292 9449 400 9504
rect 767 9449 845 9530
rect 1817 9526 1838 9572
rect 1868 9572 1885 9592
rect 1868 9542 1887 9572
rect 1868 9526 1888 9542
rect 1817 9510 1888 9526
rect 1467 9499 1539 9500
rect 1466 9491 1565 9499
rect 1466 9488 1518 9491
rect 1466 9453 1474 9488
rect 1499 9453 1518 9488
rect 1543 9453 1565 9491
rect 292 9020 399 9449
rect 771 9208 843 9449
rect 1466 9441 1565 9453
rect 1467 9422 1535 9441
rect 1468 9419 1501 9422
rect 1703 9419 1735 9420
rect 878 9358 1081 9371
rect 878 9325 902 9358
rect 938 9357 1081 9358
rect 938 9354 1049 9357
rect 938 9327 975 9354
rect 1004 9330 1049 9354
rect 1078 9330 1081 9357
rect 1004 9327 1081 9330
rect 938 9325 1081 9327
rect 878 9312 1081 9325
rect 878 9311 979 9312
rect 771 9166 780 9208
rect 829 9166 843 9208
rect 771 9145 843 9166
rect 771 9103 781 9145
rect 830 9103 843 9145
rect 771 9085 843 9103
rect 1256 9249 1288 9256
rect 1256 9229 1263 9249
rect 1284 9229 1288 9249
rect 1256 9164 1288 9229
rect 1468 9220 1499 9419
rect 1700 9414 1735 9419
rect 1700 9394 1707 9414
rect 1727 9394 1735 9414
rect 1700 9386 1735 9394
rect 1468 9190 1474 9220
rect 1495 9190 1499 9220
rect 1468 9182 1499 9190
rect 1626 9164 1666 9165
rect 1256 9162 1668 9164
rect 1256 9136 1636 9162
rect 1662 9136 1668 9162
rect 1256 9128 1668 9136
rect 1256 9100 1288 9128
rect 1701 9108 1735 9386
rect 1817 9199 1887 9510
rect 2514 9501 3856 9506
rect 2514 9499 3813 9501
rect 2511 9473 3813 9499
rect 3841 9473 3856 9501
rect 2511 9465 3856 9473
rect 2511 9440 2550 9465
rect 2511 9423 2552 9440
rect 2511 9416 2550 9423
rect 1926 9354 2129 9367
rect 1926 9321 1950 9354
rect 1986 9353 2129 9354
rect 1986 9350 2097 9353
rect 1986 9323 2023 9350
rect 2052 9326 2097 9350
rect 2126 9326 2129 9353
rect 2052 9323 2129 9326
rect 1986 9321 2129 9323
rect 1926 9308 2129 9321
rect 1926 9307 2027 9308
rect 1256 9080 1261 9100
rect 1282 9080 1288 9100
rect 1256 9073 1288 9080
rect 1679 9103 1735 9108
rect 1679 9083 1686 9103
rect 1706 9083 1735 9103
rect 1812 9193 1887 9199
rect 1812 9160 1820 9193
rect 1873 9160 1887 9193
rect 1812 9135 1887 9160
rect 1812 9102 1825 9135
rect 1878 9102 1887 9135
rect 1812 9093 1887 9102
rect 2304 9245 2336 9252
rect 2304 9225 2311 9245
rect 2332 9225 2336 9245
rect 2304 9160 2336 9225
rect 2516 9216 2547 9416
rect 2751 9415 2783 9416
rect 2748 9410 2783 9415
rect 2748 9390 2755 9410
rect 2775 9390 2783 9410
rect 2748 9382 2783 9390
rect 2516 9186 2522 9216
rect 2543 9186 2547 9216
rect 2516 9178 2547 9186
rect 2674 9160 2714 9161
rect 2304 9158 2716 9160
rect 2304 9132 2684 9158
rect 2710 9132 2716 9158
rect 2304 9124 2716 9132
rect 2304 9096 2336 9124
rect 2749 9104 2783 9382
rect 1812 9088 1870 9093
rect 1679 9076 1735 9083
rect 2304 9076 2309 9096
rect 2330 9076 2336 9096
rect 1679 9075 1714 9076
rect 2304 9069 2336 9076
rect 2727 9099 2783 9104
rect 2727 9079 2734 9099
rect 2754 9079 2783 9099
rect 2727 9072 2783 9079
rect 2727 9071 2762 9072
rect 970 9020 1081 9024
rect 2845 9020 3835 9021
rect 292 9002 3835 9020
rect 292 8982 978 9002
rect 997 8982 1055 9002
rect 1074 8998 3835 9002
rect 1074 8982 2026 8998
rect 292 8978 2026 8982
rect 2045 8978 2103 8998
rect 2122 8978 3835 8998
rect 292 8964 3835 8978
rect 292 8341 399 8964
rect 2018 8961 2129 8964
rect 778 8915 842 8919
rect 774 8909 842 8915
rect 774 8876 791 8909
rect 831 8876 842 8909
rect 774 8864 842 8876
rect 1825 8878 1890 8900
rect 774 8862 831 8864
rect 778 8501 829 8862
rect 1825 8839 1842 8878
rect 1887 8839 1890 8878
rect 1466 8794 1501 8796
rect 1466 8785 1570 8794
rect 1466 8784 1517 8785
rect 1466 8764 1469 8784
rect 1494 8765 1517 8784
rect 1549 8765 1570 8785
rect 1494 8764 1570 8765
rect 1466 8757 1570 8764
rect 1466 8745 1501 8757
rect 878 8679 1081 8692
rect 878 8646 902 8679
rect 938 8678 1081 8679
rect 938 8675 1049 8678
rect 938 8648 975 8675
rect 1004 8651 1049 8675
rect 1078 8651 1081 8678
rect 1004 8648 1081 8651
rect 938 8646 1081 8648
rect 878 8633 1081 8646
rect 878 8632 979 8633
rect 1256 8570 1288 8577
rect 1256 8550 1263 8570
rect 1284 8550 1288 8570
rect 767 8492 832 8501
rect 767 8455 777 8492
rect 817 8458 832 8492
rect 1256 8485 1288 8550
rect 1468 8541 1499 8745
rect 1703 8740 1735 8741
rect 1700 8735 1735 8740
rect 1700 8715 1707 8735
rect 1727 8715 1735 8735
rect 1700 8707 1735 8715
rect 1468 8511 1474 8541
rect 1495 8511 1499 8541
rect 1468 8503 1499 8511
rect 1626 8485 1666 8486
rect 1256 8483 1668 8485
rect 817 8455 834 8458
rect 767 8436 834 8455
rect 767 8415 781 8436
rect 817 8415 834 8436
rect 767 8408 834 8415
rect 1256 8457 1636 8483
rect 1662 8457 1668 8483
rect 1256 8449 1668 8457
rect 1256 8421 1288 8449
rect 1701 8429 1735 8707
rect 1825 8539 1890 8839
rect 1256 8401 1261 8421
rect 1282 8401 1288 8421
rect 1256 8394 1288 8401
rect 1679 8424 1735 8429
rect 1679 8404 1686 8424
rect 1706 8404 1735 8424
rect 1679 8397 1735 8404
rect 1815 8528 1895 8539
rect 1815 8502 1832 8528
rect 1872 8502 1895 8528
rect 1815 8475 1895 8502
rect 4367 8478 4416 13664
rect 4864 13661 5022 13664
rect 4884 13653 5022 13661
rect 5404 13106 5512 14236
rect 16123 14233 16143 14285
rect 16221 14233 16234 14291
rect 16123 14220 16234 14233
rect 27077 14292 27185 14320
rect 27077 14234 27097 14292
rect 27175 14234 27185 14292
rect 37799 14289 37907 14309
rect 37799 14283 37816 14289
rect 15066 14152 15153 14170
rect 15066 14108 15083 14152
rect 15135 14108 15153 14152
rect 15066 14091 15153 14108
rect 13808 14048 13889 14049
rect 13802 14034 13901 14048
rect 13802 13984 13822 14034
rect 13874 13984 13901 14034
rect 13802 13964 13901 13984
rect 10005 13851 10070 13934
rect 9955 13833 10076 13851
rect 9955 13831 10026 13833
rect 9955 13790 9970 13831
rect 10007 13792 10026 13831
rect 10063 13792 10076 13833
rect 10007 13790 10076 13792
rect 9955 13780 10076 13790
rect 6471 13751 7949 13753
rect 10436 13751 11113 13775
rect 6471 13746 9631 13751
rect 9889 13746 11113 13751
rect 6471 13733 11113 13746
rect 6471 13713 9762 13733
rect 9781 13713 9839 13733
rect 9858 13713 11113 13733
rect 6471 13695 11113 13713
rect 7904 13694 8111 13695
rect 9755 13691 9866 13695
rect 10436 13687 11113 13695
rect 8941 13632 9021 13644
rect 9122 13639 9157 13640
rect 8941 13606 8957 13632
rect 8997 13606 9021 13632
rect 8941 13587 9021 13606
rect 8941 13561 8960 13587
rect 9000 13561 9021 13587
rect 8941 13534 9021 13561
rect 8941 13508 8964 13534
rect 9004 13508 9021 13534
rect 8941 13497 9021 13508
rect 9101 13632 9157 13639
rect 9101 13612 9130 13632
rect 9150 13612 9157 13632
rect 9101 13607 9157 13612
rect 9548 13635 9580 13642
rect 9548 13615 9554 13635
rect 9575 13615 9580 13635
rect 8946 13197 9011 13497
rect 9101 13329 9135 13607
rect 9548 13587 9580 13615
rect 9168 13579 9580 13587
rect 9168 13553 9174 13579
rect 9200 13553 9580 13579
rect 10002 13621 10069 13628
rect 10002 13600 10019 13621
rect 10055 13600 10069 13621
rect 10002 13581 10069 13600
rect 10002 13578 10019 13581
rect 9168 13551 9580 13553
rect 9170 13550 9210 13551
rect 9337 13525 9368 13533
rect 9337 13495 9341 13525
rect 9362 13495 9368 13525
rect 9101 13321 9136 13329
rect 9101 13301 9109 13321
rect 9129 13301 9136 13321
rect 9101 13296 9136 13301
rect 9101 13295 9133 13296
rect 9337 13291 9368 13495
rect 9548 13486 9580 13551
rect 10004 13544 10019 13578
rect 10059 13544 10069 13581
rect 10004 13535 10069 13544
rect 9548 13466 9552 13486
rect 9573 13466 9580 13486
rect 9548 13459 9580 13466
rect 9857 13403 9958 13404
rect 9755 13390 9958 13403
rect 9755 13388 9898 13390
rect 9755 13385 9832 13388
rect 9755 13358 9758 13385
rect 9787 13361 9832 13385
rect 9861 13361 9898 13388
rect 9787 13358 9898 13361
rect 9755 13357 9898 13358
rect 9934 13357 9958 13390
rect 9755 13344 9958 13357
rect 9335 13279 9370 13291
rect 9266 13272 9370 13279
rect 9266 13271 9342 13272
rect 9266 13251 9287 13271
rect 9319 13252 9342 13271
rect 9367 13252 9370 13272
rect 9319 13251 9370 13252
rect 9266 13242 9370 13251
rect 9335 13240 9370 13242
rect 8946 13158 8949 13197
rect 8994 13158 9011 13197
rect 10007 13174 10058 13535
rect 10005 13172 10062 13174
rect 8946 13136 9011 13158
rect 9994 13160 10062 13172
rect 9994 13127 10005 13160
rect 10045 13127 10062 13160
rect 9994 13121 10062 13127
rect 9994 13117 10058 13121
rect 4481 8670 4684 8683
rect 4481 8637 4505 8670
rect 4541 8669 4684 8670
rect 4541 8666 4652 8669
rect 4541 8639 4578 8666
rect 4607 8642 4652 8666
rect 4681 8642 4684 8669
rect 4607 8639 4684 8642
rect 4541 8637 4684 8639
rect 4481 8624 4684 8637
rect 4481 8623 4582 8624
rect 4859 8561 4891 8568
rect 4859 8541 4866 8561
rect 4887 8541 4891 8561
rect 1815 8449 1836 8475
rect 1876 8449 1895 8475
rect 1815 8430 1895 8449
rect 4366 8468 4477 8478
rect 4366 8467 4431 8468
rect 4366 8443 4374 8467
rect 4398 8444 4431 8467
rect 4455 8444 4477 8468
rect 4398 8443 4477 8444
rect 4366 8436 4477 8443
rect 4859 8476 4891 8541
rect 5071 8532 5102 8732
rect 5306 8731 5338 8732
rect 5303 8726 5338 8731
rect 5303 8706 5310 8726
rect 5330 8706 5338 8726
rect 5303 8698 5338 8706
rect 5071 8502 5077 8532
rect 5098 8502 5102 8532
rect 5071 8494 5102 8502
rect 5229 8476 5269 8477
rect 4859 8474 5271 8476
rect 4859 8448 5239 8474
rect 5265 8448 5271 8474
rect 4859 8440 5271 8448
rect 1815 8404 1839 8430
rect 1879 8404 1895 8430
rect 1679 8396 1714 8397
rect 1815 8392 1895 8404
rect 4859 8412 4891 8440
rect 5304 8420 5338 8698
rect 4859 8392 4864 8412
rect 4885 8392 4891 8412
rect 4859 8385 4891 8392
rect 5070 8412 5104 8419
rect 5070 8390 5077 8412
rect 5101 8390 5104 8412
rect 970 8341 1081 8345
rect 2725 8341 2932 8342
rect 290 8336 4365 8341
rect 290 8323 4684 8336
rect 290 8303 978 8323
rect 997 8303 1055 8323
rect 1074 8314 4684 8323
rect 1074 8303 4581 8314
rect 290 8294 4581 8303
rect 4600 8294 4658 8314
rect 4677 8294 4684 8314
rect 290 8285 4684 8294
rect 292 8112 399 8285
rect 2887 8283 4684 8285
rect 4573 8277 4684 8283
rect 760 8246 881 8256
rect 760 8244 829 8246
rect 760 8203 773 8244
rect 810 8205 829 8244
rect 866 8205 881 8246
rect 810 8203 881 8205
rect 760 8185 881 8203
rect 4908 8235 4960 8266
rect 4908 8201 4917 8235
rect 4946 8201 4960 8235
rect 283 8085 399 8112
rect 766 8093 831 8185
rect 4908 8175 4960 8201
rect 5070 8184 5104 8390
rect 5282 8415 5338 8420
rect 5282 8395 5289 8415
rect 5309 8395 5338 8415
rect 5282 8388 5338 8395
rect 5282 8387 5317 8388
rect 283 7946 394 8085
rect 764 8047 831 8093
rect 1816 8131 1888 8153
rect 1816 8083 1830 8131
rect 1876 8126 1888 8131
rect 4908 8141 4916 8175
rect 4945 8141 4960 8175
rect 1876 8083 1893 8126
rect 764 7946 829 8047
rect 283 7886 396 7946
rect 764 7908 840 7946
rect 289 7426 396 7886
rect 768 7614 840 7908
rect 1464 7905 1536 7906
rect 1463 7897 1562 7905
rect 1816 7900 1893 8083
rect 3104 8084 3188 8095
rect 3104 8056 3132 8084
rect 3176 8056 3188 8084
rect 2918 8005 2992 8033
rect 2918 7957 2941 8005
rect 2978 7957 2992 8005
rect 3104 8027 3188 8056
rect 3104 7999 3129 8027
rect 3173 7999 3188 8027
rect 3104 7966 3188 7999
rect 2918 7948 2992 7957
rect 2514 7906 2586 7907
rect 1463 7894 1515 7897
rect 1463 7859 1471 7894
rect 1496 7859 1515 7894
rect 1540 7859 1562 7897
rect 1463 7847 1562 7859
rect 1814 7871 1893 7900
rect 2513 7898 2602 7906
rect 2513 7895 2565 7898
rect 1464 7828 1532 7847
rect 1465 7825 1498 7828
rect 1700 7825 1732 7826
rect 875 7764 1078 7777
rect 875 7731 899 7764
rect 935 7763 1078 7764
rect 935 7760 1046 7763
rect 935 7733 972 7760
rect 1001 7736 1046 7760
rect 1075 7736 1078 7763
rect 1001 7733 1078 7736
rect 935 7731 1078 7733
rect 875 7718 1078 7731
rect 875 7717 976 7718
rect 768 7572 777 7614
rect 826 7572 840 7614
rect 768 7551 840 7572
rect 768 7509 778 7551
rect 827 7509 840 7551
rect 768 7491 840 7509
rect 1253 7655 1285 7662
rect 1253 7635 1260 7655
rect 1281 7635 1285 7655
rect 1253 7570 1285 7635
rect 1465 7626 1496 7825
rect 1697 7820 1732 7825
rect 1697 7800 1704 7820
rect 1724 7800 1732 7820
rect 1697 7792 1732 7800
rect 1465 7596 1471 7626
rect 1492 7596 1496 7626
rect 1465 7588 1496 7596
rect 1623 7570 1663 7571
rect 1253 7568 1665 7570
rect 1253 7542 1633 7568
rect 1659 7542 1665 7568
rect 1253 7534 1665 7542
rect 1253 7506 1285 7534
rect 1698 7514 1732 7792
rect 1814 7605 1884 7871
rect 2513 7860 2521 7895
rect 2546 7860 2565 7895
rect 2590 7860 2602 7898
rect 2513 7848 2602 7860
rect 2513 7847 2582 7848
rect 2513 7829 2549 7847
rect 1923 7760 2126 7773
rect 1923 7727 1947 7760
rect 1983 7759 2126 7760
rect 1983 7756 2094 7759
rect 1983 7729 2020 7756
rect 2049 7732 2094 7756
rect 2123 7732 2126 7759
rect 2049 7729 2126 7732
rect 1983 7727 2126 7729
rect 1923 7714 2126 7727
rect 1923 7713 2024 7714
rect 1253 7486 1258 7506
rect 1279 7486 1285 7506
rect 1253 7479 1285 7486
rect 1676 7509 1732 7514
rect 1676 7489 1683 7509
rect 1703 7489 1732 7509
rect 1809 7599 1884 7605
rect 1809 7566 1817 7599
rect 1870 7566 1884 7599
rect 1809 7541 1884 7566
rect 1809 7508 1822 7541
rect 1875 7508 1884 7541
rect 1809 7499 1884 7508
rect 2301 7651 2333 7658
rect 2301 7631 2308 7651
rect 2329 7631 2333 7651
rect 2301 7566 2333 7631
rect 2513 7622 2544 7829
rect 2748 7821 2780 7822
rect 2745 7816 2780 7821
rect 2745 7796 2752 7816
rect 2772 7796 2780 7816
rect 2745 7788 2780 7796
rect 2513 7592 2519 7622
rect 2540 7592 2544 7622
rect 2513 7584 2544 7592
rect 2671 7566 2711 7567
rect 2301 7564 2713 7566
rect 2301 7538 2681 7564
rect 2707 7538 2713 7564
rect 2301 7530 2713 7538
rect 2301 7502 2333 7530
rect 2746 7510 2780 7788
rect 2929 7603 2991 7948
rect 3098 7921 3188 7966
rect 3098 7606 3180 7921
rect 2929 7584 2993 7603
rect 2929 7545 2942 7584
rect 2976 7545 2993 7584
rect 2929 7526 2993 7545
rect 3098 7565 3119 7606
rect 3155 7565 3180 7606
rect 3098 7536 3180 7565
rect 1809 7494 1867 7499
rect 1676 7482 1732 7489
rect 2301 7482 2306 7502
rect 2327 7482 2333 7502
rect 1676 7481 1711 7482
rect 2301 7475 2333 7482
rect 2724 7505 2780 7510
rect 2724 7485 2731 7505
rect 2751 7485 2780 7505
rect 2724 7478 2780 7485
rect 2724 7477 2759 7478
rect 967 7426 1078 7430
rect 2750 7426 4320 7427
rect 289 7408 4320 7426
rect 289 7388 975 7408
rect 994 7388 1052 7408
rect 1071 7404 4320 7408
rect 1071 7388 2023 7404
rect 289 7384 2023 7388
rect 2042 7384 2100 7404
rect 2119 7384 4320 7404
rect 289 7370 4320 7384
rect 289 6747 396 7370
rect 2015 7367 2126 7370
rect 775 7321 839 7325
rect 771 7315 839 7321
rect 771 7282 788 7315
rect 828 7282 839 7315
rect 771 7270 839 7282
rect 1822 7284 1887 7306
rect 771 7268 828 7270
rect 775 6907 826 7268
rect 1822 7245 1839 7284
rect 1884 7245 1887 7284
rect 1463 7200 1498 7202
rect 1463 7191 1567 7200
rect 1463 7190 1514 7191
rect 1463 7170 1466 7190
rect 1491 7171 1514 7190
rect 1546 7171 1567 7191
rect 1491 7170 1567 7171
rect 1463 7163 1567 7170
rect 1463 7151 1498 7163
rect 875 7085 1078 7098
rect 875 7052 899 7085
rect 935 7084 1078 7085
rect 935 7081 1046 7084
rect 935 7054 972 7081
rect 1001 7057 1046 7081
rect 1075 7057 1078 7084
rect 1001 7054 1078 7057
rect 935 7052 1078 7054
rect 875 7039 1078 7052
rect 875 7038 976 7039
rect 1253 6976 1285 6983
rect 1253 6956 1260 6976
rect 1281 6956 1285 6976
rect 764 6898 829 6907
rect 764 6861 774 6898
rect 814 6864 829 6898
rect 1253 6891 1285 6956
rect 1465 6947 1496 7151
rect 1700 7146 1732 7147
rect 1697 7141 1732 7146
rect 1697 7121 1704 7141
rect 1724 7121 1732 7141
rect 1697 7113 1732 7121
rect 1465 6917 1471 6947
rect 1492 6917 1496 6947
rect 1465 6909 1496 6917
rect 1623 6891 1663 6892
rect 1253 6889 1665 6891
rect 814 6861 831 6864
rect 764 6842 831 6861
rect 764 6821 778 6842
rect 814 6821 831 6842
rect 764 6814 831 6821
rect 1253 6863 1633 6889
rect 1659 6863 1665 6889
rect 1253 6855 1665 6863
rect 1253 6827 1285 6855
rect 1698 6835 1732 7113
rect 1822 6945 1887 7245
rect 3093 7269 3186 7284
rect 3093 7225 3108 7269
rect 3168 7225 3186 7269
rect 1253 6807 1258 6827
rect 1279 6807 1285 6827
rect 1253 6800 1285 6807
rect 1676 6830 1732 6835
rect 1676 6810 1683 6830
rect 1703 6810 1732 6830
rect 1676 6803 1732 6810
rect 1812 6934 1892 6945
rect 1812 6908 1829 6934
rect 1869 6908 1892 6934
rect 1812 6881 1892 6908
rect 1812 6855 1833 6881
rect 1873 6855 1892 6881
rect 1812 6836 1892 6855
rect 1812 6810 1836 6836
rect 1876 6810 1892 6836
rect 1676 6802 1711 6803
rect 1812 6798 1892 6810
rect 3093 6852 3186 7225
rect 3370 7080 3573 7093
rect 3370 7047 3394 7080
rect 3430 7079 3573 7080
rect 3430 7076 3541 7079
rect 3430 7049 3467 7076
rect 3496 7052 3541 7076
rect 3570 7052 3573 7079
rect 3496 7049 3573 7052
rect 3430 7047 3573 7049
rect 3370 7034 3573 7047
rect 3370 7033 3471 7034
rect 3093 6811 3108 6852
rect 3162 6811 3186 6852
rect 3093 6804 3186 6811
rect 3748 6971 3780 6978
rect 3748 6951 3755 6971
rect 3776 6951 3780 6971
rect 3748 6886 3780 6951
rect 3960 6942 3991 7143
rect 4195 7141 4227 7142
rect 4192 7136 4227 7141
rect 4192 7116 4199 7136
rect 4219 7116 4227 7136
rect 4192 7108 4227 7116
rect 3960 6912 3966 6942
rect 3987 6912 3991 6942
rect 3960 6904 3991 6912
rect 4118 6886 4158 6887
rect 3748 6884 4160 6886
rect 3748 6858 4128 6884
rect 4154 6858 4160 6884
rect 3748 6850 4160 6858
rect 3748 6822 3780 6850
rect 4193 6830 4227 7108
rect 3748 6802 3753 6822
rect 3774 6802 3780 6822
rect 3748 6795 3780 6802
rect 4171 6825 4227 6830
rect 4171 6805 4178 6825
rect 4198 6805 4227 6825
rect 4171 6798 4227 6805
rect 4171 6797 4206 6798
rect 967 6747 1078 6751
rect 2709 6747 4353 6750
rect 287 6729 4353 6747
rect 287 6709 975 6729
rect 994 6709 1052 6729
rect 1071 6724 4353 6729
rect 1071 6709 3470 6724
rect 287 6704 3470 6709
rect 3489 6704 3547 6724
rect 3566 6704 4353 6724
rect 287 6694 4353 6704
rect 287 6691 912 6694
rect 1099 6691 4353 6694
rect 289 6463 396 6691
rect 2709 6690 4353 6691
rect 3462 6687 3573 6690
rect 757 6652 878 6662
rect 757 6650 826 6652
rect 757 6609 770 6650
rect 807 6611 826 6650
rect 863 6611 878 6652
rect 807 6609 878 6611
rect 757 6591 878 6609
rect 3962 6632 4048 6636
rect 3962 6614 3977 6632
rect 4029 6614 4048 6632
rect 3962 6605 4048 6614
rect 763 6489 842 6591
rect 1815 6551 1882 6570
rect 1815 6531 1835 6551
rect 289 6408 397 6463
rect 764 6408 842 6489
rect 1814 6485 1835 6531
rect 1865 6531 1882 6551
rect 1865 6501 1884 6531
rect 1865 6485 1885 6501
rect 1814 6469 1885 6485
rect 1464 6458 1536 6459
rect 1463 6450 1562 6458
rect 1463 6447 1515 6450
rect 1463 6412 1471 6447
rect 1496 6412 1515 6447
rect 1540 6412 1562 6450
rect 289 5979 396 6408
rect 768 6167 840 6408
rect 1463 6400 1562 6412
rect 1464 6381 1532 6400
rect 1465 6378 1498 6381
rect 1700 6378 1732 6379
rect 875 6317 1078 6330
rect 875 6284 899 6317
rect 935 6316 1078 6317
rect 935 6313 1046 6316
rect 935 6286 972 6313
rect 1001 6289 1046 6313
rect 1075 6289 1078 6316
rect 1001 6286 1078 6289
rect 935 6284 1078 6286
rect 875 6271 1078 6284
rect 875 6270 976 6271
rect 768 6125 777 6167
rect 826 6125 840 6167
rect 768 6104 840 6125
rect 768 6062 778 6104
rect 827 6062 840 6104
rect 768 6044 840 6062
rect 1253 6208 1285 6215
rect 1253 6188 1260 6208
rect 1281 6188 1285 6208
rect 1253 6123 1285 6188
rect 1465 6179 1496 6378
rect 1697 6373 1732 6378
rect 1697 6353 1704 6373
rect 1724 6353 1732 6373
rect 1697 6345 1732 6353
rect 1465 6149 1471 6179
rect 1492 6149 1496 6179
rect 1465 6141 1496 6149
rect 1623 6123 1663 6124
rect 1253 6121 1665 6123
rect 1253 6095 1633 6121
rect 1659 6095 1665 6121
rect 1253 6087 1665 6095
rect 1253 6059 1285 6087
rect 1698 6067 1732 6345
rect 1814 6158 1884 6469
rect 3739 6459 3811 6460
rect 3738 6456 3827 6459
rect 2510 6454 3827 6456
rect 2507 6451 3827 6454
rect 2507 6448 3790 6451
rect 2507 6413 3746 6448
rect 3771 6413 3790 6448
rect 3815 6413 3827 6451
rect 2507 6403 3827 6413
rect 4003 6452 4039 6605
rect 4003 6429 4009 6452
rect 4033 6429 4039 6452
rect 4003 6408 4039 6429
rect 2507 6401 3792 6403
rect 2507 6391 2604 6401
rect 2513 6382 2549 6391
rect 4003 6385 4009 6408
rect 4033 6385 4039 6408
rect 1923 6313 2126 6326
rect 1923 6280 1947 6313
rect 1983 6312 2126 6313
rect 1983 6309 2094 6312
rect 1983 6282 2020 6309
rect 2049 6285 2094 6309
rect 2123 6285 2126 6312
rect 2049 6282 2126 6285
rect 1983 6280 2126 6282
rect 1923 6267 2126 6280
rect 1923 6266 2024 6267
rect 1253 6039 1258 6059
rect 1279 6039 1285 6059
rect 1253 6032 1285 6039
rect 1676 6062 1732 6067
rect 1676 6042 1683 6062
rect 1703 6042 1732 6062
rect 1809 6152 1884 6158
rect 1809 6119 1817 6152
rect 1870 6119 1884 6152
rect 1809 6094 1884 6119
rect 1809 6061 1822 6094
rect 1875 6061 1884 6094
rect 1809 6052 1884 6061
rect 2301 6204 2333 6211
rect 2301 6184 2308 6204
rect 2329 6184 2333 6204
rect 2301 6119 2333 6184
rect 2513 6175 2544 6382
rect 2748 6374 2780 6375
rect 4003 6374 4039 6385
rect 2745 6369 2780 6374
rect 2745 6349 2752 6369
rect 2772 6349 2780 6369
rect 2745 6341 2780 6349
rect 2513 6145 2519 6175
rect 2540 6145 2544 6175
rect 2513 6137 2544 6145
rect 2671 6119 2711 6120
rect 2301 6117 2713 6119
rect 2301 6091 2681 6117
rect 2707 6091 2713 6117
rect 2301 6083 2713 6091
rect 2301 6055 2333 6083
rect 2746 6063 2780 6341
rect 1809 6047 1867 6052
rect 1676 6035 1732 6042
rect 2301 6035 2306 6055
rect 2327 6035 2333 6055
rect 1676 6034 1711 6035
rect 2301 6028 2333 6035
rect 2724 6058 2780 6063
rect 2724 6038 2731 6058
rect 2751 6038 2780 6058
rect 2724 6031 2780 6038
rect 2724 6030 2759 6031
rect 967 5979 1078 5983
rect 2842 5979 4001 5980
rect 289 5961 4001 5979
rect 289 5941 975 5961
rect 994 5941 1052 5961
rect 1071 5957 4001 5961
rect 1071 5941 2023 5957
rect 289 5937 2023 5941
rect 2042 5937 2100 5957
rect 2119 5937 4001 5957
rect 289 5923 4001 5937
rect 289 5300 396 5923
rect 2015 5920 2126 5923
rect 775 5874 839 5878
rect 771 5868 839 5874
rect 771 5835 788 5868
rect 828 5835 839 5868
rect 771 5823 839 5835
rect 1822 5837 1887 5859
rect 771 5821 828 5823
rect 775 5460 826 5821
rect 1822 5798 1839 5837
rect 1884 5798 1887 5837
rect 4908 5835 4960 8141
rect 5069 8118 5104 8184
rect 5069 6802 5103 8118
rect 5407 7971 5512 13106
rect 8707 13072 8818 13075
rect 10437 13072 10544 13687
rect 6471 13058 10544 13072
rect 6471 13038 8714 13058
rect 8733 13038 8791 13058
rect 8810 13054 10544 13058
rect 8810 13038 9762 13054
rect 6471 13034 9762 13038
rect 9781 13034 9839 13054
rect 9858 13034 10544 13054
rect 6471 13016 10544 13034
rect 6471 13015 7991 13016
rect 9755 13012 9866 13016
rect 8074 12964 8109 12965
rect 8053 12957 8109 12964
rect 8053 12937 8082 12957
rect 8102 12937 8109 12957
rect 8053 12932 8109 12937
rect 8500 12960 8532 12967
rect 9122 12960 9157 12961
rect 8500 12940 8506 12960
rect 8527 12940 8532 12960
rect 9101 12953 9157 12960
rect 8966 12943 9024 12948
rect 8053 12654 8087 12932
rect 8500 12912 8532 12940
rect 8120 12904 8532 12912
rect 8120 12878 8126 12904
rect 8152 12878 8532 12904
rect 8120 12876 8532 12878
rect 8122 12875 8162 12876
rect 8289 12850 8320 12858
rect 8289 12820 8293 12850
rect 8314 12820 8320 12850
rect 8053 12646 8088 12654
rect 8053 12626 8061 12646
rect 8081 12626 8088 12646
rect 8053 12621 8088 12626
rect 8053 12620 8085 12621
rect 8289 12620 8320 12820
rect 8500 12811 8532 12876
rect 8500 12791 8504 12811
rect 8525 12791 8532 12811
rect 8500 12784 8532 12791
rect 8949 12934 9024 12943
rect 8949 12901 8958 12934
rect 9011 12901 9024 12934
rect 8949 12876 9024 12901
rect 8949 12843 8963 12876
rect 9016 12843 9024 12876
rect 8949 12837 9024 12843
rect 9101 12933 9130 12953
rect 9150 12933 9157 12953
rect 9101 12928 9157 12933
rect 9548 12956 9580 12963
rect 9548 12936 9554 12956
rect 9575 12936 9580 12956
rect 8809 12728 8910 12729
rect 8707 12715 8910 12728
rect 8707 12713 8850 12715
rect 8707 12710 8784 12713
rect 8707 12683 8710 12710
rect 8739 12686 8784 12710
rect 8813 12686 8850 12713
rect 8739 12683 8850 12686
rect 8707 12682 8850 12683
rect 8886 12682 8910 12715
rect 8707 12669 8910 12682
rect 8286 12613 8325 12620
rect 8284 12596 8325 12613
rect 8286 12571 8325 12596
rect 6980 12563 8325 12571
rect 6980 12535 6995 12563
rect 7023 12537 8325 12563
rect 7023 12535 8322 12537
rect 6980 12530 8322 12535
rect 8949 12526 9019 12837
rect 9101 12650 9135 12928
rect 9548 12908 9580 12936
rect 9168 12900 9580 12908
rect 9168 12874 9174 12900
rect 9200 12874 9580 12900
rect 9168 12872 9580 12874
rect 9170 12871 9210 12872
rect 9337 12846 9368 12854
rect 9337 12816 9341 12846
rect 9362 12816 9368 12846
rect 9101 12642 9136 12650
rect 9101 12622 9109 12642
rect 9129 12622 9136 12642
rect 9101 12617 9136 12622
rect 9337 12617 9368 12816
rect 9548 12807 9580 12872
rect 9548 12787 9552 12807
rect 9573 12787 9580 12807
rect 9548 12780 9580 12787
rect 9993 12933 10065 12951
rect 9993 12891 10006 12933
rect 10055 12891 10065 12933
rect 9993 12870 10065 12891
rect 9993 12828 10007 12870
rect 10056 12828 10065 12870
rect 9857 12724 9958 12725
rect 9755 12711 9958 12724
rect 9755 12709 9898 12711
rect 9755 12706 9832 12709
rect 9755 12679 9758 12706
rect 9787 12682 9832 12706
rect 9861 12682 9898 12709
rect 9787 12679 9898 12682
rect 9755 12678 9898 12679
rect 9934 12678 9958 12711
rect 9755 12665 9958 12678
rect 9101 12616 9133 12617
rect 9335 12614 9368 12617
rect 9301 12595 9369 12614
rect 9271 12583 9370 12595
rect 9993 12587 10065 12828
rect 10437 12587 10544 13016
rect 10999 13428 11106 13687
rect 11478 13616 11550 13917
rect 12174 13907 12246 13908
rect 12173 13899 12272 13907
rect 12173 13896 12225 13899
rect 12173 13861 12181 13896
rect 12206 13861 12225 13896
rect 12250 13861 12272 13899
rect 12173 13849 12272 13861
rect 12174 13830 12242 13849
rect 12175 13827 12208 13830
rect 12410 13827 12442 13828
rect 11585 13766 11788 13779
rect 11585 13733 11609 13766
rect 11645 13765 11788 13766
rect 11645 13762 11756 13765
rect 11645 13735 11682 13762
rect 11711 13738 11756 13762
rect 11785 13738 11788 13765
rect 11711 13735 11788 13738
rect 11645 13733 11788 13735
rect 11585 13720 11788 13733
rect 11585 13719 11686 13720
rect 11478 13574 11487 13616
rect 11536 13574 11550 13616
rect 11478 13553 11550 13574
rect 11478 13511 11488 13553
rect 11537 13511 11550 13553
rect 11478 13493 11550 13511
rect 11963 13657 11995 13664
rect 11963 13637 11970 13657
rect 11991 13637 11995 13657
rect 11963 13572 11995 13637
rect 12175 13628 12206 13827
rect 12407 13822 12442 13827
rect 12407 13802 12414 13822
rect 12434 13802 12442 13822
rect 12407 13794 12442 13802
rect 12175 13598 12181 13628
rect 12202 13598 12206 13628
rect 12175 13590 12206 13598
rect 12333 13572 12373 13573
rect 11963 13570 12375 13572
rect 11963 13544 12343 13570
rect 12369 13544 12375 13570
rect 11963 13536 12375 13544
rect 11963 13508 11995 13536
rect 12408 13516 12442 13794
rect 12524 13607 12594 13907
rect 13223 13900 13312 13907
rect 13223 13897 13275 13900
rect 13223 13862 13231 13897
rect 13256 13862 13275 13897
rect 13300 13862 13312 13900
rect 13223 13850 13312 13862
rect 13223 13849 13292 13850
rect 13223 13831 13259 13849
rect 12633 13762 12836 13775
rect 12633 13729 12657 13762
rect 12693 13761 12836 13762
rect 12693 13758 12804 13761
rect 12693 13731 12730 13758
rect 12759 13734 12804 13758
rect 12833 13734 12836 13761
rect 12759 13731 12836 13734
rect 12693 13729 12836 13731
rect 12633 13716 12836 13729
rect 12633 13715 12734 13716
rect 11963 13488 11968 13508
rect 11989 13488 11995 13508
rect 11963 13481 11995 13488
rect 12386 13511 12442 13516
rect 12386 13491 12393 13511
rect 12413 13491 12442 13511
rect 12519 13601 12594 13607
rect 12519 13568 12527 13601
rect 12580 13568 12594 13601
rect 12519 13543 12594 13568
rect 12519 13510 12532 13543
rect 12585 13510 12594 13543
rect 12519 13501 12594 13510
rect 13011 13653 13043 13660
rect 13011 13633 13018 13653
rect 13039 13633 13043 13653
rect 13011 13568 13043 13633
rect 13223 13624 13254 13831
rect 13458 13823 13490 13824
rect 13455 13818 13490 13823
rect 13455 13798 13462 13818
rect 13482 13798 13490 13818
rect 13455 13790 13490 13798
rect 13223 13594 13229 13624
rect 13250 13594 13254 13624
rect 13223 13586 13254 13594
rect 13381 13568 13421 13569
rect 13011 13566 13423 13568
rect 13011 13540 13391 13566
rect 13417 13540 13423 13566
rect 13011 13532 13423 13540
rect 13011 13504 13043 13532
rect 13456 13512 13490 13790
rect 13639 13605 13701 13907
rect 13808 13608 13890 13964
rect 15075 13804 15124 14091
rect 15075 13772 15244 13804
rect 15075 13766 15190 13772
rect 15075 13757 15130 13766
rect 15065 13669 15130 13757
rect 15168 13675 15190 13766
rect 15228 13675 15244 13772
rect 15168 13669 15244 13675
rect 15065 13658 15244 13669
rect 13639 13586 13703 13605
rect 13639 13547 13652 13586
rect 13686 13547 13703 13586
rect 13639 13528 13703 13547
rect 13808 13567 13829 13608
rect 13865 13567 13890 13608
rect 13808 13538 13890 13567
rect 15075 13653 15244 13658
rect 12519 13496 12577 13501
rect 12386 13484 12442 13491
rect 13011 13484 13016 13504
rect 13037 13484 13043 13504
rect 12386 13483 12421 13484
rect 13011 13477 13043 13484
rect 13434 13507 13490 13512
rect 13434 13487 13441 13507
rect 13461 13487 13490 13507
rect 13434 13480 13490 13487
rect 13434 13479 13469 13480
rect 11677 13428 11788 13432
rect 13460 13428 14573 13429
rect 10999 13410 14573 13428
rect 10999 13390 11685 13410
rect 11704 13390 11762 13410
rect 11781 13406 14573 13410
rect 11781 13390 12733 13406
rect 10999 13386 12733 13390
rect 12752 13386 12810 13406
rect 12829 13386 14573 13406
rect 10999 13372 14573 13386
rect 10999 12749 11106 13372
rect 12725 13369 12836 13372
rect 11485 13323 11549 13327
rect 11481 13317 11549 13323
rect 11481 13284 11498 13317
rect 11538 13284 11549 13317
rect 11481 13272 11549 13284
rect 12532 13286 12597 13308
rect 11481 13270 11538 13272
rect 11485 12909 11536 13270
rect 12532 13247 12549 13286
rect 12594 13247 12597 13286
rect 12173 13202 12208 13204
rect 12173 13193 12277 13202
rect 12173 13192 12224 13193
rect 12173 13172 12176 13192
rect 12201 13173 12224 13192
rect 12256 13173 12277 13193
rect 12201 13172 12277 13173
rect 12173 13165 12277 13172
rect 12173 13153 12208 13165
rect 11585 13087 11788 13100
rect 11585 13054 11609 13087
rect 11645 13086 11788 13087
rect 11645 13083 11756 13086
rect 11645 13056 11682 13083
rect 11711 13059 11756 13083
rect 11785 13059 11788 13086
rect 11711 13056 11788 13059
rect 11645 13054 11788 13056
rect 11585 13041 11788 13054
rect 11585 13040 11686 13041
rect 11963 12978 11995 12985
rect 11963 12958 11970 12978
rect 11991 12958 11995 12978
rect 11474 12900 11539 12909
rect 11474 12863 11484 12900
rect 11524 12866 11539 12900
rect 11963 12893 11995 12958
rect 12175 12949 12206 13153
rect 12410 13148 12442 13149
rect 12407 13143 12442 13148
rect 12407 13123 12414 13143
rect 12434 13123 12442 13143
rect 12407 13115 12442 13123
rect 12175 12919 12181 12949
rect 12202 12919 12206 12949
rect 12175 12911 12206 12919
rect 12333 12893 12373 12894
rect 11963 12891 12375 12893
rect 11524 12863 11541 12866
rect 11474 12844 11541 12863
rect 11474 12823 11488 12844
rect 11524 12823 11541 12844
rect 11474 12816 11541 12823
rect 11963 12865 12343 12891
rect 12369 12865 12375 12891
rect 11963 12857 12375 12865
rect 11963 12829 11995 12857
rect 12408 12837 12442 13115
rect 12532 12947 12597 13247
rect 13803 13271 13896 13286
rect 13803 13227 13818 13271
rect 13878 13227 13896 13271
rect 11963 12809 11968 12829
rect 11989 12809 11995 12829
rect 11963 12802 11995 12809
rect 12386 12832 12442 12837
rect 12386 12812 12393 12832
rect 12413 12812 12442 12832
rect 12386 12805 12442 12812
rect 12522 12936 12602 12947
rect 12522 12910 12539 12936
rect 12579 12910 12602 12936
rect 12522 12883 12602 12910
rect 12522 12857 12543 12883
rect 12583 12857 12602 12883
rect 12522 12838 12602 12857
rect 12522 12812 12546 12838
rect 12586 12812 12602 12838
rect 12386 12804 12421 12805
rect 12522 12800 12602 12812
rect 13803 12854 13896 13227
rect 14080 13082 14283 13095
rect 14080 13049 14104 13082
rect 14140 13081 14283 13082
rect 14140 13078 14251 13081
rect 14140 13051 14177 13078
rect 14206 13054 14251 13078
rect 14280 13054 14283 13081
rect 14206 13051 14283 13054
rect 14140 13049 14283 13051
rect 14080 13036 14283 13049
rect 14080 13035 14181 13036
rect 13803 12813 13818 12854
rect 13872 12813 13896 12854
rect 13803 12806 13896 12813
rect 14458 12973 14490 12980
rect 14458 12953 14465 12973
rect 14486 12953 14490 12973
rect 14458 12888 14490 12953
rect 14670 12944 14701 13145
rect 14905 13143 14937 13144
rect 14902 13138 14937 13143
rect 14902 13118 14909 13138
rect 14929 13118 14937 13138
rect 14902 13110 14937 13118
rect 14670 12914 14676 12944
rect 14697 12914 14701 12944
rect 14670 12906 14701 12914
rect 14828 12888 14868 12889
rect 14458 12886 14870 12888
rect 14458 12860 14838 12886
rect 14864 12860 14870 12886
rect 14458 12852 14870 12860
rect 14458 12824 14490 12852
rect 14903 12832 14937 13110
rect 14458 12804 14463 12824
rect 14484 12804 14490 12824
rect 14458 12797 14490 12804
rect 14881 12827 14937 12832
rect 14881 12807 14888 12827
rect 14908 12807 14937 12827
rect 14881 12800 14937 12807
rect 14881 12799 14916 12800
rect 11677 12749 11788 12753
rect 13419 12749 14968 12752
rect 10997 12731 14968 12749
rect 10997 12711 11685 12731
rect 11704 12711 11762 12731
rect 11781 12726 14968 12731
rect 11781 12711 14180 12726
rect 10997 12706 14180 12711
rect 14199 12706 14257 12726
rect 14276 12706 14968 12726
rect 10997 12696 14968 12706
rect 10997 12693 11622 12696
rect 11809 12693 14968 12696
rect 9271 12545 9293 12583
rect 9318 12548 9337 12583
rect 9362 12548 9370 12583
rect 9318 12545 9370 12548
rect 9271 12537 9370 12545
rect 9297 12536 9369 12537
rect 8948 12510 9019 12526
rect 8948 12494 8968 12510
rect 8949 12464 8968 12494
rect 8951 12444 8968 12464
rect 8998 12464 9019 12510
rect 9991 12506 10069 12587
rect 10436 12532 10544 12587
rect 8998 12444 9018 12464
rect 8951 12425 9018 12444
rect 9991 12404 10070 12506
rect 9955 12386 10076 12404
rect 9955 12384 10026 12386
rect 9955 12343 9970 12384
rect 10007 12345 10026 12384
rect 10063 12345 10076 12386
rect 10007 12343 10076 12345
rect 9955 12333 10076 12343
rect 7260 12305 7371 12308
rect 6471 12304 8124 12305
rect 10437 12304 10544 12532
rect 10999 12465 11106 12693
rect 13419 12692 14968 12693
rect 14172 12689 14283 12692
rect 11467 12654 11588 12664
rect 11467 12652 11536 12654
rect 11467 12611 11480 12652
rect 11517 12613 11536 12652
rect 11573 12613 11588 12654
rect 11517 12611 11588 12613
rect 11467 12593 11588 12611
rect 14672 12634 14758 12638
rect 14672 12616 14687 12634
rect 14739 12616 14758 12634
rect 14672 12607 14758 12616
rect 11473 12491 11552 12593
rect 12525 12553 12592 12572
rect 12525 12533 12545 12553
rect 10999 12410 11107 12465
rect 11474 12410 11552 12491
rect 12524 12487 12545 12533
rect 12575 12533 12592 12553
rect 12575 12503 12594 12533
rect 12575 12487 12595 12503
rect 12524 12471 12595 12487
rect 12174 12460 12246 12461
rect 12173 12452 12272 12460
rect 12173 12449 12225 12452
rect 12173 12414 12181 12449
rect 12206 12414 12225 12449
rect 12250 12414 12272 12452
rect 6471 12301 9734 12304
rect 9921 12301 10546 12304
rect 6471 12291 10546 12301
rect 6471 12271 7267 12291
rect 7286 12271 7344 12291
rect 7363 12286 10546 12291
rect 7363 12271 9762 12286
rect 6471 12266 9762 12271
rect 9781 12266 9839 12286
rect 9858 12266 10546 12286
rect 6471 12248 10546 12266
rect 6471 12245 8124 12248
rect 9755 12244 9866 12248
rect 6627 12197 6662 12198
rect 6606 12190 6662 12197
rect 6606 12170 6635 12190
rect 6655 12170 6662 12190
rect 6606 12165 6662 12170
rect 7053 12193 7085 12200
rect 7053 12173 7059 12193
rect 7080 12173 7085 12193
rect 6606 11887 6640 12165
rect 7053 12145 7085 12173
rect 8941 12185 9021 12197
rect 9122 12192 9157 12193
rect 6673 12137 7085 12145
rect 6673 12111 6679 12137
rect 6705 12111 7085 12137
rect 7471 12151 7908 12164
rect 7471 12128 7484 12151
rect 7510 12144 7908 12151
rect 7510 12128 7864 12144
rect 7471 12121 7864 12128
rect 7890 12121 7908 12144
rect 7471 12115 7908 12121
rect 8941 12159 8957 12185
rect 8997 12159 9021 12185
rect 8941 12140 9021 12159
rect 6673 12109 7085 12111
rect 6675 12108 6715 12109
rect 6842 12083 6873 12091
rect 6842 12053 6846 12083
rect 6867 12053 6873 12083
rect 6606 11879 6641 11887
rect 6606 11859 6614 11879
rect 6634 11859 6641 11879
rect 6606 11854 6641 11859
rect 6606 11853 6638 11854
rect 6842 11846 6873 12053
rect 7053 12044 7085 12109
rect 8941 12114 8960 12140
rect 9000 12114 9021 12140
rect 8941 12087 9021 12114
rect 8941 12061 8964 12087
rect 9004 12061 9021 12087
rect 8941 12050 9021 12061
rect 9101 12185 9157 12192
rect 9101 12165 9130 12185
rect 9150 12165 9157 12185
rect 9101 12160 9157 12165
rect 9548 12188 9580 12195
rect 9548 12168 9554 12188
rect 9575 12168 9580 12188
rect 7053 12024 7057 12044
rect 7078 12024 7085 12044
rect 7053 12017 7085 12024
rect 7362 11961 7463 11962
rect 7260 11948 7463 11961
rect 7260 11946 7403 11948
rect 7260 11943 7337 11946
rect 7260 11916 7263 11943
rect 7292 11919 7337 11943
rect 7366 11919 7403 11946
rect 7292 11916 7403 11919
rect 7260 11915 7403 11916
rect 7439 11915 7463 11948
rect 7260 11902 7463 11915
rect 6840 11840 6873 11846
rect 6836 11836 6873 11840
rect 6836 11826 6874 11836
rect 6836 11813 6846 11826
rect 6837 11789 6846 11813
rect 6863 11789 6874 11826
rect 6837 11768 6874 11789
rect 8946 11750 9011 12050
rect 9101 11882 9135 12160
rect 9548 12140 9580 12168
rect 9168 12132 9580 12140
rect 9168 12106 9174 12132
rect 9200 12106 9580 12132
rect 10002 12174 10069 12181
rect 10002 12153 10019 12174
rect 10055 12153 10069 12174
rect 10002 12134 10069 12153
rect 10002 12131 10019 12134
rect 9168 12104 9580 12106
rect 9170 12103 9210 12104
rect 9337 12078 9368 12086
rect 9337 12048 9341 12078
rect 9362 12048 9368 12078
rect 9101 11874 9136 11882
rect 9101 11854 9109 11874
rect 9129 11854 9136 11874
rect 9101 11849 9136 11854
rect 9101 11848 9133 11849
rect 9337 11844 9368 12048
rect 9548 12039 9580 12104
rect 10004 12097 10019 12131
rect 10059 12097 10069 12134
rect 10004 12088 10069 12097
rect 9548 12019 9552 12039
rect 9573 12019 9580 12039
rect 9548 12012 9580 12019
rect 9857 11956 9958 11957
rect 9755 11943 9958 11956
rect 9755 11941 9898 11943
rect 9755 11938 9832 11941
rect 9755 11911 9758 11938
rect 9787 11914 9832 11938
rect 9861 11914 9898 11941
rect 9787 11911 9898 11914
rect 9755 11910 9898 11911
rect 9934 11910 9958 11943
rect 9755 11897 9958 11910
rect 9335 11832 9370 11844
rect 9266 11825 9370 11832
rect 9266 11824 9342 11825
rect 9266 11804 9287 11824
rect 9319 11805 9342 11824
rect 9367 11805 9370 11825
rect 9319 11804 9370 11805
rect 9266 11795 9370 11804
rect 9335 11793 9370 11795
rect 8946 11711 8949 11750
rect 8994 11711 9011 11750
rect 10007 11727 10058 12088
rect 10005 11725 10062 11727
rect 8946 11689 9011 11711
rect 9994 11713 10062 11725
rect 9994 11680 10005 11713
rect 10045 11680 10062 11713
rect 9994 11674 10062 11680
rect 9994 11670 10058 11674
rect 8707 11625 8818 11628
rect 10437 11625 10544 12248
rect 6094 11611 10544 11625
rect 6094 11591 8714 11611
rect 8733 11591 8791 11611
rect 8810 11607 10544 11611
rect 8810 11591 9762 11607
rect 6094 11587 9762 11591
rect 9781 11587 9839 11607
rect 9858 11587 10544 11607
rect 6094 11573 10544 11587
rect 6513 11569 10544 11573
rect 6513 11568 8083 11569
rect 9755 11565 9866 11569
rect 8074 11517 8109 11518
rect 8053 11510 8109 11517
rect 8053 11490 8082 11510
rect 8102 11490 8109 11510
rect 8053 11485 8109 11490
rect 8500 11513 8532 11520
rect 9122 11513 9157 11514
rect 8500 11493 8506 11513
rect 8527 11493 8532 11513
rect 9101 11506 9157 11513
rect 8966 11496 9024 11501
rect 8053 11207 8087 11485
rect 8500 11465 8532 11493
rect 8120 11457 8532 11465
rect 8120 11431 8126 11457
rect 8152 11431 8532 11457
rect 8120 11429 8532 11431
rect 8122 11428 8162 11429
rect 8289 11403 8320 11411
rect 8289 11373 8293 11403
rect 8314 11373 8320 11403
rect 8053 11199 8088 11207
rect 8053 11179 8061 11199
rect 8081 11179 8088 11199
rect 8053 11174 8088 11179
rect 8053 11173 8085 11174
rect 8289 11166 8320 11373
rect 8500 11364 8532 11429
rect 8500 11344 8504 11364
rect 8525 11344 8532 11364
rect 8500 11337 8532 11344
rect 8949 11487 9024 11496
rect 8949 11454 8958 11487
rect 9011 11454 9024 11487
rect 8949 11429 9024 11454
rect 8949 11396 8963 11429
rect 9016 11396 9024 11429
rect 8949 11390 9024 11396
rect 9101 11486 9130 11506
rect 9150 11486 9157 11506
rect 9101 11481 9157 11486
rect 9548 11509 9580 11516
rect 9548 11489 9554 11509
rect 9575 11489 9580 11509
rect 8809 11281 8910 11282
rect 8707 11268 8910 11281
rect 8707 11266 8850 11268
rect 8707 11263 8784 11266
rect 8707 11236 8710 11263
rect 8739 11239 8784 11263
rect 8813 11239 8850 11266
rect 8739 11236 8850 11239
rect 8707 11235 8850 11236
rect 8886 11235 8910 11268
rect 8707 11222 8910 11235
rect 7787 11153 7951 11156
rect 8284 11153 8320 11166
rect 6986 11135 8325 11153
rect 6986 11097 6996 11135
rect 7021 11120 8325 11135
rect 7021 11097 7031 11120
rect 7787 11113 7951 11120
rect 6986 11089 7031 11097
rect 7000 11088 7031 11089
rect 8949 11074 9019 11390
rect 9101 11203 9135 11481
rect 9548 11461 9580 11489
rect 9168 11453 9580 11461
rect 9168 11427 9174 11453
rect 9200 11427 9580 11453
rect 9168 11425 9580 11427
rect 9170 11424 9210 11425
rect 9337 11399 9368 11407
rect 9337 11369 9341 11399
rect 9362 11369 9368 11399
rect 9101 11195 9136 11203
rect 9101 11175 9109 11195
rect 9129 11175 9136 11195
rect 9101 11170 9136 11175
rect 9337 11170 9368 11369
rect 9548 11360 9580 11425
rect 9548 11340 9552 11360
rect 9573 11340 9580 11360
rect 9548 11333 9580 11340
rect 9993 11486 10065 11504
rect 9993 11444 10006 11486
rect 10055 11444 10065 11486
rect 9993 11423 10065 11444
rect 9993 11381 10007 11423
rect 10056 11381 10065 11423
rect 9857 11277 9958 11278
rect 9755 11264 9958 11277
rect 9755 11262 9898 11264
rect 9755 11259 9832 11262
rect 9755 11232 9758 11259
rect 9787 11235 9832 11259
rect 9861 11235 9898 11262
rect 9787 11232 9898 11235
rect 9755 11231 9898 11232
rect 9934 11231 9958 11264
rect 9755 11218 9958 11231
rect 9101 11169 9133 11170
rect 9335 11167 9368 11170
rect 9301 11148 9369 11167
rect 9271 11136 9370 11148
rect 9271 11098 9293 11136
rect 9318 11101 9337 11136
rect 9362 11101 9370 11136
rect 9318 11098 9370 11101
rect 9271 11090 9370 11098
rect 9297 11089 9369 11090
rect 8949 11055 9028 11074
rect 8952 11035 9028 11055
rect 8945 11011 9028 11035
rect 9993 11070 10065 11381
rect 9993 11027 10069 11070
rect 8945 10945 8957 11011
rect 9011 10945 9028 11011
rect 8945 10925 9028 10945
rect 8945 10888 8962 10925
rect 9006 10911 9028 10925
rect 9994 10976 10069 11027
rect 10437 10976 10544 11569
rect 10999 11981 11106 12410
rect 11478 12169 11550 12410
rect 12173 12402 12272 12414
rect 12174 12383 12242 12402
rect 12175 12380 12208 12383
rect 12410 12380 12442 12381
rect 11585 12319 11788 12332
rect 11585 12286 11609 12319
rect 11645 12318 11788 12319
rect 11645 12315 11756 12318
rect 11645 12288 11682 12315
rect 11711 12291 11756 12315
rect 11785 12291 11788 12318
rect 11711 12288 11788 12291
rect 11645 12286 11788 12288
rect 11585 12273 11788 12286
rect 11585 12272 11686 12273
rect 11478 12127 11487 12169
rect 11536 12127 11550 12169
rect 11478 12106 11550 12127
rect 11478 12064 11488 12106
rect 11537 12064 11550 12106
rect 11478 12046 11550 12064
rect 11963 12210 11995 12217
rect 11963 12190 11970 12210
rect 11991 12190 11995 12210
rect 11963 12125 11995 12190
rect 12175 12181 12206 12380
rect 12407 12375 12442 12380
rect 12407 12355 12414 12375
rect 12434 12355 12442 12375
rect 12407 12347 12442 12355
rect 12175 12151 12181 12181
rect 12202 12151 12206 12181
rect 12175 12143 12206 12151
rect 12333 12125 12373 12126
rect 11963 12123 12375 12125
rect 11963 12097 12343 12123
rect 12369 12097 12375 12123
rect 11963 12089 12375 12097
rect 11963 12061 11995 12089
rect 12408 12069 12442 12347
rect 12524 12160 12594 12471
rect 14449 12461 14521 12462
rect 14448 12458 14537 12461
rect 13220 12456 14537 12458
rect 13217 12453 14537 12456
rect 13217 12450 14500 12453
rect 13217 12415 14456 12450
rect 14481 12415 14500 12450
rect 14525 12415 14537 12453
rect 13217 12405 14537 12415
rect 14713 12454 14749 12607
rect 14713 12431 14719 12454
rect 14743 12431 14749 12454
rect 14713 12410 14749 12431
rect 13217 12403 14502 12405
rect 13217 12393 13314 12403
rect 13223 12384 13259 12393
rect 14713 12387 14719 12410
rect 14743 12387 14749 12410
rect 12633 12315 12836 12328
rect 12633 12282 12657 12315
rect 12693 12314 12836 12315
rect 12693 12311 12804 12314
rect 12693 12284 12730 12311
rect 12759 12287 12804 12311
rect 12833 12287 12836 12314
rect 12759 12284 12836 12287
rect 12693 12282 12836 12284
rect 12633 12269 12836 12282
rect 12633 12268 12734 12269
rect 11963 12041 11968 12061
rect 11989 12041 11995 12061
rect 11963 12034 11995 12041
rect 12386 12064 12442 12069
rect 12386 12044 12393 12064
rect 12413 12044 12442 12064
rect 12519 12154 12594 12160
rect 12519 12121 12527 12154
rect 12580 12121 12594 12154
rect 12519 12096 12594 12121
rect 12519 12063 12532 12096
rect 12585 12063 12594 12096
rect 12519 12054 12594 12063
rect 13011 12206 13043 12213
rect 13011 12186 13018 12206
rect 13039 12186 13043 12206
rect 13011 12121 13043 12186
rect 13223 12177 13254 12384
rect 13458 12376 13490 12377
rect 14713 12376 14749 12387
rect 13455 12371 13490 12376
rect 13455 12351 13462 12371
rect 13482 12351 13490 12371
rect 13455 12343 13490 12351
rect 13223 12147 13229 12177
rect 13250 12147 13254 12177
rect 13223 12139 13254 12147
rect 13381 12121 13421 12122
rect 13011 12119 13423 12121
rect 13011 12093 13391 12119
rect 13417 12093 13423 12119
rect 13011 12085 13423 12093
rect 13011 12057 13043 12085
rect 13456 12065 13490 12343
rect 12519 12049 12577 12054
rect 12386 12037 12442 12044
rect 13011 12037 13016 12057
rect 13037 12037 13043 12057
rect 12386 12036 12421 12037
rect 13011 12030 13043 12037
rect 13434 12060 13490 12065
rect 13434 12040 13441 12060
rect 13461 12040 13490 12060
rect 13434 12033 13490 12040
rect 13434 12032 13469 12033
rect 11677 11981 11788 11985
rect 13552 11981 14793 11982
rect 10999 11963 14793 11981
rect 10999 11943 11685 11963
rect 11704 11943 11762 11963
rect 11781 11959 14793 11963
rect 11781 11943 12733 11959
rect 10999 11939 12733 11943
rect 12752 11939 12810 11959
rect 12829 11939 14793 11959
rect 10999 11925 14793 11939
rect 10999 11302 11106 11925
rect 12725 11922 12836 11925
rect 11485 11876 11549 11880
rect 11481 11870 11549 11876
rect 11481 11837 11498 11870
rect 11538 11837 11549 11870
rect 11481 11825 11549 11837
rect 12532 11839 12597 11861
rect 11481 11823 11538 11825
rect 11485 11462 11536 11823
rect 12532 11800 12549 11839
rect 12594 11800 12597 11839
rect 12173 11755 12208 11757
rect 12173 11746 12277 11755
rect 12173 11745 12224 11746
rect 12173 11725 12176 11745
rect 12201 11726 12224 11745
rect 12256 11726 12277 11746
rect 12201 11725 12277 11726
rect 12173 11718 12277 11725
rect 12173 11706 12208 11718
rect 11585 11640 11788 11653
rect 11585 11607 11609 11640
rect 11645 11639 11788 11640
rect 11645 11636 11756 11639
rect 11645 11609 11682 11636
rect 11711 11612 11756 11636
rect 11785 11612 11788 11639
rect 11711 11609 11788 11612
rect 11645 11607 11788 11609
rect 11585 11594 11788 11607
rect 11585 11593 11686 11594
rect 11963 11531 11995 11538
rect 11963 11511 11970 11531
rect 11991 11511 11995 11531
rect 11474 11453 11539 11462
rect 11474 11416 11484 11453
rect 11524 11419 11539 11453
rect 11963 11446 11995 11511
rect 12175 11502 12206 11706
rect 12410 11701 12442 11702
rect 12407 11696 12442 11701
rect 12407 11676 12414 11696
rect 12434 11676 12442 11696
rect 12407 11668 12442 11676
rect 12175 11472 12181 11502
rect 12202 11472 12206 11502
rect 12175 11464 12206 11472
rect 12333 11446 12373 11447
rect 11963 11444 12375 11446
rect 11524 11416 11541 11419
rect 11474 11397 11541 11416
rect 11474 11376 11488 11397
rect 11524 11376 11541 11397
rect 11474 11369 11541 11376
rect 11963 11418 12343 11444
rect 12369 11418 12375 11444
rect 11963 11410 12375 11418
rect 11963 11382 11995 11410
rect 12408 11390 12442 11668
rect 12532 11500 12597 11800
rect 14711 11794 14816 11803
rect 14711 11789 14765 11794
rect 14711 11768 14724 11789
rect 14744 11773 14765 11789
rect 14785 11773 14816 11794
rect 14744 11768 14816 11773
rect 14711 11737 14816 11768
rect 14714 11720 14749 11737
rect 14713 11702 14749 11720
rect 14123 11637 14326 11650
rect 14123 11604 14147 11637
rect 14183 11636 14326 11637
rect 14183 11633 14294 11636
rect 14183 11606 14220 11633
rect 14249 11609 14294 11633
rect 14323 11609 14326 11636
rect 14249 11606 14326 11609
rect 14183 11604 14326 11606
rect 14123 11591 14326 11604
rect 14123 11590 14224 11591
rect 14501 11528 14533 11535
rect 14501 11508 14508 11528
rect 14529 11508 14533 11528
rect 11963 11362 11968 11382
rect 11989 11362 11995 11382
rect 11963 11355 11995 11362
rect 12386 11385 12442 11390
rect 12386 11365 12393 11385
rect 12413 11365 12442 11385
rect 12386 11358 12442 11365
rect 12522 11489 12602 11500
rect 12522 11463 12539 11489
rect 12579 11463 12602 11489
rect 12522 11436 12602 11463
rect 12522 11410 12543 11436
rect 12583 11410 12602 11436
rect 12522 11391 12602 11410
rect 12522 11365 12546 11391
rect 12586 11365 12602 11391
rect 12386 11357 12421 11358
rect 12522 11353 12602 11365
rect 14501 11443 14533 11508
rect 14713 11499 14744 11702
rect 14948 11698 14980 11699
rect 14945 11693 14980 11698
rect 14945 11673 14952 11693
rect 14972 11673 14980 11693
rect 14945 11665 14980 11673
rect 14713 11469 14719 11499
rect 14740 11469 14744 11499
rect 14713 11461 14744 11469
rect 14871 11443 14911 11444
rect 14501 11441 14913 11443
rect 14501 11415 14881 11441
rect 14907 11415 14913 11441
rect 14501 11407 14913 11415
rect 14501 11379 14533 11407
rect 14946 11387 14980 11665
rect 14501 11359 14506 11379
rect 14527 11359 14533 11379
rect 14501 11352 14533 11359
rect 14924 11382 14980 11387
rect 14924 11362 14931 11382
rect 14951 11362 14980 11382
rect 14924 11355 14980 11362
rect 14924 11354 14959 11355
rect 11677 11302 11788 11306
rect 13432 11302 13639 11303
rect 14215 11302 14326 11303
rect 10997 11284 15017 11302
rect 10997 11264 11685 11284
rect 11704 11264 11762 11284
rect 11781 11281 15017 11284
rect 11781 11264 14223 11281
rect 10997 11261 14223 11264
rect 14242 11261 14300 11281
rect 14319 11261 15017 11281
rect 10997 11246 15017 11261
rect 10999 11058 11106 11246
rect 13594 11244 15017 11246
rect 11467 11207 11588 11217
rect 11467 11205 11536 11207
rect 11467 11164 11480 11205
rect 11517 11166 11536 11205
rect 11573 11166 11588 11207
rect 11517 11164 11588 11166
rect 11467 11146 11588 11164
rect 10999 11054 11107 11058
rect 11473 11054 11550 11146
rect 12523 11142 12599 11158
rect 12523 11119 12538 11142
rect 9006 10888 9021 10911
rect 8945 10872 9021 10888
rect 9994 10884 10071 10976
rect 10437 10972 10545 10976
rect 9956 10866 10077 10884
rect 9956 10864 10027 10866
rect 9956 10823 9971 10864
rect 10008 10825 10027 10864
rect 10064 10825 10077 10866
rect 10008 10823 10077 10825
rect 9956 10813 10077 10823
rect 6481 10784 7950 10786
rect 10438 10784 10545 10972
rect 6481 10769 10547 10784
rect 6481 10749 7225 10769
rect 7244 10749 7302 10769
rect 7321 10766 10547 10769
rect 7321 10749 9763 10766
rect 6481 10746 9763 10749
rect 9782 10746 9840 10766
rect 9859 10746 10547 10766
rect 6481 10728 10547 10746
rect 7218 10727 7329 10728
rect 7905 10727 8112 10728
rect 9756 10724 9867 10728
rect 6585 10675 6620 10676
rect 6564 10668 6620 10675
rect 6564 10648 6593 10668
rect 6613 10648 6620 10668
rect 6564 10643 6620 10648
rect 7011 10671 7043 10678
rect 7011 10651 7017 10671
rect 7038 10651 7043 10671
rect 6564 10365 6598 10643
rect 7011 10623 7043 10651
rect 6631 10615 7043 10623
rect 6631 10589 6637 10615
rect 6663 10589 7043 10615
rect 6631 10587 7043 10589
rect 6633 10586 6673 10587
rect 6800 10561 6831 10569
rect 6800 10531 6804 10561
rect 6825 10531 6831 10561
rect 6564 10357 6599 10365
rect 6564 10337 6572 10357
rect 6592 10337 6599 10357
rect 6564 10332 6599 10337
rect 6800 10335 6831 10531
rect 7011 10522 7043 10587
rect 8942 10665 9022 10677
rect 9123 10672 9158 10673
rect 8942 10639 8958 10665
rect 8998 10639 9022 10665
rect 8942 10620 9022 10639
rect 8942 10594 8961 10620
rect 9001 10594 9022 10620
rect 8942 10567 9022 10594
rect 8942 10541 8965 10567
rect 9005 10541 9022 10567
rect 8942 10530 9022 10541
rect 9102 10665 9158 10672
rect 9102 10645 9131 10665
rect 9151 10645 9158 10665
rect 9102 10640 9158 10645
rect 9549 10668 9581 10675
rect 9549 10648 9555 10668
rect 9576 10648 9581 10668
rect 7011 10502 7015 10522
rect 7036 10502 7043 10522
rect 7011 10495 7043 10502
rect 7320 10439 7421 10440
rect 7218 10426 7421 10439
rect 7218 10424 7361 10426
rect 7218 10421 7295 10424
rect 7218 10394 7221 10421
rect 7250 10397 7295 10421
rect 7324 10397 7361 10424
rect 7250 10394 7361 10397
rect 7218 10393 7361 10394
rect 7397 10393 7421 10426
rect 7218 10380 7421 10393
rect 6564 10331 6596 10332
rect 6800 10246 6834 10335
rect 6421 10242 6834 10246
rect 5407 7917 5424 7971
rect 5487 7917 5512 7971
rect 5407 7896 5512 7917
rect 5874 10197 6834 10242
rect 8947 10230 9012 10530
rect 9102 10362 9136 10640
rect 9549 10620 9581 10648
rect 9169 10612 9581 10620
rect 9169 10586 9175 10612
rect 9201 10586 9581 10612
rect 10003 10654 10070 10661
rect 10003 10633 10020 10654
rect 10056 10633 10070 10654
rect 10003 10614 10070 10633
rect 10003 10611 10020 10614
rect 9169 10584 9581 10586
rect 9171 10583 9211 10584
rect 9338 10558 9369 10566
rect 9338 10528 9342 10558
rect 9363 10528 9369 10558
rect 9102 10354 9137 10362
rect 9102 10334 9110 10354
rect 9130 10334 9137 10354
rect 9102 10329 9137 10334
rect 9102 10328 9134 10329
rect 9338 10324 9369 10528
rect 9549 10519 9581 10584
rect 10005 10577 10020 10611
rect 10060 10577 10070 10614
rect 10005 10568 10070 10577
rect 9549 10499 9553 10519
rect 9574 10499 9581 10519
rect 9549 10492 9581 10499
rect 9858 10436 9959 10437
rect 9756 10423 9959 10436
rect 9756 10421 9899 10423
rect 9756 10418 9833 10421
rect 9756 10391 9759 10418
rect 9788 10394 9833 10418
rect 9862 10394 9899 10421
rect 9788 10391 9899 10394
rect 9756 10390 9899 10391
rect 9935 10390 9959 10423
rect 9756 10377 9959 10390
rect 9336 10312 9371 10324
rect 9267 10305 9371 10312
rect 9267 10304 9343 10305
rect 9267 10284 9288 10304
rect 9320 10285 9343 10304
rect 9368 10285 9371 10305
rect 9320 10284 9371 10285
rect 9267 10275 9371 10284
rect 9336 10273 9371 10275
rect 5874 10193 6471 10197
rect 5874 7887 5926 10193
rect 8947 10191 8950 10230
rect 8995 10191 9012 10230
rect 10008 10207 10059 10568
rect 10006 10205 10063 10207
rect 8947 10169 9012 10191
rect 9995 10193 10063 10205
rect 9995 10160 10006 10193
rect 10046 10160 10063 10193
rect 9995 10154 10063 10160
rect 9995 10150 10059 10154
rect 8708 10105 8819 10108
rect 10438 10105 10545 10728
rect 6833 10091 10545 10105
rect 6833 10071 8715 10091
rect 8734 10071 8792 10091
rect 8811 10087 10545 10091
rect 8811 10071 9763 10087
rect 6833 10067 9763 10071
rect 9782 10067 9840 10087
rect 9859 10067 10545 10087
rect 6833 10049 10545 10067
rect 6833 10048 7992 10049
rect 9756 10045 9867 10049
rect 8075 9997 8110 9998
rect 8054 9990 8110 9997
rect 8054 9970 8083 9990
rect 8103 9970 8110 9990
rect 8054 9965 8110 9970
rect 8501 9993 8533 10000
rect 9123 9993 9158 9994
rect 8501 9973 8507 9993
rect 8528 9973 8533 9993
rect 9102 9986 9158 9993
rect 8967 9976 9025 9981
rect 8054 9687 8088 9965
rect 8501 9945 8533 9973
rect 8121 9937 8533 9945
rect 8121 9911 8127 9937
rect 8153 9911 8533 9937
rect 8121 9909 8533 9911
rect 8123 9908 8163 9909
rect 8290 9883 8321 9891
rect 8290 9853 8294 9883
rect 8315 9853 8321 9883
rect 8054 9679 8089 9687
rect 8054 9659 8062 9679
rect 8082 9659 8089 9679
rect 8054 9654 8089 9659
rect 6795 9643 6831 9654
rect 8054 9653 8086 9654
rect 8290 9646 8321 9853
rect 8501 9844 8533 9909
rect 8501 9824 8505 9844
rect 8526 9824 8533 9844
rect 8501 9817 8533 9824
rect 8950 9967 9025 9976
rect 8950 9934 8959 9967
rect 9012 9934 9025 9967
rect 8950 9909 9025 9934
rect 8950 9876 8964 9909
rect 9017 9876 9025 9909
rect 8950 9870 9025 9876
rect 9102 9966 9131 9986
rect 9151 9966 9158 9986
rect 9102 9961 9158 9966
rect 9549 9989 9581 9996
rect 9549 9969 9555 9989
rect 9576 9969 9581 9989
rect 8810 9761 8911 9762
rect 8708 9748 8911 9761
rect 8708 9746 8851 9748
rect 8708 9743 8785 9746
rect 8708 9716 8711 9743
rect 8740 9719 8785 9743
rect 8814 9719 8851 9746
rect 8740 9716 8851 9719
rect 8708 9715 8851 9716
rect 8887 9715 8911 9748
rect 8708 9702 8911 9715
rect 6795 9620 6801 9643
rect 6825 9620 6831 9643
rect 8285 9637 8321 9646
rect 8230 9627 8327 9637
rect 7042 9625 8327 9627
rect 6795 9599 6831 9620
rect 6795 9576 6801 9599
rect 6825 9576 6831 9599
rect 6795 9423 6831 9576
rect 7007 9615 8327 9625
rect 7007 9577 7019 9615
rect 7044 9580 7063 9615
rect 7088 9580 8327 9615
rect 7044 9577 8327 9580
rect 7007 9574 8327 9577
rect 7007 9572 8324 9574
rect 7007 9569 7096 9572
rect 7023 9568 7095 9569
rect 8950 9559 9020 9870
rect 9102 9683 9136 9961
rect 9549 9941 9581 9969
rect 9169 9933 9581 9941
rect 9169 9907 9175 9933
rect 9201 9907 9581 9933
rect 9169 9905 9581 9907
rect 9171 9904 9211 9905
rect 9338 9879 9369 9887
rect 9338 9849 9342 9879
rect 9363 9849 9369 9879
rect 9102 9675 9137 9683
rect 9102 9655 9110 9675
rect 9130 9655 9137 9675
rect 9102 9650 9137 9655
rect 9338 9650 9369 9849
rect 9549 9840 9581 9905
rect 9549 9820 9553 9840
rect 9574 9820 9581 9840
rect 9549 9813 9581 9820
rect 9994 9966 10066 9984
rect 9994 9924 10007 9966
rect 10056 9924 10066 9966
rect 9994 9903 10066 9924
rect 9994 9861 10008 9903
rect 10057 9861 10066 9903
rect 9858 9757 9959 9758
rect 9756 9744 9959 9757
rect 9756 9742 9899 9744
rect 9756 9739 9833 9742
rect 9756 9712 9759 9739
rect 9788 9715 9833 9739
rect 9862 9715 9899 9742
rect 9788 9712 9899 9715
rect 9756 9711 9899 9712
rect 9935 9711 9959 9744
rect 9756 9698 9959 9711
rect 9102 9649 9134 9650
rect 9336 9647 9369 9650
rect 9302 9628 9370 9647
rect 9272 9616 9371 9628
rect 9994 9620 10066 9861
rect 10438 9620 10545 10049
rect 11000 10461 11107 11054
rect 11475 11003 11550 11054
rect 12516 11105 12538 11119
rect 12582 11105 12599 11142
rect 12516 11085 12599 11105
rect 12516 11019 12533 11085
rect 12587 11019 12599 11085
rect 11475 10960 11551 11003
rect 11479 10649 11551 10960
rect 12516 10995 12599 11019
rect 12516 10975 12592 10995
rect 12516 10956 12595 10975
rect 12175 10940 12247 10941
rect 12174 10932 12273 10940
rect 12174 10929 12226 10932
rect 12174 10894 12182 10929
rect 12207 10894 12226 10929
rect 12251 10894 12273 10932
rect 12174 10882 12273 10894
rect 12175 10863 12243 10882
rect 12176 10860 12209 10863
rect 12411 10860 12443 10861
rect 11586 10799 11789 10812
rect 11586 10766 11610 10799
rect 11646 10798 11789 10799
rect 11646 10795 11757 10798
rect 11646 10768 11683 10795
rect 11712 10771 11757 10795
rect 11786 10771 11789 10798
rect 11712 10768 11789 10771
rect 11646 10766 11789 10768
rect 11586 10753 11789 10766
rect 11586 10752 11687 10753
rect 11479 10607 11488 10649
rect 11537 10607 11551 10649
rect 11479 10586 11551 10607
rect 11479 10544 11489 10586
rect 11538 10544 11551 10586
rect 11479 10526 11551 10544
rect 11964 10690 11996 10697
rect 11964 10670 11971 10690
rect 11992 10670 11996 10690
rect 11964 10605 11996 10670
rect 12176 10661 12207 10860
rect 12408 10855 12443 10860
rect 12408 10835 12415 10855
rect 12435 10835 12443 10855
rect 12408 10827 12443 10835
rect 12176 10631 12182 10661
rect 12203 10631 12207 10661
rect 12176 10623 12207 10631
rect 12334 10605 12374 10606
rect 11964 10603 12376 10605
rect 11964 10577 12344 10603
rect 12370 10577 12376 10603
rect 11964 10569 12376 10577
rect 11964 10541 11996 10569
rect 12409 10549 12443 10827
rect 12525 10640 12595 10956
rect 14513 10941 14544 10942
rect 14513 10933 14558 10941
rect 13593 10910 13757 10917
rect 14513 10910 14523 10933
rect 13219 10895 14523 10910
rect 14548 10895 14558 10933
rect 13219 10877 14558 10895
rect 13224 10864 13260 10877
rect 13593 10874 13757 10877
rect 12634 10795 12837 10808
rect 12634 10762 12658 10795
rect 12694 10794 12837 10795
rect 12694 10791 12805 10794
rect 12694 10764 12731 10791
rect 12760 10767 12805 10791
rect 12834 10767 12837 10794
rect 12760 10764 12837 10767
rect 12694 10762 12837 10764
rect 12634 10749 12837 10762
rect 12634 10748 12735 10749
rect 11964 10521 11969 10541
rect 11990 10521 11996 10541
rect 11964 10514 11996 10521
rect 12387 10544 12443 10549
rect 12387 10524 12394 10544
rect 12414 10524 12443 10544
rect 12520 10634 12595 10640
rect 12520 10601 12528 10634
rect 12581 10601 12595 10634
rect 12520 10576 12595 10601
rect 12520 10543 12533 10576
rect 12586 10543 12595 10576
rect 12520 10534 12595 10543
rect 13012 10686 13044 10693
rect 13012 10666 13019 10686
rect 13040 10666 13044 10686
rect 13012 10601 13044 10666
rect 13224 10657 13255 10864
rect 13459 10856 13491 10857
rect 13456 10851 13491 10856
rect 13456 10831 13463 10851
rect 13483 10831 13491 10851
rect 13456 10823 13491 10831
rect 13224 10627 13230 10657
rect 13251 10627 13255 10657
rect 13224 10619 13255 10627
rect 13382 10601 13422 10602
rect 13012 10599 13424 10601
rect 13012 10573 13392 10599
rect 13418 10573 13424 10599
rect 13012 10565 13424 10573
rect 13012 10537 13044 10565
rect 13457 10545 13491 10823
rect 12520 10529 12578 10534
rect 12387 10517 12443 10524
rect 13012 10517 13017 10537
rect 13038 10517 13044 10537
rect 12387 10516 12422 10517
rect 13012 10510 13044 10517
rect 13435 10540 13491 10545
rect 13435 10520 13442 10540
rect 13462 10520 13491 10540
rect 13435 10513 13491 10520
rect 13435 10512 13470 10513
rect 11678 10461 11789 10465
rect 13461 10461 14761 10462
rect 11000 10443 14761 10461
rect 11000 10423 11686 10443
rect 11705 10423 11763 10443
rect 11782 10439 14761 10443
rect 11782 10423 12734 10439
rect 11000 10419 12734 10423
rect 12753 10419 12811 10439
rect 12830 10419 14761 10439
rect 11000 10405 14761 10419
rect 11000 9782 11107 10405
rect 12726 10402 12837 10405
rect 11486 10356 11550 10360
rect 11482 10350 11550 10356
rect 11482 10317 11499 10350
rect 11539 10317 11550 10350
rect 11482 10305 11550 10317
rect 12533 10319 12598 10341
rect 11482 10303 11539 10305
rect 11486 9942 11537 10303
rect 12533 10280 12550 10319
rect 12595 10280 12598 10319
rect 12174 10235 12209 10237
rect 12174 10226 12278 10235
rect 12174 10225 12225 10226
rect 12174 10205 12177 10225
rect 12202 10206 12225 10225
rect 12257 10206 12278 10226
rect 12202 10205 12278 10206
rect 12174 10198 12278 10205
rect 12174 10186 12209 10198
rect 11586 10120 11789 10133
rect 11586 10087 11610 10120
rect 11646 10119 11789 10120
rect 11646 10116 11757 10119
rect 11646 10089 11683 10116
rect 11712 10092 11757 10116
rect 11786 10092 11789 10119
rect 11712 10089 11789 10092
rect 11646 10087 11789 10089
rect 11586 10074 11789 10087
rect 11586 10073 11687 10074
rect 11964 10011 11996 10018
rect 11964 9991 11971 10011
rect 11992 9991 11996 10011
rect 11475 9933 11540 9942
rect 11475 9896 11485 9933
rect 11525 9899 11540 9933
rect 11964 9926 11996 9991
rect 12176 9982 12207 10186
rect 12411 10181 12443 10182
rect 12408 10176 12443 10181
rect 12408 10156 12415 10176
rect 12435 10156 12443 10176
rect 12408 10148 12443 10156
rect 12176 9952 12182 9982
rect 12203 9952 12207 9982
rect 12176 9944 12207 9952
rect 12334 9926 12374 9927
rect 11964 9924 12376 9926
rect 11525 9896 11542 9899
rect 11475 9877 11542 9896
rect 11475 9856 11489 9877
rect 11525 9856 11542 9877
rect 11475 9849 11542 9856
rect 11964 9898 12344 9924
rect 12370 9898 12376 9924
rect 11964 9890 12376 9898
rect 11964 9862 11996 9890
rect 12409 9870 12443 10148
rect 12533 9980 12598 10280
rect 14670 10241 14707 10262
rect 14670 10204 14681 10241
rect 14698 10217 14707 10241
rect 14698 10204 14708 10217
rect 14670 10194 14708 10204
rect 14671 10190 14708 10194
rect 14671 10184 14704 10190
rect 14081 10115 14284 10128
rect 14081 10082 14105 10115
rect 14141 10114 14284 10115
rect 14141 10111 14252 10114
rect 14141 10084 14178 10111
rect 14207 10087 14252 10111
rect 14281 10087 14284 10114
rect 14207 10084 14284 10087
rect 14141 10082 14284 10084
rect 14081 10069 14284 10082
rect 14081 10068 14182 10069
rect 14459 10006 14491 10013
rect 14459 9986 14466 10006
rect 14487 9986 14491 10006
rect 11964 9842 11969 9862
rect 11990 9842 11996 9862
rect 11964 9835 11996 9842
rect 12387 9865 12443 9870
rect 12387 9845 12394 9865
rect 12414 9845 12443 9865
rect 12387 9838 12443 9845
rect 12523 9969 12603 9980
rect 12523 9943 12540 9969
rect 12580 9943 12603 9969
rect 12523 9916 12603 9943
rect 12523 9890 12544 9916
rect 12584 9890 12603 9916
rect 14459 9921 14491 9986
rect 14671 9977 14702 10184
rect 14906 10176 14938 10177
rect 14903 10171 14938 10176
rect 14903 10151 14910 10171
rect 14930 10151 14938 10171
rect 14903 10143 14938 10151
rect 14671 9947 14677 9977
rect 14698 9947 14702 9977
rect 14671 9939 14702 9947
rect 14829 9921 14869 9922
rect 14459 9919 14871 9921
rect 12523 9871 12603 9890
rect 12523 9845 12547 9871
rect 12587 9845 12603 9871
rect 13636 9909 14073 9915
rect 13636 9886 13654 9909
rect 13680 9902 14073 9909
rect 13680 9886 14034 9902
rect 13636 9879 14034 9886
rect 14060 9879 14073 9902
rect 13636 9866 14073 9879
rect 14459 9893 14839 9919
rect 14865 9893 14871 9919
rect 14459 9885 14871 9893
rect 12387 9837 12422 9838
rect 12523 9833 12603 9845
rect 14459 9857 14491 9885
rect 14904 9865 14938 10143
rect 14459 9837 14464 9857
rect 14485 9837 14491 9857
rect 14459 9830 14491 9837
rect 14882 9860 14938 9865
rect 14882 9840 14889 9860
rect 14909 9840 14938 9860
rect 14882 9833 14938 9840
rect 14882 9832 14917 9833
rect 11678 9782 11789 9786
rect 13420 9782 14970 9785
rect 10998 9764 14970 9782
rect 10998 9744 11686 9764
rect 11705 9744 11763 9764
rect 11782 9759 14970 9764
rect 11782 9744 14181 9759
rect 10998 9739 14181 9744
rect 14200 9739 14258 9759
rect 14277 9739 14970 9759
rect 10998 9729 14970 9739
rect 10998 9726 11623 9729
rect 11810 9726 14970 9729
rect 9272 9578 9294 9616
rect 9319 9581 9338 9616
rect 9363 9581 9371 9616
rect 9319 9578 9371 9581
rect 9272 9570 9371 9578
rect 9298 9569 9370 9570
rect 8949 9543 9020 9559
rect 8949 9527 8969 9543
rect 8950 9497 8969 9527
rect 8952 9477 8969 9497
rect 8999 9497 9020 9543
rect 9992 9539 10070 9620
rect 10437 9565 10545 9620
rect 8999 9477 9019 9497
rect 8952 9458 9019 9477
rect 9992 9437 10071 9539
rect 6786 9414 6872 9423
rect 6786 9396 6805 9414
rect 6857 9396 6872 9414
rect 6786 9392 6872 9396
rect 9956 9419 10077 9437
rect 9956 9417 10027 9419
rect 9956 9376 9971 9417
rect 10008 9378 10027 9417
rect 10064 9378 10077 9419
rect 10008 9376 10077 9378
rect 9956 9366 10077 9376
rect 7261 9338 7372 9341
rect 6481 9337 8125 9338
rect 10438 9337 10545 9565
rect 11000 9498 11107 9726
rect 13420 9725 14970 9726
rect 14173 9722 14284 9725
rect 11468 9687 11589 9697
rect 11468 9685 11537 9687
rect 11468 9644 11481 9685
rect 11518 9646 11537 9685
rect 11574 9646 11589 9687
rect 11518 9644 11589 9646
rect 11468 9626 11589 9644
rect 11474 9524 11553 9626
rect 12526 9586 12593 9605
rect 12526 9566 12546 9586
rect 11000 9443 11108 9498
rect 11475 9443 11553 9524
rect 12525 9520 12546 9566
rect 12576 9566 12593 9586
rect 12576 9536 12595 9566
rect 12576 9520 12596 9536
rect 12525 9504 12596 9520
rect 12175 9493 12247 9494
rect 12174 9485 12273 9493
rect 12174 9482 12226 9485
rect 12174 9447 12182 9482
rect 12207 9447 12226 9482
rect 12251 9447 12273 9485
rect 6481 9334 9735 9337
rect 9922 9334 10547 9337
rect 6481 9324 10547 9334
rect 6481 9304 7268 9324
rect 7287 9304 7345 9324
rect 7364 9319 10547 9324
rect 7364 9304 9763 9319
rect 6481 9299 9763 9304
rect 9782 9299 9840 9319
rect 9859 9299 10547 9319
rect 6481 9281 10547 9299
rect 6481 9278 8125 9281
rect 9756 9277 9867 9281
rect 6628 9230 6663 9231
rect 6607 9223 6663 9230
rect 6607 9203 6636 9223
rect 6656 9203 6663 9223
rect 6607 9198 6663 9203
rect 7054 9226 7086 9233
rect 7054 9206 7060 9226
rect 7081 9206 7086 9226
rect 6607 8920 6641 9198
rect 7054 9178 7086 9206
rect 6674 9170 7086 9178
rect 6674 9144 6680 9170
rect 6706 9144 7086 9170
rect 6674 9142 7086 9144
rect 6676 9141 6716 9142
rect 6843 9116 6874 9124
rect 6843 9086 6847 9116
rect 6868 9086 6874 9116
rect 6607 8912 6642 8920
rect 6607 8892 6615 8912
rect 6635 8892 6642 8912
rect 6607 8887 6642 8892
rect 6607 8886 6639 8887
rect 6843 8885 6874 9086
rect 7054 9077 7086 9142
rect 7054 9057 7058 9077
rect 7079 9057 7086 9077
rect 7054 9050 7086 9057
rect 7648 9217 7741 9224
rect 7648 9176 7672 9217
rect 7726 9176 7741 9217
rect 7363 8994 7464 8995
rect 7261 8981 7464 8994
rect 7261 8979 7404 8981
rect 7261 8976 7338 8979
rect 7261 8949 7264 8976
rect 7293 8952 7338 8976
rect 7367 8952 7404 8979
rect 7293 8949 7404 8952
rect 7261 8948 7404 8949
rect 7440 8948 7464 8981
rect 7261 8935 7464 8948
rect 7648 8803 7741 9176
rect 8942 9218 9022 9230
rect 9123 9225 9158 9226
rect 8942 9192 8958 9218
rect 8998 9192 9022 9218
rect 8942 9173 9022 9192
rect 8942 9147 8961 9173
rect 9001 9147 9022 9173
rect 8942 9120 9022 9147
rect 8942 9094 8965 9120
rect 9005 9094 9022 9120
rect 8942 9083 9022 9094
rect 9102 9218 9158 9225
rect 9102 9198 9131 9218
rect 9151 9198 9158 9218
rect 9102 9193 9158 9198
rect 9549 9221 9581 9228
rect 9549 9201 9555 9221
rect 9576 9201 9581 9221
rect 7648 8759 7666 8803
rect 7726 8759 7741 8803
rect 7648 8744 7741 8759
rect 8947 8783 9012 9083
rect 9102 8915 9136 9193
rect 9549 9173 9581 9201
rect 9169 9165 9581 9173
rect 9169 9139 9175 9165
rect 9201 9139 9581 9165
rect 10003 9207 10070 9214
rect 10003 9186 10020 9207
rect 10056 9186 10070 9207
rect 10003 9167 10070 9186
rect 10003 9164 10020 9167
rect 9169 9137 9581 9139
rect 9171 9136 9211 9137
rect 9338 9111 9369 9119
rect 9338 9081 9342 9111
rect 9363 9081 9369 9111
rect 9102 8907 9137 8915
rect 9102 8887 9110 8907
rect 9130 8887 9137 8907
rect 9102 8882 9137 8887
rect 9102 8881 9134 8882
rect 9338 8877 9369 9081
rect 9549 9072 9581 9137
rect 10005 9130 10020 9164
rect 10060 9130 10070 9167
rect 10005 9121 10070 9130
rect 9549 9052 9553 9072
rect 9574 9052 9581 9072
rect 9549 9045 9581 9052
rect 9858 8989 9959 8990
rect 9756 8976 9959 8989
rect 9756 8974 9899 8976
rect 9756 8971 9833 8974
rect 9756 8944 9759 8971
rect 9788 8947 9833 8971
rect 9862 8947 9899 8974
rect 9788 8944 9899 8947
rect 9756 8943 9899 8944
rect 9935 8943 9959 8976
rect 9756 8930 9959 8943
rect 9336 8865 9371 8877
rect 9267 8858 9371 8865
rect 9267 8857 9343 8858
rect 9267 8837 9288 8857
rect 9320 8838 9343 8857
rect 9368 8838 9371 8858
rect 9320 8837 9371 8838
rect 9267 8828 9371 8837
rect 9336 8826 9371 8828
rect 8947 8744 8950 8783
rect 8995 8744 9012 8783
rect 10008 8760 10059 9121
rect 10006 8758 10063 8760
rect 8947 8722 9012 8744
rect 9995 8746 10063 8758
rect 9995 8713 10006 8746
rect 10046 8713 10063 8746
rect 9995 8707 10063 8713
rect 9995 8703 10059 8707
rect 8708 8658 8819 8661
rect 10438 8658 10545 9281
rect 6514 8644 10545 8658
rect 6514 8624 8715 8644
rect 8734 8624 8792 8644
rect 8811 8640 10545 8644
rect 8811 8624 9763 8640
rect 6514 8620 9763 8624
rect 9782 8620 9840 8640
rect 9859 8620 10545 8640
rect 6514 8602 10545 8620
rect 6514 8601 8084 8602
rect 9756 8598 9867 8602
rect 8075 8550 8110 8551
rect 8054 8543 8110 8550
rect 8054 8523 8083 8543
rect 8103 8523 8110 8543
rect 8054 8518 8110 8523
rect 8501 8546 8533 8553
rect 9123 8546 9158 8547
rect 8501 8526 8507 8546
rect 8528 8526 8533 8546
rect 9102 8539 9158 8546
rect 8967 8529 9025 8534
rect 7654 8463 7736 8492
rect 7654 8422 7679 8463
rect 7715 8422 7736 8463
rect 7841 8483 7905 8502
rect 7841 8444 7858 8483
rect 7892 8444 7905 8483
rect 7841 8425 7905 8444
rect 7654 8107 7736 8422
rect 7646 8062 7736 8107
rect 7843 8080 7905 8425
rect 8054 8240 8088 8518
rect 8501 8498 8533 8526
rect 8121 8490 8533 8498
rect 8121 8464 8127 8490
rect 8153 8464 8533 8490
rect 8121 8462 8533 8464
rect 8123 8461 8163 8462
rect 8290 8436 8321 8444
rect 8290 8406 8294 8436
rect 8315 8406 8321 8436
rect 8054 8232 8089 8240
rect 8054 8212 8062 8232
rect 8082 8212 8089 8232
rect 8054 8207 8089 8212
rect 8054 8206 8086 8207
rect 8290 8199 8321 8406
rect 8501 8397 8533 8462
rect 8501 8377 8505 8397
rect 8526 8377 8533 8397
rect 8501 8370 8533 8377
rect 8950 8520 9025 8529
rect 8950 8487 8959 8520
rect 9012 8487 9025 8520
rect 8950 8462 9025 8487
rect 8950 8429 8964 8462
rect 9017 8429 9025 8462
rect 8950 8423 9025 8429
rect 9102 8519 9131 8539
rect 9151 8519 9158 8539
rect 9102 8514 9158 8519
rect 9549 8542 9581 8549
rect 9549 8522 9555 8542
rect 9576 8522 9581 8542
rect 8810 8314 8911 8315
rect 8708 8301 8911 8314
rect 8708 8299 8851 8301
rect 8708 8296 8785 8299
rect 8708 8269 8711 8296
rect 8740 8272 8785 8296
rect 8814 8272 8851 8299
rect 8740 8269 8851 8272
rect 8708 8268 8851 8269
rect 8887 8268 8911 8301
rect 8708 8255 8911 8268
rect 8285 8181 8321 8199
rect 8252 8180 8321 8181
rect 8232 8168 8321 8180
rect 8232 8130 8244 8168
rect 8269 8133 8288 8168
rect 8313 8133 8321 8168
rect 8950 8157 9020 8423
rect 9102 8236 9136 8514
rect 9549 8494 9581 8522
rect 9169 8486 9581 8494
rect 9169 8460 9175 8486
rect 9201 8460 9581 8486
rect 9169 8458 9581 8460
rect 9171 8457 9211 8458
rect 9338 8432 9369 8440
rect 9338 8402 9342 8432
rect 9363 8402 9369 8432
rect 9102 8228 9137 8236
rect 9102 8208 9110 8228
rect 9130 8208 9137 8228
rect 9102 8203 9137 8208
rect 9338 8203 9369 8402
rect 9549 8393 9581 8458
rect 9549 8373 9553 8393
rect 9574 8373 9581 8393
rect 9549 8366 9581 8373
rect 9994 8519 10066 8537
rect 9994 8477 10007 8519
rect 10056 8477 10066 8519
rect 9994 8456 10066 8477
rect 9994 8414 10008 8456
rect 10057 8414 10066 8456
rect 9858 8310 9959 8311
rect 9756 8297 9959 8310
rect 9756 8295 9899 8297
rect 9756 8292 9833 8295
rect 9756 8265 9759 8292
rect 9788 8268 9833 8292
rect 9862 8268 9899 8295
rect 9788 8265 9899 8268
rect 9756 8264 9899 8265
rect 9935 8264 9959 8297
rect 9756 8251 9959 8264
rect 9102 8202 9134 8203
rect 9336 8200 9369 8203
rect 9302 8181 9370 8200
rect 8269 8130 8321 8133
rect 8232 8122 8321 8130
rect 8941 8128 9020 8157
rect 9272 8169 9371 8181
rect 9272 8131 9294 8169
rect 9319 8134 9338 8169
rect 9363 8134 9371 8169
rect 9319 8131 9371 8134
rect 8248 8121 8320 8122
rect 7842 8071 7916 8080
rect 7646 8029 7730 8062
rect 7646 8001 7661 8029
rect 7705 8001 7730 8029
rect 7646 7972 7730 8001
rect 7842 8023 7856 8071
rect 7893 8023 7916 8071
rect 7842 7995 7916 8023
rect 7646 7944 7658 7972
rect 7702 7944 7730 7972
rect 7646 7933 7730 7944
rect 8941 7945 9018 8128
rect 9272 8123 9371 8131
rect 9298 8122 9370 8123
rect 9994 8120 10066 8414
rect 10438 8142 10545 8602
rect 11000 9014 11107 9443
rect 11479 9202 11551 9443
rect 12174 9435 12273 9447
rect 12175 9416 12243 9435
rect 12176 9413 12209 9416
rect 12411 9413 12443 9414
rect 11586 9352 11789 9365
rect 11586 9319 11610 9352
rect 11646 9351 11789 9352
rect 11646 9348 11757 9351
rect 11646 9321 11683 9348
rect 11712 9324 11757 9348
rect 11786 9324 11789 9351
rect 11712 9321 11789 9324
rect 11646 9319 11789 9321
rect 11586 9306 11789 9319
rect 11586 9305 11687 9306
rect 11479 9160 11488 9202
rect 11537 9160 11551 9202
rect 11479 9139 11551 9160
rect 11479 9097 11489 9139
rect 11538 9097 11551 9139
rect 11479 9079 11551 9097
rect 11964 9243 11996 9250
rect 11964 9223 11971 9243
rect 11992 9223 11996 9243
rect 11964 9158 11996 9223
rect 12176 9214 12207 9413
rect 12408 9408 12443 9413
rect 12408 9388 12415 9408
rect 12435 9388 12443 9408
rect 12408 9380 12443 9388
rect 12176 9184 12182 9214
rect 12203 9184 12207 9214
rect 12176 9176 12207 9184
rect 12334 9158 12374 9159
rect 11964 9156 12376 9158
rect 11964 9130 12344 9156
rect 12370 9130 12376 9156
rect 11964 9122 12376 9130
rect 11964 9094 11996 9122
rect 12409 9102 12443 9380
rect 12525 9193 12595 9504
rect 13222 9495 14564 9500
rect 13222 9493 14521 9495
rect 13219 9467 14521 9493
rect 14549 9467 14564 9495
rect 13219 9459 14564 9467
rect 13219 9434 13258 9459
rect 13219 9417 13260 9434
rect 13219 9410 13258 9417
rect 12634 9348 12837 9361
rect 12634 9315 12658 9348
rect 12694 9347 12837 9348
rect 12694 9344 12805 9347
rect 12694 9317 12731 9344
rect 12760 9320 12805 9344
rect 12834 9320 12837 9347
rect 12760 9317 12837 9320
rect 12694 9315 12837 9317
rect 12634 9302 12837 9315
rect 12634 9301 12735 9302
rect 11964 9074 11969 9094
rect 11990 9074 11996 9094
rect 11964 9067 11996 9074
rect 12387 9097 12443 9102
rect 12387 9077 12394 9097
rect 12414 9077 12443 9097
rect 12520 9187 12595 9193
rect 12520 9154 12528 9187
rect 12581 9154 12595 9187
rect 12520 9129 12595 9154
rect 12520 9096 12533 9129
rect 12586 9096 12595 9129
rect 12520 9087 12595 9096
rect 13012 9239 13044 9246
rect 13012 9219 13019 9239
rect 13040 9219 13044 9239
rect 13012 9154 13044 9219
rect 13224 9210 13255 9410
rect 13459 9409 13491 9410
rect 13456 9404 13491 9409
rect 13456 9384 13463 9404
rect 13483 9384 13491 9404
rect 13456 9376 13491 9384
rect 13224 9180 13230 9210
rect 13251 9180 13255 9210
rect 13224 9172 13255 9180
rect 13382 9154 13422 9155
rect 13012 9152 13424 9154
rect 13012 9126 13392 9152
rect 13418 9126 13424 9152
rect 13012 9118 13424 9126
rect 13012 9090 13044 9118
rect 13457 9098 13491 9376
rect 12520 9082 12578 9087
rect 12387 9070 12443 9077
rect 13012 9070 13017 9090
rect 13038 9070 13044 9090
rect 12387 9069 12422 9070
rect 13012 9063 13044 9070
rect 13435 9093 13491 9098
rect 13435 9073 13442 9093
rect 13462 9073 13491 9093
rect 13435 9066 13491 9073
rect 13435 9065 13470 9066
rect 11678 9014 11789 9018
rect 13553 9014 14543 9015
rect 11000 8996 14543 9014
rect 11000 8976 11686 8996
rect 11705 8976 11763 8996
rect 11782 8992 14543 8996
rect 11782 8976 12734 8992
rect 11000 8972 12734 8976
rect 12753 8972 12811 8992
rect 12830 8972 14543 8992
rect 11000 8958 14543 8972
rect 11000 8335 11107 8958
rect 12726 8955 12837 8958
rect 11486 8909 11550 8913
rect 11482 8903 11550 8909
rect 11482 8870 11499 8903
rect 11539 8870 11550 8903
rect 11482 8858 11550 8870
rect 12533 8872 12598 8894
rect 11482 8856 11539 8858
rect 11486 8495 11537 8856
rect 12533 8833 12550 8872
rect 12595 8833 12598 8872
rect 12174 8788 12209 8790
rect 12174 8779 12278 8788
rect 12174 8778 12225 8779
rect 12174 8758 12177 8778
rect 12202 8759 12225 8778
rect 12257 8759 12278 8779
rect 12202 8758 12278 8759
rect 12174 8751 12278 8758
rect 12174 8739 12209 8751
rect 11586 8673 11789 8686
rect 11586 8640 11610 8673
rect 11646 8672 11789 8673
rect 11646 8669 11757 8672
rect 11646 8642 11683 8669
rect 11712 8645 11757 8669
rect 11786 8645 11789 8672
rect 11712 8642 11789 8645
rect 11646 8640 11789 8642
rect 11586 8627 11789 8640
rect 11586 8626 11687 8627
rect 11964 8564 11996 8571
rect 11964 8544 11971 8564
rect 11992 8544 11996 8564
rect 11475 8486 11540 8495
rect 11475 8449 11485 8486
rect 11525 8452 11540 8486
rect 11964 8479 11996 8544
rect 12176 8535 12207 8739
rect 12411 8734 12443 8735
rect 12408 8729 12443 8734
rect 12408 8709 12415 8729
rect 12435 8709 12443 8729
rect 12408 8701 12443 8709
rect 12176 8505 12182 8535
rect 12203 8505 12207 8535
rect 12176 8497 12207 8505
rect 12334 8479 12374 8480
rect 11964 8477 12376 8479
rect 11525 8449 11542 8452
rect 11475 8430 11542 8449
rect 11475 8409 11489 8430
rect 11525 8409 11542 8430
rect 11475 8402 11542 8409
rect 11964 8451 12344 8477
rect 12370 8451 12376 8477
rect 11964 8443 12376 8451
rect 11964 8415 11996 8443
rect 12409 8423 12443 8701
rect 12533 8533 12598 8833
rect 11964 8395 11969 8415
rect 11990 8395 11996 8415
rect 11964 8388 11996 8395
rect 12387 8418 12443 8423
rect 12387 8398 12394 8418
rect 12414 8398 12443 8418
rect 12387 8391 12443 8398
rect 12523 8522 12603 8533
rect 12523 8496 12540 8522
rect 12580 8496 12603 8522
rect 12523 8469 12603 8496
rect 15075 8472 15124 13653
rect 16123 13065 16210 14220
rect 26018 14167 26117 14174
rect 26018 14112 26034 14167
rect 26100 14112 26117 14167
rect 26018 14098 26117 14112
rect 24758 14056 24879 14074
rect 24758 13983 24772 14056
rect 24842 13983 24879 14056
rect 20713 13845 20778 13983
rect 20663 13827 20784 13845
rect 20663 13825 20734 13827
rect 20663 13784 20678 13825
rect 20715 13786 20734 13825
rect 20771 13786 20784 13827
rect 20715 13784 20784 13786
rect 20663 13774 20784 13784
rect 17179 13745 18657 13747
rect 21145 13745 21252 13748
rect 17179 13727 21254 13745
rect 17179 13707 20470 13727
rect 20489 13707 20547 13727
rect 20566 13707 21254 13727
rect 17179 13689 21254 13707
rect 18612 13688 18819 13689
rect 20463 13685 20574 13689
rect 19649 13626 19729 13638
rect 19830 13633 19865 13634
rect 19649 13600 19665 13626
rect 19705 13600 19729 13626
rect 19649 13581 19729 13600
rect 19649 13555 19668 13581
rect 19708 13555 19729 13581
rect 19649 13528 19729 13555
rect 19649 13502 19672 13528
rect 19712 13502 19729 13528
rect 19649 13491 19729 13502
rect 19809 13626 19865 13633
rect 19809 13606 19838 13626
rect 19858 13606 19865 13626
rect 19809 13601 19865 13606
rect 20256 13629 20288 13636
rect 20256 13609 20262 13629
rect 20283 13609 20288 13629
rect 19654 13191 19719 13491
rect 19809 13323 19843 13601
rect 20256 13581 20288 13609
rect 19876 13573 20288 13581
rect 19876 13547 19882 13573
rect 19908 13547 20288 13573
rect 20710 13615 20777 13622
rect 20710 13594 20727 13615
rect 20763 13594 20777 13615
rect 20710 13575 20777 13594
rect 20710 13572 20727 13575
rect 19876 13545 20288 13547
rect 19878 13544 19918 13545
rect 20045 13519 20076 13527
rect 20045 13489 20049 13519
rect 20070 13489 20076 13519
rect 19809 13315 19844 13323
rect 19809 13295 19817 13315
rect 19837 13295 19844 13315
rect 19809 13290 19844 13295
rect 19809 13289 19841 13290
rect 20045 13285 20076 13489
rect 20256 13480 20288 13545
rect 20712 13538 20727 13572
rect 20767 13538 20777 13575
rect 20712 13529 20777 13538
rect 20256 13460 20260 13480
rect 20281 13460 20288 13480
rect 20256 13453 20288 13460
rect 20565 13397 20666 13398
rect 20463 13384 20666 13397
rect 20463 13382 20606 13384
rect 20463 13379 20540 13382
rect 20463 13352 20466 13379
rect 20495 13355 20540 13379
rect 20569 13355 20606 13382
rect 20495 13352 20606 13355
rect 20463 13351 20606 13352
rect 20642 13351 20666 13384
rect 20463 13338 20666 13351
rect 20043 13273 20078 13285
rect 19974 13266 20078 13273
rect 19974 13265 20050 13266
rect 19974 13245 19995 13265
rect 20027 13246 20050 13265
rect 20075 13246 20078 13266
rect 20027 13245 20078 13246
rect 19974 13236 20078 13245
rect 20043 13234 20078 13236
rect 19654 13152 19657 13191
rect 19702 13152 19719 13191
rect 20715 13168 20766 13529
rect 20713 13166 20770 13168
rect 19654 13130 19719 13152
rect 20702 13154 20770 13166
rect 20702 13121 20713 13154
rect 20753 13121 20770 13154
rect 20702 13115 20770 13121
rect 20702 13111 20766 13115
rect 19415 13066 19526 13069
rect 21145 13066 21252 13689
rect 15189 8664 15392 8677
rect 15189 8631 15213 8664
rect 15249 8663 15392 8664
rect 15249 8660 15360 8663
rect 15249 8633 15286 8660
rect 15315 8636 15360 8660
rect 15389 8636 15392 8663
rect 15315 8633 15392 8636
rect 15249 8631 15392 8633
rect 15189 8618 15392 8631
rect 15189 8617 15290 8618
rect 15567 8555 15599 8562
rect 15567 8535 15574 8555
rect 15595 8535 15599 8555
rect 12523 8443 12544 8469
rect 12584 8443 12603 8469
rect 12523 8424 12603 8443
rect 15074 8462 15185 8472
rect 15074 8461 15139 8462
rect 15074 8437 15082 8461
rect 15106 8438 15139 8461
rect 15163 8438 15185 8462
rect 15106 8437 15185 8438
rect 15074 8430 15185 8437
rect 15567 8470 15599 8535
rect 15779 8526 15810 8726
rect 16014 8725 16046 8726
rect 16011 8720 16046 8725
rect 16011 8700 16018 8720
rect 16038 8700 16046 8720
rect 16011 8692 16046 8700
rect 15779 8496 15785 8526
rect 15806 8496 15810 8526
rect 15779 8488 15810 8496
rect 15937 8470 15977 8471
rect 15567 8468 15979 8470
rect 15567 8442 15947 8468
rect 15973 8442 15979 8468
rect 15567 8434 15979 8442
rect 12523 8398 12547 8424
rect 12587 8398 12603 8424
rect 12387 8390 12422 8391
rect 12523 8386 12603 8398
rect 15567 8406 15599 8434
rect 16012 8414 16046 8692
rect 15567 8386 15572 8406
rect 15593 8386 15599 8406
rect 15567 8379 15599 8386
rect 15778 8406 15812 8413
rect 15778 8384 15785 8406
rect 15809 8384 15812 8406
rect 11678 8335 11789 8339
rect 13433 8335 13640 8336
rect 10998 8330 15073 8335
rect 10998 8317 15392 8330
rect 10998 8297 11686 8317
rect 11705 8297 11763 8317
rect 11782 8308 15392 8317
rect 11782 8297 15289 8308
rect 10998 8288 15289 8297
rect 15308 8288 15366 8308
rect 15385 8288 15392 8308
rect 10998 8279 15392 8288
rect 9994 8082 10070 8120
rect 10438 8082 10551 8142
rect 11000 8106 11107 8279
rect 13595 8277 15392 8279
rect 15281 8271 15392 8277
rect 11468 8240 11589 8250
rect 11468 8238 11537 8240
rect 11468 8197 11481 8238
rect 11518 8199 11537 8238
rect 11574 8199 11589 8240
rect 11518 8197 11589 8199
rect 11468 8179 11589 8197
rect 15616 8229 15668 8260
rect 15616 8195 15625 8229
rect 15654 8195 15668 8229
rect 10005 7981 10070 8082
rect 8941 7902 8958 7945
rect 5874 7853 5889 7887
rect 5918 7853 5926 7887
rect 8946 7897 8958 7902
rect 9004 7897 9018 7945
rect 8946 7875 9018 7897
rect 10003 7935 10070 7981
rect 10440 7943 10551 8082
rect 5874 7827 5926 7853
rect 10003 7843 10068 7935
rect 10435 7916 10551 7943
rect 10991 8079 11107 8106
rect 11474 8087 11539 8179
rect 15616 8169 15668 8195
rect 15778 8178 15812 8384
rect 15990 8409 16046 8414
rect 15990 8389 15997 8409
rect 16017 8389 16046 8409
rect 15990 8382 16046 8389
rect 15990 8381 16025 8382
rect 10991 7940 11102 8079
rect 11472 8041 11539 8087
rect 12524 8125 12596 8147
rect 12524 8077 12538 8125
rect 12584 8120 12596 8125
rect 15616 8135 15624 8169
rect 15653 8135 15668 8169
rect 12584 8077 12601 8120
rect 11472 7940 11537 8041
rect 5874 7793 5888 7827
rect 5917 7793 5926 7827
rect 5874 7762 5926 7793
rect 9953 7825 10074 7843
rect 9953 7823 10024 7825
rect 9953 7782 9968 7823
rect 10005 7784 10024 7823
rect 10061 7784 10074 7825
rect 10005 7782 10074 7784
rect 9953 7772 10074 7782
rect 6150 7745 6261 7751
rect 6150 7743 7947 7745
rect 10435 7743 10542 7916
rect 10991 7880 11104 7940
rect 11472 7902 11548 7940
rect 6150 7734 10544 7743
rect 6150 7714 6157 7734
rect 6176 7714 6234 7734
rect 6253 7725 10544 7734
rect 6253 7714 9760 7725
rect 6150 7705 9760 7714
rect 9779 7705 9837 7725
rect 9856 7705 10544 7725
rect 6150 7692 10544 7705
rect 6469 7687 10544 7692
rect 7902 7686 8109 7687
rect 9753 7683 9864 7687
rect 5517 7640 5552 7641
rect 5496 7633 5552 7640
rect 5496 7613 5525 7633
rect 5545 7613 5552 7633
rect 5496 7608 5552 7613
rect 5943 7636 5975 7643
rect 5943 7616 5949 7636
rect 5970 7616 5975 7636
rect 5496 7330 5530 7608
rect 5943 7588 5975 7616
rect 8939 7624 9019 7636
rect 9120 7631 9155 7632
rect 8939 7598 8955 7624
rect 8995 7598 9019 7624
rect 5563 7580 5975 7588
rect 5563 7554 5569 7580
rect 5595 7554 5975 7580
rect 5563 7552 5975 7554
rect 5565 7551 5605 7552
rect 5732 7526 5763 7534
rect 5732 7496 5736 7526
rect 5757 7496 5763 7526
rect 5496 7322 5531 7330
rect 5496 7302 5504 7322
rect 5524 7302 5531 7322
rect 5732 7311 5763 7496
rect 5943 7487 5975 7552
rect 6357 7585 6468 7592
rect 6357 7584 6436 7585
rect 6357 7560 6379 7584
rect 6403 7561 6436 7584
rect 6460 7561 6468 7585
rect 6403 7560 6468 7561
rect 6357 7550 6468 7560
rect 8939 7579 9019 7598
rect 8939 7553 8958 7579
rect 8998 7553 9019 7579
rect 6418 7533 6467 7550
rect 8939 7526 9019 7553
rect 8939 7500 8962 7526
rect 9002 7500 9019 7526
rect 8939 7489 9019 7500
rect 9099 7624 9155 7631
rect 9099 7604 9128 7624
rect 9148 7604 9155 7624
rect 9099 7599 9155 7604
rect 9546 7627 9578 7634
rect 9546 7607 9552 7627
rect 9573 7607 9578 7627
rect 5943 7467 5947 7487
rect 5968 7467 5975 7487
rect 5943 7460 5975 7467
rect 6252 7404 6353 7405
rect 6150 7391 6353 7404
rect 6150 7389 6293 7391
rect 6150 7386 6227 7389
rect 6150 7359 6153 7386
rect 6182 7362 6227 7386
rect 6256 7362 6293 7389
rect 6182 7359 6293 7362
rect 6150 7358 6293 7359
rect 6329 7358 6353 7391
rect 6150 7345 6353 7358
rect 5496 7297 5531 7302
rect 5496 7296 5528 7297
rect 5730 7234 5764 7311
rect 4363 5831 4960 5835
rect 1463 5753 1498 5755
rect 1463 5744 1567 5753
rect 1463 5743 1514 5744
rect 1463 5723 1466 5743
rect 1491 5724 1514 5743
rect 1546 5724 1567 5744
rect 1491 5723 1567 5724
rect 1463 5716 1567 5723
rect 1463 5704 1498 5716
rect 875 5638 1078 5651
rect 875 5605 899 5638
rect 935 5637 1078 5638
rect 935 5634 1046 5637
rect 935 5607 972 5634
rect 1001 5610 1046 5634
rect 1075 5610 1078 5637
rect 1001 5607 1078 5610
rect 935 5605 1078 5607
rect 875 5592 1078 5605
rect 875 5591 976 5592
rect 1253 5529 1285 5536
rect 1253 5509 1260 5529
rect 1281 5509 1285 5529
rect 764 5451 829 5460
rect 764 5414 774 5451
rect 814 5417 829 5451
rect 1253 5444 1285 5509
rect 1465 5500 1496 5704
rect 1700 5699 1732 5700
rect 1697 5694 1732 5699
rect 1697 5674 1704 5694
rect 1724 5674 1732 5694
rect 1697 5666 1732 5674
rect 1465 5470 1471 5500
rect 1492 5470 1496 5500
rect 1465 5462 1496 5470
rect 1623 5444 1663 5445
rect 1253 5442 1665 5444
rect 814 5414 831 5417
rect 764 5395 831 5414
rect 764 5374 778 5395
rect 814 5374 831 5395
rect 764 5367 831 5374
rect 1253 5416 1633 5442
rect 1659 5416 1665 5442
rect 1253 5408 1665 5416
rect 1253 5380 1285 5408
rect 1698 5388 1732 5666
rect 1822 5498 1887 5798
rect 4000 5786 4960 5831
rect 5067 6174 5103 6802
rect 4000 5782 4413 5786
rect 4000 5693 4034 5782
rect 4238 5696 4270 5697
rect 3413 5635 3616 5648
rect 3413 5602 3437 5635
rect 3473 5634 3616 5635
rect 3473 5631 3584 5634
rect 3473 5604 3510 5631
rect 3539 5607 3584 5631
rect 3613 5607 3616 5634
rect 3539 5604 3616 5607
rect 3473 5602 3616 5604
rect 3413 5589 3616 5602
rect 3413 5588 3514 5589
rect 3791 5526 3823 5533
rect 3791 5506 3798 5526
rect 3819 5506 3823 5526
rect 1253 5360 1258 5380
rect 1279 5360 1285 5380
rect 1253 5353 1285 5360
rect 1676 5383 1732 5388
rect 1676 5363 1683 5383
rect 1703 5363 1732 5383
rect 1676 5356 1732 5363
rect 1812 5487 1892 5498
rect 1812 5461 1829 5487
rect 1869 5461 1892 5487
rect 1812 5434 1892 5461
rect 1812 5408 1833 5434
rect 1873 5408 1892 5434
rect 1812 5389 1892 5408
rect 1812 5363 1836 5389
rect 1876 5363 1892 5389
rect 1676 5355 1711 5356
rect 1812 5351 1892 5363
rect 3791 5441 3823 5506
rect 4003 5497 4034 5693
rect 4235 5691 4270 5696
rect 4235 5671 4242 5691
rect 4262 5671 4270 5691
rect 4235 5663 4270 5671
rect 4003 5467 4009 5497
rect 4030 5467 4034 5497
rect 4003 5459 4034 5467
rect 4161 5441 4201 5442
rect 3791 5439 4203 5441
rect 3791 5413 4171 5439
rect 4197 5413 4203 5439
rect 3791 5405 4203 5413
rect 3791 5377 3823 5405
rect 4236 5385 4270 5663
rect 3791 5357 3796 5377
rect 3817 5357 3823 5377
rect 3791 5350 3823 5357
rect 4214 5380 4270 5385
rect 4214 5360 4221 5380
rect 4241 5360 4270 5380
rect 4214 5353 4270 5360
rect 4214 5352 4249 5353
rect 967 5300 1078 5304
rect 2722 5300 2929 5301
rect 3505 5300 3616 5301
rect 287 5282 4353 5300
rect 287 5262 975 5282
rect 994 5262 1052 5282
rect 1071 5279 4353 5282
rect 1071 5262 3513 5279
rect 287 5259 3513 5262
rect 3532 5259 3590 5279
rect 3609 5259 4353 5279
rect 287 5244 4353 5259
rect 289 5056 396 5244
rect 2884 5242 4353 5244
rect 757 5205 878 5215
rect 757 5203 826 5205
rect 757 5162 770 5203
rect 807 5164 826 5203
rect 863 5164 878 5205
rect 807 5162 878 5164
rect 757 5144 878 5162
rect 289 5052 397 5056
rect 763 5052 840 5144
rect 1813 5140 1889 5156
rect 1813 5117 1828 5140
rect 290 4459 397 5052
rect 765 5001 840 5052
rect 1806 5103 1828 5117
rect 1872 5103 1889 5140
rect 1806 5083 1889 5103
rect 1806 5017 1823 5083
rect 1877 5017 1889 5083
rect 765 4958 841 5001
rect 769 4647 841 4958
rect 1806 4993 1889 5017
rect 1806 4973 1882 4993
rect 1806 4954 1885 4973
rect 1465 4938 1537 4939
rect 1464 4930 1563 4938
rect 1464 4927 1516 4930
rect 1464 4892 1472 4927
rect 1497 4892 1516 4927
rect 1541 4892 1563 4930
rect 1464 4880 1563 4892
rect 1465 4861 1533 4880
rect 1466 4858 1499 4861
rect 1701 4858 1733 4859
rect 876 4797 1079 4810
rect 876 4764 900 4797
rect 936 4796 1079 4797
rect 936 4793 1047 4796
rect 936 4766 973 4793
rect 1002 4769 1047 4793
rect 1076 4769 1079 4796
rect 1002 4766 1079 4769
rect 936 4764 1079 4766
rect 876 4751 1079 4764
rect 876 4750 977 4751
rect 769 4605 778 4647
rect 827 4605 841 4647
rect 769 4584 841 4605
rect 769 4542 779 4584
rect 828 4542 841 4584
rect 769 4524 841 4542
rect 1254 4688 1286 4695
rect 1254 4668 1261 4688
rect 1282 4668 1286 4688
rect 1254 4603 1286 4668
rect 1466 4659 1497 4858
rect 1698 4853 1733 4858
rect 1698 4833 1705 4853
rect 1725 4833 1733 4853
rect 1698 4825 1733 4833
rect 1466 4629 1472 4659
rect 1493 4629 1497 4659
rect 1466 4621 1497 4629
rect 1624 4603 1664 4604
rect 1254 4601 1666 4603
rect 1254 4575 1634 4601
rect 1660 4575 1666 4601
rect 1254 4567 1666 4575
rect 1254 4539 1286 4567
rect 1699 4547 1733 4825
rect 1815 4638 1885 4954
rect 3803 4939 3834 4940
rect 3803 4931 3848 4939
rect 2883 4908 3047 4915
rect 3803 4908 3813 4931
rect 2509 4893 3813 4908
rect 3838 4893 3848 4931
rect 5067 4934 5101 6174
rect 5067 4930 5297 4934
rect 5067 4904 5266 4930
rect 5291 4904 5297 4930
rect 5067 4896 5297 4904
rect 2509 4875 3848 4893
rect 2514 4862 2550 4875
rect 2883 4872 3047 4875
rect 1924 4793 2127 4806
rect 1924 4760 1948 4793
rect 1984 4792 2127 4793
rect 1984 4789 2095 4792
rect 1984 4762 2021 4789
rect 2050 4765 2095 4789
rect 2124 4765 2127 4792
rect 2050 4762 2127 4765
rect 1984 4760 2127 4762
rect 1924 4747 2127 4760
rect 1924 4746 2025 4747
rect 1254 4519 1259 4539
rect 1280 4519 1286 4539
rect 1254 4512 1286 4519
rect 1677 4542 1733 4547
rect 1677 4522 1684 4542
rect 1704 4522 1733 4542
rect 1810 4632 1885 4638
rect 1810 4599 1818 4632
rect 1871 4599 1885 4632
rect 1810 4574 1885 4599
rect 1810 4541 1823 4574
rect 1876 4541 1885 4574
rect 1810 4532 1885 4541
rect 2302 4684 2334 4691
rect 2302 4664 2309 4684
rect 2330 4664 2334 4684
rect 2302 4599 2334 4664
rect 2514 4655 2545 4862
rect 2749 4854 2781 4855
rect 2746 4849 2781 4854
rect 2746 4829 2753 4849
rect 2773 4829 2781 4849
rect 2746 4821 2781 4829
rect 2514 4625 2520 4655
rect 2541 4625 2545 4655
rect 2514 4617 2545 4625
rect 2672 4599 2712 4600
rect 2302 4597 2714 4599
rect 2302 4571 2682 4597
rect 2708 4571 2714 4597
rect 2302 4563 2714 4571
rect 2302 4535 2334 4563
rect 2747 4543 2781 4821
rect 4826 4799 5029 4812
rect 4826 4766 4850 4799
rect 4886 4798 5029 4799
rect 4886 4795 4997 4798
rect 4886 4768 4923 4795
rect 4952 4771 4997 4795
rect 5026 4771 5029 4798
rect 4952 4768 5029 4771
rect 4886 4766 5029 4768
rect 4826 4753 5029 4766
rect 4826 4752 4927 4753
rect 1810 4527 1868 4532
rect 1677 4515 1733 4522
rect 2302 4515 2307 4535
rect 2328 4515 2334 4535
rect 1677 4514 1712 4515
rect 2302 4508 2334 4515
rect 2725 4538 2781 4543
rect 2725 4518 2732 4538
rect 2752 4518 2781 4538
rect 2725 4511 2781 4518
rect 5204 4690 5236 4697
rect 5204 4670 5211 4690
rect 5232 4670 5236 4690
rect 5204 4605 5236 4670
rect 5416 4661 5447 4861
rect 5651 4860 5683 4861
rect 5648 4855 5683 4860
rect 5648 4835 5655 4855
rect 5675 4835 5683 4855
rect 5648 4827 5683 4835
rect 5416 4631 5422 4661
rect 5443 4631 5447 4661
rect 5416 4623 5447 4631
rect 5574 4605 5614 4606
rect 5204 4603 5616 4605
rect 5204 4577 5584 4603
rect 5610 4577 5616 4603
rect 5204 4569 5616 4577
rect 5204 4541 5236 4569
rect 5204 4521 5209 4541
rect 5230 4521 5236 4541
rect 5204 4514 5236 4521
rect 5406 4543 5454 4550
rect 5649 4549 5683 4827
rect 5406 4523 5413 4543
rect 5446 4523 5454 4543
rect 2725 4510 2760 4511
rect 968 4459 1079 4463
rect 2751 4459 4321 4460
rect 290 4455 4321 4459
rect 4646 4455 5064 4468
rect 290 4443 5064 4455
rect 290 4441 4926 4443
rect 290 4421 976 4441
rect 995 4421 1053 4441
rect 1072 4437 4926 4441
rect 1072 4421 2024 4437
rect 290 4417 2024 4421
rect 2043 4417 2101 4437
rect 2120 4423 4926 4437
rect 4945 4423 5003 4443
rect 5022 4423 5064 4443
rect 2120 4417 5064 4423
rect 290 4403 5064 4417
rect 290 3780 397 4403
rect 2016 4400 2127 4403
rect 4646 4397 5064 4403
rect 776 4354 840 4358
rect 772 4348 840 4354
rect 772 4315 789 4348
rect 829 4315 840 4348
rect 772 4303 840 4315
rect 1823 4317 1888 4339
rect 772 4301 829 4303
rect 776 3940 827 4301
rect 1823 4278 1840 4317
rect 1885 4278 1888 4317
rect 1464 4233 1499 4235
rect 1464 4224 1568 4233
rect 1464 4223 1515 4224
rect 1464 4203 1467 4223
rect 1492 4204 1515 4223
rect 1547 4204 1568 4224
rect 1492 4203 1568 4204
rect 1464 4196 1568 4203
rect 1464 4184 1499 4196
rect 876 4118 1079 4131
rect 876 4085 900 4118
rect 936 4117 1079 4118
rect 936 4114 1047 4117
rect 936 4087 973 4114
rect 1002 4090 1047 4114
rect 1076 4090 1079 4117
rect 1002 4087 1079 4090
rect 936 4085 1079 4087
rect 876 4072 1079 4085
rect 876 4071 977 4072
rect 1254 4009 1286 4016
rect 1254 3989 1261 4009
rect 1282 3989 1286 4009
rect 765 3931 830 3940
rect 765 3894 775 3931
rect 815 3897 830 3931
rect 1254 3924 1286 3989
rect 1466 3980 1497 4184
rect 1701 4179 1733 4180
rect 1698 4174 1733 4179
rect 1698 4154 1705 4174
rect 1725 4154 1733 4174
rect 1698 4146 1733 4154
rect 1466 3950 1472 3980
rect 1493 3950 1497 3980
rect 1466 3942 1497 3950
rect 1624 3924 1664 3925
rect 1254 3922 1666 3924
rect 815 3894 832 3897
rect 765 3875 832 3894
rect 765 3854 779 3875
rect 815 3854 832 3875
rect 765 3847 832 3854
rect 1254 3896 1634 3922
rect 1660 3896 1666 3922
rect 1254 3888 1666 3896
rect 1254 3860 1286 3888
rect 1699 3868 1733 4146
rect 1823 3978 1888 4278
rect 3960 4239 3997 4260
rect 3960 4202 3971 4239
rect 3988 4215 3997 4239
rect 3988 4202 3998 4215
rect 3960 4192 3998 4202
rect 3961 4188 3998 4192
rect 3961 4182 3994 4188
rect 3371 4113 3574 4126
rect 3371 4080 3395 4113
rect 3431 4112 3574 4113
rect 3431 4109 3542 4112
rect 3431 4082 3468 4109
rect 3497 4085 3542 4109
rect 3571 4085 3574 4112
rect 3497 4082 3574 4085
rect 3431 4080 3574 4082
rect 3371 4067 3574 4080
rect 3371 4066 3472 4067
rect 3749 4004 3781 4011
rect 3749 3984 3756 4004
rect 3777 3984 3781 4004
rect 1254 3840 1259 3860
rect 1280 3840 1286 3860
rect 1254 3833 1286 3840
rect 1677 3863 1733 3868
rect 1677 3843 1684 3863
rect 1704 3843 1733 3863
rect 1677 3836 1733 3843
rect 1813 3967 1893 3978
rect 1813 3941 1830 3967
rect 1870 3941 1893 3967
rect 1813 3914 1893 3941
rect 1813 3888 1834 3914
rect 1874 3888 1893 3914
rect 1813 3869 1893 3888
rect 1813 3843 1837 3869
rect 1877 3843 1893 3869
rect 2887 3913 2992 3934
rect 3749 3919 3781 3984
rect 3961 3975 3992 4182
rect 4196 4174 4228 4175
rect 4193 4169 4228 4174
rect 4193 4149 4200 4169
rect 4220 4149 4228 4169
rect 4193 4141 4228 4149
rect 3961 3945 3967 3975
rect 3988 3945 3992 3975
rect 3961 3937 3992 3945
rect 4119 3919 4159 3920
rect 3749 3917 4161 3919
rect 2887 3907 3363 3913
rect 2887 3905 2944 3907
rect 2887 3874 2899 3905
rect 2924 3884 2944 3905
rect 2970 3900 3363 3907
rect 2970 3884 3324 3900
rect 2924 3877 3324 3884
rect 3350 3877 3363 3900
rect 2924 3874 3363 3877
rect 2887 3864 3363 3874
rect 3749 3891 4129 3917
rect 4155 3891 4161 3917
rect 3749 3883 4161 3891
rect 2887 3862 2992 3864
rect 1677 3835 1712 3836
rect 1813 3831 1893 3843
rect 3749 3855 3781 3883
rect 4194 3863 4228 4141
rect 3749 3835 3754 3855
rect 3775 3835 3781 3855
rect 3749 3828 3781 3835
rect 4172 3858 4228 3863
rect 4172 3838 4179 3858
rect 4199 3838 4228 3858
rect 4172 3831 4228 3838
rect 4172 3830 4207 3831
rect 968 3780 1079 3784
rect 2710 3780 4363 3783
rect 288 3762 4363 3780
rect 288 3742 976 3762
rect 995 3742 1053 3762
rect 1072 3757 4363 3762
rect 1072 3742 3471 3757
rect 288 3737 3471 3742
rect 3490 3737 3548 3757
rect 3567 3737 4363 3757
rect 288 3727 4363 3737
rect 288 3724 913 3727
rect 1100 3724 4363 3727
rect 290 3496 397 3724
rect 2710 3723 4363 3724
rect 3463 3720 3574 3723
rect 758 3685 879 3695
rect 758 3683 827 3685
rect 758 3642 771 3683
rect 808 3644 827 3683
rect 864 3644 879 3685
rect 808 3642 879 3644
rect 758 3624 879 3642
rect 764 3522 843 3624
rect 1816 3584 1883 3603
rect 1816 3564 1836 3584
rect 290 3441 398 3496
rect 765 3441 843 3522
rect 1815 3518 1836 3564
rect 1866 3564 1883 3584
rect 1866 3534 1885 3564
rect 1866 3518 1886 3534
rect 1815 3502 1886 3518
rect 1465 3491 1537 3492
rect 1464 3483 1563 3491
rect 1464 3480 1516 3483
rect 1464 3445 1472 3480
rect 1497 3445 1516 3480
rect 1541 3445 1563 3483
rect 290 3012 397 3441
rect 769 3200 841 3441
rect 1464 3433 1563 3445
rect 1465 3414 1533 3433
rect 1466 3411 1499 3414
rect 1701 3411 1733 3412
rect 876 3350 1079 3363
rect 876 3317 900 3350
rect 936 3349 1079 3350
rect 936 3346 1047 3349
rect 936 3319 973 3346
rect 1002 3322 1047 3346
rect 1076 3322 1079 3349
rect 1002 3319 1079 3322
rect 936 3317 1079 3319
rect 876 3304 1079 3317
rect 876 3303 977 3304
rect 769 3158 778 3200
rect 827 3158 841 3200
rect 769 3137 841 3158
rect 769 3095 779 3137
rect 828 3095 841 3137
rect 769 3077 841 3095
rect 1254 3241 1286 3248
rect 1254 3221 1261 3241
rect 1282 3221 1286 3241
rect 1254 3156 1286 3221
rect 1466 3212 1497 3411
rect 1698 3406 1733 3411
rect 1698 3386 1705 3406
rect 1725 3386 1733 3406
rect 1698 3378 1733 3386
rect 1466 3182 1472 3212
rect 1493 3182 1497 3212
rect 1466 3174 1497 3182
rect 1624 3156 1664 3157
rect 1254 3154 1666 3156
rect 1254 3128 1634 3154
rect 1660 3128 1666 3154
rect 1254 3120 1666 3128
rect 1254 3092 1286 3120
rect 1699 3100 1733 3378
rect 1815 3191 1885 3502
rect 2512 3493 3854 3498
rect 2512 3491 3811 3493
rect 2509 3465 3811 3491
rect 3839 3465 3854 3493
rect 2509 3457 3854 3465
rect 2509 3432 2548 3457
rect 2509 3415 2550 3432
rect 2509 3408 2548 3415
rect 1924 3346 2127 3359
rect 1924 3313 1948 3346
rect 1984 3345 2127 3346
rect 1984 3342 2095 3345
rect 1984 3315 2021 3342
rect 2050 3318 2095 3342
rect 2124 3318 2127 3345
rect 2050 3315 2127 3318
rect 1984 3313 2127 3315
rect 1924 3300 2127 3313
rect 1924 3299 2025 3300
rect 1254 3072 1259 3092
rect 1280 3072 1286 3092
rect 1254 3065 1286 3072
rect 1677 3095 1733 3100
rect 1677 3075 1684 3095
rect 1704 3075 1733 3095
rect 1810 3185 1885 3191
rect 1810 3152 1818 3185
rect 1871 3152 1885 3185
rect 1810 3127 1885 3152
rect 1810 3094 1823 3127
rect 1876 3094 1885 3127
rect 1810 3085 1885 3094
rect 2302 3237 2334 3244
rect 2302 3217 2309 3237
rect 2330 3217 2334 3237
rect 2302 3152 2334 3217
rect 2514 3208 2545 3408
rect 2749 3407 2781 3408
rect 2746 3402 2781 3407
rect 2746 3382 2753 3402
rect 2773 3382 2781 3402
rect 2746 3374 2781 3382
rect 2514 3178 2520 3208
rect 2541 3178 2545 3208
rect 2514 3170 2545 3178
rect 2672 3152 2712 3153
rect 2302 3150 2714 3152
rect 2302 3124 2682 3150
rect 2708 3124 2714 3150
rect 2302 3116 2714 3124
rect 2302 3088 2334 3116
rect 2747 3096 2781 3374
rect 1810 3080 1868 3085
rect 1677 3068 1733 3075
rect 2302 3068 2307 3088
rect 2328 3068 2334 3088
rect 1677 3067 1712 3068
rect 2302 3061 2334 3068
rect 2725 3091 2781 3096
rect 2725 3071 2732 3091
rect 2752 3071 2781 3091
rect 2725 3064 2781 3071
rect 2725 3063 2760 3064
rect 968 3012 1079 3016
rect 2843 3012 4363 3013
rect 290 2994 4363 3012
rect 290 2974 976 2994
rect 995 2974 1053 2994
rect 1072 2990 4363 2994
rect 1072 2974 2024 2990
rect 290 2970 2024 2974
rect 2043 2970 2101 2990
rect 2120 2970 4363 2990
rect 290 2956 4363 2970
rect 290 2333 397 2956
rect 2016 2953 2127 2956
rect 776 2907 840 2911
rect 772 2901 840 2907
rect 772 2868 789 2901
rect 829 2868 840 2901
rect 772 2856 840 2868
rect 1823 2870 1888 2892
rect 772 2854 829 2856
rect 776 2493 827 2854
rect 1823 2831 1840 2870
rect 1885 2831 1888 2870
rect 1464 2786 1499 2788
rect 1464 2777 1568 2786
rect 1464 2776 1515 2777
rect 1464 2756 1467 2776
rect 1492 2757 1515 2776
rect 1547 2757 1568 2777
rect 1492 2756 1568 2757
rect 1464 2749 1568 2756
rect 1464 2737 1499 2749
rect 876 2671 1079 2684
rect 876 2638 900 2671
rect 936 2670 1079 2671
rect 936 2667 1047 2670
rect 936 2640 973 2667
rect 1002 2643 1047 2667
rect 1076 2643 1079 2670
rect 1002 2640 1079 2643
rect 936 2638 1079 2640
rect 876 2625 1079 2638
rect 876 2624 977 2625
rect 1254 2562 1286 2569
rect 1254 2542 1261 2562
rect 1282 2542 1286 2562
rect 765 2484 830 2493
rect 765 2447 775 2484
rect 815 2450 830 2484
rect 1254 2477 1286 2542
rect 1466 2533 1497 2737
rect 1701 2732 1733 2733
rect 1698 2727 1733 2732
rect 1698 2707 1705 2727
rect 1725 2707 1733 2727
rect 1698 2699 1733 2707
rect 1466 2503 1472 2533
rect 1493 2503 1497 2533
rect 1466 2495 1497 2503
rect 1624 2477 1664 2478
rect 1254 2475 1666 2477
rect 815 2447 832 2450
rect 765 2428 832 2447
rect 765 2407 779 2428
rect 815 2407 832 2428
rect 765 2400 832 2407
rect 1254 2449 1634 2475
rect 1660 2449 1666 2475
rect 1254 2441 1666 2449
rect 1254 2413 1286 2441
rect 1699 2421 1733 2699
rect 1823 2568 1888 2831
rect 1823 2564 1884 2568
rect 1254 2393 1259 2413
rect 1280 2393 1286 2413
rect 1254 2386 1286 2393
rect 1677 2416 1733 2421
rect 1677 2396 1684 2416
rect 1704 2396 1733 2416
rect 1677 2389 1733 2396
rect 1677 2388 1712 2389
rect 968 2333 1079 2337
rect 288 2315 1607 2333
rect 288 2295 976 2315
rect 995 2295 1053 2315
rect 1072 2295 1607 2315
rect 288 2277 1607 2295
rect 290 2157 397 2277
rect 758 2238 879 2248
rect 758 2236 827 2238
rect 758 2195 771 2236
rect 808 2197 827 2236
rect 864 2197 879 2238
rect 808 2195 879 2197
rect 758 2177 879 2195
rect 89 2084 223 2113
rect 89 1972 127 2084
rect 206 1972 223 2084
rect 290 2077 398 2157
rect 89 1019 223 1972
rect 291 1265 398 2077
rect 764 2105 829 2177
rect 764 2039 832 2105
rect 765 1493 832 2039
rect 1819 1677 1884 2564
rect 2862 2294 2999 2298
rect 2849 2290 3006 2294
rect 2849 2183 2886 2290
rect 2986 2183 3006 2290
rect 2849 2141 3006 2183
rect 2862 1893 2999 2141
rect 2852 1851 3018 1893
rect 2852 1776 2881 1851
rect 2998 1776 3018 1851
rect 2852 1760 3018 1776
rect 1808 1656 1945 1677
rect 1808 1581 1833 1656
rect 1903 1581 1945 1656
rect 1808 1550 1945 1581
rect 751 1444 926 1493
rect 751 1365 784 1444
rect 884 1365 926 1444
rect 751 1360 926 1365
rect 291 1223 439 1265
rect 291 1215 331 1223
rect 293 1136 331 1215
rect 401 1136 439 1223
rect 293 1098 439 1136
rect 85 983 224 1019
rect 85 888 99 983
rect 189 888 224 983
rect 85 870 224 888
rect 5406 793 5454 4523
rect 5627 4544 5683 4549
rect 5627 4524 5634 4544
rect 5654 4524 5683 4544
rect 5627 4517 5683 4524
rect 5627 4516 5662 4517
rect 5731 4426 5759 7234
rect 8944 7189 9009 7489
rect 9099 7321 9133 7599
rect 9546 7579 9578 7607
rect 9166 7571 9578 7579
rect 9166 7545 9172 7571
rect 9198 7545 9578 7571
rect 10000 7613 10067 7620
rect 10000 7592 10017 7613
rect 10053 7592 10067 7613
rect 10000 7573 10067 7592
rect 10000 7570 10017 7573
rect 9166 7543 9578 7545
rect 9168 7542 9208 7543
rect 9335 7517 9366 7525
rect 9335 7487 9339 7517
rect 9360 7487 9366 7517
rect 9099 7313 9134 7321
rect 9099 7293 9107 7313
rect 9127 7293 9134 7313
rect 9099 7288 9134 7293
rect 9099 7287 9131 7288
rect 9335 7283 9366 7487
rect 9546 7478 9578 7543
rect 10002 7536 10017 7570
rect 10057 7536 10067 7573
rect 10002 7527 10067 7536
rect 9546 7458 9550 7478
rect 9571 7458 9578 7478
rect 9546 7451 9578 7458
rect 9855 7395 9956 7396
rect 9753 7382 9956 7395
rect 9753 7380 9896 7382
rect 9753 7377 9830 7380
rect 9753 7350 9756 7377
rect 9785 7353 9830 7377
rect 9859 7353 9896 7380
rect 9785 7350 9896 7353
rect 9753 7349 9896 7350
rect 9932 7349 9956 7382
rect 9753 7336 9956 7349
rect 9333 7271 9368 7283
rect 9264 7264 9368 7271
rect 9264 7263 9340 7264
rect 9264 7243 9285 7263
rect 9317 7244 9340 7263
rect 9365 7244 9368 7264
rect 9317 7243 9368 7244
rect 9264 7234 9368 7243
rect 9333 7232 9368 7234
rect 8944 7150 8947 7189
rect 8992 7150 9009 7189
rect 10005 7166 10056 7527
rect 10003 7164 10060 7166
rect 8944 7128 9009 7150
rect 9992 7152 10060 7164
rect 9992 7119 10003 7152
rect 10043 7119 10060 7152
rect 9992 7113 10060 7119
rect 9992 7109 10056 7113
rect 8705 7064 8816 7067
rect 10435 7064 10542 7687
rect 6999 7050 10542 7064
rect 6999 7030 8712 7050
rect 8731 7030 8789 7050
rect 8808 7046 10542 7050
rect 8808 7030 9760 7046
rect 6999 7026 9760 7030
rect 9779 7026 9837 7046
rect 9856 7026 10542 7046
rect 6999 7008 10542 7026
rect 6999 7007 7989 7008
rect 9753 7004 9864 7008
rect 8072 6956 8107 6957
rect 8051 6949 8107 6956
rect 8051 6929 8080 6949
rect 8100 6929 8107 6949
rect 8051 6924 8107 6929
rect 8498 6952 8530 6959
rect 9120 6952 9155 6953
rect 8498 6932 8504 6952
rect 8525 6932 8530 6952
rect 9099 6945 9155 6952
rect 8964 6935 9022 6940
rect 8051 6646 8085 6924
rect 8498 6904 8530 6932
rect 8118 6896 8530 6904
rect 8118 6870 8124 6896
rect 8150 6870 8530 6896
rect 8118 6868 8530 6870
rect 8120 6867 8160 6868
rect 8287 6842 8318 6850
rect 8287 6812 8291 6842
rect 8312 6812 8318 6842
rect 8051 6638 8086 6646
rect 8051 6618 8059 6638
rect 8079 6618 8086 6638
rect 8051 6613 8086 6618
rect 8051 6612 8083 6613
rect 8287 6612 8318 6812
rect 8498 6803 8530 6868
rect 8498 6783 8502 6803
rect 8523 6783 8530 6803
rect 8498 6776 8530 6783
rect 8947 6926 9022 6935
rect 8947 6893 8956 6926
rect 9009 6893 9022 6926
rect 8947 6868 9022 6893
rect 8947 6835 8961 6868
rect 9014 6835 9022 6868
rect 8947 6829 9022 6835
rect 9099 6925 9128 6945
rect 9148 6925 9155 6945
rect 9099 6920 9155 6925
rect 9546 6948 9578 6955
rect 9546 6928 9552 6948
rect 9573 6928 9578 6948
rect 8807 6720 8908 6721
rect 8705 6707 8908 6720
rect 8705 6705 8848 6707
rect 8705 6702 8782 6705
rect 8705 6675 8708 6702
rect 8737 6678 8782 6702
rect 8811 6678 8848 6705
rect 8737 6675 8848 6678
rect 8705 6674 8848 6675
rect 8884 6674 8908 6707
rect 8705 6661 8908 6674
rect 8284 6605 8323 6612
rect 8282 6588 8323 6605
rect 8284 6563 8323 6588
rect 6978 6555 8323 6563
rect 6978 6527 6993 6555
rect 7021 6529 8323 6555
rect 7021 6527 8320 6529
rect 6978 6522 8320 6527
rect 8947 6518 9017 6829
rect 9099 6642 9133 6920
rect 9546 6900 9578 6928
rect 9166 6892 9578 6900
rect 9166 6866 9172 6892
rect 9198 6866 9578 6892
rect 9166 6864 9578 6866
rect 9168 6863 9208 6864
rect 9335 6838 9366 6846
rect 9335 6808 9339 6838
rect 9360 6808 9366 6838
rect 9099 6634 9134 6642
rect 9099 6614 9107 6634
rect 9127 6614 9134 6634
rect 9099 6609 9134 6614
rect 9335 6609 9366 6808
rect 9546 6799 9578 6864
rect 9546 6779 9550 6799
rect 9571 6779 9578 6799
rect 9546 6772 9578 6779
rect 9991 6925 10063 6943
rect 9991 6883 10004 6925
rect 10053 6883 10063 6925
rect 9991 6862 10063 6883
rect 9991 6820 10005 6862
rect 10054 6820 10063 6862
rect 9855 6716 9956 6717
rect 9753 6703 9956 6716
rect 9753 6701 9896 6703
rect 9753 6698 9830 6701
rect 9753 6671 9756 6698
rect 9785 6674 9830 6698
rect 9859 6674 9896 6701
rect 9785 6671 9896 6674
rect 9753 6670 9896 6671
rect 9932 6670 9956 6703
rect 9753 6657 9956 6670
rect 9099 6608 9131 6609
rect 9333 6606 9366 6609
rect 9299 6587 9367 6606
rect 9269 6575 9368 6587
rect 9991 6579 10063 6820
rect 10435 6579 10542 7008
rect 10997 7420 11104 7880
rect 11476 7608 11548 7902
rect 12172 7899 12244 7900
rect 12171 7891 12270 7899
rect 12524 7894 12601 8077
rect 13812 8078 13896 8089
rect 13812 8050 13840 8078
rect 13884 8050 13896 8078
rect 13626 7999 13700 8027
rect 13626 7951 13649 7999
rect 13686 7951 13700 7999
rect 13812 8021 13896 8050
rect 13812 7993 13837 8021
rect 13881 7993 13896 8021
rect 13812 7960 13896 7993
rect 13626 7942 13700 7951
rect 13222 7900 13294 7901
rect 12171 7888 12223 7891
rect 12171 7853 12179 7888
rect 12204 7853 12223 7888
rect 12248 7853 12270 7891
rect 12171 7841 12270 7853
rect 12522 7865 12601 7894
rect 13221 7892 13310 7900
rect 13221 7889 13273 7892
rect 12172 7822 12240 7841
rect 12173 7819 12206 7822
rect 12408 7819 12440 7820
rect 11583 7758 11786 7771
rect 11583 7725 11607 7758
rect 11643 7757 11786 7758
rect 11643 7754 11754 7757
rect 11643 7727 11680 7754
rect 11709 7730 11754 7754
rect 11783 7730 11786 7757
rect 11709 7727 11786 7730
rect 11643 7725 11786 7727
rect 11583 7712 11786 7725
rect 11583 7711 11684 7712
rect 11476 7566 11485 7608
rect 11534 7566 11548 7608
rect 11476 7545 11548 7566
rect 11476 7503 11486 7545
rect 11535 7503 11548 7545
rect 11476 7485 11548 7503
rect 11961 7649 11993 7656
rect 11961 7629 11968 7649
rect 11989 7629 11993 7649
rect 11961 7564 11993 7629
rect 12173 7620 12204 7819
rect 12405 7814 12440 7819
rect 12405 7794 12412 7814
rect 12432 7794 12440 7814
rect 12405 7786 12440 7794
rect 12173 7590 12179 7620
rect 12200 7590 12204 7620
rect 12173 7582 12204 7590
rect 12331 7564 12371 7565
rect 11961 7562 12373 7564
rect 11961 7536 12341 7562
rect 12367 7536 12373 7562
rect 11961 7528 12373 7536
rect 11961 7500 11993 7528
rect 12406 7508 12440 7786
rect 12522 7599 12592 7865
rect 13221 7854 13229 7889
rect 13254 7854 13273 7889
rect 13298 7854 13310 7892
rect 13221 7842 13310 7854
rect 13221 7841 13290 7842
rect 13221 7823 13257 7841
rect 12631 7754 12834 7767
rect 12631 7721 12655 7754
rect 12691 7753 12834 7754
rect 12691 7750 12802 7753
rect 12691 7723 12728 7750
rect 12757 7726 12802 7750
rect 12831 7726 12834 7753
rect 12757 7723 12834 7726
rect 12691 7721 12834 7723
rect 12631 7708 12834 7721
rect 12631 7707 12732 7708
rect 11961 7480 11966 7500
rect 11987 7480 11993 7500
rect 11961 7473 11993 7480
rect 12384 7503 12440 7508
rect 12384 7483 12391 7503
rect 12411 7483 12440 7503
rect 12517 7593 12592 7599
rect 12517 7560 12525 7593
rect 12578 7560 12592 7593
rect 12517 7535 12592 7560
rect 12517 7502 12530 7535
rect 12583 7502 12592 7535
rect 12517 7493 12592 7502
rect 13009 7645 13041 7652
rect 13009 7625 13016 7645
rect 13037 7625 13041 7645
rect 13009 7560 13041 7625
rect 13221 7616 13252 7823
rect 13456 7815 13488 7816
rect 13453 7810 13488 7815
rect 13453 7790 13460 7810
rect 13480 7790 13488 7810
rect 13453 7782 13488 7790
rect 13221 7586 13227 7616
rect 13248 7586 13252 7616
rect 13221 7578 13252 7586
rect 13379 7560 13419 7561
rect 13009 7558 13421 7560
rect 13009 7532 13389 7558
rect 13415 7532 13421 7558
rect 13009 7524 13421 7532
rect 13009 7496 13041 7524
rect 13454 7504 13488 7782
rect 13637 7597 13699 7942
rect 13806 7915 13896 7960
rect 13806 7600 13888 7915
rect 13637 7578 13701 7597
rect 13637 7539 13650 7578
rect 13684 7539 13701 7578
rect 13637 7520 13701 7539
rect 13806 7559 13827 7600
rect 13863 7559 13888 7600
rect 13806 7530 13888 7559
rect 12517 7488 12575 7493
rect 12384 7476 12440 7483
rect 13009 7476 13014 7496
rect 13035 7476 13041 7496
rect 12384 7475 12419 7476
rect 13009 7469 13041 7476
rect 13432 7499 13488 7504
rect 13432 7479 13439 7499
rect 13459 7479 13488 7499
rect 13432 7472 13488 7479
rect 13432 7471 13467 7472
rect 11675 7420 11786 7424
rect 13458 7420 15028 7421
rect 10997 7402 15028 7420
rect 10997 7382 11683 7402
rect 11702 7382 11760 7402
rect 11779 7398 15028 7402
rect 11779 7382 12731 7398
rect 10997 7378 12731 7382
rect 12750 7378 12808 7398
rect 12827 7378 15028 7398
rect 10997 7364 15028 7378
rect 10997 6741 11104 7364
rect 12723 7361 12834 7364
rect 11483 7315 11547 7319
rect 11479 7309 11547 7315
rect 11479 7276 11496 7309
rect 11536 7276 11547 7309
rect 11479 7264 11547 7276
rect 12530 7278 12595 7300
rect 11479 7262 11536 7264
rect 11483 6901 11534 7262
rect 12530 7239 12547 7278
rect 12592 7239 12595 7278
rect 12171 7194 12206 7196
rect 12171 7185 12275 7194
rect 12171 7184 12222 7185
rect 12171 7164 12174 7184
rect 12199 7165 12222 7184
rect 12254 7165 12275 7185
rect 12199 7164 12275 7165
rect 12171 7157 12275 7164
rect 12171 7145 12206 7157
rect 11583 7079 11786 7092
rect 11583 7046 11607 7079
rect 11643 7078 11786 7079
rect 11643 7075 11754 7078
rect 11643 7048 11680 7075
rect 11709 7051 11754 7075
rect 11783 7051 11786 7078
rect 11709 7048 11786 7051
rect 11643 7046 11786 7048
rect 11583 7033 11786 7046
rect 11583 7032 11684 7033
rect 11961 6970 11993 6977
rect 11961 6950 11968 6970
rect 11989 6950 11993 6970
rect 11472 6892 11537 6901
rect 11472 6855 11482 6892
rect 11522 6858 11537 6892
rect 11961 6885 11993 6950
rect 12173 6941 12204 7145
rect 12408 7140 12440 7141
rect 12405 7135 12440 7140
rect 12405 7115 12412 7135
rect 12432 7115 12440 7135
rect 12405 7107 12440 7115
rect 12173 6911 12179 6941
rect 12200 6911 12204 6941
rect 12173 6903 12204 6911
rect 12331 6885 12371 6886
rect 11961 6883 12373 6885
rect 11522 6855 11539 6858
rect 11472 6836 11539 6855
rect 11472 6815 11486 6836
rect 11522 6815 11539 6836
rect 11472 6808 11539 6815
rect 11961 6857 12341 6883
rect 12367 6857 12373 6883
rect 11961 6849 12373 6857
rect 11961 6821 11993 6849
rect 12406 6829 12440 7107
rect 12530 6939 12595 7239
rect 13801 7263 13894 7278
rect 13801 7219 13816 7263
rect 13876 7219 13894 7263
rect 11961 6801 11966 6821
rect 11987 6801 11993 6821
rect 11961 6794 11993 6801
rect 12384 6824 12440 6829
rect 12384 6804 12391 6824
rect 12411 6804 12440 6824
rect 12384 6797 12440 6804
rect 12520 6928 12600 6939
rect 12520 6902 12537 6928
rect 12577 6902 12600 6928
rect 12520 6875 12600 6902
rect 12520 6849 12541 6875
rect 12581 6849 12600 6875
rect 12520 6830 12600 6849
rect 12520 6804 12544 6830
rect 12584 6804 12600 6830
rect 12384 6796 12419 6797
rect 12520 6792 12600 6804
rect 13801 6846 13894 7219
rect 14078 7074 14281 7087
rect 14078 7041 14102 7074
rect 14138 7073 14281 7074
rect 14138 7070 14249 7073
rect 14138 7043 14175 7070
rect 14204 7046 14249 7070
rect 14278 7046 14281 7073
rect 14204 7043 14281 7046
rect 14138 7041 14281 7043
rect 14078 7028 14281 7041
rect 14078 7027 14179 7028
rect 13801 6805 13816 6846
rect 13870 6805 13894 6846
rect 13801 6798 13894 6805
rect 14456 6965 14488 6972
rect 14456 6945 14463 6965
rect 14484 6945 14488 6965
rect 14456 6880 14488 6945
rect 14668 6936 14699 7137
rect 14903 7135 14935 7136
rect 14900 7130 14935 7135
rect 14900 7110 14907 7130
rect 14927 7110 14935 7130
rect 14900 7102 14935 7110
rect 14668 6906 14674 6936
rect 14695 6906 14699 6936
rect 14668 6898 14699 6906
rect 14826 6880 14866 6881
rect 14456 6878 14868 6880
rect 14456 6852 14836 6878
rect 14862 6852 14868 6878
rect 14456 6844 14868 6852
rect 14456 6816 14488 6844
rect 14901 6824 14935 7102
rect 14456 6796 14461 6816
rect 14482 6796 14488 6816
rect 14456 6789 14488 6796
rect 14879 6819 14935 6824
rect 14879 6799 14886 6819
rect 14906 6799 14935 6819
rect 14879 6792 14935 6799
rect 14879 6791 14914 6792
rect 11675 6741 11786 6745
rect 13417 6741 15061 6744
rect 10995 6723 15061 6741
rect 10995 6703 11683 6723
rect 11702 6703 11760 6723
rect 11779 6718 15061 6723
rect 11779 6703 14178 6718
rect 10995 6698 14178 6703
rect 14197 6698 14255 6718
rect 14274 6698 15061 6718
rect 10995 6688 15061 6698
rect 10995 6685 11620 6688
rect 11807 6685 15061 6688
rect 9269 6537 9291 6575
rect 9316 6540 9335 6575
rect 9360 6540 9368 6575
rect 9316 6537 9368 6540
rect 9269 6529 9368 6537
rect 9295 6528 9367 6529
rect 8946 6502 9017 6518
rect 8946 6486 8966 6502
rect 8947 6456 8966 6486
rect 8949 6436 8966 6456
rect 8996 6456 9017 6502
rect 9989 6498 10067 6579
rect 10434 6524 10542 6579
rect 8996 6436 9016 6456
rect 8949 6417 9016 6436
rect 9989 6396 10068 6498
rect 9953 6378 10074 6396
rect 9953 6376 10024 6378
rect 9953 6335 9968 6376
rect 10005 6337 10024 6376
rect 10061 6337 10074 6378
rect 10005 6335 10074 6337
rect 9953 6325 10074 6335
rect 7258 6297 7369 6300
rect 6572 6296 8122 6297
rect 10435 6296 10542 6524
rect 10997 6457 11104 6685
rect 13417 6684 15061 6685
rect 14170 6681 14281 6684
rect 11465 6646 11586 6656
rect 11465 6644 11534 6646
rect 11465 6603 11478 6644
rect 11515 6605 11534 6644
rect 11571 6605 11586 6646
rect 11515 6603 11586 6605
rect 11465 6585 11586 6603
rect 14670 6626 14756 6630
rect 14670 6608 14685 6626
rect 14737 6608 14756 6626
rect 14670 6599 14756 6608
rect 11471 6483 11550 6585
rect 12523 6545 12590 6564
rect 12523 6525 12543 6545
rect 10997 6402 11105 6457
rect 11472 6402 11550 6483
rect 12522 6479 12543 6525
rect 12573 6525 12590 6545
rect 12573 6495 12592 6525
rect 12573 6479 12593 6495
rect 12522 6463 12593 6479
rect 12172 6452 12244 6453
rect 12171 6444 12270 6452
rect 12171 6441 12223 6444
rect 12171 6406 12179 6441
rect 12204 6406 12223 6441
rect 12248 6406 12270 6444
rect 6572 6293 9732 6296
rect 9919 6293 10544 6296
rect 6572 6283 10544 6293
rect 6572 6263 7265 6283
rect 7284 6263 7342 6283
rect 7361 6278 10544 6283
rect 7361 6263 9760 6278
rect 6572 6258 9760 6263
rect 9779 6258 9837 6278
rect 9856 6258 10544 6278
rect 6572 6240 10544 6258
rect 6572 6237 8122 6240
rect 9753 6236 9864 6240
rect 6625 6189 6660 6190
rect 6604 6182 6660 6189
rect 6604 6162 6633 6182
rect 6653 6162 6660 6182
rect 6604 6157 6660 6162
rect 7051 6185 7083 6192
rect 7051 6165 7057 6185
rect 7078 6165 7083 6185
rect 6604 5879 6638 6157
rect 7051 6137 7083 6165
rect 8939 6177 9019 6189
rect 9120 6184 9155 6185
rect 6671 6129 7083 6137
rect 6671 6103 6677 6129
rect 6703 6103 7083 6129
rect 7469 6143 7906 6156
rect 7469 6120 7482 6143
rect 7508 6136 7906 6143
rect 7508 6120 7862 6136
rect 7469 6113 7862 6120
rect 7888 6113 7906 6136
rect 7469 6107 7906 6113
rect 8939 6151 8955 6177
rect 8995 6151 9019 6177
rect 8939 6132 9019 6151
rect 6671 6101 7083 6103
rect 6673 6100 6713 6101
rect 6840 6075 6871 6083
rect 6840 6045 6844 6075
rect 6865 6045 6871 6075
rect 6604 5871 6639 5879
rect 6604 5851 6612 5871
rect 6632 5851 6639 5871
rect 6604 5846 6639 5851
rect 6604 5845 6636 5846
rect 6840 5838 6871 6045
rect 7051 6036 7083 6101
rect 8939 6106 8958 6132
rect 8998 6106 9019 6132
rect 8939 6079 9019 6106
rect 8939 6053 8962 6079
rect 9002 6053 9019 6079
rect 8939 6042 9019 6053
rect 9099 6177 9155 6184
rect 9099 6157 9128 6177
rect 9148 6157 9155 6177
rect 9099 6152 9155 6157
rect 9546 6180 9578 6187
rect 9546 6160 9552 6180
rect 9573 6160 9578 6180
rect 7051 6016 7055 6036
rect 7076 6016 7083 6036
rect 7051 6009 7083 6016
rect 7360 5953 7461 5954
rect 7258 5940 7461 5953
rect 7258 5938 7401 5940
rect 7258 5935 7335 5938
rect 7258 5908 7261 5935
rect 7290 5911 7335 5935
rect 7364 5911 7401 5938
rect 7290 5908 7401 5911
rect 7258 5907 7401 5908
rect 7437 5907 7461 5940
rect 7258 5894 7461 5907
rect 6838 5832 6871 5838
rect 6834 5828 6871 5832
rect 6834 5818 6872 5828
rect 6834 5805 6844 5818
rect 6835 5781 6844 5805
rect 6861 5781 6872 5818
rect 6835 5760 6872 5781
rect 8944 5742 9009 6042
rect 9099 5874 9133 6152
rect 9546 6132 9578 6160
rect 9166 6124 9578 6132
rect 9166 6098 9172 6124
rect 9198 6098 9578 6124
rect 10000 6166 10067 6173
rect 10000 6145 10017 6166
rect 10053 6145 10067 6166
rect 10000 6126 10067 6145
rect 10000 6123 10017 6126
rect 9166 6096 9578 6098
rect 9168 6095 9208 6096
rect 9335 6070 9366 6078
rect 9335 6040 9339 6070
rect 9360 6040 9366 6070
rect 9099 5866 9134 5874
rect 9099 5846 9107 5866
rect 9127 5846 9134 5866
rect 9099 5841 9134 5846
rect 9099 5840 9131 5841
rect 9335 5836 9366 6040
rect 9546 6031 9578 6096
rect 10002 6089 10017 6123
rect 10057 6089 10067 6126
rect 10002 6080 10067 6089
rect 9546 6011 9550 6031
rect 9571 6011 9578 6031
rect 9546 6004 9578 6011
rect 9855 5948 9956 5949
rect 9753 5935 9956 5948
rect 9753 5933 9896 5935
rect 9753 5930 9830 5933
rect 9753 5903 9756 5930
rect 9785 5906 9830 5930
rect 9859 5906 9896 5933
rect 9785 5903 9896 5906
rect 9753 5902 9896 5903
rect 9932 5902 9956 5935
rect 9753 5889 9956 5902
rect 9333 5824 9368 5836
rect 9264 5817 9368 5824
rect 9264 5816 9340 5817
rect 9264 5796 9285 5816
rect 9317 5797 9340 5816
rect 9365 5797 9368 5817
rect 9317 5796 9368 5797
rect 9264 5787 9368 5796
rect 9333 5785 9368 5787
rect 8944 5703 8947 5742
rect 8992 5703 9009 5742
rect 10005 5719 10056 6080
rect 10003 5717 10060 5719
rect 8944 5681 9009 5703
rect 9992 5705 10060 5717
rect 9992 5672 10003 5705
rect 10043 5672 10060 5705
rect 9992 5666 10060 5672
rect 9992 5662 10056 5666
rect 8705 5617 8816 5620
rect 10435 5617 10542 6240
rect 6781 5603 10542 5617
rect 6781 5583 8712 5603
rect 8731 5583 8789 5603
rect 8808 5599 10542 5603
rect 8808 5583 9760 5599
rect 6781 5579 9760 5583
rect 9779 5579 9837 5599
rect 9856 5579 10542 5599
rect 6781 5561 10542 5579
rect 6781 5560 8081 5561
rect 9753 5557 9864 5561
rect 8072 5509 8107 5510
rect 8051 5502 8107 5509
rect 8051 5482 8080 5502
rect 8100 5482 8107 5502
rect 8051 5477 8107 5482
rect 8498 5505 8530 5512
rect 9120 5505 9155 5506
rect 8498 5485 8504 5505
rect 8525 5485 8530 5505
rect 9099 5498 9155 5505
rect 8964 5488 9022 5493
rect 8051 5199 8085 5477
rect 8498 5457 8530 5485
rect 8118 5449 8530 5457
rect 8118 5423 8124 5449
rect 8150 5423 8530 5449
rect 8118 5421 8530 5423
rect 8120 5420 8160 5421
rect 8287 5395 8318 5403
rect 8287 5365 8291 5395
rect 8312 5365 8318 5395
rect 8051 5191 8086 5199
rect 8051 5171 8059 5191
rect 8079 5171 8086 5191
rect 8051 5166 8086 5171
rect 8051 5165 8083 5166
rect 8287 5158 8318 5365
rect 8498 5356 8530 5421
rect 8498 5336 8502 5356
rect 8523 5336 8530 5356
rect 8498 5329 8530 5336
rect 8947 5479 9022 5488
rect 8947 5446 8956 5479
rect 9009 5446 9022 5479
rect 8947 5421 9022 5446
rect 8947 5388 8961 5421
rect 9014 5388 9022 5421
rect 8947 5382 9022 5388
rect 9099 5478 9128 5498
rect 9148 5478 9155 5498
rect 9099 5473 9155 5478
rect 9546 5501 9578 5508
rect 9546 5481 9552 5501
rect 9573 5481 9578 5501
rect 8807 5273 8908 5274
rect 8705 5260 8908 5273
rect 8705 5258 8848 5260
rect 8705 5255 8782 5258
rect 8705 5228 8708 5255
rect 8737 5231 8782 5255
rect 8811 5231 8848 5258
rect 8737 5228 8848 5231
rect 8705 5227 8848 5228
rect 8884 5227 8908 5260
rect 8705 5214 8908 5227
rect 7785 5145 7949 5148
rect 8282 5145 8318 5158
rect 6984 5127 8323 5145
rect 6984 5089 6994 5127
rect 7019 5112 8323 5127
rect 7019 5089 7029 5112
rect 7785 5105 7949 5112
rect 6984 5081 7029 5089
rect 6998 5080 7029 5081
rect 8947 5066 9017 5382
rect 9099 5195 9133 5473
rect 9546 5453 9578 5481
rect 9166 5445 9578 5453
rect 9166 5419 9172 5445
rect 9198 5419 9578 5445
rect 9166 5417 9578 5419
rect 9168 5416 9208 5417
rect 9335 5391 9366 5399
rect 9335 5361 9339 5391
rect 9360 5361 9366 5391
rect 9099 5187 9134 5195
rect 9099 5167 9107 5187
rect 9127 5167 9134 5187
rect 9099 5162 9134 5167
rect 9335 5162 9366 5361
rect 9546 5352 9578 5417
rect 9546 5332 9550 5352
rect 9571 5332 9578 5352
rect 9546 5325 9578 5332
rect 9991 5478 10063 5496
rect 9991 5436 10004 5478
rect 10053 5436 10063 5478
rect 9991 5415 10063 5436
rect 9991 5373 10005 5415
rect 10054 5373 10063 5415
rect 9855 5269 9956 5270
rect 9753 5256 9956 5269
rect 9753 5254 9896 5256
rect 9753 5251 9830 5254
rect 9753 5224 9756 5251
rect 9785 5227 9830 5251
rect 9859 5227 9896 5254
rect 9785 5224 9896 5227
rect 9753 5223 9896 5224
rect 9932 5223 9956 5256
rect 9753 5210 9956 5223
rect 9099 5161 9131 5162
rect 9333 5159 9366 5162
rect 9299 5140 9367 5159
rect 9269 5128 9368 5140
rect 9269 5090 9291 5128
rect 9316 5093 9335 5128
rect 9360 5093 9368 5128
rect 9316 5090 9368 5093
rect 9269 5082 9368 5090
rect 9295 5081 9367 5082
rect 8947 5047 9026 5066
rect 8950 5027 9026 5047
rect 8943 5003 9026 5027
rect 9991 5062 10063 5373
rect 9991 5019 10067 5062
rect 8943 4937 8955 5003
rect 9009 4937 9026 5003
rect 8943 4917 9026 4937
rect 8943 4880 8960 4917
rect 9004 4903 9026 4917
rect 9992 4968 10067 5019
rect 10435 4968 10542 5561
rect 10997 5973 11104 6402
rect 11476 6161 11548 6402
rect 12171 6394 12270 6406
rect 12172 6375 12240 6394
rect 12173 6372 12206 6375
rect 12408 6372 12440 6373
rect 11583 6311 11786 6324
rect 11583 6278 11607 6311
rect 11643 6310 11786 6311
rect 11643 6307 11754 6310
rect 11643 6280 11680 6307
rect 11709 6283 11754 6307
rect 11783 6283 11786 6310
rect 11709 6280 11786 6283
rect 11643 6278 11786 6280
rect 11583 6265 11786 6278
rect 11583 6264 11684 6265
rect 11476 6119 11485 6161
rect 11534 6119 11548 6161
rect 11476 6098 11548 6119
rect 11476 6056 11486 6098
rect 11535 6056 11548 6098
rect 11476 6038 11548 6056
rect 11961 6202 11993 6209
rect 11961 6182 11968 6202
rect 11989 6182 11993 6202
rect 11961 6117 11993 6182
rect 12173 6173 12204 6372
rect 12405 6367 12440 6372
rect 12405 6347 12412 6367
rect 12432 6347 12440 6367
rect 12405 6339 12440 6347
rect 12173 6143 12179 6173
rect 12200 6143 12204 6173
rect 12173 6135 12204 6143
rect 12331 6117 12371 6118
rect 11961 6115 12373 6117
rect 11961 6089 12341 6115
rect 12367 6089 12373 6115
rect 11961 6081 12373 6089
rect 11961 6053 11993 6081
rect 12406 6061 12440 6339
rect 12522 6152 12592 6463
rect 14447 6453 14519 6454
rect 14446 6450 14535 6453
rect 13218 6448 14535 6450
rect 13215 6445 14535 6448
rect 13215 6442 14498 6445
rect 13215 6407 14454 6442
rect 14479 6407 14498 6442
rect 14523 6407 14535 6445
rect 13215 6397 14535 6407
rect 14711 6446 14747 6599
rect 14711 6423 14717 6446
rect 14741 6423 14747 6446
rect 14711 6402 14747 6423
rect 13215 6395 14500 6397
rect 13215 6385 13312 6395
rect 13221 6376 13257 6385
rect 14711 6379 14717 6402
rect 14741 6379 14747 6402
rect 12631 6307 12834 6320
rect 12631 6274 12655 6307
rect 12691 6306 12834 6307
rect 12691 6303 12802 6306
rect 12691 6276 12728 6303
rect 12757 6279 12802 6303
rect 12831 6279 12834 6306
rect 12757 6276 12834 6279
rect 12691 6274 12834 6276
rect 12631 6261 12834 6274
rect 12631 6260 12732 6261
rect 11961 6033 11966 6053
rect 11987 6033 11993 6053
rect 11961 6026 11993 6033
rect 12384 6056 12440 6061
rect 12384 6036 12391 6056
rect 12411 6036 12440 6056
rect 12517 6146 12592 6152
rect 12517 6113 12525 6146
rect 12578 6113 12592 6146
rect 12517 6088 12592 6113
rect 12517 6055 12530 6088
rect 12583 6055 12592 6088
rect 12517 6046 12592 6055
rect 13009 6198 13041 6205
rect 13009 6178 13016 6198
rect 13037 6178 13041 6198
rect 13009 6113 13041 6178
rect 13221 6169 13252 6376
rect 13456 6368 13488 6369
rect 14711 6368 14747 6379
rect 13453 6363 13488 6368
rect 13453 6343 13460 6363
rect 13480 6343 13488 6363
rect 13453 6335 13488 6343
rect 13221 6139 13227 6169
rect 13248 6139 13252 6169
rect 13221 6131 13252 6139
rect 13379 6113 13419 6114
rect 13009 6111 13421 6113
rect 13009 6085 13389 6111
rect 13415 6085 13421 6111
rect 13009 6077 13421 6085
rect 13009 6049 13041 6077
rect 13454 6057 13488 6335
rect 12517 6041 12575 6046
rect 12384 6029 12440 6036
rect 13009 6029 13014 6049
rect 13035 6029 13041 6049
rect 12384 6028 12419 6029
rect 13009 6022 13041 6029
rect 13432 6052 13488 6057
rect 13432 6032 13439 6052
rect 13459 6032 13488 6052
rect 13432 6025 13488 6032
rect 13432 6024 13467 6025
rect 11675 5973 11786 5977
rect 13550 5973 14709 5974
rect 10997 5955 14709 5973
rect 10997 5935 11683 5955
rect 11702 5935 11760 5955
rect 11779 5951 14709 5955
rect 11779 5935 12731 5951
rect 10997 5931 12731 5935
rect 12750 5931 12808 5951
rect 12827 5931 14709 5951
rect 10997 5917 14709 5931
rect 10997 5294 11104 5917
rect 12723 5914 12834 5917
rect 11483 5868 11547 5872
rect 11479 5862 11547 5868
rect 11479 5829 11496 5862
rect 11536 5829 11547 5862
rect 11479 5817 11547 5829
rect 12530 5831 12595 5853
rect 11479 5815 11536 5817
rect 11483 5454 11534 5815
rect 12530 5792 12547 5831
rect 12592 5792 12595 5831
rect 15616 5829 15668 8135
rect 15777 8112 15812 8178
rect 15777 6796 15811 8112
rect 16115 7965 16220 13065
rect 17179 13052 21252 13066
rect 17179 13032 19422 13052
rect 19441 13032 19499 13052
rect 19518 13048 21252 13052
rect 19518 13032 20470 13048
rect 17179 13028 20470 13032
rect 20489 13028 20547 13048
rect 20566 13028 21252 13048
rect 17179 13010 21252 13028
rect 17179 13009 18699 13010
rect 20463 13006 20574 13010
rect 18782 12958 18817 12959
rect 18761 12951 18817 12958
rect 18761 12931 18790 12951
rect 18810 12931 18817 12951
rect 18761 12926 18817 12931
rect 19208 12954 19240 12961
rect 19830 12954 19865 12955
rect 19208 12934 19214 12954
rect 19235 12934 19240 12954
rect 19809 12947 19865 12954
rect 19674 12937 19732 12942
rect 18761 12648 18795 12926
rect 19208 12906 19240 12934
rect 18828 12898 19240 12906
rect 18828 12872 18834 12898
rect 18860 12872 19240 12898
rect 18828 12870 19240 12872
rect 18830 12869 18870 12870
rect 18997 12844 19028 12852
rect 18997 12814 19001 12844
rect 19022 12814 19028 12844
rect 18761 12640 18796 12648
rect 18761 12620 18769 12640
rect 18789 12620 18796 12640
rect 18761 12615 18796 12620
rect 18761 12614 18793 12615
rect 18997 12614 19028 12814
rect 19208 12805 19240 12870
rect 19208 12785 19212 12805
rect 19233 12785 19240 12805
rect 19208 12778 19240 12785
rect 19657 12928 19732 12937
rect 19657 12895 19666 12928
rect 19719 12895 19732 12928
rect 19657 12870 19732 12895
rect 19657 12837 19671 12870
rect 19724 12837 19732 12870
rect 19657 12831 19732 12837
rect 19809 12927 19838 12947
rect 19858 12927 19865 12947
rect 19809 12922 19865 12927
rect 20256 12950 20288 12957
rect 20256 12930 20262 12950
rect 20283 12930 20288 12950
rect 19517 12722 19618 12723
rect 19415 12709 19618 12722
rect 19415 12707 19558 12709
rect 19415 12704 19492 12707
rect 19415 12677 19418 12704
rect 19447 12680 19492 12704
rect 19521 12680 19558 12707
rect 19447 12677 19558 12680
rect 19415 12676 19558 12677
rect 19594 12676 19618 12709
rect 19415 12663 19618 12676
rect 18994 12607 19033 12614
rect 18992 12590 19033 12607
rect 18994 12565 19033 12590
rect 17688 12557 19033 12565
rect 17688 12529 17703 12557
rect 17731 12531 19033 12557
rect 17731 12529 19030 12531
rect 17688 12524 19030 12529
rect 19657 12520 19727 12831
rect 19809 12644 19843 12922
rect 20256 12902 20288 12930
rect 19876 12894 20288 12902
rect 19876 12868 19882 12894
rect 19908 12868 20288 12894
rect 19876 12866 20288 12868
rect 19878 12865 19918 12866
rect 20045 12840 20076 12848
rect 20045 12810 20049 12840
rect 20070 12810 20076 12840
rect 19809 12636 19844 12644
rect 19809 12616 19817 12636
rect 19837 12616 19844 12636
rect 19809 12611 19844 12616
rect 20045 12611 20076 12810
rect 20256 12801 20288 12866
rect 20256 12781 20260 12801
rect 20281 12781 20288 12801
rect 20256 12774 20288 12781
rect 20701 12927 20773 12945
rect 20701 12885 20714 12927
rect 20763 12885 20773 12927
rect 20701 12864 20773 12885
rect 20701 12822 20715 12864
rect 20764 12822 20773 12864
rect 20565 12718 20666 12719
rect 20463 12705 20666 12718
rect 20463 12703 20606 12705
rect 20463 12700 20540 12703
rect 20463 12673 20466 12700
rect 20495 12676 20540 12700
rect 20569 12676 20606 12703
rect 20495 12673 20606 12676
rect 20463 12672 20606 12673
rect 20642 12672 20666 12705
rect 20463 12659 20666 12672
rect 19809 12610 19841 12611
rect 20043 12608 20076 12611
rect 20009 12589 20077 12608
rect 19979 12577 20078 12589
rect 20701 12581 20773 12822
rect 21145 12581 21252 13010
rect 21964 13432 22071 13792
rect 22443 13620 22515 13972
rect 23139 13911 23211 13912
rect 23138 13903 23237 13911
rect 23138 13900 23190 13903
rect 23138 13865 23146 13900
rect 23171 13865 23190 13900
rect 23215 13865 23237 13903
rect 23138 13853 23237 13865
rect 23139 13834 23207 13853
rect 23140 13831 23173 13834
rect 23375 13831 23407 13832
rect 22550 13770 22753 13783
rect 22550 13737 22574 13770
rect 22610 13769 22753 13770
rect 22610 13766 22721 13769
rect 22610 13739 22647 13766
rect 22676 13742 22721 13766
rect 22750 13742 22753 13769
rect 22676 13739 22753 13742
rect 22610 13737 22753 13739
rect 22550 13724 22753 13737
rect 22550 13723 22651 13724
rect 22443 13578 22452 13620
rect 22501 13578 22515 13620
rect 22443 13557 22515 13578
rect 22443 13515 22453 13557
rect 22502 13515 22515 13557
rect 22443 13497 22515 13515
rect 22928 13661 22960 13668
rect 22928 13641 22935 13661
rect 22956 13641 22960 13661
rect 22928 13576 22960 13641
rect 23140 13632 23171 13831
rect 23372 13826 23407 13831
rect 23372 13806 23379 13826
rect 23399 13806 23407 13826
rect 23372 13798 23407 13806
rect 23140 13602 23146 13632
rect 23167 13602 23171 13632
rect 23140 13594 23171 13602
rect 23298 13576 23338 13577
rect 22928 13574 23340 13576
rect 22928 13548 23308 13574
rect 23334 13548 23340 13574
rect 22928 13540 23340 13548
rect 22928 13512 22960 13540
rect 23373 13520 23407 13798
rect 23489 13611 23559 13972
rect 24189 13912 24261 13913
rect 24188 13904 24277 13912
rect 24188 13901 24240 13904
rect 24188 13866 24196 13901
rect 24221 13866 24240 13901
rect 24265 13866 24277 13904
rect 24188 13854 24277 13866
rect 24188 13853 24257 13854
rect 24188 13835 24224 13853
rect 23598 13766 23801 13779
rect 23598 13733 23622 13766
rect 23658 13765 23801 13766
rect 23658 13762 23769 13765
rect 23658 13735 23695 13762
rect 23724 13738 23769 13762
rect 23798 13738 23801 13765
rect 23724 13735 23801 13738
rect 23658 13733 23801 13735
rect 23598 13720 23801 13733
rect 23598 13719 23699 13720
rect 22928 13492 22933 13512
rect 22954 13492 22960 13512
rect 22928 13485 22960 13492
rect 23351 13515 23407 13520
rect 23351 13495 23358 13515
rect 23378 13495 23407 13515
rect 23484 13605 23559 13611
rect 23484 13572 23492 13605
rect 23545 13572 23559 13605
rect 23484 13547 23559 13572
rect 23484 13514 23497 13547
rect 23550 13514 23559 13547
rect 23484 13505 23559 13514
rect 23976 13657 24008 13664
rect 23976 13637 23983 13657
rect 24004 13637 24008 13657
rect 23976 13572 24008 13637
rect 24188 13628 24219 13835
rect 24423 13827 24455 13828
rect 24420 13822 24455 13827
rect 24420 13802 24427 13822
rect 24447 13802 24455 13822
rect 24420 13794 24455 13802
rect 24188 13598 24194 13628
rect 24215 13598 24219 13628
rect 24188 13590 24219 13598
rect 24346 13572 24386 13573
rect 23976 13570 24388 13572
rect 23976 13544 24356 13570
rect 24382 13544 24388 13570
rect 23976 13536 24388 13544
rect 23976 13508 24008 13536
rect 24421 13516 24455 13794
rect 24604 13609 24666 13972
rect 24758 13967 24879 13983
rect 24773 13612 24855 13967
rect 26040 13761 26089 14098
rect 26557 13773 26695 13777
rect 26537 13761 26695 13773
rect 26030 13745 26695 13761
rect 26030 13678 26589 13745
rect 26675 13678 26695 13745
rect 26030 13662 26695 13678
rect 24604 13590 24668 13609
rect 24604 13551 24617 13590
rect 24651 13551 24668 13590
rect 24604 13532 24668 13551
rect 24773 13571 24794 13612
rect 24830 13571 24855 13612
rect 24773 13542 24855 13571
rect 23484 13500 23542 13505
rect 23351 13488 23407 13495
rect 23976 13488 23981 13508
rect 24002 13488 24008 13508
rect 23351 13487 23386 13488
rect 23976 13481 24008 13488
rect 24399 13511 24455 13516
rect 24399 13491 24406 13511
rect 24426 13491 24455 13511
rect 24399 13484 24455 13491
rect 24399 13483 24434 13484
rect 22642 13432 22753 13436
rect 24425 13432 25538 13433
rect 21964 13414 25538 13432
rect 21964 13394 22650 13414
rect 22669 13394 22727 13414
rect 22746 13410 25538 13414
rect 22746 13394 23698 13410
rect 21964 13390 23698 13394
rect 23717 13390 23775 13410
rect 23794 13390 25538 13410
rect 21964 13376 25538 13390
rect 21964 12753 22071 13376
rect 23690 13373 23801 13376
rect 22450 13327 22514 13331
rect 22446 13321 22514 13327
rect 22446 13288 22463 13321
rect 22503 13288 22514 13321
rect 22446 13276 22514 13288
rect 23497 13290 23562 13312
rect 22446 13274 22503 13276
rect 22450 12913 22501 13274
rect 23497 13251 23514 13290
rect 23559 13251 23562 13290
rect 23138 13206 23173 13208
rect 23138 13197 23242 13206
rect 23138 13196 23189 13197
rect 23138 13176 23141 13196
rect 23166 13177 23189 13196
rect 23221 13177 23242 13197
rect 23166 13176 23242 13177
rect 23138 13169 23242 13176
rect 23138 13157 23173 13169
rect 22550 13091 22753 13104
rect 22550 13058 22574 13091
rect 22610 13090 22753 13091
rect 22610 13087 22721 13090
rect 22610 13060 22647 13087
rect 22676 13063 22721 13087
rect 22750 13063 22753 13090
rect 22676 13060 22753 13063
rect 22610 13058 22753 13060
rect 22550 13045 22753 13058
rect 22550 13044 22651 13045
rect 22928 12982 22960 12989
rect 22928 12962 22935 12982
rect 22956 12962 22960 12982
rect 22439 12904 22504 12913
rect 22439 12867 22449 12904
rect 22489 12870 22504 12904
rect 22928 12897 22960 12962
rect 23140 12953 23171 13157
rect 23375 13152 23407 13153
rect 23372 13147 23407 13152
rect 23372 13127 23379 13147
rect 23399 13127 23407 13147
rect 23372 13119 23407 13127
rect 23140 12923 23146 12953
rect 23167 12923 23171 12953
rect 23140 12915 23171 12923
rect 23298 12897 23338 12898
rect 22928 12895 23340 12897
rect 22489 12867 22506 12870
rect 22439 12848 22506 12867
rect 22439 12827 22453 12848
rect 22489 12827 22506 12848
rect 22439 12820 22506 12827
rect 22928 12869 23308 12895
rect 23334 12869 23340 12895
rect 22928 12861 23340 12869
rect 22928 12833 22960 12861
rect 23373 12841 23407 13119
rect 23497 12951 23562 13251
rect 24768 13275 24861 13290
rect 24768 13231 24783 13275
rect 24843 13231 24861 13275
rect 22928 12813 22933 12833
rect 22954 12813 22960 12833
rect 22928 12806 22960 12813
rect 23351 12836 23407 12841
rect 23351 12816 23358 12836
rect 23378 12816 23407 12836
rect 23351 12809 23407 12816
rect 23487 12940 23567 12951
rect 23487 12914 23504 12940
rect 23544 12914 23567 12940
rect 23487 12887 23567 12914
rect 23487 12861 23508 12887
rect 23548 12861 23567 12887
rect 23487 12842 23567 12861
rect 23487 12816 23511 12842
rect 23551 12816 23567 12842
rect 23351 12808 23386 12809
rect 23487 12804 23567 12816
rect 24768 12858 24861 13231
rect 25045 13086 25248 13099
rect 25045 13053 25069 13086
rect 25105 13085 25248 13086
rect 25105 13082 25216 13085
rect 25105 13055 25142 13082
rect 25171 13058 25216 13082
rect 25245 13058 25248 13085
rect 25171 13055 25248 13058
rect 25105 13053 25248 13055
rect 25045 13040 25248 13053
rect 25045 13039 25146 13040
rect 24768 12817 24783 12858
rect 24837 12817 24861 12858
rect 24768 12810 24861 12817
rect 25423 12977 25455 12984
rect 25423 12957 25430 12977
rect 25451 12957 25455 12977
rect 25423 12892 25455 12957
rect 25635 12948 25666 13149
rect 25870 13147 25902 13148
rect 25867 13142 25902 13147
rect 25867 13122 25874 13142
rect 25894 13122 25902 13142
rect 25867 13114 25902 13122
rect 25635 12918 25641 12948
rect 25662 12918 25666 12948
rect 25635 12910 25666 12918
rect 25793 12892 25833 12893
rect 25423 12890 25835 12892
rect 25423 12864 25803 12890
rect 25829 12864 25835 12890
rect 25423 12856 25835 12864
rect 25423 12828 25455 12856
rect 25868 12836 25902 13114
rect 25423 12808 25428 12828
rect 25449 12808 25455 12828
rect 25423 12801 25455 12808
rect 25846 12831 25902 12836
rect 25846 12811 25853 12831
rect 25873 12811 25902 12831
rect 25846 12804 25902 12811
rect 25846 12803 25881 12804
rect 22642 12753 22753 12757
rect 24384 12753 25933 12756
rect 21962 12735 25933 12753
rect 21962 12715 22650 12735
rect 22669 12715 22727 12735
rect 22746 12730 25933 12735
rect 22746 12715 25145 12730
rect 21962 12710 25145 12715
rect 25164 12710 25222 12730
rect 25241 12710 25933 12730
rect 21962 12700 25933 12710
rect 21962 12697 22587 12700
rect 22774 12697 25933 12700
rect 19979 12539 20001 12577
rect 20026 12542 20045 12577
rect 20070 12542 20078 12577
rect 20026 12539 20078 12542
rect 19979 12531 20078 12539
rect 20005 12530 20077 12531
rect 19656 12504 19727 12520
rect 19656 12488 19676 12504
rect 19657 12458 19676 12488
rect 19659 12438 19676 12458
rect 19706 12458 19727 12504
rect 20699 12500 20777 12581
rect 21144 12526 21252 12581
rect 19706 12438 19726 12458
rect 19659 12419 19726 12438
rect 20699 12398 20778 12500
rect 20663 12380 20784 12398
rect 20663 12378 20734 12380
rect 20663 12337 20678 12378
rect 20715 12339 20734 12378
rect 20771 12339 20784 12380
rect 20715 12337 20784 12339
rect 20663 12327 20784 12337
rect 17968 12299 18079 12302
rect 17179 12298 18832 12299
rect 21145 12298 21252 12526
rect 21964 12469 22071 12697
rect 24384 12696 25933 12697
rect 25137 12693 25248 12696
rect 22432 12658 22553 12668
rect 22432 12656 22501 12658
rect 22432 12615 22445 12656
rect 22482 12617 22501 12656
rect 22538 12617 22553 12658
rect 22482 12615 22553 12617
rect 22432 12597 22553 12615
rect 25637 12638 25723 12642
rect 25637 12620 25652 12638
rect 25704 12620 25723 12638
rect 25637 12611 25723 12620
rect 22438 12495 22517 12597
rect 23490 12557 23557 12576
rect 23490 12537 23510 12557
rect 21964 12414 22072 12469
rect 22439 12414 22517 12495
rect 23489 12491 23510 12537
rect 23540 12537 23557 12557
rect 23540 12507 23559 12537
rect 23540 12491 23560 12507
rect 23489 12475 23560 12491
rect 23139 12464 23211 12465
rect 23138 12456 23237 12464
rect 23138 12453 23190 12456
rect 23138 12418 23146 12453
rect 23171 12418 23190 12453
rect 23215 12418 23237 12456
rect 17179 12295 20442 12298
rect 20629 12295 21254 12298
rect 17179 12285 21254 12295
rect 17179 12265 17975 12285
rect 17994 12265 18052 12285
rect 18071 12280 21254 12285
rect 18071 12265 20470 12280
rect 17179 12260 20470 12265
rect 20489 12260 20547 12280
rect 20566 12260 21254 12280
rect 17179 12242 21254 12260
rect 17179 12239 18832 12242
rect 20463 12238 20574 12242
rect 17335 12191 17370 12192
rect 17314 12184 17370 12191
rect 17314 12164 17343 12184
rect 17363 12164 17370 12184
rect 17314 12159 17370 12164
rect 17761 12187 17793 12194
rect 17761 12167 17767 12187
rect 17788 12167 17793 12187
rect 17314 11881 17348 12159
rect 17761 12139 17793 12167
rect 19649 12179 19729 12191
rect 19830 12186 19865 12187
rect 17381 12131 17793 12139
rect 17381 12105 17387 12131
rect 17413 12105 17793 12131
rect 18179 12145 18616 12158
rect 18179 12122 18192 12145
rect 18218 12138 18616 12145
rect 18218 12122 18572 12138
rect 18179 12115 18572 12122
rect 18598 12115 18616 12138
rect 18179 12109 18616 12115
rect 19649 12153 19665 12179
rect 19705 12153 19729 12179
rect 19649 12134 19729 12153
rect 17381 12103 17793 12105
rect 17383 12102 17423 12103
rect 17550 12077 17581 12085
rect 17550 12047 17554 12077
rect 17575 12047 17581 12077
rect 17314 11873 17349 11881
rect 17314 11853 17322 11873
rect 17342 11853 17349 11873
rect 17314 11848 17349 11853
rect 17314 11847 17346 11848
rect 17550 11840 17581 12047
rect 17761 12038 17793 12103
rect 19649 12108 19668 12134
rect 19708 12108 19729 12134
rect 19649 12081 19729 12108
rect 19649 12055 19672 12081
rect 19712 12055 19729 12081
rect 19649 12044 19729 12055
rect 19809 12179 19865 12186
rect 19809 12159 19838 12179
rect 19858 12159 19865 12179
rect 19809 12154 19865 12159
rect 20256 12182 20288 12189
rect 20256 12162 20262 12182
rect 20283 12162 20288 12182
rect 17761 12018 17765 12038
rect 17786 12018 17793 12038
rect 17761 12011 17793 12018
rect 18070 11955 18171 11956
rect 17968 11942 18171 11955
rect 17968 11940 18111 11942
rect 17968 11937 18045 11940
rect 17968 11910 17971 11937
rect 18000 11913 18045 11937
rect 18074 11913 18111 11940
rect 18000 11910 18111 11913
rect 17968 11909 18111 11910
rect 18147 11909 18171 11942
rect 17968 11896 18171 11909
rect 17548 11834 17581 11840
rect 17544 11830 17581 11834
rect 17544 11820 17582 11830
rect 17544 11807 17554 11820
rect 17545 11783 17554 11807
rect 17571 11783 17582 11820
rect 17545 11762 17582 11783
rect 19654 11744 19719 12044
rect 19809 11876 19843 12154
rect 20256 12134 20288 12162
rect 19876 12126 20288 12134
rect 19876 12100 19882 12126
rect 19908 12100 20288 12126
rect 20710 12168 20777 12175
rect 20710 12147 20727 12168
rect 20763 12147 20777 12168
rect 20710 12128 20777 12147
rect 20710 12125 20727 12128
rect 19876 12098 20288 12100
rect 19878 12097 19918 12098
rect 20045 12072 20076 12080
rect 20045 12042 20049 12072
rect 20070 12042 20076 12072
rect 19809 11868 19844 11876
rect 19809 11848 19817 11868
rect 19837 11848 19844 11868
rect 19809 11843 19844 11848
rect 19809 11842 19841 11843
rect 20045 11838 20076 12042
rect 20256 12033 20288 12098
rect 20712 12091 20727 12125
rect 20767 12091 20777 12128
rect 20712 12082 20777 12091
rect 20256 12013 20260 12033
rect 20281 12013 20288 12033
rect 20256 12006 20288 12013
rect 20565 11950 20666 11951
rect 20463 11937 20666 11950
rect 20463 11935 20606 11937
rect 20463 11932 20540 11935
rect 20463 11905 20466 11932
rect 20495 11908 20540 11932
rect 20569 11908 20606 11935
rect 20495 11905 20606 11908
rect 20463 11904 20606 11905
rect 20642 11904 20666 11937
rect 20463 11891 20666 11904
rect 20043 11826 20078 11838
rect 19974 11819 20078 11826
rect 19974 11818 20050 11819
rect 19974 11798 19995 11818
rect 20027 11799 20050 11818
rect 20075 11799 20078 11819
rect 20027 11798 20078 11799
rect 19974 11789 20078 11798
rect 20043 11787 20078 11789
rect 19654 11705 19657 11744
rect 19702 11705 19719 11744
rect 20715 11721 20766 12082
rect 20713 11719 20770 11721
rect 19654 11683 19719 11705
rect 20702 11707 20770 11719
rect 20702 11674 20713 11707
rect 20753 11674 20770 11707
rect 20702 11668 20770 11674
rect 20702 11664 20766 11668
rect 19415 11619 19526 11622
rect 21145 11619 21252 12242
rect 16802 11605 21252 11619
rect 16802 11585 19422 11605
rect 19441 11585 19499 11605
rect 19518 11601 21252 11605
rect 19518 11585 20470 11601
rect 16802 11581 20470 11585
rect 20489 11581 20547 11601
rect 20566 11581 21252 11601
rect 16802 11567 21252 11581
rect 17221 11563 21252 11567
rect 17221 11562 18791 11563
rect 20463 11559 20574 11563
rect 18782 11511 18817 11512
rect 18761 11504 18817 11511
rect 18761 11484 18790 11504
rect 18810 11484 18817 11504
rect 18761 11479 18817 11484
rect 19208 11507 19240 11514
rect 19830 11507 19865 11508
rect 19208 11487 19214 11507
rect 19235 11487 19240 11507
rect 19809 11500 19865 11507
rect 19674 11490 19732 11495
rect 18761 11201 18795 11479
rect 19208 11459 19240 11487
rect 18828 11451 19240 11459
rect 18828 11425 18834 11451
rect 18860 11425 19240 11451
rect 18828 11423 19240 11425
rect 18830 11422 18870 11423
rect 18997 11397 19028 11405
rect 18997 11367 19001 11397
rect 19022 11367 19028 11397
rect 18761 11193 18796 11201
rect 18761 11173 18769 11193
rect 18789 11173 18796 11193
rect 18761 11168 18796 11173
rect 18761 11167 18793 11168
rect 18997 11160 19028 11367
rect 19208 11358 19240 11423
rect 19208 11338 19212 11358
rect 19233 11338 19240 11358
rect 19208 11331 19240 11338
rect 19657 11481 19732 11490
rect 19657 11448 19666 11481
rect 19719 11448 19732 11481
rect 19657 11423 19732 11448
rect 19657 11390 19671 11423
rect 19724 11390 19732 11423
rect 19657 11384 19732 11390
rect 19809 11480 19838 11500
rect 19858 11480 19865 11500
rect 19809 11475 19865 11480
rect 20256 11503 20288 11510
rect 20256 11483 20262 11503
rect 20283 11483 20288 11503
rect 19517 11275 19618 11276
rect 19415 11262 19618 11275
rect 19415 11260 19558 11262
rect 19415 11257 19492 11260
rect 19415 11230 19418 11257
rect 19447 11233 19492 11257
rect 19521 11233 19558 11260
rect 19447 11230 19558 11233
rect 19415 11229 19558 11230
rect 19594 11229 19618 11262
rect 19415 11216 19618 11229
rect 18495 11147 18659 11150
rect 18992 11147 19028 11160
rect 17694 11129 19033 11147
rect 17694 11091 17704 11129
rect 17729 11114 19033 11129
rect 17729 11091 17739 11114
rect 18495 11107 18659 11114
rect 17694 11083 17739 11091
rect 17708 11082 17739 11083
rect 19657 11068 19727 11384
rect 19809 11197 19843 11475
rect 20256 11455 20288 11483
rect 19876 11447 20288 11455
rect 19876 11421 19882 11447
rect 19908 11421 20288 11447
rect 19876 11419 20288 11421
rect 19878 11418 19918 11419
rect 20045 11393 20076 11401
rect 20045 11363 20049 11393
rect 20070 11363 20076 11393
rect 19809 11189 19844 11197
rect 19809 11169 19817 11189
rect 19837 11169 19844 11189
rect 19809 11164 19844 11169
rect 20045 11164 20076 11363
rect 20256 11354 20288 11419
rect 20256 11334 20260 11354
rect 20281 11334 20288 11354
rect 20256 11327 20288 11334
rect 20701 11480 20773 11498
rect 20701 11438 20714 11480
rect 20763 11438 20773 11480
rect 20701 11417 20773 11438
rect 20701 11375 20715 11417
rect 20764 11375 20773 11417
rect 20565 11271 20666 11272
rect 20463 11258 20666 11271
rect 20463 11256 20606 11258
rect 20463 11253 20540 11256
rect 20463 11226 20466 11253
rect 20495 11229 20540 11253
rect 20569 11229 20606 11256
rect 20495 11226 20606 11229
rect 20463 11225 20606 11226
rect 20642 11225 20666 11258
rect 20463 11212 20666 11225
rect 19809 11163 19841 11164
rect 20043 11161 20076 11164
rect 20009 11142 20077 11161
rect 19979 11130 20078 11142
rect 19979 11092 20001 11130
rect 20026 11095 20045 11130
rect 20070 11095 20078 11130
rect 20026 11092 20078 11095
rect 19979 11084 20078 11092
rect 20005 11083 20077 11084
rect 19657 11049 19736 11068
rect 19660 11029 19736 11049
rect 19653 11005 19736 11029
rect 20701 11064 20773 11375
rect 20701 11021 20777 11064
rect 19653 10939 19665 11005
rect 19719 10939 19736 11005
rect 19653 10919 19736 10939
rect 19653 10882 19670 10919
rect 19714 10905 19736 10919
rect 20702 10970 20777 11021
rect 21145 10970 21252 11563
rect 21964 11985 22071 12414
rect 22443 12173 22515 12414
rect 23138 12406 23237 12418
rect 23139 12387 23207 12406
rect 23140 12384 23173 12387
rect 23375 12384 23407 12385
rect 22550 12323 22753 12336
rect 22550 12290 22574 12323
rect 22610 12322 22753 12323
rect 22610 12319 22721 12322
rect 22610 12292 22647 12319
rect 22676 12295 22721 12319
rect 22750 12295 22753 12322
rect 22676 12292 22753 12295
rect 22610 12290 22753 12292
rect 22550 12277 22753 12290
rect 22550 12276 22651 12277
rect 22443 12131 22452 12173
rect 22501 12131 22515 12173
rect 22443 12110 22515 12131
rect 22443 12068 22453 12110
rect 22502 12068 22515 12110
rect 22443 12050 22515 12068
rect 22928 12214 22960 12221
rect 22928 12194 22935 12214
rect 22956 12194 22960 12214
rect 22928 12129 22960 12194
rect 23140 12185 23171 12384
rect 23372 12379 23407 12384
rect 23372 12359 23379 12379
rect 23399 12359 23407 12379
rect 23372 12351 23407 12359
rect 23140 12155 23146 12185
rect 23167 12155 23171 12185
rect 23140 12147 23171 12155
rect 23298 12129 23338 12130
rect 22928 12127 23340 12129
rect 22928 12101 23308 12127
rect 23334 12101 23340 12127
rect 22928 12093 23340 12101
rect 22928 12065 22960 12093
rect 23373 12073 23407 12351
rect 23489 12164 23559 12475
rect 25414 12465 25486 12466
rect 25413 12462 25502 12465
rect 24185 12460 25502 12462
rect 24182 12457 25502 12460
rect 24182 12454 25465 12457
rect 24182 12419 25421 12454
rect 25446 12419 25465 12454
rect 25490 12419 25502 12457
rect 24182 12409 25502 12419
rect 25678 12458 25714 12611
rect 25678 12435 25684 12458
rect 25708 12435 25714 12458
rect 25678 12414 25714 12435
rect 24182 12407 25467 12409
rect 24182 12397 24279 12407
rect 24188 12388 24224 12397
rect 25678 12391 25684 12414
rect 25708 12391 25714 12414
rect 23598 12319 23801 12332
rect 23598 12286 23622 12319
rect 23658 12318 23801 12319
rect 23658 12315 23769 12318
rect 23658 12288 23695 12315
rect 23724 12291 23769 12315
rect 23798 12291 23801 12318
rect 23724 12288 23801 12291
rect 23658 12286 23801 12288
rect 23598 12273 23801 12286
rect 23598 12272 23699 12273
rect 22928 12045 22933 12065
rect 22954 12045 22960 12065
rect 22928 12038 22960 12045
rect 23351 12068 23407 12073
rect 23351 12048 23358 12068
rect 23378 12048 23407 12068
rect 23484 12158 23559 12164
rect 23484 12125 23492 12158
rect 23545 12125 23559 12158
rect 23484 12100 23559 12125
rect 23484 12067 23497 12100
rect 23550 12067 23559 12100
rect 23484 12058 23559 12067
rect 23976 12210 24008 12217
rect 23976 12190 23983 12210
rect 24004 12190 24008 12210
rect 23976 12125 24008 12190
rect 24188 12181 24219 12388
rect 24423 12380 24455 12381
rect 25678 12380 25714 12391
rect 24420 12375 24455 12380
rect 24420 12355 24427 12375
rect 24447 12355 24455 12375
rect 24420 12347 24455 12355
rect 24188 12151 24194 12181
rect 24215 12151 24219 12181
rect 24188 12143 24219 12151
rect 24346 12125 24386 12126
rect 23976 12123 24388 12125
rect 23976 12097 24356 12123
rect 24382 12097 24388 12123
rect 23976 12089 24388 12097
rect 23976 12061 24008 12089
rect 24421 12069 24455 12347
rect 23484 12053 23542 12058
rect 23351 12041 23407 12048
rect 23976 12041 23981 12061
rect 24002 12041 24008 12061
rect 23351 12040 23386 12041
rect 23976 12034 24008 12041
rect 24399 12064 24455 12069
rect 24399 12044 24406 12064
rect 24426 12044 24455 12064
rect 24399 12037 24455 12044
rect 24399 12036 24434 12037
rect 22642 11985 22753 11989
rect 24517 11985 25758 11986
rect 21964 11967 25758 11985
rect 21964 11947 22650 11967
rect 22669 11947 22727 11967
rect 22746 11963 25758 11967
rect 22746 11947 23698 11963
rect 21964 11943 23698 11947
rect 23717 11943 23775 11963
rect 23794 11943 25758 11963
rect 21964 11929 25758 11943
rect 21964 11306 22071 11929
rect 23690 11926 23801 11929
rect 22450 11880 22514 11884
rect 22446 11874 22514 11880
rect 22446 11841 22463 11874
rect 22503 11841 22514 11874
rect 22446 11829 22514 11841
rect 23497 11843 23562 11865
rect 22446 11827 22503 11829
rect 22450 11466 22501 11827
rect 23497 11804 23514 11843
rect 23559 11804 23562 11843
rect 23138 11759 23173 11761
rect 23138 11750 23242 11759
rect 23138 11749 23189 11750
rect 23138 11729 23141 11749
rect 23166 11730 23189 11749
rect 23221 11730 23242 11750
rect 23166 11729 23242 11730
rect 23138 11722 23242 11729
rect 23138 11710 23173 11722
rect 22550 11644 22753 11657
rect 22550 11611 22574 11644
rect 22610 11643 22753 11644
rect 22610 11640 22721 11643
rect 22610 11613 22647 11640
rect 22676 11616 22721 11640
rect 22750 11616 22753 11643
rect 22676 11613 22753 11616
rect 22610 11611 22753 11613
rect 22550 11598 22753 11611
rect 22550 11597 22651 11598
rect 22928 11535 22960 11542
rect 22928 11515 22935 11535
rect 22956 11515 22960 11535
rect 22439 11457 22504 11466
rect 22439 11420 22449 11457
rect 22489 11423 22504 11457
rect 22928 11450 22960 11515
rect 23140 11506 23171 11710
rect 23375 11705 23407 11706
rect 23372 11700 23407 11705
rect 23372 11680 23379 11700
rect 23399 11680 23407 11700
rect 23372 11672 23407 11680
rect 23140 11476 23146 11506
rect 23167 11476 23171 11506
rect 23140 11468 23171 11476
rect 23298 11450 23338 11451
rect 22928 11448 23340 11450
rect 22489 11420 22506 11423
rect 22439 11401 22506 11420
rect 22439 11380 22453 11401
rect 22489 11380 22506 11401
rect 22439 11373 22506 11380
rect 22928 11422 23308 11448
rect 23334 11422 23340 11448
rect 22928 11414 23340 11422
rect 22928 11386 22960 11414
rect 23373 11394 23407 11672
rect 23497 11504 23562 11804
rect 25676 11798 25781 11807
rect 25676 11793 25730 11798
rect 25676 11772 25689 11793
rect 25709 11777 25730 11793
rect 25750 11777 25781 11798
rect 25709 11772 25781 11777
rect 25676 11741 25781 11772
rect 25679 11724 25714 11741
rect 25678 11706 25714 11724
rect 25088 11641 25291 11654
rect 25088 11608 25112 11641
rect 25148 11640 25291 11641
rect 25148 11637 25259 11640
rect 25148 11610 25185 11637
rect 25214 11613 25259 11637
rect 25288 11613 25291 11640
rect 25214 11610 25291 11613
rect 25148 11608 25291 11610
rect 25088 11595 25291 11608
rect 25088 11594 25189 11595
rect 25466 11532 25498 11539
rect 25466 11512 25473 11532
rect 25494 11512 25498 11532
rect 22928 11366 22933 11386
rect 22954 11366 22960 11386
rect 22928 11359 22960 11366
rect 23351 11389 23407 11394
rect 23351 11369 23358 11389
rect 23378 11369 23407 11389
rect 23351 11362 23407 11369
rect 23487 11493 23567 11504
rect 23487 11467 23504 11493
rect 23544 11467 23567 11493
rect 23487 11440 23567 11467
rect 23487 11414 23508 11440
rect 23548 11414 23567 11440
rect 23487 11395 23567 11414
rect 23487 11369 23511 11395
rect 23551 11369 23567 11395
rect 23351 11361 23386 11362
rect 23487 11357 23567 11369
rect 25466 11447 25498 11512
rect 25678 11503 25709 11706
rect 25913 11702 25945 11703
rect 25910 11697 25945 11702
rect 25910 11677 25917 11697
rect 25937 11677 25945 11697
rect 25910 11669 25945 11677
rect 25678 11473 25684 11503
rect 25705 11473 25709 11503
rect 25678 11465 25709 11473
rect 25836 11447 25876 11448
rect 25466 11445 25878 11447
rect 25466 11419 25846 11445
rect 25872 11419 25878 11445
rect 25466 11411 25878 11419
rect 25466 11383 25498 11411
rect 25911 11391 25945 11669
rect 25466 11363 25471 11383
rect 25492 11363 25498 11383
rect 25466 11356 25498 11363
rect 25889 11386 25945 11391
rect 25889 11366 25896 11386
rect 25916 11366 25945 11386
rect 25889 11359 25945 11366
rect 25889 11358 25924 11359
rect 22642 11306 22753 11310
rect 24397 11306 24604 11307
rect 25180 11306 25291 11307
rect 21962 11288 25982 11306
rect 21962 11268 22650 11288
rect 22669 11268 22727 11288
rect 22746 11285 25982 11288
rect 22746 11268 25188 11285
rect 21962 11265 25188 11268
rect 25207 11265 25265 11285
rect 25284 11265 25982 11285
rect 21962 11250 25982 11265
rect 21964 11062 22071 11250
rect 24559 11248 25982 11250
rect 22432 11211 22553 11221
rect 22432 11209 22501 11211
rect 22432 11168 22445 11209
rect 22482 11170 22501 11209
rect 22538 11170 22553 11211
rect 22482 11168 22553 11170
rect 22432 11150 22553 11168
rect 21964 11058 22072 11062
rect 22438 11058 22515 11150
rect 23488 11146 23564 11162
rect 23488 11123 23503 11146
rect 19714 10882 19729 10905
rect 19653 10866 19729 10882
rect 20702 10878 20779 10970
rect 21145 10966 21253 10970
rect 20664 10860 20785 10878
rect 20664 10858 20735 10860
rect 20664 10817 20679 10858
rect 20716 10819 20735 10858
rect 20772 10819 20785 10860
rect 20716 10817 20785 10819
rect 20664 10807 20785 10817
rect 17189 10778 18658 10780
rect 21146 10778 21253 10966
rect 17189 10763 21255 10778
rect 17189 10743 17933 10763
rect 17952 10743 18010 10763
rect 18029 10760 21255 10763
rect 18029 10743 20471 10760
rect 17189 10740 20471 10743
rect 20490 10740 20548 10760
rect 20567 10740 21255 10760
rect 17189 10722 21255 10740
rect 17926 10721 18037 10722
rect 18613 10721 18820 10722
rect 20464 10718 20575 10722
rect 17293 10669 17328 10670
rect 17272 10662 17328 10669
rect 17272 10642 17301 10662
rect 17321 10642 17328 10662
rect 17272 10637 17328 10642
rect 17719 10665 17751 10672
rect 17719 10645 17725 10665
rect 17746 10645 17751 10665
rect 17272 10359 17306 10637
rect 17719 10617 17751 10645
rect 17339 10609 17751 10617
rect 17339 10583 17345 10609
rect 17371 10583 17751 10609
rect 17339 10581 17751 10583
rect 17341 10580 17381 10581
rect 17508 10555 17539 10563
rect 17508 10525 17512 10555
rect 17533 10525 17539 10555
rect 17272 10351 17307 10359
rect 17272 10331 17280 10351
rect 17300 10331 17307 10351
rect 17272 10326 17307 10331
rect 17508 10329 17539 10525
rect 17719 10516 17751 10581
rect 19650 10659 19730 10671
rect 19831 10666 19866 10667
rect 19650 10633 19666 10659
rect 19706 10633 19730 10659
rect 19650 10614 19730 10633
rect 19650 10588 19669 10614
rect 19709 10588 19730 10614
rect 19650 10561 19730 10588
rect 19650 10535 19673 10561
rect 19713 10535 19730 10561
rect 19650 10524 19730 10535
rect 19810 10659 19866 10666
rect 19810 10639 19839 10659
rect 19859 10639 19866 10659
rect 19810 10634 19866 10639
rect 20257 10662 20289 10669
rect 20257 10642 20263 10662
rect 20284 10642 20289 10662
rect 17719 10496 17723 10516
rect 17744 10496 17751 10516
rect 17719 10489 17751 10496
rect 18028 10433 18129 10434
rect 17926 10420 18129 10433
rect 17926 10418 18069 10420
rect 17926 10415 18003 10418
rect 17926 10388 17929 10415
rect 17958 10391 18003 10415
rect 18032 10391 18069 10418
rect 17958 10388 18069 10391
rect 17926 10387 18069 10388
rect 18105 10387 18129 10420
rect 17926 10374 18129 10387
rect 17272 10325 17304 10326
rect 17508 10240 17542 10329
rect 17129 10236 17542 10240
rect 16115 7911 16132 7965
rect 16195 7911 16220 7965
rect 16115 7890 16220 7911
rect 16582 10191 17542 10236
rect 19655 10224 19720 10524
rect 19810 10356 19844 10634
rect 20257 10614 20289 10642
rect 19877 10606 20289 10614
rect 19877 10580 19883 10606
rect 19909 10580 20289 10606
rect 20711 10648 20778 10655
rect 20711 10627 20728 10648
rect 20764 10627 20778 10648
rect 20711 10608 20778 10627
rect 20711 10605 20728 10608
rect 19877 10578 20289 10580
rect 19879 10577 19919 10578
rect 20046 10552 20077 10560
rect 20046 10522 20050 10552
rect 20071 10522 20077 10552
rect 19810 10348 19845 10356
rect 19810 10328 19818 10348
rect 19838 10328 19845 10348
rect 19810 10323 19845 10328
rect 19810 10322 19842 10323
rect 20046 10318 20077 10522
rect 20257 10513 20289 10578
rect 20713 10571 20728 10605
rect 20768 10571 20778 10608
rect 20713 10562 20778 10571
rect 20257 10493 20261 10513
rect 20282 10493 20289 10513
rect 20257 10486 20289 10493
rect 20566 10430 20667 10431
rect 20464 10417 20667 10430
rect 20464 10415 20607 10417
rect 20464 10412 20541 10415
rect 20464 10385 20467 10412
rect 20496 10388 20541 10412
rect 20570 10388 20607 10415
rect 20496 10385 20607 10388
rect 20464 10384 20607 10385
rect 20643 10384 20667 10417
rect 20464 10371 20667 10384
rect 20044 10306 20079 10318
rect 19975 10299 20079 10306
rect 19975 10298 20051 10299
rect 19975 10278 19996 10298
rect 20028 10279 20051 10298
rect 20076 10279 20079 10299
rect 20028 10278 20079 10279
rect 19975 10269 20079 10278
rect 20044 10267 20079 10269
rect 16582 10187 17179 10191
rect 16582 7881 16634 10187
rect 19655 10185 19658 10224
rect 19703 10185 19720 10224
rect 20716 10201 20767 10562
rect 20714 10199 20771 10201
rect 19655 10163 19720 10185
rect 20703 10187 20771 10199
rect 20703 10154 20714 10187
rect 20754 10154 20771 10187
rect 20703 10148 20771 10154
rect 20703 10144 20767 10148
rect 19416 10099 19527 10102
rect 21146 10099 21253 10722
rect 17541 10085 21253 10099
rect 17541 10065 19423 10085
rect 19442 10065 19500 10085
rect 19519 10081 21253 10085
rect 19519 10065 20471 10081
rect 17541 10061 20471 10065
rect 20490 10061 20548 10081
rect 20567 10061 21253 10081
rect 17541 10043 21253 10061
rect 17541 10042 18700 10043
rect 20464 10039 20575 10043
rect 18783 9991 18818 9992
rect 18762 9984 18818 9991
rect 18762 9964 18791 9984
rect 18811 9964 18818 9984
rect 18762 9959 18818 9964
rect 19209 9987 19241 9994
rect 19831 9987 19866 9988
rect 19209 9967 19215 9987
rect 19236 9967 19241 9987
rect 19810 9980 19866 9987
rect 19675 9970 19733 9975
rect 18762 9681 18796 9959
rect 19209 9939 19241 9967
rect 18829 9931 19241 9939
rect 18829 9905 18835 9931
rect 18861 9905 19241 9931
rect 18829 9903 19241 9905
rect 18831 9902 18871 9903
rect 18998 9877 19029 9885
rect 18998 9847 19002 9877
rect 19023 9847 19029 9877
rect 18762 9673 18797 9681
rect 18762 9653 18770 9673
rect 18790 9653 18797 9673
rect 18762 9648 18797 9653
rect 17503 9637 17539 9648
rect 18762 9647 18794 9648
rect 18998 9640 19029 9847
rect 19209 9838 19241 9903
rect 19209 9818 19213 9838
rect 19234 9818 19241 9838
rect 19209 9811 19241 9818
rect 19658 9961 19733 9970
rect 19658 9928 19667 9961
rect 19720 9928 19733 9961
rect 19658 9903 19733 9928
rect 19658 9870 19672 9903
rect 19725 9870 19733 9903
rect 19658 9864 19733 9870
rect 19810 9960 19839 9980
rect 19859 9960 19866 9980
rect 19810 9955 19866 9960
rect 20257 9983 20289 9990
rect 20257 9963 20263 9983
rect 20284 9963 20289 9983
rect 19518 9755 19619 9756
rect 19416 9742 19619 9755
rect 19416 9740 19559 9742
rect 19416 9737 19493 9740
rect 19416 9710 19419 9737
rect 19448 9713 19493 9737
rect 19522 9713 19559 9740
rect 19448 9710 19559 9713
rect 19416 9709 19559 9710
rect 19595 9709 19619 9742
rect 19416 9696 19619 9709
rect 17503 9614 17509 9637
rect 17533 9614 17539 9637
rect 18993 9631 19029 9640
rect 18938 9621 19035 9631
rect 17750 9619 19035 9621
rect 17503 9593 17539 9614
rect 17503 9570 17509 9593
rect 17533 9570 17539 9593
rect 17503 9417 17539 9570
rect 17715 9609 19035 9619
rect 17715 9571 17727 9609
rect 17752 9574 17771 9609
rect 17796 9574 19035 9609
rect 17752 9571 19035 9574
rect 17715 9568 19035 9571
rect 17715 9566 19032 9568
rect 17715 9563 17804 9566
rect 17731 9562 17803 9563
rect 19658 9553 19728 9864
rect 19810 9677 19844 9955
rect 20257 9935 20289 9963
rect 19877 9927 20289 9935
rect 19877 9901 19883 9927
rect 19909 9901 20289 9927
rect 19877 9899 20289 9901
rect 19879 9898 19919 9899
rect 20046 9873 20077 9881
rect 20046 9843 20050 9873
rect 20071 9843 20077 9873
rect 19810 9669 19845 9677
rect 19810 9649 19818 9669
rect 19838 9649 19845 9669
rect 19810 9644 19845 9649
rect 20046 9644 20077 9843
rect 20257 9834 20289 9899
rect 20257 9814 20261 9834
rect 20282 9814 20289 9834
rect 20257 9807 20289 9814
rect 20702 9960 20774 9978
rect 20702 9918 20715 9960
rect 20764 9918 20774 9960
rect 20702 9897 20774 9918
rect 20702 9855 20716 9897
rect 20765 9855 20774 9897
rect 20566 9751 20667 9752
rect 20464 9738 20667 9751
rect 20464 9736 20607 9738
rect 20464 9733 20541 9736
rect 20464 9706 20467 9733
rect 20496 9709 20541 9733
rect 20570 9709 20607 9736
rect 20496 9706 20607 9709
rect 20464 9705 20607 9706
rect 20643 9705 20667 9738
rect 20464 9692 20667 9705
rect 19810 9643 19842 9644
rect 20044 9641 20077 9644
rect 20010 9622 20078 9641
rect 19980 9610 20079 9622
rect 20702 9614 20774 9855
rect 21146 9614 21253 10043
rect 21965 10465 22072 11058
rect 22440 11007 22515 11058
rect 23481 11109 23503 11123
rect 23547 11109 23564 11146
rect 23481 11089 23564 11109
rect 23481 11023 23498 11089
rect 23552 11023 23564 11089
rect 22440 10964 22516 11007
rect 22444 10653 22516 10964
rect 23481 10999 23564 11023
rect 23481 10979 23557 10999
rect 23481 10960 23560 10979
rect 23140 10944 23212 10945
rect 23139 10936 23238 10944
rect 23139 10933 23191 10936
rect 23139 10898 23147 10933
rect 23172 10898 23191 10933
rect 23216 10898 23238 10936
rect 23139 10886 23238 10898
rect 23140 10867 23208 10886
rect 23141 10864 23174 10867
rect 23376 10864 23408 10865
rect 22551 10803 22754 10816
rect 22551 10770 22575 10803
rect 22611 10802 22754 10803
rect 22611 10799 22722 10802
rect 22611 10772 22648 10799
rect 22677 10775 22722 10799
rect 22751 10775 22754 10802
rect 22677 10772 22754 10775
rect 22611 10770 22754 10772
rect 22551 10757 22754 10770
rect 22551 10756 22652 10757
rect 22444 10611 22453 10653
rect 22502 10611 22516 10653
rect 22444 10590 22516 10611
rect 22444 10548 22454 10590
rect 22503 10548 22516 10590
rect 22444 10530 22516 10548
rect 22929 10694 22961 10701
rect 22929 10674 22936 10694
rect 22957 10674 22961 10694
rect 22929 10609 22961 10674
rect 23141 10665 23172 10864
rect 23373 10859 23408 10864
rect 23373 10839 23380 10859
rect 23400 10839 23408 10859
rect 23373 10831 23408 10839
rect 23141 10635 23147 10665
rect 23168 10635 23172 10665
rect 23141 10627 23172 10635
rect 23299 10609 23339 10610
rect 22929 10607 23341 10609
rect 22929 10581 23309 10607
rect 23335 10581 23341 10607
rect 22929 10573 23341 10581
rect 22929 10545 22961 10573
rect 23374 10553 23408 10831
rect 23490 10644 23560 10960
rect 25478 10945 25509 10946
rect 25478 10937 25523 10945
rect 24558 10914 24722 10921
rect 25478 10914 25488 10937
rect 24184 10899 25488 10914
rect 25513 10899 25523 10937
rect 24184 10881 25523 10899
rect 24189 10868 24225 10881
rect 24558 10878 24722 10881
rect 23599 10799 23802 10812
rect 23599 10766 23623 10799
rect 23659 10798 23802 10799
rect 23659 10795 23770 10798
rect 23659 10768 23696 10795
rect 23725 10771 23770 10795
rect 23799 10771 23802 10798
rect 23725 10768 23802 10771
rect 23659 10766 23802 10768
rect 23599 10753 23802 10766
rect 23599 10752 23700 10753
rect 22929 10525 22934 10545
rect 22955 10525 22961 10545
rect 22929 10518 22961 10525
rect 23352 10548 23408 10553
rect 23352 10528 23359 10548
rect 23379 10528 23408 10548
rect 23485 10638 23560 10644
rect 23485 10605 23493 10638
rect 23546 10605 23560 10638
rect 23485 10580 23560 10605
rect 23485 10547 23498 10580
rect 23551 10547 23560 10580
rect 23485 10538 23560 10547
rect 23977 10690 24009 10697
rect 23977 10670 23984 10690
rect 24005 10670 24009 10690
rect 23977 10605 24009 10670
rect 24189 10661 24220 10868
rect 24424 10860 24456 10861
rect 24421 10855 24456 10860
rect 24421 10835 24428 10855
rect 24448 10835 24456 10855
rect 24421 10827 24456 10835
rect 24189 10631 24195 10661
rect 24216 10631 24220 10661
rect 24189 10623 24220 10631
rect 24347 10605 24387 10606
rect 23977 10603 24389 10605
rect 23977 10577 24357 10603
rect 24383 10577 24389 10603
rect 23977 10569 24389 10577
rect 23977 10541 24009 10569
rect 24422 10549 24456 10827
rect 23485 10533 23543 10538
rect 23352 10521 23408 10528
rect 23977 10521 23982 10541
rect 24003 10521 24009 10541
rect 23352 10520 23387 10521
rect 23977 10514 24009 10521
rect 24400 10544 24456 10549
rect 24400 10524 24407 10544
rect 24427 10524 24456 10544
rect 24400 10517 24456 10524
rect 24400 10516 24435 10517
rect 22643 10465 22754 10469
rect 24426 10465 25726 10466
rect 21965 10447 25726 10465
rect 21965 10427 22651 10447
rect 22670 10427 22728 10447
rect 22747 10443 25726 10447
rect 22747 10427 23699 10443
rect 21965 10423 23699 10427
rect 23718 10423 23776 10443
rect 23795 10423 25726 10443
rect 21965 10409 25726 10423
rect 21965 9786 22072 10409
rect 23691 10406 23802 10409
rect 22451 10360 22515 10364
rect 22447 10354 22515 10360
rect 22447 10321 22464 10354
rect 22504 10321 22515 10354
rect 22447 10309 22515 10321
rect 23498 10323 23563 10345
rect 22447 10307 22504 10309
rect 22451 9946 22502 10307
rect 23498 10284 23515 10323
rect 23560 10284 23563 10323
rect 23139 10239 23174 10241
rect 23139 10230 23243 10239
rect 23139 10229 23190 10230
rect 23139 10209 23142 10229
rect 23167 10210 23190 10229
rect 23222 10210 23243 10230
rect 23167 10209 23243 10210
rect 23139 10202 23243 10209
rect 23139 10190 23174 10202
rect 22551 10124 22754 10137
rect 22551 10091 22575 10124
rect 22611 10123 22754 10124
rect 22611 10120 22722 10123
rect 22611 10093 22648 10120
rect 22677 10096 22722 10120
rect 22751 10096 22754 10123
rect 22677 10093 22754 10096
rect 22611 10091 22754 10093
rect 22551 10078 22754 10091
rect 22551 10077 22652 10078
rect 22929 10015 22961 10022
rect 22929 9995 22936 10015
rect 22957 9995 22961 10015
rect 22440 9937 22505 9946
rect 22440 9900 22450 9937
rect 22490 9903 22505 9937
rect 22929 9930 22961 9995
rect 23141 9986 23172 10190
rect 23376 10185 23408 10186
rect 23373 10180 23408 10185
rect 23373 10160 23380 10180
rect 23400 10160 23408 10180
rect 23373 10152 23408 10160
rect 23141 9956 23147 9986
rect 23168 9956 23172 9986
rect 23141 9948 23172 9956
rect 23299 9930 23339 9931
rect 22929 9928 23341 9930
rect 22490 9900 22507 9903
rect 22440 9881 22507 9900
rect 22440 9860 22454 9881
rect 22490 9860 22507 9881
rect 22440 9853 22507 9860
rect 22929 9902 23309 9928
rect 23335 9902 23341 9928
rect 22929 9894 23341 9902
rect 22929 9866 22961 9894
rect 23374 9874 23408 10152
rect 23498 9984 23563 10284
rect 25635 10245 25672 10266
rect 25635 10208 25646 10245
rect 25663 10221 25672 10245
rect 25663 10208 25673 10221
rect 25635 10198 25673 10208
rect 25636 10194 25673 10198
rect 25636 10188 25669 10194
rect 25046 10119 25249 10132
rect 25046 10086 25070 10119
rect 25106 10118 25249 10119
rect 25106 10115 25217 10118
rect 25106 10088 25143 10115
rect 25172 10091 25217 10115
rect 25246 10091 25249 10118
rect 25172 10088 25249 10091
rect 25106 10086 25249 10088
rect 25046 10073 25249 10086
rect 25046 10072 25147 10073
rect 25424 10010 25456 10017
rect 25424 9990 25431 10010
rect 25452 9990 25456 10010
rect 22929 9846 22934 9866
rect 22955 9846 22961 9866
rect 22929 9839 22961 9846
rect 23352 9869 23408 9874
rect 23352 9849 23359 9869
rect 23379 9849 23408 9869
rect 23352 9842 23408 9849
rect 23488 9973 23568 9984
rect 23488 9947 23505 9973
rect 23545 9947 23568 9973
rect 23488 9920 23568 9947
rect 23488 9894 23509 9920
rect 23549 9894 23568 9920
rect 25424 9925 25456 9990
rect 25636 9981 25667 10188
rect 25871 10180 25903 10181
rect 25868 10175 25903 10180
rect 25868 10155 25875 10175
rect 25895 10155 25903 10175
rect 25868 10147 25903 10155
rect 25636 9951 25642 9981
rect 25663 9951 25667 9981
rect 25636 9943 25667 9951
rect 25794 9925 25834 9926
rect 25424 9923 25836 9925
rect 23488 9875 23568 9894
rect 23488 9849 23512 9875
rect 23552 9849 23568 9875
rect 24601 9913 25038 9919
rect 24601 9890 24619 9913
rect 24645 9906 25038 9913
rect 24645 9890 24999 9906
rect 24601 9883 24999 9890
rect 25025 9883 25038 9906
rect 24601 9870 25038 9883
rect 25424 9897 25804 9923
rect 25830 9897 25836 9923
rect 25424 9889 25836 9897
rect 23352 9841 23387 9842
rect 23488 9837 23568 9849
rect 25424 9861 25456 9889
rect 25869 9869 25903 10147
rect 25424 9841 25429 9861
rect 25450 9841 25456 9861
rect 25424 9834 25456 9841
rect 25847 9864 25903 9869
rect 25847 9844 25854 9864
rect 25874 9844 25903 9864
rect 25847 9837 25903 9844
rect 25847 9836 25882 9837
rect 22643 9786 22754 9790
rect 24385 9786 25935 9789
rect 21963 9768 25935 9786
rect 21963 9748 22651 9768
rect 22670 9748 22728 9768
rect 22747 9763 25935 9768
rect 22747 9748 25146 9763
rect 21963 9743 25146 9748
rect 25165 9743 25223 9763
rect 25242 9743 25935 9763
rect 21963 9733 25935 9743
rect 21963 9730 22588 9733
rect 22775 9730 25935 9733
rect 19980 9572 20002 9610
rect 20027 9575 20046 9610
rect 20071 9575 20079 9610
rect 20027 9572 20079 9575
rect 19980 9564 20079 9572
rect 20006 9563 20078 9564
rect 19657 9537 19728 9553
rect 19657 9521 19677 9537
rect 19658 9491 19677 9521
rect 19660 9471 19677 9491
rect 19707 9491 19728 9537
rect 20700 9533 20778 9614
rect 21145 9559 21253 9614
rect 19707 9471 19727 9491
rect 19660 9452 19727 9471
rect 20700 9431 20779 9533
rect 17494 9408 17580 9417
rect 17494 9390 17513 9408
rect 17565 9390 17580 9408
rect 17494 9386 17580 9390
rect 20664 9413 20785 9431
rect 20664 9411 20735 9413
rect 20664 9370 20679 9411
rect 20716 9372 20735 9411
rect 20772 9372 20785 9413
rect 20716 9370 20785 9372
rect 20664 9360 20785 9370
rect 17969 9332 18080 9335
rect 17189 9331 18833 9332
rect 21146 9331 21253 9559
rect 21965 9502 22072 9730
rect 24385 9729 25935 9730
rect 25138 9726 25249 9729
rect 22433 9691 22554 9701
rect 22433 9689 22502 9691
rect 22433 9648 22446 9689
rect 22483 9650 22502 9689
rect 22539 9650 22554 9691
rect 22483 9648 22554 9650
rect 22433 9630 22554 9648
rect 22439 9528 22518 9630
rect 23491 9590 23558 9609
rect 23491 9570 23511 9590
rect 21965 9447 22073 9502
rect 22440 9447 22518 9528
rect 23490 9524 23511 9570
rect 23541 9570 23558 9590
rect 23541 9540 23560 9570
rect 23541 9524 23561 9540
rect 23490 9508 23561 9524
rect 23140 9497 23212 9498
rect 23139 9489 23238 9497
rect 23139 9486 23191 9489
rect 23139 9451 23147 9486
rect 23172 9451 23191 9486
rect 23216 9451 23238 9489
rect 17189 9328 20443 9331
rect 20630 9328 21255 9331
rect 17189 9318 21255 9328
rect 17189 9298 17976 9318
rect 17995 9298 18053 9318
rect 18072 9313 21255 9318
rect 18072 9298 20471 9313
rect 17189 9293 20471 9298
rect 20490 9293 20548 9313
rect 20567 9293 21255 9313
rect 17189 9275 21255 9293
rect 17189 9272 18833 9275
rect 20464 9271 20575 9275
rect 17336 9224 17371 9225
rect 17315 9217 17371 9224
rect 17315 9197 17344 9217
rect 17364 9197 17371 9217
rect 17315 9192 17371 9197
rect 17762 9220 17794 9227
rect 17762 9200 17768 9220
rect 17789 9200 17794 9220
rect 17315 8914 17349 9192
rect 17762 9172 17794 9200
rect 17382 9164 17794 9172
rect 17382 9138 17388 9164
rect 17414 9138 17794 9164
rect 17382 9136 17794 9138
rect 17384 9135 17424 9136
rect 17551 9110 17582 9118
rect 17551 9080 17555 9110
rect 17576 9080 17582 9110
rect 17315 8906 17350 8914
rect 17315 8886 17323 8906
rect 17343 8886 17350 8906
rect 17315 8881 17350 8886
rect 17315 8880 17347 8881
rect 17551 8879 17582 9080
rect 17762 9071 17794 9136
rect 17762 9051 17766 9071
rect 17787 9051 17794 9071
rect 17762 9044 17794 9051
rect 18356 9211 18449 9218
rect 18356 9170 18380 9211
rect 18434 9170 18449 9211
rect 18071 8988 18172 8989
rect 17969 8975 18172 8988
rect 17969 8973 18112 8975
rect 17969 8970 18046 8973
rect 17969 8943 17972 8970
rect 18001 8946 18046 8970
rect 18075 8946 18112 8973
rect 18001 8943 18112 8946
rect 17969 8942 18112 8943
rect 18148 8942 18172 8975
rect 17969 8929 18172 8942
rect 18356 8797 18449 9170
rect 19650 9212 19730 9224
rect 19831 9219 19866 9220
rect 19650 9186 19666 9212
rect 19706 9186 19730 9212
rect 19650 9167 19730 9186
rect 19650 9141 19669 9167
rect 19709 9141 19730 9167
rect 19650 9114 19730 9141
rect 19650 9088 19673 9114
rect 19713 9088 19730 9114
rect 19650 9077 19730 9088
rect 19810 9212 19866 9219
rect 19810 9192 19839 9212
rect 19859 9192 19866 9212
rect 19810 9187 19866 9192
rect 20257 9215 20289 9222
rect 20257 9195 20263 9215
rect 20284 9195 20289 9215
rect 18356 8753 18374 8797
rect 18434 8753 18449 8797
rect 18356 8738 18449 8753
rect 19655 8777 19720 9077
rect 19810 8909 19844 9187
rect 20257 9167 20289 9195
rect 19877 9159 20289 9167
rect 19877 9133 19883 9159
rect 19909 9133 20289 9159
rect 20711 9201 20778 9208
rect 20711 9180 20728 9201
rect 20764 9180 20778 9201
rect 20711 9161 20778 9180
rect 20711 9158 20728 9161
rect 19877 9131 20289 9133
rect 19879 9130 19919 9131
rect 20046 9105 20077 9113
rect 20046 9075 20050 9105
rect 20071 9075 20077 9105
rect 19810 8901 19845 8909
rect 19810 8881 19818 8901
rect 19838 8881 19845 8901
rect 19810 8876 19845 8881
rect 19810 8875 19842 8876
rect 20046 8871 20077 9075
rect 20257 9066 20289 9131
rect 20713 9124 20728 9158
rect 20768 9124 20778 9161
rect 20713 9115 20778 9124
rect 20257 9046 20261 9066
rect 20282 9046 20289 9066
rect 20257 9039 20289 9046
rect 20566 8983 20667 8984
rect 20464 8970 20667 8983
rect 20464 8968 20607 8970
rect 20464 8965 20541 8968
rect 20464 8938 20467 8965
rect 20496 8941 20541 8965
rect 20570 8941 20607 8968
rect 20496 8938 20607 8941
rect 20464 8937 20607 8938
rect 20643 8937 20667 8970
rect 20464 8924 20667 8937
rect 20044 8859 20079 8871
rect 19975 8852 20079 8859
rect 19975 8851 20051 8852
rect 19975 8831 19996 8851
rect 20028 8832 20051 8851
rect 20076 8832 20079 8852
rect 20028 8831 20079 8832
rect 19975 8822 20079 8831
rect 20044 8820 20079 8822
rect 19655 8738 19658 8777
rect 19703 8738 19720 8777
rect 20716 8754 20767 9115
rect 20714 8752 20771 8754
rect 19655 8716 19720 8738
rect 20703 8740 20771 8752
rect 20703 8707 20714 8740
rect 20754 8707 20771 8740
rect 20703 8701 20771 8707
rect 20703 8697 20767 8701
rect 19416 8652 19527 8655
rect 21146 8652 21253 9275
rect 17222 8638 21253 8652
rect 17222 8618 19423 8638
rect 19442 8618 19500 8638
rect 19519 8634 21253 8638
rect 19519 8618 20471 8634
rect 17222 8614 20471 8618
rect 20490 8614 20548 8634
rect 20567 8614 21253 8634
rect 17222 8596 21253 8614
rect 17222 8595 18792 8596
rect 20464 8592 20575 8596
rect 18783 8544 18818 8545
rect 18762 8537 18818 8544
rect 18762 8517 18791 8537
rect 18811 8517 18818 8537
rect 18762 8512 18818 8517
rect 19209 8540 19241 8547
rect 19831 8540 19866 8541
rect 19209 8520 19215 8540
rect 19236 8520 19241 8540
rect 19810 8533 19866 8540
rect 19675 8523 19733 8528
rect 18362 8457 18444 8486
rect 18362 8416 18387 8457
rect 18423 8416 18444 8457
rect 18549 8477 18613 8496
rect 18549 8438 18566 8477
rect 18600 8438 18613 8477
rect 18549 8419 18613 8438
rect 18362 8101 18444 8416
rect 18354 8056 18444 8101
rect 18551 8074 18613 8419
rect 18762 8234 18796 8512
rect 19209 8492 19241 8520
rect 18829 8484 19241 8492
rect 18829 8458 18835 8484
rect 18861 8458 19241 8484
rect 18829 8456 19241 8458
rect 18831 8455 18871 8456
rect 18998 8430 19029 8438
rect 18998 8400 19002 8430
rect 19023 8400 19029 8430
rect 18762 8226 18797 8234
rect 18762 8206 18770 8226
rect 18790 8206 18797 8226
rect 18762 8201 18797 8206
rect 18762 8200 18794 8201
rect 18998 8193 19029 8400
rect 19209 8391 19241 8456
rect 19209 8371 19213 8391
rect 19234 8371 19241 8391
rect 19209 8364 19241 8371
rect 19658 8514 19733 8523
rect 19658 8481 19667 8514
rect 19720 8481 19733 8514
rect 19658 8456 19733 8481
rect 19658 8423 19672 8456
rect 19725 8423 19733 8456
rect 19658 8417 19733 8423
rect 19810 8513 19839 8533
rect 19859 8513 19866 8533
rect 19810 8508 19866 8513
rect 20257 8536 20289 8543
rect 20257 8516 20263 8536
rect 20284 8516 20289 8536
rect 19518 8308 19619 8309
rect 19416 8295 19619 8308
rect 19416 8293 19559 8295
rect 19416 8290 19493 8293
rect 19416 8263 19419 8290
rect 19448 8266 19493 8290
rect 19522 8266 19559 8293
rect 19448 8263 19559 8266
rect 19416 8262 19559 8263
rect 19595 8262 19619 8295
rect 19416 8249 19619 8262
rect 18993 8175 19029 8193
rect 18960 8174 19029 8175
rect 18940 8162 19029 8174
rect 18940 8124 18952 8162
rect 18977 8127 18996 8162
rect 19021 8127 19029 8162
rect 19658 8151 19728 8417
rect 19810 8230 19844 8508
rect 20257 8488 20289 8516
rect 19877 8480 20289 8488
rect 19877 8454 19883 8480
rect 19909 8454 20289 8480
rect 19877 8452 20289 8454
rect 19879 8451 19919 8452
rect 20046 8426 20077 8434
rect 20046 8396 20050 8426
rect 20071 8396 20077 8426
rect 19810 8222 19845 8230
rect 19810 8202 19818 8222
rect 19838 8202 19845 8222
rect 19810 8197 19845 8202
rect 20046 8197 20077 8396
rect 20257 8387 20289 8452
rect 20257 8367 20261 8387
rect 20282 8367 20289 8387
rect 20257 8360 20289 8367
rect 20702 8513 20774 8531
rect 20702 8471 20715 8513
rect 20764 8471 20774 8513
rect 20702 8450 20774 8471
rect 20702 8408 20716 8450
rect 20765 8408 20774 8450
rect 20566 8304 20667 8305
rect 20464 8291 20667 8304
rect 20464 8289 20607 8291
rect 20464 8286 20541 8289
rect 20464 8259 20467 8286
rect 20496 8262 20541 8286
rect 20570 8262 20607 8289
rect 20496 8259 20607 8262
rect 20464 8258 20607 8259
rect 20643 8258 20667 8291
rect 20464 8245 20667 8258
rect 19810 8196 19842 8197
rect 20044 8194 20077 8197
rect 20010 8175 20078 8194
rect 18977 8124 19029 8127
rect 18940 8116 19029 8124
rect 19649 8122 19728 8151
rect 19980 8163 20079 8175
rect 19980 8125 20002 8163
rect 20027 8128 20046 8163
rect 20071 8128 20079 8163
rect 20027 8125 20079 8128
rect 18956 8115 19028 8116
rect 18550 8065 18624 8074
rect 18354 8023 18438 8056
rect 18354 7995 18369 8023
rect 18413 7995 18438 8023
rect 18354 7966 18438 7995
rect 18550 8017 18564 8065
rect 18601 8017 18624 8065
rect 18550 7989 18624 8017
rect 18354 7938 18366 7966
rect 18410 7938 18438 7966
rect 18354 7927 18438 7938
rect 19649 7939 19726 8122
rect 19980 8117 20079 8125
rect 20006 8116 20078 8117
rect 20702 8114 20774 8408
rect 21146 8136 21253 8596
rect 21965 9018 22072 9447
rect 22444 9206 22516 9447
rect 23139 9439 23238 9451
rect 23140 9420 23208 9439
rect 23141 9417 23174 9420
rect 23376 9417 23408 9418
rect 22551 9356 22754 9369
rect 22551 9323 22575 9356
rect 22611 9355 22754 9356
rect 22611 9352 22722 9355
rect 22611 9325 22648 9352
rect 22677 9328 22722 9352
rect 22751 9328 22754 9355
rect 22677 9325 22754 9328
rect 22611 9323 22754 9325
rect 22551 9310 22754 9323
rect 22551 9309 22652 9310
rect 22444 9164 22453 9206
rect 22502 9164 22516 9206
rect 22444 9143 22516 9164
rect 22444 9101 22454 9143
rect 22503 9101 22516 9143
rect 22444 9083 22516 9101
rect 22929 9247 22961 9254
rect 22929 9227 22936 9247
rect 22957 9227 22961 9247
rect 22929 9162 22961 9227
rect 23141 9218 23172 9417
rect 23373 9412 23408 9417
rect 23373 9392 23380 9412
rect 23400 9392 23408 9412
rect 23373 9384 23408 9392
rect 23141 9188 23147 9218
rect 23168 9188 23172 9218
rect 23141 9180 23172 9188
rect 23299 9162 23339 9163
rect 22929 9160 23341 9162
rect 22929 9134 23309 9160
rect 23335 9134 23341 9160
rect 22929 9126 23341 9134
rect 22929 9098 22961 9126
rect 23374 9106 23408 9384
rect 23490 9197 23560 9508
rect 24187 9499 25529 9504
rect 24187 9497 25486 9499
rect 24184 9471 25486 9497
rect 25514 9471 25529 9499
rect 24184 9463 25529 9471
rect 24184 9438 24223 9463
rect 24184 9421 24225 9438
rect 24184 9414 24223 9421
rect 23599 9352 23802 9365
rect 23599 9319 23623 9352
rect 23659 9351 23802 9352
rect 23659 9348 23770 9351
rect 23659 9321 23696 9348
rect 23725 9324 23770 9348
rect 23799 9324 23802 9351
rect 23725 9321 23802 9324
rect 23659 9319 23802 9321
rect 23599 9306 23802 9319
rect 23599 9305 23700 9306
rect 22929 9078 22934 9098
rect 22955 9078 22961 9098
rect 22929 9071 22961 9078
rect 23352 9101 23408 9106
rect 23352 9081 23359 9101
rect 23379 9081 23408 9101
rect 23485 9191 23560 9197
rect 23485 9158 23493 9191
rect 23546 9158 23560 9191
rect 23485 9133 23560 9158
rect 23485 9100 23498 9133
rect 23551 9100 23560 9133
rect 23485 9091 23560 9100
rect 23977 9243 24009 9250
rect 23977 9223 23984 9243
rect 24005 9223 24009 9243
rect 23977 9158 24009 9223
rect 24189 9214 24220 9414
rect 24424 9413 24456 9414
rect 24421 9408 24456 9413
rect 24421 9388 24428 9408
rect 24448 9388 24456 9408
rect 24421 9380 24456 9388
rect 24189 9184 24195 9214
rect 24216 9184 24220 9214
rect 24189 9176 24220 9184
rect 24347 9158 24387 9159
rect 23977 9156 24389 9158
rect 23977 9130 24357 9156
rect 24383 9130 24389 9156
rect 23977 9122 24389 9130
rect 23977 9094 24009 9122
rect 24422 9102 24456 9380
rect 23485 9086 23543 9091
rect 23352 9074 23408 9081
rect 23977 9074 23982 9094
rect 24003 9074 24009 9094
rect 23352 9073 23387 9074
rect 23977 9067 24009 9074
rect 24400 9097 24456 9102
rect 24400 9077 24407 9097
rect 24427 9077 24456 9097
rect 24400 9070 24456 9077
rect 24400 9069 24435 9070
rect 22643 9018 22754 9022
rect 24518 9018 24961 9019
rect 21965 9000 24961 9018
rect 21965 8980 22651 9000
rect 22670 8980 22728 9000
rect 22747 8996 24961 9000
rect 22747 8980 23699 8996
rect 21965 8976 23699 8980
rect 23718 8976 23776 8996
rect 23795 8976 24961 8996
rect 21965 8962 24961 8976
rect 21965 8339 22072 8962
rect 23691 8959 23802 8962
rect 22451 8913 22515 8917
rect 22447 8907 22515 8913
rect 22447 8874 22464 8907
rect 22504 8874 22515 8907
rect 22447 8862 22515 8874
rect 23498 8876 23563 8898
rect 22447 8860 22504 8862
rect 22451 8499 22502 8860
rect 23498 8837 23515 8876
rect 23560 8837 23563 8876
rect 23139 8792 23174 8794
rect 23139 8783 23243 8792
rect 23139 8782 23190 8783
rect 23139 8762 23142 8782
rect 23167 8763 23190 8782
rect 23222 8763 23243 8783
rect 23167 8762 23243 8763
rect 23139 8755 23243 8762
rect 23139 8743 23174 8755
rect 22551 8677 22754 8690
rect 22551 8644 22575 8677
rect 22611 8676 22754 8677
rect 22611 8673 22722 8676
rect 22611 8646 22648 8673
rect 22677 8649 22722 8673
rect 22751 8649 22754 8676
rect 22677 8646 22754 8649
rect 22611 8644 22754 8646
rect 22551 8631 22754 8644
rect 22551 8630 22652 8631
rect 22929 8568 22961 8575
rect 22929 8548 22936 8568
rect 22957 8548 22961 8568
rect 22440 8490 22505 8499
rect 22440 8453 22450 8490
rect 22490 8456 22505 8490
rect 22929 8483 22961 8548
rect 23141 8539 23172 8743
rect 23376 8738 23408 8739
rect 23373 8733 23408 8738
rect 23373 8713 23380 8733
rect 23400 8713 23408 8733
rect 23373 8705 23408 8713
rect 23141 8509 23147 8539
rect 23168 8509 23172 8539
rect 23141 8501 23172 8509
rect 23299 8483 23339 8484
rect 22929 8481 23341 8483
rect 22490 8453 22507 8456
rect 22440 8434 22507 8453
rect 22440 8413 22454 8434
rect 22490 8413 22507 8434
rect 22440 8406 22507 8413
rect 22929 8455 23309 8481
rect 23335 8455 23341 8481
rect 22929 8447 23341 8455
rect 22929 8419 22961 8447
rect 23374 8427 23408 8705
rect 23498 8537 23563 8837
rect 22929 8399 22934 8419
rect 22955 8399 22961 8419
rect 22929 8392 22961 8399
rect 23352 8422 23408 8427
rect 23352 8402 23359 8422
rect 23379 8402 23408 8422
rect 23352 8395 23408 8402
rect 23488 8526 23568 8537
rect 23488 8500 23505 8526
rect 23545 8500 23568 8526
rect 23488 8473 23568 8500
rect 26040 8476 26089 13662
rect 26537 13659 26695 13662
rect 26557 13651 26695 13659
rect 27077 13104 27185 14234
rect 37796 14231 37816 14283
rect 37894 14231 37907 14289
rect 37796 14218 37907 14231
rect 36739 14150 36826 14168
rect 36739 14106 36756 14150
rect 36808 14106 36826 14150
rect 36739 14089 36826 14106
rect 35481 14046 35562 14047
rect 35475 14032 35574 14046
rect 35475 13982 35495 14032
rect 35547 13982 35574 14032
rect 35475 13962 35574 13982
rect 31678 13849 31743 13932
rect 31628 13831 31749 13849
rect 31628 13829 31699 13831
rect 31628 13788 31643 13829
rect 31680 13790 31699 13829
rect 31736 13790 31749 13831
rect 31680 13788 31749 13790
rect 31628 13778 31749 13788
rect 32109 13749 32786 13773
rect 29633 13744 31304 13749
rect 31562 13744 32786 13749
rect 29633 13731 32786 13744
rect 29633 13711 31435 13731
rect 31454 13711 31512 13731
rect 31531 13711 32786 13731
rect 29633 13693 32786 13711
rect 29633 13692 29784 13693
rect 31428 13689 31539 13693
rect 32109 13685 32786 13693
rect 30614 13630 30694 13642
rect 30795 13637 30830 13638
rect 30614 13604 30630 13630
rect 30670 13604 30694 13630
rect 30614 13585 30694 13604
rect 30614 13559 30633 13585
rect 30673 13559 30694 13585
rect 30614 13532 30694 13559
rect 30614 13506 30637 13532
rect 30677 13506 30694 13532
rect 30614 13495 30694 13506
rect 30774 13630 30830 13637
rect 30774 13610 30803 13630
rect 30823 13610 30830 13630
rect 30774 13605 30830 13610
rect 31221 13633 31253 13640
rect 31221 13613 31227 13633
rect 31248 13613 31253 13633
rect 30619 13195 30684 13495
rect 30774 13327 30808 13605
rect 31221 13585 31253 13613
rect 30841 13577 31253 13585
rect 30841 13551 30847 13577
rect 30873 13551 31253 13577
rect 31675 13619 31742 13626
rect 31675 13598 31692 13619
rect 31728 13598 31742 13619
rect 31675 13579 31742 13598
rect 31675 13576 31692 13579
rect 30841 13549 31253 13551
rect 30843 13548 30883 13549
rect 31010 13523 31041 13531
rect 31010 13493 31014 13523
rect 31035 13493 31041 13523
rect 30774 13319 30809 13327
rect 30774 13299 30782 13319
rect 30802 13299 30809 13319
rect 30774 13294 30809 13299
rect 30774 13293 30806 13294
rect 31010 13289 31041 13493
rect 31221 13484 31253 13549
rect 31677 13542 31692 13576
rect 31732 13542 31742 13579
rect 31677 13533 31742 13542
rect 31221 13464 31225 13484
rect 31246 13464 31253 13484
rect 31221 13457 31253 13464
rect 31530 13401 31631 13402
rect 31428 13388 31631 13401
rect 31428 13386 31571 13388
rect 31428 13383 31505 13386
rect 31428 13356 31431 13383
rect 31460 13359 31505 13383
rect 31534 13359 31571 13386
rect 31460 13356 31571 13359
rect 31428 13355 31571 13356
rect 31607 13355 31631 13388
rect 31428 13342 31631 13355
rect 31008 13277 31043 13289
rect 30939 13270 31043 13277
rect 30939 13269 31015 13270
rect 30939 13249 30960 13269
rect 30992 13250 31015 13269
rect 31040 13250 31043 13270
rect 30992 13249 31043 13250
rect 30939 13240 31043 13249
rect 31008 13238 31043 13240
rect 30619 13156 30622 13195
rect 30667 13156 30684 13195
rect 31680 13172 31731 13533
rect 31678 13170 31735 13172
rect 30619 13134 30684 13156
rect 31667 13158 31735 13170
rect 31667 13125 31678 13158
rect 31718 13125 31735 13158
rect 31667 13119 31735 13125
rect 31667 13115 31731 13119
rect 26154 8668 26357 8681
rect 26154 8635 26178 8668
rect 26214 8667 26357 8668
rect 26214 8664 26325 8667
rect 26214 8637 26251 8664
rect 26280 8640 26325 8664
rect 26354 8640 26357 8667
rect 26280 8637 26357 8640
rect 26214 8635 26357 8637
rect 26154 8622 26357 8635
rect 26154 8621 26255 8622
rect 26532 8559 26564 8566
rect 26532 8539 26539 8559
rect 26560 8539 26564 8559
rect 23488 8447 23509 8473
rect 23549 8447 23568 8473
rect 23488 8428 23568 8447
rect 26039 8466 26150 8476
rect 26039 8465 26104 8466
rect 26039 8441 26047 8465
rect 26071 8442 26104 8465
rect 26128 8442 26150 8466
rect 26071 8441 26150 8442
rect 26039 8434 26150 8441
rect 26532 8474 26564 8539
rect 26744 8530 26775 8730
rect 26979 8729 27011 8730
rect 26976 8724 27011 8729
rect 26976 8704 26983 8724
rect 27003 8704 27011 8724
rect 26976 8696 27011 8704
rect 26744 8500 26750 8530
rect 26771 8500 26775 8530
rect 26744 8492 26775 8500
rect 26902 8474 26942 8475
rect 26532 8472 26944 8474
rect 26532 8446 26912 8472
rect 26938 8446 26944 8472
rect 26532 8438 26944 8446
rect 23488 8402 23512 8428
rect 23552 8402 23568 8428
rect 23352 8394 23387 8395
rect 23488 8390 23568 8402
rect 26532 8410 26564 8438
rect 26977 8418 27011 8696
rect 26532 8390 26537 8410
rect 26558 8390 26564 8410
rect 26532 8383 26564 8390
rect 26743 8410 26777 8417
rect 26743 8388 26750 8410
rect 26774 8388 26777 8410
rect 22643 8339 22754 8343
rect 24398 8339 24605 8340
rect 21963 8334 26038 8339
rect 21963 8321 26357 8334
rect 21963 8301 22651 8321
rect 22670 8301 22728 8321
rect 22747 8312 26357 8321
rect 22747 8301 26254 8312
rect 21963 8292 26254 8301
rect 26273 8292 26331 8312
rect 26350 8292 26357 8312
rect 21963 8283 26357 8292
rect 20702 8076 20778 8114
rect 21146 8076 21259 8136
rect 21965 8110 22072 8283
rect 24560 8281 26357 8283
rect 26246 8275 26357 8281
rect 22433 8244 22554 8254
rect 22433 8242 22502 8244
rect 22433 8201 22446 8242
rect 22483 8203 22502 8242
rect 22539 8203 22554 8244
rect 22483 8201 22554 8203
rect 22433 8183 22554 8201
rect 26581 8233 26633 8264
rect 26581 8199 26590 8233
rect 26619 8199 26633 8233
rect 20713 7975 20778 8076
rect 19649 7896 19666 7939
rect 16582 7847 16597 7881
rect 16626 7847 16634 7881
rect 19654 7891 19666 7896
rect 19712 7891 19726 7939
rect 19654 7869 19726 7891
rect 20711 7929 20778 7975
rect 21148 7937 21259 8076
rect 16582 7821 16634 7847
rect 20711 7837 20776 7929
rect 21143 7910 21259 7937
rect 21956 8083 22072 8110
rect 22439 8091 22504 8183
rect 26581 8173 26633 8199
rect 26743 8182 26777 8388
rect 26955 8413 27011 8418
rect 26955 8393 26962 8413
rect 26982 8393 27011 8413
rect 26955 8386 27011 8393
rect 26955 8385 26990 8386
rect 21956 7944 22067 8083
rect 22437 8045 22504 8091
rect 23489 8129 23561 8151
rect 23489 8081 23503 8129
rect 23549 8124 23561 8129
rect 26581 8139 26589 8173
rect 26618 8139 26633 8173
rect 23549 8081 23566 8124
rect 22437 7944 22502 8045
rect 16582 7787 16596 7821
rect 16625 7787 16634 7821
rect 16582 7756 16634 7787
rect 20661 7819 20782 7837
rect 20661 7817 20732 7819
rect 20661 7776 20676 7817
rect 20713 7778 20732 7817
rect 20769 7778 20782 7819
rect 20713 7776 20782 7778
rect 20661 7766 20782 7776
rect 16858 7739 16969 7745
rect 16858 7737 18655 7739
rect 21143 7737 21250 7910
rect 21956 7884 22069 7944
rect 22437 7906 22513 7944
rect 16858 7728 21252 7737
rect 16858 7708 16865 7728
rect 16884 7708 16942 7728
rect 16961 7719 21252 7728
rect 16961 7708 20468 7719
rect 16858 7699 20468 7708
rect 20487 7699 20545 7719
rect 20564 7699 21252 7719
rect 16858 7686 21252 7699
rect 17177 7681 21252 7686
rect 18610 7680 18817 7681
rect 20461 7677 20572 7681
rect 16225 7634 16260 7635
rect 16204 7627 16260 7634
rect 16204 7607 16233 7627
rect 16253 7607 16260 7627
rect 16204 7602 16260 7607
rect 16651 7630 16683 7637
rect 16651 7610 16657 7630
rect 16678 7610 16683 7630
rect 16204 7324 16238 7602
rect 16651 7582 16683 7610
rect 19647 7618 19727 7630
rect 19828 7625 19863 7626
rect 19647 7592 19663 7618
rect 19703 7592 19727 7618
rect 16271 7574 16683 7582
rect 16271 7548 16277 7574
rect 16303 7548 16683 7574
rect 16271 7546 16683 7548
rect 16273 7545 16313 7546
rect 16440 7520 16471 7528
rect 16440 7490 16444 7520
rect 16465 7490 16471 7520
rect 16204 7316 16239 7324
rect 16204 7296 16212 7316
rect 16232 7296 16239 7316
rect 16440 7305 16471 7490
rect 16651 7481 16683 7546
rect 17065 7579 17176 7586
rect 17065 7578 17144 7579
rect 17065 7554 17087 7578
rect 17111 7555 17144 7578
rect 17168 7555 17176 7579
rect 17111 7554 17176 7555
rect 17065 7544 17176 7554
rect 19647 7573 19727 7592
rect 19647 7547 19666 7573
rect 19706 7547 19727 7573
rect 17126 7527 17175 7544
rect 19647 7520 19727 7547
rect 19647 7494 19670 7520
rect 19710 7494 19727 7520
rect 19647 7483 19727 7494
rect 19807 7618 19863 7625
rect 19807 7598 19836 7618
rect 19856 7598 19863 7618
rect 19807 7593 19863 7598
rect 20254 7621 20286 7628
rect 20254 7601 20260 7621
rect 20281 7601 20286 7621
rect 16651 7461 16655 7481
rect 16676 7461 16683 7481
rect 16651 7454 16683 7461
rect 16960 7398 17061 7399
rect 16858 7385 17061 7398
rect 16858 7383 17001 7385
rect 16858 7380 16935 7383
rect 16858 7353 16861 7380
rect 16890 7356 16935 7380
rect 16964 7356 17001 7383
rect 16890 7353 17001 7356
rect 16858 7352 17001 7353
rect 17037 7352 17061 7385
rect 16858 7339 17061 7352
rect 16204 7291 16239 7296
rect 16204 7290 16236 7291
rect 16438 7228 16472 7305
rect 15071 5825 15668 5829
rect 12171 5747 12206 5749
rect 12171 5738 12275 5747
rect 12171 5737 12222 5738
rect 12171 5717 12174 5737
rect 12199 5718 12222 5737
rect 12254 5718 12275 5738
rect 12199 5717 12275 5718
rect 12171 5710 12275 5717
rect 12171 5698 12206 5710
rect 11583 5632 11786 5645
rect 11583 5599 11607 5632
rect 11643 5631 11786 5632
rect 11643 5628 11754 5631
rect 11643 5601 11680 5628
rect 11709 5604 11754 5628
rect 11783 5604 11786 5631
rect 11709 5601 11786 5604
rect 11643 5599 11786 5601
rect 11583 5586 11786 5599
rect 11583 5585 11684 5586
rect 11961 5523 11993 5530
rect 11961 5503 11968 5523
rect 11989 5503 11993 5523
rect 11472 5445 11537 5454
rect 11472 5408 11482 5445
rect 11522 5411 11537 5445
rect 11961 5438 11993 5503
rect 12173 5494 12204 5698
rect 12408 5693 12440 5694
rect 12405 5688 12440 5693
rect 12405 5668 12412 5688
rect 12432 5668 12440 5688
rect 12405 5660 12440 5668
rect 12173 5464 12179 5494
rect 12200 5464 12204 5494
rect 12173 5456 12204 5464
rect 12331 5438 12371 5439
rect 11961 5436 12373 5438
rect 11522 5408 11539 5411
rect 11472 5389 11539 5408
rect 11472 5368 11486 5389
rect 11522 5368 11539 5389
rect 11472 5361 11539 5368
rect 11961 5410 12341 5436
rect 12367 5410 12373 5436
rect 11961 5402 12373 5410
rect 11961 5374 11993 5402
rect 12406 5382 12440 5660
rect 12530 5492 12595 5792
rect 14708 5780 15668 5825
rect 15775 6168 15811 6796
rect 14708 5776 15121 5780
rect 14708 5687 14742 5776
rect 14946 5690 14978 5691
rect 14121 5629 14324 5642
rect 14121 5596 14145 5629
rect 14181 5628 14324 5629
rect 14181 5625 14292 5628
rect 14181 5598 14218 5625
rect 14247 5601 14292 5625
rect 14321 5601 14324 5628
rect 14247 5598 14324 5601
rect 14181 5596 14324 5598
rect 14121 5583 14324 5596
rect 14121 5582 14222 5583
rect 14499 5520 14531 5527
rect 14499 5500 14506 5520
rect 14527 5500 14531 5520
rect 11961 5354 11966 5374
rect 11987 5354 11993 5374
rect 11961 5347 11993 5354
rect 12384 5377 12440 5382
rect 12384 5357 12391 5377
rect 12411 5357 12440 5377
rect 12384 5350 12440 5357
rect 12520 5481 12600 5492
rect 12520 5455 12537 5481
rect 12577 5455 12600 5481
rect 12520 5428 12600 5455
rect 12520 5402 12541 5428
rect 12581 5402 12600 5428
rect 12520 5383 12600 5402
rect 12520 5357 12544 5383
rect 12584 5357 12600 5383
rect 12384 5349 12419 5350
rect 12520 5345 12600 5357
rect 14499 5435 14531 5500
rect 14711 5491 14742 5687
rect 14943 5685 14978 5690
rect 14943 5665 14950 5685
rect 14970 5665 14978 5685
rect 14943 5657 14978 5665
rect 14711 5461 14717 5491
rect 14738 5461 14742 5491
rect 14711 5453 14742 5461
rect 14869 5435 14909 5436
rect 14499 5433 14911 5435
rect 14499 5407 14879 5433
rect 14905 5407 14911 5433
rect 14499 5399 14911 5407
rect 14499 5371 14531 5399
rect 14944 5379 14978 5657
rect 14499 5351 14504 5371
rect 14525 5351 14531 5371
rect 14499 5344 14531 5351
rect 14922 5374 14978 5379
rect 14922 5354 14929 5374
rect 14949 5354 14978 5374
rect 14922 5347 14978 5354
rect 14922 5346 14957 5347
rect 11675 5294 11786 5298
rect 13430 5294 13637 5295
rect 14213 5294 14324 5295
rect 10995 5276 15061 5294
rect 10995 5256 11683 5276
rect 11702 5256 11760 5276
rect 11779 5273 15061 5276
rect 11779 5256 14221 5273
rect 10995 5253 14221 5256
rect 14240 5253 14298 5273
rect 14317 5253 15061 5273
rect 10995 5238 15061 5253
rect 10997 5050 11104 5238
rect 13592 5236 15061 5238
rect 11465 5199 11586 5209
rect 11465 5197 11534 5199
rect 11465 5156 11478 5197
rect 11515 5158 11534 5197
rect 11571 5158 11586 5199
rect 11515 5156 11586 5158
rect 11465 5138 11586 5156
rect 10997 5046 11105 5050
rect 11471 5046 11548 5138
rect 12521 5134 12597 5150
rect 12521 5111 12536 5134
rect 9004 4880 9019 4903
rect 8943 4864 9019 4880
rect 9992 4876 10069 4968
rect 10435 4964 10543 4968
rect 9954 4858 10075 4876
rect 9954 4856 10025 4858
rect 9954 4815 9969 4856
rect 10006 4817 10025 4856
rect 10062 4817 10075 4858
rect 10006 4815 10075 4817
rect 9954 4805 10075 4815
rect 6525 4776 7948 4778
rect 10436 4776 10543 4964
rect 6525 4761 10545 4776
rect 6525 4741 7223 4761
rect 7242 4741 7300 4761
rect 7319 4758 10545 4761
rect 7319 4741 9761 4758
rect 6525 4738 9761 4741
rect 9780 4738 9838 4758
rect 9857 4738 10545 4758
rect 6525 4720 10545 4738
rect 7216 4719 7327 4720
rect 7903 4719 8110 4720
rect 9754 4716 9865 4720
rect 6583 4667 6618 4668
rect 6562 4660 6618 4667
rect 6562 4640 6591 4660
rect 6611 4640 6618 4660
rect 6562 4635 6618 4640
rect 7009 4663 7041 4670
rect 7009 4643 7015 4663
rect 7036 4643 7041 4663
rect 5731 4411 5757 4426
rect 5728 4404 5764 4411
rect 5728 4366 5734 4404
rect 5757 4366 5764 4404
rect 5728 4360 5764 4366
rect 6562 4357 6596 4635
rect 7009 4615 7041 4643
rect 6629 4607 7041 4615
rect 6629 4581 6635 4607
rect 6661 4581 7041 4607
rect 6629 4579 7041 4581
rect 6631 4578 6671 4579
rect 6798 4553 6829 4561
rect 6798 4523 6802 4553
rect 6823 4523 6829 4553
rect 6562 4349 6597 4357
rect 6562 4329 6570 4349
rect 6590 4329 6597 4349
rect 6562 4324 6597 4329
rect 6562 4323 6594 4324
rect 6798 4320 6829 4523
rect 7009 4514 7041 4579
rect 8940 4657 9020 4669
rect 9121 4664 9156 4665
rect 8940 4631 8956 4657
rect 8996 4631 9020 4657
rect 8940 4612 9020 4631
rect 8940 4586 8959 4612
rect 8999 4586 9020 4612
rect 8940 4559 9020 4586
rect 8940 4533 8963 4559
rect 9003 4533 9020 4559
rect 8940 4522 9020 4533
rect 9100 4657 9156 4664
rect 9100 4637 9129 4657
rect 9149 4637 9156 4657
rect 9100 4632 9156 4637
rect 9547 4660 9579 4667
rect 9547 4640 9553 4660
rect 9574 4640 9579 4660
rect 7009 4494 7013 4514
rect 7034 4494 7041 4514
rect 7009 4487 7041 4494
rect 7318 4431 7419 4432
rect 7216 4418 7419 4431
rect 7216 4416 7359 4418
rect 7216 4413 7293 4416
rect 7216 4386 7219 4413
rect 7248 4389 7293 4413
rect 7322 4389 7359 4416
rect 7248 4386 7359 4389
rect 7216 4385 7359 4386
rect 7395 4385 7419 4418
rect 7216 4372 7419 4385
rect 6793 4302 6829 4320
rect 6793 4285 6828 4302
rect 6726 4254 6831 4285
rect 6726 4249 6798 4254
rect 6726 4228 6757 4249
rect 6777 4233 6798 4249
rect 6818 4233 6831 4254
rect 6777 4228 6831 4233
rect 6726 4219 6831 4228
rect 8945 4222 9010 4522
rect 9100 4354 9134 4632
rect 9547 4612 9579 4640
rect 9167 4604 9579 4612
rect 9167 4578 9173 4604
rect 9199 4578 9579 4604
rect 10001 4646 10068 4653
rect 10001 4625 10018 4646
rect 10054 4625 10068 4646
rect 10001 4606 10068 4625
rect 10001 4603 10018 4606
rect 9167 4576 9579 4578
rect 9169 4575 9209 4576
rect 9336 4550 9367 4558
rect 9336 4520 9340 4550
rect 9361 4520 9367 4550
rect 9100 4346 9135 4354
rect 9100 4326 9108 4346
rect 9128 4326 9135 4346
rect 9100 4321 9135 4326
rect 9100 4320 9132 4321
rect 9336 4316 9367 4520
rect 9547 4511 9579 4576
rect 10003 4569 10018 4603
rect 10058 4569 10068 4606
rect 10003 4560 10068 4569
rect 9547 4491 9551 4511
rect 9572 4491 9579 4511
rect 9547 4484 9579 4491
rect 9856 4428 9957 4429
rect 9754 4415 9957 4428
rect 9754 4413 9897 4415
rect 9754 4410 9831 4413
rect 9754 4383 9757 4410
rect 9786 4386 9831 4410
rect 9860 4386 9897 4413
rect 9786 4383 9897 4386
rect 9754 4382 9897 4383
rect 9933 4382 9957 4415
rect 9754 4369 9957 4382
rect 9334 4304 9369 4316
rect 9265 4297 9369 4304
rect 9265 4296 9341 4297
rect 9265 4276 9286 4296
rect 9318 4277 9341 4296
rect 9366 4277 9369 4297
rect 9318 4276 9369 4277
rect 9265 4267 9369 4276
rect 9334 4265 9369 4267
rect 8945 4183 8948 4222
rect 8993 4183 9010 4222
rect 10006 4199 10057 4560
rect 10004 4197 10061 4199
rect 8945 4161 9010 4183
rect 9993 4185 10061 4197
rect 9993 4152 10004 4185
rect 10044 4152 10061 4185
rect 9993 4146 10061 4152
rect 9993 4142 10057 4146
rect 8706 4097 8817 4100
rect 10436 4097 10543 4720
rect 6749 4083 10543 4097
rect 6749 4063 8713 4083
rect 8732 4063 8790 4083
rect 8809 4079 10543 4083
rect 8809 4063 9761 4079
rect 6749 4059 9761 4063
rect 9780 4059 9838 4079
rect 9857 4059 10543 4079
rect 6749 4041 10543 4059
rect 6749 4040 7990 4041
rect 9754 4037 9865 4041
rect 8073 3989 8108 3990
rect 8052 3982 8108 3989
rect 8052 3962 8081 3982
rect 8101 3962 8108 3982
rect 8052 3957 8108 3962
rect 8499 3985 8531 3992
rect 9121 3985 9156 3986
rect 8499 3965 8505 3985
rect 8526 3965 8531 3985
rect 9100 3978 9156 3985
rect 8965 3968 9023 3973
rect 8052 3679 8086 3957
rect 8499 3937 8531 3965
rect 8119 3929 8531 3937
rect 8119 3903 8125 3929
rect 8151 3903 8531 3929
rect 8119 3901 8531 3903
rect 8121 3900 8161 3901
rect 8288 3875 8319 3883
rect 8288 3845 8292 3875
rect 8313 3845 8319 3875
rect 8052 3671 8087 3679
rect 8052 3651 8060 3671
rect 8080 3651 8087 3671
rect 8052 3646 8087 3651
rect 6793 3635 6829 3646
rect 8052 3645 8084 3646
rect 8288 3638 8319 3845
rect 8499 3836 8531 3901
rect 8499 3816 8503 3836
rect 8524 3816 8531 3836
rect 8499 3809 8531 3816
rect 8948 3959 9023 3968
rect 8948 3926 8957 3959
rect 9010 3926 9023 3959
rect 8948 3901 9023 3926
rect 8948 3868 8962 3901
rect 9015 3868 9023 3901
rect 8948 3862 9023 3868
rect 9100 3958 9129 3978
rect 9149 3958 9156 3978
rect 9100 3953 9156 3958
rect 9547 3981 9579 3988
rect 9547 3961 9553 3981
rect 9574 3961 9579 3981
rect 8808 3753 8909 3754
rect 8706 3740 8909 3753
rect 8706 3738 8849 3740
rect 8706 3735 8783 3738
rect 8706 3708 8709 3735
rect 8738 3711 8783 3735
rect 8812 3711 8849 3738
rect 8738 3708 8849 3711
rect 8706 3707 8849 3708
rect 8885 3707 8909 3740
rect 8706 3694 8909 3707
rect 6793 3612 6799 3635
rect 6823 3612 6829 3635
rect 8283 3629 8319 3638
rect 8228 3619 8325 3629
rect 7040 3617 8325 3619
rect 6793 3591 6829 3612
rect 6793 3568 6799 3591
rect 6823 3568 6829 3591
rect 6793 3415 6829 3568
rect 7005 3607 8325 3617
rect 7005 3569 7017 3607
rect 7042 3572 7061 3607
rect 7086 3572 8325 3607
rect 7042 3569 8325 3572
rect 7005 3566 8325 3569
rect 7005 3564 8322 3566
rect 7005 3561 7094 3564
rect 7021 3560 7093 3561
rect 8948 3551 9018 3862
rect 9100 3675 9134 3953
rect 9547 3933 9579 3961
rect 9167 3925 9579 3933
rect 9167 3899 9173 3925
rect 9199 3899 9579 3925
rect 9167 3897 9579 3899
rect 9169 3896 9209 3897
rect 9336 3871 9367 3879
rect 9336 3841 9340 3871
rect 9361 3841 9367 3871
rect 9100 3667 9135 3675
rect 9100 3647 9108 3667
rect 9128 3647 9135 3667
rect 9100 3642 9135 3647
rect 9336 3642 9367 3841
rect 9547 3832 9579 3897
rect 9547 3812 9551 3832
rect 9572 3812 9579 3832
rect 9547 3805 9579 3812
rect 9992 3958 10064 3976
rect 9992 3916 10005 3958
rect 10054 3916 10064 3958
rect 9992 3895 10064 3916
rect 9992 3853 10006 3895
rect 10055 3853 10064 3895
rect 9856 3749 9957 3750
rect 9754 3736 9957 3749
rect 9754 3734 9897 3736
rect 9754 3731 9831 3734
rect 9754 3704 9757 3731
rect 9786 3707 9831 3731
rect 9860 3707 9897 3734
rect 9786 3704 9897 3707
rect 9754 3703 9897 3704
rect 9933 3703 9957 3736
rect 9754 3690 9957 3703
rect 9100 3641 9132 3642
rect 9334 3639 9367 3642
rect 9300 3620 9368 3639
rect 9270 3608 9369 3620
rect 9992 3612 10064 3853
rect 10436 3612 10543 4041
rect 10998 4453 11105 5046
rect 11473 4995 11548 5046
rect 12514 5097 12536 5111
rect 12580 5097 12597 5134
rect 12514 5077 12597 5097
rect 12514 5011 12531 5077
rect 12585 5011 12597 5077
rect 11473 4952 11549 4995
rect 11477 4641 11549 4952
rect 12514 4987 12597 5011
rect 12514 4967 12590 4987
rect 12514 4948 12593 4967
rect 12173 4932 12245 4933
rect 12172 4924 12271 4932
rect 12172 4921 12224 4924
rect 12172 4886 12180 4921
rect 12205 4886 12224 4921
rect 12249 4886 12271 4924
rect 12172 4874 12271 4886
rect 12173 4855 12241 4874
rect 12174 4852 12207 4855
rect 12409 4852 12441 4853
rect 11584 4791 11787 4804
rect 11584 4758 11608 4791
rect 11644 4790 11787 4791
rect 11644 4787 11755 4790
rect 11644 4760 11681 4787
rect 11710 4763 11755 4787
rect 11784 4763 11787 4790
rect 11710 4760 11787 4763
rect 11644 4758 11787 4760
rect 11584 4745 11787 4758
rect 11584 4744 11685 4745
rect 11477 4599 11486 4641
rect 11535 4599 11549 4641
rect 11477 4578 11549 4599
rect 11477 4536 11487 4578
rect 11536 4536 11549 4578
rect 11477 4518 11549 4536
rect 11962 4682 11994 4689
rect 11962 4662 11969 4682
rect 11990 4662 11994 4682
rect 11962 4597 11994 4662
rect 12174 4653 12205 4852
rect 12406 4847 12441 4852
rect 12406 4827 12413 4847
rect 12433 4827 12441 4847
rect 12406 4819 12441 4827
rect 12174 4623 12180 4653
rect 12201 4623 12205 4653
rect 12174 4615 12205 4623
rect 12332 4597 12372 4598
rect 11962 4595 12374 4597
rect 11962 4569 12342 4595
rect 12368 4569 12374 4595
rect 11962 4561 12374 4569
rect 11962 4533 11994 4561
rect 12407 4541 12441 4819
rect 12523 4632 12593 4948
rect 14511 4933 14542 4934
rect 14511 4925 14556 4933
rect 13591 4902 13755 4909
rect 14511 4902 14521 4925
rect 13217 4887 14521 4902
rect 14546 4887 14556 4925
rect 15775 4928 15809 6168
rect 15775 4924 16005 4928
rect 15775 4898 15974 4924
rect 15999 4898 16005 4924
rect 15775 4890 16005 4898
rect 13217 4869 14556 4887
rect 13222 4856 13258 4869
rect 13591 4866 13755 4869
rect 12632 4787 12835 4800
rect 12632 4754 12656 4787
rect 12692 4786 12835 4787
rect 12692 4783 12803 4786
rect 12692 4756 12729 4783
rect 12758 4759 12803 4783
rect 12832 4759 12835 4786
rect 12758 4756 12835 4759
rect 12692 4754 12835 4756
rect 12632 4741 12835 4754
rect 12632 4740 12733 4741
rect 11962 4513 11967 4533
rect 11988 4513 11994 4533
rect 11962 4506 11994 4513
rect 12385 4536 12441 4541
rect 12385 4516 12392 4536
rect 12412 4516 12441 4536
rect 12518 4626 12593 4632
rect 12518 4593 12526 4626
rect 12579 4593 12593 4626
rect 12518 4568 12593 4593
rect 12518 4535 12531 4568
rect 12584 4535 12593 4568
rect 12518 4526 12593 4535
rect 13010 4678 13042 4685
rect 13010 4658 13017 4678
rect 13038 4658 13042 4678
rect 13010 4593 13042 4658
rect 13222 4649 13253 4856
rect 16359 4854 16391 4855
rect 13457 4848 13489 4849
rect 13454 4843 13489 4848
rect 13454 4823 13461 4843
rect 13481 4823 13489 4843
rect 13454 4815 13489 4823
rect 13222 4619 13228 4649
rect 13249 4619 13253 4649
rect 13222 4611 13253 4619
rect 13380 4593 13420 4594
rect 13010 4591 13422 4593
rect 13010 4565 13390 4591
rect 13416 4565 13422 4591
rect 13010 4557 13422 4565
rect 13010 4529 13042 4557
rect 13455 4537 13489 4815
rect 15534 4793 15737 4806
rect 15534 4760 15558 4793
rect 15594 4792 15737 4793
rect 15594 4789 15705 4792
rect 15594 4762 15631 4789
rect 15660 4765 15705 4789
rect 15734 4765 15737 4792
rect 15660 4762 15737 4765
rect 15594 4760 15737 4762
rect 15534 4747 15737 4760
rect 15534 4746 15635 4747
rect 12518 4521 12576 4526
rect 12385 4509 12441 4516
rect 13010 4509 13015 4529
rect 13036 4509 13042 4529
rect 12385 4508 12420 4509
rect 13010 4502 13042 4509
rect 13433 4532 13489 4537
rect 13433 4512 13440 4532
rect 13460 4512 13489 4532
rect 13433 4505 13489 4512
rect 15912 4684 15944 4691
rect 15912 4664 15919 4684
rect 15940 4664 15944 4684
rect 15912 4599 15944 4664
rect 16124 4655 16155 4852
rect 16356 4849 16391 4854
rect 16356 4829 16363 4849
rect 16383 4829 16391 4849
rect 16356 4821 16391 4829
rect 16124 4625 16130 4655
rect 16151 4625 16155 4655
rect 16124 4617 16155 4625
rect 16282 4599 16322 4600
rect 15912 4597 16324 4599
rect 15912 4571 16292 4597
rect 16318 4571 16324 4597
rect 15912 4563 16324 4571
rect 15912 4535 15944 4563
rect 15912 4515 15917 4535
rect 15938 4515 15944 4535
rect 15912 4508 15944 4515
rect 16114 4537 16162 4544
rect 16357 4543 16391 4821
rect 16114 4517 16121 4537
rect 16154 4517 16162 4537
rect 13433 4504 13468 4505
rect 11676 4453 11787 4457
rect 13459 4453 15029 4454
rect 10998 4449 15029 4453
rect 15354 4449 15772 4462
rect 10998 4437 15772 4449
rect 10998 4435 15634 4437
rect 10998 4415 11684 4435
rect 11703 4415 11761 4435
rect 11780 4431 15634 4435
rect 11780 4415 12732 4431
rect 10998 4411 12732 4415
rect 12751 4411 12809 4431
rect 12828 4417 15634 4431
rect 15653 4417 15711 4437
rect 15730 4417 15772 4437
rect 12828 4411 15772 4417
rect 10998 4397 15772 4411
rect 10998 3774 11105 4397
rect 12724 4394 12835 4397
rect 15354 4391 15772 4397
rect 11484 4348 11548 4352
rect 11480 4342 11548 4348
rect 11480 4309 11497 4342
rect 11537 4309 11548 4342
rect 11480 4297 11548 4309
rect 12531 4311 12596 4333
rect 11480 4295 11537 4297
rect 11484 3934 11535 4295
rect 12531 4272 12548 4311
rect 12593 4272 12596 4311
rect 12172 4227 12207 4229
rect 12172 4218 12276 4227
rect 12172 4217 12223 4218
rect 12172 4197 12175 4217
rect 12200 4198 12223 4217
rect 12255 4198 12276 4218
rect 12200 4197 12276 4198
rect 12172 4190 12276 4197
rect 12172 4178 12207 4190
rect 11584 4112 11787 4125
rect 11584 4079 11608 4112
rect 11644 4111 11787 4112
rect 11644 4108 11755 4111
rect 11644 4081 11681 4108
rect 11710 4084 11755 4108
rect 11784 4084 11787 4111
rect 11710 4081 11787 4084
rect 11644 4079 11787 4081
rect 11584 4066 11787 4079
rect 11584 4065 11685 4066
rect 11962 4003 11994 4010
rect 11962 3983 11969 4003
rect 11990 3983 11994 4003
rect 11473 3925 11538 3934
rect 11473 3888 11483 3925
rect 11523 3891 11538 3925
rect 11962 3918 11994 3983
rect 12174 3974 12205 4178
rect 12409 4173 12441 4174
rect 12406 4168 12441 4173
rect 12406 4148 12413 4168
rect 12433 4148 12441 4168
rect 12406 4140 12441 4148
rect 12174 3944 12180 3974
rect 12201 3944 12205 3974
rect 12174 3936 12205 3944
rect 12332 3918 12372 3919
rect 11962 3916 12374 3918
rect 11523 3888 11540 3891
rect 11473 3869 11540 3888
rect 11473 3848 11487 3869
rect 11523 3848 11540 3869
rect 11473 3841 11540 3848
rect 11962 3890 12342 3916
rect 12368 3890 12374 3916
rect 11962 3882 12374 3890
rect 11962 3854 11994 3882
rect 12407 3862 12441 4140
rect 12531 3972 12596 4272
rect 14668 4233 14705 4254
rect 14668 4196 14679 4233
rect 14696 4209 14705 4233
rect 14696 4196 14706 4209
rect 14668 4186 14706 4196
rect 14669 4182 14706 4186
rect 14669 4176 14702 4182
rect 14079 4107 14282 4120
rect 14079 4074 14103 4107
rect 14139 4106 14282 4107
rect 14139 4103 14250 4106
rect 14139 4076 14176 4103
rect 14205 4079 14250 4103
rect 14279 4079 14282 4106
rect 14205 4076 14282 4079
rect 14139 4074 14282 4076
rect 14079 4061 14282 4074
rect 14079 4060 14180 4061
rect 14457 3998 14489 4005
rect 14457 3978 14464 3998
rect 14485 3978 14489 3998
rect 11962 3834 11967 3854
rect 11988 3834 11994 3854
rect 11962 3827 11994 3834
rect 12385 3857 12441 3862
rect 12385 3837 12392 3857
rect 12412 3837 12441 3857
rect 12385 3830 12441 3837
rect 12521 3961 12601 3972
rect 12521 3935 12538 3961
rect 12578 3935 12601 3961
rect 12521 3908 12601 3935
rect 12521 3882 12542 3908
rect 12582 3882 12601 3908
rect 12521 3863 12601 3882
rect 12521 3837 12545 3863
rect 12585 3837 12601 3863
rect 13595 3907 13700 3928
rect 14457 3913 14489 3978
rect 14669 3969 14700 4176
rect 14904 4168 14936 4169
rect 14901 4163 14936 4168
rect 14901 4143 14908 4163
rect 14928 4143 14936 4163
rect 14901 4135 14936 4143
rect 14669 3939 14675 3969
rect 14696 3939 14700 3969
rect 14669 3931 14700 3939
rect 14827 3913 14867 3914
rect 14457 3911 14869 3913
rect 13595 3901 14071 3907
rect 13595 3899 13652 3901
rect 13595 3868 13607 3899
rect 13632 3878 13652 3899
rect 13678 3894 14071 3901
rect 13678 3878 14032 3894
rect 13632 3871 14032 3878
rect 14058 3871 14071 3894
rect 13632 3868 14071 3871
rect 13595 3858 14071 3868
rect 14457 3885 14837 3911
rect 14863 3885 14869 3911
rect 14457 3877 14869 3885
rect 13595 3856 13700 3858
rect 12385 3829 12420 3830
rect 12521 3825 12601 3837
rect 14457 3849 14489 3877
rect 14902 3857 14936 4135
rect 14457 3829 14462 3849
rect 14483 3829 14489 3849
rect 14457 3822 14489 3829
rect 14880 3852 14936 3857
rect 14880 3832 14887 3852
rect 14907 3832 14936 3852
rect 14880 3825 14936 3832
rect 14880 3824 14915 3825
rect 11676 3774 11787 3778
rect 13418 3774 15071 3777
rect 10996 3756 15071 3774
rect 10996 3736 11684 3756
rect 11703 3736 11761 3756
rect 11780 3751 15071 3756
rect 11780 3736 14179 3751
rect 10996 3731 14179 3736
rect 14198 3731 14256 3751
rect 14275 3731 15071 3751
rect 10996 3721 15071 3731
rect 10996 3718 11621 3721
rect 11808 3718 15071 3721
rect 9270 3570 9292 3608
rect 9317 3573 9336 3608
rect 9361 3573 9369 3608
rect 9317 3570 9369 3573
rect 9270 3562 9369 3570
rect 9296 3561 9368 3562
rect 8947 3535 9018 3551
rect 8947 3519 8967 3535
rect 8948 3489 8967 3519
rect 8950 3469 8967 3489
rect 8997 3489 9018 3535
rect 9990 3531 10068 3612
rect 10435 3557 10543 3612
rect 8997 3469 9017 3489
rect 8950 3450 9017 3469
rect 9990 3429 10069 3531
rect 6784 3406 6870 3415
rect 6784 3388 6803 3406
rect 6855 3388 6870 3406
rect 6784 3384 6870 3388
rect 9954 3411 10075 3429
rect 9954 3409 10025 3411
rect 9954 3368 9969 3409
rect 10006 3370 10025 3409
rect 10062 3370 10075 3411
rect 10006 3368 10075 3370
rect 9954 3358 10075 3368
rect 7259 3330 7370 3333
rect 6574 3329 8123 3330
rect 10436 3329 10543 3557
rect 10998 3490 11105 3718
rect 13418 3717 15071 3718
rect 14171 3714 14282 3717
rect 11466 3679 11587 3689
rect 11466 3677 11535 3679
rect 11466 3636 11479 3677
rect 11516 3638 11535 3677
rect 11572 3638 11587 3679
rect 11516 3636 11587 3638
rect 11466 3618 11587 3636
rect 11472 3516 11551 3618
rect 12524 3578 12591 3597
rect 12524 3558 12544 3578
rect 10998 3435 11106 3490
rect 11473 3435 11551 3516
rect 12523 3512 12544 3558
rect 12574 3558 12591 3578
rect 12574 3528 12593 3558
rect 12574 3512 12594 3528
rect 12523 3496 12594 3512
rect 12173 3485 12245 3486
rect 12172 3477 12271 3485
rect 12172 3474 12224 3477
rect 12172 3439 12180 3474
rect 12205 3439 12224 3474
rect 12249 3439 12271 3477
rect 6574 3326 9733 3329
rect 9920 3326 10545 3329
rect 6574 3316 10545 3326
rect 6574 3296 7266 3316
rect 7285 3296 7343 3316
rect 7362 3311 10545 3316
rect 7362 3296 9761 3311
rect 6574 3291 9761 3296
rect 9780 3291 9838 3311
rect 9857 3291 10545 3311
rect 6574 3273 10545 3291
rect 6574 3270 8123 3273
rect 9754 3269 9865 3273
rect 6626 3222 6661 3223
rect 6605 3215 6661 3222
rect 6605 3195 6634 3215
rect 6654 3195 6661 3215
rect 6605 3190 6661 3195
rect 7052 3218 7084 3225
rect 7052 3198 7058 3218
rect 7079 3198 7084 3218
rect 6605 2912 6639 3190
rect 7052 3170 7084 3198
rect 6672 3162 7084 3170
rect 6672 3136 6678 3162
rect 6704 3136 7084 3162
rect 6672 3134 7084 3136
rect 6674 3133 6714 3134
rect 6841 3108 6872 3116
rect 6841 3078 6845 3108
rect 6866 3078 6872 3108
rect 6605 2904 6640 2912
rect 6605 2884 6613 2904
rect 6633 2884 6640 2904
rect 6605 2879 6640 2884
rect 6605 2878 6637 2879
rect 6841 2877 6872 3078
rect 7052 3069 7084 3134
rect 7052 3049 7056 3069
rect 7077 3049 7084 3069
rect 7052 3042 7084 3049
rect 7646 3209 7739 3216
rect 7646 3168 7670 3209
rect 7724 3168 7739 3209
rect 7361 2986 7462 2987
rect 7259 2973 7462 2986
rect 7259 2971 7402 2973
rect 7259 2968 7336 2971
rect 7259 2941 7262 2968
rect 7291 2944 7336 2968
rect 7365 2944 7402 2971
rect 7291 2941 7402 2944
rect 7259 2940 7402 2941
rect 7438 2940 7462 2973
rect 7259 2927 7462 2940
rect 7646 2795 7739 3168
rect 8940 3210 9020 3222
rect 9121 3217 9156 3218
rect 8940 3184 8956 3210
rect 8996 3184 9020 3210
rect 8940 3165 9020 3184
rect 8940 3139 8959 3165
rect 8999 3139 9020 3165
rect 8940 3112 9020 3139
rect 8940 3086 8963 3112
rect 9003 3086 9020 3112
rect 8940 3075 9020 3086
rect 9100 3210 9156 3217
rect 9100 3190 9129 3210
rect 9149 3190 9156 3210
rect 9100 3185 9156 3190
rect 9547 3213 9579 3220
rect 9547 3193 9553 3213
rect 9574 3193 9579 3213
rect 7646 2751 7664 2795
rect 7724 2751 7739 2795
rect 7646 2736 7739 2751
rect 8945 2775 9010 3075
rect 9100 2907 9134 3185
rect 9547 3165 9579 3193
rect 9167 3157 9579 3165
rect 9167 3131 9173 3157
rect 9199 3131 9579 3157
rect 10001 3199 10068 3206
rect 10001 3178 10018 3199
rect 10054 3178 10068 3199
rect 10001 3159 10068 3178
rect 10001 3156 10018 3159
rect 9167 3129 9579 3131
rect 9169 3128 9209 3129
rect 9336 3103 9367 3111
rect 9336 3073 9340 3103
rect 9361 3073 9367 3103
rect 9100 2899 9135 2907
rect 9100 2879 9108 2899
rect 9128 2879 9135 2899
rect 9100 2874 9135 2879
rect 9100 2873 9132 2874
rect 9336 2869 9367 3073
rect 9547 3064 9579 3129
rect 10003 3122 10018 3156
rect 10058 3122 10068 3159
rect 10003 3113 10068 3122
rect 9547 3044 9551 3064
rect 9572 3044 9579 3064
rect 9547 3037 9579 3044
rect 9856 2981 9957 2982
rect 9754 2968 9957 2981
rect 9754 2966 9897 2968
rect 9754 2963 9831 2966
rect 9754 2936 9757 2963
rect 9786 2939 9831 2963
rect 9860 2939 9897 2966
rect 9786 2936 9897 2939
rect 9754 2935 9897 2936
rect 9933 2935 9957 2968
rect 9754 2922 9957 2935
rect 9334 2857 9369 2869
rect 9265 2850 9369 2857
rect 9265 2849 9341 2850
rect 9265 2829 9286 2849
rect 9318 2830 9341 2849
rect 9366 2830 9369 2850
rect 9318 2829 9369 2830
rect 9265 2820 9369 2829
rect 9334 2818 9369 2820
rect 8945 2736 8948 2775
rect 8993 2736 9010 2775
rect 10006 2752 10057 3113
rect 10004 2750 10061 2752
rect 8945 2714 9010 2736
rect 9993 2738 10061 2750
rect 9993 2705 10004 2738
rect 10044 2705 10061 2738
rect 9993 2699 10061 2705
rect 9993 2695 10057 2699
rect 8706 2650 8817 2653
rect 10436 2650 10543 3273
rect 6969 2636 10543 2650
rect 6969 2616 8713 2636
rect 8732 2616 8790 2636
rect 8809 2632 10543 2636
rect 8809 2616 9761 2632
rect 6969 2612 9761 2616
rect 9780 2612 9838 2632
rect 9857 2612 10543 2632
rect 6969 2594 10543 2612
rect 6969 2593 8082 2594
rect 9754 2590 9865 2594
rect 8073 2542 8108 2543
rect 8052 2535 8108 2542
rect 8052 2515 8081 2535
rect 8101 2515 8108 2535
rect 8052 2510 8108 2515
rect 8499 2538 8531 2545
rect 9121 2538 9156 2539
rect 8499 2518 8505 2538
rect 8526 2518 8531 2538
rect 9100 2531 9156 2538
rect 8965 2521 9023 2526
rect 5888 2475 7741 2508
rect 5888 2410 5953 2475
rect 6084 2455 7741 2475
rect 6084 2414 7677 2455
rect 7713 2414 7741 2455
rect 7839 2475 7903 2494
rect 7839 2436 7856 2475
rect 7890 2436 7903 2475
rect 7839 2417 7903 2436
rect 6084 2410 7741 2414
rect 5888 2385 7741 2410
rect 7652 2382 7734 2385
rect 7841 1905 7903 2417
rect 8052 2232 8086 2510
rect 8499 2490 8531 2518
rect 8119 2482 8531 2490
rect 8119 2456 8125 2482
rect 8151 2456 8531 2482
rect 8119 2454 8531 2456
rect 8121 2453 8161 2454
rect 8288 2428 8319 2436
rect 8288 2398 8292 2428
rect 8313 2398 8319 2428
rect 8052 2224 8087 2232
rect 8052 2204 8060 2224
rect 8080 2204 8087 2224
rect 8052 2199 8087 2204
rect 8052 2198 8084 2199
rect 8288 2191 8319 2398
rect 8499 2389 8531 2454
rect 8499 2369 8503 2389
rect 8524 2369 8531 2389
rect 8499 2362 8531 2369
rect 8948 2512 9023 2521
rect 8948 2479 8957 2512
rect 9010 2479 9023 2512
rect 8948 2454 9023 2479
rect 8948 2421 8962 2454
rect 9015 2421 9023 2454
rect 8948 2415 9023 2421
rect 9100 2511 9129 2531
rect 9149 2511 9156 2531
rect 9100 2506 9156 2511
rect 9547 2534 9579 2541
rect 9547 2514 9553 2534
rect 9574 2514 9579 2534
rect 8808 2306 8909 2307
rect 8706 2293 8909 2306
rect 8706 2291 8849 2293
rect 8706 2288 8783 2291
rect 8706 2261 8709 2288
rect 8738 2264 8783 2288
rect 8812 2264 8849 2291
rect 8738 2261 8849 2264
rect 8706 2260 8849 2261
rect 8885 2260 8909 2293
rect 8706 2247 8909 2260
rect 8283 2173 8319 2191
rect 8250 2172 8319 2173
rect 8230 2160 8319 2172
rect 8230 2122 8242 2160
rect 8267 2125 8286 2160
rect 8311 2125 8319 2160
rect 8267 2122 8319 2125
rect 8230 2114 8319 2122
rect 8246 2113 8318 2114
rect 7799 1847 7915 1905
rect 8948 1894 9018 2415
rect 9100 2228 9134 2506
rect 9547 2486 9579 2514
rect 9167 2478 9579 2486
rect 9167 2452 9173 2478
rect 9199 2452 9579 2478
rect 9167 2450 9579 2452
rect 9169 2449 9209 2450
rect 9336 2424 9367 2432
rect 9336 2394 9340 2424
rect 9361 2394 9367 2424
rect 9100 2220 9135 2228
rect 9100 2200 9108 2220
rect 9128 2200 9135 2220
rect 9100 2195 9135 2200
rect 9336 2195 9367 2394
rect 9547 2385 9579 2450
rect 9547 2365 9551 2385
rect 9572 2365 9579 2385
rect 9547 2358 9579 2365
rect 9992 2511 10064 2529
rect 9992 2469 10005 2511
rect 10054 2469 10064 2511
rect 9992 2448 10064 2469
rect 9992 2406 10006 2448
rect 10055 2406 10064 2448
rect 9856 2302 9957 2303
rect 9754 2289 9957 2302
rect 9754 2287 9897 2289
rect 9754 2284 9831 2287
rect 9754 2257 9757 2284
rect 9786 2260 9831 2284
rect 9860 2260 9897 2287
rect 9786 2257 9897 2260
rect 9754 2256 9897 2257
rect 9933 2256 9957 2289
rect 9754 2243 9957 2256
rect 9100 2194 9132 2195
rect 9334 2192 9367 2195
rect 9300 2173 9368 2192
rect 9270 2161 9369 2173
rect 9270 2123 9292 2161
rect 9317 2126 9336 2161
rect 9361 2126 9369 2161
rect 9317 2123 9369 2126
rect 9270 2115 9369 2123
rect 9296 2114 9368 2115
rect 7799 1776 7811 1847
rect 7890 1776 7915 1847
rect 7799 1756 7915 1776
rect 8929 1693 9031 1894
rect 9992 1886 10064 2406
rect 10436 1982 10543 2594
rect 10998 3006 11105 3435
rect 11477 3194 11549 3435
rect 12172 3427 12271 3439
rect 12173 3408 12241 3427
rect 12174 3405 12207 3408
rect 12409 3405 12441 3406
rect 11584 3344 11787 3357
rect 11584 3311 11608 3344
rect 11644 3343 11787 3344
rect 11644 3340 11755 3343
rect 11644 3313 11681 3340
rect 11710 3316 11755 3340
rect 11784 3316 11787 3343
rect 11710 3313 11787 3316
rect 11644 3311 11787 3313
rect 11584 3298 11787 3311
rect 11584 3297 11685 3298
rect 11477 3152 11486 3194
rect 11535 3152 11549 3194
rect 11477 3131 11549 3152
rect 11477 3089 11487 3131
rect 11536 3089 11549 3131
rect 11477 3071 11549 3089
rect 11962 3235 11994 3242
rect 11962 3215 11969 3235
rect 11990 3215 11994 3235
rect 11962 3150 11994 3215
rect 12174 3206 12205 3405
rect 12406 3400 12441 3405
rect 12406 3380 12413 3400
rect 12433 3380 12441 3400
rect 12406 3372 12441 3380
rect 12174 3176 12180 3206
rect 12201 3176 12205 3206
rect 12174 3168 12205 3176
rect 12332 3150 12372 3151
rect 11962 3148 12374 3150
rect 11962 3122 12342 3148
rect 12368 3122 12374 3148
rect 11962 3114 12374 3122
rect 11962 3086 11994 3114
rect 12407 3094 12441 3372
rect 12523 3185 12593 3496
rect 13220 3487 14562 3492
rect 13220 3485 14519 3487
rect 13217 3459 14519 3485
rect 14547 3459 14562 3487
rect 13217 3451 14562 3459
rect 13217 3426 13256 3451
rect 13217 3409 13258 3426
rect 13217 3402 13256 3409
rect 12632 3340 12835 3353
rect 12632 3307 12656 3340
rect 12692 3339 12835 3340
rect 12692 3336 12803 3339
rect 12692 3309 12729 3336
rect 12758 3312 12803 3336
rect 12832 3312 12835 3339
rect 12758 3309 12835 3312
rect 12692 3307 12835 3309
rect 12632 3294 12835 3307
rect 12632 3293 12733 3294
rect 11962 3066 11967 3086
rect 11988 3066 11994 3086
rect 11962 3059 11994 3066
rect 12385 3089 12441 3094
rect 12385 3069 12392 3089
rect 12412 3069 12441 3089
rect 12518 3179 12593 3185
rect 12518 3146 12526 3179
rect 12579 3146 12593 3179
rect 12518 3121 12593 3146
rect 12518 3088 12531 3121
rect 12584 3088 12593 3121
rect 12518 3079 12593 3088
rect 13010 3231 13042 3238
rect 13010 3211 13017 3231
rect 13038 3211 13042 3231
rect 13010 3146 13042 3211
rect 13222 3202 13253 3402
rect 13457 3401 13489 3402
rect 13454 3396 13489 3401
rect 13454 3376 13461 3396
rect 13481 3376 13489 3396
rect 13454 3368 13489 3376
rect 13222 3172 13228 3202
rect 13249 3172 13253 3202
rect 13222 3164 13253 3172
rect 13380 3146 13420 3147
rect 13010 3144 13422 3146
rect 13010 3118 13390 3144
rect 13416 3118 13422 3144
rect 13010 3110 13422 3118
rect 13010 3082 13042 3110
rect 13455 3090 13489 3368
rect 12518 3074 12576 3079
rect 12385 3062 12441 3069
rect 13010 3062 13015 3082
rect 13036 3062 13042 3082
rect 12385 3061 12420 3062
rect 13010 3055 13042 3062
rect 13433 3085 13489 3090
rect 13433 3065 13440 3085
rect 13460 3065 13489 3085
rect 13433 3058 13489 3065
rect 13433 3057 13468 3058
rect 11676 3006 11787 3010
rect 13551 3006 15071 3007
rect 10998 2988 15071 3006
rect 10998 2968 11684 2988
rect 11703 2968 11761 2988
rect 11780 2984 15071 2988
rect 11780 2968 12732 2984
rect 10998 2964 12732 2968
rect 12751 2964 12809 2984
rect 12828 2964 15071 2984
rect 10998 2950 15071 2964
rect 10998 2327 11105 2950
rect 12724 2947 12835 2950
rect 11484 2901 11548 2905
rect 11480 2895 11548 2901
rect 11480 2862 11497 2895
rect 11537 2862 11548 2895
rect 11480 2850 11548 2862
rect 12531 2864 12596 2886
rect 11480 2848 11537 2850
rect 11484 2487 11535 2848
rect 12531 2825 12548 2864
rect 12593 2825 12596 2864
rect 12172 2780 12207 2782
rect 12172 2771 12276 2780
rect 12172 2770 12223 2771
rect 12172 2750 12175 2770
rect 12200 2751 12223 2770
rect 12255 2751 12276 2771
rect 12200 2750 12276 2751
rect 12172 2743 12276 2750
rect 12172 2731 12207 2743
rect 11584 2665 11787 2678
rect 11584 2632 11608 2665
rect 11644 2664 11787 2665
rect 11644 2661 11755 2664
rect 11644 2634 11681 2661
rect 11710 2637 11755 2661
rect 11784 2637 11787 2664
rect 11710 2634 11787 2637
rect 11644 2632 11787 2634
rect 11584 2619 11787 2632
rect 11584 2618 11685 2619
rect 11962 2556 11994 2563
rect 11962 2536 11969 2556
rect 11990 2536 11994 2556
rect 11473 2478 11538 2487
rect 11473 2441 11483 2478
rect 11523 2444 11538 2478
rect 11962 2471 11994 2536
rect 12174 2527 12205 2731
rect 12409 2726 12441 2727
rect 12406 2721 12441 2726
rect 12406 2701 12413 2721
rect 12433 2701 12441 2721
rect 12406 2693 12441 2701
rect 12174 2497 12180 2527
rect 12201 2497 12205 2527
rect 12174 2489 12205 2497
rect 12332 2471 12372 2472
rect 11962 2469 12374 2471
rect 11523 2441 11540 2444
rect 11473 2422 11540 2441
rect 11473 2401 11487 2422
rect 11523 2401 11540 2422
rect 11473 2394 11540 2401
rect 11962 2443 12342 2469
rect 12368 2443 12374 2469
rect 11962 2435 12374 2443
rect 11962 2407 11994 2435
rect 12407 2415 12441 2693
rect 12531 2562 12596 2825
rect 12531 2558 12592 2562
rect 11962 2387 11967 2407
rect 11988 2387 11994 2407
rect 11962 2380 11994 2387
rect 12385 2410 12441 2415
rect 12385 2390 12392 2410
rect 12412 2390 12441 2410
rect 12385 2383 12441 2390
rect 12385 2382 12420 2383
rect 11676 2327 11787 2331
rect 10996 2309 12315 2327
rect 10996 2289 11684 2309
rect 11703 2289 11761 2309
rect 11780 2289 12315 2309
rect 10996 2271 12315 2289
rect 10998 2151 11105 2271
rect 11466 2232 11587 2242
rect 11466 2230 11535 2232
rect 11466 2189 11479 2230
rect 11516 2191 11535 2230
rect 11572 2191 11587 2232
rect 11516 2189 11587 2191
rect 11466 2171 11587 2189
rect 10435 1946 10543 1982
rect 10590 2105 10744 2130
rect 10590 1993 10603 2105
rect 10724 1993 10744 2105
rect 8893 1656 9059 1693
rect 8893 1577 8930 1656
rect 9014 1577 9059 1656
rect 8893 1539 9059 1577
rect 9970 1485 10067 1886
rect 10428 1810 10548 1946
rect 10435 1804 10543 1810
rect 9900 1456 10075 1485
rect 9900 1377 9946 1456
rect 10046 1377 10075 1456
rect 9900 1352 10075 1377
rect 10435 1261 10539 1804
rect 10278 1231 10549 1261
rect 10278 1144 10312 1231
rect 10382 1223 10549 1231
rect 10382 1144 10445 1223
rect 10278 1136 10445 1144
rect 10515 1136 10549 1223
rect 10278 1090 10549 1136
rect 5402 775 10311 793
rect 5402 729 10213 775
rect 10289 729 10311 775
rect 5402 718 10311 729
rect 10163 333 10292 340
rect 10163 329 10187 333
rect 0 274 10187 329
rect 10218 274 10249 333
rect 10280 274 10292 333
rect 0 265 10292 274
rect 10163 261 10292 265
rect 10383 157 10455 1090
rect 10590 1019 10744 1993
rect 10588 1003 10744 1019
rect 10797 2078 10931 2107
rect 10797 1966 10835 2078
rect 10914 1966 10931 2078
rect 10998 2071 11106 2151
rect 10797 1013 10931 1966
rect 10999 1259 11106 2071
rect 11472 2099 11537 2171
rect 11472 2033 11540 2099
rect 11473 1487 11540 2033
rect 12527 1671 12592 2558
rect 13570 2288 13707 2292
rect 13557 2284 13714 2288
rect 13557 2177 13594 2284
rect 13694 2177 13714 2284
rect 13557 2135 13714 2177
rect 13570 1887 13707 2135
rect 13560 1845 13726 1887
rect 13560 1770 13589 1845
rect 13706 1770 13726 1845
rect 13560 1754 13726 1770
rect 12516 1650 12653 1671
rect 12516 1575 12541 1650
rect 12611 1575 12653 1650
rect 12516 1544 12653 1575
rect 11459 1438 11634 1487
rect 11459 1359 11492 1438
rect 11592 1359 11634 1438
rect 11459 1354 11634 1359
rect 10999 1217 11147 1259
rect 10999 1209 11039 1217
rect 11001 1130 11039 1209
rect 11109 1130 11147 1217
rect 11001 1092 11147 1130
rect 10588 978 10740 1003
rect 10588 883 10618 978
rect 10708 883 10740 978
rect 10588 870 10740 883
rect 10793 977 10932 1013
rect 10793 882 10807 977
rect 10897 882 10932 977
rect 10793 864 10932 882
rect 16114 797 16162 4517
rect 16335 4538 16391 4543
rect 16335 4518 16342 4538
rect 16362 4518 16391 4538
rect 16335 4511 16391 4518
rect 16335 4510 16370 4511
rect 16439 4420 16467 7228
rect 19652 7183 19717 7483
rect 19807 7315 19841 7593
rect 20254 7573 20286 7601
rect 19874 7565 20286 7573
rect 19874 7539 19880 7565
rect 19906 7539 20286 7565
rect 20708 7607 20775 7614
rect 20708 7586 20725 7607
rect 20761 7586 20775 7607
rect 20708 7567 20775 7586
rect 20708 7564 20725 7567
rect 19874 7537 20286 7539
rect 19876 7536 19916 7537
rect 20043 7511 20074 7519
rect 20043 7481 20047 7511
rect 20068 7481 20074 7511
rect 19807 7307 19842 7315
rect 19807 7287 19815 7307
rect 19835 7287 19842 7307
rect 19807 7282 19842 7287
rect 19807 7281 19839 7282
rect 20043 7277 20074 7481
rect 20254 7472 20286 7537
rect 20710 7530 20725 7564
rect 20765 7530 20775 7567
rect 20710 7521 20775 7530
rect 20254 7452 20258 7472
rect 20279 7452 20286 7472
rect 20254 7445 20286 7452
rect 20563 7389 20664 7390
rect 20461 7376 20664 7389
rect 20461 7374 20604 7376
rect 20461 7371 20538 7374
rect 20461 7344 20464 7371
rect 20493 7347 20538 7371
rect 20567 7347 20604 7374
rect 20493 7344 20604 7347
rect 20461 7343 20604 7344
rect 20640 7343 20664 7376
rect 20461 7330 20664 7343
rect 20041 7265 20076 7277
rect 19972 7258 20076 7265
rect 19972 7257 20048 7258
rect 19972 7237 19993 7257
rect 20025 7238 20048 7257
rect 20073 7238 20076 7258
rect 20025 7237 20076 7238
rect 19972 7228 20076 7237
rect 20041 7226 20076 7228
rect 19652 7144 19655 7183
rect 19700 7144 19717 7183
rect 20713 7160 20764 7521
rect 20711 7158 20768 7160
rect 19652 7122 19717 7144
rect 20700 7146 20768 7158
rect 20700 7113 20711 7146
rect 20751 7113 20768 7146
rect 20700 7107 20768 7113
rect 20700 7103 20764 7107
rect 19413 7058 19524 7061
rect 21143 7058 21250 7681
rect 17707 7044 21250 7058
rect 17707 7024 19420 7044
rect 19439 7024 19497 7044
rect 19516 7040 21250 7044
rect 19516 7024 20468 7040
rect 17707 7020 20468 7024
rect 20487 7020 20545 7040
rect 20564 7020 21250 7040
rect 17707 7002 21250 7020
rect 17707 7001 18697 7002
rect 20461 6998 20572 7002
rect 18780 6950 18815 6951
rect 18759 6943 18815 6950
rect 18759 6923 18788 6943
rect 18808 6923 18815 6943
rect 18759 6918 18815 6923
rect 19206 6946 19238 6953
rect 19828 6946 19863 6947
rect 19206 6926 19212 6946
rect 19233 6926 19238 6946
rect 19807 6939 19863 6946
rect 19672 6929 19730 6934
rect 18759 6640 18793 6918
rect 19206 6898 19238 6926
rect 18826 6890 19238 6898
rect 18826 6864 18832 6890
rect 18858 6864 19238 6890
rect 18826 6862 19238 6864
rect 18828 6861 18868 6862
rect 18995 6836 19026 6844
rect 18995 6806 18999 6836
rect 19020 6806 19026 6836
rect 18759 6632 18794 6640
rect 18759 6612 18767 6632
rect 18787 6612 18794 6632
rect 18759 6607 18794 6612
rect 18759 6606 18791 6607
rect 18995 6606 19026 6806
rect 19206 6797 19238 6862
rect 19206 6777 19210 6797
rect 19231 6777 19238 6797
rect 19206 6770 19238 6777
rect 19655 6920 19730 6929
rect 19655 6887 19664 6920
rect 19717 6887 19730 6920
rect 19655 6862 19730 6887
rect 19655 6829 19669 6862
rect 19722 6829 19730 6862
rect 19655 6823 19730 6829
rect 19807 6919 19836 6939
rect 19856 6919 19863 6939
rect 19807 6914 19863 6919
rect 20254 6942 20286 6949
rect 20254 6922 20260 6942
rect 20281 6922 20286 6942
rect 19515 6714 19616 6715
rect 19413 6701 19616 6714
rect 19413 6699 19556 6701
rect 19413 6696 19490 6699
rect 19413 6669 19416 6696
rect 19445 6672 19490 6696
rect 19519 6672 19556 6699
rect 19445 6669 19556 6672
rect 19413 6668 19556 6669
rect 19592 6668 19616 6701
rect 19413 6655 19616 6668
rect 18992 6599 19031 6606
rect 18990 6582 19031 6599
rect 18992 6557 19031 6582
rect 17686 6549 19031 6557
rect 17686 6521 17701 6549
rect 17729 6523 19031 6549
rect 17729 6521 19028 6523
rect 17686 6516 19028 6521
rect 19655 6512 19725 6823
rect 19807 6636 19841 6914
rect 20254 6894 20286 6922
rect 19874 6886 20286 6894
rect 19874 6860 19880 6886
rect 19906 6860 20286 6886
rect 19874 6858 20286 6860
rect 19876 6857 19916 6858
rect 20043 6832 20074 6840
rect 20043 6802 20047 6832
rect 20068 6802 20074 6832
rect 19807 6628 19842 6636
rect 19807 6608 19815 6628
rect 19835 6608 19842 6628
rect 19807 6603 19842 6608
rect 20043 6603 20074 6802
rect 20254 6793 20286 6858
rect 20254 6773 20258 6793
rect 20279 6773 20286 6793
rect 20254 6766 20286 6773
rect 20699 6919 20771 6937
rect 20699 6877 20712 6919
rect 20761 6877 20771 6919
rect 20699 6856 20771 6877
rect 20699 6814 20713 6856
rect 20762 6814 20771 6856
rect 20563 6710 20664 6711
rect 20461 6697 20664 6710
rect 20461 6695 20604 6697
rect 20461 6692 20538 6695
rect 20461 6665 20464 6692
rect 20493 6668 20538 6692
rect 20567 6668 20604 6695
rect 20493 6665 20604 6668
rect 20461 6664 20604 6665
rect 20640 6664 20664 6697
rect 20461 6651 20664 6664
rect 19807 6602 19839 6603
rect 20041 6600 20074 6603
rect 20007 6581 20075 6600
rect 19977 6569 20076 6581
rect 20699 6573 20771 6814
rect 21143 6573 21250 7002
rect 21962 7424 22069 7884
rect 22441 7612 22513 7906
rect 23137 7903 23209 7904
rect 23136 7895 23235 7903
rect 23489 7898 23566 8081
rect 24777 8082 24861 8093
rect 24777 8054 24805 8082
rect 24849 8054 24861 8082
rect 24591 8003 24665 8031
rect 24591 7955 24614 8003
rect 24651 7955 24665 8003
rect 24777 8025 24861 8054
rect 24777 7997 24802 8025
rect 24846 7997 24861 8025
rect 24777 7964 24861 7997
rect 24591 7946 24665 7955
rect 24187 7904 24259 7905
rect 23136 7892 23188 7895
rect 23136 7857 23144 7892
rect 23169 7857 23188 7892
rect 23213 7857 23235 7895
rect 23136 7845 23235 7857
rect 23487 7869 23566 7898
rect 24186 7896 24275 7904
rect 24186 7893 24238 7896
rect 23137 7826 23205 7845
rect 23138 7823 23171 7826
rect 23373 7823 23405 7824
rect 22548 7762 22751 7775
rect 22548 7729 22572 7762
rect 22608 7761 22751 7762
rect 22608 7758 22719 7761
rect 22608 7731 22645 7758
rect 22674 7734 22719 7758
rect 22748 7734 22751 7761
rect 22674 7731 22751 7734
rect 22608 7729 22751 7731
rect 22548 7716 22751 7729
rect 22548 7715 22649 7716
rect 22441 7570 22450 7612
rect 22499 7570 22513 7612
rect 22441 7549 22513 7570
rect 22441 7507 22451 7549
rect 22500 7507 22513 7549
rect 22441 7489 22513 7507
rect 22926 7653 22958 7660
rect 22926 7633 22933 7653
rect 22954 7633 22958 7653
rect 22926 7568 22958 7633
rect 23138 7624 23169 7823
rect 23370 7818 23405 7823
rect 23370 7798 23377 7818
rect 23397 7798 23405 7818
rect 23370 7790 23405 7798
rect 23138 7594 23144 7624
rect 23165 7594 23169 7624
rect 23138 7586 23169 7594
rect 23296 7568 23336 7569
rect 22926 7566 23338 7568
rect 22926 7540 23306 7566
rect 23332 7540 23338 7566
rect 22926 7532 23338 7540
rect 22926 7504 22958 7532
rect 23371 7512 23405 7790
rect 23487 7603 23557 7869
rect 24186 7858 24194 7893
rect 24219 7858 24238 7893
rect 24263 7858 24275 7896
rect 24186 7846 24275 7858
rect 24186 7845 24255 7846
rect 24186 7827 24222 7845
rect 23596 7758 23799 7771
rect 23596 7725 23620 7758
rect 23656 7757 23799 7758
rect 23656 7754 23767 7757
rect 23656 7727 23693 7754
rect 23722 7730 23767 7754
rect 23796 7730 23799 7757
rect 23722 7727 23799 7730
rect 23656 7725 23799 7727
rect 23596 7712 23799 7725
rect 23596 7711 23697 7712
rect 22926 7484 22931 7504
rect 22952 7484 22958 7504
rect 22926 7477 22958 7484
rect 23349 7507 23405 7512
rect 23349 7487 23356 7507
rect 23376 7487 23405 7507
rect 23482 7597 23557 7603
rect 23482 7564 23490 7597
rect 23543 7564 23557 7597
rect 23482 7539 23557 7564
rect 23482 7506 23495 7539
rect 23548 7506 23557 7539
rect 23482 7497 23557 7506
rect 23974 7649 24006 7656
rect 23974 7629 23981 7649
rect 24002 7629 24006 7649
rect 23974 7564 24006 7629
rect 24186 7620 24217 7827
rect 24421 7819 24453 7820
rect 24418 7814 24453 7819
rect 24418 7794 24425 7814
rect 24445 7794 24453 7814
rect 24418 7786 24453 7794
rect 24186 7590 24192 7620
rect 24213 7590 24217 7620
rect 24186 7582 24217 7590
rect 24344 7564 24384 7565
rect 23974 7562 24386 7564
rect 23974 7536 24354 7562
rect 24380 7536 24386 7562
rect 23974 7528 24386 7536
rect 23974 7500 24006 7528
rect 24419 7508 24453 7786
rect 24602 7601 24664 7946
rect 24771 7919 24861 7964
rect 24771 7604 24853 7919
rect 24602 7582 24666 7601
rect 24602 7543 24615 7582
rect 24649 7543 24666 7582
rect 24602 7524 24666 7543
rect 24771 7563 24792 7604
rect 24828 7563 24853 7604
rect 24771 7534 24853 7563
rect 23482 7492 23540 7497
rect 23349 7480 23405 7487
rect 23974 7480 23979 7500
rect 24000 7480 24006 7500
rect 23349 7479 23384 7480
rect 23974 7473 24006 7480
rect 24397 7503 24453 7508
rect 24397 7483 24404 7503
rect 24424 7483 24453 7503
rect 24397 7476 24453 7483
rect 24397 7475 24432 7476
rect 22640 7424 22751 7428
rect 24423 7424 25993 7425
rect 21962 7406 25993 7424
rect 21962 7386 22648 7406
rect 22667 7386 22725 7406
rect 22744 7402 25993 7406
rect 22744 7386 23696 7402
rect 21962 7382 23696 7386
rect 23715 7382 23773 7402
rect 23792 7382 25993 7402
rect 21962 7368 25993 7382
rect 21962 6745 22069 7368
rect 23688 7365 23799 7368
rect 22448 7319 22512 7323
rect 22444 7313 22512 7319
rect 22444 7280 22461 7313
rect 22501 7280 22512 7313
rect 22444 7268 22512 7280
rect 23495 7282 23560 7304
rect 22444 7266 22501 7268
rect 22448 6905 22499 7266
rect 23495 7243 23512 7282
rect 23557 7243 23560 7282
rect 23136 7198 23171 7200
rect 23136 7189 23240 7198
rect 23136 7188 23187 7189
rect 23136 7168 23139 7188
rect 23164 7169 23187 7188
rect 23219 7169 23240 7189
rect 23164 7168 23240 7169
rect 23136 7161 23240 7168
rect 23136 7149 23171 7161
rect 22548 7083 22751 7096
rect 22548 7050 22572 7083
rect 22608 7082 22751 7083
rect 22608 7079 22719 7082
rect 22608 7052 22645 7079
rect 22674 7055 22719 7079
rect 22748 7055 22751 7082
rect 22674 7052 22751 7055
rect 22608 7050 22751 7052
rect 22548 7037 22751 7050
rect 22548 7036 22649 7037
rect 22926 6974 22958 6981
rect 22926 6954 22933 6974
rect 22954 6954 22958 6974
rect 22437 6896 22502 6905
rect 22437 6859 22447 6896
rect 22487 6862 22502 6896
rect 22926 6889 22958 6954
rect 23138 6945 23169 7149
rect 23373 7144 23405 7145
rect 23370 7139 23405 7144
rect 23370 7119 23377 7139
rect 23397 7119 23405 7139
rect 23370 7111 23405 7119
rect 23138 6915 23144 6945
rect 23165 6915 23169 6945
rect 23138 6907 23169 6915
rect 23296 6889 23336 6890
rect 22926 6887 23338 6889
rect 22487 6859 22504 6862
rect 22437 6840 22504 6859
rect 22437 6819 22451 6840
rect 22487 6819 22504 6840
rect 22437 6812 22504 6819
rect 22926 6861 23306 6887
rect 23332 6861 23338 6887
rect 22926 6853 23338 6861
rect 22926 6825 22958 6853
rect 23371 6833 23405 7111
rect 23495 6943 23560 7243
rect 24766 7267 24859 7282
rect 24766 7223 24781 7267
rect 24841 7223 24859 7267
rect 22926 6805 22931 6825
rect 22952 6805 22958 6825
rect 22926 6798 22958 6805
rect 23349 6828 23405 6833
rect 23349 6808 23356 6828
rect 23376 6808 23405 6828
rect 23349 6801 23405 6808
rect 23485 6932 23565 6943
rect 23485 6906 23502 6932
rect 23542 6906 23565 6932
rect 23485 6879 23565 6906
rect 23485 6853 23506 6879
rect 23546 6853 23565 6879
rect 23485 6834 23565 6853
rect 23485 6808 23509 6834
rect 23549 6808 23565 6834
rect 23349 6800 23384 6801
rect 23485 6796 23565 6808
rect 24766 6850 24859 7223
rect 25043 7078 25246 7091
rect 25043 7045 25067 7078
rect 25103 7077 25246 7078
rect 25103 7074 25214 7077
rect 25103 7047 25140 7074
rect 25169 7050 25214 7074
rect 25243 7050 25246 7077
rect 25169 7047 25246 7050
rect 25103 7045 25246 7047
rect 25043 7032 25246 7045
rect 25043 7031 25144 7032
rect 24766 6809 24781 6850
rect 24835 6809 24859 6850
rect 24766 6802 24859 6809
rect 25421 6969 25453 6976
rect 25421 6949 25428 6969
rect 25449 6949 25453 6969
rect 25421 6884 25453 6949
rect 25633 6940 25664 7141
rect 25868 7139 25900 7140
rect 25865 7134 25900 7139
rect 25865 7114 25872 7134
rect 25892 7114 25900 7134
rect 25865 7106 25900 7114
rect 25633 6910 25639 6940
rect 25660 6910 25664 6940
rect 25633 6902 25664 6910
rect 25791 6884 25831 6885
rect 25421 6882 25833 6884
rect 25421 6856 25801 6882
rect 25827 6856 25833 6882
rect 25421 6848 25833 6856
rect 25421 6820 25453 6848
rect 25866 6828 25900 7106
rect 25421 6800 25426 6820
rect 25447 6800 25453 6820
rect 25421 6793 25453 6800
rect 25844 6823 25900 6828
rect 25844 6803 25851 6823
rect 25871 6803 25900 6823
rect 25844 6796 25900 6803
rect 25844 6795 25879 6796
rect 22640 6745 22751 6749
rect 24382 6745 26026 6748
rect 21960 6727 26026 6745
rect 21960 6707 22648 6727
rect 22667 6707 22725 6727
rect 22744 6722 26026 6727
rect 22744 6707 25143 6722
rect 21960 6702 25143 6707
rect 25162 6702 25220 6722
rect 25239 6702 26026 6722
rect 21960 6692 26026 6702
rect 21960 6689 22585 6692
rect 22772 6689 26026 6692
rect 19977 6531 19999 6569
rect 20024 6534 20043 6569
rect 20068 6534 20076 6569
rect 20024 6531 20076 6534
rect 19977 6523 20076 6531
rect 20003 6522 20075 6523
rect 19654 6496 19725 6512
rect 19654 6480 19674 6496
rect 19655 6450 19674 6480
rect 19657 6430 19674 6450
rect 19704 6450 19725 6496
rect 20697 6492 20775 6573
rect 21142 6518 21250 6573
rect 19704 6430 19724 6450
rect 19657 6411 19724 6430
rect 20697 6390 20776 6492
rect 20661 6372 20782 6390
rect 20661 6370 20732 6372
rect 20661 6329 20676 6370
rect 20713 6331 20732 6370
rect 20769 6331 20782 6372
rect 20713 6329 20782 6331
rect 20661 6319 20782 6329
rect 17966 6291 18077 6294
rect 17280 6290 18830 6291
rect 21143 6290 21250 6518
rect 21962 6461 22069 6689
rect 24382 6688 26026 6689
rect 25135 6685 25246 6688
rect 22430 6650 22551 6660
rect 22430 6648 22499 6650
rect 22430 6607 22443 6648
rect 22480 6609 22499 6648
rect 22536 6609 22551 6650
rect 22480 6607 22551 6609
rect 22430 6589 22551 6607
rect 25635 6630 25721 6634
rect 25635 6612 25650 6630
rect 25702 6612 25721 6630
rect 25635 6603 25721 6612
rect 22436 6487 22515 6589
rect 23488 6549 23555 6568
rect 23488 6529 23508 6549
rect 21962 6406 22070 6461
rect 22437 6406 22515 6487
rect 23487 6483 23508 6529
rect 23538 6529 23555 6549
rect 23538 6499 23557 6529
rect 23538 6483 23558 6499
rect 23487 6467 23558 6483
rect 23137 6456 23209 6457
rect 23136 6448 23235 6456
rect 23136 6445 23188 6448
rect 23136 6410 23144 6445
rect 23169 6410 23188 6445
rect 23213 6410 23235 6448
rect 17280 6287 20440 6290
rect 20627 6287 21252 6290
rect 17280 6277 21252 6287
rect 17280 6257 17973 6277
rect 17992 6257 18050 6277
rect 18069 6272 21252 6277
rect 18069 6257 20468 6272
rect 17280 6252 20468 6257
rect 20487 6252 20545 6272
rect 20564 6252 21252 6272
rect 17280 6234 21252 6252
rect 17280 6231 18830 6234
rect 20461 6230 20572 6234
rect 17333 6183 17368 6184
rect 17312 6176 17368 6183
rect 17312 6156 17341 6176
rect 17361 6156 17368 6176
rect 17312 6151 17368 6156
rect 17759 6179 17791 6186
rect 17759 6159 17765 6179
rect 17786 6159 17791 6179
rect 17312 5873 17346 6151
rect 17759 6131 17791 6159
rect 19647 6171 19727 6183
rect 19828 6178 19863 6179
rect 17379 6123 17791 6131
rect 17379 6097 17385 6123
rect 17411 6097 17791 6123
rect 18177 6137 18614 6150
rect 18177 6114 18190 6137
rect 18216 6130 18614 6137
rect 18216 6114 18570 6130
rect 18177 6107 18570 6114
rect 18596 6107 18614 6130
rect 18177 6101 18614 6107
rect 19647 6145 19663 6171
rect 19703 6145 19727 6171
rect 19647 6126 19727 6145
rect 17379 6095 17791 6097
rect 17381 6094 17421 6095
rect 17548 6069 17579 6077
rect 17548 6039 17552 6069
rect 17573 6039 17579 6069
rect 17312 5865 17347 5873
rect 17312 5845 17320 5865
rect 17340 5845 17347 5865
rect 17312 5840 17347 5845
rect 17312 5839 17344 5840
rect 17548 5832 17579 6039
rect 17759 6030 17791 6095
rect 19647 6100 19666 6126
rect 19706 6100 19727 6126
rect 19647 6073 19727 6100
rect 19647 6047 19670 6073
rect 19710 6047 19727 6073
rect 19647 6036 19727 6047
rect 19807 6171 19863 6178
rect 19807 6151 19836 6171
rect 19856 6151 19863 6171
rect 19807 6146 19863 6151
rect 20254 6174 20286 6181
rect 20254 6154 20260 6174
rect 20281 6154 20286 6174
rect 17759 6010 17763 6030
rect 17784 6010 17791 6030
rect 17759 6003 17791 6010
rect 18068 5947 18169 5948
rect 17966 5934 18169 5947
rect 17966 5932 18109 5934
rect 17966 5929 18043 5932
rect 17966 5902 17969 5929
rect 17998 5905 18043 5929
rect 18072 5905 18109 5932
rect 17998 5902 18109 5905
rect 17966 5901 18109 5902
rect 18145 5901 18169 5934
rect 17966 5888 18169 5901
rect 17546 5826 17579 5832
rect 17542 5822 17579 5826
rect 17542 5812 17580 5822
rect 17542 5799 17552 5812
rect 17543 5775 17552 5799
rect 17569 5775 17580 5812
rect 17543 5754 17580 5775
rect 19652 5736 19717 6036
rect 19807 5868 19841 6146
rect 20254 6126 20286 6154
rect 19874 6118 20286 6126
rect 19874 6092 19880 6118
rect 19906 6092 20286 6118
rect 20708 6160 20775 6167
rect 20708 6139 20725 6160
rect 20761 6139 20775 6160
rect 20708 6120 20775 6139
rect 20708 6117 20725 6120
rect 19874 6090 20286 6092
rect 19876 6089 19916 6090
rect 20043 6064 20074 6072
rect 20043 6034 20047 6064
rect 20068 6034 20074 6064
rect 19807 5860 19842 5868
rect 19807 5840 19815 5860
rect 19835 5840 19842 5860
rect 19807 5835 19842 5840
rect 19807 5834 19839 5835
rect 20043 5830 20074 6034
rect 20254 6025 20286 6090
rect 20710 6083 20725 6117
rect 20765 6083 20775 6120
rect 20710 6074 20775 6083
rect 20254 6005 20258 6025
rect 20279 6005 20286 6025
rect 20254 5998 20286 6005
rect 20563 5942 20664 5943
rect 20461 5929 20664 5942
rect 20461 5927 20604 5929
rect 20461 5924 20538 5927
rect 20461 5897 20464 5924
rect 20493 5900 20538 5924
rect 20567 5900 20604 5927
rect 20493 5897 20604 5900
rect 20461 5896 20604 5897
rect 20640 5896 20664 5929
rect 20461 5883 20664 5896
rect 20041 5818 20076 5830
rect 19972 5811 20076 5818
rect 19972 5810 20048 5811
rect 19972 5790 19993 5810
rect 20025 5791 20048 5810
rect 20073 5791 20076 5811
rect 20025 5790 20076 5791
rect 19972 5781 20076 5790
rect 20041 5779 20076 5781
rect 19652 5697 19655 5736
rect 19700 5697 19717 5736
rect 20713 5713 20764 6074
rect 20711 5711 20768 5713
rect 19652 5675 19717 5697
rect 20700 5699 20768 5711
rect 20700 5666 20711 5699
rect 20751 5666 20768 5699
rect 20700 5660 20768 5666
rect 20700 5656 20764 5660
rect 19413 5611 19524 5614
rect 21143 5611 21250 6234
rect 17489 5597 21250 5611
rect 17489 5577 19420 5597
rect 19439 5577 19497 5597
rect 19516 5593 21250 5597
rect 19516 5577 20468 5593
rect 17489 5573 20468 5577
rect 20487 5573 20545 5593
rect 20564 5573 21250 5593
rect 17489 5555 21250 5573
rect 17489 5554 18789 5555
rect 20461 5551 20572 5555
rect 18780 5503 18815 5504
rect 18759 5496 18815 5503
rect 18759 5476 18788 5496
rect 18808 5476 18815 5496
rect 18759 5471 18815 5476
rect 19206 5499 19238 5506
rect 19828 5499 19863 5500
rect 19206 5479 19212 5499
rect 19233 5479 19238 5499
rect 19807 5492 19863 5499
rect 19672 5482 19730 5487
rect 18759 5193 18793 5471
rect 19206 5451 19238 5479
rect 18826 5443 19238 5451
rect 18826 5417 18832 5443
rect 18858 5417 19238 5443
rect 18826 5415 19238 5417
rect 18828 5414 18868 5415
rect 18995 5389 19026 5397
rect 18995 5359 18999 5389
rect 19020 5359 19026 5389
rect 18759 5185 18794 5193
rect 18759 5165 18767 5185
rect 18787 5165 18794 5185
rect 18759 5160 18794 5165
rect 18759 5159 18791 5160
rect 18995 5152 19026 5359
rect 19206 5350 19238 5415
rect 19206 5330 19210 5350
rect 19231 5330 19238 5350
rect 19206 5323 19238 5330
rect 19655 5473 19730 5482
rect 19655 5440 19664 5473
rect 19717 5440 19730 5473
rect 19655 5415 19730 5440
rect 19655 5382 19669 5415
rect 19722 5382 19730 5415
rect 19655 5376 19730 5382
rect 19807 5472 19836 5492
rect 19856 5472 19863 5492
rect 19807 5467 19863 5472
rect 20254 5495 20286 5502
rect 20254 5475 20260 5495
rect 20281 5475 20286 5495
rect 19515 5267 19616 5268
rect 19413 5254 19616 5267
rect 19413 5252 19556 5254
rect 19413 5249 19490 5252
rect 19413 5222 19416 5249
rect 19445 5225 19490 5249
rect 19519 5225 19556 5252
rect 19445 5222 19556 5225
rect 19413 5221 19556 5222
rect 19592 5221 19616 5254
rect 19413 5208 19616 5221
rect 18493 5139 18657 5142
rect 18990 5139 19026 5152
rect 17692 5121 19031 5139
rect 17692 5083 17702 5121
rect 17727 5106 19031 5121
rect 17727 5083 17737 5106
rect 18493 5099 18657 5106
rect 17692 5075 17737 5083
rect 17706 5074 17737 5075
rect 19655 5060 19725 5376
rect 19807 5189 19841 5467
rect 20254 5447 20286 5475
rect 19874 5439 20286 5447
rect 19874 5413 19880 5439
rect 19906 5413 20286 5439
rect 19874 5411 20286 5413
rect 19876 5410 19916 5411
rect 20043 5385 20074 5393
rect 20043 5355 20047 5385
rect 20068 5355 20074 5385
rect 19807 5181 19842 5189
rect 19807 5161 19815 5181
rect 19835 5161 19842 5181
rect 19807 5156 19842 5161
rect 20043 5156 20074 5355
rect 20254 5346 20286 5411
rect 20254 5326 20258 5346
rect 20279 5326 20286 5346
rect 20254 5319 20286 5326
rect 20699 5472 20771 5490
rect 20699 5430 20712 5472
rect 20761 5430 20771 5472
rect 20699 5409 20771 5430
rect 20699 5367 20713 5409
rect 20762 5367 20771 5409
rect 20563 5263 20664 5264
rect 20461 5250 20664 5263
rect 20461 5248 20604 5250
rect 20461 5245 20538 5248
rect 20461 5218 20464 5245
rect 20493 5221 20538 5245
rect 20567 5221 20604 5248
rect 20493 5218 20604 5221
rect 20461 5217 20604 5218
rect 20640 5217 20664 5250
rect 20461 5204 20664 5217
rect 19807 5155 19839 5156
rect 20041 5153 20074 5156
rect 20007 5134 20075 5153
rect 19977 5122 20076 5134
rect 19977 5084 19999 5122
rect 20024 5087 20043 5122
rect 20068 5087 20076 5122
rect 20024 5084 20076 5087
rect 19977 5076 20076 5084
rect 20003 5075 20075 5076
rect 19655 5041 19734 5060
rect 19658 5021 19734 5041
rect 19651 4997 19734 5021
rect 20699 5056 20771 5367
rect 20699 5013 20775 5056
rect 19651 4931 19663 4997
rect 19717 4931 19734 4997
rect 19651 4911 19734 4931
rect 19651 4874 19668 4911
rect 19712 4897 19734 4911
rect 20700 4962 20775 5013
rect 21143 4962 21250 5555
rect 21962 5977 22069 6406
rect 22441 6165 22513 6406
rect 23136 6398 23235 6410
rect 23137 6379 23205 6398
rect 23138 6376 23171 6379
rect 23373 6376 23405 6377
rect 22548 6315 22751 6328
rect 22548 6282 22572 6315
rect 22608 6314 22751 6315
rect 22608 6311 22719 6314
rect 22608 6284 22645 6311
rect 22674 6287 22719 6311
rect 22748 6287 22751 6314
rect 22674 6284 22751 6287
rect 22608 6282 22751 6284
rect 22548 6269 22751 6282
rect 22548 6268 22649 6269
rect 22441 6123 22450 6165
rect 22499 6123 22513 6165
rect 22441 6102 22513 6123
rect 22441 6060 22451 6102
rect 22500 6060 22513 6102
rect 22441 6042 22513 6060
rect 22926 6206 22958 6213
rect 22926 6186 22933 6206
rect 22954 6186 22958 6206
rect 22926 6121 22958 6186
rect 23138 6177 23169 6376
rect 23370 6371 23405 6376
rect 23370 6351 23377 6371
rect 23397 6351 23405 6371
rect 23370 6343 23405 6351
rect 23138 6147 23144 6177
rect 23165 6147 23169 6177
rect 23138 6139 23169 6147
rect 23296 6121 23336 6122
rect 22926 6119 23338 6121
rect 22926 6093 23306 6119
rect 23332 6093 23338 6119
rect 22926 6085 23338 6093
rect 22926 6057 22958 6085
rect 23371 6065 23405 6343
rect 23487 6156 23557 6467
rect 25412 6457 25484 6458
rect 25411 6454 25500 6457
rect 24183 6452 25500 6454
rect 24180 6449 25500 6452
rect 24180 6446 25463 6449
rect 24180 6411 25419 6446
rect 25444 6411 25463 6446
rect 25488 6411 25500 6449
rect 24180 6401 25500 6411
rect 25676 6450 25712 6603
rect 25676 6427 25682 6450
rect 25706 6427 25712 6450
rect 25676 6406 25712 6427
rect 24180 6399 25465 6401
rect 24180 6389 24277 6399
rect 24186 6380 24222 6389
rect 25676 6383 25682 6406
rect 25706 6383 25712 6406
rect 23596 6311 23799 6324
rect 23596 6278 23620 6311
rect 23656 6310 23799 6311
rect 23656 6307 23767 6310
rect 23656 6280 23693 6307
rect 23722 6283 23767 6307
rect 23796 6283 23799 6310
rect 23722 6280 23799 6283
rect 23656 6278 23799 6280
rect 23596 6265 23799 6278
rect 23596 6264 23697 6265
rect 22926 6037 22931 6057
rect 22952 6037 22958 6057
rect 22926 6030 22958 6037
rect 23349 6060 23405 6065
rect 23349 6040 23356 6060
rect 23376 6040 23405 6060
rect 23482 6150 23557 6156
rect 23482 6117 23490 6150
rect 23543 6117 23557 6150
rect 23482 6092 23557 6117
rect 23482 6059 23495 6092
rect 23548 6059 23557 6092
rect 23482 6050 23557 6059
rect 23974 6202 24006 6209
rect 23974 6182 23981 6202
rect 24002 6182 24006 6202
rect 23974 6117 24006 6182
rect 24186 6173 24217 6380
rect 24421 6372 24453 6373
rect 25676 6372 25712 6383
rect 24418 6367 24453 6372
rect 24418 6347 24425 6367
rect 24445 6347 24453 6367
rect 24418 6339 24453 6347
rect 24186 6143 24192 6173
rect 24213 6143 24217 6173
rect 24186 6135 24217 6143
rect 24344 6117 24384 6118
rect 23974 6115 24386 6117
rect 23974 6089 24354 6115
rect 24380 6089 24386 6115
rect 23974 6081 24386 6089
rect 23974 6053 24006 6081
rect 24419 6061 24453 6339
rect 23482 6045 23540 6050
rect 23349 6033 23405 6040
rect 23974 6033 23979 6053
rect 24000 6033 24006 6053
rect 23349 6032 23384 6033
rect 23974 6026 24006 6033
rect 24397 6056 24453 6061
rect 24397 6036 24404 6056
rect 24424 6036 24453 6056
rect 24397 6029 24453 6036
rect 24397 6028 24432 6029
rect 22640 5977 22751 5981
rect 24515 5977 25674 5978
rect 21962 5959 25674 5977
rect 21962 5939 22648 5959
rect 22667 5939 22725 5959
rect 22744 5955 25674 5959
rect 22744 5939 23696 5955
rect 21962 5935 23696 5939
rect 23715 5935 23773 5955
rect 23792 5935 25674 5955
rect 21962 5921 25674 5935
rect 21962 5298 22069 5921
rect 23688 5918 23799 5921
rect 22448 5872 22512 5876
rect 22444 5866 22512 5872
rect 22444 5833 22461 5866
rect 22501 5833 22512 5866
rect 22444 5821 22512 5833
rect 23495 5835 23560 5857
rect 22444 5819 22501 5821
rect 22448 5458 22499 5819
rect 23495 5796 23512 5835
rect 23557 5796 23560 5835
rect 26581 5833 26633 8139
rect 26742 8116 26777 8182
rect 26742 6800 26776 8116
rect 27080 7969 27185 13104
rect 30380 13070 30491 13073
rect 32110 13070 32217 13685
rect 29633 13056 32217 13070
rect 29633 13036 30387 13056
rect 30406 13036 30464 13056
rect 30483 13052 32217 13056
rect 30483 13036 31435 13052
rect 29633 13032 31435 13036
rect 31454 13032 31512 13052
rect 31531 13032 32217 13052
rect 29633 13014 32217 13032
rect 29633 13013 29664 13014
rect 31428 13010 31539 13014
rect 29747 12962 29782 12963
rect 29726 12955 29782 12962
rect 29726 12935 29755 12955
rect 29775 12935 29782 12955
rect 29726 12930 29782 12935
rect 30173 12958 30205 12965
rect 30795 12958 30830 12959
rect 30173 12938 30179 12958
rect 30200 12938 30205 12958
rect 30774 12951 30830 12958
rect 30639 12941 30697 12946
rect 29726 12652 29760 12930
rect 30173 12910 30205 12938
rect 29793 12902 30205 12910
rect 29793 12876 29799 12902
rect 29825 12876 30205 12902
rect 29793 12874 30205 12876
rect 29795 12873 29835 12874
rect 29962 12848 29993 12856
rect 29962 12818 29966 12848
rect 29987 12818 29993 12848
rect 29726 12644 29761 12652
rect 29726 12624 29734 12644
rect 29754 12624 29761 12644
rect 29726 12619 29761 12624
rect 29726 12618 29758 12619
rect 29962 12618 29993 12818
rect 30173 12809 30205 12874
rect 30173 12789 30177 12809
rect 30198 12789 30205 12809
rect 30173 12782 30205 12789
rect 30622 12932 30697 12941
rect 30622 12899 30631 12932
rect 30684 12899 30697 12932
rect 30622 12874 30697 12899
rect 30622 12841 30636 12874
rect 30689 12841 30697 12874
rect 30622 12835 30697 12841
rect 30774 12931 30803 12951
rect 30823 12931 30830 12951
rect 30774 12926 30830 12931
rect 31221 12954 31253 12961
rect 31221 12934 31227 12954
rect 31248 12934 31253 12954
rect 30482 12726 30583 12727
rect 30380 12713 30583 12726
rect 30380 12711 30523 12713
rect 30380 12708 30457 12711
rect 30380 12681 30383 12708
rect 30412 12684 30457 12708
rect 30486 12684 30523 12711
rect 30412 12681 30523 12684
rect 30380 12680 30523 12681
rect 30559 12680 30583 12713
rect 30380 12667 30583 12680
rect 29959 12611 29998 12618
rect 29957 12594 29998 12611
rect 29959 12569 29998 12594
rect 28653 12561 29998 12569
rect 28653 12533 28668 12561
rect 28696 12535 29998 12561
rect 28696 12533 29995 12535
rect 28653 12528 29995 12533
rect 30622 12524 30692 12835
rect 30774 12648 30808 12926
rect 31221 12906 31253 12934
rect 30841 12898 31253 12906
rect 30841 12872 30847 12898
rect 30873 12872 31253 12898
rect 30841 12870 31253 12872
rect 30843 12869 30883 12870
rect 31010 12844 31041 12852
rect 31010 12814 31014 12844
rect 31035 12814 31041 12844
rect 30774 12640 30809 12648
rect 30774 12620 30782 12640
rect 30802 12620 30809 12640
rect 30774 12615 30809 12620
rect 31010 12615 31041 12814
rect 31221 12805 31253 12870
rect 31221 12785 31225 12805
rect 31246 12785 31253 12805
rect 31221 12778 31253 12785
rect 31666 12931 31738 12949
rect 31666 12889 31679 12931
rect 31728 12889 31738 12931
rect 31666 12868 31738 12889
rect 31666 12826 31680 12868
rect 31729 12826 31738 12868
rect 31530 12722 31631 12723
rect 31428 12709 31631 12722
rect 31428 12707 31571 12709
rect 31428 12704 31505 12707
rect 31428 12677 31431 12704
rect 31460 12680 31505 12704
rect 31534 12680 31571 12707
rect 31460 12677 31571 12680
rect 31428 12676 31571 12677
rect 31607 12676 31631 12709
rect 31428 12663 31631 12676
rect 30774 12614 30806 12615
rect 31008 12612 31041 12615
rect 30974 12593 31042 12612
rect 30944 12581 31043 12593
rect 31666 12585 31738 12826
rect 32110 12585 32217 13014
rect 32672 13426 32779 13685
rect 33151 13614 33223 13915
rect 33847 13905 33919 13906
rect 33846 13897 33945 13905
rect 33846 13894 33898 13897
rect 33846 13859 33854 13894
rect 33879 13859 33898 13894
rect 33923 13859 33945 13897
rect 33846 13847 33945 13859
rect 33847 13828 33915 13847
rect 33848 13825 33881 13828
rect 34083 13825 34115 13826
rect 33258 13764 33461 13777
rect 33258 13731 33282 13764
rect 33318 13763 33461 13764
rect 33318 13760 33429 13763
rect 33318 13733 33355 13760
rect 33384 13736 33429 13760
rect 33458 13736 33461 13763
rect 33384 13733 33461 13736
rect 33318 13731 33461 13733
rect 33258 13718 33461 13731
rect 33258 13717 33359 13718
rect 33151 13572 33160 13614
rect 33209 13572 33223 13614
rect 33151 13551 33223 13572
rect 33151 13509 33161 13551
rect 33210 13509 33223 13551
rect 33151 13491 33223 13509
rect 33636 13655 33668 13662
rect 33636 13635 33643 13655
rect 33664 13635 33668 13655
rect 33636 13570 33668 13635
rect 33848 13626 33879 13825
rect 34080 13820 34115 13825
rect 34080 13800 34087 13820
rect 34107 13800 34115 13820
rect 34080 13792 34115 13800
rect 33848 13596 33854 13626
rect 33875 13596 33879 13626
rect 33848 13588 33879 13596
rect 34006 13570 34046 13571
rect 33636 13568 34048 13570
rect 33636 13542 34016 13568
rect 34042 13542 34048 13568
rect 33636 13534 34048 13542
rect 33636 13506 33668 13534
rect 34081 13514 34115 13792
rect 34197 13605 34267 13905
rect 34896 13898 34985 13905
rect 34896 13895 34948 13898
rect 34896 13860 34904 13895
rect 34929 13860 34948 13895
rect 34973 13860 34985 13898
rect 34896 13848 34985 13860
rect 34896 13847 34965 13848
rect 34896 13829 34932 13847
rect 34306 13760 34509 13773
rect 34306 13727 34330 13760
rect 34366 13759 34509 13760
rect 34366 13756 34477 13759
rect 34366 13729 34403 13756
rect 34432 13732 34477 13756
rect 34506 13732 34509 13759
rect 34432 13729 34509 13732
rect 34366 13727 34509 13729
rect 34306 13714 34509 13727
rect 34306 13713 34407 13714
rect 33636 13486 33641 13506
rect 33662 13486 33668 13506
rect 33636 13479 33668 13486
rect 34059 13509 34115 13514
rect 34059 13489 34066 13509
rect 34086 13489 34115 13509
rect 34192 13599 34267 13605
rect 34192 13566 34200 13599
rect 34253 13566 34267 13599
rect 34192 13541 34267 13566
rect 34192 13508 34205 13541
rect 34258 13508 34267 13541
rect 34192 13499 34267 13508
rect 34684 13651 34716 13658
rect 34684 13631 34691 13651
rect 34712 13631 34716 13651
rect 34684 13566 34716 13631
rect 34896 13622 34927 13829
rect 35131 13821 35163 13822
rect 35128 13816 35163 13821
rect 35128 13796 35135 13816
rect 35155 13796 35163 13816
rect 35128 13788 35163 13796
rect 34896 13592 34902 13622
rect 34923 13592 34927 13622
rect 34896 13584 34927 13592
rect 35054 13566 35094 13567
rect 34684 13564 35096 13566
rect 34684 13538 35064 13564
rect 35090 13538 35096 13564
rect 34684 13530 35096 13538
rect 34684 13502 34716 13530
rect 35129 13510 35163 13788
rect 35312 13603 35374 13905
rect 35481 13606 35563 13962
rect 36748 13802 36797 14089
rect 36748 13770 36917 13802
rect 36748 13764 36863 13770
rect 36748 13755 36803 13764
rect 36738 13667 36803 13755
rect 36841 13673 36863 13764
rect 36901 13673 36917 13770
rect 36841 13667 36917 13673
rect 36738 13656 36917 13667
rect 35312 13584 35376 13603
rect 35312 13545 35325 13584
rect 35359 13545 35376 13584
rect 35312 13526 35376 13545
rect 35481 13565 35502 13606
rect 35538 13565 35563 13606
rect 35481 13536 35563 13565
rect 36748 13651 36917 13656
rect 34192 13494 34250 13499
rect 34059 13482 34115 13489
rect 34684 13482 34689 13502
rect 34710 13482 34716 13502
rect 34059 13481 34094 13482
rect 34684 13475 34716 13482
rect 35107 13505 35163 13510
rect 35107 13485 35114 13505
rect 35134 13485 35163 13505
rect 35107 13478 35163 13485
rect 35107 13477 35142 13478
rect 33350 13426 33461 13430
rect 35133 13426 36246 13427
rect 32672 13408 36246 13426
rect 32672 13388 33358 13408
rect 33377 13388 33435 13408
rect 33454 13404 36246 13408
rect 33454 13388 34406 13404
rect 32672 13384 34406 13388
rect 34425 13384 34483 13404
rect 34502 13384 36246 13404
rect 32672 13370 36246 13384
rect 32672 12747 32779 13370
rect 34398 13367 34509 13370
rect 33158 13321 33222 13325
rect 33154 13315 33222 13321
rect 33154 13282 33171 13315
rect 33211 13282 33222 13315
rect 33154 13270 33222 13282
rect 34205 13284 34270 13306
rect 33154 13268 33211 13270
rect 33158 12907 33209 13268
rect 34205 13245 34222 13284
rect 34267 13245 34270 13284
rect 33846 13200 33881 13202
rect 33846 13191 33950 13200
rect 33846 13190 33897 13191
rect 33846 13170 33849 13190
rect 33874 13171 33897 13190
rect 33929 13171 33950 13191
rect 33874 13170 33950 13171
rect 33846 13163 33950 13170
rect 33846 13151 33881 13163
rect 33258 13085 33461 13098
rect 33258 13052 33282 13085
rect 33318 13084 33461 13085
rect 33318 13081 33429 13084
rect 33318 13054 33355 13081
rect 33384 13057 33429 13081
rect 33458 13057 33461 13084
rect 33384 13054 33461 13057
rect 33318 13052 33461 13054
rect 33258 13039 33461 13052
rect 33258 13038 33359 13039
rect 33636 12976 33668 12983
rect 33636 12956 33643 12976
rect 33664 12956 33668 12976
rect 33147 12898 33212 12907
rect 33147 12861 33157 12898
rect 33197 12864 33212 12898
rect 33636 12891 33668 12956
rect 33848 12947 33879 13151
rect 34083 13146 34115 13147
rect 34080 13141 34115 13146
rect 34080 13121 34087 13141
rect 34107 13121 34115 13141
rect 34080 13113 34115 13121
rect 33848 12917 33854 12947
rect 33875 12917 33879 12947
rect 33848 12909 33879 12917
rect 34006 12891 34046 12892
rect 33636 12889 34048 12891
rect 33197 12861 33214 12864
rect 33147 12842 33214 12861
rect 33147 12821 33161 12842
rect 33197 12821 33214 12842
rect 33147 12814 33214 12821
rect 33636 12863 34016 12889
rect 34042 12863 34048 12889
rect 33636 12855 34048 12863
rect 33636 12827 33668 12855
rect 34081 12835 34115 13113
rect 34205 12945 34270 13245
rect 35476 13269 35569 13284
rect 35476 13225 35491 13269
rect 35551 13225 35569 13269
rect 33636 12807 33641 12827
rect 33662 12807 33668 12827
rect 33636 12800 33668 12807
rect 34059 12830 34115 12835
rect 34059 12810 34066 12830
rect 34086 12810 34115 12830
rect 34059 12803 34115 12810
rect 34195 12934 34275 12945
rect 34195 12908 34212 12934
rect 34252 12908 34275 12934
rect 34195 12881 34275 12908
rect 34195 12855 34216 12881
rect 34256 12855 34275 12881
rect 34195 12836 34275 12855
rect 34195 12810 34219 12836
rect 34259 12810 34275 12836
rect 34059 12802 34094 12803
rect 34195 12798 34275 12810
rect 35476 12852 35569 13225
rect 35753 13080 35956 13093
rect 35753 13047 35777 13080
rect 35813 13079 35956 13080
rect 35813 13076 35924 13079
rect 35813 13049 35850 13076
rect 35879 13052 35924 13076
rect 35953 13052 35956 13079
rect 35879 13049 35956 13052
rect 35813 13047 35956 13049
rect 35753 13034 35956 13047
rect 35753 13033 35854 13034
rect 35476 12811 35491 12852
rect 35545 12811 35569 12852
rect 35476 12804 35569 12811
rect 36131 12971 36163 12978
rect 36131 12951 36138 12971
rect 36159 12951 36163 12971
rect 36131 12886 36163 12951
rect 36343 12942 36374 13143
rect 36578 13141 36610 13142
rect 36575 13136 36610 13141
rect 36575 13116 36582 13136
rect 36602 13116 36610 13136
rect 36575 13108 36610 13116
rect 36343 12912 36349 12942
rect 36370 12912 36374 12942
rect 36343 12904 36374 12912
rect 36501 12886 36541 12887
rect 36131 12884 36543 12886
rect 36131 12858 36511 12884
rect 36537 12858 36543 12884
rect 36131 12850 36543 12858
rect 36131 12822 36163 12850
rect 36576 12830 36610 13108
rect 36131 12802 36136 12822
rect 36157 12802 36163 12822
rect 36131 12795 36163 12802
rect 36554 12825 36610 12830
rect 36554 12805 36561 12825
rect 36581 12805 36610 12825
rect 36554 12798 36610 12805
rect 36554 12797 36589 12798
rect 33350 12747 33461 12751
rect 35092 12747 36641 12750
rect 32670 12729 36641 12747
rect 32670 12709 33358 12729
rect 33377 12709 33435 12729
rect 33454 12724 36641 12729
rect 33454 12709 35853 12724
rect 32670 12704 35853 12709
rect 35872 12704 35930 12724
rect 35949 12704 36641 12724
rect 32670 12694 36641 12704
rect 32670 12691 33295 12694
rect 33482 12691 36641 12694
rect 30944 12543 30966 12581
rect 30991 12546 31010 12581
rect 31035 12546 31043 12581
rect 30991 12543 31043 12546
rect 30944 12535 31043 12543
rect 30970 12534 31042 12535
rect 30621 12508 30692 12524
rect 30621 12492 30641 12508
rect 30622 12462 30641 12492
rect 30624 12442 30641 12462
rect 30671 12462 30692 12508
rect 31664 12504 31742 12585
rect 32109 12530 32217 12585
rect 30671 12442 30691 12462
rect 30624 12423 30691 12442
rect 31664 12402 31743 12504
rect 31628 12384 31749 12402
rect 31628 12382 31699 12384
rect 31628 12341 31643 12382
rect 31680 12343 31699 12382
rect 31736 12343 31749 12384
rect 31680 12341 31749 12343
rect 31628 12331 31749 12341
rect 28933 12303 29044 12306
rect 28144 12302 29797 12303
rect 32110 12302 32217 12530
rect 32672 12463 32779 12691
rect 35092 12690 36641 12691
rect 35845 12687 35956 12690
rect 33140 12652 33261 12662
rect 33140 12650 33209 12652
rect 33140 12609 33153 12650
rect 33190 12611 33209 12650
rect 33246 12611 33261 12652
rect 33190 12609 33261 12611
rect 33140 12591 33261 12609
rect 36345 12632 36431 12636
rect 36345 12614 36360 12632
rect 36412 12614 36431 12632
rect 36345 12605 36431 12614
rect 33146 12489 33225 12591
rect 34198 12551 34265 12570
rect 34198 12531 34218 12551
rect 32672 12408 32780 12463
rect 33147 12408 33225 12489
rect 34197 12485 34218 12531
rect 34248 12531 34265 12551
rect 34248 12501 34267 12531
rect 34248 12485 34268 12501
rect 34197 12469 34268 12485
rect 33847 12458 33919 12459
rect 33846 12450 33945 12458
rect 33846 12447 33898 12450
rect 33846 12412 33854 12447
rect 33879 12412 33898 12447
rect 33923 12412 33945 12450
rect 28144 12299 31407 12302
rect 31594 12299 32219 12302
rect 28144 12289 32219 12299
rect 28144 12269 28940 12289
rect 28959 12269 29017 12289
rect 29036 12284 32219 12289
rect 29036 12269 31435 12284
rect 28144 12264 31435 12269
rect 31454 12264 31512 12284
rect 31531 12264 32219 12284
rect 28144 12246 32219 12264
rect 28144 12243 29797 12246
rect 31428 12242 31539 12246
rect 28300 12195 28335 12196
rect 28279 12188 28335 12195
rect 28279 12168 28308 12188
rect 28328 12168 28335 12188
rect 28279 12163 28335 12168
rect 28726 12191 28758 12198
rect 28726 12171 28732 12191
rect 28753 12171 28758 12191
rect 28279 11885 28313 12163
rect 28726 12143 28758 12171
rect 30614 12183 30694 12195
rect 30795 12190 30830 12191
rect 28346 12135 28758 12143
rect 28346 12109 28352 12135
rect 28378 12109 28758 12135
rect 29144 12149 29581 12162
rect 29144 12126 29157 12149
rect 29183 12142 29581 12149
rect 29183 12126 29537 12142
rect 29144 12119 29537 12126
rect 29563 12119 29581 12142
rect 29144 12113 29581 12119
rect 30614 12157 30630 12183
rect 30670 12157 30694 12183
rect 30614 12138 30694 12157
rect 28346 12107 28758 12109
rect 28348 12106 28388 12107
rect 28515 12081 28546 12089
rect 28515 12051 28519 12081
rect 28540 12051 28546 12081
rect 28279 11877 28314 11885
rect 28279 11857 28287 11877
rect 28307 11857 28314 11877
rect 28279 11852 28314 11857
rect 28279 11851 28311 11852
rect 28515 11844 28546 12051
rect 28726 12042 28758 12107
rect 30614 12112 30633 12138
rect 30673 12112 30694 12138
rect 30614 12085 30694 12112
rect 30614 12059 30637 12085
rect 30677 12059 30694 12085
rect 30614 12048 30694 12059
rect 30774 12183 30830 12190
rect 30774 12163 30803 12183
rect 30823 12163 30830 12183
rect 30774 12158 30830 12163
rect 31221 12186 31253 12193
rect 31221 12166 31227 12186
rect 31248 12166 31253 12186
rect 28726 12022 28730 12042
rect 28751 12022 28758 12042
rect 28726 12015 28758 12022
rect 29035 11959 29136 11960
rect 28933 11946 29136 11959
rect 28933 11944 29076 11946
rect 28933 11941 29010 11944
rect 28933 11914 28936 11941
rect 28965 11917 29010 11941
rect 29039 11917 29076 11944
rect 28965 11914 29076 11917
rect 28933 11913 29076 11914
rect 29112 11913 29136 11946
rect 28933 11900 29136 11913
rect 28513 11838 28546 11844
rect 28509 11834 28546 11838
rect 28509 11824 28547 11834
rect 28509 11811 28519 11824
rect 28510 11787 28519 11811
rect 28536 11787 28547 11824
rect 28510 11766 28547 11787
rect 30619 11748 30684 12048
rect 30774 11880 30808 12158
rect 31221 12138 31253 12166
rect 30841 12130 31253 12138
rect 30841 12104 30847 12130
rect 30873 12104 31253 12130
rect 31675 12172 31742 12179
rect 31675 12151 31692 12172
rect 31728 12151 31742 12172
rect 31675 12132 31742 12151
rect 31675 12129 31692 12132
rect 30841 12102 31253 12104
rect 30843 12101 30883 12102
rect 31010 12076 31041 12084
rect 31010 12046 31014 12076
rect 31035 12046 31041 12076
rect 30774 11872 30809 11880
rect 30774 11852 30782 11872
rect 30802 11852 30809 11872
rect 30774 11847 30809 11852
rect 30774 11846 30806 11847
rect 31010 11842 31041 12046
rect 31221 12037 31253 12102
rect 31677 12095 31692 12129
rect 31732 12095 31742 12132
rect 31677 12086 31742 12095
rect 31221 12017 31225 12037
rect 31246 12017 31253 12037
rect 31221 12010 31253 12017
rect 31530 11954 31631 11955
rect 31428 11941 31631 11954
rect 31428 11939 31571 11941
rect 31428 11936 31505 11939
rect 31428 11909 31431 11936
rect 31460 11912 31505 11936
rect 31534 11912 31571 11939
rect 31460 11909 31571 11912
rect 31428 11908 31571 11909
rect 31607 11908 31631 11941
rect 31428 11895 31631 11908
rect 31008 11830 31043 11842
rect 30939 11823 31043 11830
rect 30939 11822 31015 11823
rect 30939 11802 30960 11822
rect 30992 11803 31015 11822
rect 31040 11803 31043 11823
rect 30992 11802 31043 11803
rect 30939 11793 31043 11802
rect 31008 11791 31043 11793
rect 30619 11709 30622 11748
rect 30667 11709 30684 11748
rect 31680 11725 31731 12086
rect 31678 11723 31735 11725
rect 30619 11687 30684 11709
rect 31667 11711 31735 11723
rect 31667 11678 31678 11711
rect 31718 11678 31735 11711
rect 31667 11672 31735 11678
rect 31667 11668 31731 11672
rect 30380 11623 30491 11626
rect 32110 11623 32217 12246
rect 27767 11609 32217 11623
rect 27767 11589 30387 11609
rect 30406 11589 30464 11609
rect 30483 11605 32217 11609
rect 30483 11589 31435 11605
rect 27767 11585 31435 11589
rect 31454 11585 31512 11605
rect 31531 11585 32217 11605
rect 27767 11571 32217 11585
rect 28186 11567 32217 11571
rect 28186 11566 29756 11567
rect 31428 11563 31539 11567
rect 29747 11515 29782 11516
rect 29726 11508 29782 11515
rect 29726 11488 29755 11508
rect 29775 11488 29782 11508
rect 29726 11483 29782 11488
rect 30173 11511 30205 11518
rect 30795 11511 30830 11512
rect 30173 11491 30179 11511
rect 30200 11491 30205 11511
rect 30774 11504 30830 11511
rect 30639 11494 30697 11499
rect 29726 11205 29760 11483
rect 30173 11463 30205 11491
rect 29793 11455 30205 11463
rect 29793 11429 29799 11455
rect 29825 11429 30205 11455
rect 29793 11427 30205 11429
rect 29795 11426 29835 11427
rect 29962 11401 29993 11409
rect 29962 11371 29966 11401
rect 29987 11371 29993 11401
rect 29726 11197 29761 11205
rect 29726 11177 29734 11197
rect 29754 11177 29761 11197
rect 29726 11172 29761 11177
rect 29726 11171 29758 11172
rect 29962 11164 29993 11371
rect 30173 11362 30205 11427
rect 30173 11342 30177 11362
rect 30198 11342 30205 11362
rect 30173 11335 30205 11342
rect 30622 11485 30697 11494
rect 30622 11452 30631 11485
rect 30684 11452 30697 11485
rect 30622 11427 30697 11452
rect 30622 11394 30636 11427
rect 30689 11394 30697 11427
rect 30622 11388 30697 11394
rect 30774 11484 30803 11504
rect 30823 11484 30830 11504
rect 30774 11479 30830 11484
rect 31221 11507 31253 11514
rect 31221 11487 31227 11507
rect 31248 11487 31253 11507
rect 30482 11279 30583 11280
rect 30380 11266 30583 11279
rect 30380 11264 30523 11266
rect 30380 11261 30457 11264
rect 30380 11234 30383 11261
rect 30412 11237 30457 11261
rect 30486 11237 30523 11264
rect 30412 11234 30523 11237
rect 30380 11233 30523 11234
rect 30559 11233 30583 11266
rect 30380 11220 30583 11233
rect 29460 11151 29624 11154
rect 29957 11151 29993 11164
rect 28659 11133 29998 11151
rect 28659 11095 28669 11133
rect 28694 11118 29998 11133
rect 28694 11095 28704 11118
rect 29460 11111 29624 11118
rect 28659 11087 28704 11095
rect 28673 11086 28704 11087
rect 30622 11072 30692 11388
rect 30774 11201 30808 11479
rect 31221 11459 31253 11487
rect 30841 11451 31253 11459
rect 30841 11425 30847 11451
rect 30873 11425 31253 11451
rect 30841 11423 31253 11425
rect 30843 11422 30883 11423
rect 31010 11397 31041 11405
rect 31010 11367 31014 11397
rect 31035 11367 31041 11397
rect 30774 11193 30809 11201
rect 30774 11173 30782 11193
rect 30802 11173 30809 11193
rect 30774 11168 30809 11173
rect 31010 11168 31041 11367
rect 31221 11358 31253 11423
rect 31221 11338 31225 11358
rect 31246 11338 31253 11358
rect 31221 11331 31253 11338
rect 31666 11484 31738 11502
rect 31666 11442 31679 11484
rect 31728 11442 31738 11484
rect 31666 11421 31738 11442
rect 31666 11379 31680 11421
rect 31729 11379 31738 11421
rect 31530 11275 31631 11276
rect 31428 11262 31631 11275
rect 31428 11260 31571 11262
rect 31428 11257 31505 11260
rect 31428 11230 31431 11257
rect 31460 11233 31505 11257
rect 31534 11233 31571 11260
rect 31460 11230 31571 11233
rect 31428 11229 31571 11230
rect 31607 11229 31631 11262
rect 31428 11216 31631 11229
rect 30774 11167 30806 11168
rect 31008 11165 31041 11168
rect 30974 11146 31042 11165
rect 30944 11134 31043 11146
rect 30944 11096 30966 11134
rect 30991 11099 31010 11134
rect 31035 11099 31043 11134
rect 30991 11096 31043 11099
rect 30944 11088 31043 11096
rect 30970 11087 31042 11088
rect 30622 11053 30701 11072
rect 30625 11033 30701 11053
rect 30618 11009 30701 11033
rect 31666 11068 31738 11379
rect 31666 11025 31742 11068
rect 30618 10943 30630 11009
rect 30684 10943 30701 11009
rect 30618 10923 30701 10943
rect 30618 10886 30635 10923
rect 30679 10909 30701 10923
rect 31667 10974 31742 11025
rect 32110 10974 32217 11567
rect 32672 11979 32779 12408
rect 33151 12167 33223 12408
rect 33846 12400 33945 12412
rect 33847 12381 33915 12400
rect 33848 12378 33881 12381
rect 34083 12378 34115 12379
rect 33258 12317 33461 12330
rect 33258 12284 33282 12317
rect 33318 12316 33461 12317
rect 33318 12313 33429 12316
rect 33318 12286 33355 12313
rect 33384 12289 33429 12313
rect 33458 12289 33461 12316
rect 33384 12286 33461 12289
rect 33318 12284 33461 12286
rect 33258 12271 33461 12284
rect 33258 12270 33359 12271
rect 33151 12125 33160 12167
rect 33209 12125 33223 12167
rect 33151 12104 33223 12125
rect 33151 12062 33161 12104
rect 33210 12062 33223 12104
rect 33151 12044 33223 12062
rect 33636 12208 33668 12215
rect 33636 12188 33643 12208
rect 33664 12188 33668 12208
rect 33636 12123 33668 12188
rect 33848 12179 33879 12378
rect 34080 12373 34115 12378
rect 34080 12353 34087 12373
rect 34107 12353 34115 12373
rect 34080 12345 34115 12353
rect 33848 12149 33854 12179
rect 33875 12149 33879 12179
rect 33848 12141 33879 12149
rect 34006 12123 34046 12124
rect 33636 12121 34048 12123
rect 33636 12095 34016 12121
rect 34042 12095 34048 12121
rect 33636 12087 34048 12095
rect 33636 12059 33668 12087
rect 34081 12067 34115 12345
rect 34197 12158 34267 12469
rect 36122 12459 36194 12460
rect 36121 12456 36210 12459
rect 34893 12454 36210 12456
rect 34890 12451 36210 12454
rect 34890 12448 36173 12451
rect 34890 12413 36129 12448
rect 36154 12413 36173 12448
rect 36198 12413 36210 12451
rect 34890 12403 36210 12413
rect 36386 12452 36422 12605
rect 36386 12429 36392 12452
rect 36416 12429 36422 12452
rect 36386 12408 36422 12429
rect 34890 12401 36175 12403
rect 34890 12391 34987 12401
rect 34896 12382 34932 12391
rect 36386 12385 36392 12408
rect 36416 12385 36422 12408
rect 34306 12313 34509 12326
rect 34306 12280 34330 12313
rect 34366 12312 34509 12313
rect 34366 12309 34477 12312
rect 34366 12282 34403 12309
rect 34432 12285 34477 12309
rect 34506 12285 34509 12312
rect 34432 12282 34509 12285
rect 34366 12280 34509 12282
rect 34306 12267 34509 12280
rect 34306 12266 34407 12267
rect 33636 12039 33641 12059
rect 33662 12039 33668 12059
rect 33636 12032 33668 12039
rect 34059 12062 34115 12067
rect 34059 12042 34066 12062
rect 34086 12042 34115 12062
rect 34192 12152 34267 12158
rect 34192 12119 34200 12152
rect 34253 12119 34267 12152
rect 34192 12094 34267 12119
rect 34192 12061 34205 12094
rect 34258 12061 34267 12094
rect 34192 12052 34267 12061
rect 34684 12204 34716 12211
rect 34684 12184 34691 12204
rect 34712 12184 34716 12204
rect 34684 12119 34716 12184
rect 34896 12175 34927 12382
rect 35131 12374 35163 12375
rect 36386 12374 36422 12385
rect 35128 12369 35163 12374
rect 35128 12349 35135 12369
rect 35155 12349 35163 12369
rect 35128 12341 35163 12349
rect 34896 12145 34902 12175
rect 34923 12145 34927 12175
rect 34896 12137 34927 12145
rect 35054 12119 35094 12120
rect 34684 12117 35096 12119
rect 34684 12091 35064 12117
rect 35090 12091 35096 12117
rect 34684 12083 35096 12091
rect 34684 12055 34716 12083
rect 35129 12063 35163 12341
rect 34192 12047 34250 12052
rect 34059 12035 34115 12042
rect 34684 12035 34689 12055
rect 34710 12035 34716 12055
rect 34059 12034 34094 12035
rect 34684 12028 34716 12035
rect 35107 12058 35163 12063
rect 35107 12038 35114 12058
rect 35134 12038 35163 12058
rect 35107 12031 35163 12038
rect 35107 12030 35142 12031
rect 33350 11979 33461 11983
rect 35225 11979 36466 11980
rect 32672 11961 36466 11979
rect 32672 11941 33358 11961
rect 33377 11941 33435 11961
rect 33454 11957 36466 11961
rect 33454 11941 34406 11957
rect 32672 11937 34406 11941
rect 34425 11937 34483 11957
rect 34502 11937 36466 11957
rect 32672 11923 36466 11937
rect 32672 11300 32779 11923
rect 34398 11920 34509 11923
rect 33158 11874 33222 11878
rect 33154 11868 33222 11874
rect 33154 11835 33171 11868
rect 33211 11835 33222 11868
rect 33154 11823 33222 11835
rect 34205 11837 34270 11859
rect 33154 11821 33211 11823
rect 33158 11460 33209 11821
rect 34205 11798 34222 11837
rect 34267 11798 34270 11837
rect 33846 11753 33881 11755
rect 33846 11744 33950 11753
rect 33846 11743 33897 11744
rect 33846 11723 33849 11743
rect 33874 11724 33897 11743
rect 33929 11724 33950 11744
rect 33874 11723 33950 11724
rect 33846 11716 33950 11723
rect 33846 11704 33881 11716
rect 33258 11638 33461 11651
rect 33258 11605 33282 11638
rect 33318 11637 33461 11638
rect 33318 11634 33429 11637
rect 33318 11607 33355 11634
rect 33384 11610 33429 11634
rect 33458 11610 33461 11637
rect 33384 11607 33461 11610
rect 33318 11605 33461 11607
rect 33258 11592 33461 11605
rect 33258 11591 33359 11592
rect 33636 11529 33668 11536
rect 33636 11509 33643 11529
rect 33664 11509 33668 11529
rect 33147 11451 33212 11460
rect 33147 11414 33157 11451
rect 33197 11417 33212 11451
rect 33636 11444 33668 11509
rect 33848 11500 33879 11704
rect 34083 11699 34115 11700
rect 34080 11694 34115 11699
rect 34080 11674 34087 11694
rect 34107 11674 34115 11694
rect 34080 11666 34115 11674
rect 33848 11470 33854 11500
rect 33875 11470 33879 11500
rect 33848 11462 33879 11470
rect 34006 11444 34046 11445
rect 33636 11442 34048 11444
rect 33197 11414 33214 11417
rect 33147 11395 33214 11414
rect 33147 11374 33161 11395
rect 33197 11374 33214 11395
rect 33147 11367 33214 11374
rect 33636 11416 34016 11442
rect 34042 11416 34048 11442
rect 33636 11408 34048 11416
rect 33636 11380 33668 11408
rect 34081 11388 34115 11666
rect 34205 11498 34270 11798
rect 36384 11792 36489 11801
rect 36384 11787 36438 11792
rect 36384 11766 36397 11787
rect 36417 11771 36438 11787
rect 36458 11771 36489 11792
rect 36417 11766 36489 11771
rect 36384 11735 36489 11766
rect 36387 11718 36422 11735
rect 36386 11700 36422 11718
rect 35796 11635 35999 11648
rect 35796 11602 35820 11635
rect 35856 11634 35999 11635
rect 35856 11631 35967 11634
rect 35856 11604 35893 11631
rect 35922 11607 35967 11631
rect 35996 11607 35999 11634
rect 35922 11604 35999 11607
rect 35856 11602 35999 11604
rect 35796 11589 35999 11602
rect 35796 11588 35897 11589
rect 36174 11526 36206 11533
rect 36174 11506 36181 11526
rect 36202 11506 36206 11526
rect 33636 11360 33641 11380
rect 33662 11360 33668 11380
rect 33636 11353 33668 11360
rect 34059 11383 34115 11388
rect 34059 11363 34066 11383
rect 34086 11363 34115 11383
rect 34059 11356 34115 11363
rect 34195 11487 34275 11498
rect 34195 11461 34212 11487
rect 34252 11461 34275 11487
rect 34195 11434 34275 11461
rect 34195 11408 34216 11434
rect 34256 11408 34275 11434
rect 34195 11389 34275 11408
rect 34195 11363 34219 11389
rect 34259 11363 34275 11389
rect 34059 11355 34094 11356
rect 34195 11351 34275 11363
rect 36174 11441 36206 11506
rect 36386 11497 36417 11700
rect 36621 11696 36653 11697
rect 36618 11691 36653 11696
rect 36618 11671 36625 11691
rect 36645 11671 36653 11691
rect 36618 11663 36653 11671
rect 36386 11467 36392 11497
rect 36413 11467 36417 11497
rect 36386 11459 36417 11467
rect 36544 11441 36584 11442
rect 36174 11439 36586 11441
rect 36174 11413 36554 11439
rect 36580 11413 36586 11439
rect 36174 11405 36586 11413
rect 36174 11377 36206 11405
rect 36619 11385 36653 11663
rect 36174 11357 36179 11377
rect 36200 11357 36206 11377
rect 36174 11350 36206 11357
rect 36597 11380 36653 11385
rect 36597 11360 36604 11380
rect 36624 11360 36653 11380
rect 36597 11353 36653 11360
rect 36597 11352 36632 11353
rect 33350 11300 33461 11304
rect 35105 11300 35312 11301
rect 35888 11300 35999 11301
rect 32670 11282 36690 11300
rect 32670 11262 33358 11282
rect 33377 11262 33435 11282
rect 33454 11279 36690 11282
rect 33454 11262 35896 11279
rect 32670 11259 35896 11262
rect 35915 11259 35973 11279
rect 35992 11259 36690 11279
rect 32670 11244 36690 11259
rect 32672 11056 32779 11244
rect 35267 11242 36690 11244
rect 33140 11205 33261 11215
rect 33140 11203 33209 11205
rect 33140 11162 33153 11203
rect 33190 11164 33209 11203
rect 33246 11164 33261 11205
rect 33190 11162 33261 11164
rect 33140 11144 33261 11162
rect 32672 11052 32780 11056
rect 33146 11052 33223 11144
rect 34196 11140 34272 11156
rect 34196 11117 34211 11140
rect 30679 10886 30694 10909
rect 30618 10870 30694 10886
rect 31667 10882 31744 10974
rect 32110 10970 32218 10974
rect 31629 10864 31750 10882
rect 31629 10862 31700 10864
rect 31629 10821 31644 10862
rect 31681 10823 31700 10862
rect 31737 10823 31750 10864
rect 31681 10821 31750 10823
rect 31629 10811 31750 10821
rect 28154 10782 29623 10784
rect 32111 10782 32218 10970
rect 28154 10767 32220 10782
rect 28154 10747 28898 10767
rect 28917 10747 28975 10767
rect 28994 10764 32220 10767
rect 28994 10747 31436 10764
rect 28154 10744 31436 10747
rect 31455 10744 31513 10764
rect 31532 10744 32220 10764
rect 28154 10726 32220 10744
rect 28891 10725 29002 10726
rect 29578 10725 29785 10726
rect 31429 10722 31540 10726
rect 28258 10673 28293 10674
rect 28237 10666 28293 10673
rect 28237 10646 28266 10666
rect 28286 10646 28293 10666
rect 28237 10641 28293 10646
rect 28684 10669 28716 10676
rect 28684 10649 28690 10669
rect 28711 10649 28716 10669
rect 28237 10363 28271 10641
rect 28684 10621 28716 10649
rect 28304 10613 28716 10621
rect 28304 10587 28310 10613
rect 28336 10587 28716 10613
rect 28304 10585 28716 10587
rect 28306 10584 28346 10585
rect 28473 10559 28504 10567
rect 28473 10529 28477 10559
rect 28498 10529 28504 10559
rect 28237 10355 28272 10363
rect 28237 10335 28245 10355
rect 28265 10335 28272 10355
rect 28237 10330 28272 10335
rect 28473 10333 28504 10529
rect 28684 10520 28716 10585
rect 30615 10663 30695 10675
rect 30796 10670 30831 10671
rect 30615 10637 30631 10663
rect 30671 10637 30695 10663
rect 30615 10618 30695 10637
rect 30615 10592 30634 10618
rect 30674 10592 30695 10618
rect 30615 10565 30695 10592
rect 30615 10539 30638 10565
rect 30678 10539 30695 10565
rect 30615 10528 30695 10539
rect 30775 10663 30831 10670
rect 30775 10643 30804 10663
rect 30824 10643 30831 10663
rect 30775 10638 30831 10643
rect 31222 10666 31254 10673
rect 31222 10646 31228 10666
rect 31249 10646 31254 10666
rect 28684 10500 28688 10520
rect 28709 10500 28716 10520
rect 28684 10493 28716 10500
rect 28993 10437 29094 10438
rect 28891 10424 29094 10437
rect 28891 10422 29034 10424
rect 28891 10419 28968 10422
rect 28891 10392 28894 10419
rect 28923 10395 28968 10419
rect 28997 10395 29034 10422
rect 28923 10392 29034 10395
rect 28891 10391 29034 10392
rect 29070 10391 29094 10424
rect 28891 10378 29094 10391
rect 28237 10329 28269 10330
rect 28473 10244 28507 10333
rect 28094 10240 28507 10244
rect 27080 7915 27097 7969
rect 27160 7915 27185 7969
rect 27080 7894 27185 7915
rect 27547 10195 28507 10240
rect 30620 10228 30685 10528
rect 30775 10360 30809 10638
rect 31222 10618 31254 10646
rect 30842 10610 31254 10618
rect 30842 10584 30848 10610
rect 30874 10584 31254 10610
rect 31676 10652 31743 10659
rect 31676 10631 31693 10652
rect 31729 10631 31743 10652
rect 31676 10612 31743 10631
rect 31676 10609 31693 10612
rect 30842 10582 31254 10584
rect 30844 10581 30884 10582
rect 31011 10556 31042 10564
rect 31011 10526 31015 10556
rect 31036 10526 31042 10556
rect 30775 10352 30810 10360
rect 30775 10332 30783 10352
rect 30803 10332 30810 10352
rect 30775 10327 30810 10332
rect 30775 10326 30807 10327
rect 31011 10322 31042 10526
rect 31222 10517 31254 10582
rect 31678 10575 31693 10609
rect 31733 10575 31743 10612
rect 31678 10566 31743 10575
rect 31222 10497 31226 10517
rect 31247 10497 31254 10517
rect 31222 10490 31254 10497
rect 31531 10434 31632 10435
rect 31429 10421 31632 10434
rect 31429 10419 31572 10421
rect 31429 10416 31506 10419
rect 31429 10389 31432 10416
rect 31461 10392 31506 10416
rect 31535 10392 31572 10419
rect 31461 10389 31572 10392
rect 31429 10388 31572 10389
rect 31608 10388 31632 10421
rect 31429 10375 31632 10388
rect 31009 10310 31044 10322
rect 30940 10303 31044 10310
rect 30940 10302 31016 10303
rect 30940 10282 30961 10302
rect 30993 10283 31016 10302
rect 31041 10283 31044 10303
rect 30993 10282 31044 10283
rect 30940 10273 31044 10282
rect 31009 10271 31044 10273
rect 27547 10191 28144 10195
rect 27547 7885 27599 10191
rect 30620 10189 30623 10228
rect 30668 10189 30685 10228
rect 31681 10205 31732 10566
rect 31679 10203 31736 10205
rect 30620 10167 30685 10189
rect 31668 10191 31736 10203
rect 31668 10158 31679 10191
rect 31719 10158 31736 10191
rect 31668 10152 31736 10158
rect 31668 10148 31732 10152
rect 30381 10103 30492 10106
rect 32111 10103 32218 10726
rect 28506 10089 32218 10103
rect 28506 10069 30388 10089
rect 30407 10069 30465 10089
rect 30484 10085 32218 10089
rect 30484 10069 31436 10085
rect 28506 10065 31436 10069
rect 31455 10065 31513 10085
rect 31532 10065 32218 10085
rect 28506 10047 32218 10065
rect 28506 10046 29665 10047
rect 31429 10043 31540 10047
rect 29748 9995 29783 9996
rect 29727 9988 29783 9995
rect 29727 9968 29756 9988
rect 29776 9968 29783 9988
rect 29727 9963 29783 9968
rect 30174 9991 30206 9998
rect 30796 9991 30831 9992
rect 30174 9971 30180 9991
rect 30201 9971 30206 9991
rect 30775 9984 30831 9991
rect 30640 9974 30698 9979
rect 29727 9685 29761 9963
rect 30174 9943 30206 9971
rect 29794 9935 30206 9943
rect 29794 9909 29800 9935
rect 29826 9909 30206 9935
rect 29794 9907 30206 9909
rect 29796 9906 29836 9907
rect 29963 9881 29994 9889
rect 29963 9851 29967 9881
rect 29988 9851 29994 9881
rect 29727 9677 29762 9685
rect 29727 9657 29735 9677
rect 29755 9657 29762 9677
rect 29727 9652 29762 9657
rect 28468 9641 28504 9652
rect 29727 9651 29759 9652
rect 29963 9644 29994 9851
rect 30174 9842 30206 9907
rect 30174 9822 30178 9842
rect 30199 9822 30206 9842
rect 30174 9815 30206 9822
rect 30623 9965 30698 9974
rect 30623 9932 30632 9965
rect 30685 9932 30698 9965
rect 30623 9907 30698 9932
rect 30623 9874 30637 9907
rect 30690 9874 30698 9907
rect 30623 9868 30698 9874
rect 30775 9964 30804 9984
rect 30824 9964 30831 9984
rect 30775 9959 30831 9964
rect 31222 9987 31254 9994
rect 31222 9967 31228 9987
rect 31249 9967 31254 9987
rect 30483 9759 30584 9760
rect 30381 9746 30584 9759
rect 30381 9744 30524 9746
rect 30381 9741 30458 9744
rect 30381 9714 30384 9741
rect 30413 9717 30458 9741
rect 30487 9717 30524 9744
rect 30413 9714 30524 9717
rect 30381 9713 30524 9714
rect 30560 9713 30584 9746
rect 30381 9700 30584 9713
rect 28468 9618 28474 9641
rect 28498 9618 28504 9641
rect 29958 9635 29994 9644
rect 29903 9625 30000 9635
rect 28715 9623 30000 9625
rect 28468 9597 28504 9618
rect 28468 9574 28474 9597
rect 28498 9574 28504 9597
rect 28468 9421 28504 9574
rect 28680 9613 30000 9623
rect 28680 9575 28692 9613
rect 28717 9578 28736 9613
rect 28761 9578 30000 9613
rect 28717 9575 30000 9578
rect 28680 9572 30000 9575
rect 28680 9570 29997 9572
rect 28680 9567 28769 9570
rect 28696 9566 28768 9567
rect 30623 9557 30693 9868
rect 30775 9681 30809 9959
rect 31222 9939 31254 9967
rect 30842 9931 31254 9939
rect 30842 9905 30848 9931
rect 30874 9905 31254 9931
rect 30842 9903 31254 9905
rect 30844 9902 30884 9903
rect 31011 9877 31042 9885
rect 31011 9847 31015 9877
rect 31036 9847 31042 9877
rect 30775 9673 30810 9681
rect 30775 9653 30783 9673
rect 30803 9653 30810 9673
rect 30775 9648 30810 9653
rect 31011 9648 31042 9847
rect 31222 9838 31254 9903
rect 31222 9818 31226 9838
rect 31247 9818 31254 9838
rect 31222 9811 31254 9818
rect 31667 9964 31739 9982
rect 31667 9922 31680 9964
rect 31729 9922 31739 9964
rect 31667 9901 31739 9922
rect 31667 9859 31681 9901
rect 31730 9859 31739 9901
rect 31531 9755 31632 9756
rect 31429 9742 31632 9755
rect 31429 9740 31572 9742
rect 31429 9737 31506 9740
rect 31429 9710 31432 9737
rect 31461 9713 31506 9737
rect 31535 9713 31572 9740
rect 31461 9710 31572 9713
rect 31429 9709 31572 9710
rect 31608 9709 31632 9742
rect 31429 9696 31632 9709
rect 30775 9647 30807 9648
rect 31009 9645 31042 9648
rect 30975 9626 31043 9645
rect 30945 9614 31044 9626
rect 31667 9618 31739 9859
rect 32111 9618 32218 10047
rect 32673 10459 32780 11052
rect 33148 11001 33223 11052
rect 34189 11103 34211 11117
rect 34255 11103 34272 11140
rect 34189 11083 34272 11103
rect 34189 11017 34206 11083
rect 34260 11017 34272 11083
rect 33148 10958 33224 11001
rect 33152 10647 33224 10958
rect 34189 10993 34272 11017
rect 34189 10973 34265 10993
rect 34189 10954 34268 10973
rect 33848 10938 33920 10939
rect 33847 10930 33946 10938
rect 33847 10927 33899 10930
rect 33847 10892 33855 10927
rect 33880 10892 33899 10927
rect 33924 10892 33946 10930
rect 33847 10880 33946 10892
rect 33848 10861 33916 10880
rect 33849 10858 33882 10861
rect 34084 10858 34116 10859
rect 33259 10797 33462 10810
rect 33259 10764 33283 10797
rect 33319 10796 33462 10797
rect 33319 10793 33430 10796
rect 33319 10766 33356 10793
rect 33385 10769 33430 10793
rect 33459 10769 33462 10796
rect 33385 10766 33462 10769
rect 33319 10764 33462 10766
rect 33259 10751 33462 10764
rect 33259 10750 33360 10751
rect 33152 10605 33161 10647
rect 33210 10605 33224 10647
rect 33152 10584 33224 10605
rect 33152 10542 33162 10584
rect 33211 10542 33224 10584
rect 33152 10524 33224 10542
rect 33637 10688 33669 10695
rect 33637 10668 33644 10688
rect 33665 10668 33669 10688
rect 33637 10603 33669 10668
rect 33849 10659 33880 10858
rect 34081 10853 34116 10858
rect 34081 10833 34088 10853
rect 34108 10833 34116 10853
rect 34081 10825 34116 10833
rect 33849 10629 33855 10659
rect 33876 10629 33880 10659
rect 33849 10621 33880 10629
rect 34007 10603 34047 10604
rect 33637 10601 34049 10603
rect 33637 10575 34017 10601
rect 34043 10575 34049 10601
rect 33637 10567 34049 10575
rect 33637 10539 33669 10567
rect 34082 10547 34116 10825
rect 34198 10638 34268 10954
rect 36186 10939 36217 10940
rect 36186 10931 36231 10939
rect 35266 10908 35430 10915
rect 36186 10908 36196 10931
rect 34892 10893 36196 10908
rect 36221 10893 36231 10931
rect 34892 10875 36231 10893
rect 34897 10862 34933 10875
rect 35266 10872 35430 10875
rect 34307 10793 34510 10806
rect 34307 10760 34331 10793
rect 34367 10792 34510 10793
rect 34367 10789 34478 10792
rect 34367 10762 34404 10789
rect 34433 10765 34478 10789
rect 34507 10765 34510 10792
rect 34433 10762 34510 10765
rect 34367 10760 34510 10762
rect 34307 10747 34510 10760
rect 34307 10746 34408 10747
rect 33637 10519 33642 10539
rect 33663 10519 33669 10539
rect 33637 10512 33669 10519
rect 34060 10542 34116 10547
rect 34060 10522 34067 10542
rect 34087 10522 34116 10542
rect 34193 10632 34268 10638
rect 34193 10599 34201 10632
rect 34254 10599 34268 10632
rect 34193 10574 34268 10599
rect 34193 10541 34206 10574
rect 34259 10541 34268 10574
rect 34193 10532 34268 10541
rect 34685 10684 34717 10691
rect 34685 10664 34692 10684
rect 34713 10664 34717 10684
rect 34685 10599 34717 10664
rect 34897 10655 34928 10862
rect 35132 10854 35164 10855
rect 35129 10849 35164 10854
rect 35129 10829 35136 10849
rect 35156 10829 35164 10849
rect 35129 10821 35164 10829
rect 34897 10625 34903 10655
rect 34924 10625 34928 10655
rect 34897 10617 34928 10625
rect 35055 10599 35095 10600
rect 34685 10597 35097 10599
rect 34685 10571 35065 10597
rect 35091 10571 35097 10597
rect 34685 10563 35097 10571
rect 34685 10535 34717 10563
rect 35130 10543 35164 10821
rect 34193 10527 34251 10532
rect 34060 10515 34116 10522
rect 34685 10515 34690 10535
rect 34711 10515 34717 10535
rect 34060 10514 34095 10515
rect 34685 10508 34717 10515
rect 35108 10538 35164 10543
rect 35108 10518 35115 10538
rect 35135 10518 35164 10538
rect 35108 10511 35164 10518
rect 35108 10510 35143 10511
rect 33351 10459 33462 10463
rect 35134 10459 36434 10460
rect 32673 10441 36434 10459
rect 32673 10421 33359 10441
rect 33378 10421 33436 10441
rect 33455 10437 36434 10441
rect 33455 10421 34407 10437
rect 32673 10417 34407 10421
rect 34426 10417 34484 10437
rect 34503 10417 36434 10437
rect 32673 10403 36434 10417
rect 32673 9780 32780 10403
rect 34399 10400 34510 10403
rect 33159 10354 33223 10358
rect 33155 10348 33223 10354
rect 33155 10315 33172 10348
rect 33212 10315 33223 10348
rect 33155 10303 33223 10315
rect 34206 10317 34271 10339
rect 33155 10301 33212 10303
rect 33159 9940 33210 10301
rect 34206 10278 34223 10317
rect 34268 10278 34271 10317
rect 33847 10233 33882 10235
rect 33847 10224 33951 10233
rect 33847 10223 33898 10224
rect 33847 10203 33850 10223
rect 33875 10204 33898 10223
rect 33930 10204 33951 10224
rect 33875 10203 33951 10204
rect 33847 10196 33951 10203
rect 33847 10184 33882 10196
rect 33259 10118 33462 10131
rect 33259 10085 33283 10118
rect 33319 10117 33462 10118
rect 33319 10114 33430 10117
rect 33319 10087 33356 10114
rect 33385 10090 33430 10114
rect 33459 10090 33462 10117
rect 33385 10087 33462 10090
rect 33319 10085 33462 10087
rect 33259 10072 33462 10085
rect 33259 10071 33360 10072
rect 33637 10009 33669 10016
rect 33637 9989 33644 10009
rect 33665 9989 33669 10009
rect 33148 9931 33213 9940
rect 33148 9894 33158 9931
rect 33198 9897 33213 9931
rect 33637 9924 33669 9989
rect 33849 9980 33880 10184
rect 34084 10179 34116 10180
rect 34081 10174 34116 10179
rect 34081 10154 34088 10174
rect 34108 10154 34116 10174
rect 34081 10146 34116 10154
rect 33849 9950 33855 9980
rect 33876 9950 33880 9980
rect 33849 9942 33880 9950
rect 34007 9924 34047 9925
rect 33637 9922 34049 9924
rect 33198 9894 33215 9897
rect 33148 9875 33215 9894
rect 33148 9854 33162 9875
rect 33198 9854 33215 9875
rect 33148 9847 33215 9854
rect 33637 9896 34017 9922
rect 34043 9896 34049 9922
rect 33637 9888 34049 9896
rect 33637 9860 33669 9888
rect 34082 9868 34116 10146
rect 34206 9978 34271 10278
rect 36343 10239 36380 10260
rect 36343 10202 36354 10239
rect 36371 10215 36380 10239
rect 36371 10202 36381 10215
rect 36343 10192 36381 10202
rect 36344 10188 36381 10192
rect 36344 10182 36377 10188
rect 35754 10113 35957 10126
rect 35754 10080 35778 10113
rect 35814 10112 35957 10113
rect 35814 10109 35925 10112
rect 35814 10082 35851 10109
rect 35880 10085 35925 10109
rect 35954 10085 35957 10112
rect 35880 10082 35957 10085
rect 35814 10080 35957 10082
rect 35754 10067 35957 10080
rect 35754 10066 35855 10067
rect 36132 10004 36164 10011
rect 36132 9984 36139 10004
rect 36160 9984 36164 10004
rect 33637 9840 33642 9860
rect 33663 9840 33669 9860
rect 33637 9833 33669 9840
rect 34060 9863 34116 9868
rect 34060 9843 34067 9863
rect 34087 9843 34116 9863
rect 34060 9836 34116 9843
rect 34196 9967 34276 9978
rect 34196 9941 34213 9967
rect 34253 9941 34276 9967
rect 34196 9914 34276 9941
rect 34196 9888 34217 9914
rect 34257 9888 34276 9914
rect 36132 9919 36164 9984
rect 36344 9975 36375 10182
rect 36579 10174 36611 10175
rect 36576 10169 36611 10174
rect 36576 10149 36583 10169
rect 36603 10149 36611 10169
rect 36576 10141 36611 10149
rect 36344 9945 36350 9975
rect 36371 9945 36375 9975
rect 36344 9937 36375 9945
rect 36502 9919 36542 9920
rect 36132 9917 36544 9919
rect 34196 9869 34276 9888
rect 34196 9843 34220 9869
rect 34260 9843 34276 9869
rect 35309 9907 35746 9913
rect 35309 9884 35327 9907
rect 35353 9900 35746 9907
rect 35353 9884 35707 9900
rect 35309 9877 35707 9884
rect 35733 9877 35746 9900
rect 35309 9864 35746 9877
rect 36132 9891 36512 9917
rect 36538 9891 36544 9917
rect 36132 9883 36544 9891
rect 34060 9835 34095 9836
rect 34196 9831 34276 9843
rect 36132 9855 36164 9883
rect 36577 9863 36611 10141
rect 36132 9835 36137 9855
rect 36158 9835 36164 9855
rect 36132 9828 36164 9835
rect 36555 9858 36611 9863
rect 36555 9838 36562 9858
rect 36582 9838 36611 9858
rect 36555 9831 36611 9838
rect 36555 9830 36590 9831
rect 33351 9780 33462 9784
rect 35093 9780 36643 9783
rect 32671 9762 36643 9780
rect 32671 9742 33359 9762
rect 33378 9742 33436 9762
rect 33455 9757 36643 9762
rect 33455 9742 35854 9757
rect 32671 9737 35854 9742
rect 35873 9737 35931 9757
rect 35950 9737 36643 9757
rect 32671 9727 36643 9737
rect 32671 9724 33296 9727
rect 33483 9724 36643 9727
rect 30945 9576 30967 9614
rect 30992 9579 31011 9614
rect 31036 9579 31044 9614
rect 30992 9576 31044 9579
rect 30945 9568 31044 9576
rect 30971 9567 31043 9568
rect 30622 9541 30693 9557
rect 30622 9525 30642 9541
rect 30623 9495 30642 9525
rect 30625 9475 30642 9495
rect 30672 9495 30693 9541
rect 31665 9537 31743 9618
rect 32110 9563 32218 9618
rect 30672 9475 30692 9495
rect 30625 9456 30692 9475
rect 31665 9435 31744 9537
rect 28459 9412 28545 9421
rect 28459 9394 28478 9412
rect 28530 9394 28545 9412
rect 28459 9390 28545 9394
rect 31629 9417 31750 9435
rect 31629 9415 31700 9417
rect 31629 9374 31644 9415
rect 31681 9376 31700 9415
rect 31737 9376 31750 9417
rect 31681 9374 31750 9376
rect 31629 9364 31750 9374
rect 28934 9336 29045 9339
rect 28154 9335 29798 9336
rect 32111 9335 32218 9563
rect 32673 9496 32780 9724
rect 35093 9723 36643 9724
rect 35846 9720 35957 9723
rect 33141 9685 33262 9695
rect 33141 9683 33210 9685
rect 33141 9642 33154 9683
rect 33191 9644 33210 9683
rect 33247 9644 33262 9685
rect 33191 9642 33262 9644
rect 33141 9624 33262 9642
rect 33147 9522 33226 9624
rect 34199 9584 34266 9603
rect 34199 9564 34219 9584
rect 32673 9441 32781 9496
rect 33148 9441 33226 9522
rect 34198 9518 34219 9564
rect 34249 9564 34266 9584
rect 34249 9534 34268 9564
rect 34249 9518 34269 9534
rect 34198 9502 34269 9518
rect 33848 9491 33920 9492
rect 33847 9483 33946 9491
rect 33847 9480 33899 9483
rect 33847 9445 33855 9480
rect 33880 9445 33899 9480
rect 33924 9445 33946 9483
rect 28154 9332 31408 9335
rect 31595 9332 32220 9335
rect 28154 9322 32220 9332
rect 28154 9302 28941 9322
rect 28960 9302 29018 9322
rect 29037 9317 32220 9322
rect 29037 9302 31436 9317
rect 28154 9297 31436 9302
rect 31455 9297 31513 9317
rect 31532 9297 32220 9317
rect 28154 9279 32220 9297
rect 28154 9276 29798 9279
rect 31429 9275 31540 9279
rect 28301 9228 28336 9229
rect 28280 9221 28336 9228
rect 28280 9201 28309 9221
rect 28329 9201 28336 9221
rect 28280 9196 28336 9201
rect 28727 9224 28759 9231
rect 28727 9204 28733 9224
rect 28754 9204 28759 9224
rect 28280 8918 28314 9196
rect 28727 9176 28759 9204
rect 28347 9168 28759 9176
rect 28347 9142 28353 9168
rect 28379 9142 28759 9168
rect 28347 9140 28759 9142
rect 28349 9139 28389 9140
rect 28516 9114 28547 9122
rect 28516 9084 28520 9114
rect 28541 9084 28547 9114
rect 28280 8910 28315 8918
rect 28280 8890 28288 8910
rect 28308 8890 28315 8910
rect 28280 8885 28315 8890
rect 28280 8884 28312 8885
rect 28516 8883 28547 9084
rect 28727 9075 28759 9140
rect 28727 9055 28731 9075
rect 28752 9055 28759 9075
rect 28727 9048 28759 9055
rect 29321 9215 29414 9222
rect 29321 9174 29345 9215
rect 29399 9174 29414 9215
rect 29036 8992 29137 8993
rect 28934 8979 29137 8992
rect 28934 8977 29077 8979
rect 28934 8974 29011 8977
rect 28934 8947 28937 8974
rect 28966 8950 29011 8974
rect 29040 8950 29077 8977
rect 28966 8947 29077 8950
rect 28934 8946 29077 8947
rect 29113 8946 29137 8979
rect 28934 8933 29137 8946
rect 29321 8801 29414 9174
rect 30615 9216 30695 9228
rect 30796 9223 30831 9224
rect 30615 9190 30631 9216
rect 30671 9190 30695 9216
rect 30615 9171 30695 9190
rect 30615 9145 30634 9171
rect 30674 9145 30695 9171
rect 30615 9118 30695 9145
rect 30615 9092 30638 9118
rect 30678 9092 30695 9118
rect 30615 9081 30695 9092
rect 30775 9216 30831 9223
rect 30775 9196 30804 9216
rect 30824 9196 30831 9216
rect 30775 9191 30831 9196
rect 31222 9219 31254 9226
rect 31222 9199 31228 9219
rect 31249 9199 31254 9219
rect 29321 8757 29339 8801
rect 29399 8757 29414 8801
rect 29321 8742 29414 8757
rect 30620 8781 30685 9081
rect 30775 8913 30809 9191
rect 31222 9171 31254 9199
rect 30842 9163 31254 9171
rect 30842 9137 30848 9163
rect 30874 9137 31254 9163
rect 31676 9205 31743 9212
rect 31676 9184 31693 9205
rect 31729 9184 31743 9205
rect 31676 9165 31743 9184
rect 31676 9162 31693 9165
rect 30842 9135 31254 9137
rect 30844 9134 30884 9135
rect 31011 9109 31042 9117
rect 31011 9079 31015 9109
rect 31036 9079 31042 9109
rect 30775 8905 30810 8913
rect 30775 8885 30783 8905
rect 30803 8885 30810 8905
rect 30775 8880 30810 8885
rect 30775 8879 30807 8880
rect 31011 8875 31042 9079
rect 31222 9070 31254 9135
rect 31678 9128 31693 9162
rect 31733 9128 31743 9165
rect 31678 9119 31743 9128
rect 31222 9050 31226 9070
rect 31247 9050 31254 9070
rect 31222 9043 31254 9050
rect 31531 8987 31632 8988
rect 31429 8974 31632 8987
rect 31429 8972 31572 8974
rect 31429 8969 31506 8972
rect 31429 8942 31432 8969
rect 31461 8945 31506 8969
rect 31535 8945 31572 8972
rect 31461 8942 31572 8945
rect 31429 8941 31572 8942
rect 31608 8941 31632 8974
rect 31429 8928 31632 8941
rect 31009 8863 31044 8875
rect 30940 8856 31044 8863
rect 30940 8855 31016 8856
rect 30940 8835 30961 8855
rect 30993 8836 31016 8855
rect 31041 8836 31044 8856
rect 30993 8835 31044 8836
rect 30940 8826 31044 8835
rect 31009 8824 31044 8826
rect 30620 8742 30623 8781
rect 30668 8742 30685 8781
rect 31681 8758 31732 9119
rect 31679 8756 31736 8758
rect 30620 8720 30685 8742
rect 31668 8744 31736 8756
rect 31668 8711 31679 8744
rect 31719 8711 31736 8744
rect 31668 8705 31736 8711
rect 31668 8701 31732 8705
rect 30381 8656 30492 8659
rect 32111 8656 32218 9279
rect 28187 8642 32218 8656
rect 28187 8622 30388 8642
rect 30407 8622 30465 8642
rect 30484 8638 32218 8642
rect 30484 8622 31436 8638
rect 28187 8618 31436 8622
rect 31455 8618 31513 8638
rect 31532 8618 32218 8638
rect 28187 8600 32218 8618
rect 28187 8599 29757 8600
rect 31429 8596 31540 8600
rect 29748 8548 29783 8549
rect 29727 8541 29783 8548
rect 29727 8521 29756 8541
rect 29776 8521 29783 8541
rect 29727 8516 29783 8521
rect 30174 8544 30206 8551
rect 30796 8544 30831 8545
rect 30174 8524 30180 8544
rect 30201 8524 30206 8544
rect 30775 8537 30831 8544
rect 30640 8527 30698 8532
rect 29327 8461 29409 8490
rect 29327 8420 29352 8461
rect 29388 8420 29409 8461
rect 29514 8481 29578 8500
rect 29514 8442 29531 8481
rect 29565 8442 29578 8481
rect 29514 8423 29578 8442
rect 29327 8105 29409 8420
rect 29319 8060 29409 8105
rect 29516 8078 29578 8423
rect 29727 8238 29761 8516
rect 30174 8496 30206 8524
rect 29794 8488 30206 8496
rect 29794 8462 29800 8488
rect 29826 8462 30206 8488
rect 29794 8460 30206 8462
rect 29796 8459 29836 8460
rect 29963 8434 29994 8442
rect 29963 8404 29967 8434
rect 29988 8404 29994 8434
rect 29727 8230 29762 8238
rect 29727 8210 29735 8230
rect 29755 8210 29762 8230
rect 29727 8205 29762 8210
rect 29727 8204 29759 8205
rect 29963 8197 29994 8404
rect 30174 8395 30206 8460
rect 30174 8375 30178 8395
rect 30199 8375 30206 8395
rect 30174 8368 30206 8375
rect 30623 8518 30698 8527
rect 30623 8485 30632 8518
rect 30685 8485 30698 8518
rect 30623 8460 30698 8485
rect 30623 8427 30637 8460
rect 30690 8427 30698 8460
rect 30623 8421 30698 8427
rect 30775 8517 30804 8537
rect 30824 8517 30831 8537
rect 30775 8512 30831 8517
rect 31222 8540 31254 8547
rect 31222 8520 31228 8540
rect 31249 8520 31254 8540
rect 30483 8312 30584 8313
rect 30381 8299 30584 8312
rect 30381 8297 30524 8299
rect 30381 8294 30458 8297
rect 30381 8267 30384 8294
rect 30413 8270 30458 8294
rect 30487 8270 30524 8297
rect 30413 8267 30524 8270
rect 30381 8266 30524 8267
rect 30560 8266 30584 8299
rect 30381 8253 30584 8266
rect 29958 8179 29994 8197
rect 29925 8178 29994 8179
rect 29905 8166 29994 8178
rect 29905 8128 29917 8166
rect 29942 8131 29961 8166
rect 29986 8131 29994 8166
rect 30623 8155 30693 8421
rect 30775 8234 30809 8512
rect 31222 8492 31254 8520
rect 30842 8484 31254 8492
rect 30842 8458 30848 8484
rect 30874 8458 31254 8484
rect 30842 8456 31254 8458
rect 30844 8455 30884 8456
rect 31011 8430 31042 8438
rect 31011 8400 31015 8430
rect 31036 8400 31042 8430
rect 30775 8226 30810 8234
rect 30775 8206 30783 8226
rect 30803 8206 30810 8226
rect 30775 8201 30810 8206
rect 31011 8201 31042 8400
rect 31222 8391 31254 8456
rect 31222 8371 31226 8391
rect 31247 8371 31254 8391
rect 31222 8364 31254 8371
rect 31667 8517 31739 8535
rect 31667 8475 31680 8517
rect 31729 8475 31739 8517
rect 31667 8454 31739 8475
rect 31667 8412 31681 8454
rect 31730 8412 31739 8454
rect 31531 8308 31632 8309
rect 31429 8295 31632 8308
rect 31429 8293 31572 8295
rect 31429 8290 31506 8293
rect 31429 8263 31432 8290
rect 31461 8266 31506 8290
rect 31535 8266 31572 8293
rect 31461 8263 31572 8266
rect 31429 8262 31572 8263
rect 31608 8262 31632 8295
rect 31429 8249 31632 8262
rect 30775 8200 30807 8201
rect 31009 8198 31042 8201
rect 30975 8179 31043 8198
rect 29942 8128 29994 8131
rect 29905 8120 29994 8128
rect 30614 8126 30693 8155
rect 30945 8167 31044 8179
rect 30945 8129 30967 8167
rect 30992 8132 31011 8167
rect 31036 8132 31044 8167
rect 30992 8129 31044 8132
rect 29921 8119 29993 8120
rect 29515 8069 29589 8078
rect 29319 8027 29403 8060
rect 29319 7999 29334 8027
rect 29378 7999 29403 8027
rect 29319 7970 29403 7999
rect 29515 8021 29529 8069
rect 29566 8021 29589 8069
rect 29515 7993 29589 8021
rect 29319 7942 29331 7970
rect 29375 7942 29403 7970
rect 29319 7931 29403 7942
rect 30614 7943 30691 8126
rect 30945 8121 31044 8129
rect 30971 8120 31043 8121
rect 31667 8118 31739 8412
rect 32111 8140 32218 8600
rect 32673 9012 32780 9441
rect 33152 9200 33224 9441
rect 33847 9433 33946 9445
rect 33848 9414 33916 9433
rect 33849 9411 33882 9414
rect 34084 9411 34116 9412
rect 33259 9350 33462 9363
rect 33259 9317 33283 9350
rect 33319 9349 33462 9350
rect 33319 9346 33430 9349
rect 33319 9319 33356 9346
rect 33385 9322 33430 9346
rect 33459 9322 33462 9349
rect 33385 9319 33462 9322
rect 33319 9317 33462 9319
rect 33259 9304 33462 9317
rect 33259 9303 33360 9304
rect 33152 9158 33161 9200
rect 33210 9158 33224 9200
rect 33152 9137 33224 9158
rect 33152 9095 33162 9137
rect 33211 9095 33224 9137
rect 33152 9077 33224 9095
rect 33637 9241 33669 9248
rect 33637 9221 33644 9241
rect 33665 9221 33669 9241
rect 33637 9156 33669 9221
rect 33849 9212 33880 9411
rect 34081 9406 34116 9411
rect 34081 9386 34088 9406
rect 34108 9386 34116 9406
rect 34081 9378 34116 9386
rect 33849 9182 33855 9212
rect 33876 9182 33880 9212
rect 33849 9174 33880 9182
rect 34007 9156 34047 9157
rect 33637 9154 34049 9156
rect 33637 9128 34017 9154
rect 34043 9128 34049 9154
rect 33637 9120 34049 9128
rect 33637 9092 33669 9120
rect 34082 9100 34116 9378
rect 34198 9191 34268 9502
rect 34895 9493 36237 9498
rect 34895 9491 36194 9493
rect 34892 9465 36194 9491
rect 36222 9465 36237 9493
rect 34892 9457 36237 9465
rect 34892 9432 34931 9457
rect 34892 9415 34933 9432
rect 34892 9408 34931 9415
rect 34307 9346 34510 9359
rect 34307 9313 34331 9346
rect 34367 9345 34510 9346
rect 34367 9342 34478 9345
rect 34367 9315 34404 9342
rect 34433 9318 34478 9342
rect 34507 9318 34510 9345
rect 34433 9315 34510 9318
rect 34367 9313 34510 9315
rect 34307 9300 34510 9313
rect 34307 9299 34408 9300
rect 33637 9072 33642 9092
rect 33663 9072 33669 9092
rect 33637 9065 33669 9072
rect 34060 9095 34116 9100
rect 34060 9075 34067 9095
rect 34087 9075 34116 9095
rect 34193 9185 34268 9191
rect 34193 9152 34201 9185
rect 34254 9152 34268 9185
rect 34193 9127 34268 9152
rect 34193 9094 34206 9127
rect 34259 9094 34268 9127
rect 34193 9085 34268 9094
rect 34685 9237 34717 9244
rect 34685 9217 34692 9237
rect 34713 9217 34717 9237
rect 34685 9152 34717 9217
rect 34897 9208 34928 9408
rect 35132 9407 35164 9408
rect 35129 9402 35164 9407
rect 35129 9382 35136 9402
rect 35156 9382 35164 9402
rect 35129 9374 35164 9382
rect 34897 9178 34903 9208
rect 34924 9178 34928 9208
rect 34897 9170 34928 9178
rect 35055 9152 35095 9153
rect 34685 9150 35097 9152
rect 34685 9124 35065 9150
rect 35091 9124 35097 9150
rect 34685 9116 35097 9124
rect 34685 9088 34717 9116
rect 35130 9096 35164 9374
rect 34193 9080 34251 9085
rect 34060 9068 34116 9075
rect 34685 9068 34690 9088
rect 34711 9068 34717 9088
rect 34060 9067 34095 9068
rect 34685 9061 34717 9068
rect 35108 9091 35164 9096
rect 35108 9071 35115 9091
rect 35135 9071 35164 9091
rect 35108 9064 35164 9071
rect 35108 9063 35143 9064
rect 33351 9012 33462 9016
rect 35226 9012 35665 9013
rect 32673 8994 35665 9012
rect 32673 8974 33359 8994
rect 33378 8974 33436 8994
rect 33455 8990 35665 8994
rect 33455 8974 34407 8990
rect 32673 8970 34407 8974
rect 34426 8970 34484 8990
rect 34503 8970 35665 8990
rect 32673 8956 35665 8970
rect 32673 8333 32780 8956
rect 34399 8953 34510 8956
rect 33159 8907 33223 8911
rect 33155 8901 33223 8907
rect 33155 8868 33172 8901
rect 33212 8868 33223 8901
rect 33155 8856 33223 8868
rect 34206 8870 34271 8892
rect 33155 8854 33212 8856
rect 33159 8493 33210 8854
rect 34206 8831 34223 8870
rect 34268 8831 34271 8870
rect 33847 8786 33882 8788
rect 33847 8777 33951 8786
rect 33847 8776 33898 8777
rect 33847 8756 33850 8776
rect 33875 8757 33898 8776
rect 33930 8757 33951 8777
rect 33875 8756 33951 8757
rect 33847 8749 33951 8756
rect 33847 8737 33882 8749
rect 33259 8671 33462 8684
rect 33259 8638 33283 8671
rect 33319 8670 33462 8671
rect 33319 8667 33430 8670
rect 33319 8640 33356 8667
rect 33385 8643 33430 8667
rect 33459 8643 33462 8670
rect 33385 8640 33462 8643
rect 33319 8638 33462 8640
rect 33259 8625 33462 8638
rect 33259 8624 33360 8625
rect 33637 8562 33669 8569
rect 33637 8542 33644 8562
rect 33665 8542 33669 8562
rect 33148 8484 33213 8493
rect 33148 8447 33158 8484
rect 33198 8450 33213 8484
rect 33637 8477 33669 8542
rect 33849 8533 33880 8737
rect 34084 8732 34116 8733
rect 34081 8727 34116 8732
rect 34081 8707 34088 8727
rect 34108 8707 34116 8727
rect 34081 8699 34116 8707
rect 33849 8503 33855 8533
rect 33876 8503 33880 8533
rect 33849 8495 33880 8503
rect 34007 8477 34047 8478
rect 33637 8475 34049 8477
rect 33198 8447 33215 8450
rect 33148 8428 33215 8447
rect 33148 8407 33162 8428
rect 33198 8407 33215 8428
rect 33148 8400 33215 8407
rect 33637 8449 34017 8475
rect 34043 8449 34049 8475
rect 33637 8441 34049 8449
rect 33637 8413 33669 8441
rect 34082 8421 34116 8699
rect 34206 8531 34271 8831
rect 33637 8393 33642 8413
rect 33663 8393 33669 8413
rect 33637 8386 33669 8393
rect 34060 8416 34116 8421
rect 34060 8396 34067 8416
rect 34087 8396 34116 8416
rect 34060 8389 34116 8396
rect 34196 8520 34276 8531
rect 34196 8494 34213 8520
rect 34253 8494 34276 8520
rect 34196 8467 34276 8494
rect 36748 8470 36797 13651
rect 37796 13063 37883 14218
rect 42386 13843 42451 13981
rect 42336 13825 42457 13843
rect 42336 13823 42407 13825
rect 42336 13782 42351 13823
rect 42388 13784 42407 13823
rect 42444 13784 42457 13825
rect 42388 13782 42457 13784
rect 42336 13772 42457 13782
rect 40271 13743 40330 13745
rect 42818 13743 42925 13943
rect 40271 13725 42927 13743
rect 40271 13705 42143 13725
rect 42162 13705 42220 13725
rect 42239 13705 42927 13725
rect 40271 13687 42927 13705
rect 40285 13686 40492 13687
rect 42136 13683 42247 13687
rect 41322 13624 41402 13636
rect 41503 13631 41538 13632
rect 41322 13598 41338 13624
rect 41378 13598 41402 13624
rect 41322 13579 41402 13598
rect 41322 13553 41341 13579
rect 41381 13553 41402 13579
rect 41322 13526 41402 13553
rect 41322 13500 41345 13526
rect 41385 13500 41402 13526
rect 41322 13489 41402 13500
rect 41482 13624 41538 13631
rect 41482 13604 41511 13624
rect 41531 13604 41538 13624
rect 41482 13599 41538 13604
rect 41929 13627 41961 13634
rect 41929 13607 41935 13627
rect 41956 13607 41961 13627
rect 41327 13189 41392 13489
rect 41482 13321 41516 13599
rect 41929 13579 41961 13607
rect 41549 13571 41961 13579
rect 41549 13545 41555 13571
rect 41581 13545 41961 13571
rect 42383 13613 42450 13620
rect 42383 13592 42400 13613
rect 42436 13592 42450 13613
rect 42383 13573 42450 13592
rect 42383 13570 42400 13573
rect 41549 13543 41961 13545
rect 41551 13542 41591 13543
rect 41718 13517 41749 13525
rect 41718 13487 41722 13517
rect 41743 13487 41749 13517
rect 41482 13313 41517 13321
rect 41482 13293 41490 13313
rect 41510 13293 41517 13313
rect 41482 13288 41517 13293
rect 41482 13287 41514 13288
rect 41718 13283 41749 13487
rect 41929 13478 41961 13543
rect 42385 13536 42400 13570
rect 42440 13536 42450 13573
rect 42385 13527 42450 13536
rect 41929 13458 41933 13478
rect 41954 13458 41961 13478
rect 41929 13451 41961 13458
rect 42238 13395 42339 13396
rect 42136 13382 42339 13395
rect 42136 13380 42279 13382
rect 42136 13377 42213 13380
rect 42136 13350 42139 13377
rect 42168 13353 42213 13377
rect 42242 13353 42279 13380
rect 42168 13350 42279 13353
rect 42136 13349 42279 13350
rect 42315 13349 42339 13382
rect 42136 13336 42339 13349
rect 41716 13271 41751 13283
rect 41647 13264 41751 13271
rect 41647 13263 41723 13264
rect 41647 13243 41668 13263
rect 41700 13244 41723 13263
rect 41748 13244 41751 13264
rect 41700 13243 41751 13244
rect 41647 13234 41751 13243
rect 41716 13232 41751 13234
rect 41327 13150 41330 13189
rect 41375 13150 41392 13189
rect 42388 13166 42439 13527
rect 42386 13164 42443 13166
rect 41327 13128 41392 13150
rect 42375 13152 42443 13164
rect 42375 13119 42386 13152
rect 42426 13119 42443 13152
rect 42375 13113 42443 13119
rect 42375 13109 42439 13113
rect 41088 13064 41199 13067
rect 42818 13064 42925 13687
rect 36862 8662 37065 8675
rect 36862 8629 36886 8662
rect 36922 8661 37065 8662
rect 36922 8658 37033 8661
rect 36922 8631 36959 8658
rect 36988 8634 37033 8658
rect 37062 8634 37065 8661
rect 36988 8631 37065 8634
rect 36922 8629 37065 8631
rect 36862 8616 37065 8629
rect 36862 8615 36963 8616
rect 37240 8553 37272 8560
rect 37240 8533 37247 8553
rect 37268 8533 37272 8553
rect 34196 8441 34217 8467
rect 34257 8441 34276 8467
rect 34196 8422 34276 8441
rect 36747 8460 36858 8470
rect 36747 8459 36812 8460
rect 36747 8435 36755 8459
rect 36779 8436 36812 8459
rect 36836 8436 36858 8460
rect 36779 8435 36858 8436
rect 36747 8428 36858 8435
rect 37240 8468 37272 8533
rect 37452 8524 37483 8724
rect 37687 8723 37719 8724
rect 37684 8718 37719 8723
rect 37684 8698 37691 8718
rect 37711 8698 37719 8718
rect 37684 8690 37719 8698
rect 37452 8494 37458 8524
rect 37479 8494 37483 8524
rect 37452 8486 37483 8494
rect 37610 8468 37650 8469
rect 37240 8466 37652 8468
rect 37240 8440 37620 8466
rect 37646 8440 37652 8466
rect 37240 8432 37652 8440
rect 34196 8396 34220 8422
rect 34260 8396 34276 8422
rect 34060 8388 34095 8389
rect 34196 8384 34276 8396
rect 37240 8404 37272 8432
rect 37685 8412 37719 8690
rect 37240 8384 37245 8404
rect 37266 8384 37272 8404
rect 37240 8377 37272 8384
rect 37451 8404 37485 8411
rect 37451 8382 37458 8404
rect 37482 8382 37485 8404
rect 33351 8333 33462 8337
rect 35106 8333 35313 8334
rect 32671 8328 36746 8333
rect 32671 8315 37065 8328
rect 32671 8295 33359 8315
rect 33378 8295 33436 8315
rect 33455 8306 37065 8315
rect 33455 8295 36962 8306
rect 32671 8286 36962 8295
rect 36981 8286 37039 8306
rect 37058 8286 37065 8306
rect 32671 8277 37065 8286
rect 31667 8080 31743 8118
rect 32111 8080 32224 8140
rect 32673 8104 32780 8277
rect 35268 8275 37065 8277
rect 36954 8269 37065 8275
rect 33141 8238 33262 8248
rect 33141 8236 33210 8238
rect 33141 8195 33154 8236
rect 33191 8197 33210 8236
rect 33247 8197 33262 8238
rect 33191 8195 33262 8197
rect 33141 8177 33262 8195
rect 37289 8227 37341 8258
rect 37289 8193 37298 8227
rect 37327 8193 37341 8227
rect 31678 7979 31743 8080
rect 30614 7900 30631 7943
rect 27547 7851 27562 7885
rect 27591 7851 27599 7885
rect 30619 7895 30631 7900
rect 30677 7895 30691 7943
rect 30619 7873 30691 7895
rect 31676 7933 31743 7979
rect 32113 7941 32224 8080
rect 27547 7825 27599 7851
rect 31676 7841 31741 7933
rect 32108 7914 32224 7941
rect 32664 8077 32780 8104
rect 33147 8085 33212 8177
rect 37289 8167 37341 8193
rect 37451 8176 37485 8382
rect 37663 8407 37719 8412
rect 37663 8387 37670 8407
rect 37690 8387 37719 8407
rect 37663 8380 37719 8387
rect 37663 8379 37698 8380
rect 32664 7938 32775 8077
rect 33145 8039 33212 8085
rect 34197 8123 34269 8145
rect 34197 8075 34211 8123
rect 34257 8118 34269 8123
rect 37289 8133 37297 8167
rect 37326 8133 37341 8167
rect 34257 8075 34274 8118
rect 33145 7938 33210 8039
rect 27547 7791 27561 7825
rect 27590 7791 27599 7825
rect 27547 7760 27599 7791
rect 31626 7823 31747 7841
rect 31626 7821 31697 7823
rect 31626 7780 31641 7821
rect 31678 7782 31697 7821
rect 31734 7782 31747 7823
rect 31678 7780 31747 7782
rect 31626 7770 31747 7780
rect 27823 7743 27934 7749
rect 27823 7741 29620 7743
rect 32108 7741 32215 7914
rect 32664 7878 32777 7938
rect 33145 7900 33221 7938
rect 27823 7732 32217 7741
rect 27823 7712 27830 7732
rect 27849 7712 27907 7732
rect 27926 7723 32217 7732
rect 27926 7712 31433 7723
rect 27823 7703 31433 7712
rect 31452 7703 31510 7723
rect 31529 7703 32217 7723
rect 27823 7690 32217 7703
rect 28142 7685 32217 7690
rect 29575 7684 29782 7685
rect 31426 7681 31537 7685
rect 27190 7638 27225 7639
rect 27169 7631 27225 7638
rect 27169 7611 27198 7631
rect 27218 7611 27225 7631
rect 27169 7606 27225 7611
rect 27616 7634 27648 7641
rect 27616 7614 27622 7634
rect 27643 7614 27648 7634
rect 27169 7328 27203 7606
rect 27616 7586 27648 7614
rect 30612 7622 30692 7634
rect 30793 7629 30828 7630
rect 30612 7596 30628 7622
rect 30668 7596 30692 7622
rect 27236 7578 27648 7586
rect 27236 7552 27242 7578
rect 27268 7552 27648 7578
rect 27236 7550 27648 7552
rect 27238 7549 27278 7550
rect 27405 7524 27436 7532
rect 27405 7494 27409 7524
rect 27430 7494 27436 7524
rect 27169 7320 27204 7328
rect 27169 7300 27177 7320
rect 27197 7300 27204 7320
rect 27405 7309 27436 7494
rect 27616 7485 27648 7550
rect 28030 7583 28141 7590
rect 28030 7582 28109 7583
rect 28030 7558 28052 7582
rect 28076 7559 28109 7582
rect 28133 7559 28141 7583
rect 28076 7558 28141 7559
rect 28030 7548 28141 7558
rect 30612 7577 30692 7596
rect 30612 7551 30631 7577
rect 30671 7551 30692 7577
rect 28091 7531 28140 7548
rect 30612 7524 30692 7551
rect 30612 7498 30635 7524
rect 30675 7498 30692 7524
rect 30612 7487 30692 7498
rect 30772 7622 30828 7629
rect 30772 7602 30801 7622
rect 30821 7602 30828 7622
rect 30772 7597 30828 7602
rect 31219 7625 31251 7632
rect 31219 7605 31225 7625
rect 31246 7605 31251 7625
rect 27616 7465 27620 7485
rect 27641 7465 27648 7485
rect 27616 7458 27648 7465
rect 27925 7402 28026 7403
rect 27823 7389 28026 7402
rect 27823 7387 27966 7389
rect 27823 7384 27900 7387
rect 27823 7357 27826 7384
rect 27855 7360 27900 7384
rect 27929 7360 27966 7387
rect 27855 7357 27966 7360
rect 27823 7356 27966 7357
rect 28002 7356 28026 7389
rect 27823 7343 28026 7356
rect 27169 7295 27204 7300
rect 27169 7294 27201 7295
rect 27403 7232 27437 7309
rect 26036 5829 26633 5833
rect 23136 5751 23171 5753
rect 23136 5742 23240 5751
rect 23136 5741 23187 5742
rect 23136 5721 23139 5741
rect 23164 5722 23187 5741
rect 23219 5722 23240 5742
rect 23164 5721 23240 5722
rect 23136 5714 23240 5721
rect 23136 5702 23171 5714
rect 22548 5636 22751 5649
rect 22548 5603 22572 5636
rect 22608 5635 22751 5636
rect 22608 5632 22719 5635
rect 22608 5605 22645 5632
rect 22674 5608 22719 5632
rect 22748 5608 22751 5635
rect 22674 5605 22751 5608
rect 22608 5603 22751 5605
rect 22548 5590 22751 5603
rect 22548 5589 22649 5590
rect 22926 5527 22958 5534
rect 22926 5507 22933 5527
rect 22954 5507 22958 5527
rect 22437 5449 22502 5458
rect 22437 5412 22447 5449
rect 22487 5415 22502 5449
rect 22926 5442 22958 5507
rect 23138 5498 23169 5702
rect 23373 5697 23405 5698
rect 23370 5692 23405 5697
rect 23370 5672 23377 5692
rect 23397 5672 23405 5692
rect 23370 5664 23405 5672
rect 23138 5468 23144 5498
rect 23165 5468 23169 5498
rect 23138 5460 23169 5468
rect 23296 5442 23336 5443
rect 22926 5440 23338 5442
rect 22487 5412 22504 5415
rect 22437 5393 22504 5412
rect 22437 5372 22451 5393
rect 22487 5372 22504 5393
rect 22437 5365 22504 5372
rect 22926 5414 23306 5440
rect 23332 5414 23338 5440
rect 22926 5406 23338 5414
rect 22926 5378 22958 5406
rect 23371 5386 23405 5664
rect 23495 5496 23560 5796
rect 25673 5784 26633 5829
rect 26740 6172 26776 6800
rect 25673 5780 26086 5784
rect 25673 5691 25707 5780
rect 25911 5694 25943 5695
rect 25086 5633 25289 5646
rect 25086 5600 25110 5633
rect 25146 5632 25289 5633
rect 25146 5629 25257 5632
rect 25146 5602 25183 5629
rect 25212 5605 25257 5629
rect 25286 5605 25289 5632
rect 25212 5602 25289 5605
rect 25146 5600 25289 5602
rect 25086 5587 25289 5600
rect 25086 5586 25187 5587
rect 25464 5524 25496 5531
rect 25464 5504 25471 5524
rect 25492 5504 25496 5524
rect 22926 5358 22931 5378
rect 22952 5358 22958 5378
rect 22926 5351 22958 5358
rect 23349 5381 23405 5386
rect 23349 5361 23356 5381
rect 23376 5361 23405 5381
rect 23349 5354 23405 5361
rect 23485 5485 23565 5496
rect 23485 5459 23502 5485
rect 23542 5459 23565 5485
rect 23485 5432 23565 5459
rect 23485 5406 23506 5432
rect 23546 5406 23565 5432
rect 23485 5387 23565 5406
rect 23485 5361 23509 5387
rect 23549 5361 23565 5387
rect 23349 5353 23384 5354
rect 23485 5349 23565 5361
rect 25464 5439 25496 5504
rect 25676 5495 25707 5691
rect 25908 5689 25943 5694
rect 25908 5669 25915 5689
rect 25935 5669 25943 5689
rect 25908 5661 25943 5669
rect 25676 5465 25682 5495
rect 25703 5465 25707 5495
rect 25676 5457 25707 5465
rect 25834 5439 25874 5440
rect 25464 5437 25876 5439
rect 25464 5411 25844 5437
rect 25870 5411 25876 5437
rect 25464 5403 25876 5411
rect 25464 5375 25496 5403
rect 25909 5383 25943 5661
rect 25464 5355 25469 5375
rect 25490 5355 25496 5375
rect 25464 5348 25496 5355
rect 25887 5378 25943 5383
rect 25887 5358 25894 5378
rect 25914 5358 25943 5378
rect 25887 5351 25943 5358
rect 25887 5350 25922 5351
rect 22640 5298 22751 5302
rect 24395 5298 24602 5299
rect 25178 5298 25289 5299
rect 21960 5280 26026 5298
rect 21960 5260 22648 5280
rect 22667 5260 22725 5280
rect 22744 5277 26026 5280
rect 22744 5260 25186 5277
rect 21960 5257 25186 5260
rect 25205 5257 25263 5277
rect 25282 5257 26026 5277
rect 21960 5242 26026 5257
rect 21962 5054 22069 5242
rect 24557 5240 26026 5242
rect 22430 5203 22551 5213
rect 22430 5201 22499 5203
rect 22430 5160 22443 5201
rect 22480 5162 22499 5201
rect 22536 5162 22551 5203
rect 22480 5160 22551 5162
rect 22430 5142 22551 5160
rect 21962 5050 22070 5054
rect 22436 5050 22513 5142
rect 23486 5138 23562 5154
rect 23486 5115 23501 5138
rect 19712 4874 19727 4897
rect 19651 4858 19727 4874
rect 20700 4870 20777 4962
rect 21143 4958 21251 4962
rect 20662 4852 20783 4870
rect 20662 4850 20733 4852
rect 20662 4809 20677 4850
rect 20714 4811 20733 4850
rect 20770 4811 20783 4852
rect 20714 4809 20783 4811
rect 20662 4799 20783 4809
rect 17233 4770 18656 4772
rect 21144 4770 21251 4958
rect 17233 4755 21253 4770
rect 17233 4735 17931 4755
rect 17950 4735 18008 4755
rect 18027 4752 21253 4755
rect 18027 4735 20469 4752
rect 17233 4732 20469 4735
rect 20488 4732 20546 4752
rect 20565 4732 21253 4752
rect 17233 4714 21253 4732
rect 17924 4713 18035 4714
rect 18611 4713 18818 4714
rect 20462 4710 20573 4714
rect 17291 4661 17326 4662
rect 17270 4654 17326 4661
rect 17270 4634 17299 4654
rect 17319 4634 17326 4654
rect 17270 4629 17326 4634
rect 17717 4657 17749 4664
rect 17717 4637 17723 4657
rect 17744 4637 17749 4657
rect 16439 4405 16465 4420
rect 16436 4398 16472 4405
rect 16436 4360 16442 4398
rect 16465 4360 16472 4398
rect 16436 4354 16472 4360
rect 17270 4351 17304 4629
rect 17717 4609 17749 4637
rect 17337 4601 17749 4609
rect 17337 4575 17343 4601
rect 17369 4575 17749 4601
rect 17337 4573 17749 4575
rect 17339 4572 17379 4573
rect 17506 4547 17537 4555
rect 17506 4517 17510 4547
rect 17531 4517 17537 4547
rect 17270 4343 17305 4351
rect 17270 4323 17278 4343
rect 17298 4323 17305 4343
rect 17270 4318 17305 4323
rect 17270 4317 17302 4318
rect 17506 4314 17537 4517
rect 17717 4508 17749 4573
rect 19648 4651 19728 4663
rect 19829 4658 19864 4659
rect 19648 4625 19664 4651
rect 19704 4625 19728 4651
rect 19648 4606 19728 4625
rect 19648 4580 19667 4606
rect 19707 4580 19728 4606
rect 19648 4553 19728 4580
rect 19648 4527 19671 4553
rect 19711 4527 19728 4553
rect 19648 4516 19728 4527
rect 19808 4651 19864 4658
rect 19808 4631 19837 4651
rect 19857 4631 19864 4651
rect 19808 4626 19864 4631
rect 20255 4654 20287 4661
rect 20255 4634 20261 4654
rect 20282 4634 20287 4654
rect 17717 4488 17721 4508
rect 17742 4488 17749 4508
rect 17717 4481 17749 4488
rect 18026 4425 18127 4426
rect 17924 4412 18127 4425
rect 17924 4410 18067 4412
rect 17924 4407 18001 4410
rect 17924 4380 17927 4407
rect 17956 4383 18001 4407
rect 18030 4383 18067 4410
rect 17956 4380 18067 4383
rect 17924 4379 18067 4380
rect 18103 4379 18127 4412
rect 17924 4366 18127 4379
rect 17501 4296 17537 4314
rect 17501 4279 17536 4296
rect 17434 4248 17539 4279
rect 17434 4243 17506 4248
rect 17434 4222 17465 4243
rect 17485 4227 17506 4243
rect 17526 4227 17539 4248
rect 17485 4222 17539 4227
rect 17434 4213 17539 4222
rect 19653 4216 19718 4516
rect 19808 4348 19842 4626
rect 20255 4606 20287 4634
rect 19875 4598 20287 4606
rect 19875 4572 19881 4598
rect 19907 4572 20287 4598
rect 20709 4640 20776 4647
rect 20709 4619 20726 4640
rect 20762 4619 20776 4640
rect 20709 4600 20776 4619
rect 20709 4597 20726 4600
rect 19875 4570 20287 4572
rect 19877 4569 19917 4570
rect 20044 4544 20075 4552
rect 20044 4514 20048 4544
rect 20069 4514 20075 4544
rect 19808 4340 19843 4348
rect 19808 4320 19816 4340
rect 19836 4320 19843 4340
rect 19808 4315 19843 4320
rect 19808 4314 19840 4315
rect 20044 4310 20075 4514
rect 20255 4505 20287 4570
rect 20711 4563 20726 4597
rect 20766 4563 20776 4600
rect 20711 4554 20776 4563
rect 20255 4485 20259 4505
rect 20280 4485 20287 4505
rect 20255 4478 20287 4485
rect 20564 4422 20665 4423
rect 20462 4409 20665 4422
rect 20462 4407 20605 4409
rect 20462 4404 20539 4407
rect 20462 4377 20465 4404
rect 20494 4380 20539 4404
rect 20568 4380 20605 4407
rect 20494 4377 20605 4380
rect 20462 4376 20605 4377
rect 20641 4376 20665 4409
rect 20462 4363 20665 4376
rect 20042 4298 20077 4310
rect 19973 4291 20077 4298
rect 19973 4290 20049 4291
rect 19973 4270 19994 4290
rect 20026 4271 20049 4290
rect 20074 4271 20077 4291
rect 20026 4270 20077 4271
rect 19973 4261 20077 4270
rect 20042 4259 20077 4261
rect 19653 4177 19656 4216
rect 19701 4177 19718 4216
rect 20714 4193 20765 4554
rect 20712 4191 20769 4193
rect 19653 4155 19718 4177
rect 20701 4179 20769 4191
rect 20701 4146 20712 4179
rect 20752 4146 20769 4179
rect 20701 4140 20769 4146
rect 20701 4136 20765 4140
rect 19414 4091 19525 4094
rect 21144 4091 21251 4714
rect 17457 4077 21251 4091
rect 17457 4057 19421 4077
rect 19440 4057 19498 4077
rect 19517 4073 21251 4077
rect 19517 4057 20469 4073
rect 17457 4053 20469 4057
rect 20488 4053 20546 4073
rect 20565 4053 21251 4073
rect 17457 4035 21251 4053
rect 17457 4034 18698 4035
rect 20462 4031 20573 4035
rect 18781 3983 18816 3984
rect 18760 3976 18816 3983
rect 18760 3956 18789 3976
rect 18809 3956 18816 3976
rect 18760 3951 18816 3956
rect 19207 3979 19239 3986
rect 19829 3979 19864 3980
rect 19207 3959 19213 3979
rect 19234 3959 19239 3979
rect 19808 3972 19864 3979
rect 19673 3962 19731 3967
rect 18760 3673 18794 3951
rect 19207 3931 19239 3959
rect 18827 3923 19239 3931
rect 18827 3897 18833 3923
rect 18859 3897 19239 3923
rect 18827 3895 19239 3897
rect 18829 3894 18869 3895
rect 18996 3869 19027 3877
rect 18996 3839 19000 3869
rect 19021 3839 19027 3869
rect 18760 3665 18795 3673
rect 18760 3645 18768 3665
rect 18788 3645 18795 3665
rect 18760 3640 18795 3645
rect 17501 3629 17537 3640
rect 18760 3639 18792 3640
rect 18996 3632 19027 3839
rect 19207 3830 19239 3895
rect 19207 3810 19211 3830
rect 19232 3810 19239 3830
rect 19207 3803 19239 3810
rect 19656 3953 19731 3962
rect 19656 3920 19665 3953
rect 19718 3920 19731 3953
rect 19656 3895 19731 3920
rect 19656 3862 19670 3895
rect 19723 3862 19731 3895
rect 19656 3856 19731 3862
rect 19808 3952 19837 3972
rect 19857 3952 19864 3972
rect 19808 3947 19864 3952
rect 20255 3975 20287 3982
rect 20255 3955 20261 3975
rect 20282 3955 20287 3975
rect 19516 3747 19617 3748
rect 19414 3734 19617 3747
rect 19414 3732 19557 3734
rect 19414 3729 19491 3732
rect 19414 3702 19417 3729
rect 19446 3705 19491 3729
rect 19520 3705 19557 3732
rect 19446 3702 19557 3705
rect 19414 3701 19557 3702
rect 19593 3701 19617 3734
rect 19414 3688 19617 3701
rect 17501 3606 17507 3629
rect 17531 3606 17537 3629
rect 18991 3623 19027 3632
rect 18936 3613 19033 3623
rect 17748 3611 19033 3613
rect 17501 3585 17537 3606
rect 17501 3562 17507 3585
rect 17531 3562 17537 3585
rect 17501 3409 17537 3562
rect 17713 3601 19033 3611
rect 17713 3563 17725 3601
rect 17750 3566 17769 3601
rect 17794 3566 19033 3601
rect 17750 3563 19033 3566
rect 17713 3560 19033 3563
rect 17713 3558 19030 3560
rect 17713 3555 17802 3558
rect 17729 3554 17801 3555
rect 19656 3545 19726 3856
rect 19808 3669 19842 3947
rect 20255 3927 20287 3955
rect 19875 3919 20287 3927
rect 19875 3893 19881 3919
rect 19907 3893 20287 3919
rect 19875 3891 20287 3893
rect 19877 3890 19917 3891
rect 20044 3865 20075 3873
rect 20044 3835 20048 3865
rect 20069 3835 20075 3865
rect 19808 3661 19843 3669
rect 19808 3641 19816 3661
rect 19836 3641 19843 3661
rect 19808 3636 19843 3641
rect 20044 3636 20075 3835
rect 20255 3826 20287 3891
rect 20255 3806 20259 3826
rect 20280 3806 20287 3826
rect 20255 3799 20287 3806
rect 20700 3952 20772 3970
rect 20700 3910 20713 3952
rect 20762 3910 20772 3952
rect 20700 3889 20772 3910
rect 20700 3847 20714 3889
rect 20763 3847 20772 3889
rect 20564 3743 20665 3744
rect 20462 3730 20665 3743
rect 20462 3728 20605 3730
rect 20462 3725 20539 3728
rect 20462 3698 20465 3725
rect 20494 3701 20539 3725
rect 20568 3701 20605 3728
rect 20494 3698 20605 3701
rect 20462 3697 20605 3698
rect 20641 3697 20665 3730
rect 20462 3684 20665 3697
rect 19808 3635 19840 3636
rect 20042 3633 20075 3636
rect 20008 3614 20076 3633
rect 19978 3602 20077 3614
rect 20700 3606 20772 3847
rect 21144 3606 21251 4035
rect 21963 4457 22070 5050
rect 22438 4999 22513 5050
rect 23479 5101 23501 5115
rect 23545 5101 23562 5138
rect 23479 5081 23562 5101
rect 23479 5015 23496 5081
rect 23550 5015 23562 5081
rect 22438 4956 22514 4999
rect 22442 4645 22514 4956
rect 23479 4991 23562 5015
rect 23479 4971 23555 4991
rect 23479 4952 23558 4971
rect 23138 4936 23210 4937
rect 23137 4928 23236 4936
rect 23137 4925 23189 4928
rect 23137 4890 23145 4925
rect 23170 4890 23189 4925
rect 23214 4890 23236 4928
rect 23137 4878 23236 4890
rect 23138 4859 23206 4878
rect 23139 4856 23172 4859
rect 23374 4856 23406 4857
rect 22549 4795 22752 4808
rect 22549 4762 22573 4795
rect 22609 4794 22752 4795
rect 22609 4791 22720 4794
rect 22609 4764 22646 4791
rect 22675 4767 22720 4791
rect 22749 4767 22752 4794
rect 22675 4764 22752 4767
rect 22609 4762 22752 4764
rect 22549 4749 22752 4762
rect 22549 4748 22650 4749
rect 22442 4603 22451 4645
rect 22500 4603 22514 4645
rect 22442 4582 22514 4603
rect 22442 4540 22452 4582
rect 22501 4540 22514 4582
rect 22442 4522 22514 4540
rect 22927 4686 22959 4693
rect 22927 4666 22934 4686
rect 22955 4666 22959 4686
rect 22927 4601 22959 4666
rect 23139 4657 23170 4856
rect 23371 4851 23406 4856
rect 23371 4831 23378 4851
rect 23398 4831 23406 4851
rect 23371 4823 23406 4831
rect 23139 4627 23145 4657
rect 23166 4627 23170 4657
rect 23139 4619 23170 4627
rect 23297 4601 23337 4602
rect 22927 4599 23339 4601
rect 22927 4573 23307 4599
rect 23333 4573 23339 4599
rect 22927 4565 23339 4573
rect 22927 4537 22959 4565
rect 23372 4545 23406 4823
rect 23488 4636 23558 4952
rect 25476 4937 25507 4938
rect 25476 4929 25521 4937
rect 24556 4906 24720 4913
rect 25476 4906 25486 4929
rect 24182 4891 25486 4906
rect 25511 4891 25521 4929
rect 26740 4932 26774 6172
rect 26740 4928 26970 4932
rect 26740 4902 26939 4928
rect 26964 4902 26970 4928
rect 26740 4894 26970 4902
rect 24182 4873 25521 4891
rect 24187 4860 24223 4873
rect 24556 4870 24720 4873
rect 23597 4791 23800 4804
rect 23597 4758 23621 4791
rect 23657 4790 23800 4791
rect 23657 4787 23768 4790
rect 23657 4760 23694 4787
rect 23723 4763 23768 4787
rect 23797 4763 23800 4790
rect 23723 4760 23800 4763
rect 23657 4758 23800 4760
rect 23597 4745 23800 4758
rect 23597 4744 23698 4745
rect 22927 4517 22932 4537
rect 22953 4517 22959 4537
rect 22927 4510 22959 4517
rect 23350 4540 23406 4545
rect 23350 4520 23357 4540
rect 23377 4520 23406 4540
rect 23483 4630 23558 4636
rect 23483 4597 23491 4630
rect 23544 4597 23558 4630
rect 23483 4572 23558 4597
rect 23483 4539 23496 4572
rect 23549 4539 23558 4572
rect 23483 4530 23558 4539
rect 23975 4682 24007 4689
rect 23975 4662 23982 4682
rect 24003 4662 24007 4682
rect 23975 4597 24007 4662
rect 24187 4653 24218 4860
rect 24422 4852 24454 4853
rect 24419 4847 24454 4852
rect 24419 4827 24426 4847
rect 24446 4827 24454 4847
rect 24419 4819 24454 4827
rect 24187 4623 24193 4653
rect 24214 4623 24218 4653
rect 24187 4615 24218 4623
rect 24345 4597 24385 4598
rect 23975 4595 24387 4597
rect 23975 4569 24355 4595
rect 24381 4569 24387 4595
rect 23975 4561 24387 4569
rect 23975 4533 24007 4561
rect 24420 4541 24454 4819
rect 26499 4797 26702 4810
rect 26499 4764 26523 4797
rect 26559 4796 26702 4797
rect 26559 4793 26670 4796
rect 26559 4766 26596 4793
rect 26625 4769 26670 4793
rect 26699 4769 26702 4796
rect 26625 4766 26702 4769
rect 26559 4764 26702 4766
rect 26499 4751 26702 4764
rect 26499 4750 26600 4751
rect 23483 4525 23541 4530
rect 23350 4513 23406 4520
rect 23975 4513 23980 4533
rect 24001 4513 24007 4533
rect 23350 4512 23385 4513
rect 23975 4506 24007 4513
rect 24398 4536 24454 4541
rect 24398 4516 24405 4536
rect 24425 4516 24454 4536
rect 24398 4509 24454 4516
rect 26877 4688 26909 4695
rect 26877 4668 26884 4688
rect 26905 4668 26909 4688
rect 26877 4603 26909 4668
rect 27089 4659 27120 4859
rect 27324 4858 27356 4859
rect 27321 4853 27356 4858
rect 27321 4833 27328 4853
rect 27348 4833 27356 4853
rect 27321 4825 27356 4833
rect 27089 4629 27095 4659
rect 27116 4629 27120 4659
rect 27089 4621 27120 4629
rect 27247 4603 27287 4604
rect 26877 4601 27289 4603
rect 26877 4575 27257 4601
rect 27283 4575 27289 4601
rect 26877 4567 27289 4575
rect 26877 4539 26909 4567
rect 26877 4519 26882 4539
rect 26903 4519 26909 4539
rect 26877 4512 26909 4519
rect 27079 4541 27127 4548
rect 27322 4547 27356 4825
rect 27079 4521 27086 4541
rect 27119 4521 27127 4541
rect 24398 4508 24433 4509
rect 22641 4457 22752 4461
rect 24424 4457 25994 4458
rect 21963 4453 25994 4457
rect 26319 4453 26737 4466
rect 21963 4441 26737 4453
rect 21963 4439 26599 4441
rect 21963 4419 22649 4439
rect 22668 4419 22726 4439
rect 22745 4435 26599 4439
rect 22745 4419 23697 4435
rect 21963 4415 23697 4419
rect 23716 4415 23774 4435
rect 23793 4421 26599 4435
rect 26618 4421 26676 4441
rect 26695 4421 26737 4441
rect 23793 4415 26737 4421
rect 21963 4401 26737 4415
rect 21963 3778 22070 4401
rect 23689 4398 23800 4401
rect 26319 4395 26737 4401
rect 22449 4352 22513 4356
rect 22445 4346 22513 4352
rect 22445 4313 22462 4346
rect 22502 4313 22513 4346
rect 22445 4301 22513 4313
rect 23496 4315 23561 4337
rect 22445 4299 22502 4301
rect 22449 3938 22500 4299
rect 23496 4276 23513 4315
rect 23558 4276 23561 4315
rect 23137 4231 23172 4233
rect 23137 4222 23241 4231
rect 23137 4221 23188 4222
rect 23137 4201 23140 4221
rect 23165 4202 23188 4221
rect 23220 4202 23241 4222
rect 23165 4201 23241 4202
rect 23137 4194 23241 4201
rect 23137 4182 23172 4194
rect 22549 4116 22752 4129
rect 22549 4083 22573 4116
rect 22609 4115 22752 4116
rect 22609 4112 22720 4115
rect 22609 4085 22646 4112
rect 22675 4088 22720 4112
rect 22749 4088 22752 4115
rect 22675 4085 22752 4088
rect 22609 4083 22752 4085
rect 22549 4070 22752 4083
rect 22549 4069 22650 4070
rect 22927 4007 22959 4014
rect 22927 3987 22934 4007
rect 22955 3987 22959 4007
rect 22438 3929 22503 3938
rect 22438 3892 22448 3929
rect 22488 3895 22503 3929
rect 22927 3922 22959 3987
rect 23139 3978 23170 4182
rect 23374 4177 23406 4178
rect 23371 4172 23406 4177
rect 23371 4152 23378 4172
rect 23398 4152 23406 4172
rect 23371 4144 23406 4152
rect 23139 3948 23145 3978
rect 23166 3948 23170 3978
rect 23139 3940 23170 3948
rect 23297 3922 23337 3923
rect 22927 3920 23339 3922
rect 22488 3892 22505 3895
rect 22438 3873 22505 3892
rect 22438 3852 22452 3873
rect 22488 3852 22505 3873
rect 22438 3845 22505 3852
rect 22927 3894 23307 3920
rect 23333 3894 23339 3920
rect 22927 3886 23339 3894
rect 22927 3858 22959 3886
rect 23372 3866 23406 4144
rect 23496 3976 23561 4276
rect 25633 4237 25670 4258
rect 25633 4200 25644 4237
rect 25661 4213 25670 4237
rect 25661 4200 25671 4213
rect 25633 4190 25671 4200
rect 25634 4186 25671 4190
rect 25634 4180 25667 4186
rect 25044 4111 25247 4124
rect 25044 4078 25068 4111
rect 25104 4110 25247 4111
rect 25104 4107 25215 4110
rect 25104 4080 25141 4107
rect 25170 4083 25215 4107
rect 25244 4083 25247 4110
rect 25170 4080 25247 4083
rect 25104 4078 25247 4080
rect 25044 4065 25247 4078
rect 25044 4064 25145 4065
rect 25422 4002 25454 4009
rect 25422 3982 25429 4002
rect 25450 3982 25454 4002
rect 22927 3838 22932 3858
rect 22953 3838 22959 3858
rect 22927 3831 22959 3838
rect 23350 3861 23406 3866
rect 23350 3841 23357 3861
rect 23377 3841 23406 3861
rect 23350 3834 23406 3841
rect 23486 3965 23566 3976
rect 23486 3939 23503 3965
rect 23543 3939 23566 3965
rect 23486 3912 23566 3939
rect 23486 3886 23507 3912
rect 23547 3886 23566 3912
rect 23486 3867 23566 3886
rect 23486 3841 23510 3867
rect 23550 3841 23566 3867
rect 24560 3911 24665 3932
rect 25422 3917 25454 3982
rect 25634 3973 25665 4180
rect 25869 4172 25901 4173
rect 25866 4167 25901 4172
rect 25866 4147 25873 4167
rect 25893 4147 25901 4167
rect 25866 4139 25901 4147
rect 25634 3943 25640 3973
rect 25661 3943 25665 3973
rect 25634 3935 25665 3943
rect 25792 3917 25832 3918
rect 25422 3915 25834 3917
rect 24560 3905 25036 3911
rect 24560 3903 24617 3905
rect 24560 3872 24572 3903
rect 24597 3882 24617 3903
rect 24643 3898 25036 3905
rect 24643 3882 24997 3898
rect 24597 3875 24997 3882
rect 25023 3875 25036 3898
rect 24597 3872 25036 3875
rect 24560 3862 25036 3872
rect 25422 3889 25802 3915
rect 25828 3889 25834 3915
rect 25422 3881 25834 3889
rect 24560 3860 24665 3862
rect 23350 3833 23385 3834
rect 23486 3829 23566 3841
rect 25422 3853 25454 3881
rect 25867 3861 25901 4139
rect 25422 3833 25427 3853
rect 25448 3833 25454 3853
rect 25422 3826 25454 3833
rect 25845 3856 25901 3861
rect 25845 3836 25852 3856
rect 25872 3836 25901 3856
rect 25845 3829 25901 3836
rect 25845 3828 25880 3829
rect 22641 3778 22752 3782
rect 24383 3778 26036 3781
rect 21961 3760 26036 3778
rect 21961 3740 22649 3760
rect 22668 3740 22726 3760
rect 22745 3755 26036 3760
rect 22745 3740 25144 3755
rect 21961 3735 25144 3740
rect 25163 3735 25221 3755
rect 25240 3735 26036 3755
rect 21961 3725 26036 3735
rect 21961 3722 22586 3725
rect 22773 3722 26036 3725
rect 19978 3564 20000 3602
rect 20025 3567 20044 3602
rect 20069 3567 20077 3602
rect 20025 3564 20077 3567
rect 19978 3556 20077 3564
rect 20004 3555 20076 3556
rect 19655 3529 19726 3545
rect 19655 3513 19675 3529
rect 19656 3483 19675 3513
rect 19658 3463 19675 3483
rect 19705 3483 19726 3529
rect 20698 3525 20776 3606
rect 21143 3551 21251 3606
rect 19705 3463 19725 3483
rect 19658 3444 19725 3463
rect 20698 3423 20777 3525
rect 17492 3400 17578 3409
rect 17492 3382 17511 3400
rect 17563 3382 17578 3400
rect 17492 3378 17578 3382
rect 20662 3405 20783 3423
rect 20662 3403 20733 3405
rect 20662 3362 20677 3403
rect 20714 3364 20733 3403
rect 20770 3364 20783 3405
rect 20714 3362 20783 3364
rect 20662 3352 20783 3362
rect 17967 3324 18078 3327
rect 17282 3323 18831 3324
rect 21144 3323 21251 3551
rect 21963 3494 22070 3722
rect 24383 3721 26036 3722
rect 25136 3718 25247 3721
rect 22431 3683 22552 3693
rect 22431 3681 22500 3683
rect 22431 3640 22444 3681
rect 22481 3642 22500 3681
rect 22537 3642 22552 3683
rect 22481 3640 22552 3642
rect 22431 3622 22552 3640
rect 22437 3520 22516 3622
rect 23489 3582 23556 3601
rect 23489 3562 23509 3582
rect 21963 3439 22071 3494
rect 22438 3439 22516 3520
rect 23488 3516 23509 3562
rect 23539 3562 23556 3582
rect 23539 3532 23558 3562
rect 23539 3516 23559 3532
rect 23488 3500 23559 3516
rect 23138 3489 23210 3490
rect 23137 3481 23236 3489
rect 23137 3478 23189 3481
rect 23137 3443 23145 3478
rect 23170 3443 23189 3478
rect 23214 3443 23236 3481
rect 17282 3320 20441 3323
rect 20628 3320 21253 3323
rect 17282 3310 21253 3320
rect 17282 3290 17974 3310
rect 17993 3290 18051 3310
rect 18070 3305 21253 3310
rect 18070 3290 20469 3305
rect 17282 3285 20469 3290
rect 20488 3285 20546 3305
rect 20565 3285 21253 3305
rect 17282 3267 21253 3285
rect 17282 3264 18831 3267
rect 20462 3263 20573 3267
rect 17334 3216 17369 3217
rect 17313 3209 17369 3216
rect 17313 3189 17342 3209
rect 17362 3189 17369 3209
rect 17313 3184 17369 3189
rect 17760 3212 17792 3219
rect 17760 3192 17766 3212
rect 17787 3192 17792 3212
rect 17313 2906 17347 3184
rect 17760 3164 17792 3192
rect 17380 3156 17792 3164
rect 17380 3130 17386 3156
rect 17412 3130 17792 3156
rect 17380 3128 17792 3130
rect 17382 3127 17422 3128
rect 17549 3102 17580 3110
rect 17549 3072 17553 3102
rect 17574 3072 17580 3102
rect 17313 2898 17348 2906
rect 17313 2878 17321 2898
rect 17341 2878 17348 2898
rect 17313 2873 17348 2878
rect 17313 2872 17345 2873
rect 17549 2871 17580 3072
rect 17760 3063 17792 3128
rect 17760 3043 17764 3063
rect 17785 3043 17792 3063
rect 17760 3036 17792 3043
rect 18354 3203 18447 3210
rect 18354 3162 18378 3203
rect 18432 3162 18447 3203
rect 18069 2980 18170 2981
rect 17967 2967 18170 2980
rect 17967 2965 18110 2967
rect 17967 2962 18044 2965
rect 17967 2935 17970 2962
rect 17999 2938 18044 2962
rect 18073 2938 18110 2965
rect 17999 2935 18110 2938
rect 17967 2934 18110 2935
rect 18146 2934 18170 2967
rect 17967 2921 18170 2934
rect 18354 2789 18447 3162
rect 19648 3204 19728 3216
rect 19829 3211 19864 3212
rect 19648 3178 19664 3204
rect 19704 3178 19728 3204
rect 19648 3159 19728 3178
rect 19648 3133 19667 3159
rect 19707 3133 19728 3159
rect 19648 3106 19728 3133
rect 19648 3080 19671 3106
rect 19711 3080 19728 3106
rect 19648 3069 19728 3080
rect 19808 3204 19864 3211
rect 19808 3184 19837 3204
rect 19857 3184 19864 3204
rect 19808 3179 19864 3184
rect 20255 3207 20287 3214
rect 20255 3187 20261 3207
rect 20282 3187 20287 3207
rect 18354 2745 18372 2789
rect 18432 2745 18447 2789
rect 18354 2730 18447 2745
rect 19653 2769 19718 3069
rect 19808 2901 19842 3179
rect 20255 3159 20287 3187
rect 19875 3151 20287 3159
rect 19875 3125 19881 3151
rect 19907 3125 20287 3151
rect 20709 3193 20776 3200
rect 20709 3172 20726 3193
rect 20762 3172 20776 3193
rect 20709 3153 20776 3172
rect 20709 3150 20726 3153
rect 19875 3123 20287 3125
rect 19877 3122 19917 3123
rect 20044 3097 20075 3105
rect 20044 3067 20048 3097
rect 20069 3067 20075 3097
rect 19808 2893 19843 2901
rect 19808 2873 19816 2893
rect 19836 2873 19843 2893
rect 19808 2868 19843 2873
rect 19808 2867 19840 2868
rect 20044 2863 20075 3067
rect 20255 3058 20287 3123
rect 20711 3116 20726 3150
rect 20766 3116 20776 3153
rect 20711 3107 20776 3116
rect 20255 3038 20259 3058
rect 20280 3038 20287 3058
rect 20255 3031 20287 3038
rect 20564 2975 20665 2976
rect 20462 2962 20665 2975
rect 20462 2960 20605 2962
rect 20462 2957 20539 2960
rect 20462 2930 20465 2957
rect 20494 2933 20539 2957
rect 20568 2933 20605 2960
rect 20494 2930 20605 2933
rect 20462 2929 20605 2930
rect 20641 2929 20665 2962
rect 20462 2916 20665 2929
rect 20042 2851 20077 2863
rect 19973 2844 20077 2851
rect 19973 2843 20049 2844
rect 19973 2823 19994 2843
rect 20026 2824 20049 2843
rect 20074 2824 20077 2844
rect 20026 2823 20077 2824
rect 19973 2814 20077 2823
rect 20042 2812 20077 2814
rect 19653 2730 19656 2769
rect 19701 2730 19718 2769
rect 20714 2746 20765 3107
rect 20712 2744 20769 2746
rect 19653 2708 19718 2730
rect 20701 2732 20769 2744
rect 20701 2699 20712 2732
rect 20752 2699 20769 2732
rect 20701 2693 20769 2699
rect 20701 2689 20765 2693
rect 19414 2644 19525 2647
rect 21144 2644 21251 3267
rect 17677 2630 21251 2644
rect 17677 2610 19421 2630
rect 19440 2610 19498 2630
rect 19517 2626 21251 2630
rect 19517 2610 20469 2626
rect 17677 2606 20469 2610
rect 20488 2606 20546 2626
rect 20565 2606 21251 2626
rect 17677 2588 21251 2606
rect 17677 2587 18790 2588
rect 20462 2584 20573 2588
rect 18781 2536 18816 2537
rect 18760 2529 18816 2536
rect 18760 2509 18789 2529
rect 18809 2509 18816 2529
rect 18760 2504 18816 2509
rect 19207 2532 19239 2539
rect 19829 2532 19864 2533
rect 19207 2512 19213 2532
rect 19234 2512 19239 2532
rect 19808 2525 19864 2532
rect 19673 2515 19731 2520
rect 16596 2469 18449 2502
rect 16596 2404 16661 2469
rect 16792 2449 18449 2469
rect 16792 2408 18385 2449
rect 18421 2408 18449 2449
rect 18547 2469 18611 2488
rect 18547 2430 18564 2469
rect 18598 2430 18611 2469
rect 18547 2411 18611 2430
rect 16792 2404 18449 2408
rect 16596 2379 18449 2404
rect 18360 2376 18442 2379
rect 18549 1899 18611 2411
rect 18760 2226 18794 2504
rect 19207 2484 19239 2512
rect 18827 2476 19239 2484
rect 18827 2450 18833 2476
rect 18859 2450 19239 2476
rect 18827 2448 19239 2450
rect 18829 2447 18869 2448
rect 18996 2422 19027 2430
rect 18996 2392 19000 2422
rect 19021 2392 19027 2422
rect 18760 2218 18795 2226
rect 18760 2198 18768 2218
rect 18788 2198 18795 2218
rect 18760 2193 18795 2198
rect 18760 2192 18792 2193
rect 18996 2185 19027 2392
rect 19207 2383 19239 2448
rect 19207 2363 19211 2383
rect 19232 2363 19239 2383
rect 19207 2356 19239 2363
rect 19656 2506 19731 2515
rect 19656 2473 19665 2506
rect 19718 2473 19731 2506
rect 19656 2448 19731 2473
rect 19656 2415 19670 2448
rect 19723 2415 19731 2448
rect 19656 2409 19731 2415
rect 19808 2505 19837 2525
rect 19857 2505 19864 2525
rect 19808 2500 19864 2505
rect 20255 2528 20287 2535
rect 20255 2508 20261 2528
rect 20282 2508 20287 2528
rect 19516 2300 19617 2301
rect 19414 2287 19617 2300
rect 19414 2285 19557 2287
rect 19414 2282 19491 2285
rect 19414 2255 19417 2282
rect 19446 2258 19491 2282
rect 19520 2258 19557 2285
rect 19446 2255 19557 2258
rect 19414 2254 19557 2255
rect 19593 2254 19617 2287
rect 19414 2241 19617 2254
rect 18991 2167 19027 2185
rect 18958 2166 19027 2167
rect 18938 2154 19027 2166
rect 18938 2116 18950 2154
rect 18975 2119 18994 2154
rect 19019 2119 19027 2154
rect 18975 2116 19027 2119
rect 18938 2108 19027 2116
rect 18954 2107 19026 2108
rect 18507 1841 18623 1899
rect 19656 1888 19726 2409
rect 19808 2222 19842 2500
rect 20255 2480 20287 2508
rect 19875 2472 20287 2480
rect 19875 2446 19881 2472
rect 19907 2446 20287 2472
rect 19875 2444 20287 2446
rect 19877 2443 19917 2444
rect 20044 2418 20075 2426
rect 20044 2388 20048 2418
rect 20069 2388 20075 2418
rect 19808 2214 19843 2222
rect 19808 2194 19816 2214
rect 19836 2194 19843 2214
rect 19808 2189 19843 2194
rect 20044 2189 20075 2388
rect 20255 2379 20287 2444
rect 20255 2359 20259 2379
rect 20280 2359 20287 2379
rect 20255 2352 20287 2359
rect 20700 2505 20772 2523
rect 20700 2463 20713 2505
rect 20762 2463 20772 2505
rect 20700 2442 20772 2463
rect 20700 2400 20714 2442
rect 20763 2400 20772 2442
rect 20564 2296 20665 2297
rect 20462 2283 20665 2296
rect 20462 2281 20605 2283
rect 20462 2278 20539 2281
rect 20462 2251 20465 2278
rect 20494 2254 20539 2278
rect 20568 2254 20605 2281
rect 20494 2251 20605 2254
rect 20462 2250 20605 2251
rect 20641 2250 20665 2283
rect 20462 2237 20665 2250
rect 19808 2188 19840 2189
rect 20042 2186 20075 2189
rect 20008 2167 20076 2186
rect 19978 2155 20077 2167
rect 19978 2117 20000 2155
rect 20025 2120 20044 2155
rect 20069 2120 20077 2155
rect 20025 2117 20077 2120
rect 19978 2109 20077 2117
rect 20004 2108 20076 2109
rect 18507 1770 18519 1841
rect 18598 1770 18623 1841
rect 18507 1750 18623 1770
rect 19637 1687 19739 1888
rect 20700 1880 20772 2400
rect 21144 1976 21251 2588
rect 21963 3010 22070 3439
rect 22442 3198 22514 3439
rect 23137 3431 23236 3443
rect 23138 3412 23206 3431
rect 23139 3409 23172 3412
rect 23374 3409 23406 3410
rect 22549 3348 22752 3361
rect 22549 3315 22573 3348
rect 22609 3347 22752 3348
rect 22609 3344 22720 3347
rect 22609 3317 22646 3344
rect 22675 3320 22720 3344
rect 22749 3320 22752 3347
rect 22675 3317 22752 3320
rect 22609 3315 22752 3317
rect 22549 3302 22752 3315
rect 22549 3301 22650 3302
rect 22442 3156 22451 3198
rect 22500 3156 22514 3198
rect 22442 3135 22514 3156
rect 22442 3093 22452 3135
rect 22501 3093 22514 3135
rect 22442 3075 22514 3093
rect 22927 3239 22959 3246
rect 22927 3219 22934 3239
rect 22955 3219 22959 3239
rect 22927 3154 22959 3219
rect 23139 3210 23170 3409
rect 23371 3404 23406 3409
rect 23371 3384 23378 3404
rect 23398 3384 23406 3404
rect 23371 3376 23406 3384
rect 23139 3180 23145 3210
rect 23166 3180 23170 3210
rect 23139 3172 23170 3180
rect 23297 3154 23337 3155
rect 22927 3152 23339 3154
rect 22927 3126 23307 3152
rect 23333 3126 23339 3152
rect 22927 3118 23339 3126
rect 22927 3090 22959 3118
rect 23372 3098 23406 3376
rect 23488 3189 23558 3500
rect 24185 3491 25527 3496
rect 24185 3489 25484 3491
rect 24182 3463 25484 3489
rect 25512 3463 25527 3491
rect 24182 3455 25527 3463
rect 24182 3430 24221 3455
rect 24182 3413 24223 3430
rect 24182 3406 24221 3413
rect 23597 3344 23800 3357
rect 23597 3311 23621 3344
rect 23657 3343 23800 3344
rect 23657 3340 23768 3343
rect 23657 3313 23694 3340
rect 23723 3316 23768 3340
rect 23797 3316 23800 3343
rect 23723 3313 23800 3316
rect 23657 3311 23800 3313
rect 23597 3298 23800 3311
rect 23597 3297 23698 3298
rect 22927 3070 22932 3090
rect 22953 3070 22959 3090
rect 22927 3063 22959 3070
rect 23350 3093 23406 3098
rect 23350 3073 23357 3093
rect 23377 3073 23406 3093
rect 23483 3183 23558 3189
rect 23483 3150 23491 3183
rect 23544 3150 23558 3183
rect 23483 3125 23558 3150
rect 23483 3092 23496 3125
rect 23549 3092 23558 3125
rect 23483 3083 23558 3092
rect 23975 3235 24007 3242
rect 23975 3215 23982 3235
rect 24003 3215 24007 3235
rect 23975 3150 24007 3215
rect 24187 3206 24218 3406
rect 24422 3405 24454 3406
rect 24419 3400 24454 3405
rect 24419 3380 24426 3400
rect 24446 3380 24454 3400
rect 24419 3372 24454 3380
rect 24187 3176 24193 3206
rect 24214 3176 24218 3206
rect 24187 3168 24218 3176
rect 24345 3150 24385 3151
rect 23975 3148 24387 3150
rect 23975 3122 24355 3148
rect 24381 3122 24387 3148
rect 23975 3114 24387 3122
rect 23975 3086 24007 3114
rect 24420 3094 24454 3372
rect 23483 3078 23541 3083
rect 23350 3066 23406 3073
rect 23975 3066 23980 3086
rect 24001 3066 24007 3086
rect 23350 3065 23385 3066
rect 23975 3059 24007 3066
rect 24398 3089 24454 3094
rect 24398 3069 24405 3089
rect 24425 3069 24454 3089
rect 24398 3062 24454 3069
rect 24398 3061 24433 3062
rect 22641 3010 22752 3014
rect 24516 3010 25111 3011
rect 21963 2992 25111 3010
rect 21963 2972 22649 2992
rect 22668 2972 22726 2992
rect 22745 2988 25111 2992
rect 22745 2972 23697 2988
rect 21963 2968 23697 2972
rect 23716 2968 23774 2988
rect 23793 2968 25111 2988
rect 21963 2954 25111 2968
rect 21963 2331 22070 2954
rect 23689 2951 23800 2954
rect 22449 2905 22513 2909
rect 22445 2899 22513 2905
rect 22445 2866 22462 2899
rect 22502 2866 22513 2899
rect 22445 2854 22513 2866
rect 23496 2868 23561 2890
rect 22445 2852 22502 2854
rect 22449 2491 22500 2852
rect 23496 2829 23513 2868
rect 23558 2829 23561 2868
rect 23137 2784 23172 2786
rect 23137 2775 23241 2784
rect 23137 2774 23188 2775
rect 23137 2754 23140 2774
rect 23165 2755 23188 2774
rect 23220 2755 23241 2775
rect 23165 2754 23241 2755
rect 23137 2747 23241 2754
rect 23137 2735 23172 2747
rect 22549 2669 22752 2682
rect 22549 2636 22573 2669
rect 22609 2668 22752 2669
rect 22609 2665 22720 2668
rect 22609 2638 22646 2665
rect 22675 2641 22720 2665
rect 22749 2641 22752 2668
rect 22675 2638 22752 2641
rect 22609 2636 22752 2638
rect 22549 2623 22752 2636
rect 22549 2622 22650 2623
rect 22927 2560 22959 2567
rect 22927 2540 22934 2560
rect 22955 2540 22959 2560
rect 22438 2482 22503 2491
rect 22438 2445 22448 2482
rect 22488 2448 22503 2482
rect 22927 2475 22959 2540
rect 23139 2531 23170 2735
rect 23374 2730 23406 2731
rect 23371 2725 23406 2730
rect 23371 2705 23378 2725
rect 23398 2705 23406 2725
rect 23371 2697 23406 2705
rect 23139 2501 23145 2531
rect 23166 2501 23170 2531
rect 23139 2493 23170 2501
rect 23297 2475 23337 2476
rect 22927 2473 23339 2475
rect 22488 2445 22505 2448
rect 22438 2426 22505 2445
rect 22438 2405 22452 2426
rect 22488 2405 22505 2426
rect 22438 2398 22505 2405
rect 22927 2447 23307 2473
rect 23333 2447 23339 2473
rect 22927 2439 23339 2447
rect 22927 2411 22959 2439
rect 23372 2419 23406 2697
rect 23496 2566 23561 2829
rect 23496 2562 23557 2566
rect 22927 2391 22932 2411
rect 22953 2391 22959 2411
rect 22927 2384 22959 2391
rect 23350 2414 23406 2419
rect 23350 2394 23357 2414
rect 23377 2394 23406 2414
rect 23350 2387 23406 2394
rect 23350 2386 23385 2387
rect 22641 2331 22752 2335
rect 21961 2313 23280 2331
rect 21961 2293 22649 2313
rect 22668 2293 22726 2313
rect 22745 2293 23280 2313
rect 21961 2275 23280 2293
rect 21963 2155 22070 2275
rect 22431 2236 22552 2246
rect 22431 2234 22500 2236
rect 22431 2193 22444 2234
rect 22481 2195 22500 2234
rect 22537 2195 22552 2236
rect 22481 2193 22552 2195
rect 22431 2175 22552 2193
rect 21143 1940 21251 1976
rect 21298 2099 21452 2124
rect 21298 1987 21311 2099
rect 21432 1987 21452 2099
rect 19601 1650 19767 1687
rect 19601 1571 19638 1650
rect 19722 1571 19767 1650
rect 19601 1533 19767 1571
rect 20678 1479 20775 1880
rect 21136 1804 21256 1940
rect 21143 1798 21251 1804
rect 20608 1450 20783 1479
rect 20608 1371 20654 1450
rect 20754 1371 20783 1450
rect 20608 1346 20783 1371
rect 20955 1255 21018 1261
rect 21143 1255 21247 1798
rect 20955 1225 21257 1255
rect 20955 1138 21020 1225
rect 21090 1217 21257 1225
rect 21090 1138 21153 1217
rect 20955 1130 21153 1138
rect 21223 1130 21257 1217
rect 20955 1084 21257 1130
rect 16114 757 16166 797
rect 16116 710 16166 757
rect 11660 699 16166 710
rect 11660 651 11675 699
rect 11716 651 16166 699
rect 11660 646 16166 651
rect 11660 631 11725 646
rect 16116 644 16166 646
rect 10587 512 10790 525
rect 10587 479 10611 512
rect 10647 511 10790 512
rect 10647 508 10758 511
rect 10647 481 10684 508
rect 10713 484 10758 508
rect 10787 484 10790 511
rect 10713 481 10790 484
rect 10647 479 10790 481
rect 10587 466 10790 479
rect 10587 465 10688 466
rect 10965 403 10997 410
rect 10965 383 10972 403
rect 10993 383 10997 403
rect 10965 318 10997 383
rect 11177 374 11208 600
rect 11412 573 11444 574
rect 11409 568 11444 573
rect 11409 548 11416 568
rect 11436 548 11444 568
rect 11409 540 11444 548
rect 11177 344 11183 374
rect 11204 344 11208 374
rect 11177 336 11208 344
rect 11335 318 11375 319
rect 10965 316 11377 318
rect 10965 290 11345 316
rect 11371 290 11377 316
rect 10965 282 11377 290
rect 10965 254 10997 282
rect 11410 262 11444 540
rect 20148 572 20217 582
rect 20148 547 20162 572
rect 20203 547 20217 572
rect 20148 539 20217 547
rect 20150 432 20215 539
rect 10965 234 10970 254
rect 10991 234 10997 254
rect 10965 227 10997 234
rect 11176 255 11209 262
rect 11176 232 11184 255
rect 11204 232 11209 255
rect 10679 157 10790 178
rect 10383 156 10790 157
rect 10383 136 10687 156
rect 10706 136 10764 156
rect 10783 136 10790 156
rect 10383 119 10790 136
rect 11176 124 11209 232
rect 11388 257 11444 262
rect 11388 237 11395 257
rect 11415 237 11444 257
rect 11388 230 11444 237
rect 20145 403 20215 432
rect 11388 229 11423 230
rect 20145 124 20213 403
rect 20470 337 20571 352
rect 20470 319 20816 337
rect 20470 266 20556 319
rect 20753 266 20816 319
rect 20470 246 20816 266
rect 10383 85 10784 119
rect 11176 59 20220 124
rect 11176 56 11209 59
rect 20470 13 20571 246
rect 20955 154 21054 1084
rect 21298 1013 21452 1987
rect 21762 2082 21896 2111
rect 21762 1970 21800 2082
rect 21879 1970 21896 2082
rect 21963 2075 22071 2155
rect 21762 1017 21896 1970
rect 21964 1263 22071 2075
rect 22437 2103 22502 2175
rect 22437 2037 22505 2103
rect 22438 1491 22505 2037
rect 23492 1675 23557 2562
rect 24535 2292 24672 2296
rect 24522 2288 24679 2292
rect 24522 2181 24559 2288
rect 24659 2181 24679 2288
rect 24522 2139 24679 2181
rect 24535 1891 24672 2139
rect 24525 1849 24691 1891
rect 24525 1774 24554 1849
rect 24671 1774 24691 1849
rect 24525 1758 24691 1774
rect 23481 1654 23618 1675
rect 23481 1579 23506 1654
rect 23576 1579 23618 1654
rect 23481 1548 23618 1579
rect 22424 1442 22599 1491
rect 22424 1363 22457 1442
rect 22557 1363 22599 1442
rect 22424 1358 22599 1363
rect 21964 1221 22112 1263
rect 21964 1213 22004 1221
rect 21966 1134 22004 1213
rect 22074 1134 22112 1221
rect 21966 1096 22112 1134
rect 21296 997 21452 1013
rect 21296 972 21448 997
rect 21296 877 21326 972
rect 21416 877 21448 972
rect 21296 864 21448 877
rect 21758 981 21897 1017
rect 21758 886 21772 981
rect 21862 886 21897 981
rect 21758 868 21897 886
rect 27079 791 27127 4521
rect 27300 4542 27356 4547
rect 27300 4522 27307 4542
rect 27327 4522 27356 4542
rect 27300 4515 27356 4522
rect 27300 4514 27335 4515
rect 27404 4424 27432 7232
rect 30617 7187 30682 7487
rect 30772 7319 30806 7597
rect 31219 7577 31251 7605
rect 30839 7569 31251 7577
rect 30839 7543 30845 7569
rect 30871 7543 31251 7569
rect 31673 7611 31740 7618
rect 31673 7590 31690 7611
rect 31726 7590 31740 7611
rect 31673 7571 31740 7590
rect 31673 7568 31690 7571
rect 30839 7541 31251 7543
rect 30841 7540 30881 7541
rect 31008 7515 31039 7523
rect 31008 7485 31012 7515
rect 31033 7485 31039 7515
rect 30772 7311 30807 7319
rect 30772 7291 30780 7311
rect 30800 7291 30807 7311
rect 30772 7286 30807 7291
rect 30772 7285 30804 7286
rect 31008 7281 31039 7485
rect 31219 7476 31251 7541
rect 31675 7534 31690 7568
rect 31730 7534 31740 7571
rect 31675 7525 31740 7534
rect 31219 7456 31223 7476
rect 31244 7456 31251 7476
rect 31219 7449 31251 7456
rect 31528 7393 31629 7394
rect 31426 7380 31629 7393
rect 31426 7378 31569 7380
rect 31426 7375 31503 7378
rect 31426 7348 31429 7375
rect 31458 7351 31503 7375
rect 31532 7351 31569 7378
rect 31458 7348 31569 7351
rect 31426 7347 31569 7348
rect 31605 7347 31629 7380
rect 31426 7334 31629 7347
rect 31006 7269 31041 7281
rect 30937 7262 31041 7269
rect 30937 7261 31013 7262
rect 30937 7241 30958 7261
rect 30990 7242 31013 7261
rect 31038 7242 31041 7262
rect 30990 7241 31041 7242
rect 30937 7232 31041 7241
rect 31006 7230 31041 7232
rect 30617 7148 30620 7187
rect 30665 7148 30682 7187
rect 31678 7164 31729 7525
rect 31676 7162 31733 7164
rect 30617 7126 30682 7148
rect 31665 7150 31733 7162
rect 31665 7117 31676 7150
rect 31716 7117 31733 7150
rect 31665 7111 31733 7117
rect 31665 7107 31729 7111
rect 30378 7062 30489 7065
rect 32108 7062 32215 7685
rect 28672 7048 32215 7062
rect 28672 7028 30385 7048
rect 30404 7028 30462 7048
rect 30481 7044 32215 7048
rect 30481 7028 31433 7044
rect 28672 7024 31433 7028
rect 31452 7024 31510 7044
rect 31529 7024 32215 7044
rect 28672 7006 32215 7024
rect 28672 7005 29662 7006
rect 31426 7002 31537 7006
rect 29745 6954 29780 6955
rect 29724 6947 29780 6954
rect 29724 6927 29753 6947
rect 29773 6927 29780 6947
rect 29724 6922 29780 6927
rect 30171 6950 30203 6957
rect 30793 6950 30828 6951
rect 30171 6930 30177 6950
rect 30198 6930 30203 6950
rect 30772 6943 30828 6950
rect 30637 6933 30695 6938
rect 29724 6644 29758 6922
rect 30171 6902 30203 6930
rect 29791 6894 30203 6902
rect 29791 6868 29797 6894
rect 29823 6868 30203 6894
rect 29791 6866 30203 6868
rect 29793 6865 29833 6866
rect 29960 6840 29991 6848
rect 29960 6810 29964 6840
rect 29985 6810 29991 6840
rect 29724 6636 29759 6644
rect 29724 6616 29732 6636
rect 29752 6616 29759 6636
rect 29724 6611 29759 6616
rect 29724 6610 29756 6611
rect 29960 6610 29991 6810
rect 30171 6801 30203 6866
rect 30171 6781 30175 6801
rect 30196 6781 30203 6801
rect 30171 6774 30203 6781
rect 30620 6924 30695 6933
rect 30620 6891 30629 6924
rect 30682 6891 30695 6924
rect 30620 6866 30695 6891
rect 30620 6833 30634 6866
rect 30687 6833 30695 6866
rect 30620 6827 30695 6833
rect 30772 6923 30801 6943
rect 30821 6923 30828 6943
rect 30772 6918 30828 6923
rect 31219 6946 31251 6953
rect 31219 6926 31225 6946
rect 31246 6926 31251 6946
rect 30480 6718 30581 6719
rect 30378 6705 30581 6718
rect 30378 6703 30521 6705
rect 30378 6700 30455 6703
rect 30378 6673 30381 6700
rect 30410 6676 30455 6700
rect 30484 6676 30521 6703
rect 30410 6673 30521 6676
rect 30378 6672 30521 6673
rect 30557 6672 30581 6705
rect 30378 6659 30581 6672
rect 29957 6603 29996 6610
rect 29955 6586 29996 6603
rect 29957 6561 29996 6586
rect 28651 6553 29996 6561
rect 28651 6525 28666 6553
rect 28694 6527 29996 6553
rect 28694 6525 29993 6527
rect 28651 6520 29993 6525
rect 30620 6516 30690 6827
rect 30772 6640 30806 6918
rect 31219 6898 31251 6926
rect 30839 6890 31251 6898
rect 30839 6864 30845 6890
rect 30871 6864 31251 6890
rect 30839 6862 31251 6864
rect 30841 6861 30881 6862
rect 31008 6836 31039 6844
rect 31008 6806 31012 6836
rect 31033 6806 31039 6836
rect 30772 6632 30807 6640
rect 30772 6612 30780 6632
rect 30800 6612 30807 6632
rect 30772 6607 30807 6612
rect 31008 6607 31039 6806
rect 31219 6797 31251 6862
rect 31219 6777 31223 6797
rect 31244 6777 31251 6797
rect 31219 6770 31251 6777
rect 31664 6923 31736 6941
rect 31664 6881 31677 6923
rect 31726 6881 31736 6923
rect 31664 6860 31736 6881
rect 31664 6818 31678 6860
rect 31727 6818 31736 6860
rect 31528 6714 31629 6715
rect 31426 6701 31629 6714
rect 31426 6699 31569 6701
rect 31426 6696 31503 6699
rect 31426 6669 31429 6696
rect 31458 6672 31503 6696
rect 31532 6672 31569 6699
rect 31458 6669 31569 6672
rect 31426 6668 31569 6669
rect 31605 6668 31629 6701
rect 31426 6655 31629 6668
rect 30772 6606 30804 6607
rect 31006 6604 31039 6607
rect 30972 6585 31040 6604
rect 30942 6573 31041 6585
rect 31664 6577 31736 6818
rect 32108 6577 32215 7006
rect 32670 7418 32777 7878
rect 33149 7606 33221 7900
rect 33845 7897 33917 7898
rect 33844 7889 33943 7897
rect 34197 7892 34274 8075
rect 35485 8076 35569 8087
rect 35485 8048 35513 8076
rect 35557 8048 35569 8076
rect 35299 7997 35373 8025
rect 35299 7949 35322 7997
rect 35359 7949 35373 7997
rect 35485 8019 35569 8048
rect 35485 7991 35510 8019
rect 35554 7991 35569 8019
rect 35485 7958 35569 7991
rect 35299 7940 35373 7949
rect 34895 7898 34967 7899
rect 33844 7886 33896 7889
rect 33844 7851 33852 7886
rect 33877 7851 33896 7886
rect 33921 7851 33943 7889
rect 33844 7839 33943 7851
rect 34195 7863 34274 7892
rect 34894 7890 34983 7898
rect 34894 7887 34946 7890
rect 33845 7820 33913 7839
rect 33846 7817 33879 7820
rect 34081 7817 34113 7818
rect 33256 7756 33459 7769
rect 33256 7723 33280 7756
rect 33316 7755 33459 7756
rect 33316 7752 33427 7755
rect 33316 7725 33353 7752
rect 33382 7728 33427 7752
rect 33456 7728 33459 7755
rect 33382 7725 33459 7728
rect 33316 7723 33459 7725
rect 33256 7710 33459 7723
rect 33256 7709 33357 7710
rect 33149 7564 33158 7606
rect 33207 7564 33221 7606
rect 33149 7543 33221 7564
rect 33149 7501 33159 7543
rect 33208 7501 33221 7543
rect 33149 7483 33221 7501
rect 33634 7647 33666 7654
rect 33634 7627 33641 7647
rect 33662 7627 33666 7647
rect 33634 7562 33666 7627
rect 33846 7618 33877 7817
rect 34078 7812 34113 7817
rect 34078 7792 34085 7812
rect 34105 7792 34113 7812
rect 34078 7784 34113 7792
rect 33846 7588 33852 7618
rect 33873 7588 33877 7618
rect 33846 7580 33877 7588
rect 34004 7562 34044 7563
rect 33634 7560 34046 7562
rect 33634 7534 34014 7560
rect 34040 7534 34046 7560
rect 33634 7526 34046 7534
rect 33634 7498 33666 7526
rect 34079 7506 34113 7784
rect 34195 7597 34265 7863
rect 34894 7852 34902 7887
rect 34927 7852 34946 7887
rect 34971 7852 34983 7890
rect 34894 7840 34983 7852
rect 34894 7839 34963 7840
rect 34894 7821 34930 7839
rect 34304 7752 34507 7765
rect 34304 7719 34328 7752
rect 34364 7751 34507 7752
rect 34364 7748 34475 7751
rect 34364 7721 34401 7748
rect 34430 7724 34475 7748
rect 34504 7724 34507 7751
rect 34430 7721 34507 7724
rect 34364 7719 34507 7721
rect 34304 7706 34507 7719
rect 34304 7705 34405 7706
rect 33634 7478 33639 7498
rect 33660 7478 33666 7498
rect 33634 7471 33666 7478
rect 34057 7501 34113 7506
rect 34057 7481 34064 7501
rect 34084 7481 34113 7501
rect 34190 7591 34265 7597
rect 34190 7558 34198 7591
rect 34251 7558 34265 7591
rect 34190 7533 34265 7558
rect 34190 7500 34203 7533
rect 34256 7500 34265 7533
rect 34190 7491 34265 7500
rect 34682 7643 34714 7650
rect 34682 7623 34689 7643
rect 34710 7623 34714 7643
rect 34682 7558 34714 7623
rect 34894 7614 34925 7821
rect 35129 7813 35161 7814
rect 35126 7808 35161 7813
rect 35126 7788 35133 7808
rect 35153 7788 35161 7808
rect 35126 7780 35161 7788
rect 34894 7584 34900 7614
rect 34921 7584 34925 7614
rect 34894 7576 34925 7584
rect 35052 7558 35092 7559
rect 34682 7556 35094 7558
rect 34682 7530 35062 7556
rect 35088 7530 35094 7556
rect 34682 7522 35094 7530
rect 34682 7494 34714 7522
rect 35127 7502 35161 7780
rect 35310 7595 35372 7940
rect 35479 7913 35569 7958
rect 35479 7598 35561 7913
rect 35310 7576 35374 7595
rect 35310 7537 35323 7576
rect 35357 7537 35374 7576
rect 35310 7518 35374 7537
rect 35479 7557 35500 7598
rect 35536 7557 35561 7598
rect 35479 7528 35561 7557
rect 34190 7486 34248 7491
rect 34057 7474 34113 7481
rect 34682 7474 34687 7494
rect 34708 7474 34714 7494
rect 34057 7473 34092 7474
rect 34682 7467 34714 7474
rect 35105 7497 35161 7502
rect 35105 7477 35112 7497
rect 35132 7477 35161 7497
rect 35105 7470 35161 7477
rect 35105 7469 35140 7470
rect 33348 7418 33459 7422
rect 35131 7418 36701 7419
rect 32670 7400 36701 7418
rect 32670 7380 33356 7400
rect 33375 7380 33433 7400
rect 33452 7396 36701 7400
rect 33452 7380 34404 7396
rect 32670 7376 34404 7380
rect 34423 7376 34481 7396
rect 34500 7376 36701 7396
rect 32670 7362 36701 7376
rect 32670 6739 32777 7362
rect 34396 7359 34507 7362
rect 33156 7313 33220 7317
rect 33152 7307 33220 7313
rect 33152 7274 33169 7307
rect 33209 7274 33220 7307
rect 33152 7262 33220 7274
rect 34203 7276 34268 7298
rect 33152 7260 33209 7262
rect 33156 6899 33207 7260
rect 34203 7237 34220 7276
rect 34265 7237 34268 7276
rect 33844 7192 33879 7194
rect 33844 7183 33948 7192
rect 33844 7182 33895 7183
rect 33844 7162 33847 7182
rect 33872 7163 33895 7182
rect 33927 7163 33948 7183
rect 33872 7162 33948 7163
rect 33844 7155 33948 7162
rect 33844 7143 33879 7155
rect 33256 7077 33459 7090
rect 33256 7044 33280 7077
rect 33316 7076 33459 7077
rect 33316 7073 33427 7076
rect 33316 7046 33353 7073
rect 33382 7049 33427 7073
rect 33456 7049 33459 7076
rect 33382 7046 33459 7049
rect 33316 7044 33459 7046
rect 33256 7031 33459 7044
rect 33256 7030 33357 7031
rect 33634 6968 33666 6975
rect 33634 6948 33641 6968
rect 33662 6948 33666 6968
rect 33145 6890 33210 6899
rect 33145 6853 33155 6890
rect 33195 6856 33210 6890
rect 33634 6883 33666 6948
rect 33846 6939 33877 7143
rect 34081 7138 34113 7139
rect 34078 7133 34113 7138
rect 34078 7113 34085 7133
rect 34105 7113 34113 7133
rect 34078 7105 34113 7113
rect 33846 6909 33852 6939
rect 33873 6909 33877 6939
rect 33846 6901 33877 6909
rect 34004 6883 34044 6884
rect 33634 6881 34046 6883
rect 33195 6853 33212 6856
rect 33145 6834 33212 6853
rect 33145 6813 33159 6834
rect 33195 6813 33212 6834
rect 33145 6806 33212 6813
rect 33634 6855 34014 6881
rect 34040 6855 34046 6881
rect 33634 6847 34046 6855
rect 33634 6819 33666 6847
rect 34079 6827 34113 7105
rect 34203 6937 34268 7237
rect 35474 7261 35567 7276
rect 35474 7217 35489 7261
rect 35549 7217 35567 7261
rect 33634 6799 33639 6819
rect 33660 6799 33666 6819
rect 33634 6792 33666 6799
rect 34057 6822 34113 6827
rect 34057 6802 34064 6822
rect 34084 6802 34113 6822
rect 34057 6795 34113 6802
rect 34193 6926 34273 6937
rect 34193 6900 34210 6926
rect 34250 6900 34273 6926
rect 34193 6873 34273 6900
rect 34193 6847 34214 6873
rect 34254 6847 34273 6873
rect 34193 6828 34273 6847
rect 34193 6802 34217 6828
rect 34257 6802 34273 6828
rect 34057 6794 34092 6795
rect 34193 6790 34273 6802
rect 35474 6844 35567 7217
rect 35751 7072 35954 7085
rect 35751 7039 35775 7072
rect 35811 7071 35954 7072
rect 35811 7068 35922 7071
rect 35811 7041 35848 7068
rect 35877 7044 35922 7068
rect 35951 7044 35954 7071
rect 35877 7041 35954 7044
rect 35811 7039 35954 7041
rect 35751 7026 35954 7039
rect 35751 7025 35852 7026
rect 35474 6803 35489 6844
rect 35543 6803 35567 6844
rect 35474 6796 35567 6803
rect 36129 6963 36161 6970
rect 36129 6943 36136 6963
rect 36157 6943 36161 6963
rect 36129 6878 36161 6943
rect 36341 6934 36372 7135
rect 36576 7133 36608 7134
rect 36573 7128 36608 7133
rect 36573 7108 36580 7128
rect 36600 7108 36608 7128
rect 36573 7100 36608 7108
rect 36341 6904 36347 6934
rect 36368 6904 36372 6934
rect 36341 6896 36372 6904
rect 36499 6878 36539 6879
rect 36129 6876 36541 6878
rect 36129 6850 36509 6876
rect 36535 6850 36541 6876
rect 36129 6842 36541 6850
rect 36129 6814 36161 6842
rect 36574 6822 36608 7100
rect 36129 6794 36134 6814
rect 36155 6794 36161 6814
rect 36129 6787 36161 6794
rect 36552 6817 36608 6822
rect 36552 6797 36559 6817
rect 36579 6797 36608 6817
rect 36552 6790 36608 6797
rect 36552 6789 36587 6790
rect 33348 6739 33459 6743
rect 35090 6739 36734 6742
rect 32668 6721 36734 6739
rect 32668 6701 33356 6721
rect 33375 6701 33433 6721
rect 33452 6716 36734 6721
rect 33452 6701 35851 6716
rect 32668 6696 35851 6701
rect 35870 6696 35928 6716
rect 35947 6696 36734 6716
rect 32668 6686 36734 6696
rect 32668 6683 33293 6686
rect 33480 6683 36734 6686
rect 30942 6535 30964 6573
rect 30989 6538 31008 6573
rect 31033 6538 31041 6573
rect 30989 6535 31041 6538
rect 30942 6527 31041 6535
rect 30968 6526 31040 6527
rect 30619 6500 30690 6516
rect 30619 6484 30639 6500
rect 30620 6454 30639 6484
rect 30622 6434 30639 6454
rect 30669 6454 30690 6500
rect 31662 6496 31740 6577
rect 32107 6522 32215 6577
rect 30669 6434 30689 6454
rect 30622 6415 30689 6434
rect 31662 6394 31741 6496
rect 31626 6376 31747 6394
rect 31626 6374 31697 6376
rect 31626 6333 31641 6374
rect 31678 6335 31697 6374
rect 31734 6335 31747 6376
rect 31678 6333 31747 6335
rect 31626 6323 31747 6333
rect 28931 6295 29042 6298
rect 28245 6294 29795 6295
rect 32108 6294 32215 6522
rect 32670 6455 32777 6683
rect 35090 6682 36734 6683
rect 35843 6679 35954 6682
rect 33138 6644 33259 6654
rect 33138 6642 33207 6644
rect 33138 6601 33151 6642
rect 33188 6603 33207 6642
rect 33244 6603 33259 6644
rect 33188 6601 33259 6603
rect 33138 6583 33259 6601
rect 36343 6624 36429 6628
rect 36343 6606 36358 6624
rect 36410 6606 36429 6624
rect 36343 6597 36429 6606
rect 33144 6481 33223 6583
rect 34196 6543 34263 6562
rect 34196 6523 34216 6543
rect 32670 6400 32778 6455
rect 33145 6400 33223 6481
rect 34195 6477 34216 6523
rect 34246 6523 34263 6543
rect 34246 6493 34265 6523
rect 34246 6477 34266 6493
rect 34195 6461 34266 6477
rect 33845 6450 33917 6451
rect 33844 6442 33943 6450
rect 33844 6439 33896 6442
rect 33844 6404 33852 6439
rect 33877 6404 33896 6439
rect 33921 6404 33943 6442
rect 28245 6291 31405 6294
rect 31592 6291 32217 6294
rect 28245 6281 32217 6291
rect 28245 6261 28938 6281
rect 28957 6261 29015 6281
rect 29034 6276 32217 6281
rect 29034 6261 31433 6276
rect 28245 6256 31433 6261
rect 31452 6256 31510 6276
rect 31529 6256 32217 6276
rect 28245 6238 32217 6256
rect 28245 6235 29795 6238
rect 31426 6234 31537 6238
rect 28298 6187 28333 6188
rect 28277 6180 28333 6187
rect 28277 6160 28306 6180
rect 28326 6160 28333 6180
rect 28277 6155 28333 6160
rect 28724 6183 28756 6190
rect 28724 6163 28730 6183
rect 28751 6163 28756 6183
rect 28277 5877 28311 6155
rect 28724 6135 28756 6163
rect 30612 6175 30692 6187
rect 30793 6182 30828 6183
rect 28344 6127 28756 6135
rect 28344 6101 28350 6127
rect 28376 6101 28756 6127
rect 29142 6141 29579 6154
rect 29142 6118 29155 6141
rect 29181 6134 29579 6141
rect 29181 6118 29535 6134
rect 29142 6111 29535 6118
rect 29561 6111 29579 6134
rect 29142 6105 29579 6111
rect 30612 6149 30628 6175
rect 30668 6149 30692 6175
rect 30612 6130 30692 6149
rect 28344 6099 28756 6101
rect 28346 6098 28386 6099
rect 28513 6073 28544 6081
rect 28513 6043 28517 6073
rect 28538 6043 28544 6073
rect 28277 5869 28312 5877
rect 28277 5849 28285 5869
rect 28305 5849 28312 5869
rect 28277 5844 28312 5849
rect 28277 5843 28309 5844
rect 28513 5836 28544 6043
rect 28724 6034 28756 6099
rect 30612 6104 30631 6130
rect 30671 6104 30692 6130
rect 30612 6077 30692 6104
rect 30612 6051 30635 6077
rect 30675 6051 30692 6077
rect 30612 6040 30692 6051
rect 30772 6175 30828 6182
rect 30772 6155 30801 6175
rect 30821 6155 30828 6175
rect 30772 6150 30828 6155
rect 31219 6178 31251 6185
rect 31219 6158 31225 6178
rect 31246 6158 31251 6178
rect 28724 6014 28728 6034
rect 28749 6014 28756 6034
rect 28724 6007 28756 6014
rect 29033 5951 29134 5952
rect 28931 5938 29134 5951
rect 28931 5936 29074 5938
rect 28931 5933 29008 5936
rect 28931 5906 28934 5933
rect 28963 5909 29008 5933
rect 29037 5909 29074 5936
rect 28963 5906 29074 5909
rect 28931 5905 29074 5906
rect 29110 5905 29134 5938
rect 28931 5892 29134 5905
rect 28511 5830 28544 5836
rect 28507 5826 28544 5830
rect 28507 5816 28545 5826
rect 28507 5803 28517 5816
rect 28508 5779 28517 5803
rect 28534 5779 28545 5816
rect 28508 5758 28545 5779
rect 30617 5740 30682 6040
rect 30772 5872 30806 6150
rect 31219 6130 31251 6158
rect 30839 6122 31251 6130
rect 30839 6096 30845 6122
rect 30871 6096 31251 6122
rect 31673 6164 31740 6171
rect 31673 6143 31690 6164
rect 31726 6143 31740 6164
rect 31673 6124 31740 6143
rect 31673 6121 31690 6124
rect 30839 6094 31251 6096
rect 30841 6093 30881 6094
rect 31008 6068 31039 6076
rect 31008 6038 31012 6068
rect 31033 6038 31039 6068
rect 30772 5864 30807 5872
rect 30772 5844 30780 5864
rect 30800 5844 30807 5864
rect 30772 5839 30807 5844
rect 30772 5838 30804 5839
rect 31008 5834 31039 6038
rect 31219 6029 31251 6094
rect 31675 6087 31690 6121
rect 31730 6087 31740 6124
rect 31675 6078 31740 6087
rect 31219 6009 31223 6029
rect 31244 6009 31251 6029
rect 31219 6002 31251 6009
rect 31528 5946 31629 5947
rect 31426 5933 31629 5946
rect 31426 5931 31569 5933
rect 31426 5928 31503 5931
rect 31426 5901 31429 5928
rect 31458 5904 31503 5928
rect 31532 5904 31569 5931
rect 31458 5901 31569 5904
rect 31426 5900 31569 5901
rect 31605 5900 31629 5933
rect 31426 5887 31629 5900
rect 31006 5822 31041 5834
rect 30937 5815 31041 5822
rect 30937 5814 31013 5815
rect 30937 5794 30958 5814
rect 30990 5795 31013 5814
rect 31038 5795 31041 5815
rect 30990 5794 31041 5795
rect 30937 5785 31041 5794
rect 31006 5783 31041 5785
rect 30617 5701 30620 5740
rect 30665 5701 30682 5740
rect 31678 5717 31729 6078
rect 31676 5715 31733 5717
rect 30617 5679 30682 5701
rect 31665 5703 31733 5715
rect 31665 5670 31676 5703
rect 31716 5670 31733 5703
rect 31665 5664 31733 5670
rect 31665 5660 31729 5664
rect 30378 5615 30489 5618
rect 32108 5615 32215 6238
rect 28454 5601 32215 5615
rect 28454 5581 30385 5601
rect 30404 5581 30462 5601
rect 30481 5597 32215 5601
rect 30481 5581 31433 5597
rect 28454 5577 31433 5581
rect 31452 5577 31510 5597
rect 31529 5577 32215 5597
rect 28454 5559 32215 5577
rect 28454 5558 29754 5559
rect 31426 5555 31537 5559
rect 29745 5507 29780 5508
rect 29724 5500 29780 5507
rect 29724 5480 29753 5500
rect 29773 5480 29780 5500
rect 29724 5475 29780 5480
rect 30171 5503 30203 5510
rect 30793 5503 30828 5504
rect 30171 5483 30177 5503
rect 30198 5483 30203 5503
rect 30772 5496 30828 5503
rect 30637 5486 30695 5491
rect 29724 5197 29758 5475
rect 30171 5455 30203 5483
rect 29791 5447 30203 5455
rect 29791 5421 29797 5447
rect 29823 5421 30203 5447
rect 29791 5419 30203 5421
rect 29793 5418 29833 5419
rect 29960 5393 29991 5401
rect 29960 5363 29964 5393
rect 29985 5363 29991 5393
rect 29724 5189 29759 5197
rect 29724 5169 29732 5189
rect 29752 5169 29759 5189
rect 29724 5164 29759 5169
rect 29724 5163 29756 5164
rect 29960 5156 29991 5363
rect 30171 5354 30203 5419
rect 30171 5334 30175 5354
rect 30196 5334 30203 5354
rect 30171 5327 30203 5334
rect 30620 5477 30695 5486
rect 30620 5444 30629 5477
rect 30682 5444 30695 5477
rect 30620 5419 30695 5444
rect 30620 5386 30634 5419
rect 30687 5386 30695 5419
rect 30620 5380 30695 5386
rect 30772 5476 30801 5496
rect 30821 5476 30828 5496
rect 30772 5471 30828 5476
rect 31219 5499 31251 5506
rect 31219 5479 31225 5499
rect 31246 5479 31251 5499
rect 30480 5271 30581 5272
rect 30378 5258 30581 5271
rect 30378 5256 30521 5258
rect 30378 5253 30455 5256
rect 30378 5226 30381 5253
rect 30410 5229 30455 5253
rect 30484 5229 30521 5256
rect 30410 5226 30521 5229
rect 30378 5225 30521 5226
rect 30557 5225 30581 5258
rect 30378 5212 30581 5225
rect 29458 5143 29622 5146
rect 29955 5143 29991 5156
rect 28657 5125 29996 5143
rect 28657 5087 28667 5125
rect 28692 5110 29996 5125
rect 28692 5087 28702 5110
rect 29458 5103 29622 5110
rect 28657 5079 28702 5087
rect 28671 5078 28702 5079
rect 30620 5064 30690 5380
rect 30772 5193 30806 5471
rect 31219 5451 31251 5479
rect 30839 5443 31251 5451
rect 30839 5417 30845 5443
rect 30871 5417 31251 5443
rect 30839 5415 31251 5417
rect 30841 5414 30881 5415
rect 31008 5389 31039 5397
rect 31008 5359 31012 5389
rect 31033 5359 31039 5389
rect 30772 5185 30807 5193
rect 30772 5165 30780 5185
rect 30800 5165 30807 5185
rect 30772 5160 30807 5165
rect 31008 5160 31039 5359
rect 31219 5350 31251 5415
rect 31219 5330 31223 5350
rect 31244 5330 31251 5350
rect 31219 5323 31251 5330
rect 31664 5476 31736 5494
rect 31664 5434 31677 5476
rect 31726 5434 31736 5476
rect 31664 5413 31736 5434
rect 31664 5371 31678 5413
rect 31727 5371 31736 5413
rect 31528 5267 31629 5268
rect 31426 5254 31629 5267
rect 31426 5252 31569 5254
rect 31426 5249 31503 5252
rect 31426 5222 31429 5249
rect 31458 5225 31503 5249
rect 31532 5225 31569 5252
rect 31458 5222 31569 5225
rect 31426 5221 31569 5222
rect 31605 5221 31629 5254
rect 31426 5208 31629 5221
rect 30772 5159 30804 5160
rect 31006 5157 31039 5160
rect 30972 5138 31040 5157
rect 30942 5126 31041 5138
rect 30942 5088 30964 5126
rect 30989 5091 31008 5126
rect 31033 5091 31041 5126
rect 30989 5088 31041 5091
rect 30942 5080 31041 5088
rect 30968 5079 31040 5080
rect 30620 5045 30699 5064
rect 30623 5025 30699 5045
rect 30616 5001 30699 5025
rect 31664 5060 31736 5371
rect 31664 5017 31740 5060
rect 30616 4935 30628 5001
rect 30682 4935 30699 5001
rect 30616 4915 30699 4935
rect 30616 4878 30633 4915
rect 30677 4901 30699 4915
rect 31665 4966 31740 5017
rect 32108 4966 32215 5559
rect 32670 5971 32777 6400
rect 33149 6159 33221 6400
rect 33844 6392 33943 6404
rect 33845 6373 33913 6392
rect 33846 6370 33879 6373
rect 34081 6370 34113 6371
rect 33256 6309 33459 6322
rect 33256 6276 33280 6309
rect 33316 6308 33459 6309
rect 33316 6305 33427 6308
rect 33316 6278 33353 6305
rect 33382 6281 33427 6305
rect 33456 6281 33459 6308
rect 33382 6278 33459 6281
rect 33316 6276 33459 6278
rect 33256 6263 33459 6276
rect 33256 6262 33357 6263
rect 33149 6117 33158 6159
rect 33207 6117 33221 6159
rect 33149 6096 33221 6117
rect 33149 6054 33159 6096
rect 33208 6054 33221 6096
rect 33149 6036 33221 6054
rect 33634 6200 33666 6207
rect 33634 6180 33641 6200
rect 33662 6180 33666 6200
rect 33634 6115 33666 6180
rect 33846 6171 33877 6370
rect 34078 6365 34113 6370
rect 34078 6345 34085 6365
rect 34105 6345 34113 6365
rect 34078 6337 34113 6345
rect 33846 6141 33852 6171
rect 33873 6141 33877 6171
rect 33846 6133 33877 6141
rect 34004 6115 34044 6116
rect 33634 6113 34046 6115
rect 33634 6087 34014 6113
rect 34040 6087 34046 6113
rect 33634 6079 34046 6087
rect 33634 6051 33666 6079
rect 34079 6059 34113 6337
rect 34195 6150 34265 6461
rect 36120 6451 36192 6452
rect 36119 6448 36208 6451
rect 34891 6446 36208 6448
rect 34888 6443 36208 6446
rect 34888 6440 36171 6443
rect 34888 6405 36127 6440
rect 36152 6405 36171 6440
rect 36196 6405 36208 6443
rect 34888 6395 36208 6405
rect 36384 6444 36420 6597
rect 36384 6421 36390 6444
rect 36414 6421 36420 6444
rect 36384 6400 36420 6421
rect 34888 6393 36173 6395
rect 34888 6383 34985 6393
rect 34894 6374 34930 6383
rect 36384 6377 36390 6400
rect 36414 6377 36420 6400
rect 34304 6305 34507 6318
rect 34304 6272 34328 6305
rect 34364 6304 34507 6305
rect 34364 6301 34475 6304
rect 34364 6274 34401 6301
rect 34430 6277 34475 6301
rect 34504 6277 34507 6304
rect 34430 6274 34507 6277
rect 34364 6272 34507 6274
rect 34304 6259 34507 6272
rect 34304 6258 34405 6259
rect 33634 6031 33639 6051
rect 33660 6031 33666 6051
rect 33634 6024 33666 6031
rect 34057 6054 34113 6059
rect 34057 6034 34064 6054
rect 34084 6034 34113 6054
rect 34190 6144 34265 6150
rect 34190 6111 34198 6144
rect 34251 6111 34265 6144
rect 34190 6086 34265 6111
rect 34190 6053 34203 6086
rect 34256 6053 34265 6086
rect 34190 6044 34265 6053
rect 34682 6196 34714 6203
rect 34682 6176 34689 6196
rect 34710 6176 34714 6196
rect 34682 6111 34714 6176
rect 34894 6167 34925 6374
rect 35129 6366 35161 6367
rect 36384 6366 36420 6377
rect 35126 6361 35161 6366
rect 35126 6341 35133 6361
rect 35153 6341 35161 6361
rect 35126 6333 35161 6341
rect 34894 6137 34900 6167
rect 34921 6137 34925 6167
rect 34894 6129 34925 6137
rect 35052 6111 35092 6112
rect 34682 6109 35094 6111
rect 34682 6083 35062 6109
rect 35088 6083 35094 6109
rect 34682 6075 35094 6083
rect 34682 6047 34714 6075
rect 35127 6055 35161 6333
rect 34190 6039 34248 6044
rect 34057 6027 34113 6034
rect 34682 6027 34687 6047
rect 34708 6027 34714 6047
rect 34057 6026 34092 6027
rect 34682 6020 34714 6027
rect 35105 6050 35161 6055
rect 35105 6030 35112 6050
rect 35132 6030 35161 6050
rect 35105 6023 35161 6030
rect 35105 6022 35140 6023
rect 33348 5971 33459 5975
rect 35223 5971 36382 5972
rect 32670 5953 36382 5971
rect 32670 5933 33356 5953
rect 33375 5933 33433 5953
rect 33452 5949 36382 5953
rect 33452 5933 34404 5949
rect 32670 5929 34404 5933
rect 34423 5929 34481 5949
rect 34500 5929 36382 5949
rect 32670 5915 36382 5929
rect 32670 5292 32777 5915
rect 34396 5912 34507 5915
rect 33156 5866 33220 5870
rect 33152 5860 33220 5866
rect 33152 5827 33169 5860
rect 33209 5827 33220 5860
rect 33152 5815 33220 5827
rect 34203 5829 34268 5851
rect 33152 5813 33209 5815
rect 33156 5452 33207 5813
rect 34203 5790 34220 5829
rect 34265 5790 34268 5829
rect 37289 5827 37341 8133
rect 37450 8110 37485 8176
rect 37450 6794 37484 8110
rect 37788 7963 37893 13063
rect 40271 13050 42925 13064
rect 40271 13030 41095 13050
rect 41114 13030 41172 13050
rect 41191 13046 42925 13050
rect 41191 13030 42143 13046
rect 40271 13026 42143 13030
rect 42162 13026 42220 13046
rect 42239 13026 42925 13046
rect 40271 13008 42925 13026
rect 40271 13007 40372 13008
rect 42136 13004 42247 13008
rect 40455 12956 40490 12957
rect 40434 12949 40490 12956
rect 40434 12929 40463 12949
rect 40483 12929 40490 12949
rect 40434 12924 40490 12929
rect 40881 12952 40913 12959
rect 41503 12952 41538 12953
rect 40881 12932 40887 12952
rect 40908 12932 40913 12952
rect 41482 12945 41538 12952
rect 41347 12935 41405 12940
rect 40434 12646 40468 12924
rect 40881 12904 40913 12932
rect 40501 12896 40913 12904
rect 40501 12870 40507 12896
rect 40533 12870 40913 12896
rect 40501 12868 40913 12870
rect 40503 12867 40543 12868
rect 40670 12842 40701 12850
rect 40670 12812 40674 12842
rect 40695 12812 40701 12842
rect 40434 12638 40469 12646
rect 40434 12618 40442 12638
rect 40462 12618 40469 12638
rect 40434 12613 40469 12618
rect 40434 12612 40466 12613
rect 40670 12612 40701 12812
rect 40881 12803 40913 12868
rect 40881 12783 40885 12803
rect 40906 12783 40913 12803
rect 40881 12776 40913 12783
rect 41330 12926 41405 12935
rect 41330 12893 41339 12926
rect 41392 12893 41405 12926
rect 41330 12868 41405 12893
rect 41330 12835 41344 12868
rect 41397 12835 41405 12868
rect 41330 12829 41405 12835
rect 41482 12925 41511 12945
rect 41531 12925 41538 12945
rect 41482 12920 41538 12925
rect 41929 12948 41961 12955
rect 41929 12928 41935 12948
rect 41956 12928 41961 12948
rect 41190 12720 41291 12721
rect 41088 12707 41291 12720
rect 41088 12705 41231 12707
rect 41088 12702 41165 12705
rect 41088 12675 41091 12702
rect 41120 12678 41165 12702
rect 41194 12678 41231 12705
rect 41120 12675 41231 12678
rect 41088 12674 41231 12675
rect 41267 12674 41291 12707
rect 41088 12661 41291 12674
rect 40667 12605 40706 12612
rect 40665 12588 40706 12605
rect 40667 12563 40706 12588
rect 39361 12555 40706 12563
rect 39361 12527 39376 12555
rect 39404 12529 40706 12555
rect 39404 12527 40703 12529
rect 39361 12522 40703 12527
rect 41330 12518 41400 12829
rect 41482 12642 41516 12920
rect 41929 12900 41961 12928
rect 41549 12892 41961 12900
rect 41549 12866 41555 12892
rect 41581 12866 41961 12892
rect 41549 12864 41961 12866
rect 41551 12863 41591 12864
rect 41718 12838 41749 12846
rect 41718 12808 41722 12838
rect 41743 12808 41749 12838
rect 41482 12634 41517 12642
rect 41482 12614 41490 12634
rect 41510 12614 41517 12634
rect 41482 12609 41517 12614
rect 41718 12609 41749 12808
rect 41929 12799 41961 12864
rect 41929 12779 41933 12799
rect 41954 12779 41961 12799
rect 41929 12772 41961 12779
rect 42374 12925 42446 12943
rect 42374 12883 42387 12925
rect 42436 12883 42446 12925
rect 42374 12862 42446 12883
rect 42374 12820 42388 12862
rect 42437 12820 42446 12862
rect 42238 12716 42339 12717
rect 42136 12703 42339 12716
rect 42136 12701 42279 12703
rect 42136 12698 42213 12701
rect 42136 12671 42139 12698
rect 42168 12674 42213 12698
rect 42242 12674 42279 12701
rect 42168 12671 42279 12674
rect 42136 12670 42279 12671
rect 42315 12670 42339 12703
rect 42136 12657 42339 12670
rect 41482 12608 41514 12609
rect 41716 12606 41749 12609
rect 41682 12587 41750 12606
rect 41652 12575 41751 12587
rect 42374 12579 42446 12820
rect 42818 12579 42925 13008
rect 41652 12537 41674 12575
rect 41699 12540 41718 12575
rect 41743 12540 41751 12575
rect 41699 12537 41751 12540
rect 41652 12529 41751 12537
rect 41678 12528 41750 12529
rect 41329 12502 41400 12518
rect 41329 12486 41349 12502
rect 41330 12456 41349 12486
rect 41332 12436 41349 12456
rect 41379 12456 41400 12502
rect 42372 12498 42450 12579
rect 42817 12524 42925 12579
rect 41379 12436 41399 12456
rect 41332 12417 41399 12436
rect 42372 12396 42451 12498
rect 42336 12378 42457 12396
rect 42336 12376 42407 12378
rect 42336 12335 42351 12376
rect 42388 12337 42407 12376
rect 42444 12337 42457 12378
rect 42388 12335 42457 12337
rect 42336 12325 42457 12335
rect 39641 12297 39752 12300
rect 38852 12296 40505 12297
rect 42818 12296 42925 12524
rect 38852 12293 42115 12296
rect 42302 12293 42927 12296
rect 38852 12283 42927 12293
rect 38852 12263 39648 12283
rect 39667 12263 39725 12283
rect 39744 12278 42927 12283
rect 39744 12263 42143 12278
rect 38852 12258 42143 12263
rect 42162 12258 42220 12278
rect 42239 12258 42927 12278
rect 38852 12240 42927 12258
rect 38852 12237 40505 12240
rect 42136 12236 42247 12240
rect 39008 12189 39043 12190
rect 38987 12182 39043 12189
rect 38987 12162 39016 12182
rect 39036 12162 39043 12182
rect 38987 12157 39043 12162
rect 39434 12185 39466 12192
rect 39434 12165 39440 12185
rect 39461 12165 39466 12185
rect 38987 11879 39021 12157
rect 39434 12137 39466 12165
rect 41322 12177 41402 12189
rect 41503 12184 41538 12185
rect 39054 12129 39466 12137
rect 39054 12103 39060 12129
rect 39086 12103 39466 12129
rect 39852 12143 40289 12156
rect 39852 12120 39865 12143
rect 39891 12136 40289 12143
rect 39891 12120 40245 12136
rect 39852 12113 40245 12120
rect 40271 12113 40289 12136
rect 39852 12107 40289 12113
rect 41322 12151 41338 12177
rect 41378 12151 41402 12177
rect 41322 12132 41402 12151
rect 39054 12101 39466 12103
rect 39056 12100 39096 12101
rect 39223 12075 39254 12083
rect 39223 12045 39227 12075
rect 39248 12045 39254 12075
rect 38987 11871 39022 11879
rect 38987 11851 38995 11871
rect 39015 11851 39022 11871
rect 38987 11846 39022 11851
rect 38987 11845 39019 11846
rect 39223 11838 39254 12045
rect 39434 12036 39466 12101
rect 41322 12106 41341 12132
rect 41381 12106 41402 12132
rect 41322 12079 41402 12106
rect 41322 12053 41345 12079
rect 41385 12053 41402 12079
rect 41322 12042 41402 12053
rect 41482 12177 41538 12184
rect 41482 12157 41511 12177
rect 41531 12157 41538 12177
rect 41482 12152 41538 12157
rect 41929 12180 41961 12187
rect 41929 12160 41935 12180
rect 41956 12160 41961 12180
rect 39434 12016 39438 12036
rect 39459 12016 39466 12036
rect 39434 12009 39466 12016
rect 39743 11953 39844 11954
rect 39641 11940 39844 11953
rect 39641 11938 39784 11940
rect 39641 11935 39718 11938
rect 39641 11908 39644 11935
rect 39673 11911 39718 11935
rect 39747 11911 39784 11938
rect 39673 11908 39784 11911
rect 39641 11907 39784 11908
rect 39820 11907 39844 11940
rect 39641 11894 39844 11907
rect 39221 11832 39254 11838
rect 39217 11828 39254 11832
rect 39217 11818 39255 11828
rect 39217 11805 39227 11818
rect 39218 11781 39227 11805
rect 39244 11781 39255 11818
rect 39218 11760 39255 11781
rect 41327 11742 41392 12042
rect 41482 11874 41516 12152
rect 41929 12132 41961 12160
rect 41549 12124 41961 12132
rect 41549 12098 41555 12124
rect 41581 12098 41961 12124
rect 42383 12166 42450 12173
rect 42383 12145 42400 12166
rect 42436 12145 42450 12166
rect 42383 12126 42450 12145
rect 42383 12123 42400 12126
rect 41549 12096 41961 12098
rect 41551 12095 41591 12096
rect 41718 12070 41749 12078
rect 41718 12040 41722 12070
rect 41743 12040 41749 12070
rect 41482 11866 41517 11874
rect 41482 11846 41490 11866
rect 41510 11846 41517 11866
rect 41482 11841 41517 11846
rect 41482 11840 41514 11841
rect 41718 11836 41749 12040
rect 41929 12031 41961 12096
rect 42385 12089 42400 12123
rect 42440 12089 42450 12126
rect 42385 12080 42450 12089
rect 41929 12011 41933 12031
rect 41954 12011 41961 12031
rect 41929 12004 41961 12011
rect 42238 11948 42339 11949
rect 42136 11935 42339 11948
rect 42136 11933 42279 11935
rect 42136 11930 42213 11933
rect 42136 11903 42139 11930
rect 42168 11906 42213 11930
rect 42242 11906 42279 11933
rect 42168 11903 42279 11906
rect 42136 11902 42279 11903
rect 42315 11902 42339 11935
rect 42136 11889 42339 11902
rect 41716 11824 41751 11836
rect 41647 11817 41751 11824
rect 41647 11816 41723 11817
rect 41647 11796 41668 11816
rect 41700 11797 41723 11816
rect 41748 11797 41751 11817
rect 41700 11796 41751 11797
rect 41647 11787 41751 11796
rect 41716 11785 41751 11787
rect 41327 11703 41330 11742
rect 41375 11703 41392 11742
rect 42388 11719 42439 12080
rect 42386 11717 42443 11719
rect 41327 11681 41392 11703
rect 42375 11705 42443 11717
rect 42375 11672 42386 11705
rect 42426 11672 42443 11705
rect 42375 11666 42443 11672
rect 42375 11662 42439 11666
rect 41088 11617 41199 11620
rect 42818 11617 42925 12240
rect 39173 11603 42925 11617
rect 39173 11583 41095 11603
rect 41114 11583 41172 11603
rect 41191 11599 42925 11603
rect 41191 11583 42143 11599
rect 39173 11579 42143 11583
rect 42162 11579 42220 11599
rect 42239 11579 42925 11599
rect 39173 11561 42925 11579
rect 39173 11560 40464 11561
rect 42136 11557 42247 11561
rect 40455 11509 40490 11510
rect 40434 11502 40490 11509
rect 40434 11482 40463 11502
rect 40483 11482 40490 11502
rect 40434 11477 40490 11482
rect 40881 11505 40913 11512
rect 41503 11505 41538 11506
rect 40881 11485 40887 11505
rect 40908 11485 40913 11505
rect 41482 11498 41538 11505
rect 41347 11488 41405 11493
rect 40434 11199 40468 11477
rect 40881 11457 40913 11485
rect 40501 11449 40913 11457
rect 40501 11423 40507 11449
rect 40533 11423 40913 11449
rect 40501 11421 40913 11423
rect 40503 11420 40543 11421
rect 40670 11395 40701 11403
rect 40670 11365 40674 11395
rect 40695 11365 40701 11395
rect 40434 11191 40469 11199
rect 40434 11171 40442 11191
rect 40462 11171 40469 11191
rect 40434 11166 40469 11171
rect 40434 11165 40466 11166
rect 40670 11158 40701 11365
rect 40881 11356 40913 11421
rect 40881 11336 40885 11356
rect 40906 11336 40913 11356
rect 40881 11329 40913 11336
rect 41330 11479 41405 11488
rect 41330 11446 41339 11479
rect 41392 11446 41405 11479
rect 41330 11421 41405 11446
rect 41330 11388 41344 11421
rect 41397 11388 41405 11421
rect 41330 11382 41405 11388
rect 41482 11478 41511 11498
rect 41531 11478 41538 11498
rect 41482 11473 41538 11478
rect 41929 11501 41961 11508
rect 41929 11481 41935 11501
rect 41956 11481 41961 11501
rect 41190 11273 41291 11274
rect 41088 11260 41291 11273
rect 41088 11258 41231 11260
rect 41088 11255 41165 11258
rect 41088 11228 41091 11255
rect 41120 11231 41165 11255
rect 41194 11231 41231 11258
rect 41120 11228 41231 11231
rect 41088 11227 41231 11228
rect 41267 11227 41291 11260
rect 41088 11214 41291 11227
rect 40168 11145 40332 11148
rect 40665 11145 40701 11158
rect 39367 11127 40706 11145
rect 39367 11089 39377 11127
rect 39402 11112 40706 11127
rect 39402 11089 39412 11112
rect 40168 11105 40332 11112
rect 39367 11081 39412 11089
rect 39381 11080 39412 11081
rect 41330 11066 41400 11382
rect 41482 11195 41516 11473
rect 41929 11453 41961 11481
rect 41549 11445 41961 11453
rect 41549 11419 41555 11445
rect 41581 11419 41961 11445
rect 41549 11417 41961 11419
rect 41551 11416 41591 11417
rect 41718 11391 41749 11399
rect 41718 11361 41722 11391
rect 41743 11361 41749 11391
rect 41482 11187 41517 11195
rect 41482 11167 41490 11187
rect 41510 11167 41517 11187
rect 41482 11162 41517 11167
rect 41718 11162 41749 11361
rect 41929 11352 41961 11417
rect 41929 11332 41933 11352
rect 41954 11332 41961 11352
rect 41929 11325 41961 11332
rect 42374 11478 42446 11496
rect 42374 11436 42387 11478
rect 42436 11436 42446 11478
rect 42374 11415 42446 11436
rect 42374 11373 42388 11415
rect 42437 11373 42446 11415
rect 42238 11269 42339 11270
rect 42136 11256 42339 11269
rect 42136 11254 42279 11256
rect 42136 11251 42213 11254
rect 42136 11224 42139 11251
rect 42168 11227 42213 11251
rect 42242 11227 42279 11254
rect 42168 11224 42279 11227
rect 42136 11223 42279 11224
rect 42315 11223 42339 11256
rect 42136 11210 42339 11223
rect 41482 11161 41514 11162
rect 41716 11159 41749 11162
rect 41682 11140 41750 11159
rect 41652 11128 41751 11140
rect 41652 11090 41674 11128
rect 41699 11093 41718 11128
rect 41743 11093 41751 11128
rect 41699 11090 41751 11093
rect 41652 11082 41751 11090
rect 41678 11081 41750 11082
rect 41330 11047 41409 11066
rect 41333 11027 41409 11047
rect 41326 11003 41409 11027
rect 42374 11062 42446 11373
rect 42374 11019 42450 11062
rect 41326 10937 41338 11003
rect 41392 10937 41409 11003
rect 41326 10917 41409 10937
rect 41326 10880 41343 10917
rect 41387 10903 41409 10917
rect 42375 10968 42450 11019
rect 42818 10968 42925 11561
rect 41387 10880 41402 10903
rect 41326 10864 41402 10880
rect 42375 10876 42452 10968
rect 42818 10964 42926 10968
rect 42337 10858 42458 10876
rect 42337 10856 42408 10858
rect 42337 10815 42352 10856
rect 42389 10817 42408 10856
rect 42445 10817 42458 10858
rect 42389 10815 42458 10817
rect 42337 10805 42458 10815
rect 38862 10776 40331 10778
rect 42819 10776 42926 10964
rect 38862 10761 42928 10776
rect 38862 10741 39606 10761
rect 39625 10741 39683 10761
rect 39702 10758 42928 10761
rect 39702 10741 42144 10758
rect 38862 10738 42144 10741
rect 42163 10738 42221 10758
rect 42240 10738 42928 10758
rect 38862 10720 42928 10738
rect 39599 10719 39710 10720
rect 40286 10719 40493 10720
rect 42137 10716 42248 10720
rect 38966 10667 39001 10668
rect 38945 10660 39001 10667
rect 38945 10640 38974 10660
rect 38994 10640 39001 10660
rect 38945 10635 39001 10640
rect 39392 10663 39424 10670
rect 39392 10643 39398 10663
rect 39419 10643 39424 10663
rect 38945 10357 38979 10635
rect 39392 10615 39424 10643
rect 39012 10607 39424 10615
rect 39012 10581 39018 10607
rect 39044 10581 39424 10607
rect 39012 10579 39424 10581
rect 39014 10578 39054 10579
rect 39181 10553 39212 10561
rect 39181 10523 39185 10553
rect 39206 10523 39212 10553
rect 38945 10349 38980 10357
rect 38945 10329 38953 10349
rect 38973 10329 38980 10349
rect 38945 10324 38980 10329
rect 39181 10327 39212 10523
rect 39392 10514 39424 10579
rect 41323 10657 41403 10669
rect 41504 10664 41539 10665
rect 41323 10631 41339 10657
rect 41379 10631 41403 10657
rect 41323 10612 41403 10631
rect 41323 10586 41342 10612
rect 41382 10586 41403 10612
rect 41323 10559 41403 10586
rect 41323 10533 41346 10559
rect 41386 10533 41403 10559
rect 41323 10522 41403 10533
rect 41483 10657 41539 10664
rect 41483 10637 41512 10657
rect 41532 10637 41539 10657
rect 41483 10632 41539 10637
rect 41930 10660 41962 10667
rect 41930 10640 41936 10660
rect 41957 10640 41962 10660
rect 39392 10494 39396 10514
rect 39417 10494 39424 10514
rect 39392 10487 39424 10494
rect 39701 10431 39802 10432
rect 39599 10418 39802 10431
rect 39599 10416 39742 10418
rect 39599 10413 39676 10416
rect 39599 10386 39602 10413
rect 39631 10389 39676 10413
rect 39705 10389 39742 10416
rect 39631 10386 39742 10389
rect 39599 10385 39742 10386
rect 39778 10385 39802 10418
rect 39599 10372 39802 10385
rect 38945 10323 38977 10324
rect 39181 10238 39215 10327
rect 38802 10234 39215 10238
rect 37788 7909 37805 7963
rect 37868 7909 37893 7963
rect 37788 7888 37893 7909
rect 38255 10189 39215 10234
rect 41328 10222 41393 10522
rect 41483 10354 41517 10632
rect 41930 10612 41962 10640
rect 41550 10604 41962 10612
rect 41550 10578 41556 10604
rect 41582 10578 41962 10604
rect 42384 10646 42451 10653
rect 42384 10625 42401 10646
rect 42437 10625 42451 10646
rect 42384 10606 42451 10625
rect 42384 10603 42401 10606
rect 41550 10576 41962 10578
rect 41552 10575 41592 10576
rect 41719 10550 41750 10558
rect 41719 10520 41723 10550
rect 41744 10520 41750 10550
rect 41483 10346 41518 10354
rect 41483 10326 41491 10346
rect 41511 10326 41518 10346
rect 41483 10321 41518 10326
rect 41483 10320 41515 10321
rect 41719 10316 41750 10520
rect 41930 10511 41962 10576
rect 42386 10569 42401 10603
rect 42441 10569 42451 10606
rect 42386 10560 42451 10569
rect 41930 10491 41934 10511
rect 41955 10491 41962 10511
rect 41930 10484 41962 10491
rect 42239 10428 42340 10429
rect 42137 10415 42340 10428
rect 42137 10413 42280 10415
rect 42137 10410 42214 10413
rect 42137 10383 42140 10410
rect 42169 10386 42214 10410
rect 42243 10386 42280 10413
rect 42169 10383 42280 10386
rect 42137 10382 42280 10383
rect 42316 10382 42340 10415
rect 42137 10369 42340 10382
rect 41717 10304 41752 10316
rect 41648 10297 41752 10304
rect 41648 10296 41724 10297
rect 41648 10276 41669 10296
rect 41701 10277 41724 10296
rect 41749 10277 41752 10297
rect 41701 10276 41752 10277
rect 41648 10267 41752 10276
rect 41717 10265 41752 10267
rect 38255 10185 38852 10189
rect 38255 7879 38307 10185
rect 41328 10183 41331 10222
rect 41376 10183 41393 10222
rect 42389 10199 42440 10560
rect 42387 10197 42444 10199
rect 41328 10161 41393 10183
rect 42376 10185 42444 10197
rect 42376 10152 42387 10185
rect 42427 10152 42444 10185
rect 42376 10146 42444 10152
rect 42376 10142 42440 10146
rect 41089 10097 41200 10100
rect 42819 10097 42926 10720
rect 39214 10083 42926 10097
rect 39214 10063 41096 10083
rect 41115 10063 41173 10083
rect 41192 10079 42926 10083
rect 41192 10063 42144 10079
rect 39214 10059 42144 10063
rect 42163 10059 42221 10079
rect 42240 10059 42926 10079
rect 39214 10041 42926 10059
rect 39214 10040 40373 10041
rect 42137 10037 42248 10041
rect 40456 9989 40491 9990
rect 40435 9982 40491 9989
rect 40435 9962 40464 9982
rect 40484 9962 40491 9982
rect 40435 9957 40491 9962
rect 40882 9985 40914 9992
rect 41504 9985 41539 9986
rect 40882 9965 40888 9985
rect 40909 9965 40914 9985
rect 41483 9978 41539 9985
rect 41348 9968 41406 9973
rect 40435 9679 40469 9957
rect 40882 9937 40914 9965
rect 40502 9929 40914 9937
rect 40502 9903 40508 9929
rect 40534 9903 40914 9929
rect 40502 9901 40914 9903
rect 40504 9900 40544 9901
rect 40671 9875 40702 9883
rect 40671 9845 40675 9875
rect 40696 9845 40702 9875
rect 40435 9671 40470 9679
rect 40435 9651 40443 9671
rect 40463 9651 40470 9671
rect 40435 9646 40470 9651
rect 39176 9635 39212 9646
rect 40435 9645 40467 9646
rect 40671 9638 40702 9845
rect 40882 9836 40914 9901
rect 40882 9816 40886 9836
rect 40907 9816 40914 9836
rect 40882 9809 40914 9816
rect 41331 9959 41406 9968
rect 41331 9926 41340 9959
rect 41393 9926 41406 9959
rect 41331 9901 41406 9926
rect 41331 9868 41345 9901
rect 41398 9868 41406 9901
rect 41331 9862 41406 9868
rect 41483 9958 41512 9978
rect 41532 9958 41539 9978
rect 41483 9953 41539 9958
rect 41930 9981 41962 9988
rect 41930 9961 41936 9981
rect 41957 9961 41962 9981
rect 41191 9753 41292 9754
rect 41089 9740 41292 9753
rect 41089 9738 41232 9740
rect 41089 9735 41166 9738
rect 41089 9708 41092 9735
rect 41121 9711 41166 9735
rect 41195 9711 41232 9738
rect 41121 9708 41232 9711
rect 41089 9707 41232 9708
rect 41268 9707 41292 9740
rect 41089 9694 41292 9707
rect 39176 9612 39182 9635
rect 39206 9612 39212 9635
rect 40666 9629 40702 9638
rect 40611 9619 40708 9629
rect 39423 9617 40708 9619
rect 39176 9591 39212 9612
rect 39176 9568 39182 9591
rect 39206 9568 39212 9591
rect 39176 9415 39212 9568
rect 39388 9607 40708 9617
rect 39388 9569 39400 9607
rect 39425 9572 39444 9607
rect 39469 9572 40708 9607
rect 39425 9569 40708 9572
rect 39388 9566 40708 9569
rect 39388 9564 40705 9566
rect 39388 9561 39477 9564
rect 39404 9560 39476 9561
rect 41331 9551 41401 9862
rect 41483 9675 41517 9953
rect 41930 9933 41962 9961
rect 41550 9925 41962 9933
rect 41550 9899 41556 9925
rect 41582 9899 41962 9925
rect 41550 9897 41962 9899
rect 41552 9896 41592 9897
rect 41719 9871 41750 9879
rect 41719 9841 41723 9871
rect 41744 9841 41750 9871
rect 41483 9667 41518 9675
rect 41483 9647 41491 9667
rect 41511 9647 41518 9667
rect 41483 9642 41518 9647
rect 41719 9642 41750 9841
rect 41930 9832 41962 9897
rect 41930 9812 41934 9832
rect 41955 9812 41962 9832
rect 41930 9805 41962 9812
rect 42375 9958 42447 9976
rect 42375 9916 42388 9958
rect 42437 9916 42447 9958
rect 42375 9895 42447 9916
rect 42375 9853 42389 9895
rect 42438 9853 42447 9895
rect 42239 9749 42340 9750
rect 42137 9736 42340 9749
rect 42137 9734 42280 9736
rect 42137 9731 42214 9734
rect 42137 9704 42140 9731
rect 42169 9707 42214 9731
rect 42243 9707 42280 9734
rect 42169 9704 42280 9707
rect 42137 9703 42280 9704
rect 42316 9703 42340 9736
rect 42137 9690 42340 9703
rect 41483 9641 41515 9642
rect 41717 9639 41750 9642
rect 41683 9620 41751 9639
rect 41653 9608 41752 9620
rect 42375 9612 42447 9853
rect 42819 9612 42926 10041
rect 41653 9570 41675 9608
rect 41700 9573 41719 9608
rect 41744 9573 41752 9608
rect 41700 9570 41752 9573
rect 41653 9562 41752 9570
rect 41679 9561 41751 9562
rect 41330 9535 41401 9551
rect 41330 9519 41350 9535
rect 41331 9489 41350 9519
rect 41333 9469 41350 9489
rect 41380 9489 41401 9535
rect 42373 9531 42451 9612
rect 42818 9557 42926 9612
rect 41380 9469 41400 9489
rect 41333 9450 41400 9469
rect 42373 9429 42452 9531
rect 39167 9406 39253 9415
rect 39167 9388 39186 9406
rect 39238 9388 39253 9406
rect 39167 9384 39253 9388
rect 42337 9411 42458 9429
rect 42337 9409 42408 9411
rect 42337 9368 42352 9409
rect 42389 9370 42408 9409
rect 42445 9370 42458 9411
rect 42389 9368 42458 9370
rect 42337 9358 42458 9368
rect 39642 9330 39753 9333
rect 38862 9329 40506 9330
rect 42819 9329 42926 9557
rect 38862 9326 42116 9329
rect 42303 9326 42928 9329
rect 38862 9316 42928 9326
rect 38862 9296 39649 9316
rect 39668 9296 39726 9316
rect 39745 9311 42928 9316
rect 39745 9296 42144 9311
rect 38862 9291 42144 9296
rect 42163 9291 42221 9311
rect 42240 9291 42928 9311
rect 38862 9273 42928 9291
rect 38862 9270 40506 9273
rect 42137 9269 42248 9273
rect 39009 9222 39044 9223
rect 38988 9215 39044 9222
rect 38988 9195 39017 9215
rect 39037 9195 39044 9215
rect 38988 9190 39044 9195
rect 39435 9218 39467 9225
rect 39435 9198 39441 9218
rect 39462 9198 39467 9218
rect 38988 8912 39022 9190
rect 39435 9170 39467 9198
rect 39055 9162 39467 9170
rect 39055 9136 39061 9162
rect 39087 9136 39467 9162
rect 39055 9134 39467 9136
rect 39057 9133 39097 9134
rect 39224 9108 39255 9116
rect 39224 9078 39228 9108
rect 39249 9078 39255 9108
rect 38988 8904 39023 8912
rect 38988 8884 38996 8904
rect 39016 8884 39023 8904
rect 38988 8879 39023 8884
rect 38988 8878 39020 8879
rect 39224 8877 39255 9078
rect 39435 9069 39467 9134
rect 39435 9049 39439 9069
rect 39460 9049 39467 9069
rect 39435 9042 39467 9049
rect 40029 9209 40122 9216
rect 40029 9168 40053 9209
rect 40107 9168 40122 9209
rect 39744 8986 39845 8987
rect 39642 8973 39845 8986
rect 39642 8971 39785 8973
rect 39642 8968 39719 8971
rect 39642 8941 39645 8968
rect 39674 8944 39719 8968
rect 39748 8944 39785 8971
rect 39674 8941 39785 8944
rect 39642 8940 39785 8941
rect 39821 8940 39845 8973
rect 39642 8927 39845 8940
rect 40029 8795 40122 9168
rect 41323 9210 41403 9222
rect 41504 9217 41539 9218
rect 41323 9184 41339 9210
rect 41379 9184 41403 9210
rect 41323 9165 41403 9184
rect 41323 9139 41342 9165
rect 41382 9139 41403 9165
rect 41323 9112 41403 9139
rect 41323 9086 41346 9112
rect 41386 9086 41403 9112
rect 41323 9075 41403 9086
rect 41483 9210 41539 9217
rect 41483 9190 41512 9210
rect 41532 9190 41539 9210
rect 41483 9185 41539 9190
rect 41930 9213 41962 9220
rect 41930 9193 41936 9213
rect 41957 9193 41962 9213
rect 40029 8751 40047 8795
rect 40107 8751 40122 8795
rect 40029 8736 40122 8751
rect 41328 8775 41393 9075
rect 41483 8907 41517 9185
rect 41930 9165 41962 9193
rect 41550 9157 41962 9165
rect 41550 9131 41556 9157
rect 41582 9131 41962 9157
rect 42384 9199 42451 9206
rect 42384 9178 42401 9199
rect 42437 9178 42451 9199
rect 42384 9159 42451 9178
rect 42384 9156 42401 9159
rect 41550 9129 41962 9131
rect 41552 9128 41592 9129
rect 41719 9103 41750 9111
rect 41719 9073 41723 9103
rect 41744 9073 41750 9103
rect 41483 8899 41518 8907
rect 41483 8879 41491 8899
rect 41511 8879 41518 8899
rect 41483 8874 41518 8879
rect 41483 8873 41515 8874
rect 41719 8869 41750 9073
rect 41930 9064 41962 9129
rect 42386 9122 42401 9156
rect 42441 9122 42451 9159
rect 42386 9113 42451 9122
rect 41930 9044 41934 9064
rect 41955 9044 41962 9064
rect 41930 9037 41962 9044
rect 42239 8981 42340 8982
rect 42137 8968 42340 8981
rect 42137 8966 42280 8968
rect 42137 8963 42214 8966
rect 42137 8936 42140 8963
rect 42169 8939 42214 8963
rect 42243 8939 42280 8966
rect 42169 8936 42280 8939
rect 42137 8935 42280 8936
rect 42316 8935 42340 8968
rect 42137 8922 42340 8935
rect 41717 8857 41752 8869
rect 41648 8850 41752 8857
rect 41648 8849 41724 8850
rect 41648 8829 41669 8849
rect 41701 8830 41724 8849
rect 41749 8830 41752 8850
rect 41701 8829 41752 8830
rect 41648 8820 41752 8829
rect 41717 8818 41752 8820
rect 41328 8736 41331 8775
rect 41376 8736 41393 8775
rect 42389 8752 42440 9113
rect 42387 8750 42444 8752
rect 41328 8714 41393 8736
rect 42376 8738 42444 8750
rect 42376 8705 42387 8738
rect 42427 8705 42444 8738
rect 42376 8699 42444 8705
rect 42376 8695 42440 8699
rect 41089 8650 41200 8653
rect 42819 8650 42926 9273
rect 38895 8636 42926 8650
rect 38895 8616 41096 8636
rect 41115 8616 41173 8636
rect 41192 8632 42926 8636
rect 41192 8616 42144 8632
rect 38895 8612 42144 8616
rect 42163 8612 42221 8632
rect 42240 8612 42926 8632
rect 38895 8594 42926 8612
rect 38895 8593 40465 8594
rect 42137 8590 42248 8594
rect 40456 8542 40491 8543
rect 40435 8535 40491 8542
rect 40435 8515 40464 8535
rect 40484 8515 40491 8535
rect 40435 8510 40491 8515
rect 40882 8538 40914 8545
rect 41504 8538 41539 8539
rect 40882 8518 40888 8538
rect 40909 8518 40914 8538
rect 41483 8531 41539 8538
rect 41348 8521 41406 8526
rect 40035 8455 40117 8484
rect 40035 8414 40060 8455
rect 40096 8414 40117 8455
rect 40222 8475 40286 8494
rect 40222 8436 40239 8475
rect 40273 8436 40286 8475
rect 40222 8417 40286 8436
rect 40035 8099 40117 8414
rect 40027 8054 40117 8099
rect 40224 8072 40286 8417
rect 40435 8232 40469 8510
rect 40882 8490 40914 8518
rect 40502 8482 40914 8490
rect 40502 8456 40508 8482
rect 40534 8456 40914 8482
rect 40502 8454 40914 8456
rect 40504 8453 40544 8454
rect 40671 8428 40702 8436
rect 40671 8398 40675 8428
rect 40696 8398 40702 8428
rect 40435 8224 40470 8232
rect 40435 8204 40443 8224
rect 40463 8204 40470 8224
rect 40435 8199 40470 8204
rect 40435 8198 40467 8199
rect 40671 8191 40702 8398
rect 40882 8389 40914 8454
rect 40882 8369 40886 8389
rect 40907 8369 40914 8389
rect 40882 8362 40914 8369
rect 41331 8512 41406 8521
rect 41331 8479 41340 8512
rect 41393 8479 41406 8512
rect 41331 8454 41406 8479
rect 41331 8421 41345 8454
rect 41398 8421 41406 8454
rect 41331 8415 41406 8421
rect 41483 8511 41512 8531
rect 41532 8511 41539 8531
rect 41483 8506 41539 8511
rect 41930 8534 41962 8541
rect 41930 8514 41936 8534
rect 41957 8514 41962 8534
rect 41191 8306 41292 8307
rect 41089 8293 41292 8306
rect 41089 8291 41232 8293
rect 41089 8288 41166 8291
rect 41089 8261 41092 8288
rect 41121 8264 41166 8288
rect 41195 8264 41232 8291
rect 41121 8261 41232 8264
rect 41089 8260 41232 8261
rect 41268 8260 41292 8293
rect 41089 8247 41292 8260
rect 40666 8173 40702 8191
rect 40633 8172 40702 8173
rect 40613 8160 40702 8172
rect 40613 8122 40625 8160
rect 40650 8125 40669 8160
rect 40694 8125 40702 8160
rect 41331 8149 41401 8415
rect 41483 8228 41517 8506
rect 41930 8486 41962 8514
rect 41550 8478 41962 8486
rect 41550 8452 41556 8478
rect 41582 8452 41962 8478
rect 41550 8450 41962 8452
rect 41552 8449 41592 8450
rect 41719 8424 41750 8432
rect 41719 8394 41723 8424
rect 41744 8394 41750 8424
rect 41483 8220 41518 8228
rect 41483 8200 41491 8220
rect 41511 8200 41518 8220
rect 41483 8195 41518 8200
rect 41719 8195 41750 8394
rect 41930 8385 41962 8450
rect 41930 8365 41934 8385
rect 41955 8365 41962 8385
rect 41930 8358 41962 8365
rect 42375 8511 42447 8529
rect 42375 8469 42388 8511
rect 42437 8469 42447 8511
rect 42375 8448 42447 8469
rect 42375 8406 42389 8448
rect 42438 8406 42447 8448
rect 42239 8302 42340 8303
rect 42137 8289 42340 8302
rect 42137 8287 42280 8289
rect 42137 8284 42214 8287
rect 42137 8257 42140 8284
rect 42169 8260 42214 8284
rect 42243 8260 42280 8287
rect 42169 8257 42280 8260
rect 42137 8256 42280 8257
rect 42316 8256 42340 8289
rect 42137 8243 42340 8256
rect 41483 8194 41515 8195
rect 41717 8192 41750 8195
rect 41683 8173 41751 8192
rect 40650 8122 40702 8125
rect 40613 8114 40702 8122
rect 41322 8120 41401 8149
rect 41653 8161 41752 8173
rect 41653 8123 41675 8161
rect 41700 8126 41719 8161
rect 41744 8126 41752 8161
rect 41700 8123 41752 8126
rect 40629 8113 40701 8114
rect 40223 8063 40297 8072
rect 40027 8021 40111 8054
rect 40027 7993 40042 8021
rect 40086 7993 40111 8021
rect 40027 7964 40111 7993
rect 40223 8015 40237 8063
rect 40274 8015 40297 8063
rect 40223 7987 40297 8015
rect 40027 7936 40039 7964
rect 40083 7936 40111 7964
rect 40027 7925 40111 7936
rect 41322 7937 41399 8120
rect 41653 8115 41752 8123
rect 41679 8114 41751 8115
rect 42375 8112 42447 8406
rect 42819 8134 42926 8594
rect 42375 8074 42451 8112
rect 42819 8074 42932 8134
rect 42386 7973 42451 8074
rect 41322 7894 41339 7937
rect 38255 7845 38270 7879
rect 38299 7845 38307 7879
rect 41327 7889 41339 7894
rect 41385 7889 41399 7937
rect 41327 7867 41399 7889
rect 42384 7927 42451 7973
rect 42821 7935 42932 8074
rect 38255 7819 38307 7845
rect 42384 7835 42449 7927
rect 42816 7908 42932 7935
rect 38255 7785 38269 7819
rect 38298 7785 38307 7819
rect 38255 7754 38307 7785
rect 42334 7817 42455 7835
rect 42334 7815 42405 7817
rect 42334 7774 42349 7815
rect 42386 7776 42405 7815
rect 42442 7776 42455 7817
rect 42386 7774 42455 7776
rect 42334 7764 42455 7774
rect 38531 7737 38642 7743
rect 38531 7735 40328 7737
rect 42816 7735 42923 7908
rect 38531 7726 42925 7735
rect 38531 7706 38538 7726
rect 38557 7706 38615 7726
rect 38634 7717 42925 7726
rect 38634 7706 42141 7717
rect 38531 7697 42141 7706
rect 42160 7697 42218 7717
rect 42237 7697 42925 7717
rect 38531 7684 42925 7697
rect 38850 7679 42925 7684
rect 40283 7678 40490 7679
rect 42134 7675 42245 7679
rect 37898 7632 37933 7633
rect 37877 7625 37933 7632
rect 37877 7605 37906 7625
rect 37926 7605 37933 7625
rect 37877 7600 37933 7605
rect 38324 7628 38356 7635
rect 38324 7608 38330 7628
rect 38351 7608 38356 7628
rect 37877 7322 37911 7600
rect 38324 7580 38356 7608
rect 41320 7616 41400 7628
rect 41501 7623 41536 7624
rect 41320 7590 41336 7616
rect 41376 7590 41400 7616
rect 37944 7572 38356 7580
rect 37944 7546 37950 7572
rect 37976 7546 38356 7572
rect 37944 7544 38356 7546
rect 37946 7543 37986 7544
rect 38113 7518 38144 7526
rect 38113 7488 38117 7518
rect 38138 7488 38144 7518
rect 37877 7314 37912 7322
rect 37877 7294 37885 7314
rect 37905 7294 37912 7314
rect 38113 7303 38144 7488
rect 38324 7479 38356 7544
rect 38738 7577 38849 7584
rect 38738 7576 38817 7577
rect 38738 7552 38760 7576
rect 38784 7553 38817 7576
rect 38841 7553 38849 7577
rect 38784 7552 38849 7553
rect 38738 7542 38849 7552
rect 41320 7571 41400 7590
rect 41320 7545 41339 7571
rect 41379 7545 41400 7571
rect 38799 7525 38848 7542
rect 41320 7518 41400 7545
rect 41320 7492 41343 7518
rect 41383 7492 41400 7518
rect 41320 7481 41400 7492
rect 41480 7616 41536 7623
rect 41480 7596 41509 7616
rect 41529 7596 41536 7616
rect 41480 7591 41536 7596
rect 41927 7619 41959 7626
rect 41927 7599 41933 7619
rect 41954 7599 41959 7619
rect 38324 7459 38328 7479
rect 38349 7459 38356 7479
rect 38324 7452 38356 7459
rect 38633 7396 38734 7397
rect 38531 7383 38734 7396
rect 38531 7381 38674 7383
rect 38531 7378 38608 7381
rect 38531 7351 38534 7378
rect 38563 7354 38608 7378
rect 38637 7354 38674 7381
rect 38563 7351 38674 7354
rect 38531 7350 38674 7351
rect 38710 7350 38734 7383
rect 38531 7337 38734 7350
rect 37877 7289 37912 7294
rect 37877 7288 37909 7289
rect 38111 7226 38145 7303
rect 36744 5823 37341 5827
rect 33844 5745 33879 5747
rect 33844 5736 33948 5745
rect 33844 5735 33895 5736
rect 33844 5715 33847 5735
rect 33872 5716 33895 5735
rect 33927 5716 33948 5736
rect 33872 5715 33948 5716
rect 33844 5708 33948 5715
rect 33844 5696 33879 5708
rect 33256 5630 33459 5643
rect 33256 5597 33280 5630
rect 33316 5629 33459 5630
rect 33316 5626 33427 5629
rect 33316 5599 33353 5626
rect 33382 5602 33427 5626
rect 33456 5602 33459 5629
rect 33382 5599 33459 5602
rect 33316 5597 33459 5599
rect 33256 5584 33459 5597
rect 33256 5583 33357 5584
rect 33634 5521 33666 5528
rect 33634 5501 33641 5521
rect 33662 5501 33666 5521
rect 33145 5443 33210 5452
rect 33145 5406 33155 5443
rect 33195 5409 33210 5443
rect 33634 5436 33666 5501
rect 33846 5492 33877 5696
rect 34081 5691 34113 5692
rect 34078 5686 34113 5691
rect 34078 5666 34085 5686
rect 34105 5666 34113 5686
rect 34078 5658 34113 5666
rect 33846 5462 33852 5492
rect 33873 5462 33877 5492
rect 33846 5454 33877 5462
rect 34004 5436 34044 5437
rect 33634 5434 34046 5436
rect 33195 5406 33212 5409
rect 33145 5387 33212 5406
rect 33145 5366 33159 5387
rect 33195 5366 33212 5387
rect 33145 5359 33212 5366
rect 33634 5408 34014 5434
rect 34040 5408 34046 5434
rect 33634 5400 34046 5408
rect 33634 5372 33666 5400
rect 34079 5380 34113 5658
rect 34203 5490 34268 5790
rect 36381 5778 37341 5823
rect 37448 6166 37484 6794
rect 36381 5774 36794 5778
rect 36381 5685 36415 5774
rect 36619 5688 36651 5689
rect 35794 5627 35997 5640
rect 35794 5594 35818 5627
rect 35854 5626 35997 5627
rect 35854 5623 35965 5626
rect 35854 5596 35891 5623
rect 35920 5599 35965 5623
rect 35994 5599 35997 5626
rect 35920 5596 35997 5599
rect 35854 5594 35997 5596
rect 35794 5581 35997 5594
rect 35794 5580 35895 5581
rect 36172 5518 36204 5525
rect 36172 5498 36179 5518
rect 36200 5498 36204 5518
rect 33634 5352 33639 5372
rect 33660 5352 33666 5372
rect 33634 5345 33666 5352
rect 34057 5375 34113 5380
rect 34057 5355 34064 5375
rect 34084 5355 34113 5375
rect 34057 5348 34113 5355
rect 34193 5479 34273 5490
rect 34193 5453 34210 5479
rect 34250 5453 34273 5479
rect 34193 5426 34273 5453
rect 34193 5400 34214 5426
rect 34254 5400 34273 5426
rect 34193 5381 34273 5400
rect 34193 5355 34217 5381
rect 34257 5355 34273 5381
rect 34057 5347 34092 5348
rect 34193 5343 34273 5355
rect 36172 5433 36204 5498
rect 36384 5489 36415 5685
rect 36616 5683 36651 5688
rect 36616 5663 36623 5683
rect 36643 5663 36651 5683
rect 36616 5655 36651 5663
rect 36384 5459 36390 5489
rect 36411 5459 36415 5489
rect 36384 5451 36415 5459
rect 36542 5433 36582 5434
rect 36172 5431 36584 5433
rect 36172 5405 36552 5431
rect 36578 5405 36584 5431
rect 36172 5397 36584 5405
rect 36172 5369 36204 5397
rect 36617 5377 36651 5655
rect 36172 5349 36177 5369
rect 36198 5349 36204 5369
rect 36172 5342 36204 5349
rect 36595 5372 36651 5377
rect 36595 5352 36602 5372
rect 36622 5352 36651 5372
rect 36595 5345 36651 5352
rect 36595 5344 36630 5345
rect 33348 5292 33459 5296
rect 35103 5292 35310 5293
rect 35886 5292 35997 5293
rect 32668 5274 36734 5292
rect 32668 5254 33356 5274
rect 33375 5254 33433 5274
rect 33452 5271 36734 5274
rect 33452 5254 35894 5271
rect 32668 5251 35894 5254
rect 35913 5251 35971 5271
rect 35990 5251 36734 5271
rect 32668 5236 36734 5251
rect 32670 5048 32777 5236
rect 35265 5234 36734 5236
rect 33138 5197 33259 5207
rect 33138 5195 33207 5197
rect 33138 5154 33151 5195
rect 33188 5156 33207 5195
rect 33244 5156 33259 5197
rect 33188 5154 33259 5156
rect 33138 5136 33259 5154
rect 32670 5044 32778 5048
rect 33144 5044 33221 5136
rect 34194 5132 34270 5148
rect 34194 5109 34209 5132
rect 30677 4878 30692 4901
rect 30616 4862 30692 4878
rect 31665 4874 31742 4966
rect 32108 4962 32216 4966
rect 31627 4856 31748 4874
rect 31627 4854 31698 4856
rect 31627 4813 31642 4854
rect 31679 4815 31698 4854
rect 31735 4815 31748 4856
rect 31679 4813 31748 4815
rect 31627 4803 31748 4813
rect 28198 4774 29621 4776
rect 32109 4774 32216 4962
rect 28198 4759 32218 4774
rect 28198 4739 28896 4759
rect 28915 4739 28973 4759
rect 28992 4756 32218 4759
rect 28992 4739 31434 4756
rect 28198 4736 31434 4739
rect 31453 4736 31511 4756
rect 31530 4736 32218 4756
rect 28198 4718 32218 4736
rect 28889 4717 29000 4718
rect 29576 4717 29783 4718
rect 31427 4714 31538 4718
rect 28256 4665 28291 4666
rect 28235 4658 28291 4665
rect 28235 4638 28264 4658
rect 28284 4638 28291 4658
rect 28235 4633 28291 4638
rect 28682 4661 28714 4668
rect 28682 4641 28688 4661
rect 28709 4641 28714 4661
rect 27404 4409 27430 4424
rect 27401 4402 27437 4409
rect 27401 4364 27407 4402
rect 27430 4364 27437 4402
rect 27401 4358 27437 4364
rect 28235 4355 28269 4633
rect 28682 4613 28714 4641
rect 28302 4605 28714 4613
rect 28302 4579 28308 4605
rect 28334 4579 28714 4605
rect 28302 4577 28714 4579
rect 28304 4576 28344 4577
rect 28471 4551 28502 4559
rect 28471 4521 28475 4551
rect 28496 4521 28502 4551
rect 28235 4347 28270 4355
rect 28235 4327 28243 4347
rect 28263 4327 28270 4347
rect 28235 4322 28270 4327
rect 28235 4321 28267 4322
rect 28471 4318 28502 4521
rect 28682 4512 28714 4577
rect 30613 4655 30693 4667
rect 30794 4662 30829 4663
rect 30613 4629 30629 4655
rect 30669 4629 30693 4655
rect 30613 4610 30693 4629
rect 30613 4584 30632 4610
rect 30672 4584 30693 4610
rect 30613 4557 30693 4584
rect 30613 4531 30636 4557
rect 30676 4531 30693 4557
rect 30613 4520 30693 4531
rect 30773 4655 30829 4662
rect 30773 4635 30802 4655
rect 30822 4635 30829 4655
rect 30773 4630 30829 4635
rect 31220 4658 31252 4665
rect 31220 4638 31226 4658
rect 31247 4638 31252 4658
rect 28682 4492 28686 4512
rect 28707 4492 28714 4512
rect 28682 4485 28714 4492
rect 28991 4429 29092 4430
rect 28889 4416 29092 4429
rect 28889 4414 29032 4416
rect 28889 4411 28966 4414
rect 28889 4384 28892 4411
rect 28921 4387 28966 4411
rect 28995 4387 29032 4414
rect 28921 4384 29032 4387
rect 28889 4383 29032 4384
rect 29068 4383 29092 4416
rect 28889 4370 29092 4383
rect 28466 4300 28502 4318
rect 28466 4283 28501 4300
rect 28399 4252 28504 4283
rect 28399 4247 28471 4252
rect 28399 4226 28430 4247
rect 28450 4231 28471 4247
rect 28491 4231 28504 4252
rect 28450 4226 28504 4231
rect 28399 4217 28504 4226
rect 30618 4220 30683 4520
rect 30773 4352 30807 4630
rect 31220 4610 31252 4638
rect 30840 4602 31252 4610
rect 30840 4576 30846 4602
rect 30872 4576 31252 4602
rect 31674 4644 31741 4651
rect 31674 4623 31691 4644
rect 31727 4623 31741 4644
rect 31674 4604 31741 4623
rect 31674 4601 31691 4604
rect 30840 4574 31252 4576
rect 30842 4573 30882 4574
rect 31009 4548 31040 4556
rect 31009 4518 31013 4548
rect 31034 4518 31040 4548
rect 30773 4344 30808 4352
rect 30773 4324 30781 4344
rect 30801 4324 30808 4344
rect 30773 4319 30808 4324
rect 30773 4318 30805 4319
rect 31009 4314 31040 4518
rect 31220 4509 31252 4574
rect 31676 4567 31691 4601
rect 31731 4567 31741 4604
rect 31676 4558 31741 4567
rect 31220 4489 31224 4509
rect 31245 4489 31252 4509
rect 31220 4482 31252 4489
rect 31529 4426 31630 4427
rect 31427 4413 31630 4426
rect 31427 4411 31570 4413
rect 31427 4408 31504 4411
rect 31427 4381 31430 4408
rect 31459 4384 31504 4408
rect 31533 4384 31570 4411
rect 31459 4381 31570 4384
rect 31427 4380 31570 4381
rect 31606 4380 31630 4413
rect 31427 4367 31630 4380
rect 31007 4302 31042 4314
rect 30938 4295 31042 4302
rect 30938 4294 31014 4295
rect 30938 4274 30959 4294
rect 30991 4275 31014 4294
rect 31039 4275 31042 4295
rect 30991 4274 31042 4275
rect 30938 4265 31042 4274
rect 31007 4263 31042 4265
rect 30618 4181 30621 4220
rect 30666 4181 30683 4220
rect 31679 4197 31730 4558
rect 31677 4195 31734 4197
rect 30618 4159 30683 4181
rect 31666 4183 31734 4195
rect 31666 4150 31677 4183
rect 31717 4150 31734 4183
rect 31666 4144 31734 4150
rect 31666 4140 31730 4144
rect 30379 4095 30490 4098
rect 32109 4095 32216 4718
rect 28422 4081 32216 4095
rect 28422 4061 30386 4081
rect 30405 4061 30463 4081
rect 30482 4077 32216 4081
rect 30482 4061 31434 4077
rect 28422 4057 31434 4061
rect 31453 4057 31511 4077
rect 31530 4057 32216 4077
rect 28422 4039 32216 4057
rect 28422 4038 29663 4039
rect 31427 4035 31538 4039
rect 29746 3987 29781 3988
rect 29725 3980 29781 3987
rect 29725 3960 29754 3980
rect 29774 3960 29781 3980
rect 29725 3955 29781 3960
rect 30172 3983 30204 3990
rect 30794 3983 30829 3984
rect 30172 3963 30178 3983
rect 30199 3963 30204 3983
rect 30773 3976 30829 3983
rect 30638 3966 30696 3971
rect 29725 3677 29759 3955
rect 30172 3935 30204 3963
rect 29792 3927 30204 3935
rect 29792 3901 29798 3927
rect 29824 3901 30204 3927
rect 29792 3899 30204 3901
rect 29794 3898 29834 3899
rect 29961 3873 29992 3881
rect 29961 3843 29965 3873
rect 29986 3843 29992 3873
rect 29725 3669 29760 3677
rect 29725 3649 29733 3669
rect 29753 3649 29760 3669
rect 29725 3644 29760 3649
rect 28466 3633 28502 3644
rect 29725 3643 29757 3644
rect 29961 3636 29992 3843
rect 30172 3834 30204 3899
rect 30172 3814 30176 3834
rect 30197 3814 30204 3834
rect 30172 3807 30204 3814
rect 30621 3957 30696 3966
rect 30621 3924 30630 3957
rect 30683 3924 30696 3957
rect 30621 3899 30696 3924
rect 30621 3866 30635 3899
rect 30688 3866 30696 3899
rect 30621 3860 30696 3866
rect 30773 3956 30802 3976
rect 30822 3956 30829 3976
rect 30773 3951 30829 3956
rect 31220 3979 31252 3986
rect 31220 3959 31226 3979
rect 31247 3959 31252 3979
rect 30481 3751 30582 3752
rect 30379 3738 30582 3751
rect 30379 3736 30522 3738
rect 30379 3733 30456 3736
rect 30379 3706 30382 3733
rect 30411 3709 30456 3733
rect 30485 3709 30522 3736
rect 30411 3706 30522 3709
rect 30379 3705 30522 3706
rect 30558 3705 30582 3738
rect 30379 3692 30582 3705
rect 28466 3610 28472 3633
rect 28496 3610 28502 3633
rect 29956 3627 29992 3636
rect 29901 3617 29998 3627
rect 28713 3615 29998 3617
rect 28466 3589 28502 3610
rect 28466 3566 28472 3589
rect 28496 3566 28502 3589
rect 28466 3413 28502 3566
rect 28678 3605 29998 3615
rect 28678 3567 28690 3605
rect 28715 3570 28734 3605
rect 28759 3570 29998 3605
rect 28715 3567 29998 3570
rect 28678 3564 29998 3567
rect 28678 3562 29995 3564
rect 28678 3559 28767 3562
rect 28694 3558 28766 3559
rect 30621 3549 30691 3860
rect 30773 3673 30807 3951
rect 31220 3931 31252 3959
rect 30840 3923 31252 3931
rect 30840 3897 30846 3923
rect 30872 3897 31252 3923
rect 30840 3895 31252 3897
rect 30842 3894 30882 3895
rect 31009 3869 31040 3877
rect 31009 3839 31013 3869
rect 31034 3839 31040 3869
rect 30773 3665 30808 3673
rect 30773 3645 30781 3665
rect 30801 3645 30808 3665
rect 30773 3640 30808 3645
rect 31009 3640 31040 3839
rect 31220 3830 31252 3895
rect 31220 3810 31224 3830
rect 31245 3810 31252 3830
rect 31220 3803 31252 3810
rect 31665 3956 31737 3974
rect 31665 3914 31678 3956
rect 31727 3914 31737 3956
rect 31665 3893 31737 3914
rect 31665 3851 31679 3893
rect 31728 3851 31737 3893
rect 31529 3747 31630 3748
rect 31427 3734 31630 3747
rect 31427 3732 31570 3734
rect 31427 3729 31504 3732
rect 31427 3702 31430 3729
rect 31459 3705 31504 3729
rect 31533 3705 31570 3732
rect 31459 3702 31570 3705
rect 31427 3701 31570 3702
rect 31606 3701 31630 3734
rect 31427 3688 31630 3701
rect 30773 3639 30805 3640
rect 31007 3637 31040 3640
rect 30973 3618 31041 3637
rect 30943 3606 31042 3618
rect 31665 3610 31737 3851
rect 32109 3610 32216 4039
rect 32671 4451 32778 5044
rect 33146 4993 33221 5044
rect 34187 5095 34209 5109
rect 34253 5095 34270 5132
rect 34187 5075 34270 5095
rect 34187 5009 34204 5075
rect 34258 5009 34270 5075
rect 33146 4950 33222 4993
rect 33150 4639 33222 4950
rect 34187 4985 34270 5009
rect 34187 4965 34263 4985
rect 34187 4946 34266 4965
rect 33846 4930 33918 4931
rect 33845 4922 33944 4930
rect 33845 4919 33897 4922
rect 33845 4884 33853 4919
rect 33878 4884 33897 4919
rect 33922 4884 33944 4922
rect 33845 4872 33944 4884
rect 33846 4853 33914 4872
rect 33847 4850 33880 4853
rect 34082 4850 34114 4851
rect 33257 4789 33460 4802
rect 33257 4756 33281 4789
rect 33317 4788 33460 4789
rect 33317 4785 33428 4788
rect 33317 4758 33354 4785
rect 33383 4761 33428 4785
rect 33457 4761 33460 4788
rect 33383 4758 33460 4761
rect 33317 4756 33460 4758
rect 33257 4743 33460 4756
rect 33257 4742 33358 4743
rect 33150 4597 33159 4639
rect 33208 4597 33222 4639
rect 33150 4576 33222 4597
rect 33150 4534 33160 4576
rect 33209 4534 33222 4576
rect 33150 4516 33222 4534
rect 33635 4680 33667 4687
rect 33635 4660 33642 4680
rect 33663 4660 33667 4680
rect 33635 4595 33667 4660
rect 33847 4651 33878 4850
rect 34079 4845 34114 4850
rect 34079 4825 34086 4845
rect 34106 4825 34114 4845
rect 34079 4817 34114 4825
rect 33847 4621 33853 4651
rect 33874 4621 33878 4651
rect 33847 4613 33878 4621
rect 34005 4595 34045 4596
rect 33635 4593 34047 4595
rect 33635 4567 34015 4593
rect 34041 4567 34047 4593
rect 33635 4559 34047 4567
rect 33635 4531 33667 4559
rect 34080 4539 34114 4817
rect 34196 4630 34266 4946
rect 36184 4931 36215 4932
rect 36184 4923 36229 4931
rect 35264 4900 35428 4907
rect 36184 4900 36194 4923
rect 34890 4885 36194 4900
rect 36219 4885 36229 4923
rect 37448 4926 37482 6166
rect 37448 4922 37678 4926
rect 37448 4896 37647 4922
rect 37672 4896 37678 4922
rect 37448 4888 37678 4896
rect 34890 4867 36229 4885
rect 34895 4854 34931 4867
rect 35264 4864 35428 4867
rect 34305 4785 34508 4798
rect 34305 4752 34329 4785
rect 34365 4784 34508 4785
rect 34365 4781 34476 4784
rect 34365 4754 34402 4781
rect 34431 4757 34476 4781
rect 34505 4757 34508 4784
rect 34431 4754 34508 4757
rect 34365 4752 34508 4754
rect 34305 4739 34508 4752
rect 34305 4738 34406 4739
rect 33635 4511 33640 4531
rect 33661 4511 33667 4531
rect 33635 4504 33667 4511
rect 34058 4534 34114 4539
rect 34058 4514 34065 4534
rect 34085 4514 34114 4534
rect 34191 4624 34266 4630
rect 34191 4591 34199 4624
rect 34252 4591 34266 4624
rect 34191 4566 34266 4591
rect 34191 4533 34204 4566
rect 34257 4533 34266 4566
rect 34191 4524 34266 4533
rect 34683 4676 34715 4683
rect 34683 4656 34690 4676
rect 34711 4656 34715 4676
rect 34683 4591 34715 4656
rect 34895 4647 34926 4854
rect 38032 4852 38064 4853
rect 35130 4846 35162 4847
rect 35127 4841 35162 4846
rect 35127 4821 35134 4841
rect 35154 4821 35162 4841
rect 35127 4813 35162 4821
rect 34895 4617 34901 4647
rect 34922 4617 34926 4647
rect 34895 4609 34926 4617
rect 35053 4591 35093 4592
rect 34683 4589 35095 4591
rect 34683 4563 35063 4589
rect 35089 4563 35095 4589
rect 34683 4555 35095 4563
rect 34683 4527 34715 4555
rect 35128 4535 35162 4813
rect 37207 4791 37410 4804
rect 37207 4758 37231 4791
rect 37267 4790 37410 4791
rect 37267 4787 37378 4790
rect 37267 4760 37304 4787
rect 37333 4763 37378 4787
rect 37407 4763 37410 4790
rect 37333 4760 37410 4763
rect 37267 4758 37410 4760
rect 37207 4745 37410 4758
rect 37207 4744 37308 4745
rect 34191 4519 34249 4524
rect 34058 4507 34114 4514
rect 34683 4507 34688 4527
rect 34709 4507 34715 4527
rect 34058 4506 34093 4507
rect 34683 4500 34715 4507
rect 35106 4530 35162 4535
rect 35106 4510 35113 4530
rect 35133 4510 35162 4530
rect 35106 4503 35162 4510
rect 37585 4682 37617 4689
rect 37585 4662 37592 4682
rect 37613 4662 37617 4682
rect 37585 4597 37617 4662
rect 37797 4653 37828 4850
rect 38029 4847 38064 4852
rect 38029 4827 38036 4847
rect 38056 4827 38064 4847
rect 38029 4819 38064 4827
rect 37797 4623 37803 4653
rect 37824 4623 37828 4653
rect 37797 4615 37828 4623
rect 37955 4597 37995 4598
rect 37585 4595 37997 4597
rect 37585 4569 37965 4595
rect 37991 4569 37997 4595
rect 37585 4561 37997 4569
rect 37585 4533 37617 4561
rect 37585 4513 37590 4533
rect 37611 4513 37617 4533
rect 37585 4506 37617 4513
rect 37787 4535 37835 4542
rect 38030 4541 38064 4819
rect 37787 4515 37794 4535
rect 37827 4515 37835 4535
rect 35106 4502 35141 4503
rect 33349 4451 33460 4455
rect 35132 4451 36702 4452
rect 32671 4447 36702 4451
rect 37027 4447 37445 4460
rect 32671 4435 37445 4447
rect 32671 4433 37307 4435
rect 32671 4413 33357 4433
rect 33376 4413 33434 4433
rect 33453 4429 37307 4433
rect 33453 4413 34405 4429
rect 32671 4409 34405 4413
rect 34424 4409 34482 4429
rect 34501 4415 37307 4429
rect 37326 4415 37384 4435
rect 37403 4415 37445 4435
rect 34501 4409 37445 4415
rect 32671 4395 37445 4409
rect 32671 3772 32778 4395
rect 34397 4392 34508 4395
rect 37027 4389 37445 4395
rect 33157 4346 33221 4350
rect 33153 4340 33221 4346
rect 33153 4307 33170 4340
rect 33210 4307 33221 4340
rect 33153 4295 33221 4307
rect 34204 4309 34269 4331
rect 33153 4293 33210 4295
rect 33157 3932 33208 4293
rect 34204 4270 34221 4309
rect 34266 4270 34269 4309
rect 33845 4225 33880 4227
rect 33845 4216 33949 4225
rect 33845 4215 33896 4216
rect 33845 4195 33848 4215
rect 33873 4196 33896 4215
rect 33928 4196 33949 4216
rect 33873 4195 33949 4196
rect 33845 4188 33949 4195
rect 33845 4176 33880 4188
rect 33257 4110 33460 4123
rect 33257 4077 33281 4110
rect 33317 4109 33460 4110
rect 33317 4106 33428 4109
rect 33317 4079 33354 4106
rect 33383 4082 33428 4106
rect 33457 4082 33460 4109
rect 33383 4079 33460 4082
rect 33317 4077 33460 4079
rect 33257 4064 33460 4077
rect 33257 4063 33358 4064
rect 33635 4001 33667 4008
rect 33635 3981 33642 4001
rect 33663 3981 33667 4001
rect 33146 3923 33211 3932
rect 33146 3886 33156 3923
rect 33196 3889 33211 3923
rect 33635 3916 33667 3981
rect 33847 3972 33878 4176
rect 34082 4171 34114 4172
rect 34079 4166 34114 4171
rect 34079 4146 34086 4166
rect 34106 4146 34114 4166
rect 34079 4138 34114 4146
rect 33847 3942 33853 3972
rect 33874 3942 33878 3972
rect 33847 3934 33878 3942
rect 34005 3916 34045 3917
rect 33635 3914 34047 3916
rect 33196 3886 33213 3889
rect 33146 3867 33213 3886
rect 33146 3846 33160 3867
rect 33196 3846 33213 3867
rect 33146 3839 33213 3846
rect 33635 3888 34015 3914
rect 34041 3888 34047 3914
rect 33635 3880 34047 3888
rect 33635 3852 33667 3880
rect 34080 3860 34114 4138
rect 34204 3970 34269 4270
rect 36341 4231 36378 4252
rect 36341 4194 36352 4231
rect 36369 4207 36378 4231
rect 36369 4194 36379 4207
rect 36341 4184 36379 4194
rect 36342 4180 36379 4184
rect 36342 4174 36375 4180
rect 35752 4105 35955 4118
rect 35752 4072 35776 4105
rect 35812 4104 35955 4105
rect 35812 4101 35923 4104
rect 35812 4074 35849 4101
rect 35878 4077 35923 4101
rect 35952 4077 35955 4104
rect 35878 4074 35955 4077
rect 35812 4072 35955 4074
rect 35752 4059 35955 4072
rect 35752 4058 35853 4059
rect 36130 3996 36162 4003
rect 36130 3976 36137 3996
rect 36158 3976 36162 3996
rect 33635 3832 33640 3852
rect 33661 3832 33667 3852
rect 33635 3825 33667 3832
rect 34058 3855 34114 3860
rect 34058 3835 34065 3855
rect 34085 3835 34114 3855
rect 34058 3828 34114 3835
rect 34194 3959 34274 3970
rect 34194 3933 34211 3959
rect 34251 3933 34274 3959
rect 34194 3906 34274 3933
rect 34194 3880 34215 3906
rect 34255 3880 34274 3906
rect 34194 3861 34274 3880
rect 34194 3835 34218 3861
rect 34258 3835 34274 3861
rect 35268 3905 35373 3926
rect 36130 3911 36162 3976
rect 36342 3967 36373 4174
rect 36577 4166 36609 4167
rect 36574 4161 36609 4166
rect 36574 4141 36581 4161
rect 36601 4141 36609 4161
rect 36574 4133 36609 4141
rect 36342 3937 36348 3967
rect 36369 3937 36373 3967
rect 36342 3929 36373 3937
rect 36500 3911 36540 3912
rect 36130 3909 36542 3911
rect 35268 3899 35744 3905
rect 35268 3897 35325 3899
rect 35268 3866 35280 3897
rect 35305 3876 35325 3897
rect 35351 3892 35744 3899
rect 35351 3876 35705 3892
rect 35305 3869 35705 3876
rect 35731 3869 35744 3892
rect 35305 3866 35744 3869
rect 35268 3856 35744 3866
rect 36130 3883 36510 3909
rect 36536 3883 36542 3909
rect 36130 3875 36542 3883
rect 35268 3854 35373 3856
rect 34058 3827 34093 3828
rect 34194 3823 34274 3835
rect 36130 3847 36162 3875
rect 36575 3855 36609 4133
rect 36130 3827 36135 3847
rect 36156 3827 36162 3847
rect 36130 3820 36162 3827
rect 36553 3850 36609 3855
rect 36553 3830 36560 3850
rect 36580 3830 36609 3850
rect 36553 3823 36609 3830
rect 36553 3822 36588 3823
rect 33349 3772 33460 3776
rect 35091 3772 36744 3775
rect 32669 3754 36744 3772
rect 32669 3734 33357 3754
rect 33376 3734 33434 3754
rect 33453 3749 36744 3754
rect 33453 3734 35852 3749
rect 32669 3729 35852 3734
rect 35871 3729 35929 3749
rect 35948 3729 36744 3749
rect 32669 3719 36744 3729
rect 32669 3716 33294 3719
rect 33481 3716 36744 3719
rect 30943 3568 30965 3606
rect 30990 3571 31009 3606
rect 31034 3571 31042 3606
rect 30990 3568 31042 3571
rect 30943 3560 31042 3568
rect 30969 3559 31041 3560
rect 30620 3533 30691 3549
rect 30620 3517 30640 3533
rect 30621 3487 30640 3517
rect 30623 3467 30640 3487
rect 30670 3487 30691 3533
rect 31663 3529 31741 3610
rect 32108 3555 32216 3610
rect 30670 3467 30690 3487
rect 30623 3448 30690 3467
rect 31663 3427 31742 3529
rect 28457 3404 28543 3413
rect 28457 3386 28476 3404
rect 28528 3386 28543 3404
rect 28457 3382 28543 3386
rect 31627 3409 31748 3427
rect 31627 3407 31698 3409
rect 31627 3366 31642 3407
rect 31679 3368 31698 3407
rect 31735 3368 31748 3409
rect 31679 3366 31748 3368
rect 31627 3356 31748 3366
rect 28932 3328 29043 3331
rect 28247 3327 29796 3328
rect 32109 3327 32216 3555
rect 32671 3488 32778 3716
rect 35091 3715 36744 3716
rect 35844 3712 35955 3715
rect 33139 3677 33260 3687
rect 33139 3675 33208 3677
rect 33139 3634 33152 3675
rect 33189 3636 33208 3675
rect 33245 3636 33260 3677
rect 33189 3634 33260 3636
rect 33139 3616 33260 3634
rect 33145 3514 33224 3616
rect 34197 3576 34264 3595
rect 34197 3556 34217 3576
rect 32671 3433 32779 3488
rect 33146 3433 33224 3514
rect 34196 3510 34217 3556
rect 34247 3556 34264 3576
rect 34247 3526 34266 3556
rect 34247 3510 34267 3526
rect 34196 3494 34267 3510
rect 33846 3483 33918 3484
rect 33845 3475 33944 3483
rect 33845 3472 33897 3475
rect 33845 3437 33853 3472
rect 33878 3437 33897 3472
rect 33922 3437 33944 3475
rect 28247 3324 31406 3327
rect 31593 3324 32218 3327
rect 28247 3314 32218 3324
rect 28247 3294 28939 3314
rect 28958 3294 29016 3314
rect 29035 3309 32218 3314
rect 29035 3294 31434 3309
rect 28247 3289 31434 3294
rect 31453 3289 31511 3309
rect 31530 3289 32218 3309
rect 28247 3271 32218 3289
rect 28247 3268 29796 3271
rect 31427 3267 31538 3271
rect 28299 3220 28334 3221
rect 28278 3213 28334 3220
rect 28278 3193 28307 3213
rect 28327 3193 28334 3213
rect 28278 3188 28334 3193
rect 28725 3216 28757 3223
rect 28725 3196 28731 3216
rect 28752 3196 28757 3216
rect 28278 2910 28312 3188
rect 28725 3168 28757 3196
rect 28345 3160 28757 3168
rect 28345 3134 28351 3160
rect 28377 3134 28757 3160
rect 28345 3132 28757 3134
rect 28347 3131 28387 3132
rect 28514 3106 28545 3114
rect 28514 3076 28518 3106
rect 28539 3076 28545 3106
rect 28278 2902 28313 2910
rect 28278 2882 28286 2902
rect 28306 2882 28313 2902
rect 28278 2877 28313 2882
rect 28278 2876 28310 2877
rect 28514 2875 28545 3076
rect 28725 3067 28757 3132
rect 28725 3047 28729 3067
rect 28750 3047 28757 3067
rect 28725 3040 28757 3047
rect 29319 3207 29412 3214
rect 29319 3166 29343 3207
rect 29397 3166 29412 3207
rect 29034 2984 29135 2985
rect 28932 2971 29135 2984
rect 28932 2969 29075 2971
rect 28932 2966 29009 2969
rect 28932 2939 28935 2966
rect 28964 2942 29009 2966
rect 29038 2942 29075 2969
rect 28964 2939 29075 2942
rect 28932 2938 29075 2939
rect 29111 2938 29135 2971
rect 28932 2925 29135 2938
rect 29319 2793 29412 3166
rect 30613 3208 30693 3220
rect 30794 3215 30829 3216
rect 30613 3182 30629 3208
rect 30669 3182 30693 3208
rect 30613 3163 30693 3182
rect 30613 3137 30632 3163
rect 30672 3137 30693 3163
rect 30613 3110 30693 3137
rect 30613 3084 30636 3110
rect 30676 3084 30693 3110
rect 30613 3073 30693 3084
rect 30773 3208 30829 3215
rect 30773 3188 30802 3208
rect 30822 3188 30829 3208
rect 30773 3183 30829 3188
rect 31220 3211 31252 3218
rect 31220 3191 31226 3211
rect 31247 3191 31252 3211
rect 29319 2749 29337 2793
rect 29397 2749 29412 2793
rect 29319 2734 29412 2749
rect 30618 2773 30683 3073
rect 30773 2905 30807 3183
rect 31220 3163 31252 3191
rect 30840 3155 31252 3163
rect 30840 3129 30846 3155
rect 30872 3129 31252 3155
rect 31674 3197 31741 3204
rect 31674 3176 31691 3197
rect 31727 3176 31741 3197
rect 31674 3157 31741 3176
rect 31674 3154 31691 3157
rect 30840 3127 31252 3129
rect 30842 3126 30882 3127
rect 31009 3101 31040 3109
rect 31009 3071 31013 3101
rect 31034 3071 31040 3101
rect 30773 2897 30808 2905
rect 30773 2877 30781 2897
rect 30801 2877 30808 2897
rect 30773 2872 30808 2877
rect 30773 2871 30805 2872
rect 31009 2867 31040 3071
rect 31220 3062 31252 3127
rect 31676 3120 31691 3154
rect 31731 3120 31741 3157
rect 31676 3111 31741 3120
rect 31220 3042 31224 3062
rect 31245 3042 31252 3062
rect 31220 3035 31252 3042
rect 31529 2979 31630 2980
rect 31427 2966 31630 2979
rect 31427 2964 31570 2966
rect 31427 2961 31504 2964
rect 31427 2934 31430 2961
rect 31459 2937 31504 2961
rect 31533 2937 31570 2964
rect 31459 2934 31570 2937
rect 31427 2933 31570 2934
rect 31606 2933 31630 2966
rect 31427 2920 31630 2933
rect 31007 2855 31042 2867
rect 30938 2848 31042 2855
rect 30938 2847 31014 2848
rect 30938 2827 30959 2847
rect 30991 2828 31014 2847
rect 31039 2828 31042 2848
rect 30991 2827 31042 2828
rect 30938 2818 31042 2827
rect 31007 2816 31042 2818
rect 30618 2734 30621 2773
rect 30666 2734 30683 2773
rect 31679 2750 31730 3111
rect 31677 2748 31734 2750
rect 30618 2712 30683 2734
rect 31666 2736 31734 2748
rect 31666 2703 31677 2736
rect 31717 2703 31734 2736
rect 31666 2697 31734 2703
rect 31666 2693 31730 2697
rect 30379 2648 30490 2651
rect 32109 2648 32216 3271
rect 28642 2634 32216 2648
rect 28642 2614 30386 2634
rect 30405 2614 30463 2634
rect 30482 2630 32216 2634
rect 30482 2614 31434 2630
rect 28642 2610 31434 2614
rect 31453 2610 31511 2630
rect 31530 2610 32216 2630
rect 28642 2592 32216 2610
rect 28642 2591 29755 2592
rect 31427 2588 31538 2592
rect 29746 2540 29781 2541
rect 29725 2533 29781 2540
rect 29725 2513 29754 2533
rect 29774 2513 29781 2533
rect 29725 2508 29781 2513
rect 30172 2536 30204 2543
rect 30794 2536 30829 2537
rect 30172 2516 30178 2536
rect 30199 2516 30204 2536
rect 30773 2529 30829 2536
rect 30638 2519 30696 2524
rect 27561 2473 29414 2506
rect 27561 2408 27626 2473
rect 27757 2453 29414 2473
rect 27757 2412 29350 2453
rect 29386 2412 29414 2453
rect 29512 2473 29576 2492
rect 29512 2434 29529 2473
rect 29563 2434 29576 2473
rect 29512 2415 29576 2434
rect 27757 2408 29414 2412
rect 27561 2383 29414 2408
rect 29325 2380 29407 2383
rect 29514 1903 29576 2415
rect 29725 2230 29759 2508
rect 30172 2488 30204 2516
rect 29792 2480 30204 2488
rect 29792 2454 29798 2480
rect 29824 2454 30204 2480
rect 29792 2452 30204 2454
rect 29794 2451 29834 2452
rect 29961 2426 29992 2434
rect 29961 2396 29965 2426
rect 29986 2396 29992 2426
rect 29725 2222 29760 2230
rect 29725 2202 29733 2222
rect 29753 2202 29760 2222
rect 29725 2197 29760 2202
rect 29725 2196 29757 2197
rect 29961 2189 29992 2396
rect 30172 2387 30204 2452
rect 30172 2367 30176 2387
rect 30197 2367 30204 2387
rect 30172 2360 30204 2367
rect 30621 2510 30696 2519
rect 30621 2477 30630 2510
rect 30683 2477 30696 2510
rect 30621 2452 30696 2477
rect 30621 2419 30635 2452
rect 30688 2419 30696 2452
rect 30621 2413 30696 2419
rect 30773 2509 30802 2529
rect 30822 2509 30829 2529
rect 30773 2504 30829 2509
rect 31220 2532 31252 2539
rect 31220 2512 31226 2532
rect 31247 2512 31252 2532
rect 30481 2304 30582 2305
rect 30379 2291 30582 2304
rect 30379 2289 30522 2291
rect 30379 2286 30456 2289
rect 30379 2259 30382 2286
rect 30411 2262 30456 2286
rect 30485 2262 30522 2289
rect 30411 2259 30522 2262
rect 30379 2258 30522 2259
rect 30558 2258 30582 2291
rect 30379 2245 30582 2258
rect 29956 2171 29992 2189
rect 29923 2170 29992 2171
rect 29903 2158 29992 2170
rect 29903 2120 29915 2158
rect 29940 2123 29959 2158
rect 29984 2123 29992 2158
rect 29940 2120 29992 2123
rect 29903 2112 29992 2120
rect 29919 2111 29991 2112
rect 29472 1845 29588 1903
rect 30621 1892 30691 2413
rect 30773 2226 30807 2504
rect 31220 2484 31252 2512
rect 30840 2476 31252 2484
rect 30840 2450 30846 2476
rect 30872 2450 31252 2476
rect 30840 2448 31252 2450
rect 30842 2447 30882 2448
rect 31009 2422 31040 2430
rect 31009 2392 31013 2422
rect 31034 2392 31040 2422
rect 30773 2218 30808 2226
rect 30773 2198 30781 2218
rect 30801 2198 30808 2218
rect 30773 2193 30808 2198
rect 31009 2193 31040 2392
rect 31220 2383 31252 2448
rect 31220 2363 31224 2383
rect 31245 2363 31252 2383
rect 31220 2356 31252 2363
rect 31665 2509 31737 2527
rect 31665 2467 31678 2509
rect 31727 2467 31737 2509
rect 31665 2446 31737 2467
rect 31665 2404 31679 2446
rect 31728 2404 31737 2446
rect 31529 2300 31630 2301
rect 31427 2287 31630 2300
rect 31427 2285 31570 2287
rect 31427 2282 31504 2285
rect 31427 2255 31430 2282
rect 31459 2258 31504 2282
rect 31533 2258 31570 2285
rect 31459 2255 31570 2258
rect 31427 2254 31570 2255
rect 31606 2254 31630 2287
rect 31427 2241 31630 2254
rect 30773 2192 30805 2193
rect 31007 2190 31040 2193
rect 30973 2171 31041 2190
rect 30943 2159 31042 2171
rect 30943 2121 30965 2159
rect 30990 2124 31009 2159
rect 31034 2124 31042 2159
rect 30990 2121 31042 2124
rect 30943 2113 31042 2121
rect 30969 2112 31041 2113
rect 29472 1774 29484 1845
rect 29563 1774 29588 1845
rect 29472 1754 29588 1774
rect 30602 1691 30704 1892
rect 31665 1884 31737 2404
rect 32109 1980 32216 2592
rect 32671 3004 32778 3433
rect 33150 3192 33222 3433
rect 33845 3425 33944 3437
rect 33846 3406 33914 3425
rect 33847 3403 33880 3406
rect 34082 3403 34114 3404
rect 33257 3342 33460 3355
rect 33257 3309 33281 3342
rect 33317 3341 33460 3342
rect 33317 3338 33428 3341
rect 33317 3311 33354 3338
rect 33383 3314 33428 3338
rect 33457 3314 33460 3341
rect 33383 3311 33460 3314
rect 33317 3309 33460 3311
rect 33257 3296 33460 3309
rect 33257 3295 33358 3296
rect 33150 3150 33159 3192
rect 33208 3150 33222 3192
rect 33150 3129 33222 3150
rect 33150 3087 33160 3129
rect 33209 3087 33222 3129
rect 33150 3069 33222 3087
rect 33635 3233 33667 3240
rect 33635 3213 33642 3233
rect 33663 3213 33667 3233
rect 33635 3148 33667 3213
rect 33847 3204 33878 3403
rect 34079 3398 34114 3403
rect 34079 3378 34086 3398
rect 34106 3378 34114 3398
rect 34079 3370 34114 3378
rect 33847 3174 33853 3204
rect 33874 3174 33878 3204
rect 33847 3166 33878 3174
rect 34005 3148 34045 3149
rect 33635 3146 34047 3148
rect 33635 3120 34015 3146
rect 34041 3120 34047 3146
rect 33635 3112 34047 3120
rect 33635 3084 33667 3112
rect 34080 3092 34114 3370
rect 34196 3183 34266 3494
rect 34893 3485 36235 3490
rect 34893 3483 36192 3485
rect 34890 3457 36192 3483
rect 36220 3457 36235 3485
rect 34890 3449 36235 3457
rect 34890 3424 34929 3449
rect 34890 3407 34931 3424
rect 34890 3400 34929 3407
rect 34305 3338 34508 3351
rect 34305 3305 34329 3338
rect 34365 3337 34508 3338
rect 34365 3334 34476 3337
rect 34365 3307 34402 3334
rect 34431 3310 34476 3334
rect 34505 3310 34508 3337
rect 34431 3307 34508 3310
rect 34365 3305 34508 3307
rect 34305 3292 34508 3305
rect 34305 3291 34406 3292
rect 33635 3064 33640 3084
rect 33661 3064 33667 3084
rect 33635 3057 33667 3064
rect 34058 3087 34114 3092
rect 34058 3067 34065 3087
rect 34085 3067 34114 3087
rect 34191 3177 34266 3183
rect 34191 3144 34199 3177
rect 34252 3144 34266 3177
rect 34191 3119 34266 3144
rect 34191 3086 34204 3119
rect 34257 3086 34266 3119
rect 34191 3077 34266 3086
rect 34683 3229 34715 3236
rect 34683 3209 34690 3229
rect 34711 3209 34715 3229
rect 34683 3144 34715 3209
rect 34895 3200 34926 3400
rect 35130 3399 35162 3400
rect 35127 3394 35162 3399
rect 35127 3374 35134 3394
rect 35154 3374 35162 3394
rect 35127 3366 35162 3374
rect 34895 3170 34901 3200
rect 34922 3170 34926 3200
rect 34895 3162 34926 3170
rect 35053 3144 35093 3145
rect 34683 3142 35095 3144
rect 34683 3116 35063 3142
rect 35089 3116 35095 3142
rect 34683 3108 35095 3116
rect 34683 3080 34715 3108
rect 35128 3088 35162 3366
rect 34191 3072 34249 3077
rect 34058 3060 34114 3067
rect 34683 3060 34688 3080
rect 34709 3060 34715 3080
rect 34058 3059 34093 3060
rect 34683 3053 34715 3060
rect 35106 3083 35162 3088
rect 35106 3063 35113 3083
rect 35133 3063 35162 3083
rect 35106 3056 35162 3063
rect 35106 3055 35141 3056
rect 33349 3004 33460 3008
rect 35224 3004 35655 3005
rect 32671 2986 35655 3004
rect 32671 2966 33357 2986
rect 33376 2966 33434 2986
rect 33453 2982 35655 2986
rect 33453 2966 34405 2982
rect 32671 2962 34405 2966
rect 34424 2962 34482 2982
rect 34501 2962 35655 2982
rect 32671 2948 35655 2962
rect 32671 2325 32778 2948
rect 34397 2945 34508 2948
rect 33157 2899 33221 2903
rect 33153 2893 33221 2899
rect 33153 2860 33170 2893
rect 33210 2860 33221 2893
rect 33153 2848 33221 2860
rect 34204 2862 34269 2884
rect 33153 2846 33210 2848
rect 33157 2485 33208 2846
rect 34204 2823 34221 2862
rect 34266 2823 34269 2862
rect 33845 2778 33880 2780
rect 33845 2769 33949 2778
rect 33845 2768 33896 2769
rect 33845 2748 33848 2768
rect 33873 2749 33896 2768
rect 33928 2749 33949 2769
rect 33873 2748 33949 2749
rect 33845 2741 33949 2748
rect 33845 2729 33880 2741
rect 33257 2663 33460 2676
rect 33257 2630 33281 2663
rect 33317 2662 33460 2663
rect 33317 2659 33428 2662
rect 33317 2632 33354 2659
rect 33383 2635 33428 2659
rect 33457 2635 33460 2662
rect 33383 2632 33460 2635
rect 33317 2630 33460 2632
rect 33257 2617 33460 2630
rect 33257 2616 33358 2617
rect 33635 2554 33667 2561
rect 33635 2534 33642 2554
rect 33663 2534 33667 2554
rect 33146 2476 33211 2485
rect 33146 2439 33156 2476
rect 33196 2442 33211 2476
rect 33635 2469 33667 2534
rect 33847 2525 33878 2729
rect 34082 2724 34114 2725
rect 34079 2719 34114 2724
rect 34079 2699 34086 2719
rect 34106 2699 34114 2719
rect 34079 2691 34114 2699
rect 33847 2495 33853 2525
rect 33874 2495 33878 2525
rect 33847 2487 33878 2495
rect 34005 2469 34045 2470
rect 33635 2467 34047 2469
rect 33196 2439 33213 2442
rect 33146 2420 33213 2439
rect 33146 2399 33160 2420
rect 33196 2399 33213 2420
rect 33146 2392 33213 2399
rect 33635 2441 34015 2467
rect 34041 2441 34047 2467
rect 33635 2433 34047 2441
rect 33635 2405 33667 2433
rect 34080 2413 34114 2691
rect 34204 2560 34269 2823
rect 34204 2556 34265 2560
rect 33635 2385 33640 2405
rect 33661 2385 33667 2405
rect 33635 2378 33667 2385
rect 34058 2408 34114 2413
rect 34058 2388 34065 2408
rect 34085 2388 34114 2408
rect 34058 2381 34114 2388
rect 34058 2380 34093 2381
rect 33349 2325 33460 2329
rect 32669 2307 33988 2325
rect 32669 2287 33357 2307
rect 33376 2287 33434 2307
rect 33453 2287 33988 2307
rect 32669 2269 33988 2287
rect 32671 2149 32778 2269
rect 33139 2230 33260 2240
rect 33139 2228 33208 2230
rect 33139 2187 33152 2228
rect 33189 2189 33208 2228
rect 33245 2189 33260 2230
rect 33189 2187 33260 2189
rect 33139 2169 33260 2187
rect 32108 1944 32216 1980
rect 32263 2103 32417 2128
rect 32263 1991 32276 2103
rect 32397 1991 32417 2103
rect 30566 1654 30732 1691
rect 30566 1575 30603 1654
rect 30687 1575 30732 1654
rect 30566 1537 30732 1575
rect 31643 1483 31740 1884
rect 32101 1808 32221 1944
rect 32108 1802 32216 1808
rect 31573 1454 31748 1483
rect 31573 1375 31619 1454
rect 31719 1375 31748 1454
rect 31573 1350 31748 1375
rect 32108 1259 32212 1802
rect 31951 1229 32222 1259
rect 31951 1142 31985 1229
rect 32055 1221 32222 1229
rect 32055 1142 32118 1221
rect 31951 1134 32118 1142
rect 32188 1134 32222 1221
rect 31951 1088 32222 1134
rect 27075 773 31984 791
rect 22320 733 22528 745
rect 26679 733 26790 743
rect 22287 718 26790 733
rect 22287 662 22334 718
rect 22413 708 26790 718
rect 27075 727 31886 773
rect 31962 727 31984 773
rect 27075 716 31984 727
rect 22413 662 22464 708
rect 22287 657 22464 662
rect 22510 657 26790 708
rect 22287 636 26790 657
rect 22417 630 22519 636
rect 21224 499 21427 512
rect 21224 466 21248 499
rect 21284 498 21427 499
rect 21284 495 21395 498
rect 21284 468 21321 495
rect 21350 471 21395 495
rect 21424 471 21427 498
rect 21350 468 21427 471
rect 21284 466 21427 468
rect 21224 453 21427 466
rect 21224 452 21325 453
rect 21602 390 21634 397
rect 21602 370 21609 390
rect 21630 370 21634 390
rect 21602 305 21634 370
rect 21814 361 21845 587
rect 22049 560 22081 561
rect 22046 555 22081 560
rect 22046 535 22053 555
rect 22073 535 22081 555
rect 22046 527 22081 535
rect 21814 331 21820 361
rect 21841 331 21845 361
rect 21814 323 21845 331
rect 21972 305 22012 306
rect 21602 303 22014 305
rect 21602 277 21982 303
rect 22008 277 22014 303
rect 21602 269 22014 277
rect 21602 241 21634 269
rect 21602 221 21607 241
rect 21628 221 21634 241
rect 21602 214 21634 221
rect 21816 243 21847 253
rect 22047 249 22081 527
rect 26679 327 26790 636
rect 31836 331 31965 338
rect 31836 327 31860 331
rect 26675 272 31860 327
rect 31891 272 31922 331
rect 31953 272 31965 331
rect 26675 263 31965 272
rect 26679 257 26790 263
rect 31836 259 31965 263
rect 21816 221 21823 243
rect 21841 221 21847 243
rect 21316 154 21427 165
rect 20955 143 21427 154
rect 20955 123 21324 143
rect 21343 123 21401 143
rect 21420 123 21427 143
rect 20955 111 21427 123
rect 20955 109 21054 111
rect 21316 106 21427 111
rect 19378 3 20571 13
rect 19167 -16 20571 3
rect 19167 -98 19210 -16
rect 19368 -83 20571 -16
rect 19368 -98 19411 -83
rect 19167 -117 19411 -98
rect 21816 -170 21847 221
rect 22025 244 22081 249
rect 22025 224 22032 244
rect 22052 224 22081 244
rect 22025 217 22081 224
rect 22025 216 22060 217
rect 32056 155 32128 1088
rect 32263 1017 32417 1991
rect 32261 1001 32417 1017
rect 32470 2076 32604 2105
rect 32470 1964 32508 2076
rect 32587 1964 32604 2076
rect 32671 2069 32779 2149
rect 32470 1011 32604 1964
rect 32672 1257 32779 2069
rect 33145 2097 33210 2169
rect 33145 2031 33213 2097
rect 33146 1485 33213 2031
rect 34200 1669 34265 2556
rect 35243 2286 35380 2290
rect 35230 2282 35387 2286
rect 35230 2175 35267 2282
rect 35367 2175 35387 2282
rect 35230 2133 35387 2175
rect 35243 1885 35380 2133
rect 35233 1843 35399 1885
rect 35233 1768 35262 1843
rect 35379 1768 35399 1843
rect 35233 1752 35399 1768
rect 34189 1648 34326 1669
rect 34189 1573 34214 1648
rect 34284 1573 34326 1648
rect 34189 1542 34326 1573
rect 33132 1436 33307 1485
rect 33132 1357 33165 1436
rect 33265 1357 33307 1436
rect 33132 1352 33307 1357
rect 32672 1215 32820 1257
rect 32672 1207 32712 1215
rect 32674 1128 32712 1207
rect 32782 1128 32820 1215
rect 32674 1090 32820 1128
rect 32261 976 32413 1001
rect 32261 881 32291 976
rect 32381 881 32413 976
rect 32261 868 32413 881
rect 32466 975 32605 1011
rect 32466 880 32480 975
rect 32570 880 32605 975
rect 32466 862 32605 880
rect 37787 795 37835 4515
rect 38008 4536 38064 4541
rect 38008 4516 38015 4536
rect 38035 4516 38064 4536
rect 38008 4509 38064 4516
rect 38008 4508 38043 4509
rect 38112 4418 38140 7226
rect 41325 7181 41390 7481
rect 41480 7313 41514 7591
rect 41927 7571 41959 7599
rect 41547 7563 41959 7571
rect 41547 7537 41553 7563
rect 41579 7537 41959 7563
rect 42381 7605 42448 7612
rect 42381 7584 42398 7605
rect 42434 7584 42448 7605
rect 42381 7565 42448 7584
rect 42381 7562 42398 7565
rect 41547 7535 41959 7537
rect 41549 7534 41589 7535
rect 41716 7509 41747 7517
rect 41716 7479 41720 7509
rect 41741 7479 41747 7509
rect 41480 7305 41515 7313
rect 41480 7285 41488 7305
rect 41508 7285 41515 7305
rect 41480 7280 41515 7285
rect 41480 7279 41512 7280
rect 41716 7275 41747 7479
rect 41927 7470 41959 7535
rect 42383 7528 42398 7562
rect 42438 7528 42448 7565
rect 42383 7519 42448 7528
rect 41927 7450 41931 7470
rect 41952 7450 41959 7470
rect 41927 7443 41959 7450
rect 42236 7387 42337 7388
rect 42134 7374 42337 7387
rect 42134 7372 42277 7374
rect 42134 7369 42211 7372
rect 42134 7342 42137 7369
rect 42166 7345 42211 7369
rect 42240 7345 42277 7372
rect 42166 7342 42277 7345
rect 42134 7341 42277 7342
rect 42313 7341 42337 7374
rect 42134 7328 42337 7341
rect 41714 7263 41749 7275
rect 41645 7256 41749 7263
rect 41645 7255 41721 7256
rect 41645 7235 41666 7255
rect 41698 7236 41721 7255
rect 41746 7236 41749 7256
rect 41698 7235 41749 7236
rect 41645 7226 41749 7235
rect 41714 7224 41749 7226
rect 41325 7142 41328 7181
rect 41373 7142 41390 7181
rect 42386 7158 42437 7519
rect 42384 7156 42441 7158
rect 41325 7120 41390 7142
rect 42373 7144 42441 7156
rect 42373 7111 42384 7144
rect 42424 7111 42441 7144
rect 42373 7105 42441 7111
rect 42373 7101 42437 7105
rect 41086 7056 41197 7059
rect 42816 7056 42923 7679
rect 39877 7042 42923 7056
rect 39877 7022 41093 7042
rect 41112 7022 41170 7042
rect 41189 7038 42923 7042
rect 41189 7022 42141 7038
rect 39877 7018 42141 7022
rect 42160 7018 42218 7038
rect 42237 7018 42923 7038
rect 39877 7000 42923 7018
rect 39877 6999 40370 7000
rect 42134 6996 42245 7000
rect 40453 6948 40488 6949
rect 40432 6941 40488 6948
rect 40432 6921 40461 6941
rect 40481 6921 40488 6941
rect 40432 6916 40488 6921
rect 40879 6944 40911 6951
rect 41501 6944 41536 6945
rect 40879 6924 40885 6944
rect 40906 6924 40911 6944
rect 41480 6937 41536 6944
rect 41345 6927 41403 6932
rect 40432 6638 40466 6916
rect 40879 6896 40911 6924
rect 40499 6888 40911 6896
rect 40499 6862 40505 6888
rect 40531 6862 40911 6888
rect 40499 6860 40911 6862
rect 40501 6859 40541 6860
rect 40668 6834 40699 6842
rect 40668 6804 40672 6834
rect 40693 6804 40699 6834
rect 40432 6630 40467 6638
rect 40432 6610 40440 6630
rect 40460 6610 40467 6630
rect 40432 6605 40467 6610
rect 40432 6604 40464 6605
rect 40668 6604 40699 6804
rect 40879 6795 40911 6860
rect 40879 6775 40883 6795
rect 40904 6775 40911 6795
rect 40879 6768 40911 6775
rect 41328 6918 41403 6927
rect 41328 6885 41337 6918
rect 41390 6885 41403 6918
rect 41328 6860 41403 6885
rect 41328 6827 41342 6860
rect 41395 6827 41403 6860
rect 41328 6821 41403 6827
rect 41480 6917 41509 6937
rect 41529 6917 41536 6937
rect 41480 6912 41536 6917
rect 41927 6940 41959 6947
rect 41927 6920 41933 6940
rect 41954 6920 41959 6940
rect 41188 6712 41289 6713
rect 41086 6699 41289 6712
rect 41086 6697 41229 6699
rect 41086 6694 41163 6697
rect 41086 6667 41089 6694
rect 41118 6670 41163 6694
rect 41192 6670 41229 6697
rect 41118 6667 41229 6670
rect 41086 6666 41229 6667
rect 41265 6666 41289 6699
rect 41086 6653 41289 6666
rect 40665 6597 40704 6604
rect 40663 6580 40704 6597
rect 40665 6555 40704 6580
rect 39359 6547 40704 6555
rect 39359 6519 39374 6547
rect 39402 6521 40704 6547
rect 39402 6519 40701 6521
rect 39359 6514 40701 6519
rect 41328 6510 41398 6821
rect 41480 6634 41514 6912
rect 41927 6892 41959 6920
rect 41547 6884 41959 6892
rect 41547 6858 41553 6884
rect 41579 6858 41959 6884
rect 41547 6856 41959 6858
rect 41549 6855 41589 6856
rect 41716 6830 41747 6838
rect 41716 6800 41720 6830
rect 41741 6800 41747 6830
rect 41480 6626 41515 6634
rect 41480 6606 41488 6626
rect 41508 6606 41515 6626
rect 41480 6601 41515 6606
rect 41716 6601 41747 6800
rect 41927 6791 41959 6856
rect 41927 6771 41931 6791
rect 41952 6771 41959 6791
rect 41927 6764 41959 6771
rect 42372 6917 42444 6935
rect 42372 6875 42385 6917
rect 42434 6875 42444 6917
rect 42372 6854 42444 6875
rect 42372 6812 42386 6854
rect 42435 6812 42444 6854
rect 42236 6708 42337 6709
rect 42134 6695 42337 6708
rect 42134 6693 42277 6695
rect 42134 6690 42211 6693
rect 42134 6663 42137 6690
rect 42166 6666 42211 6690
rect 42240 6666 42277 6693
rect 42166 6663 42277 6666
rect 42134 6662 42277 6663
rect 42313 6662 42337 6695
rect 42134 6649 42337 6662
rect 41480 6600 41512 6601
rect 41714 6598 41747 6601
rect 41680 6579 41748 6598
rect 41650 6567 41749 6579
rect 42372 6571 42444 6812
rect 42816 6571 42923 7000
rect 41650 6529 41672 6567
rect 41697 6532 41716 6567
rect 41741 6532 41749 6567
rect 41697 6529 41749 6532
rect 41650 6521 41749 6529
rect 41676 6520 41748 6521
rect 41327 6494 41398 6510
rect 41327 6478 41347 6494
rect 41328 6448 41347 6478
rect 41330 6428 41347 6448
rect 41377 6448 41398 6494
rect 42370 6490 42448 6571
rect 42815 6516 42923 6571
rect 41377 6428 41397 6448
rect 41330 6409 41397 6428
rect 42370 6388 42449 6490
rect 42334 6370 42455 6388
rect 42334 6368 42405 6370
rect 42334 6327 42349 6368
rect 42386 6329 42405 6368
rect 42442 6329 42455 6370
rect 42386 6327 42455 6329
rect 42334 6317 42455 6327
rect 39639 6289 39750 6292
rect 38953 6288 40503 6289
rect 42816 6288 42923 6516
rect 38953 6285 42113 6288
rect 42300 6285 42925 6288
rect 38953 6275 42925 6285
rect 38953 6255 39646 6275
rect 39665 6255 39723 6275
rect 39742 6270 42925 6275
rect 39742 6255 42141 6270
rect 38953 6250 42141 6255
rect 42160 6250 42218 6270
rect 42237 6250 42925 6270
rect 38953 6232 42925 6250
rect 38953 6229 40503 6232
rect 42134 6228 42245 6232
rect 39006 6181 39041 6182
rect 38985 6174 39041 6181
rect 38985 6154 39014 6174
rect 39034 6154 39041 6174
rect 38985 6149 39041 6154
rect 39432 6177 39464 6184
rect 39432 6157 39438 6177
rect 39459 6157 39464 6177
rect 38985 5871 39019 6149
rect 39432 6129 39464 6157
rect 41320 6169 41400 6181
rect 41501 6176 41536 6177
rect 39052 6121 39464 6129
rect 39052 6095 39058 6121
rect 39084 6095 39464 6121
rect 39850 6135 40287 6148
rect 39850 6112 39863 6135
rect 39889 6128 40287 6135
rect 39889 6112 40243 6128
rect 39850 6105 40243 6112
rect 40269 6105 40287 6128
rect 39850 6099 40287 6105
rect 41320 6143 41336 6169
rect 41376 6143 41400 6169
rect 41320 6124 41400 6143
rect 39052 6093 39464 6095
rect 39054 6092 39094 6093
rect 39221 6067 39252 6075
rect 39221 6037 39225 6067
rect 39246 6037 39252 6067
rect 38985 5863 39020 5871
rect 38985 5843 38993 5863
rect 39013 5843 39020 5863
rect 38985 5838 39020 5843
rect 38985 5837 39017 5838
rect 39221 5830 39252 6037
rect 39432 6028 39464 6093
rect 41320 6098 41339 6124
rect 41379 6098 41400 6124
rect 41320 6071 41400 6098
rect 41320 6045 41343 6071
rect 41383 6045 41400 6071
rect 41320 6034 41400 6045
rect 41480 6169 41536 6176
rect 41480 6149 41509 6169
rect 41529 6149 41536 6169
rect 41480 6144 41536 6149
rect 41927 6172 41959 6179
rect 41927 6152 41933 6172
rect 41954 6152 41959 6172
rect 39432 6008 39436 6028
rect 39457 6008 39464 6028
rect 39432 6001 39464 6008
rect 39741 5945 39842 5946
rect 39639 5932 39842 5945
rect 39639 5930 39782 5932
rect 39639 5927 39716 5930
rect 39639 5900 39642 5927
rect 39671 5903 39716 5927
rect 39745 5903 39782 5930
rect 39671 5900 39782 5903
rect 39639 5899 39782 5900
rect 39818 5899 39842 5932
rect 39639 5886 39842 5899
rect 39219 5824 39252 5830
rect 39215 5820 39252 5824
rect 39215 5810 39253 5820
rect 39215 5797 39225 5810
rect 39216 5773 39225 5797
rect 39242 5773 39253 5810
rect 39216 5752 39253 5773
rect 41325 5734 41390 6034
rect 41480 5866 41514 6144
rect 41927 6124 41959 6152
rect 41547 6116 41959 6124
rect 41547 6090 41553 6116
rect 41579 6090 41959 6116
rect 42381 6158 42448 6165
rect 42381 6137 42398 6158
rect 42434 6137 42448 6158
rect 42381 6118 42448 6137
rect 42381 6115 42398 6118
rect 41547 6088 41959 6090
rect 41549 6087 41589 6088
rect 41716 6062 41747 6070
rect 41716 6032 41720 6062
rect 41741 6032 41747 6062
rect 41480 5858 41515 5866
rect 41480 5838 41488 5858
rect 41508 5838 41515 5858
rect 41480 5833 41515 5838
rect 41480 5832 41512 5833
rect 41716 5828 41747 6032
rect 41927 6023 41959 6088
rect 42383 6081 42398 6115
rect 42438 6081 42448 6118
rect 42383 6072 42448 6081
rect 41927 6003 41931 6023
rect 41952 6003 41959 6023
rect 41927 5996 41959 6003
rect 42236 5940 42337 5941
rect 42134 5927 42337 5940
rect 42134 5925 42277 5927
rect 42134 5922 42211 5925
rect 42134 5895 42137 5922
rect 42166 5898 42211 5922
rect 42240 5898 42277 5925
rect 42166 5895 42277 5898
rect 42134 5894 42277 5895
rect 42313 5894 42337 5927
rect 42134 5881 42337 5894
rect 41714 5816 41749 5828
rect 41645 5809 41749 5816
rect 41645 5808 41721 5809
rect 41645 5788 41666 5808
rect 41698 5789 41721 5808
rect 41746 5789 41749 5809
rect 41698 5788 41749 5789
rect 41645 5779 41749 5788
rect 41714 5777 41749 5779
rect 41325 5695 41328 5734
rect 41373 5695 41390 5734
rect 42386 5711 42437 6072
rect 42384 5709 42441 5711
rect 41325 5673 41390 5695
rect 42373 5697 42441 5709
rect 42373 5664 42384 5697
rect 42424 5664 42441 5697
rect 42373 5658 42441 5664
rect 42373 5654 42437 5658
rect 41086 5609 41197 5612
rect 42816 5609 42923 6232
rect 39162 5595 42923 5609
rect 39162 5575 41093 5595
rect 41112 5575 41170 5595
rect 41189 5591 42923 5595
rect 41189 5575 42141 5591
rect 39162 5571 42141 5575
rect 42160 5571 42218 5591
rect 42237 5571 42923 5591
rect 39162 5553 42923 5571
rect 39162 5552 40462 5553
rect 42134 5549 42245 5553
rect 40453 5501 40488 5502
rect 40432 5494 40488 5501
rect 40432 5474 40461 5494
rect 40481 5474 40488 5494
rect 40432 5469 40488 5474
rect 40879 5497 40911 5504
rect 41501 5497 41536 5498
rect 40879 5477 40885 5497
rect 40906 5477 40911 5497
rect 41480 5490 41536 5497
rect 41345 5480 41403 5485
rect 40432 5191 40466 5469
rect 40879 5449 40911 5477
rect 40499 5441 40911 5449
rect 40499 5415 40505 5441
rect 40531 5415 40911 5441
rect 40499 5413 40911 5415
rect 40501 5412 40541 5413
rect 40668 5387 40699 5395
rect 40668 5357 40672 5387
rect 40693 5357 40699 5387
rect 40432 5183 40467 5191
rect 40432 5163 40440 5183
rect 40460 5163 40467 5183
rect 40432 5158 40467 5163
rect 40432 5157 40464 5158
rect 40668 5150 40699 5357
rect 40879 5348 40911 5413
rect 40879 5328 40883 5348
rect 40904 5328 40911 5348
rect 40879 5321 40911 5328
rect 41328 5471 41403 5480
rect 41328 5438 41337 5471
rect 41390 5438 41403 5471
rect 41328 5413 41403 5438
rect 41328 5380 41342 5413
rect 41395 5380 41403 5413
rect 41328 5374 41403 5380
rect 41480 5470 41509 5490
rect 41529 5470 41536 5490
rect 41480 5465 41536 5470
rect 41927 5493 41959 5500
rect 41927 5473 41933 5493
rect 41954 5473 41959 5493
rect 41188 5265 41289 5266
rect 41086 5252 41289 5265
rect 41086 5250 41229 5252
rect 41086 5247 41163 5250
rect 41086 5220 41089 5247
rect 41118 5223 41163 5247
rect 41192 5223 41229 5250
rect 41118 5220 41229 5223
rect 41086 5219 41229 5220
rect 41265 5219 41289 5252
rect 41086 5206 41289 5219
rect 40166 5137 40330 5140
rect 40663 5137 40699 5150
rect 39365 5119 40704 5137
rect 39365 5081 39375 5119
rect 39400 5104 40704 5119
rect 39400 5081 39410 5104
rect 40166 5097 40330 5104
rect 39365 5073 39410 5081
rect 39379 5072 39410 5073
rect 41328 5058 41398 5374
rect 41480 5187 41514 5465
rect 41927 5445 41959 5473
rect 41547 5437 41959 5445
rect 41547 5411 41553 5437
rect 41579 5411 41959 5437
rect 41547 5409 41959 5411
rect 41549 5408 41589 5409
rect 41716 5383 41747 5391
rect 41716 5353 41720 5383
rect 41741 5353 41747 5383
rect 41480 5179 41515 5187
rect 41480 5159 41488 5179
rect 41508 5159 41515 5179
rect 41480 5154 41515 5159
rect 41716 5154 41747 5353
rect 41927 5344 41959 5409
rect 41927 5324 41931 5344
rect 41952 5324 41959 5344
rect 41927 5317 41959 5324
rect 42372 5470 42444 5488
rect 42372 5428 42385 5470
rect 42434 5428 42444 5470
rect 42372 5407 42444 5428
rect 42372 5365 42386 5407
rect 42435 5365 42444 5407
rect 42236 5261 42337 5262
rect 42134 5248 42337 5261
rect 42134 5246 42277 5248
rect 42134 5243 42211 5246
rect 42134 5216 42137 5243
rect 42166 5219 42211 5243
rect 42240 5219 42277 5246
rect 42166 5216 42277 5219
rect 42134 5215 42277 5216
rect 42313 5215 42337 5248
rect 42134 5202 42337 5215
rect 41480 5153 41512 5154
rect 41714 5151 41747 5154
rect 41680 5132 41748 5151
rect 41650 5120 41749 5132
rect 41650 5082 41672 5120
rect 41697 5085 41716 5120
rect 41741 5085 41749 5120
rect 41697 5082 41749 5085
rect 41650 5074 41749 5082
rect 41676 5073 41748 5074
rect 41328 5039 41407 5058
rect 41331 5019 41407 5039
rect 41324 4995 41407 5019
rect 42372 5054 42444 5365
rect 42372 5011 42448 5054
rect 41324 4929 41336 4995
rect 41390 4929 41407 4995
rect 41324 4909 41407 4929
rect 41324 4872 41341 4909
rect 41385 4895 41407 4909
rect 42373 4960 42448 5011
rect 42816 4960 42923 5553
rect 41385 4872 41400 4895
rect 41324 4856 41400 4872
rect 42373 4868 42450 4960
rect 42816 4956 42924 4960
rect 42335 4850 42456 4868
rect 42335 4848 42406 4850
rect 42335 4807 42350 4848
rect 42387 4809 42406 4848
rect 42443 4809 42456 4850
rect 42387 4807 42456 4809
rect 42335 4797 42456 4807
rect 38906 4768 40329 4770
rect 42817 4768 42924 4956
rect 38906 4753 42926 4768
rect 38906 4733 39604 4753
rect 39623 4733 39681 4753
rect 39700 4750 42926 4753
rect 39700 4733 42142 4750
rect 38906 4730 42142 4733
rect 42161 4730 42219 4750
rect 42238 4730 42926 4750
rect 38906 4712 42926 4730
rect 39597 4711 39708 4712
rect 40284 4711 40491 4712
rect 42135 4708 42246 4712
rect 38964 4659 38999 4660
rect 38943 4652 38999 4659
rect 38943 4632 38972 4652
rect 38992 4632 38999 4652
rect 38943 4627 38999 4632
rect 39390 4655 39422 4662
rect 39390 4635 39396 4655
rect 39417 4635 39422 4655
rect 38112 4403 38138 4418
rect 38109 4396 38145 4403
rect 38109 4358 38115 4396
rect 38138 4358 38145 4396
rect 38109 4352 38145 4358
rect 38943 4349 38977 4627
rect 39390 4607 39422 4635
rect 39010 4599 39422 4607
rect 39010 4573 39016 4599
rect 39042 4573 39422 4599
rect 39010 4571 39422 4573
rect 39012 4570 39052 4571
rect 39179 4545 39210 4553
rect 39179 4515 39183 4545
rect 39204 4515 39210 4545
rect 38943 4341 38978 4349
rect 38943 4321 38951 4341
rect 38971 4321 38978 4341
rect 38943 4316 38978 4321
rect 38943 4315 38975 4316
rect 39179 4312 39210 4515
rect 39390 4506 39422 4571
rect 41321 4649 41401 4661
rect 41502 4656 41537 4657
rect 41321 4623 41337 4649
rect 41377 4623 41401 4649
rect 41321 4604 41401 4623
rect 41321 4578 41340 4604
rect 41380 4578 41401 4604
rect 41321 4551 41401 4578
rect 41321 4525 41344 4551
rect 41384 4525 41401 4551
rect 41321 4514 41401 4525
rect 41481 4649 41537 4656
rect 41481 4629 41510 4649
rect 41530 4629 41537 4649
rect 41481 4624 41537 4629
rect 41928 4652 41960 4659
rect 41928 4632 41934 4652
rect 41955 4632 41960 4652
rect 39390 4486 39394 4506
rect 39415 4486 39422 4506
rect 39390 4479 39422 4486
rect 39699 4423 39800 4424
rect 39597 4410 39800 4423
rect 39597 4408 39740 4410
rect 39597 4405 39674 4408
rect 39597 4378 39600 4405
rect 39629 4381 39674 4405
rect 39703 4381 39740 4408
rect 39629 4378 39740 4381
rect 39597 4377 39740 4378
rect 39776 4377 39800 4410
rect 39597 4364 39800 4377
rect 39174 4294 39210 4312
rect 39174 4277 39209 4294
rect 39107 4246 39212 4277
rect 39107 4241 39179 4246
rect 39107 4220 39138 4241
rect 39158 4225 39179 4241
rect 39199 4225 39212 4246
rect 39158 4220 39212 4225
rect 39107 4211 39212 4220
rect 41326 4214 41391 4514
rect 41481 4346 41515 4624
rect 41928 4604 41960 4632
rect 41548 4596 41960 4604
rect 41548 4570 41554 4596
rect 41580 4570 41960 4596
rect 42382 4638 42449 4645
rect 42382 4617 42399 4638
rect 42435 4617 42449 4638
rect 42382 4598 42449 4617
rect 42382 4595 42399 4598
rect 41548 4568 41960 4570
rect 41550 4567 41590 4568
rect 41717 4542 41748 4550
rect 41717 4512 41721 4542
rect 41742 4512 41748 4542
rect 41481 4338 41516 4346
rect 41481 4318 41489 4338
rect 41509 4318 41516 4338
rect 41481 4313 41516 4318
rect 41481 4312 41513 4313
rect 41717 4308 41748 4512
rect 41928 4503 41960 4568
rect 42384 4561 42399 4595
rect 42439 4561 42449 4598
rect 42384 4552 42449 4561
rect 41928 4483 41932 4503
rect 41953 4483 41960 4503
rect 41928 4476 41960 4483
rect 42237 4420 42338 4421
rect 42135 4407 42338 4420
rect 42135 4405 42278 4407
rect 42135 4402 42212 4405
rect 42135 4375 42138 4402
rect 42167 4378 42212 4402
rect 42241 4378 42278 4405
rect 42167 4375 42278 4378
rect 42135 4374 42278 4375
rect 42314 4374 42338 4407
rect 42135 4361 42338 4374
rect 41715 4296 41750 4308
rect 41646 4289 41750 4296
rect 41646 4288 41722 4289
rect 41646 4268 41667 4288
rect 41699 4269 41722 4288
rect 41747 4269 41750 4289
rect 41699 4268 41750 4269
rect 41646 4259 41750 4268
rect 41715 4257 41750 4259
rect 41326 4175 41329 4214
rect 41374 4175 41391 4214
rect 42387 4191 42438 4552
rect 42385 4189 42442 4191
rect 41326 4153 41391 4175
rect 42374 4177 42442 4189
rect 42374 4144 42385 4177
rect 42425 4144 42442 4177
rect 42374 4138 42442 4144
rect 42374 4134 42438 4138
rect 41087 4089 41198 4092
rect 42817 4089 42924 4712
rect 39130 4075 42924 4089
rect 39130 4055 41094 4075
rect 41113 4055 41171 4075
rect 41190 4071 42924 4075
rect 41190 4055 42142 4071
rect 39130 4051 42142 4055
rect 42161 4051 42219 4071
rect 42238 4051 42924 4071
rect 39130 4033 42924 4051
rect 39130 4032 40371 4033
rect 42135 4029 42246 4033
rect 40454 3981 40489 3982
rect 40433 3974 40489 3981
rect 40433 3954 40462 3974
rect 40482 3954 40489 3974
rect 40433 3949 40489 3954
rect 40880 3977 40912 3984
rect 41502 3977 41537 3978
rect 40880 3957 40886 3977
rect 40907 3957 40912 3977
rect 41481 3970 41537 3977
rect 41346 3960 41404 3965
rect 40433 3671 40467 3949
rect 40880 3929 40912 3957
rect 40500 3921 40912 3929
rect 40500 3895 40506 3921
rect 40532 3895 40912 3921
rect 40500 3893 40912 3895
rect 40502 3892 40542 3893
rect 40669 3867 40700 3875
rect 40669 3837 40673 3867
rect 40694 3837 40700 3867
rect 40433 3663 40468 3671
rect 40433 3643 40441 3663
rect 40461 3643 40468 3663
rect 40433 3638 40468 3643
rect 39174 3627 39210 3638
rect 40433 3637 40465 3638
rect 40669 3630 40700 3837
rect 40880 3828 40912 3893
rect 40880 3808 40884 3828
rect 40905 3808 40912 3828
rect 40880 3801 40912 3808
rect 41329 3951 41404 3960
rect 41329 3918 41338 3951
rect 41391 3918 41404 3951
rect 41329 3893 41404 3918
rect 41329 3860 41343 3893
rect 41396 3860 41404 3893
rect 41329 3854 41404 3860
rect 41481 3950 41510 3970
rect 41530 3950 41537 3970
rect 41481 3945 41537 3950
rect 41928 3973 41960 3980
rect 41928 3953 41934 3973
rect 41955 3953 41960 3973
rect 41189 3745 41290 3746
rect 41087 3732 41290 3745
rect 41087 3730 41230 3732
rect 41087 3727 41164 3730
rect 41087 3700 41090 3727
rect 41119 3703 41164 3727
rect 41193 3703 41230 3730
rect 41119 3700 41230 3703
rect 41087 3699 41230 3700
rect 41266 3699 41290 3732
rect 41087 3686 41290 3699
rect 39174 3604 39180 3627
rect 39204 3604 39210 3627
rect 40664 3621 40700 3630
rect 40609 3611 40706 3621
rect 39421 3609 40706 3611
rect 39174 3583 39210 3604
rect 39174 3560 39180 3583
rect 39204 3560 39210 3583
rect 39174 3407 39210 3560
rect 39386 3599 40706 3609
rect 39386 3561 39398 3599
rect 39423 3564 39442 3599
rect 39467 3564 40706 3599
rect 39423 3561 40706 3564
rect 39386 3558 40706 3561
rect 39386 3556 40703 3558
rect 39386 3553 39475 3556
rect 39402 3552 39474 3553
rect 41329 3543 41399 3854
rect 41481 3667 41515 3945
rect 41928 3925 41960 3953
rect 41548 3917 41960 3925
rect 41548 3891 41554 3917
rect 41580 3891 41960 3917
rect 41548 3889 41960 3891
rect 41550 3888 41590 3889
rect 41717 3863 41748 3871
rect 41717 3833 41721 3863
rect 41742 3833 41748 3863
rect 41481 3659 41516 3667
rect 41481 3639 41489 3659
rect 41509 3639 41516 3659
rect 41481 3634 41516 3639
rect 41717 3634 41748 3833
rect 41928 3824 41960 3889
rect 41928 3804 41932 3824
rect 41953 3804 41960 3824
rect 41928 3797 41960 3804
rect 42373 3950 42445 3968
rect 42373 3908 42386 3950
rect 42435 3908 42445 3950
rect 42373 3887 42445 3908
rect 42373 3845 42387 3887
rect 42436 3845 42445 3887
rect 42237 3741 42338 3742
rect 42135 3728 42338 3741
rect 42135 3726 42278 3728
rect 42135 3723 42212 3726
rect 42135 3696 42138 3723
rect 42167 3699 42212 3723
rect 42241 3699 42278 3726
rect 42167 3696 42278 3699
rect 42135 3695 42278 3696
rect 42314 3695 42338 3728
rect 42135 3682 42338 3695
rect 41481 3633 41513 3634
rect 41715 3631 41748 3634
rect 41681 3612 41749 3631
rect 41651 3600 41750 3612
rect 42373 3604 42445 3845
rect 42817 3604 42924 4033
rect 41651 3562 41673 3600
rect 41698 3565 41717 3600
rect 41742 3565 41750 3600
rect 41698 3562 41750 3565
rect 41651 3554 41750 3562
rect 41677 3553 41749 3554
rect 41328 3527 41399 3543
rect 41328 3511 41348 3527
rect 41329 3481 41348 3511
rect 41331 3461 41348 3481
rect 41378 3481 41399 3527
rect 42371 3523 42449 3604
rect 42816 3549 42924 3604
rect 41378 3461 41398 3481
rect 41331 3442 41398 3461
rect 42371 3421 42450 3523
rect 39165 3398 39251 3407
rect 39165 3380 39184 3398
rect 39236 3380 39251 3398
rect 39165 3376 39251 3380
rect 42335 3403 42456 3421
rect 42335 3401 42406 3403
rect 42335 3360 42350 3401
rect 42387 3362 42406 3401
rect 42443 3362 42456 3403
rect 42387 3360 42456 3362
rect 42335 3350 42456 3360
rect 39640 3322 39751 3325
rect 38955 3321 40504 3322
rect 42817 3321 42924 3549
rect 38955 3318 42114 3321
rect 42301 3318 42926 3321
rect 38955 3308 42926 3318
rect 38955 3288 39647 3308
rect 39666 3288 39724 3308
rect 39743 3303 42926 3308
rect 39743 3288 42142 3303
rect 38955 3283 42142 3288
rect 42161 3283 42219 3303
rect 42238 3283 42926 3303
rect 38955 3265 42926 3283
rect 38955 3262 40504 3265
rect 42135 3261 42246 3265
rect 39007 3214 39042 3215
rect 38986 3207 39042 3214
rect 38986 3187 39015 3207
rect 39035 3187 39042 3207
rect 38986 3182 39042 3187
rect 39433 3210 39465 3217
rect 39433 3190 39439 3210
rect 39460 3190 39465 3210
rect 38986 2904 39020 3182
rect 39433 3162 39465 3190
rect 39053 3154 39465 3162
rect 39053 3128 39059 3154
rect 39085 3128 39465 3154
rect 39053 3126 39465 3128
rect 39055 3125 39095 3126
rect 39222 3100 39253 3108
rect 39222 3070 39226 3100
rect 39247 3070 39253 3100
rect 38986 2896 39021 2904
rect 38986 2876 38994 2896
rect 39014 2876 39021 2896
rect 38986 2871 39021 2876
rect 38986 2870 39018 2871
rect 39222 2869 39253 3070
rect 39433 3061 39465 3126
rect 39433 3041 39437 3061
rect 39458 3041 39465 3061
rect 39433 3034 39465 3041
rect 40027 3201 40120 3208
rect 40027 3160 40051 3201
rect 40105 3160 40120 3201
rect 39742 2978 39843 2979
rect 39640 2965 39843 2978
rect 39640 2963 39783 2965
rect 39640 2960 39717 2963
rect 39640 2933 39643 2960
rect 39672 2936 39717 2960
rect 39746 2936 39783 2963
rect 39672 2933 39783 2936
rect 39640 2932 39783 2933
rect 39819 2932 39843 2965
rect 39640 2919 39843 2932
rect 40027 2787 40120 3160
rect 41321 3202 41401 3214
rect 41502 3209 41537 3210
rect 41321 3176 41337 3202
rect 41377 3176 41401 3202
rect 41321 3157 41401 3176
rect 41321 3131 41340 3157
rect 41380 3131 41401 3157
rect 41321 3104 41401 3131
rect 41321 3078 41344 3104
rect 41384 3078 41401 3104
rect 41321 3067 41401 3078
rect 41481 3202 41537 3209
rect 41481 3182 41510 3202
rect 41530 3182 41537 3202
rect 41481 3177 41537 3182
rect 41928 3205 41960 3212
rect 41928 3185 41934 3205
rect 41955 3185 41960 3205
rect 40027 2743 40045 2787
rect 40105 2743 40120 2787
rect 40027 2728 40120 2743
rect 41326 2767 41391 3067
rect 41481 2899 41515 3177
rect 41928 3157 41960 3185
rect 41548 3149 41960 3157
rect 41548 3123 41554 3149
rect 41580 3123 41960 3149
rect 42382 3191 42449 3198
rect 42382 3170 42399 3191
rect 42435 3170 42449 3191
rect 42382 3151 42449 3170
rect 42382 3148 42399 3151
rect 41548 3121 41960 3123
rect 41550 3120 41590 3121
rect 41717 3095 41748 3103
rect 41717 3065 41721 3095
rect 41742 3065 41748 3095
rect 41481 2891 41516 2899
rect 41481 2871 41489 2891
rect 41509 2871 41516 2891
rect 41481 2866 41516 2871
rect 41481 2865 41513 2866
rect 41717 2861 41748 3065
rect 41928 3056 41960 3121
rect 42384 3114 42399 3148
rect 42439 3114 42449 3151
rect 42384 3105 42449 3114
rect 41928 3036 41932 3056
rect 41953 3036 41960 3056
rect 41928 3029 41960 3036
rect 42237 2973 42338 2974
rect 42135 2960 42338 2973
rect 42135 2958 42278 2960
rect 42135 2955 42212 2958
rect 42135 2928 42138 2955
rect 42167 2931 42212 2955
rect 42241 2931 42278 2958
rect 42167 2928 42278 2931
rect 42135 2927 42278 2928
rect 42314 2927 42338 2960
rect 42135 2914 42338 2927
rect 41715 2849 41750 2861
rect 41646 2842 41750 2849
rect 41646 2841 41722 2842
rect 41646 2821 41667 2841
rect 41699 2822 41722 2841
rect 41747 2822 41750 2842
rect 41699 2821 41750 2822
rect 41646 2812 41750 2821
rect 41715 2810 41750 2812
rect 41326 2728 41329 2767
rect 41374 2728 41391 2767
rect 42387 2744 42438 3105
rect 42385 2742 42442 2744
rect 41326 2706 41391 2728
rect 42374 2730 42442 2742
rect 42374 2697 42385 2730
rect 42425 2697 42442 2730
rect 42374 2691 42442 2697
rect 42374 2687 42438 2691
rect 41087 2642 41198 2645
rect 42817 2642 42924 3265
rect 39350 2628 42924 2642
rect 39350 2608 41094 2628
rect 41113 2608 41171 2628
rect 41190 2624 42924 2628
rect 41190 2608 42142 2624
rect 39350 2604 42142 2608
rect 42161 2604 42219 2624
rect 42238 2604 42924 2624
rect 39350 2586 42924 2604
rect 39350 2585 40463 2586
rect 42135 2582 42246 2586
rect 40454 2534 40489 2535
rect 40433 2527 40489 2534
rect 40433 2507 40462 2527
rect 40482 2507 40489 2527
rect 40433 2502 40489 2507
rect 40880 2530 40912 2537
rect 41502 2530 41537 2531
rect 40880 2510 40886 2530
rect 40907 2510 40912 2530
rect 41481 2523 41537 2530
rect 41346 2513 41404 2518
rect 38269 2467 40122 2500
rect 38269 2402 38334 2467
rect 38465 2447 40122 2467
rect 38465 2406 40058 2447
rect 40094 2406 40122 2447
rect 40220 2467 40284 2486
rect 40220 2428 40237 2467
rect 40271 2428 40284 2467
rect 40220 2409 40284 2428
rect 38465 2402 40122 2406
rect 38269 2377 40122 2402
rect 40033 2374 40115 2377
rect 40222 1897 40284 2409
rect 40433 2224 40467 2502
rect 40880 2482 40912 2510
rect 40500 2474 40912 2482
rect 40500 2448 40506 2474
rect 40532 2448 40912 2474
rect 40500 2446 40912 2448
rect 40502 2445 40542 2446
rect 40669 2420 40700 2428
rect 40669 2390 40673 2420
rect 40694 2390 40700 2420
rect 40433 2216 40468 2224
rect 40433 2196 40441 2216
rect 40461 2196 40468 2216
rect 40433 2191 40468 2196
rect 40433 2190 40465 2191
rect 40669 2183 40700 2390
rect 40880 2381 40912 2446
rect 40880 2361 40884 2381
rect 40905 2361 40912 2381
rect 40880 2354 40912 2361
rect 41329 2504 41404 2513
rect 41329 2471 41338 2504
rect 41391 2471 41404 2504
rect 41329 2446 41404 2471
rect 41329 2413 41343 2446
rect 41396 2413 41404 2446
rect 41329 2407 41404 2413
rect 41481 2503 41510 2523
rect 41530 2503 41537 2523
rect 41481 2498 41537 2503
rect 41928 2526 41960 2533
rect 41928 2506 41934 2526
rect 41955 2506 41960 2526
rect 41189 2298 41290 2299
rect 41087 2285 41290 2298
rect 41087 2283 41230 2285
rect 41087 2280 41164 2283
rect 41087 2253 41090 2280
rect 41119 2256 41164 2280
rect 41193 2256 41230 2283
rect 41119 2253 41230 2256
rect 41087 2252 41230 2253
rect 41266 2252 41290 2285
rect 41087 2239 41290 2252
rect 40664 2165 40700 2183
rect 40631 2164 40700 2165
rect 40611 2152 40700 2164
rect 40611 2114 40623 2152
rect 40648 2117 40667 2152
rect 40692 2117 40700 2152
rect 40648 2114 40700 2117
rect 40611 2106 40700 2114
rect 40627 2105 40699 2106
rect 40180 1839 40296 1897
rect 41329 1886 41399 2407
rect 41481 2220 41515 2498
rect 41928 2478 41960 2506
rect 41548 2470 41960 2478
rect 41548 2444 41554 2470
rect 41580 2444 41960 2470
rect 41548 2442 41960 2444
rect 41550 2441 41590 2442
rect 41717 2416 41748 2424
rect 41717 2386 41721 2416
rect 41742 2386 41748 2416
rect 41481 2212 41516 2220
rect 41481 2192 41489 2212
rect 41509 2192 41516 2212
rect 41481 2187 41516 2192
rect 41717 2187 41748 2386
rect 41928 2377 41960 2442
rect 41928 2357 41932 2377
rect 41953 2357 41960 2377
rect 41928 2350 41960 2357
rect 42373 2503 42445 2521
rect 42373 2461 42386 2503
rect 42435 2461 42445 2503
rect 42373 2440 42445 2461
rect 42373 2398 42387 2440
rect 42436 2398 42445 2440
rect 42237 2294 42338 2295
rect 42135 2281 42338 2294
rect 42135 2279 42278 2281
rect 42135 2276 42212 2279
rect 42135 2249 42138 2276
rect 42167 2252 42212 2276
rect 42241 2252 42278 2279
rect 42167 2249 42278 2252
rect 42135 2248 42278 2249
rect 42314 2248 42338 2281
rect 42135 2235 42338 2248
rect 41481 2186 41513 2187
rect 41715 2184 41748 2187
rect 41681 2165 41749 2184
rect 41651 2153 41750 2165
rect 41651 2115 41673 2153
rect 41698 2118 41717 2153
rect 41742 2118 41750 2153
rect 41698 2115 41750 2118
rect 41651 2107 41750 2115
rect 41677 2106 41749 2107
rect 40180 1768 40192 1839
rect 40271 1768 40296 1839
rect 40180 1748 40296 1768
rect 41310 1685 41412 1886
rect 42373 1878 42445 2398
rect 42817 1974 42924 2586
rect 42816 1938 42924 1974
rect 42971 2097 43125 2122
rect 42971 1985 42984 2097
rect 43105 1985 43125 2097
rect 41274 1648 41440 1685
rect 41274 1569 41311 1648
rect 41395 1569 41440 1648
rect 41274 1531 41440 1569
rect 42351 1477 42448 1878
rect 42809 1802 42929 1938
rect 42816 1796 42924 1802
rect 42281 1448 42456 1477
rect 42281 1369 42327 1448
rect 42427 1369 42456 1448
rect 42281 1344 42456 1369
rect 42816 1253 42920 1796
rect 42659 1223 42930 1253
rect 42659 1136 42693 1223
rect 42763 1215 42930 1223
rect 42763 1136 42826 1215
rect 42659 1128 42826 1136
rect 42896 1128 42930 1215
rect 42659 1082 42930 1128
rect 42971 1011 43125 1985
rect 42969 995 43125 1011
rect 42969 970 43121 995
rect 42969 875 42999 970
rect 43089 875 43121 970
rect 42969 862 43121 875
rect 37787 755 37839 795
rect 37789 708 37839 755
rect 33333 697 37839 708
rect 33333 649 33348 697
rect 33389 649 37839 697
rect 33333 644 37839 649
rect 33333 629 33398 644
rect 37789 638 37839 644
rect 32260 510 32463 523
rect 32260 477 32284 510
rect 32320 509 32463 510
rect 32320 506 32431 509
rect 32320 479 32357 506
rect 32386 482 32431 506
rect 32460 482 32463 509
rect 32386 479 32463 482
rect 32320 477 32463 479
rect 32260 464 32463 477
rect 32260 463 32361 464
rect 32638 401 32670 408
rect 32638 381 32645 401
rect 32666 381 32670 401
rect 32638 316 32670 381
rect 32850 372 32881 598
rect 33085 571 33117 572
rect 33082 566 33117 571
rect 33082 546 33089 566
rect 33109 546 33117 566
rect 33082 538 33117 546
rect 32850 342 32856 372
rect 32877 342 32881 372
rect 32850 334 32881 342
rect 33008 316 33048 317
rect 32638 314 33050 316
rect 32638 288 33018 314
rect 33044 288 33050 314
rect 32638 280 33050 288
rect 32638 252 32670 280
rect 33083 260 33117 538
rect 32638 232 32643 252
rect 32664 232 32670 252
rect 32638 225 32670 232
rect 32849 253 32882 260
rect 32849 230 32857 253
rect 32877 230 32882 253
rect 32352 155 32463 176
rect 32056 154 32463 155
rect 32056 134 32360 154
rect 32379 134 32437 154
rect 32456 134 32463 154
rect 32056 117 32463 134
rect 22059 71 22117 95
rect 32056 83 32457 117
rect 22059 13 22076 71
rect 22105 32 22117 71
rect 32849 39 32882 230
rect 33061 255 33117 260
rect 33061 235 33068 255
rect 33088 235 33117 255
rect 33061 228 33117 235
rect 33061 227 33096 228
rect 22105 31 32413 32
rect 32844 31 32885 39
rect 22105 13 32885 31
rect 22059 -6 32885 13
rect 22059 -9 32413 -6
rect 32844 -9 32885 -6
<< via1 >>
rect 901 13739 937 13772
rect 1949 13735 1985 13768
rect 5424 14236 5502 14294
rect 4361 14114 4427 14169
rect 3099 13985 3169 14058
rect 901 13060 937 13093
rect 3396 13055 3432 13088
rect 901 12292 937 12325
rect 1949 12288 1985 12321
rect 901 11613 937 11646
rect 3439 11610 3475 11643
rect 902 10772 938 10805
rect 1950 10768 1986 10801
rect 902 10093 938 10126
rect 3397 10088 3433 10121
rect 902 9325 938 9358
rect 1950 9321 1986 9354
rect 902 8646 938 8679
rect 16143 14233 16221 14291
rect 27097 14234 27175 14292
rect 15083 14108 15135 14152
rect 13822 13984 13874 14034
rect 9898 13357 9934 13390
rect 4505 8637 4541 8670
rect 899 7731 935 7764
rect 1947 7727 1983 7760
rect 899 7052 935 7085
rect 3394 7047 3430 7080
rect 899 6284 935 6317
rect 1947 6280 1983 6313
rect 8850 12682 8886 12715
rect 9898 12678 9934 12711
rect 11609 13733 11645 13766
rect 12657 13729 12693 13762
rect 11609 13054 11645 13087
rect 14104 13049 14140 13082
rect 7403 11915 7439 11948
rect 9898 11910 9934 11943
rect 8850 11235 8886 11268
rect 9898 11231 9934 11264
rect 11609 12286 11645 12319
rect 12657 12282 12693 12315
rect 11609 11607 11645 11640
rect 14147 11604 14183 11637
rect 7361 10393 7397 10426
rect 9899 10390 9935 10423
rect 8851 9715 8887 9748
rect 9899 9711 9935 9744
rect 11610 10766 11646 10799
rect 12658 10762 12694 10795
rect 11610 10087 11646 10120
rect 14105 10082 14141 10115
rect 7404 8948 7440 8981
rect 9899 8943 9935 8976
rect 8851 8268 8887 8301
rect 9899 8264 9935 8297
rect 11610 9319 11646 9352
rect 12658 9315 12694 9348
rect 11610 8640 11646 8673
rect 26034 14112 26100 14167
rect 24772 13983 24842 14056
rect 20606 13351 20642 13384
rect 15213 8631 15249 8664
rect 6293 7358 6329 7391
rect 899 5605 935 5638
rect 3437 5602 3473 5635
rect 900 4764 936 4797
rect 1948 4760 1984 4793
rect 4850 4766 4886 4799
rect 900 4085 936 4118
rect 3395 4080 3431 4113
rect 900 3317 936 3350
rect 1948 3313 1984 3346
rect 900 2638 936 2671
rect 127 1972 206 2084
rect 2881 1776 2998 1851
rect 1833 1581 1903 1656
rect 784 1365 884 1444
rect 331 1136 401 1223
rect 99 888 189 983
rect 9896 7349 9932 7382
rect 8848 6674 8884 6707
rect 9896 6670 9932 6703
rect 11607 7725 11643 7758
rect 12655 7721 12691 7754
rect 11607 7046 11643 7079
rect 14102 7041 14138 7074
rect 7401 5907 7437 5940
rect 9896 5902 9932 5935
rect 8848 5227 8884 5260
rect 9896 5223 9932 5256
rect 11607 6278 11643 6311
rect 12655 6274 12691 6307
rect 19558 12676 19594 12709
rect 20606 12672 20642 12705
rect 22574 13737 22610 13770
rect 23622 13733 23658 13766
rect 22574 13058 22610 13091
rect 25069 13053 25105 13086
rect 18111 11909 18147 11942
rect 20606 11904 20642 11937
rect 19558 11229 19594 11262
rect 20606 11225 20642 11258
rect 22574 12290 22610 12323
rect 23622 12286 23658 12319
rect 22574 11611 22610 11644
rect 25112 11608 25148 11641
rect 18069 10387 18105 10420
rect 20607 10384 20643 10417
rect 19559 9709 19595 9742
rect 20607 9705 20643 9738
rect 22575 10770 22611 10803
rect 23623 10766 23659 10799
rect 22575 10091 22611 10124
rect 25070 10086 25106 10119
rect 18112 8942 18148 8975
rect 20607 8937 20643 8970
rect 19559 8262 19595 8295
rect 20607 8258 20643 8291
rect 22575 9323 22611 9356
rect 23623 9319 23659 9352
rect 22575 8644 22611 8677
rect 37816 14231 37894 14289
rect 36756 14106 36808 14150
rect 35495 13982 35547 14032
rect 31571 13355 31607 13388
rect 26178 8635 26214 8668
rect 17001 7352 17037 7385
rect 11607 5599 11643 5632
rect 14145 5596 14181 5629
rect 7359 4385 7395 4418
rect 9897 4382 9933 4415
rect 8849 3707 8885 3740
rect 9897 3703 9933 3736
rect 11608 4758 11644 4791
rect 12656 4754 12692 4787
rect 15558 4760 15594 4793
rect 11608 4079 11644 4112
rect 14103 4074 14139 4107
rect 7402 2940 7438 2973
rect 9897 2935 9933 2968
rect 8849 2260 8885 2293
rect 9897 2256 9933 2289
rect 7811 1776 7890 1847
rect 11608 3311 11644 3344
rect 12656 3307 12692 3340
rect 11608 2632 11644 2665
rect 10603 1993 10724 2105
rect 8930 1577 9014 1656
rect 9946 1377 10046 1456
rect 10312 1144 10382 1231
rect 10445 1136 10515 1223
rect 10835 1966 10914 2078
rect 13589 1770 13706 1845
rect 12541 1575 12611 1650
rect 11492 1359 11592 1438
rect 11039 1130 11109 1217
rect 10618 883 10708 978
rect 10807 882 10897 977
rect 20604 7343 20640 7376
rect 19556 6668 19592 6701
rect 20604 6664 20640 6697
rect 22572 7729 22608 7762
rect 23620 7725 23656 7758
rect 22572 7050 22608 7083
rect 25067 7045 25103 7078
rect 18109 5901 18145 5934
rect 20604 5896 20640 5929
rect 19556 5221 19592 5254
rect 20604 5217 20640 5250
rect 22572 6282 22608 6315
rect 23620 6278 23656 6311
rect 30523 12680 30559 12713
rect 31571 12676 31607 12709
rect 33282 13731 33318 13764
rect 34330 13727 34366 13760
rect 33282 13052 33318 13085
rect 35777 13047 35813 13080
rect 29076 11913 29112 11946
rect 31571 11908 31607 11941
rect 30523 11233 30559 11266
rect 31571 11229 31607 11262
rect 33282 12284 33318 12317
rect 34330 12280 34366 12313
rect 33282 11605 33318 11638
rect 35820 11602 35856 11635
rect 29034 10391 29070 10424
rect 31572 10388 31608 10421
rect 30524 9713 30560 9746
rect 31572 9709 31608 9742
rect 33283 10764 33319 10797
rect 34331 10760 34367 10793
rect 33283 10085 33319 10118
rect 35778 10080 35814 10113
rect 29077 8946 29113 8979
rect 31572 8941 31608 8974
rect 30524 8266 30560 8299
rect 31572 8262 31608 8295
rect 33283 9317 33319 9350
rect 34331 9313 34367 9346
rect 33283 8638 33319 8671
rect 42279 13349 42315 13382
rect 36886 8629 36922 8662
rect 27966 7356 28002 7389
rect 22572 5603 22608 5636
rect 25110 5600 25146 5633
rect 18067 4379 18103 4412
rect 20605 4376 20641 4409
rect 19557 3701 19593 3734
rect 20605 3697 20641 3730
rect 22573 4762 22609 4795
rect 23621 4758 23657 4791
rect 26523 4764 26559 4797
rect 22573 4083 22609 4116
rect 25068 4078 25104 4111
rect 18110 2934 18146 2967
rect 20605 2929 20641 2962
rect 19557 2254 19593 2287
rect 20605 2250 20641 2283
rect 18519 1770 18598 1841
rect 22573 3315 22609 3348
rect 23621 3311 23657 3344
rect 22573 2636 22609 2669
rect 21311 1987 21432 2099
rect 19638 1571 19722 1650
rect 20654 1371 20754 1450
rect 21020 1138 21090 1225
rect 21153 1130 21223 1217
rect 10611 479 10647 512
rect 21800 1970 21879 2082
rect 24554 1774 24671 1849
rect 23506 1579 23576 1654
rect 22457 1363 22557 1442
rect 22004 1134 22074 1221
rect 21326 877 21416 972
rect 21772 886 21862 981
rect 31569 7347 31605 7380
rect 30521 6672 30557 6705
rect 31569 6668 31605 6701
rect 33280 7723 33316 7756
rect 34328 7719 34364 7752
rect 33280 7044 33316 7077
rect 35775 7039 35811 7072
rect 29074 5905 29110 5938
rect 31569 5900 31605 5933
rect 30521 5225 30557 5258
rect 31569 5221 31605 5254
rect 33280 6276 33316 6309
rect 34328 6272 34364 6305
rect 41231 12674 41267 12707
rect 42279 12670 42315 12703
rect 39784 11907 39820 11940
rect 42279 11902 42315 11935
rect 41231 11227 41267 11260
rect 42279 11223 42315 11256
rect 39742 10385 39778 10418
rect 42280 10382 42316 10415
rect 41232 9707 41268 9740
rect 42280 9703 42316 9736
rect 39785 8940 39821 8973
rect 42280 8935 42316 8968
rect 41232 8260 41268 8293
rect 42280 8256 42316 8289
rect 38674 7350 38710 7383
rect 33280 5597 33316 5630
rect 35818 5594 35854 5627
rect 29032 4383 29068 4416
rect 31570 4380 31606 4413
rect 30522 3705 30558 3738
rect 31570 3701 31606 3734
rect 33281 4756 33317 4789
rect 34329 4752 34365 4785
rect 37231 4758 37267 4791
rect 33281 4077 33317 4110
rect 35776 4072 35812 4105
rect 29075 2938 29111 2971
rect 31570 2933 31606 2966
rect 30522 2258 30558 2291
rect 31570 2254 31606 2287
rect 29484 1774 29563 1845
rect 33281 3309 33317 3342
rect 34329 3305 34365 3338
rect 33281 2630 33317 2663
rect 32276 1991 32397 2103
rect 30603 1575 30687 1654
rect 31619 1375 31719 1454
rect 31985 1142 32055 1229
rect 32118 1134 32188 1221
rect 21248 466 21284 499
rect 19210 -98 19368 -16
rect 32508 1964 32587 2076
rect 35262 1768 35379 1843
rect 34214 1573 34284 1648
rect 33165 1357 33265 1436
rect 32712 1128 32782 1215
rect 32291 881 32381 976
rect 32480 880 32570 975
rect 42277 7341 42313 7374
rect 41229 6666 41265 6699
rect 42277 6662 42313 6695
rect 39782 5899 39818 5932
rect 42277 5894 42313 5927
rect 41229 5219 41265 5252
rect 42277 5215 42313 5248
rect 39740 4377 39776 4410
rect 42278 4374 42314 4407
rect 41230 3699 41266 3732
rect 42278 3695 42314 3728
rect 39783 2932 39819 2965
rect 42278 2927 42314 2960
rect 41230 2252 41266 2285
rect 42278 2248 42314 2281
rect 40192 1768 40271 1839
rect 42984 1985 43105 2097
rect 41311 1569 41395 1648
rect 42327 1369 42427 1448
rect 42693 1136 42763 1223
rect 42826 1128 42896 1215
rect 42999 875 43089 970
rect 32284 477 32320 510
<< metal2 >>
rect 16162 14311 27237 14315
rect 16126 14308 27237 14311
rect 5393 14306 27237 14308
rect 37799 14306 37907 14309
rect 5393 14294 37907 14306
rect 5393 14236 5424 14294
rect 5502 14292 37907 14294
rect 5502 14291 27097 14292
rect 5502 14236 16143 14291
rect 5393 14233 16143 14236
rect 16221 14251 27097 14291
rect 16221 14233 16234 14251
rect 5393 14221 16234 14233
rect 120 13787 227 14221
rect 16126 14220 16234 14221
rect 27066 14234 27097 14251
rect 27175 14289 37907 14292
rect 27175 14234 37816 14289
rect 27066 14231 37816 14234
rect 37894 14231 37907 14289
rect 27066 14219 37907 14231
rect 37799 14218 37907 14219
rect 4345 14169 4444 14180
rect 4345 14114 4361 14169
rect 4427 14156 4444 14169
rect 15066 14166 15153 14170
rect 26018 14167 26117 14174
rect 26018 14166 26034 14167
rect 15066 14156 26034 14166
rect 4427 14152 26034 14156
rect 4427 14114 15083 14152
rect 4345 14108 15083 14114
rect 15135 14112 26034 14152
rect 26100 14166 26117 14167
rect 26100 14154 26141 14166
rect 36739 14154 36826 14168
rect 26100 14150 36826 14154
rect 26100 14112 36756 14150
rect 15135 14108 36756 14112
rect 4345 14106 36756 14108
rect 36808 14106 36826 14150
rect 4345 14102 36826 14106
rect 4345 14100 15153 14102
rect 4362 14099 15153 14100
rect 15066 14091 15153 14099
rect 26018 14098 36826 14102
rect 26035 14097 36826 14098
rect 36739 14089 36826 14097
rect 3085 14058 3206 14079
rect 3085 13985 3099 14058
rect 3169 14042 3206 14058
rect 24758 14056 24879 14074
rect 13802 14045 13901 14048
rect 24758 14045 24772 14056
rect 13802 14042 24772 14045
rect 3169 14034 24772 14042
rect 3169 13985 13822 14034
rect 3085 13984 13822 13985
rect 13874 13984 24772 14034
rect 3085 13983 24772 13984
rect 24842 14040 24879 14056
rect 35475 14040 35574 14046
rect 24842 14032 35574 14040
rect 24842 13983 35495 14032
rect 3085 13982 35495 13983
rect 35547 13982 35574 14032
rect 3085 13981 35574 13982
rect 3085 13972 13901 13981
rect 3085 13969 3206 13972
rect 13802 13964 13901 13972
rect 24758 13970 35574 13981
rect 24758 13967 24879 13970
rect 35475 13962 35574 13970
rect 120 13772 3865 13787
rect 21793 13785 21900 13792
rect 120 13739 901 13772
rect 937 13768 3865 13772
rect 937 13739 1949 13768
rect 120 13735 1949 13739
rect 1985 13735 3865 13768
rect 120 13718 3865 13735
rect 120 13112 227 13718
rect 2727 13716 3865 13718
rect 10592 13781 10936 13784
rect 10592 13766 14573 13781
rect 10592 13733 11609 13766
rect 11645 13762 14573 13766
rect 11645 13733 12657 13762
rect 10592 13729 12657 13733
rect 12693 13729 14573 13762
rect 21793 13770 25538 13785
rect 10592 13712 14573 13729
rect 10592 13703 10936 13712
rect 13435 13710 14573 13712
rect 6471 13407 7976 13408
rect 10608 13407 10715 13703
rect 6471 13390 10715 13407
rect 6471 13357 9898 13390
rect 9934 13357 10715 13390
rect 6471 13338 10715 13357
rect 6471 13336 7976 13338
rect 120 13093 4260 13112
rect 120 13060 901 13093
rect 937 13088 4260 13093
rect 937 13060 3396 13088
rect 120 13055 3396 13060
rect 3432 13055 4260 13088
rect 120 13043 4260 13055
rect 120 12340 227 13043
rect 2648 13042 4260 13043
rect 10608 12732 10715 13338
rect 6471 12715 10715 12732
rect 6471 12682 8850 12715
rect 8886 12711 10715 12715
rect 8886 12682 9898 12711
rect 6471 12678 9898 12682
rect 9934 12678 10715 12711
rect 6471 12663 10715 12678
rect 6471 12660 8010 12663
rect 2877 12343 3120 12348
rect 2825 12340 4085 12343
rect 120 12325 4085 12340
rect 120 12292 901 12325
rect 937 12321 4085 12325
rect 937 12292 1949 12321
rect 120 12288 1949 12292
rect 1985 12288 4085 12321
rect 120 12271 4085 12288
rect 120 11665 227 12271
rect 2877 12262 3120 12271
rect 6472 11960 8187 11961
rect 10608 11960 10715 12663
rect 6472 11948 10715 11960
rect 6472 11915 7403 11948
rect 7439 11943 10715 11948
rect 7439 11915 9898 11943
rect 6472 11910 9898 11915
rect 9934 11910 10715 11943
rect 6472 11891 10715 11910
rect 2859 11665 4309 11667
rect 120 11646 4309 11665
rect 120 11613 901 11646
rect 937 11643 4309 11646
rect 937 11613 3439 11643
rect 120 11610 3439 11613
rect 3475 11610 4309 11643
rect 120 11596 4309 11610
rect 120 11061 227 11596
rect 2859 11595 4309 11596
rect 6094 11285 8108 11287
rect 10608 11285 10715 11891
rect 6094 11268 10715 11285
rect 6094 11235 8850 11268
rect 8886 11264 10715 11268
rect 8886 11235 9898 11264
rect 6094 11231 9898 11235
rect 9934 11231 10715 11264
rect 6094 11216 10715 11231
rect 7779 11214 7967 11216
rect 120 11060 228 11061
rect 121 11037 228 11060
rect 119 10993 228 11037
rect 121 10820 228 10993
rect 10608 11043 10715 11216
rect 10828 13106 10935 13703
rect 17179 13401 18684 13402
rect 21316 13401 21423 13748
rect 17179 13384 21423 13401
rect 17179 13351 20606 13384
rect 20642 13351 21423 13384
rect 17179 13332 21423 13351
rect 17179 13330 18684 13332
rect 10828 13087 14968 13106
rect 10828 13054 11609 13087
rect 11645 13082 14968 13087
rect 11645 13054 14104 13082
rect 10828 13049 14104 13054
rect 14140 13049 14968 13082
rect 10828 13037 14968 13049
rect 10828 12334 10935 13037
rect 13356 13036 14968 13037
rect 21316 12726 21423 13332
rect 17179 12709 21423 12726
rect 17179 12676 19558 12709
rect 19594 12705 21423 12709
rect 19594 12676 20606 12705
rect 17179 12672 20606 12676
rect 20642 12672 21423 12705
rect 17179 12657 21423 12672
rect 17179 12654 18718 12657
rect 13585 12337 13828 12342
rect 13533 12334 14793 12337
rect 10828 12319 14793 12334
rect 10828 12286 11609 12319
rect 11645 12315 14793 12319
rect 11645 12286 12657 12315
rect 10828 12282 12657 12286
rect 12693 12282 14793 12315
rect 10828 12265 14793 12282
rect 10828 11659 10935 12265
rect 13585 12256 13828 12265
rect 17180 11954 18895 11955
rect 21316 11954 21423 12657
rect 17180 11942 21423 11954
rect 17180 11909 18111 11942
rect 18147 11937 21423 11942
rect 18147 11909 20606 11937
rect 17180 11904 20606 11909
rect 20642 11904 21423 11937
rect 17180 11885 21423 11904
rect 13567 11659 15017 11661
rect 10828 11640 15017 11659
rect 10828 11607 11609 11640
rect 11645 11637 15017 11640
rect 11645 11607 14147 11637
rect 10828 11604 14147 11607
rect 14183 11604 15017 11637
rect 10828 11590 15017 11604
rect 10828 11055 10935 11590
rect 13567 11589 15017 11590
rect 16802 11279 18816 11281
rect 21316 11279 21423 11885
rect 16802 11262 21423 11279
rect 16802 11229 19558 11262
rect 19594 11258 21423 11262
rect 19594 11229 20606 11258
rect 16802 11225 20606 11229
rect 20642 11225 21423 11258
rect 16802 11210 21423 11225
rect 18487 11208 18675 11210
rect 10828 11054 10936 11055
rect 10608 10999 10717 11043
rect 10829 11031 10936 11054
rect 10608 10976 10715 10999
rect 10827 10987 10936 11031
rect 10608 10975 10716 10976
rect 2869 10820 3057 10822
rect 121 10805 4053 10820
rect 121 10772 902 10805
rect 938 10801 4053 10805
rect 938 10772 1950 10801
rect 121 10768 1950 10772
rect 1986 10768 4053 10801
rect 121 10751 4053 10768
rect 121 10145 228 10751
rect 2728 10749 4053 10751
rect 6481 10440 7977 10441
rect 10609 10440 10716 10975
rect 6481 10426 10716 10440
rect 6481 10393 7361 10426
rect 7397 10423 10716 10426
rect 7397 10393 9899 10423
rect 6481 10390 9899 10393
rect 9935 10390 10716 10423
rect 6481 10371 10716 10390
rect 6481 10369 7977 10371
rect 121 10126 4262 10145
rect 121 10093 902 10126
rect 938 10121 4262 10126
rect 938 10093 3397 10121
rect 121 10088 3397 10093
rect 3433 10088 4262 10121
rect 121 10076 4262 10088
rect 121 9373 228 10076
rect 2649 10075 4262 10076
rect 7716 9765 7959 9774
rect 10609 9765 10716 10371
rect 6481 9748 10716 9765
rect 6481 9715 8851 9748
rect 8887 9744 10716 9748
rect 8887 9715 9899 9744
rect 6481 9711 9899 9715
rect 9935 9711 10716 9744
rect 6481 9696 10716 9711
rect 6481 9693 8011 9696
rect 7716 9688 7959 9693
rect 2826 9373 3835 9376
rect 121 9358 3835 9373
rect 121 9325 902 9358
rect 938 9354 3835 9358
rect 938 9325 1950 9354
rect 121 9321 1950 9325
rect 1986 9321 3835 9354
rect 121 9304 3835 9321
rect 121 8698 228 9304
rect 6481 8993 8188 8994
rect 10609 8993 10716 9696
rect 6481 8981 10716 8993
rect 6481 8948 7404 8981
rect 7440 8976 10716 8981
rect 7440 8948 9899 8976
rect 6481 8943 9899 8948
rect 9935 8943 10716 8976
rect 6481 8924 10716 8943
rect 2860 8699 4365 8700
rect 2860 8698 4565 8699
rect 121 8683 4565 8698
rect 121 8679 4568 8683
rect 121 8646 902 8679
rect 938 8670 4568 8679
rect 938 8646 4505 8670
rect 121 8637 4505 8646
rect 4541 8637 4568 8670
rect 121 8629 4568 8637
rect 121 8112 228 8629
rect 2860 8628 4568 8629
rect 4330 8625 4568 8628
rect 6537 8318 8109 8320
rect 10609 8318 10716 8924
rect 6537 8301 10716 8318
rect 6537 8268 8851 8301
rect 8887 8297 10716 8301
rect 8887 8268 9899 8297
rect 6537 8264 9899 8268
rect 9935 8264 10716 8297
rect 6537 8249 10716 8264
rect 114 7920 230 8112
rect 10609 8108 10716 8249
rect 10829 10814 10936 10987
rect 21316 11037 21423 11210
rect 21793 13737 22574 13770
rect 22610 13766 25538 13770
rect 22610 13737 23622 13766
rect 21793 13733 23622 13737
rect 23658 13733 25538 13766
rect 21793 13716 25538 13733
rect 21793 13110 21900 13716
rect 24400 13714 25538 13716
rect 32265 13779 32609 13782
rect 32265 13764 36246 13779
rect 32265 13731 33282 13764
rect 33318 13760 36246 13764
rect 33318 13731 34330 13760
rect 32265 13727 34330 13731
rect 34366 13727 36246 13760
rect 32265 13710 36246 13727
rect 32265 13701 32609 13710
rect 35108 13708 36246 13710
rect 29633 13405 29649 13406
rect 32281 13405 32388 13701
rect 29633 13388 32388 13405
rect 29633 13355 31571 13388
rect 31607 13355 32388 13388
rect 29633 13336 32388 13355
rect 29633 13334 29649 13336
rect 21793 13091 25933 13110
rect 21793 13058 22574 13091
rect 22610 13086 25933 13091
rect 22610 13058 25069 13086
rect 21793 13053 25069 13058
rect 25105 13053 25933 13086
rect 21793 13041 25933 13053
rect 21793 12338 21900 13041
rect 24321 13040 25933 13041
rect 32281 12730 32388 13336
rect 29633 12713 32388 12730
rect 29633 12680 30523 12713
rect 30559 12709 32388 12713
rect 30559 12680 31571 12709
rect 29633 12676 31571 12680
rect 31607 12676 32388 12709
rect 29633 12661 32388 12676
rect 29633 12658 29683 12661
rect 24550 12341 24793 12346
rect 24498 12338 25758 12341
rect 21793 12323 25758 12338
rect 21793 12290 22574 12323
rect 22610 12319 25758 12323
rect 22610 12290 23622 12319
rect 21793 12286 23622 12290
rect 23658 12286 25758 12319
rect 21793 12269 25758 12286
rect 21793 11663 21900 12269
rect 24550 12260 24793 12269
rect 28145 11958 29860 11959
rect 32281 11958 32388 12661
rect 28145 11946 32388 11958
rect 28145 11913 29076 11946
rect 29112 11941 32388 11946
rect 29112 11913 31571 11941
rect 28145 11908 31571 11913
rect 31607 11908 32388 11941
rect 28145 11889 32388 11908
rect 24532 11663 25982 11665
rect 21793 11644 25982 11663
rect 21793 11611 22574 11644
rect 22610 11641 25982 11644
rect 22610 11611 25112 11641
rect 21793 11608 25112 11611
rect 25148 11608 25982 11641
rect 21793 11594 25982 11608
rect 21793 11059 21900 11594
rect 24532 11593 25982 11594
rect 27767 11283 29781 11285
rect 32281 11283 32388 11889
rect 27767 11266 32388 11283
rect 27767 11233 30523 11266
rect 30559 11262 32388 11266
rect 30559 11233 31571 11262
rect 27767 11229 31571 11233
rect 31607 11229 32388 11262
rect 27767 11214 32388 11229
rect 29452 11212 29640 11214
rect 21793 11058 21901 11059
rect 21316 10993 21425 11037
rect 21794 11035 21901 11058
rect 21316 10970 21423 10993
rect 21792 10991 21901 11035
rect 21316 10969 21424 10970
rect 13577 10814 13765 10816
rect 10829 10799 14761 10814
rect 10829 10766 11610 10799
rect 11646 10795 14761 10799
rect 11646 10766 12658 10795
rect 10829 10762 12658 10766
rect 12694 10762 14761 10795
rect 10829 10745 14761 10762
rect 10829 10139 10936 10745
rect 13436 10743 14761 10745
rect 17189 10434 18685 10435
rect 21317 10434 21424 10969
rect 17189 10420 21424 10434
rect 17189 10387 18069 10420
rect 18105 10417 21424 10420
rect 18105 10387 20607 10417
rect 17189 10384 20607 10387
rect 20643 10384 21424 10417
rect 17189 10365 21424 10384
rect 17189 10363 18685 10365
rect 10829 10120 14970 10139
rect 10829 10087 11610 10120
rect 11646 10115 14970 10120
rect 11646 10087 14105 10115
rect 10829 10082 14105 10087
rect 14141 10082 14970 10115
rect 10829 10070 14970 10082
rect 10829 9367 10936 10070
rect 13357 10069 14970 10070
rect 18424 9759 18667 9768
rect 21317 9759 21424 10365
rect 17189 9742 21424 9759
rect 17189 9709 19559 9742
rect 19595 9738 21424 9742
rect 19595 9709 20607 9738
rect 17189 9705 20607 9709
rect 20643 9705 21424 9738
rect 17189 9690 21424 9705
rect 17189 9687 18719 9690
rect 18424 9682 18667 9687
rect 13534 9367 14543 9370
rect 10829 9352 14543 9367
rect 10829 9319 11610 9352
rect 11646 9348 14543 9352
rect 11646 9319 12658 9348
rect 10829 9315 12658 9319
rect 12694 9315 14543 9348
rect 10829 9298 14543 9315
rect 10829 8692 10936 9298
rect 17189 8987 18896 8988
rect 21317 8987 21424 9690
rect 17189 8975 21424 8987
rect 17189 8942 18112 8975
rect 18148 8970 21424 8975
rect 18148 8942 20607 8970
rect 17189 8937 20607 8942
rect 20643 8937 21424 8970
rect 17189 8918 21424 8937
rect 13568 8693 15073 8694
rect 13568 8692 15273 8693
rect 10829 8677 15273 8692
rect 10829 8673 15276 8677
rect 10829 8640 11610 8673
rect 11646 8664 15276 8673
rect 11646 8640 15213 8664
rect 10829 8631 15213 8640
rect 15249 8631 15276 8664
rect 10829 8623 15276 8631
rect 118 7779 225 7920
rect 10604 7916 10720 8108
rect 10829 8106 10936 8623
rect 13568 8622 15276 8623
rect 15038 8619 15276 8622
rect 17245 8312 18817 8314
rect 21317 8312 21424 8918
rect 17245 8295 21424 8312
rect 17245 8262 19559 8295
rect 19595 8291 21424 8295
rect 19595 8262 20607 8291
rect 17245 8258 20607 8262
rect 20643 8258 21424 8291
rect 17245 8243 21424 8258
rect 118 7764 4297 7779
rect 118 7731 899 7764
rect 935 7760 4297 7764
rect 935 7731 1947 7760
rect 118 7727 1947 7731
rect 1983 7727 4297 7760
rect 118 7710 4297 7727
rect 118 7104 225 7710
rect 2725 7708 4297 7710
rect 6266 7400 6400 7403
rect 6487 7400 6504 7403
rect 6266 7399 7974 7400
rect 10606 7399 10713 7916
rect 10822 7914 10938 8106
rect 21317 8102 21424 8243
rect 21794 10818 21901 10991
rect 32281 11041 32388 11214
rect 32501 13104 32608 13701
rect 40271 13399 40357 13400
rect 42989 13399 43096 13945
rect 40271 13382 43096 13399
rect 40271 13349 42279 13382
rect 42315 13349 43096 13382
rect 40271 13330 43096 13349
rect 40271 13328 40357 13330
rect 32501 13085 36641 13104
rect 32501 13052 33282 13085
rect 33318 13080 36641 13085
rect 33318 13052 35777 13080
rect 32501 13047 35777 13052
rect 35813 13047 36641 13080
rect 32501 13035 36641 13047
rect 32501 12332 32608 13035
rect 35029 13034 36641 13035
rect 42989 12724 43096 13330
rect 40271 12707 43096 12724
rect 40271 12674 41231 12707
rect 41267 12703 43096 12707
rect 41267 12674 42279 12703
rect 40271 12670 42279 12674
rect 42315 12670 43096 12703
rect 40271 12655 43096 12670
rect 40271 12652 40391 12655
rect 35258 12335 35501 12340
rect 35206 12332 36466 12335
rect 32501 12317 36466 12332
rect 32501 12284 33282 12317
rect 33318 12313 36466 12317
rect 33318 12284 34330 12313
rect 32501 12280 34330 12284
rect 34366 12280 36466 12313
rect 32501 12263 36466 12280
rect 32501 11657 32608 12263
rect 35258 12254 35501 12263
rect 38853 11952 40568 11953
rect 42989 11952 43096 12655
rect 38853 11940 43096 11952
rect 38853 11907 39784 11940
rect 39820 11935 43096 11940
rect 39820 11907 42279 11935
rect 38853 11902 42279 11907
rect 42315 11902 43096 11935
rect 38853 11883 43096 11902
rect 35240 11657 36690 11659
rect 32501 11638 36690 11657
rect 32501 11605 33282 11638
rect 33318 11635 36690 11638
rect 33318 11605 35820 11635
rect 32501 11602 35820 11605
rect 35856 11602 36690 11635
rect 32501 11588 36690 11602
rect 32501 11053 32608 11588
rect 35240 11587 36690 11588
rect 39173 11277 40489 11279
rect 42989 11277 43096 11883
rect 39173 11260 43096 11277
rect 39173 11227 41231 11260
rect 41267 11256 43096 11260
rect 41267 11227 42279 11256
rect 39173 11223 42279 11227
rect 42315 11223 43096 11256
rect 39173 11208 43096 11223
rect 40160 11206 40348 11208
rect 32501 11052 32609 11053
rect 32281 10997 32390 11041
rect 32502 11029 32609 11052
rect 32281 10974 32388 10997
rect 32500 10985 32609 11029
rect 32281 10973 32389 10974
rect 24542 10818 24730 10820
rect 21794 10803 25726 10818
rect 21794 10770 22575 10803
rect 22611 10799 25726 10803
rect 22611 10770 23623 10799
rect 21794 10766 23623 10770
rect 23659 10766 25726 10799
rect 21794 10749 25726 10766
rect 21794 10143 21901 10749
rect 24401 10747 25726 10749
rect 28154 10438 29650 10439
rect 32282 10438 32389 10973
rect 28154 10424 32389 10438
rect 28154 10391 29034 10424
rect 29070 10421 32389 10424
rect 29070 10391 31572 10421
rect 28154 10388 31572 10391
rect 31608 10388 32389 10421
rect 28154 10369 32389 10388
rect 28154 10367 29650 10369
rect 21794 10124 25935 10143
rect 21794 10091 22575 10124
rect 22611 10119 25935 10124
rect 22611 10091 25070 10119
rect 21794 10086 25070 10091
rect 25106 10086 25935 10119
rect 21794 10074 25935 10086
rect 21794 9371 21901 10074
rect 24322 10073 25935 10074
rect 29389 9763 29632 9772
rect 32282 9763 32389 10369
rect 28154 9746 32389 9763
rect 28154 9713 30524 9746
rect 30560 9742 32389 9746
rect 30560 9713 31572 9742
rect 28154 9709 31572 9713
rect 31608 9709 32389 9742
rect 28154 9694 32389 9709
rect 28154 9691 29684 9694
rect 29389 9686 29632 9691
rect 24499 9371 24961 9374
rect 21794 9356 24961 9371
rect 21794 9323 22575 9356
rect 22611 9352 24961 9356
rect 22611 9323 23623 9352
rect 21794 9319 23623 9323
rect 23659 9319 24961 9352
rect 21794 9302 24961 9319
rect 21794 8696 21901 9302
rect 28154 8991 29861 8992
rect 32282 8991 32389 9694
rect 28154 8979 32389 8991
rect 28154 8946 29077 8979
rect 29113 8974 32389 8979
rect 29113 8946 31572 8974
rect 28154 8941 31572 8946
rect 31608 8941 32389 8974
rect 28154 8922 32389 8941
rect 24533 8697 26038 8698
rect 24533 8696 26238 8697
rect 21794 8681 26238 8696
rect 21794 8677 26241 8681
rect 21794 8644 22575 8677
rect 22611 8668 26241 8677
rect 22611 8644 26178 8668
rect 21794 8635 26178 8644
rect 26214 8635 26241 8668
rect 21794 8627 26241 8635
rect 21794 8110 21901 8627
rect 24533 8626 26241 8627
rect 26003 8623 26241 8626
rect 28210 8316 29782 8318
rect 32282 8316 32389 8922
rect 28210 8299 32389 8316
rect 28210 8266 30524 8299
rect 30560 8295 32389 8299
rect 30560 8266 31572 8295
rect 28210 8262 31572 8266
rect 31608 8262 32389 8295
rect 28210 8247 32389 8262
rect 6266 7391 10713 7399
rect 6266 7358 6293 7391
rect 6329 7382 10713 7391
rect 6329 7358 9896 7382
rect 6266 7349 9896 7358
rect 9932 7349 10713 7382
rect 6266 7345 10713 7349
rect 6269 7330 10713 7345
rect 6269 7329 7974 7330
rect 6385 7328 7974 7329
rect 6385 7313 6507 7328
rect 118 7085 4353 7104
rect 118 7052 899 7085
rect 935 7080 4353 7085
rect 935 7052 3394 7080
rect 118 7047 3394 7052
rect 3430 7047 4353 7080
rect 118 7035 4353 7047
rect 118 6332 225 7035
rect 2646 7034 4353 7035
rect 10606 6724 10713 7330
rect 6999 6707 10713 6724
rect 6999 6674 8848 6707
rect 8884 6703 10713 6707
rect 8884 6674 9896 6703
rect 6999 6670 9896 6674
rect 9932 6670 10713 6703
rect 6999 6655 10713 6670
rect 6999 6652 8008 6655
rect 2875 6335 3118 6340
rect 2823 6332 4353 6335
rect 118 6317 4353 6332
rect 118 6284 899 6317
rect 935 6313 4353 6317
rect 935 6284 1947 6313
rect 118 6280 1947 6284
rect 1983 6280 4353 6313
rect 118 6263 4353 6280
rect 118 5657 225 6263
rect 2875 6254 3118 6263
rect 6572 5952 8185 5953
rect 10606 5952 10713 6655
rect 6572 5940 10713 5952
rect 6572 5907 7401 5940
rect 7437 5935 10713 5940
rect 7437 5907 9896 5935
rect 6572 5902 9896 5907
rect 9932 5902 10713 5935
rect 6572 5883 10713 5902
rect 2857 5657 4353 5659
rect 118 5638 4353 5657
rect 118 5605 899 5638
rect 935 5635 4353 5638
rect 935 5605 3437 5635
rect 118 5602 3437 5605
rect 3473 5602 4353 5635
rect 118 5588 4353 5602
rect 118 5053 225 5588
rect 2857 5587 4353 5588
rect 6781 5277 8106 5279
rect 10606 5277 10713 5883
rect 6781 5260 10713 5277
rect 6781 5227 8848 5260
rect 8884 5256 10713 5260
rect 8884 5227 9896 5256
rect 6781 5223 9896 5227
rect 9932 5223 10713 5256
rect 6781 5208 10713 5223
rect 7777 5206 7965 5208
rect 118 5052 226 5053
rect 119 5029 226 5052
rect 117 4985 226 5029
rect 119 4812 226 4985
rect 10606 5035 10713 5208
rect 10826 7773 10933 7914
rect 21312 7910 21428 8102
rect 21787 7918 21903 8110
rect 32282 8106 32389 8247
rect 32502 10812 32609 10985
rect 42989 11035 43096 11208
rect 42989 10991 43098 11035
rect 42989 10968 43096 10991
rect 42989 10967 43097 10968
rect 35250 10812 35438 10814
rect 32502 10797 36434 10812
rect 32502 10764 33283 10797
rect 33319 10793 36434 10797
rect 33319 10764 34331 10793
rect 32502 10760 34331 10764
rect 34367 10760 36434 10793
rect 32502 10743 36434 10760
rect 32502 10137 32609 10743
rect 35109 10741 36434 10743
rect 38862 10432 40358 10433
rect 42990 10432 43097 10967
rect 38862 10418 43097 10432
rect 38862 10385 39742 10418
rect 39778 10415 43097 10418
rect 39778 10385 42280 10415
rect 38862 10382 42280 10385
rect 42316 10382 43097 10415
rect 38862 10363 43097 10382
rect 38862 10361 40358 10363
rect 32502 10118 36643 10137
rect 32502 10085 33283 10118
rect 33319 10113 36643 10118
rect 33319 10085 35778 10113
rect 32502 10080 35778 10085
rect 35814 10080 36643 10113
rect 32502 10068 36643 10080
rect 32502 9365 32609 10068
rect 35030 10067 36643 10068
rect 40097 9757 40340 9766
rect 42990 9757 43097 10363
rect 38862 9740 43097 9757
rect 38862 9707 41232 9740
rect 41268 9736 43097 9740
rect 41268 9707 42280 9736
rect 38862 9703 42280 9707
rect 42316 9703 43097 9736
rect 38862 9688 43097 9703
rect 38862 9685 40392 9688
rect 40097 9680 40340 9685
rect 35207 9365 35665 9368
rect 32502 9350 35665 9365
rect 32502 9317 33283 9350
rect 33319 9346 35665 9350
rect 33319 9317 34331 9346
rect 32502 9313 34331 9317
rect 34367 9313 35665 9346
rect 32502 9296 35665 9313
rect 32502 8690 32609 9296
rect 38862 8985 40569 8986
rect 42990 8985 43097 9688
rect 38862 8973 43097 8985
rect 38862 8940 39785 8973
rect 39821 8968 43097 8973
rect 39821 8940 42280 8968
rect 38862 8935 42280 8940
rect 42316 8935 43097 8968
rect 38862 8916 43097 8935
rect 35241 8691 36746 8692
rect 35241 8690 36946 8691
rect 32502 8675 36946 8690
rect 32502 8671 36949 8675
rect 32502 8638 33283 8671
rect 33319 8662 36949 8671
rect 33319 8638 36886 8662
rect 32502 8629 36886 8638
rect 36922 8629 36949 8662
rect 32502 8621 36949 8629
rect 10826 7758 15005 7773
rect 10826 7725 11607 7758
rect 11643 7754 15005 7758
rect 11643 7725 12655 7754
rect 10826 7721 12655 7725
rect 12691 7721 15005 7754
rect 10826 7704 15005 7721
rect 10826 7098 10933 7704
rect 13433 7702 15005 7704
rect 16974 7394 17108 7397
rect 17195 7394 17212 7397
rect 16974 7393 18682 7394
rect 21314 7393 21421 7910
rect 16974 7385 21421 7393
rect 16974 7352 17001 7385
rect 17037 7376 21421 7385
rect 17037 7352 20604 7376
rect 16974 7343 20604 7352
rect 20640 7343 21421 7376
rect 16974 7339 21421 7343
rect 16977 7324 21421 7339
rect 16977 7323 18682 7324
rect 17093 7322 18682 7323
rect 17093 7307 17215 7322
rect 10826 7079 15061 7098
rect 10826 7046 11607 7079
rect 11643 7074 15061 7079
rect 11643 7046 14102 7074
rect 10826 7041 14102 7046
rect 14138 7041 15061 7074
rect 10826 7029 15061 7041
rect 10826 6326 10933 7029
rect 13354 7028 15061 7029
rect 21314 6718 21421 7324
rect 17707 6701 21421 6718
rect 17707 6668 19556 6701
rect 19592 6697 21421 6701
rect 19592 6668 20604 6697
rect 17707 6664 20604 6668
rect 20640 6664 21421 6697
rect 17707 6649 21421 6664
rect 17707 6646 18716 6649
rect 13583 6329 13826 6334
rect 13531 6326 15061 6329
rect 10826 6311 15061 6326
rect 10826 6278 11607 6311
rect 11643 6307 15061 6311
rect 11643 6278 12655 6307
rect 10826 6274 12655 6278
rect 12691 6274 15061 6307
rect 10826 6257 15061 6274
rect 10826 5651 10933 6257
rect 13583 6248 13826 6257
rect 17280 5946 18893 5947
rect 21314 5946 21421 6649
rect 17280 5934 21421 5946
rect 17280 5901 18109 5934
rect 18145 5929 21421 5934
rect 18145 5901 20604 5929
rect 17280 5896 20604 5901
rect 20640 5896 21421 5929
rect 17280 5877 21421 5896
rect 13565 5651 15061 5653
rect 10826 5632 15061 5651
rect 10826 5599 11607 5632
rect 11643 5629 15061 5632
rect 11643 5599 14145 5629
rect 10826 5596 14145 5599
rect 14181 5596 15061 5629
rect 10826 5582 15061 5596
rect 10826 5047 10933 5582
rect 13565 5581 15061 5582
rect 17489 5271 18814 5273
rect 21314 5271 21421 5877
rect 17489 5254 21421 5271
rect 17489 5221 19556 5254
rect 19592 5250 21421 5254
rect 19592 5221 20604 5250
rect 17489 5217 20604 5221
rect 20640 5217 21421 5250
rect 17489 5202 21421 5217
rect 18485 5200 18673 5202
rect 10826 5046 10934 5047
rect 10606 4991 10715 5035
rect 10827 5023 10934 5046
rect 10606 4968 10713 4991
rect 10825 4979 10934 5023
rect 10606 4967 10714 4968
rect 2867 4812 3055 4814
rect 4646 4812 5064 4819
rect 119 4799 5064 4812
rect 119 4797 4850 4799
rect 119 4764 900 4797
rect 936 4793 4850 4797
rect 936 4764 1948 4793
rect 119 4760 1948 4764
rect 1984 4766 4850 4793
rect 4886 4766 5064 4799
rect 1984 4760 5064 4766
rect 119 4748 5064 4760
rect 119 4743 4740 4748
rect 119 4137 226 4743
rect 2726 4741 4740 4743
rect 6525 4432 7975 4433
rect 10607 4432 10714 4967
rect 6525 4418 10714 4432
rect 6525 4385 7359 4418
rect 7395 4415 10714 4418
rect 7395 4385 9897 4415
rect 6525 4382 9897 4385
rect 9933 4382 10714 4415
rect 6525 4363 10714 4382
rect 6525 4361 7975 4363
rect 119 4118 4362 4137
rect 119 4085 900 4118
rect 936 4113 4362 4118
rect 936 4085 3395 4113
rect 119 4080 3395 4085
rect 3431 4080 4362 4113
rect 119 4068 4362 4080
rect 119 3365 226 4068
rect 2647 4067 4362 4068
rect 7714 3757 7957 3766
rect 10607 3757 10714 4363
rect 6749 3740 10714 3757
rect 6749 3707 8849 3740
rect 8885 3736 10714 3740
rect 8885 3707 9897 3736
rect 6749 3703 9897 3707
rect 9933 3703 10714 3736
rect 6749 3688 10714 3703
rect 6749 3685 8009 3688
rect 7714 3680 7957 3685
rect 2824 3365 4363 3368
rect 119 3350 4363 3365
rect 119 3317 900 3350
rect 936 3346 4363 3350
rect 936 3317 1948 3346
rect 119 3313 1948 3317
rect 1984 3313 4363 3346
rect 119 3296 4363 3313
rect 119 2690 226 3296
rect 6574 2985 8186 2986
rect 10607 2985 10714 3688
rect 6574 2973 10714 2985
rect 6574 2940 7402 2973
rect 7438 2968 10714 2973
rect 7438 2940 9897 2968
rect 6574 2935 9897 2940
rect 9933 2935 10714 2968
rect 6574 2916 10714 2935
rect 2858 2690 4363 2692
rect 119 2671 4363 2690
rect 119 2638 900 2671
rect 936 2638 4363 2671
rect 119 2621 4363 2638
rect 119 2122 226 2621
rect 2858 2620 4363 2621
rect 7749 2310 8107 2312
rect 10607 2310 10714 2916
rect 7749 2293 10714 2310
rect 7749 2260 8849 2293
rect 8885 2289 10714 2293
rect 8885 2260 9897 2289
rect 7749 2256 9897 2260
rect 9933 2259 10714 2289
rect 10827 4806 10934 4979
rect 21314 5029 21421 5202
rect 21791 7777 21898 7918
rect 32277 7914 32393 8106
rect 32502 8104 32609 8621
rect 35241 8620 36949 8621
rect 36711 8617 36949 8620
rect 38918 8310 40490 8312
rect 42990 8310 43097 8916
rect 38918 8293 43097 8310
rect 38918 8260 41232 8293
rect 41268 8289 43097 8293
rect 41268 8260 42280 8289
rect 38918 8256 42280 8260
rect 42316 8256 43097 8289
rect 38918 8241 43097 8256
rect 21791 7762 25970 7777
rect 21791 7729 22572 7762
rect 22608 7758 25970 7762
rect 22608 7729 23620 7758
rect 21791 7725 23620 7729
rect 23656 7725 25970 7758
rect 21791 7708 25970 7725
rect 21791 7102 21898 7708
rect 24398 7706 25970 7708
rect 27939 7398 28073 7401
rect 28160 7398 28177 7401
rect 27939 7397 29647 7398
rect 32279 7397 32386 7914
rect 32495 7912 32611 8104
rect 42990 8100 43097 8241
rect 27939 7389 32386 7397
rect 27939 7356 27966 7389
rect 28002 7380 32386 7389
rect 28002 7356 31569 7380
rect 27939 7347 31569 7356
rect 31605 7347 32386 7380
rect 27939 7343 32386 7347
rect 27942 7328 32386 7343
rect 27942 7327 29647 7328
rect 28058 7326 29647 7327
rect 28058 7311 28180 7326
rect 21791 7083 26026 7102
rect 21791 7050 22572 7083
rect 22608 7078 26026 7083
rect 22608 7050 25067 7078
rect 21791 7045 25067 7050
rect 25103 7045 26026 7078
rect 21791 7033 26026 7045
rect 21791 6330 21898 7033
rect 24319 7032 26026 7033
rect 32279 6722 32386 7328
rect 28672 6705 32386 6722
rect 28672 6672 30521 6705
rect 30557 6701 32386 6705
rect 30557 6672 31569 6701
rect 28672 6668 31569 6672
rect 31605 6668 32386 6701
rect 28672 6653 32386 6668
rect 28672 6650 29681 6653
rect 24548 6333 24791 6338
rect 24496 6330 26026 6333
rect 21791 6315 26026 6330
rect 21791 6282 22572 6315
rect 22608 6311 26026 6315
rect 22608 6282 23620 6311
rect 21791 6278 23620 6282
rect 23656 6278 26026 6311
rect 21791 6261 26026 6278
rect 21791 5655 21898 6261
rect 24548 6252 24791 6261
rect 28245 5950 29858 5951
rect 32279 5950 32386 6653
rect 28245 5938 32386 5950
rect 28245 5905 29074 5938
rect 29110 5933 32386 5938
rect 29110 5905 31569 5933
rect 28245 5900 31569 5905
rect 31605 5900 32386 5933
rect 28245 5881 32386 5900
rect 24530 5655 26026 5657
rect 21791 5636 26026 5655
rect 21791 5603 22572 5636
rect 22608 5633 26026 5636
rect 22608 5603 25110 5633
rect 21791 5600 25110 5603
rect 25146 5600 26026 5633
rect 21791 5586 26026 5600
rect 21791 5051 21898 5586
rect 24530 5585 26026 5586
rect 28454 5275 29779 5277
rect 32279 5275 32386 5881
rect 28454 5258 32386 5275
rect 28454 5225 30521 5258
rect 30557 5254 32386 5258
rect 30557 5225 31569 5254
rect 28454 5221 31569 5225
rect 31605 5221 32386 5254
rect 28454 5206 32386 5221
rect 29450 5204 29638 5206
rect 21791 5050 21899 5051
rect 21314 4985 21423 5029
rect 21792 5027 21899 5050
rect 21314 4962 21421 4985
rect 21790 4983 21899 5027
rect 21314 4961 21422 4962
rect 13575 4806 13763 4808
rect 15354 4806 15772 4813
rect 10827 4793 15772 4806
rect 10827 4791 15558 4793
rect 10827 4758 11608 4791
rect 11644 4787 15558 4791
rect 11644 4758 12656 4787
rect 10827 4754 12656 4758
rect 12692 4760 15558 4787
rect 15594 4760 15772 4793
rect 12692 4754 15772 4760
rect 10827 4742 15772 4754
rect 10827 4737 15448 4742
rect 10827 4131 10934 4737
rect 13434 4735 15448 4737
rect 17233 4426 18683 4427
rect 21315 4426 21422 4961
rect 17233 4412 21422 4426
rect 17233 4379 18067 4412
rect 18103 4409 21422 4412
rect 18103 4379 20605 4409
rect 17233 4376 20605 4379
rect 20641 4376 21422 4409
rect 17233 4357 21422 4376
rect 17233 4355 18683 4357
rect 10827 4112 15070 4131
rect 10827 4079 11608 4112
rect 11644 4107 15070 4112
rect 11644 4079 14103 4107
rect 10827 4074 14103 4079
rect 14139 4074 15070 4107
rect 10827 4062 15070 4074
rect 10827 3359 10934 4062
rect 13355 4061 15070 4062
rect 18422 3751 18665 3760
rect 21315 3751 21422 4357
rect 17457 3734 21422 3751
rect 17457 3701 19557 3734
rect 19593 3730 21422 3734
rect 19593 3701 20605 3730
rect 17457 3697 20605 3701
rect 20641 3697 21422 3730
rect 17457 3682 21422 3697
rect 17457 3679 18717 3682
rect 18422 3674 18665 3679
rect 13532 3359 15071 3362
rect 10827 3344 15071 3359
rect 10827 3311 11608 3344
rect 11644 3340 15071 3344
rect 11644 3311 12656 3340
rect 10827 3307 12656 3311
rect 12692 3307 15071 3340
rect 10827 3290 15071 3307
rect 10827 2684 10934 3290
rect 17282 2979 18894 2980
rect 21315 2979 21422 3682
rect 17282 2967 21422 2979
rect 17282 2934 18110 2967
rect 18146 2962 21422 2967
rect 18146 2934 20605 2962
rect 17282 2929 20605 2934
rect 20641 2929 21422 2962
rect 17282 2910 21422 2929
rect 13566 2684 15071 2686
rect 10827 2665 15071 2684
rect 10827 2632 11608 2665
rect 11644 2632 15071 2665
rect 10827 2615 15071 2632
rect 9933 2256 10753 2259
rect 7749 2241 10753 2256
rect 94 2084 227 2122
rect 94 1972 127 2084
rect 206 2053 227 2084
rect 10582 2105 10753 2241
rect 10827 2116 10934 2615
rect 13566 2614 15071 2615
rect 18457 2304 18815 2306
rect 21315 2304 21422 2910
rect 18457 2287 21422 2304
rect 18457 2254 19557 2287
rect 19593 2283 21422 2287
rect 19593 2254 20605 2283
rect 18457 2250 20605 2254
rect 20641 2253 21422 2283
rect 21792 4810 21899 4983
rect 32279 5033 32386 5206
rect 32499 7771 32606 7912
rect 42985 7908 43101 8100
rect 32499 7756 36678 7771
rect 32499 7723 33280 7756
rect 33316 7752 36678 7756
rect 33316 7723 34328 7752
rect 32499 7719 34328 7723
rect 34364 7719 36678 7752
rect 32499 7702 36678 7719
rect 32499 7096 32606 7702
rect 35106 7700 36678 7702
rect 38647 7392 38781 7395
rect 38868 7392 38885 7395
rect 38647 7391 40355 7392
rect 42987 7391 43094 7908
rect 38647 7383 43094 7391
rect 38647 7350 38674 7383
rect 38710 7374 43094 7383
rect 38710 7350 42277 7374
rect 38647 7341 42277 7350
rect 42313 7341 43094 7374
rect 38647 7337 43094 7341
rect 38650 7322 43094 7337
rect 38650 7321 40355 7322
rect 38766 7320 40355 7321
rect 38766 7305 38888 7320
rect 32499 7077 36734 7096
rect 32499 7044 33280 7077
rect 33316 7072 36734 7077
rect 33316 7044 35775 7072
rect 32499 7039 35775 7044
rect 35811 7039 36734 7072
rect 32499 7027 36734 7039
rect 32499 6324 32606 7027
rect 35027 7026 36734 7027
rect 42987 6716 43094 7322
rect 39877 6699 43094 6716
rect 39877 6666 41229 6699
rect 41265 6695 43094 6699
rect 41265 6666 42277 6695
rect 39877 6662 42277 6666
rect 42313 6662 43094 6695
rect 39877 6647 43094 6662
rect 39877 6644 40389 6647
rect 35256 6327 35499 6332
rect 35204 6324 36734 6327
rect 32499 6309 36734 6324
rect 32499 6276 33280 6309
rect 33316 6305 36734 6309
rect 33316 6276 34328 6305
rect 32499 6272 34328 6276
rect 34364 6272 36734 6305
rect 32499 6255 36734 6272
rect 32499 5649 32606 6255
rect 35256 6246 35499 6255
rect 38953 5944 40566 5945
rect 42987 5944 43094 6647
rect 38953 5932 43094 5944
rect 38953 5899 39782 5932
rect 39818 5927 43094 5932
rect 39818 5899 42277 5927
rect 38953 5894 42277 5899
rect 42313 5894 43094 5927
rect 38953 5875 43094 5894
rect 35238 5649 36734 5651
rect 32499 5630 36734 5649
rect 32499 5597 33280 5630
rect 33316 5627 36734 5630
rect 33316 5597 35818 5627
rect 32499 5594 35818 5597
rect 35854 5594 36734 5627
rect 32499 5580 36734 5594
rect 32499 5045 32606 5580
rect 35238 5579 36734 5580
rect 39162 5269 40487 5271
rect 42987 5269 43094 5875
rect 39162 5252 43094 5269
rect 39162 5219 41229 5252
rect 41265 5248 43094 5252
rect 41265 5219 42277 5248
rect 39162 5215 42277 5219
rect 42313 5215 43094 5248
rect 39162 5200 43094 5215
rect 40158 5198 40346 5200
rect 32499 5044 32607 5045
rect 32279 4989 32388 5033
rect 32500 5021 32607 5044
rect 32279 4966 32386 4989
rect 32498 4977 32607 5021
rect 32279 4965 32387 4966
rect 24540 4810 24728 4812
rect 26319 4810 26737 4817
rect 21792 4797 26737 4810
rect 21792 4795 26523 4797
rect 21792 4762 22573 4795
rect 22609 4791 26523 4795
rect 22609 4762 23621 4791
rect 21792 4758 23621 4762
rect 23657 4764 26523 4791
rect 26559 4764 26737 4797
rect 23657 4758 26737 4764
rect 21792 4746 26737 4758
rect 21792 4741 26413 4746
rect 21792 4135 21899 4741
rect 24399 4739 26413 4741
rect 28198 4430 29648 4431
rect 32280 4430 32387 4965
rect 28198 4416 32387 4430
rect 28198 4383 29032 4416
rect 29068 4413 32387 4416
rect 29068 4383 31570 4413
rect 28198 4380 31570 4383
rect 31606 4380 32387 4413
rect 28198 4361 32387 4380
rect 28198 4359 29648 4361
rect 21792 4116 26035 4135
rect 21792 4083 22573 4116
rect 22609 4111 26035 4116
rect 22609 4083 25068 4111
rect 21792 4078 25068 4083
rect 25104 4078 26035 4111
rect 21792 4066 26035 4078
rect 21792 3363 21899 4066
rect 24320 4065 26035 4066
rect 29387 3755 29630 3764
rect 32280 3755 32387 4361
rect 28422 3738 32387 3755
rect 28422 3705 30522 3738
rect 30558 3734 32387 3738
rect 30558 3705 31570 3734
rect 28422 3701 31570 3705
rect 31606 3701 32387 3734
rect 28422 3686 32387 3701
rect 28422 3683 29682 3686
rect 29387 3678 29630 3683
rect 24497 3363 25111 3366
rect 21792 3348 25111 3363
rect 21792 3315 22573 3348
rect 22609 3344 25111 3348
rect 22609 3315 23621 3344
rect 21792 3311 23621 3315
rect 23657 3311 25111 3344
rect 21792 3294 25111 3311
rect 21792 2688 21899 3294
rect 28247 2983 29859 2984
rect 32280 2983 32387 3686
rect 28247 2971 32387 2983
rect 28247 2938 29075 2971
rect 29111 2966 32387 2971
rect 29111 2938 31570 2966
rect 28247 2933 31570 2938
rect 31606 2933 32387 2966
rect 28247 2914 32387 2933
rect 24531 2688 25111 2690
rect 21792 2669 25111 2688
rect 21792 2636 22573 2669
rect 22609 2636 25111 2669
rect 21792 2619 25111 2636
rect 20641 2250 21461 2253
rect 18457 2235 21461 2250
rect 206 2009 239 2053
rect 206 1972 227 2009
rect 94 1955 227 1972
rect 10582 1993 10603 2105
rect 10724 1993 10753 2105
rect 10582 1943 10753 1993
rect 10802 2078 10935 2116
rect 10802 1966 10835 2078
rect 10914 2047 10935 2078
rect 21290 2099 21461 2235
rect 21792 2120 21899 2619
rect 24531 2618 25111 2619
rect 29422 2308 29780 2310
rect 32280 2308 32387 2914
rect 29422 2291 32387 2308
rect 29422 2258 30522 2291
rect 30558 2287 32387 2291
rect 30558 2258 31570 2287
rect 29422 2254 31570 2258
rect 31606 2257 32387 2287
rect 32500 4804 32607 4977
rect 42987 5027 43094 5200
rect 42987 4983 43096 5027
rect 42987 4960 43094 4983
rect 42987 4959 43095 4960
rect 35248 4804 35436 4806
rect 37027 4804 37445 4811
rect 32500 4791 37445 4804
rect 32500 4789 37231 4791
rect 32500 4756 33281 4789
rect 33317 4785 37231 4789
rect 33317 4756 34329 4785
rect 32500 4752 34329 4756
rect 34365 4758 37231 4785
rect 37267 4758 37445 4791
rect 34365 4752 37445 4758
rect 32500 4740 37445 4752
rect 32500 4735 37121 4740
rect 32500 4129 32607 4735
rect 35107 4733 37121 4735
rect 38906 4424 40356 4425
rect 42988 4424 43095 4959
rect 38906 4410 43095 4424
rect 38906 4377 39740 4410
rect 39776 4407 43095 4410
rect 39776 4377 42278 4407
rect 38906 4374 42278 4377
rect 42314 4374 43095 4407
rect 38906 4355 43095 4374
rect 38906 4353 40356 4355
rect 32500 4110 36743 4129
rect 32500 4077 33281 4110
rect 33317 4105 36743 4110
rect 33317 4077 35776 4105
rect 32500 4072 35776 4077
rect 35812 4072 36743 4105
rect 32500 4060 36743 4072
rect 32500 3357 32607 4060
rect 35028 4059 36743 4060
rect 40095 3749 40338 3758
rect 42988 3749 43095 4355
rect 39130 3732 43095 3749
rect 39130 3699 41230 3732
rect 41266 3728 43095 3732
rect 41266 3699 42278 3728
rect 39130 3695 42278 3699
rect 42314 3695 43095 3728
rect 39130 3680 43095 3695
rect 39130 3677 40390 3680
rect 40095 3672 40338 3677
rect 35205 3357 35655 3360
rect 32500 3342 35655 3357
rect 32500 3309 33281 3342
rect 33317 3338 35655 3342
rect 33317 3309 34329 3338
rect 32500 3305 34329 3309
rect 34365 3305 35655 3338
rect 32500 3288 35655 3305
rect 32500 2682 32607 3288
rect 38955 2977 40567 2978
rect 42988 2977 43095 3680
rect 38955 2965 43095 2977
rect 38955 2932 39783 2965
rect 39819 2960 43095 2965
rect 39819 2932 42278 2960
rect 38955 2927 42278 2932
rect 42314 2927 43095 2960
rect 38955 2908 43095 2927
rect 35239 2682 35655 2684
rect 32500 2663 35655 2682
rect 32500 2630 33281 2663
rect 33317 2630 35655 2663
rect 32500 2613 35655 2630
rect 31606 2254 32426 2257
rect 29422 2239 32426 2254
rect 10914 2003 10947 2047
rect 10914 1966 10935 2003
rect 10802 1949 10935 1966
rect 21290 1987 21311 2099
rect 21432 1987 21461 2099
rect 21290 1937 21461 1987
rect 21767 2082 21900 2120
rect 21767 1970 21800 2082
rect 21879 2051 21900 2082
rect 32255 2103 32426 2239
rect 32500 2114 32607 2613
rect 35239 2612 35655 2613
rect 40130 2302 40488 2304
rect 42988 2302 43095 2908
rect 40130 2285 43095 2302
rect 40130 2252 41230 2285
rect 41266 2281 43095 2285
rect 41266 2252 42278 2281
rect 40130 2248 42278 2252
rect 42314 2251 43095 2281
rect 42314 2248 43134 2251
rect 40130 2233 43134 2248
rect 21879 2007 21912 2051
rect 21879 1970 21900 2007
rect 21767 1953 21900 1970
rect 32255 1991 32276 2103
rect 32397 1991 32426 2103
rect 32255 1941 32426 1991
rect 32475 2076 32608 2114
rect 32475 1964 32508 2076
rect 32587 2045 32608 2076
rect 42963 2097 43134 2233
rect 32587 2001 32620 2045
rect 32587 1964 32608 2001
rect 32475 1947 32608 1964
rect 42963 1985 42984 2097
rect 43105 1985 43134 2097
rect 42963 1935 43134 1985
rect 2852 1851 7915 1860
rect 24525 1856 29588 1858
rect 18484 1854 29588 1856
rect 2852 1776 2881 1851
rect 2998 1847 7915 1851
rect 2998 1776 7811 1847
rect 7890 1839 7915 1847
rect 13560 1849 29588 1854
rect 13560 1845 24554 1849
rect 13560 1839 13589 1845
rect 7890 1776 13589 1839
rect 2852 1770 13589 1776
rect 13706 1841 24554 1845
rect 13706 1770 18519 1841
rect 18598 1774 24554 1841
rect 24671 1845 29588 1849
rect 24671 1774 29484 1845
rect 29563 1837 29588 1845
rect 35233 1843 40296 1852
rect 35233 1837 35262 1843
rect 29563 1774 35262 1837
rect 18598 1771 35262 1774
rect 18598 1770 18623 1771
rect 2852 1769 18623 1770
rect 2852 1760 7915 1769
rect 13560 1754 18623 1769
rect 24525 1768 35262 1771
rect 35379 1839 40296 1843
rect 35379 1768 40192 1839
rect 40271 1768 40296 1839
rect 24525 1767 40296 1768
rect 24525 1758 29588 1767
rect 35233 1752 40296 1767
rect 1808 1657 9039 1683
rect 12516 1670 19747 1677
rect 23481 1670 30712 1681
rect 12516 1657 30712 1670
rect 1808 1656 30712 1657
rect 1808 1581 1833 1656
rect 1903 1581 8930 1656
rect 1808 1577 8930 1581
rect 9014 1655 30712 1656
rect 34189 1655 41420 1675
rect 9014 1654 41420 1655
rect 9014 1650 23506 1654
rect 9014 1577 12541 1650
rect 1808 1575 12541 1577
rect 12611 1575 19638 1650
rect 1808 1571 19638 1575
rect 19722 1579 23506 1650
rect 23576 1579 30603 1654
rect 19722 1575 30603 1579
rect 30687 1648 41420 1654
rect 30687 1575 34214 1648
rect 19722 1573 34214 1575
rect 34284 1573 41311 1648
rect 19722 1571 41311 1573
rect 1808 1550 9039 1571
rect 12516 1569 41311 1571
rect 41395 1569 41420 1648
rect 12516 1548 30712 1569
rect 12516 1544 23584 1548
rect 19633 1539 23584 1544
rect 34189 1542 41420 1569
rect 759 1463 10066 1473
rect 20567 1471 22743 1473
rect 20567 1467 31739 1471
rect 11467 1463 31739 1467
rect 759 1461 31739 1463
rect 33140 1461 42447 1465
rect 759 1456 42447 1461
rect 759 1444 9946 1456
rect 759 1365 784 1444
rect 884 1377 9946 1444
rect 10046 1454 42447 1456
rect 10046 1450 31619 1454
rect 10046 1438 20654 1450
rect 10046 1377 11492 1438
rect 884 1365 11492 1377
rect 759 1361 11492 1365
rect 759 1356 10066 1361
rect 11467 1359 11492 1361
rect 11592 1371 20654 1438
rect 20754 1442 31619 1450
rect 20754 1371 22457 1442
rect 11592 1363 22457 1371
rect 22557 1375 31619 1442
rect 31719 1448 42447 1454
rect 31719 1436 42327 1448
rect 31719 1375 33165 1436
rect 22557 1363 33165 1375
rect 11592 1359 33165 1363
rect 11467 1354 31739 1359
rect 33140 1357 33165 1359
rect 33265 1369 42327 1436
rect 42427 1369 42447 1448
rect 33265 1357 42447 1369
rect 11467 1350 22743 1354
rect 20567 1333 22743 1350
rect 33140 1348 42447 1357
rect 293 1254 10553 1256
rect 21178 1254 22124 1258
rect 293 1250 11382 1254
rect 21178 1252 32226 1254
rect 21178 1250 33055 1252
rect 293 1248 33055 1250
rect 293 1231 42934 1248
rect 293 1223 10312 1231
rect 293 1136 331 1223
rect 401 1144 10312 1223
rect 10382 1229 42934 1231
rect 10382 1225 31985 1229
rect 10382 1223 21020 1225
rect 10382 1144 10445 1223
rect 401 1136 10445 1144
rect 10515 1217 21020 1223
rect 10515 1136 11039 1217
rect 293 1130 11039 1136
rect 11109 1138 21020 1217
rect 21090 1221 31985 1225
rect 21090 1217 22004 1221
rect 21090 1138 21153 1217
rect 11109 1130 21153 1138
rect 21223 1134 22004 1217
rect 22074 1142 31985 1221
rect 32055 1223 42934 1229
rect 32055 1221 42693 1223
rect 32055 1142 32118 1221
rect 22074 1134 32118 1142
rect 32188 1215 42693 1221
rect 32188 1134 32712 1215
rect 21223 1130 32712 1134
rect 293 1128 32712 1130
rect 32782 1136 42693 1215
rect 42763 1215 42934 1223
rect 42763 1136 42826 1215
rect 32782 1128 42826 1136
rect 42896 1128 42934 1215
rect 293 1098 42934 1128
rect 293 1094 10553 1098
rect 11001 1096 42934 1098
rect 11001 1092 32226 1096
rect 11001 1088 21261 1092
rect 32674 1086 42934 1096
rect 74 1007 10747 1012
rect 21307 1010 21912 1012
rect 74 1006 11263 1007
rect 21307 1006 32420 1010
rect 74 1005 32420 1006
rect 74 1004 32936 1005
rect 74 983 43128 1004
rect 74 888 99 983
rect 189 981 43128 983
rect 189 978 21772 981
rect 189 888 10618 978
rect 74 883 10618 888
rect 10708 977 21772 978
rect 10708 883 10807 977
rect 74 882 10807 883
rect 10897 972 21772 977
rect 10897 882 21326 972
rect 74 877 21326 882
rect 21416 886 21772 972
rect 21862 976 43128 981
rect 21862 886 32291 976
rect 21416 881 32291 886
rect 32381 975 43128 976
rect 32381 881 32480 975
rect 21416 880 32480 881
rect 32570 970 43128 975
rect 32570 880 42999 970
rect 21416 877 42999 880
rect 74 875 42999 877
rect 43089 875 43128 970
rect 74 858 43128 875
rect 10307 856 43128 858
rect 10307 852 21912 856
rect 10307 851 11263 852
rect 10586 512 10695 851
rect 10586 479 10611 512
rect 10647 479 10695 512
rect 10586 466 10695 479
rect 21222 847 21912 852
rect 31980 850 43128 856
rect 31980 849 32936 850
rect 21222 499 21364 847
rect 21222 466 21248 499
rect 21284 466 21364 499
rect 21222 453 21364 466
rect 32259 510 32368 849
rect 32259 477 32284 510
rect 32320 477 32368 510
rect 32259 464 32368 477
rect -33 -16 19411 12
rect -33 -98 19210 -16
rect 19368 -98 19411 -16
rect -33 -107 19411 -98
<< labels >>
rlabel metal1 1824 14158 1877 14180 1 d1
rlabel metal1 778 14176 840 14203 1 d0
rlabel metal2 123 14161 219 14194 1 vdd
rlabel metal1 299 14161 395 14194 1 gnd
rlabel locali 563 14172 607 14194 1 vref
rlabel metal1 4372 14499 4407 14513 1 d4
rlabel metal1 3110 14454 3162 14473 1 d3
rlabel metal1 2934 14471 2984 14484 1 d2
rlabel metal1 5421 14474 5491 14518 1 d5
rlabel metal1 18 266 49 325 1 d6
rlabel metal2 6 -82 79 -4 1 d7
rlabel metal1 21820 -165 21844 -153 1 vout
<< end >>
