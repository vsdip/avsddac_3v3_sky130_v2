magic
tech sky130A
timestamp 1633150163
<< nwell >>
rect 749 2566 1560 2790
rect 1797 2562 2608 2786
rect 749 1887 1560 2111
rect 2892 1882 3703 2106
rect 749 1119 1560 1343
rect 1797 1115 2608 1339
rect 749 440 1560 664
<< nmos >>
rect 813 2465 863 2507
rect 1026 2465 1076 2507
rect 1234 2465 1284 2507
rect 1442 2465 1492 2507
rect 1861 2461 1911 2503
rect 2074 2461 2124 2503
rect 2282 2461 2332 2503
rect 2490 2461 2540 2503
rect 813 1786 863 1828
rect 1026 1786 1076 1828
rect 1234 1786 1284 1828
rect 1442 1786 1492 1828
rect 2956 1781 3006 1823
rect 3169 1781 3219 1823
rect 3377 1781 3427 1823
rect 3585 1781 3635 1823
rect 813 1018 863 1060
rect 1026 1018 1076 1060
rect 1234 1018 1284 1060
rect 1442 1018 1492 1060
rect 1861 1014 1911 1056
rect 2074 1014 2124 1056
rect 2282 1014 2332 1056
rect 2490 1014 2540 1056
rect 813 339 863 381
rect 1026 339 1076 381
rect 1234 339 1284 381
rect 1442 339 1492 381
<< pmos >>
rect 813 2584 863 2684
rect 1026 2584 1076 2684
rect 1234 2584 1284 2684
rect 1442 2584 1492 2684
rect 1861 2580 1911 2680
rect 2074 2580 2124 2680
rect 2282 2580 2332 2680
rect 2490 2580 2540 2680
rect 813 1905 863 2005
rect 1026 1905 1076 2005
rect 1234 1905 1284 2005
rect 1442 1905 1492 2005
rect 2956 1900 3006 2000
rect 3169 1900 3219 2000
rect 3377 1900 3427 2000
rect 3585 1900 3635 2000
rect 813 1137 863 1237
rect 1026 1137 1076 1237
rect 1234 1137 1284 1237
rect 1442 1137 1492 1237
rect 1861 1133 1911 1233
rect 2074 1133 2124 1233
rect 2282 1133 2332 1233
rect 2490 1133 2540 1233
rect 813 458 863 558
rect 1026 458 1076 558
rect 1234 458 1284 558
rect 1442 458 1492 558
<< ndiff >>
rect 764 2497 813 2507
rect 764 2477 775 2497
rect 795 2477 813 2497
rect 764 2465 813 2477
rect 863 2501 907 2507
rect 863 2481 878 2501
rect 898 2481 907 2501
rect 863 2465 907 2481
rect 977 2497 1026 2507
rect 977 2477 988 2497
rect 1008 2477 1026 2497
rect 977 2465 1026 2477
rect 1076 2501 1120 2507
rect 1076 2481 1091 2501
rect 1111 2481 1120 2501
rect 1076 2465 1120 2481
rect 1185 2497 1234 2507
rect 1185 2477 1196 2497
rect 1216 2477 1234 2497
rect 1185 2465 1234 2477
rect 1284 2501 1328 2507
rect 1284 2481 1299 2501
rect 1319 2481 1328 2501
rect 1284 2465 1328 2481
rect 1398 2501 1442 2507
rect 1398 2481 1407 2501
rect 1427 2481 1442 2501
rect 1398 2465 1442 2481
rect 1492 2497 1541 2507
rect 1492 2477 1510 2497
rect 1530 2477 1541 2497
rect 1492 2465 1541 2477
rect 1812 2493 1861 2503
rect 1812 2473 1823 2493
rect 1843 2473 1861 2493
rect 1812 2461 1861 2473
rect 1911 2497 1955 2503
rect 1911 2477 1926 2497
rect 1946 2477 1955 2497
rect 1911 2461 1955 2477
rect 2025 2493 2074 2503
rect 2025 2473 2036 2493
rect 2056 2473 2074 2493
rect 2025 2461 2074 2473
rect 2124 2497 2168 2503
rect 2124 2477 2139 2497
rect 2159 2477 2168 2497
rect 2124 2461 2168 2477
rect 2233 2493 2282 2503
rect 2233 2473 2244 2493
rect 2264 2473 2282 2493
rect 2233 2461 2282 2473
rect 2332 2497 2376 2503
rect 2332 2477 2347 2497
rect 2367 2477 2376 2497
rect 2332 2461 2376 2477
rect 2446 2497 2490 2503
rect 2446 2477 2455 2497
rect 2475 2477 2490 2497
rect 2446 2461 2490 2477
rect 2540 2493 2589 2503
rect 2540 2473 2558 2493
rect 2578 2473 2589 2493
rect 2540 2461 2589 2473
rect 764 1818 813 1828
rect 764 1798 775 1818
rect 795 1798 813 1818
rect 764 1786 813 1798
rect 863 1822 907 1828
rect 863 1802 878 1822
rect 898 1802 907 1822
rect 863 1786 907 1802
rect 977 1818 1026 1828
rect 977 1798 988 1818
rect 1008 1798 1026 1818
rect 977 1786 1026 1798
rect 1076 1822 1120 1828
rect 1076 1802 1091 1822
rect 1111 1802 1120 1822
rect 1076 1786 1120 1802
rect 1185 1818 1234 1828
rect 1185 1798 1196 1818
rect 1216 1798 1234 1818
rect 1185 1786 1234 1798
rect 1284 1822 1328 1828
rect 1284 1802 1299 1822
rect 1319 1802 1328 1822
rect 1284 1786 1328 1802
rect 1398 1822 1442 1828
rect 1398 1802 1407 1822
rect 1427 1802 1442 1822
rect 1398 1786 1442 1802
rect 1492 1818 1541 1828
rect 1492 1798 1510 1818
rect 1530 1798 1541 1818
rect 1492 1786 1541 1798
rect 2907 1813 2956 1823
rect 2907 1793 2918 1813
rect 2938 1793 2956 1813
rect 2907 1781 2956 1793
rect 3006 1817 3050 1823
rect 3006 1797 3021 1817
rect 3041 1797 3050 1817
rect 3006 1781 3050 1797
rect 3120 1813 3169 1823
rect 3120 1793 3131 1813
rect 3151 1793 3169 1813
rect 3120 1781 3169 1793
rect 3219 1817 3263 1823
rect 3219 1797 3234 1817
rect 3254 1797 3263 1817
rect 3219 1781 3263 1797
rect 3328 1813 3377 1823
rect 3328 1793 3339 1813
rect 3359 1793 3377 1813
rect 3328 1781 3377 1793
rect 3427 1817 3471 1823
rect 3427 1797 3442 1817
rect 3462 1797 3471 1817
rect 3427 1781 3471 1797
rect 3541 1817 3585 1823
rect 3541 1797 3550 1817
rect 3570 1797 3585 1817
rect 3541 1781 3585 1797
rect 3635 1813 3684 1823
rect 3635 1793 3653 1813
rect 3673 1793 3684 1813
rect 3635 1781 3684 1793
rect 764 1050 813 1060
rect 764 1030 775 1050
rect 795 1030 813 1050
rect 764 1018 813 1030
rect 863 1054 907 1060
rect 863 1034 878 1054
rect 898 1034 907 1054
rect 863 1018 907 1034
rect 977 1050 1026 1060
rect 977 1030 988 1050
rect 1008 1030 1026 1050
rect 977 1018 1026 1030
rect 1076 1054 1120 1060
rect 1076 1034 1091 1054
rect 1111 1034 1120 1054
rect 1076 1018 1120 1034
rect 1185 1050 1234 1060
rect 1185 1030 1196 1050
rect 1216 1030 1234 1050
rect 1185 1018 1234 1030
rect 1284 1054 1328 1060
rect 1284 1034 1299 1054
rect 1319 1034 1328 1054
rect 1284 1018 1328 1034
rect 1398 1054 1442 1060
rect 1398 1034 1407 1054
rect 1427 1034 1442 1054
rect 1398 1018 1442 1034
rect 1492 1050 1541 1060
rect 1492 1030 1510 1050
rect 1530 1030 1541 1050
rect 1492 1018 1541 1030
rect 1812 1046 1861 1056
rect 1812 1026 1823 1046
rect 1843 1026 1861 1046
rect 1812 1014 1861 1026
rect 1911 1050 1955 1056
rect 1911 1030 1926 1050
rect 1946 1030 1955 1050
rect 1911 1014 1955 1030
rect 2025 1046 2074 1056
rect 2025 1026 2036 1046
rect 2056 1026 2074 1046
rect 2025 1014 2074 1026
rect 2124 1050 2168 1056
rect 2124 1030 2139 1050
rect 2159 1030 2168 1050
rect 2124 1014 2168 1030
rect 2233 1046 2282 1056
rect 2233 1026 2244 1046
rect 2264 1026 2282 1046
rect 2233 1014 2282 1026
rect 2332 1050 2376 1056
rect 2332 1030 2347 1050
rect 2367 1030 2376 1050
rect 2332 1014 2376 1030
rect 2446 1050 2490 1056
rect 2446 1030 2455 1050
rect 2475 1030 2490 1050
rect 2446 1014 2490 1030
rect 2540 1046 2589 1056
rect 2540 1026 2558 1046
rect 2578 1026 2589 1046
rect 2540 1014 2589 1026
rect 764 371 813 381
rect 764 351 775 371
rect 795 351 813 371
rect 764 339 813 351
rect 863 375 907 381
rect 863 355 878 375
rect 898 355 907 375
rect 863 339 907 355
rect 977 371 1026 381
rect 977 351 988 371
rect 1008 351 1026 371
rect 977 339 1026 351
rect 1076 375 1120 381
rect 1076 355 1091 375
rect 1111 355 1120 375
rect 1076 339 1120 355
rect 1185 371 1234 381
rect 1185 351 1196 371
rect 1216 351 1234 371
rect 1185 339 1234 351
rect 1284 375 1328 381
rect 1284 355 1299 375
rect 1319 355 1328 375
rect 1284 339 1328 355
rect 1398 375 1442 381
rect 1398 355 1407 375
rect 1427 355 1442 375
rect 1398 339 1442 355
rect 1492 371 1541 381
rect 1492 351 1510 371
rect 1530 351 1541 371
rect 1492 339 1541 351
<< pdiff >>
rect 769 2646 813 2684
rect 769 2626 781 2646
rect 801 2626 813 2646
rect 769 2584 813 2626
rect 863 2646 905 2684
rect 863 2626 877 2646
rect 897 2626 905 2646
rect 863 2584 905 2626
rect 982 2646 1026 2684
rect 982 2626 994 2646
rect 1014 2626 1026 2646
rect 982 2584 1026 2626
rect 1076 2646 1118 2684
rect 1076 2626 1090 2646
rect 1110 2626 1118 2646
rect 1076 2584 1118 2626
rect 1190 2646 1234 2684
rect 1190 2626 1202 2646
rect 1222 2626 1234 2646
rect 1190 2584 1234 2626
rect 1284 2646 1326 2684
rect 1284 2626 1298 2646
rect 1318 2626 1326 2646
rect 1284 2584 1326 2626
rect 1400 2646 1442 2684
rect 1400 2626 1408 2646
rect 1428 2626 1442 2646
rect 1400 2584 1442 2626
rect 1492 2653 1537 2684
rect 1492 2646 1536 2653
rect 1492 2626 1504 2646
rect 1524 2626 1536 2646
rect 1492 2584 1536 2626
rect 1817 2642 1861 2680
rect 1817 2622 1829 2642
rect 1849 2622 1861 2642
rect 1817 2580 1861 2622
rect 1911 2642 1953 2680
rect 1911 2622 1925 2642
rect 1945 2622 1953 2642
rect 1911 2580 1953 2622
rect 2030 2642 2074 2680
rect 2030 2622 2042 2642
rect 2062 2622 2074 2642
rect 2030 2580 2074 2622
rect 2124 2642 2166 2680
rect 2124 2622 2138 2642
rect 2158 2622 2166 2642
rect 2124 2580 2166 2622
rect 2238 2642 2282 2680
rect 2238 2622 2250 2642
rect 2270 2622 2282 2642
rect 2238 2580 2282 2622
rect 2332 2642 2374 2680
rect 2332 2622 2346 2642
rect 2366 2622 2374 2642
rect 2332 2580 2374 2622
rect 2448 2642 2490 2680
rect 2448 2622 2456 2642
rect 2476 2622 2490 2642
rect 2448 2580 2490 2622
rect 2540 2649 2585 2680
rect 2540 2642 2584 2649
rect 2540 2622 2552 2642
rect 2572 2622 2584 2642
rect 2540 2580 2584 2622
rect 769 1967 813 2005
rect 769 1947 781 1967
rect 801 1947 813 1967
rect 769 1905 813 1947
rect 863 1967 905 2005
rect 863 1947 877 1967
rect 897 1947 905 1967
rect 863 1905 905 1947
rect 982 1967 1026 2005
rect 982 1947 994 1967
rect 1014 1947 1026 1967
rect 982 1905 1026 1947
rect 1076 1967 1118 2005
rect 1076 1947 1090 1967
rect 1110 1947 1118 1967
rect 1076 1905 1118 1947
rect 1190 1967 1234 2005
rect 1190 1947 1202 1967
rect 1222 1947 1234 1967
rect 1190 1905 1234 1947
rect 1284 1967 1326 2005
rect 1284 1947 1298 1967
rect 1318 1947 1326 1967
rect 1284 1905 1326 1947
rect 1400 1967 1442 2005
rect 1400 1947 1408 1967
rect 1428 1947 1442 1967
rect 1400 1905 1442 1947
rect 1492 1974 1537 2005
rect 1492 1967 1536 1974
rect 1492 1947 1504 1967
rect 1524 1947 1536 1967
rect 1492 1905 1536 1947
rect 2912 1962 2956 2000
rect 2912 1942 2924 1962
rect 2944 1942 2956 1962
rect 2912 1900 2956 1942
rect 3006 1962 3048 2000
rect 3006 1942 3020 1962
rect 3040 1942 3048 1962
rect 3006 1900 3048 1942
rect 3125 1962 3169 2000
rect 3125 1942 3137 1962
rect 3157 1942 3169 1962
rect 3125 1900 3169 1942
rect 3219 1962 3261 2000
rect 3219 1942 3233 1962
rect 3253 1942 3261 1962
rect 3219 1900 3261 1942
rect 3333 1962 3377 2000
rect 3333 1942 3345 1962
rect 3365 1942 3377 1962
rect 3333 1900 3377 1942
rect 3427 1962 3469 2000
rect 3427 1942 3441 1962
rect 3461 1942 3469 1962
rect 3427 1900 3469 1942
rect 3543 1962 3585 2000
rect 3543 1942 3551 1962
rect 3571 1942 3585 1962
rect 3543 1900 3585 1942
rect 3635 1969 3680 2000
rect 3635 1962 3679 1969
rect 3635 1942 3647 1962
rect 3667 1942 3679 1962
rect 3635 1900 3679 1942
rect 769 1199 813 1237
rect 769 1179 781 1199
rect 801 1179 813 1199
rect 769 1137 813 1179
rect 863 1199 905 1237
rect 863 1179 877 1199
rect 897 1179 905 1199
rect 863 1137 905 1179
rect 982 1199 1026 1237
rect 982 1179 994 1199
rect 1014 1179 1026 1199
rect 982 1137 1026 1179
rect 1076 1199 1118 1237
rect 1076 1179 1090 1199
rect 1110 1179 1118 1199
rect 1076 1137 1118 1179
rect 1190 1199 1234 1237
rect 1190 1179 1202 1199
rect 1222 1179 1234 1199
rect 1190 1137 1234 1179
rect 1284 1199 1326 1237
rect 1284 1179 1298 1199
rect 1318 1179 1326 1199
rect 1284 1137 1326 1179
rect 1400 1199 1442 1237
rect 1400 1179 1408 1199
rect 1428 1179 1442 1199
rect 1400 1137 1442 1179
rect 1492 1206 1537 1237
rect 1492 1199 1536 1206
rect 1492 1179 1504 1199
rect 1524 1179 1536 1199
rect 1492 1137 1536 1179
rect 1817 1195 1861 1233
rect 1817 1175 1829 1195
rect 1849 1175 1861 1195
rect 1817 1133 1861 1175
rect 1911 1195 1953 1233
rect 1911 1175 1925 1195
rect 1945 1175 1953 1195
rect 1911 1133 1953 1175
rect 2030 1195 2074 1233
rect 2030 1175 2042 1195
rect 2062 1175 2074 1195
rect 2030 1133 2074 1175
rect 2124 1195 2166 1233
rect 2124 1175 2138 1195
rect 2158 1175 2166 1195
rect 2124 1133 2166 1175
rect 2238 1195 2282 1233
rect 2238 1175 2250 1195
rect 2270 1175 2282 1195
rect 2238 1133 2282 1175
rect 2332 1195 2374 1233
rect 2332 1175 2346 1195
rect 2366 1175 2374 1195
rect 2332 1133 2374 1175
rect 2448 1195 2490 1233
rect 2448 1175 2456 1195
rect 2476 1175 2490 1195
rect 2448 1133 2490 1175
rect 2540 1202 2585 1233
rect 2540 1195 2584 1202
rect 2540 1175 2552 1195
rect 2572 1175 2584 1195
rect 2540 1133 2584 1175
rect 769 520 813 558
rect 769 500 781 520
rect 801 500 813 520
rect 769 458 813 500
rect 863 520 905 558
rect 863 500 877 520
rect 897 500 905 520
rect 863 458 905 500
rect 982 520 1026 558
rect 982 500 994 520
rect 1014 500 1026 520
rect 982 458 1026 500
rect 1076 520 1118 558
rect 1076 500 1090 520
rect 1110 500 1118 520
rect 1076 458 1118 500
rect 1190 520 1234 558
rect 1190 500 1202 520
rect 1222 500 1234 520
rect 1190 458 1234 500
rect 1284 520 1326 558
rect 1284 500 1298 520
rect 1318 500 1326 520
rect 1284 458 1326 500
rect 1400 520 1442 558
rect 1400 500 1408 520
rect 1428 500 1442 520
rect 1400 458 1442 500
rect 1492 527 1537 558
rect 1492 520 1536 527
rect 1492 500 1504 520
rect 1524 500 1536 520
rect 1492 458 1536 500
<< ndiffc >>
rect 455 2800 473 2818
rect 457 2701 475 2719
rect 455 2544 473 2562
rect 775 2477 795 2497
rect 878 2481 898 2501
rect 988 2477 1008 2497
rect 1091 2481 1111 2501
rect 1196 2477 1216 2497
rect 1299 2481 1319 2501
rect 1407 2481 1427 2501
rect 1510 2477 1530 2497
rect 1823 2473 1843 2493
rect 457 2445 475 2463
rect 1926 2477 1946 2497
rect 2036 2473 2056 2493
rect 2139 2477 2159 2497
rect 2244 2473 2264 2493
rect 2347 2477 2367 2497
rect 2455 2477 2475 2497
rect 2558 2473 2578 2493
rect 455 2149 473 2167
rect 457 2050 475 2068
rect 455 1894 473 1912
rect 457 1795 475 1813
rect 775 1798 795 1818
rect 878 1802 898 1822
rect 988 1798 1008 1818
rect 1091 1802 1111 1822
rect 1196 1798 1216 1818
rect 1299 1802 1319 1822
rect 1407 1802 1427 1822
rect 1510 1798 1530 1818
rect 2918 1793 2938 1813
rect 3021 1797 3041 1817
rect 3131 1793 3151 1813
rect 3234 1797 3254 1817
rect 3339 1793 3359 1813
rect 3442 1797 3462 1817
rect 3550 1797 3570 1817
rect 3653 1793 3673 1813
rect 455 1353 473 1371
rect 457 1254 475 1272
rect 455 1097 473 1115
rect 775 1030 795 1050
rect 878 1034 898 1054
rect 988 1030 1008 1050
rect 1091 1034 1111 1054
rect 1196 1030 1216 1050
rect 1299 1034 1319 1054
rect 1407 1034 1427 1054
rect 1510 1030 1530 1050
rect 1823 1026 1843 1046
rect 457 998 475 1016
rect 1926 1030 1946 1050
rect 2036 1026 2056 1046
rect 2139 1030 2159 1050
rect 2244 1026 2264 1046
rect 2347 1030 2367 1050
rect 2455 1030 2475 1050
rect 2558 1026 2578 1046
rect 455 702 473 720
rect 457 603 475 621
rect 455 447 473 465
rect 457 348 475 366
rect 775 351 795 371
rect 878 355 898 375
rect 988 351 1008 371
rect 1091 355 1111 375
rect 1196 351 1216 371
rect 1299 355 1319 375
rect 1407 355 1427 375
rect 1510 351 1530 371
<< pdiffc >>
rect 781 2626 801 2646
rect 877 2626 897 2646
rect 994 2626 1014 2646
rect 1090 2626 1110 2646
rect 1202 2626 1222 2646
rect 1298 2626 1318 2646
rect 1408 2626 1428 2646
rect 1504 2626 1524 2646
rect 1829 2622 1849 2642
rect 1925 2622 1945 2642
rect 2042 2622 2062 2642
rect 2138 2622 2158 2642
rect 2250 2622 2270 2642
rect 2346 2622 2366 2642
rect 2456 2622 2476 2642
rect 2552 2622 2572 2642
rect 781 1947 801 1967
rect 877 1947 897 1967
rect 994 1947 1014 1967
rect 1090 1947 1110 1967
rect 1202 1947 1222 1967
rect 1298 1947 1318 1967
rect 1408 1947 1428 1967
rect 1504 1947 1524 1967
rect 2924 1942 2944 1962
rect 3020 1942 3040 1962
rect 3137 1942 3157 1962
rect 3233 1942 3253 1962
rect 3345 1942 3365 1962
rect 3441 1942 3461 1962
rect 3551 1942 3571 1962
rect 3647 1942 3667 1962
rect 781 1179 801 1199
rect 877 1179 897 1199
rect 994 1179 1014 1199
rect 1090 1179 1110 1199
rect 1202 1179 1222 1199
rect 1298 1179 1318 1199
rect 1408 1179 1428 1199
rect 1504 1179 1524 1199
rect 1829 1175 1849 1195
rect 1925 1175 1945 1195
rect 2042 1175 2062 1195
rect 2138 1175 2158 1195
rect 2250 1175 2270 1195
rect 2346 1175 2366 1195
rect 2456 1175 2476 1195
rect 2552 1175 2572 1195
rect 781 500 801 520
rect 877 500 897 520
rect 994 500 1014 520
rect 1090 500 1110 520
rect 1202 500 1222 520
rect 1298 500 1318 520
rect 1408 500 1428 520
rect 1504 500 1524 520
<< psubdiff >>
rect 849 2410 960 2424
rect 849 2380 890 2410
rect 918 2380 960 2410
rect 849 2365 960 2380
rect 1897 2406 2008 2420
rect 1897 2376 1938 2406
rect 1966 2376 2008 2406
rect 1897 2361 2008 2376
rect 849 1731 960 1745
rect 849 1701 890 1731
rect 918 1701 960 1731
rect 849 1688 960 1701
rect 2992 1726 3103 1740
rect 2992 1696 3033 1726
rect 3061 1696 3103 1726
rect 2992 1681 3103 1696
rect 849 963 960 977
rect 849 933 890 963
rect 918 933 960 963
rect 849 918 960 933
rect 1897 959 2008 973
rect 1897 929 1938 959
rect 1966 929 2008 959
rect 1897 914 2008 929
rect 849 284 960 298
rect 849 254 890 284
rect 918 254 960 284
rect 849 239 960 254
<< nsubdiff >>
rect 850 2757 960 2771
rect 850 2727 893 2757
rect 921 2727 960 2757
rect 850 2712 960 2727
rect 1898 2753 2008 2767
rect 1898 2723 1941 2753
rect 1969 2723 2008 2753
rect 1898 2708 2008 2723
rect 850 2078 960 2092
rect 850 2048 893 2078
rect 921 2048 960 2078
rect 850 2033 960 2048
rect 2993 2073 3103 2087
rect 2993 2043 3036 2073
rect 3064 2043 3103 2073
rect 2993 2028 3103 2043
rect 850 1310 960 1324
rect 850 1280 893 1310
rect 921 1280 960 1310
rect 850 1265 960 1280
rect 1898 1306 2008 1320
rect 1898 1276 1941 1306
rect 1969 1276 2008 1306
rect 1898 1261 2008 1276
rect 850 631 960 645
rect 850 601 893 631
rect 921 601 960 631
rect 850 586 960 601
<< psubdiffcont >>
rect 890 2380 918 2410
rect 1938 2376 1966 2406
rect 890 1701 918 1731
rect 3033 1696 3061 1726
rect 890 933 918 963
rect 1938 929 1966 959
rect 890 254 918 284
<< nsubdiffcont >>
rect 893 2727 921 2757
rect 1941 2723 1969 2753
rect 893 2048 921 2078
rect 3036 2043 3064 2073
rect 893 1280 921 1310
rect 1941 1276 1969 1306
rect 893 601 921 631
<< poly >>
rect 813 2684 863 2697
rect 1026 2684 1076 2697
rect 1234 2684 1284 2697
rect 1442 2684 1492 2697
rect 1861 2680 1911 2693
rect 2074 2680 2124 2693
rect 2282 2680 2332 2693
rect 2490 2680 2540 2693
rect 813 2556 863 2584
rect 813 2536 826 2556
rect 846 2536 863 2556
rect 813 2507 863 2536
rect 1026 2555 1076 2584
rect 1026 2531 1037 2555
rect 1061 2531 1076 2555
rect 1026 2507 1076 2531
rect 1234 2560 1284 2584
rect 1234 2536 1246 2560
rect 1270 2536 1284 2560
rect 1234 2507 1284 2536
rect 1442 2558 1492 2584
rect 1442 2532 1460 2558
rect 1486 2532 1492 2558
rect 1442 2507 1492 2532
rect 1861 2552 1911 2580
rect 1861 2532 1874 2552
rect 1894 2532 1911 2552
rect 1861 2503 1911 2532
rect 2074 2551 2124 2580
rect 2074 2527 2085 2551
rect 2109 2527 2124 2551
rect 2074 2503 2124 2527
rect 2282 2556 2332 2580
rect 2282 2532 2294 2556
rect 2318 2532 2332 2556
rect 2282 2503 2332 2532
rect 2490 2554 2540 2580
rect 2490 2528 2508 2554
rect 2534 2528 2540 2554
rect 2490 2503 2540 2528
rect 813 2449 863 2465
rect 1026 2449 1076 2465
rect 1234 2449 1284 2465
rect 1442 2449 1492 2465
rect 1861 2445 1911 2461
rect 2074 2445 2124 2461
rect 2282 2445 2332 2461
rect 2490 2445 2540 2461
rect 813 2005 863 2018
rect 1026 2005 1076 2018
rect 1234 2005 1284 2018
rect 1442 2005 1492 2018
rect 2956 2000 3006 2013
rect 3169 2000 3219 2013
rect 3377 2000 3427 2013
rect 3585 2000 3635 2013
rect 813 1877 863 1905
rect 813 1857 826 1877
rect 846 1857 863 1877
rect 813 1828 863 1857
rect 1026 1876 1076 1905
rect 1026 1852 1037 1876
rect 1061 1852 1076 1876
rect 1026 1828 1076 1852
rect 1234 1881 1284 1905
rect 1234 1857 1246 1881
rect 1270 1857 1284 1881
rect 1234 1828 1284 1857
rect 1442 1879 1492 1905
rect 1442 1853 1460 1879
rect 1486 1853 1492 1879
rect 1442 1828 1492 1853
rect 2956 1872 3006 1900
rect 2956 1852 2969 1872
rect 2989 1852 3006 1872
rect 2956 1823 3006 1852
rect 3169 1871 3219 1900
rect 3169 1847 3180 1871
rect 3204 1847 3219 1871
rect 3169 1823 3219 1847
rect 3377 1876 3427 1900
rect 3377 1852 3389 1876
rect 3413 1852 3427 1876
rect 3377 1823 3427 1852
rect 3585 1874 3635 1900
rect 3585 1848 3603 1874
rect 3629 1848 3635 1874
rect 3585 1823 3635 1848
rect 813 1770 863 1786
rect 1026 1770 1076 1786
rect 1234 1770 1284 1786
rect 1442 1770 1492 1786
rect 2956 1765 3006 1781
rect 3169 1765 3219 1781
rect 3377 1765 3427 1781
rect 3585 1765 3635 1781
rect 813 1237 863 1250
rect 1026 1237 1076 1250
rect 1234 1237 1284 1250
rect 1442 1237 1492 1250
rect 1861 1233 1911 1246
rect 2074 1233 2124 1246
rect 2282 1233 2332 1246
rect 2490 1233 2540 1246
rect 813 1109 863 1137
rect 813 1089 826 1109
rect 846 1089 863 1109
rect 813 1060 863 1089
rect 1026 1108 1076 1137
rect 1026 1084 1037 1108
rect 1061 1084 1076 1108
rect 1026 1060 1076 1084
rect 1234 1113 1284 1137
rect 1234 1089 1246 1113
rect 1270 1089 1284 1113
rect 1234 1060 1284 1089
rect 1442 1111 1492 1137
rect 1442 1085 1460 1111
rect 1486 1085 1492 1111
rect 1442 1060 1492 1085
rect 1861 1105 1911 1133
rect 1861 1085 1874 1105
rect 1894 1085 1911 1105
rect 1861 1056 1911 1085
rect 2074 1104 2124 1133
rect 2074 1080 2085 1104
rect 2109 1080 2124 1104
rect 2074 1056 2124 1080
rect 2282 1109 2332 1133
rect 2282 1085 2294 1109
rect 2318 1085 2332 1109
rect 2282 1056 2332 1085
rect 2490 1107 2540 1133
rect 2490 1081 2508 1107
rect 2534 1081 2540 1107
rect 2490 1056 2540 1081
rect 813 1002 863 1018
rect 1026 1002 1076 1018
rect 1234 1002 1284 1018
rect 1442 1002 1492 1018
rect 1861 998 1911 1014
rect 2074 998 2124 1014
rect 2282 998 2332 1014
rect 2490 998 2540 1014
rect 813 558 863 571
rect 1026 558 1076 571
rect 1234 558 1284 571
rect 1442 558 1492 571
rect 813 430 863 458
rect 813 410 826 430
rect 846 410 863 430
rect 813 381 863 410
rect 1026 429 1076 458
rect 1026 405 1037 429
rect 1061 405 1076 429
rect 1026 381 1076 405
rect 1234 434 1284 458
rect 1234 410 1246 434
rect 1270 410 1284 434
rect 1234 381 1284 410
rect 1442 432 1492 458
rect 1442 406 1460 432
rect 1486 406 1492 432
rect 1442 381 1492 406
rect 813 323 863 339
rect 1026 323 1076 339
rect 1234 323 1284 339
rect 1442 323 1492 339
<< polycont >>
rect 826 2536 846 2556
rect 1037 2531 1061 2555
rect 1246 2536 1270 2560
rect 1460 2532 1486 2558
rect 1874 2532 1894 2552
rect 2085 2527 2109 2551
rect 2294 2532 2318 2556
rect 2508 2528 2534 2554
rect 826 1857 846 1877
rect 1037 1852 1061 1876
rect 1246 1857 1270 1881
rect 1460 1853 1486 1879
rect 2969 1852 2989 1872
rect 3180 1847 3204 1871
rect 3389 1852 3413 1876
rect 3603 1848 3629 1874
rect 826 1089 846 1109
rect 1037 1084 1061 1108
rect 1246 1089 1270 1113
rect 1460 1085 1486 1111
rect 1874 1085 1894 1105
rect 2085 1080 2109 1104
rect 2294 1085 2318 1109
rect 2508 1081 2534 1107
rect 826 410 846 430
rect 1037 405 1061 429
rect 1246 410 1270 434
rect 1460 406 1486 432
<< ndiffres >>
rect 434 2818 491 2837
rect 434 2815 455 2818
rect 340 2800 455 2815
rect 473 2800 491 2818
rect 340 2777 491 2800
rect 340 2741 382 2777
rect 339 2740 439 2741
rect 339 2719 495 2740
rect 339 2701 457 2719
rect 475 2701 495 2719
rect 339 2697 495 2701
rect 434 2681 495 2697
rect 434 2562 491 2581
rect 434 2559 455 2562
rect 340 2544 455 2559
rect 473 2544 491 2562
rect 340 2521 491 2544
rect 340 2485 382 2521
rect 339 2484 439 2485
rect 339 2463 495 2484
rect 339 2445 457 2463
rect 475 2445 495 2463
rect 339 2441 495 2445
rect 434 2425 495 2441
rect 434 2167 491 2186
rect 434 2164 455 2167
rect 340 2149 455 2164
rect 473 2149 491 2167
rect 340 2126 491 2149
rect 340 2090 382 2126
rect 339 2089 439 2090
rect 339 2068 495 2089
rect 339 2050 457 2068
rect 475 2050 495 2068
rect 339 2046 495 2050
rect 434 2030 495 2046
rect 434 1912 491 1931
rect 434 1909 455 1912
rect 340 1894 455 1909
rect 473 1894 491 1912
rect 340 1871 491 1894
rect 340 1835 382 1871
rect 339 1834 439 1835
rect 339 1813 495 1834
rect 339 1795 457 1813
rect 475 1795 495 1813
rect 339 1791 495 1795
rect 434 1775 495 1791
rect 434 1371 491 1390
rect 434 1368 455 1371
rect 340 1353 455 1368
rect 473 1353 491 1371
rect 340 1330 491 1353
rect 340 1294 382 1330
rect 339 1293 439 1294
rect 339 1272 495 1293
rect 339 1254 457 1272
rect 475 1254 495 1272
rect 339 1250 495 1254
rect 434 1234 495 1250
rect 434 1115 491 1134
rect 434 1112 455 1115
rect 340 1097 455 1112
rect 473 1097 491 1115
rect 340 1074 491 1097
rect 340 1038 382 1074
rect 339 1037 439 1038
rect 339 1016 495 1037
rect 339 998 457 1016
rect 475 998 495 1016
rect 339 994 495 998
rect 434 978 495 994
rect 434 720 491 739
rect 434 717 455 720
rect 340 702 455 717
rect 473 702 491 720
rect 340 679 491 702
rect 340 643 382 679
rect 339 642 439 643
rect 339 621 495 642
rect 339 603 457 621
rect 475 603 495 621
rect 339 599 495 603
rect 434 583 495 599
rect 434 465 491 484
rect 434 462 455 465
rect 340 447 455 462
rect 473 447 491 465
rect 340 424 491 447
rect 340 388 382 424
rect 339 387 439 388
rect 339 366 495 387
rect 339 348 457 366
rect 475 348 495 366
rect 339 344 495 348
rect 434 328 495 344
<< locali >>
rect 433 2818 492 3008
rect 2810 2999 2875 3010
rect 2810 2951 2823 2999
rect 2860 2951 2875 2999
rect 2810 2938 2875 2951
rect 2396 2900 3062 2901
rect 1346 2899 1418 2900
rect 1345 2891 1444 2899
rect 1345 2888 1397 2891
rect 1345 2853 1353 2888
rect 1378 2853 1397 2888
rect 1422 2880 1444 2891
rect 2395 2893 3062 2900
rect 3335 2893 3378 2895
rect 2395 2892 3378 2893
rect 2395 2889 2447 2892
rect 1422 2879 2289 2880
rect 1422 2853 2290 2879
rect 1345 2843 2290 2853
rect 1345 2841 1444 2843
rect 433 2800 455 2818
rect 473 2800 492 2818
rect 433 2778 492 2800
rect 700 2814 1232 2819
rect 700 2794 1586 2814
rect 1606 2794 1609 2814
rect 2245 2810 2290 2843
rect 2395 2854 2403 2889
rect 2428 2854 2447 2889
rect 2472 2854 3378 2892
rect 2395 2845 3378 2854
rect 2395 2842 2484 2845
rect 700 2790 1609 2794
rect 700 2743 743 2790
rect 1193 2789 1609 2790
rect 2241 2790 2634 2810
rect 2654 2790 2657 2810
rect 1193 2788 1534 2789
rect 850 2757 960 2771
rect 850 2754 893 2757
rect 850 2749 854 2754
rect 688 2742 743 2743
rect 432 2719 743 2742
rect 432 2701 457 2719
rect 475 2707 743 2719
rect 772 2727 854 2749
rect 883 2727 893 2754
rect 921 2730 928 2757
rect 957 2749 960 2757
rect 957 2730 1022 2749
rect 921 2727 1022 2730
rect 772 2725 1022 2727
rect 475 2701 497 2707
rect 432 2562 497 2701
rect 772 2646 809 2725
rect 850 2712 960 2725
rect 924 2656 955 2657
rect 772 2626 781 2646
rect 801 2626 809 2646
rect 432 2544 455 2562
rect 473 2544 497 2562
rect 432 2527 497 2544
rect 652 2608 720 2621
rect 772 2616 809 2626
rect 868 2646 955 2656
rect 868 2626 877 2646
rect 897 2626 955 2646
rect 868 2617 955 2626
rect 868 2616 905 2617
rect 652 2566 659 2608
rect 708 2566 720 2608
rect 652 2563 720 2566
rect 924 2564 955 2617
rect 985 2646 1022 2725
rect 1137 2656 1168 2657
rect 985 2626 994 2646
rect 1014 2626 1022 2646
rect 985 2616 1022 2626
rect 1081 2649 1168 2656
rect 1081 2646 1142 2649
rect 1081 2626 1090 2646
rect 1110 2629 1142 2646
rect 1163 2629 1168 2649
rect 1110 2626 1168 2629
rect 1081 2619 1168 2626
rect 1193 2646 1230 2788
rect 1496 2787 1533 2788
rect 2241 2785 2657 2790
rect 2241 2784 2582 2785
rect 1898 2753 2008 2767
rect 1898 2750 1941 2753
rect 1898 2745 1902 2750
rect 1820 2723 1902 2745
rect 1931 2723 1941 2750
rect 1969 2726 1976 2753
rect 2005 2745 2008 2753
rect 2005 2726 2070 2745
rect 1969 2723 2070 2726
rect 1820 2721 2070 2723
rect 1345 2656 1381 2657
rect 1193 2626 1202 2646
rect 1222 2626 1230 2646
rect 1081 2617 1137 2619
rect 1081 2616 1118 2617
rect 1193 2616 1230 2626
rect 1289 2646 1437 2656
rect 1537 2653 1633 2655
rect 1289 2626 1298 2646
rect 1318 2626 1408 2646
rect 1428 2626 1437 2646
rect 1289 2620 1437 2626
rect 1289 2617 1353 2620
rect 1289 2616 1326 2617
rect 1345 2590 1353 2617
rect 1374 2617 1437 2620
rect 1495 2646 1633 2653
rect 1495 2626 1504 2646
rect 1524 2626 1633 2646
rect 1495 2617 1633 2626
rect 1820 2642 1857 2721
rect 1898 2708 2008 2721
rect 1972 2652 2003 2653
rect 1820 2622 1829 2642
rect 1849 2622 1857 2642
rect 1374 2590 1381 2617
rect 1400 2616 1437 2617
rect 1496 2616 1533 2617
rect 1345 2565 1381 2590
rect 816 2563 857 2564
rect 652 2556 857 2563
rect 652 2545 826 2556
rect 652 2512 660 2545
rect 653 2503 660 2512
rect 709 2536 826 2545
rect 846 2536 857 2556
rect 709 2528 857 2536
rect 924 2560 1283 2564
rect 924 2555 1246 2560
rect 924 2531 1037 2555
rect 1061 2536 1246 2555
rect 1270 2536 1283 2560
rect 1061 2531 1283 2536
rect 924 2528 1283 2531
rect 1345 2528 1380 2565
rect 1448 2562 1548 2565
rect 1448 2558 1515 2562
rect 1448 2532 1460 2558
rect 1486 2536 1515 2558
rect 1541 2536 1548 2562
rect 1486 2532 1548 2536
rect 1448 2528 1548 2532
rect 709 2512 720 2528
rect 709 2503 717 2512
rect 924 2507 955 2528
rect 1345 2507 1381 2528
rect 767 2506 804 2507
rect 432 2463 497 2482
rect 432 2445 457 2463
rect 475 2445 497 2463
rect 432 2244 497 2445
rect 653 2319 717 2503
rect 766 2497 804 2506
rect 766 2477 775 2497
rect 795 2477 804 2497
rect 766 2469 804 2477
rect 870 2501 955 2507
rect 980 2506 1017 2507
rect 870 2481 878 2501
rect 898 2481 955 2501
rect 870 2473 955 2481
rect 979 2497 1017 2506
rect 979 2477 988 2497
rect 1008 2477 1017 2497
rect 870 2472 906 2473
rect 979 2469 1017 2477
rect 1083 2501 1168 2507
rect 1188 2506 1225 2507
rect 1083 2481 1091 2501
rect 1111 2500 1168 2501
rect 1111 2481 1140 2500
rect 1083 2480 1140 2481
rect 1161 2480 1168 2500
rect 1083 2473 1168 2480
rect 1187 2497 1225 2506
rect 1187 2477 1196 2497
rect 1216 2477 1225 2497
rect 1083 2472 1119 2473
rect 1187 2469 1225 2477
rect 1291 2501 1435 2507
rect 1291 2481 1299 2501
rect 1319 2481 1407 2501
rect 1427 2481 1435 2501
rect 1291 2473 1435 2481
rect 1291 2472 1327 2473
rect 1399 2472 1435 2473
rect 1501 2506 1538 2507
rect 1501 2505 1539 2506
rect 1501 2497 1565 2505
rect 1501 2477 1510 2497
rect 1530 2483 1565 2497
rect 1585 2483 1588 2503
rect 1530 2478 1588 2483
rect 1530 2477 1565 2478
rect 767 2440 804 2469
rect 768 2438 804 2440
rect 980 2438 1017 2469
rect 768 2416 1017 2438
rect 849 2410 960 2416
rect 849 2402 890 2410
rect 849 2382 857 2402
rect 876 2382 890 2402
rect 849 2380 890 2382
rect 918 2402 960 2410
rect 918 2382 934 2402
rect 953 2382 960 2402
rect 918 2380 960 2382
rect 849 2365 960 2380
rect 653 2309 721 2319
rect 653 2276 670 2309
rect 710 2276 721 2309
rect 653 2264 721 2276
rect 653 2262 717 2264
rect 1188 2245 1225 2469
rect 1501 2465 1565 2477
rect 1605 2247 1632 2617
rect 1820 2612 1857 2622
rect 1916 2642 2003 2652
rect 1916 2622 1925 2642
rect 1945 2622 2003 2642
rect 1916 2613 2003 2622
rect 1916 2612 1953 2613
rect 1696 2599 1766 2604
rect 1691 2593 1766 2599
rect 1691 2560 1699 2593
rect 1752 2560 1766 2593
rect 1972 2560 2003 2613
rect 2033 2642 2070 2721
rect 2185 2652 2216 2653
rect 2033 2622 2042 2642
rect 2062 2622 2070 2642
rect 2033 2612 2070 2622
rect 2129 2645 2216 2652
rect 2129 2642 2190 2645
rect 2129 2622 2138 2642
rect 2158 2625 2190 2642
rect 2211 2625 2216 2645
rect 2158 2622 2216 2625
rect 2129 2615 2216 2622
rect 2241 2642 2278 2784
rect 2544 2783 2581 2784
rect 2393 2652 2429 2653
rect 2241 2622 2250 2642
rect 2270 2622 2278 2642
rect 2129 2613 2185 2615
rect 2129 2612 2166 2613
rect 2241 2612 2278 2622
rect 2337 2642 2485 2652
rect 2585 2649 2681 2651
rect 2337 2622 2346 2642
rect 2366 2622 2456 2642
rect 2476 2622 2485 2642
rect 2337 2616 2485 2622
rect 2337 2613 2401 2616
rect 2337 2612 2374 2613
rect 2393 2586 2401 2613
rect 2422 2613 2485 2616
rect 2543 2642 2681 2649
rect 2543 2622 2552 2642
rect 2572 2622 2681 2642
rect 2543 2613 2681 2622
rect 2422 2586 2429 2613
rect 2448 2612 2485 2613
rect 2544 2612 2581 2613
rect 2393 2561 2429 2586
rect 1691 2559 1774 2560
rect 1864 2559 1905 2560
rect 1691 2552 1905 2559
rect 1691 2535 1874 2552
rect 1691 2502 1704 2535
rect 1757 2532 1874 2535
rect 1894 2532 1905 2552
rect 1757 2524 1905 2532
rect 1972 2556 2331 2560
rect 1972 2551 2294 2556
rect 1972 2527 2085 2551
rect 2109 2532 2294 2551
rect 2318 2532 2331 2556
rect 2109 2527 2331 2532
rect 1972 2524 2331 2527
rect 2393 2524 2428 2561
rect 2496 2558 2596 2561
rect 2496 2554 2563 2558
rect 2496 2528 2508 2554
rect 2534 2532 2563 2554
rect 2589 2532 2596 2558
rect 2534 2528 2596 2532
rect 2496 2524 2596 2528
rect 1757 2502 1774 2524
rect 1972 2503 2003 2524
rect 2393 2503 2429 2524
rect 1815 2502 1852 2503
rect 1691 2488 1774 2502
rect 1464 2245 1632 2247
rect 1188 2244 1632 2245
rect 432 2214 1632 2244
rect 1702 2278 1774 2488
rect 1814 2493 1852 2502
rect 1814 2473 1823 2493
rect 1843 2473 1852 2493
rect 1814 2465 1852 2473
rect 1918 2497 2003 2503
rect 2028 2502 2065 2503
rect 1918 2477 1926 2497
rect 1946 2477 2003 2497
rect 1918 2469 2003 2477
rect 2027 2493 2065 2502
rect 2027 2473 2036 2493
rect 2056 2473 2065 2493
rect 1918 2468 1954 2469
rect 2027 2465 2065 2473
rect 2131 2497 2216 2503
rect 2236 2502 2273 2503
rect 2131 2477 2139 2497
rect 2159 2496 2216 2497
rect 2159 2477 2188 2496
rect 2131 2476 2188 2477
rect 2209 2476 2216 2496
rect 2131 2469 2216 2476
rect 2235 2493 2273 2502
rect 2235 2473 2244 2493
rect 2264 2473 2273 2493
rect 2131 2468 2167 2469
rect 2235 2465 2273 2473
rect 2339 2497 2483 2503
rect 2339 2477 2347 2497
rect 2367 2477 2455 2497
rect 2475 2477 2483 2497
rect 2339 2469 2483 2477
rect 2339 2468 2375 2469
rect 2447 2468 2483 2469
rect 2549 2502 2586 2503
rect 2549 2501 2587 2502
rect 2549 2493 2613 2501
rect 2549 2473 2558 2493
rect 2578 2479 2613 2493
rect 2633 2479 2636 2499
rect 2578 2474 2636 2479
rect 2578 2473 2613 2474
rect 1815 2436 1852 2465
rect 1816 2434 1852 2436
rect 2028 2434 2065 2465
rect 1816 2412 2065 2434
rect 1897 2406 2008 2412
rect 1897 2398 1938 2406
rect 1897 2378 1905 2398
rect 1924 2378 1938 2398
rect 1897 2376 1938 2378
rect 1966 2398 2008 2406
rect 1966 2378 1982 2398
rect 2001 2378 2008 2398
rect 1966 2376 2008 2378
rect 1897 2361 2008 2376
rect 1702 2239 1721 2278
rect 1766 2239 1774 2278
rect 1702 2222 1774 2239
rect 2236 2266 2273 2465
rect 2549 2461 2613 2473
rect 2236 2260 2277 2266
rect 2653 2262 2680 2613
rect 2811 2578 2875 2597
rect 2811 2539 2824 2578
rect 2858 2539 2875 2578
rect 2811 2520 2875 2539
rect 2512 2260 2680 2262
rect 2236 2234 2680 2260
rect 432 2167 497 2214
rect 432 2149 455 2167
rect 473 2149 497 2167
rect 1345 2194 1380 2196
rect 1345 2192 1449 2194
rect 2238 2192 2277 2234
rect 2512 2233 2680 2234
rect 1345 2185 2279 2192
rect 1345 2184 1396 2185
rect 1345 2164 1348 2184
rect 1373 2165 1396 2184
rect 1428 2165 2279 2185
rect 1373 2164 2279 2165
rect 1345 2157 2279 2164
rect 1618 2156 2279 2157
rect 432 2128 497 2149
rect 709 2139 749 2142
rect 709 2135 1612 2139
rect 709 2115 1586 2135
rect 1606 2115 1612 2135
rect 709 2112 1612 2115
rect 433 2068 498 2088
rect 433 2050 457 2068
rect 475 2050 498 2068
rect 433 2023 498 2050
rect 709 2023 749 2112
rect 1193 2110 1609 2112
rect 1193 2109 1534 2110
rect 850 2078 960 2092
rect 850 2075 893 2078
rect 850 2070 854 2075
rect 432 1988 749 2023
rect 772 2048 854 2070
rect 883 2048 893 2075
rect 921 2051 928 2078
rect 957 2070 960 2078
rect 957 2051 1022 2070
rect 921 2048 1022 2051
rect 772 2046 1022 2048
rect 433 1912 498 1988
rect 772 1967 809 2046
rect 850 2033 960 2046
rect 924 1977 955 1978
rect 772 1947 781 1967
rect 801 1947 809 1967
rect 772 1937 809 1947
rect 868 1967 955 1977
rect 868 1947 877 1967
rect 897 1947 955 1967
rect 868 1938 955 1947
rect 868 1937 905 1938
rect 433 1894 455 1912
rect 473 1894 498 1912
rect 433 1873 498 1894
rect 646 1892 711 1901
rect 646 1855 656 1892
rect 696 1884 711 1892
rect 924 1885 955 1938
rect 985 1967 1022 2046
rect 1137 1977 1168 1978
rect 985 1947 994 1967
rect 1014 1947 1022 1967
rect 985 1937 1022 1947
rect 1081 1970 1168 1977
rect 1081 1967 1142 1970
rect 1081 1947 1090 1967
rect 1110 1950 1142 1967
rect 1163 1950 1168 1970
rect 1110 1947 1168 1950
rect 1081 1940 1168 1947
rect 1193 1967 1230 2109
rect 1496 2108 1533 2109
rect 1345 1977 1381 1978
rect 1193 1947 1202 1967
rect 1222 1947 1230 1967
rect 1081 1938 1137 1940
rect 1081 1937 1118 1938
rect 1193 1937 1230 1947
rect 1289 1967 1437 1977
rect 1537 1974 1633 1976
rect 1289 1947 1298 1967
rect 1318 1947 1408 1967
rect 1428 1947 1437 1967
rect 1289 1941 1437 1947
rect 1289 1938 1353 1941
rect 1289 1937 1326 1938
rect 1345 1911 1353 1938
rect 1374 1938 1437 1941
rect 1495 1967 1633 1974
rect 1495 1947 1504 1967
rect 1524 1947 1633 1967
rect 1495 1938 1633 1947
rect 1374 1911 1381 1938
rect 1400 1937 1437 1938
rect 1496 1937 1533 1938
rect 1345 1886 1381 1911
rect 816 1884 857 1885
rect 696 1877 857 1884
rect 696 1857 826 1877
rect 846 1857 857 1877
rect 696 1855 857 1857
rect 646 1849 857 1855
rect 924 1881 1283 1885
rect 924 1876 1246 1881
rect 924 1852 1037 1876
rect 1061 1857 1246 1876
rect 1270 1857 1283 1881
rect 1061 1852 1283 1857
rect 924 1849 1283 1852
rect 1345 1849 1380 1886
rect 1448 1883 1548 1886
rect 1448 1879 1515 1883
rect 1448 1853 1460 1879
rect 1486 1857 1515 1879
rect 1541 1857 1548 1883
rect 1486 1853 1548 1857
rect 1448 1849 1548 1853
rect 646 1836 713 1849
rect 438 1813 494 1833
rect 438 1795 457 1813
rect 475 1795 494 1813
rect 438 1682 494 1795
rect 646 1815 660 1836
rect 696 1815 713 1836
rect 924 1828 955 1849
rect 1345 1828 1381 1849
rect 767 1827 804 1828
rect 646 1808 713 1815
rect 766 1818 804 1827
rect 438 1544 493 1682
rect 646 1656 711 1808
rect 766 1798 775 1818
rect 795 1798 804 1818
rect 766 1790 804 1798
rect 870 1822 955 1828
rect 980 1827 1017 1828
rect 870 1802 878 1822
rect 898 1802 955 1822
rect 870 1794 955 1802
rect 979 1818 1017 1827
rect 979 1798 988 1818
rect 1008 1798 1017 1818
rect 870 1793 906 1794
rect 979 1790 1017 1798
rect 1083 1822 1168 1828
rect 1188 1827 1225 1828
rect 1083 1802 1091 1822
rect 1111 1821 1168 1822
rect 1111 1802 1140 1821
rect 1083 1801 1140 1802
rect 1161 1801 1168 1821
rect 1083 1794 1168 1801
rect 1187 1818 1225 1827
rect 1187 1798 1196 1818
rect 1216 1798 1225 1818
rect 1083 1793 1119 1794
rect 1187 1790 1225 1798
rect 1291 1822 1435 1828
rect 1291 1802 1299 1822
rect 1319 1802 1407 1822
rect 1427 1802 1435 1822
rect 1291 1794 1435 1802
rect 1291 1793 1327 1794
rect 1399 1793 1435 1794
rect 1501 1827 1538 1828
rect 1501 1826 1539 1827
rect 1501 1818 1565 1826
rect 1501 1798 1510 1818
rect 1530 1804 1565 1818
rect 1585 1804 1588 1824
rect 1530 1799 1588 1804
rect 1530 1798 1565 1799
rect 767 1761 804 1790
rect 768 1759 804 1761
rect 980 1759 1017 1790
rect 768 1737 1017 1759
rect 849 1731 960 1737
rect 849 1723 890 1731
rect 849 1703 857 1723
rect 876 1703 890 1723
rect 849 1701 890 1703
rect 918 1723 960 1731
rect 918 1703 934 1723
rect 953 1703 960 1723
rect 918 1701 960 1703
rect 849 1688 960 1701
rect 1188 1691 1225 1790
rect 1501 1786 1565 1798
rect 639 1646 760 1656
rect 639 1644 708 1646
rect 639 1603 652 1644
rect 689 1605 708 1644
rect 745 1605 760 1646
rect 689 1603 760 1605
rect 639 1585 760 1603
rect 431 1541 495 1544
rect 851 1541 955 1547
rect 1186 1541 1227 1691
rect 1605 1683 1632 1938
rect 1694 1928 1774 1939
rect 1694 1902 1711 1928
rect 1751 1902 1774 1928
rect 1694 1875 1774 1902
rect 1694 1849 1715 1875
rect 1755 1849 1774 1875
rect 1694 1830 1774 1849
rect 2813 1879 2875 2520
rect 3335 2130 3378 2845
rect 3489 2200 3526 2221
rect 3489 2163 3500 2200
rect 3517 2163 3526 2200
rect 3489 2153 3526 2163
rect 3335 2110 3729 2130
rect 3749 2110 3752 2130
rect 3336 2105 3752 2110
rect 3336 2104 3677 2105
rect 2993 2073 3103 2087
rect 2993 2070 3036 2073
rect 2993 2065 2997 2070
rect 2915 2043 2997 2065
rect 3026 2043 3036 2070
rect 3064 2046 3071 2073
rect 3100 2065 3103 2073
rect 3100 2046 3165 2065
rect 3064 2043 3165 2046
rect 2915 2041 3165 2043
rect 2915 1962 2952 2041
rect 2993 2028 3103 2041
rect 3067 1972 3098 1973
rect 2915 1942 2924 1962
rect 2944 1942 2952 1962
rect 2915 1932 2952 1942
rect 3011 1962 3098 1972
rect 3011 1942 3020 1962
rect 3040 1942 3098 1962
rect 3011 1933 3098 1942
rect 3011 1932 3048 1933
rect 3067 1880 3098 1933
rect 3128 1962 3165 2041
rect 3280 1972 3311 1973
rect 3128 1942 3137 1962
rect 3157 1942 3165 1962
rect 3128 1932 3165 1942
rect 3224 1965 3311 1972
rect 3224 1962 3285 1965
rect 3224 1942 3233 1962
rect 3253 1945 3285 1962
rect 3306 1945 3311 1965
rect 3253 1942 3311 1945
rect 3224 1935 3311 1942
rect 3336 1962 3373 2104
rect 3639 2103 3676 2104
rect 3488 1972 3524 1973
rect 3336 1942 3345 1962
rect 3365 1942 3373 1962
rect 3224 1933 3280 1935
rect 3224 1932 3261 1933
rect 3336 1932 3373 1942
rect 3432 1962 3580 1972
rect 3680 1969 3776 1971
rect 3432 1942 3441 1962
rect 3461 1942 3551 1962
rect 3571 1942 3580 1962
rect 3432 1936 3580 1942
rect 3432 1933 3496 1936
rect 3432 1932 3469 1933
rect 3488 1906 3496 1933
rect 3517 1933 3580 1936
rect 3638 1962 3776 1969
rect 3638 1942 3647 1962
rect 3667 1942 3776 1962
rect 3638 1933 3776 1942
rect 3517 1906 3524 1933
rect 3543 1932 3580 1933
rect 3639 1932 3676 1933
rect 3488 1881 3524 1906
rect 2959 1879 3000 1880
rect 2813 1872 3000 1879
rect 2813 1852 2969 1872
rect 2989 1852 3000 1872
rect 2813 1846 3000 1852
rect 2851 1844 3000 1846
rect 3067 1876 3426 1880
rect 3067 1871 3389 1876
rect 3067 1847 3180 1871
rect 3204 1852 3389 1871
rect 3413 1852 3426 1876
rect 3204 1847 3426 1852
rect 3067 1844 3426 1847
rect 3488 1844 3523 1881
rect 3591 1878 3691 1881
rect 3591 1874 3658 1878
rect 3591 1848 3603 1874
rect 3629 1852 3658 1874
rect 3684 1852 3691 1878
rect 3629 1848 3691 1852
rect 3591 1844 3691 1848
rect 1694 1804 1718 1830
rect 1758 1804 1774 1830
rect 3067 1823 3098 1844
rect 3488 1823 3524 1844
rect 2910 1822 2947 1823
rect 1694 1753 1774 1804
rect 2909 1813 2947 1822
rect 2909 1793 2918 1813
rect 2938 1793 2947 1813
rect 2909 1785 2947 1793
rect 3013 1817 3098 1823
rect 3123 1822 3160 1823
rect 3013 1797 3021 1817
rect 3041 1797 3098 1817
rect 3013 1789 3098 1797
rect 3122 1813 3160 1822
rect 3122 1793 3131 1813
rect 3151 1793 3160 1813
rect 3013 1788 3049 1789
rect 3122 1785 3160 1793
rect 3226 1817 3311 1823
rect 3331 1822 3368 1823
rect 3226 1797 3234 1817
rect 3254 1816 3311 1817
rect 3254 1797 3283 1816
rect 3226 1796 3283 1797
rect 3304 1796 3311 1816
rect 3226 1789 3311 1796
rect 3330 1813 3368 1822
rect 3330 1793 3339 1813
rect 3359 1793 3368 1813
rect 3226 1788 3262 1789
rect 3330 1785 3368 1793
rect 3434 1817 3578 1823
rect 3434 1797 3442 1817
rect 3462 1797 3550 1817
rect 3570 1797 3578 1817
rect 3434 1789 3578 1797
rect 3434 1788 3470 1789
rect 3542 1788 3578 1789
rect 3644 1822 3681 1823
rect 3644 1821 3682 1822
rect 3644 1813 3708 1821
rect 3644 1793 3653 1813
rect 3673 1799 3708 1813
rect 3728 1799 3731 1819
rect 3673 1794 3731 1799
rect 3673 1793 3708 1794
rect 2910 1756 2947 1785
rect 2911 1754 2947 1756
rect 3123 1754 3160 1785
rect 431 1538 1227 1541
rect 1606 1552 1632 1683
rect 1606 1538 1634 1552
rect 431 1503 1634 1538
rect 1696 1545 1766 1753
rect 2911 1732 3160 1754
rect 2992 1726 3103 1732
rect 2992 1718 3033 1726
rect 2992 1698 3000 1718
rect 3019 1698 3033 1718
rect 2992 1696 3033 1698
rect 3061 1718 3103 1726
rect 3061 1698 3077 1718
rect 3096 1698 3103 1718
rect 3061 1696 3103 1698
rect 2992 1681 3103 1696
rect 3331 1670 3368 1785
rect 3644 1781 3708 1793
rect 431 1442 495 1503
rect 851 1501 955 1503
rect 1186 1501 1227 1503
rect 1696 1500 1717 1545
rect 1697 1479 1717 1500
rect 1747 1500 1766 1545
rect 3324 1664 3371 1670
rect 3748 1666 3775 1933
rect 3607 1664 3775 1666
rect 3324 1638 3775 1664
rect 1747 1479 1764 1500
rect 1697 1460 1764 1479
rect 2396 1453 2468 1454
rect 1346 1452 1418 1453
rect 1345 1444 1444 1452
rect 433 1371 492 1442
rect 1345 1441 1397 1444
rect 1345 1406 1353 1441
rect 1378 1406 1397 1441
rect 1422 1433 1444 1444
rect 2395 1445 2484 1453
rect 2395 1442 2447 1445
rect 1422 1432 2289 1433
rect 1422 1406 2290 1432
rect 1345 1396 2290 1406
rect 1345 1394 1444 1396
rect 433 1353 455 1371
rect 473 1353 492 1371
rect 433 1331 492 1353
rect 700 1367 1232 1372
rect 700 1347 1586 1367
rect 1606 1347 1609 1367
rect 2245 1363 2290 1396
rect 2395 1407 2403 1442
rect 2428 1407 2447 1442
rect 2472 1444 2484 1445
rect 3324 1444 3371 1638
rect 3607 1637 3775 1638
rect 2472 1407 3371 1444
rect 2395 1401 3371 1407
rect 2395 1397 3367 1401
rect 2395 1395 2484 1397
rect 700 1343 1609 1347
rect 700 1296 743 1343
rect 1193 1342 1609 1343
rect 2241 1343 2634 1363
rect 2654 1343 2657 1363
rect 1193 1341 1534 1342
rect 850 1310 960 1324
rect 850 1307 893 1310
rect 850 1302 854 1307
rect 688 1295 743 1296
rect 432 1272 743 1295
rect 432 1254 457 1272
rect 475 1260 743 1272
rect 772 1280 854 1302
rect 883 1280 893 1307
rect 921 1283 928 1310
rect 957 1302 960 1310
rect 957 1283 1022 1302
rect 921 1280 1022 1283
rect 772 1278 1022 1280
rect 475 1254 497 1260
rect 432 1115 497 1254
rect 772 1199 809 1278
rect 850 1265 960 1278
rect 924 1209 955 1210
rect 772 1179 781 1199
rect 801 1179 809 1199
rect 432 1097 455 1115
rect 473 1097 497 1115
rect 432 1080 497 1097
rect 652 1161 720 1174
rect 772 1169 809 1179
rect 868 1199 955 1209
rect 868 1179 877 1199
rect 897 1179 955 1199
rect 868 1170 955 1179
rect 868 1169 905 1170
rect 652 1119 659 1161
rect 708 1119 720 1161
rect 652 1116 720 1119
rect 924 1117 955 1170
rect 985 1199 1022 1278
rect 1137 1209 1168 1210
rect 985 1179 994 1199
rect 1014 1179 1022 1199
rect 985 1169 1022 1179
rect 1081 1202 1168 1209
rect 1081 1199 1142 1202
rect 1081 1179 1090 1199
rect 1110 1182 1142 1199
rect 1163 1182 1168 1202
rect 1110 1179 1168 1182
rect 1081 1172 1168 1179
rect 1193 1199 1230 1341
rect 1496 1340 1533 1341
rect 2241 1338 2657 1343
rect 2241 1337 2582 1338
rect 1898 1306 2008 1320
rect 1898 1303 1941 1306
rect 1898 1298 1902 1303
rect 1820 1276 1902 1298
rect 1931 1276 1941 1303
rect 1969 1279 1976 1306
rect 2005 1298 2008 1306
rect 2005 1279 2070 1298
rect 1969 1276 2070 1279
rect 1820 1274 2070 1276
rect 1345 1209 1381 1210
rect 1193 1179 1202 1199
rect 1222 1179 1230 1199
rect 1081 1170 1137 1172
rect 1081 1169 1118 1170
rect 1193 1169 1230 1179
rect 1289 1199 1437 1209
rect 1537 1206 1633 1208
rect 1289 1179 1298 1199
rect 1318 1179 1408 1199
rect 1428 1179 1437 1199
rect 1289 1173 1437 1179
rect 1289 1170 1353 1173
rect 1289 1169 1326 1170
rect 1345 1143 1353 1170
rect 1374 1170 1437 1173
rect 1495 1199 1633 1206
rect 1495 1179 1504 1199
rect 1524 1179 1633 1199
rect 1495 1170 1633 1179
rect 1820 1195 1857 1274
rect 1898 1261 2008 1274
rect 1972 1205 2003 1206
rect 1820 1175 1829 1195
rect 1849 1175 1857 1195
rect 1374 1143 1381 1170
rect 1400 1169 1437 1170
rect 1496 1169 1533 1170
rect 1345 1118 1381 1143
rect 816 1116 857 1117
rect 652 1109 857 1116
rect 652 1098 826 1109
rect 652 1065 660 1098
rect 653 1056 660 1065
rect 709 1089 826 1098
rect 846 1089 857 1109
rect 709 1081 857 1089
rect 924 1113 1283 1117
rect 924 1108 1246 1113
rect 924 1084 1037 1108
rect 1061 1089 1246 1108
rect 1270 1089 1283 1113
rect 1061 1084 1283 1089
rect 924 1081 1283 1084
rect 1345 1081 1380 1118
rect 1448 1115 1548 1118
rect 1448 1111 1515 1115
rect 1448 1085 1460 1111
rect 1486 1089 1515 1111
rect 1541 1089 1548 1115
rect 1486 1085 1548 1089
rect 1448 1081 1548 1085
rect 709 1065 720 1081
rect 709 1056 717 1065
rect 924 1060 955 1081
rect 1345 1060 1381 1081
rect 767 1059 804 1060
rect 432 1016 497 1035
rect 432 998 457 1016
rect 475 998 497 1016
rect 432 797 497 998
rect 653 872 717 1056
rect 766 1050 804 1059
rect 766 1030 775 1050
rect 795 1030 804 1050
rect 766 1022 804 1030
rect 870 1054 955 1060
rect 980 1059 1017 1060
rect 870 1034 878 1054
rect 898 1034 955 1054
rect 870 1026 955 1034
rect 979 1050 1017 1059
rect 979 1030 988 1050
rect 1008 1030 1017 1050
rect 870 1025 906 1026
rect 979 1022 1017 1030
rect 1083 1054 1168 1060
rect 1188 1059 1225 1060
rect 1083 1034 1091 1054
rect 1111 1053 1168 1054
rect 1111 1034 1140 1053
rect 1083 1033 1140 1034
rect 1161 1033 1168 1053
rect 1083 1026 1168 1033
rect 1187 1050 1225 1059
rect 1187 1030 1196 1050
rect 1216 1030 1225 1050
rect 1083 1025 1119 1026
rect 1187 1022 1225 1030
rect 1291 1054 1435 1060
rect 1291 1034 1299 1054
rect 1319 1034 1407 1054
rect 1427 1034 1435 1054
rect 1291 1026 1435 1034
rect 1291 1025 1327 1026
rect 1399 1025 1435 1026
rect 1501 1059 1538 1060
rect 1501 1058 1539 1059
rect 1501 1050 1565 1058
rect 1501 1030 1510 1050
rect 1530 1036 1565 1050
rect 1585 1036 1588 1056
rect 1530 1031 1588 1036
rect 1530 1030 1565 1031
rect 767 993 804 1022
rect 768 991 804 993
rect 980 991 1017 1022
rect 768 969 1017 991
rect 849 963 960 969
rect 849 955 890 963
rect 849 935 857 955
rect 876 935 890 955
rect 849 933 890 935
rect 918 955 960 963
rect 918 935 934 955
rect 953 935 960 955
rect 918 933 960 935
rect 849 918 960 933
rect 653 862 721 872
rect 653 829 670 862
rect 710 829 721 862
rect 653 817 721 829
rect 653 815 717 817
rect 1188 798 1225 1022
rect 1501 1018 1565 1030
rect 1605 800 1632 1170
rect 1820 1165 1857 1175
rect 1916 1195 2003 1205
rect 1916 1175 1925 1195
rect 1945 1175 2003 1195
rect 1916 1166 2003 1175
rect 1916 1165 1953 1166
rect 1696 1152 1766 1157
rect 1691 1146 1766 1152
rect 1691 1113 1699 1146
rect 1752 1113 1766 1146
rect 1972 1113 2003 1166
rect 2033 1195 2070 1274
rect 2185 1205 2216 1206
rect 2033 1175 2042 1195
rect 2062 1175 2070 1195
rect 2033 1165 2070 1175
rect 2129 1198 2216 1205
rect 2129 1195 2190 1198
rect 2129 1175 2138 1195
rect 2158 1178 2190 1195
rect 2211 1178 2216 1198
rect 2158 1175 2216 1178
rect 2129 1168 2216 1175
rect 2241 1195 2278 1337
rect 2544 1336 2581 1337
rect 2393 1205 2429 1206
rect 2241 1175 2250 1195
rect 2270 1175 2278 1195
rect 2129 1166 2185 1168
rect 2129 1165 2166 1166
rect 2241 1165 2278 1175
rect 2337 1195 2485 1205
rect 2585 1202 2681 1204
rect 2337 1175 2346 1195
rect 2366 1175 2456 1195
rect 2476 1175 2485 1195
rect 2337 1169 2485 1175
rect 2337 1166 2401 1169
rect 2337 1165 2374 1166
rect 2393 1139 2401 1166
rect 2422 1166 2485 1169
rect 2543 1195 2681 1202
rect 2543 1175 2552 1195
rect 2572 1175 2681 1195
rect 2543 1166 2681 1175
rect 2422 1139 2429 1166
rect 2448 1165 2485 1166
rect 2544 1165 2581 1166
rect 2393 1114 2429 1139
rect 1691 1112 1774 1113
rect 1864 1112 1905 1113
rect 1691 1105 1905 1112
rect 1691 1088 1874 1105
rect 1691 1055 1704 1088
rect 1757 1085 1874 1088
rect 1894 1085 1905 1105
rect 1757 1077 1905 1085
rect 1972 1109 2331 1113
rect 1972 1104 2294 1109
rect 1972 1080 2085 1104
rect 2109 1085 2294 1104
rect 2318 1085 2331 1109
rect 2109 1080 2331 1085
rect 1972 1077 2331 1080
rect 2393 1077 2428 1114
rect 2496 1111 2596 1114
rect 2496 1107 2563 1111
rect 2496 1081 2508 1107
rect 2534 1085 2563 1107
rect 2589 1085 2596 1111
rect 2534 1081 2596 1085
rect 2496 1077 2596 1081
rect 1757 1055 1774 1077
rect 1972 1056 2003 1077
rect 2393 1056 2429 1077
rect 1815 1055 1852 1056
rect 1691 1041 1774 1055
rect 1464 798 1632 800
rect 1188 797 1632 798
rect 432 767 1632 797
rect 1702 831 1774 1041
rect 1814 1046 1852 1055
rect 1814 1026 1823 1046
rect 1843 1026 1852 1046
rect 1814 1018 1852 1026
rect 1918 1050 2003 1056
rect 2028 1055 2065 1056
rect 1918 1030 1926 1050
rect 1946 1030 2003 1050
rect 1918 1022 2003 1030
rect 2027 1046 2065 1055
rect 2027 1026 2036 1046
rect 2056 1026 2065 1046
rect 1918 1021 1954 1022
rect 2027 1018 2065 1026
rect 2131 1050 2216 1056
rect 2236 1055 2273 1056
rect 2131 1030 2139 1050
rect 2159 1049 2216 1050
rect 2159 1030 2188 1049
rect 2131 1029 2188 1030
rect 2209 1029 2216 1049
rect 2131 1022 2216 1029
rect 2235 1046 2273 1055
rect 2235 1026 2244 1046
rect 2264 1026 2273 1046
rect 2131 1021 2167 1022
rect 2235 1018 2273 1026
rect 2339 1050 2483 1056
rect 2339 1030 2347 1050
rect 2367 1030 2455 1050
rect 2475 1030 2483 1050
rect 2339 1022 2483 1030
rect 2339 1021 2375 1022
rect 2447 1021 2483 1022
rect 2549 1055 2586 1056
rect 2549 1054 2587 1055
rect 2549 1046 2613 1054
rect 2549 1026 2558 1046
rect 2578 1032 2613 1046
rect 2633 1032 2636 1052
rect 2578 1027 2636 1032
rect 2578 1026 2613 1027
rect 1815 989 1852 1018
rect 1816 987 1852 989
rect 2028 987 2065 1018
rect 1816 965 2065 987
rect 1897 959 2008 965
rect 1897 951 1938 959
rect 1897 931 1905 951
rect 1924 931 1938 951
rect 1897 929 1938 931
rect 1966 951 2008 959
rect 1966 931 1982 951
rect 2001 931 2008 951
rect 1966 929 2008 931
rect 1897 914 2008 929
rect 1702 792 1721 831
rect 1766 792 1774 831
rect 1702 775 1774 792
rect 2236 819 2273 1018
rect 2549 1014 2613 1026
rect 2236 813 2277 819
rect 2653 815 2680 1166
rect 2512 813 2680 815
rect 2236 787 2680 813
rect 432 720 497 767
rect 432 702 455 720
rect 473 702 497 720
rect 1345 747 1380 749
rect 1345 745 1449 747
rect 2238 745 2277 787
rect 2512 786 2680 787
rect 1345 738 2279 745
rect 1345 737 1396 738
rect 1345 717 1348 737
rect 1373 718 1396 737
rect 1428 718 2279 738
rect 1373 717 2279 718
rect 1345 710 2279 717
rect 1618 709 2279 710
rect 432 681 497 702
rect 709 692 749 695
rect 709 688 1612 692
rect 709 668 1586 688
rect 1606 668 1612 688
rect 709 665 1612 668
rect 433 621 498 641
rect 433 603 457 621
rect 475 603 498 621
rect 433 576 498 603
rect 709 576 749 665
rect 1193 663 1609 665
rect 1193 662 1534 663
rect 850 631 960 645
rect 850 628 893 631
rect 850 623 854 628
rect 432 541 749 576
rect 772 601 854 623
rect 883 601 893 628
rect 921 604 928 631
rect 957 623 960 631
rect 957 604 1022 623
rect 921 601 1022 604
rect 772 599 1022 601
rect 433 465 498 541
rect 772 520 809 599
rect 850 586 960 599
rect 924 530 955 531
rect 772 500 781 520
rect 801 500 809 520
rect 772 490 809 500
rect 868 520 955 530
rect 868 500 877 520
rect 897 500 955 520
rect 868 491 955 500
rect 868 490 905 491
rect 433 447 455 465
rect 473 447 498 465
rect 433 426 498 447
rect 646 445 711 454
rect 646 408 656 445
rect 696 437 711 445
rect 924 438 955 491
rect 985 520 1022 599
rect 1137 530 1168 531
rect 985 500 994 520
rect 1014 500 1022 520
rect 985 490 1022 500
rect 1081 523 1168 530
rect 1081 520 1142 523
rect 1081 500 1090 520
rect 1110 503 1142 520
rect 1163 503 1168 523
rect 1110 500 1168 503
rect 1081 493 1168 500
rect 1193 520 1230 662
rect 1496 661 1533 662
rect 1345 530 1381 531
rect 1193 500 1202 520
rect 1222 500 1230 520
rect 1081 491 1137 493
rect 1081 490 1118 491
rect 1193 490 1230 500
rect 1289 520 1437 530
rect 1537 527 1633 529
rect 1289 500 1298 520
rect 1318 500 1408 520
rect 1428 500 1437 520
rect 1289 494 1437 500
rect 1289 491 1353 494
rect 1289 490 1326 491
rect 1345 464 1353 491
rect 1374 491 1437 494
rect 1495 520 1633 527
rect 1495 500 1504 520
rect 1524 500 1633 520
rect 1495 491 1633 500
rect 1374 464 1381 491
rect 1400 490 1437 491
rect 1496 490 1533 491
rect 1345 439 1381 464
rect 816 437 857 438
rect 696 430 857 437
rect 696 410 826 430
rect 846 410 857 430
rect 696 408 857 410
rect 646 402 857 408
rect 924 434 1283 438
rect 924 429 1246 434
rect 924 405 1037 429
rect 1061 410 1246 429
rect 1270 410 1283 434
rect 1061 405 1283 410
rect 924 402 1283 405
rect 1345 402 1380 439
rect 1448 436 1548 439
rect 1448 432 1515 436
rect 1448 406 1460 432
rect 1486 410 1515 432
rect 1541 410 1548 436
rect 1486 406 1548 410
rect 1448 402 1548 406
rect 646 389 713 402
rect 438 366 494 386
rect 438 348 457 366
rect 475 348 494 366
rect 438 235 494 348
rect 646 368 660 389
rect 696 368 713 389
rect 924 381 955 402
rect 1345 381 1381 402
rect 767 380 804 381
rect 646 361 713 368
rect 766 371 804 380
rect 438 94 493 235
rect 646 209 711 361
rect 766 351 775 371
rect 795 351 804 371
rect 766 343 804 351
rect 870 375 955 381
rect 980 380 1017 381
rect 870 355 878 375
rect 898 355 955 375
rect 870 347 955 355
rect 979 371 1017 380
rect 979 351 988 371
rect 1008 351 1017 371
rect 870 346 906 347
rect 979 343 1017 351
rect 1083 375 1168 381
rect 1188 380 1225 381
rect 1083 355 1091 375
rect 1111 374 1168 375
rect 1111 355 1140 374
rect 1083 354 1140 355
rect 1161 354 1168 374
rect 1083 347 1168 354
rect 1187 371 1225 380
rect 1187 351 1196 371
rect 1216 351 1225 371
rect 1083 346 1119 347
rect 1187 343 1225 351
rect 1291 375 1435 381
rect 1291 355 1299 375
rect 1319 355 1407 375
rect 1427 355 1435 375
rect 1291 347 1435 355
rect 1291 346 1327 347
rect 1399 346 1435 347
rect 1501 380 1538 381
rect 1501 379 1539 380
rect 1501 371 1565 379
rect 1501 351 1510 371
rect 1530 357 1565 371
rect 1585 357 1588 377
rect 1530 352 1588 357
rect 1530 351 1565 352
rect 767 314 804 343
rect 768 312 804 314
rect 980 312 1017 343
rect 768 290 1017 312
rect 849 284 960 290
rect 849 276 890 284
rect 849 256 857 276
rect 876 256 890 276
rect 849 254 890 256
rect 918 276 960 284
rect 918 256 934 276
rect 953 256 960 276
rect 918 254 960 256
rect 849 239 960 254
rect 1188 244 1225 343
rect 1501 339 1565 351
rect 639 199 760 209
rect 639 197 708 199
rect 639 156 652 197
rect 689 158 708 197
rect 745 158 760 199
rect 689 156 760 158
rect 639 138 760 156
rect 851 94 955 239
rect 1186 94 1227 244
rect 1605 236 1632 491
rect 1694 481 1774 492
rect 1694 455 1711 481
rect 1751 455 1774 481
rect 1694 428 1774 455
rect 1694 402 1715 428
rect 1755 402 1774 428
rect 1694 383 1774 402
rect 1694 357 1718 383
rect 1758 357 1774 383
rect 1694 306 1774 357
rect 438 91 1227 94
rect 1606 105 1632 236
rect 1606 91 1634 105
rect 438 58 1634 91
rect 440 56 1634 58
rect 851 54 955 56
rect 1186 54 1227 56
rect 1696 53 1766 306
<< viali >>
rect 2823 2951 2860 2999
rect 1353 2853 1378 2888
rect 1397 2853 1422 2891
rect 1586 2794 1606 2814
rect 2403 2854 2428 2889
rect 2447 2854 2472 2892
rect 2634 2790 2654 2810
rect 854 2727 883 2754
rect 928 2730 957 2757
rect 659 2566 708 2608
rect 1142 2629 1163 2649
rect 1902 2723 1931 2750
rect 1976 2726 2005 2753
rect 1353 2590 1374 2620
rect 660 2503 709 2545
rect 1515 2536 1541 2562
rect 1140 2480 1161 2500
rect 1565 2483 1585 2503
rect 857 2382 876 2402
rect 934 2382 953 2402
rect 670 2276 710 2309
rect 1699 2560 1752 2593
rect 2190 2625 2211 2645
rect 2401 2586 2422 2616
rect 1704 2502 1757 2535
rect 2563 2532 2589 2558
rect 2188 2476 2209 2496
rect 2613 2479 2633 2499
rect 1905 2378 1924 2398
rect 1982 2378 2001 2398
rect 1721 2239 1766 2278
rect 2824 2539 2858 2578
rect 1348 2164 1373 2184
rect 1396 2165 1428 2185
rect 1586 2115 1606 2135
rect 854 2048 883 2075
rect 928 2051 957 2078
rect 656 1855 696 1892
rect 1142 1950 1163 1970
rect 1353 1911 1374 1941
rect 1515 1857 1541 1883
rect 660 1815 696 1836
rect 1140 1801 1161 1821
rect 1565 1804 1585 1824
rect 857 1703 876 1723
rect 934 1703 953 1723
rect 652 1603 689 1644
rect 708 1605 745 1646
rect 1711 1902 1751 1928
rect 1715 1849 1755 1875
rect 3500 2163 3517 2200
rect 3729 2110 3749 2130
rect 2997 2043 3026 2070
rect 3071 2046 3100 2073
rect 3285 1945 3306 1965
rect 3496 1906 3517 1936
rect 3658 1852 3684 1878
rect 1718 1804 1758 1830
rect 3283 1796 3304 1816
rect 3708 1799 3728 1819
rect 3000 1698 3019 1718
rect 3077 1698 3096 1718
rect 1717 1479 1747 1545
rect 1353 1406 1378 1441
rect 1397 1406 1422 1444
rect 1586 1347 1606 1367
rect 2403 1407 2428 1442
rect 2447 1407 2472 1445
rect 2634 1343 2654 1363
rect 854 1280 883 1307
rect 928 1283 957 1310
rect 659 1119 708 1161
rect 1142 1182 1163 1202
rect 1902 1276 1931 1303
rect 1976 1279 2005 1306
rect 1353 1143 1374 1173
rect 660 1056 709 1098
rect 1515 1089 1541 1115
rect 1140 1033 1161 1053
rect 1565 1036 1585 1056
rect 857 935 876 955
rect 934 935 953 955
rect 670 829 710 862
rect 1699 1113 1752 1146
rect 2190 1178 2211 1198
rect 2401 1139 2422 1169
rect 1704 1055 1757 1088
rect 2563 1085 2589 1111
rect 2188 1029 2209 1049
rect 2613 1032 2633 1052
rect 1905 931 1924 951
rect 1982 931 2001 951
rect 1721 792 1766 831
rect 1348 717 1373 737
rect 1396 718 1428 738
rect 1586 668 1606 688
rect 854 601 883 628
rect 928 604 957 631
rect 656 408 696 445
rect 1142 503 1163 523
rect 1353 464 1374 494
rect 1515 410 1541 436
rect 660 368 696 389
rect 1140 354 1161 374
rect 1565 357 1585 377
rect 857 256 876 276
rect 934 256 953 276
rect 652 156 689 197
rect 708 158 745 199
rect 1711 455 1751 481
rect 1715 402 1755 428
rect 1718 357 1758 383
<< metal1 >>
rect 171 2420 278 3017
rect 650 2608 722 3008
rect 1346 2899 1418 2900
rect 1345 2891 1444 2899
rect 1345 2888 1397 2891
rect 1345 2853 1353 2888
rect 1378 2853 1397 2888
rect 1422 2853 1444 2891
rect 1345 2841 1444 2853
rect 1346 2822 1414 2841
rect 1347 2819 1380 2822
rect 1582 2819 1614 2820
rect 757 2758 960 2771
rect 757 2725 781 2758
rect 817 2757 960 2758
rect 817 2754 928 2757
rect 817 2727 854 2754
rect 883 2730 928 2754
rect 957 2730 960 2757
rect 883 2727 960 2730
rect 817 2725 960 2727
rect 757 2712 960 2725
rect 757 2711 858 2712
rect 650 2566 659 2608
rect 708 2566 722 2608
rect 650 2545 722 2566
rect 650 2503 660 2545
rect 709 2503 722 2545
rect 650 2485 722 2503
rect 1135 2649 1167 2656
rect 1135 2629 1142 2649
rect 1163 2629 1167 2649
rect 1135 2564 1167 2629
rect 1347 2620 1378 2819
rect 1579 2814 1614 2819
rect 1579 2794 1586 2814
rect 1606 2794 1614 2814
rect 1579 2786 1614 2794
rect 1347 2590 1353 2620
rect 1374 2590 1378 2620
rect 1347 2582 1378 2590
rect 1505 2564 1545 2565
rect 1135 2562 1547 2564
rect 1135 2536 1515 2562
rect 1541 2536 1547 2562
rect 1135 2528 1547 2536
rect 1135 2500 1167 2528
rect 1580 2508 1614 2786
rect 1696 2599 1766 3009
rect 2810 2999 2875 3034
rect 2810 2995 2823 2999
rect 2811 2951 2823 2995
rect 2860 2995 2875 2999
rect 2860 2951 2873 2995
rect 2396 2900 2468 2901
rect 2395 2892 2484 2900
rect 2395 2889 2447 2892
rect 2395 2854 2403 2889
rect 2428 2854 2447 2889
rect 2472 2854 2484 2892
rect 2395 2842 2484 2854
rect 2395 2841 2464 2842
rect 2395 2823 2431 2841
rect 1805 2754 2008 2767
rect 1805 2721 1829 2754
rect 1865 2753 2008 2754
rect 1865 2750 1976 2753
rect 1865 2723 1902 2750
rect 1931 2726 1976 2750
rect 2005 2726 2008 2753
rect 1931 2723 2008 2726
rect 1865 2721 2008 2723
rect 1805 2708 2008 2721
rect 1805 2707 1906 2708
rect 1135 2480 1140 2500
rect 1161 2480 1167 2500
rect 1135 2473 1167 2480
rect 1558 2503 1614 2508
rect 1558 2483 1565 2503
rect 1585 2483 1614 2503
rect 1691 2593 1766 2599
rect 1691 2560 1699 2593
rect 1752 2560 1766 2593
rect 1691 2535 1766 2560
rect 1691 2502 1704 2535
rect 1757 2502 1766 2535
rect 1691 2493 1766 2502
rect 2183 2645 2215 2652
rect 2183 2625 2190 2645
rect 2211 2625 2215 2645
rect 2183 2560 2215 2625
rect 2395 2616 2426 2823
rect 2630 2815 2662 2816
rect 2627 2810 2662 2815
rect 2627 2790 2634 2810
rect 2654 2790 2662 2810
rect 2627 2782 2662 2790
rect 2395 2586 2401 2616
rect 2422 2586 2426 2616
rect 2395 2578 2426 2586
rect 2553 2560 2593 2561
rect 2183 2558 2595 2560
rect 2183 2532 2563 2558
rect 2589 2532 2595 2558
rect 2183 2524 2595 2532
rect 2183 2496 2215 2524
rect 2628 2504 2662 2782
rect 2811 2597 2873 2951
rect 2811 2578 2875 2597
rect 2811 2539 2824 2578
rect 2858 2539 2875 2578
rect 2811 2520 2875 2539
rect 1691 2488 1749 2493
rect 1558 2476 1614 2483
rect 2183 2476 2188 2496
rect 2209 2476 2215 2496
rect 1558 2475 1593 2476
rect 2183 2469 2215 2476
rect 2606 2499 2662 2504
rect 2606 2479 2613 2499
rect 2633 2479 2662 2499
rect 2606 2472 2662 2479
rect 2606 2471 2641 2472
rect 849 2420 960 2424
rect 2632 2420 3850 2421
rect 171 2402 3850 2420
rect 171 2382 857 2402
rect 876 2382 934 2402
rect 953 2398 3850 2402
rect 953 2382 1905 2398
rect 171 2378 1905 2382
rect 1924 2378 1982 2398
rect 2001 2378 3850 2398
rect 171 2364 3850 2378
rect 171 1741 278 2364
rect 1897 2361 2008 2364
rect 657 2315 721 2319
rect 653 2309 721 2315
rect 653 2276 670 2309
rect 710 2276 721 2309
rect 653 2264 721 2276
rect 1704 2278 1769 2300
rect 653 2262 710 2264
rect 657 1901 708 2262
rect 1704 2239 1721 2278
rect 1766 2239 1769 2278
rect 1345 2194 1380 2196
rect 1345 2185 1449 2194
rect 1345 2184 1396 2185
rect 1345 2164 1348 2184
rect 1373 2165 1396 2184
rect 1428 2165 1449 2185
rect 1373 2164 1449 2165
rect 1345 2157 1449 2164
rect 1345 2145 1380 2157
rect 757 2079 960 2092
rect 757 2046 781 2079
rect 817 2078 960 2079
rect 817 2075 928 2078
rect 817 2048 854 2075
rect 883 2051 928 2075
rect 957 2051 960 2078
rect 883 2048 960 2051
rect 817 2046 960 2048
rect 757 2033 960 2046
rect 757 2032 858 2033
rect 1135 1970 1167 1977
rect 1135 1950 1142 1970
rect 1163 1950 1167 1970
rect 646 1892 711 1901
rect 646 1855 656 1892
rect 696 1858 711 1892
rect 1135 1885 1167 1950
rect 1347 1941 1378 2145
rect 1582 2140 1614 2141
rect 1579 2135 1614 2140
rect 1579 2115 1586 2135
rect 1606 2115 1614 2135
rect 1579 2107 1614 2115
rect 1347 1911 1353 1941
rect 1374 1911 1378 1941
rect 1347 1903 1378 1911
rect 1505 1885 1545 1886
rect 1135 1883 1547 1885
rect 696 1855 713 1858
rect 646 1836 713 1855
rect 646 1815 660 1836
rect 696 1815 713 1836
rect 646 1808 713 1815
rect 1135 1857 1515 1883
rect 1541 1857 1547 1883
rect 1135 1849 1547 1857
rect 1135 1821 1167 1849
rect 1580 1829 1614 2107
rect 1704 1939 1769 2239
rect 3489 2200 3526 2221
rect 3489 2163 3500 2200
rect 3517 2176 3526 2200
rect 3517 2163 3547 2176
rect 3489 2153 3547 2163
rect 3490 2149 3547 2153
rect 3490 2143 3523 2149
rect 2900 2074 3103 2087
rect 2900 2041 2924 2074
rect 2960 2073 3103 2074
rect 2960 2070 3071 2073
rect 2960 2043 2997 2070
rect 3026 2046 3071 2070
rect 3100 2046 3103 2073
rect 3026 2043 3103 2046
rect 2960 2041 3103 2043
rect 2900 2028 3103 2041
rect 2900 2027 3001 2028
rect 3278 1965 3310 1972
rect 3278 1945 3285 1965
rect 3306 1945 3310 1965
rect 1135 1801 1140 1821
rect 1161 1801 1167 1821
rect 1135 1794 1167 1801
rect 1558 1824 1614 1829
rect 1558 1804 1565 1824
rect 1585 1804 1614 1824
rect 1558 1797 1614 1804
rect 1694 1928 1774 1939
rect 1694 1902 1711 1928
rect 1751 1902 1774 1928
rect 1694 1875 1774 1902
rect 1694 1849 1715 1875
rect 1755 1849 1774 1875
rect 1694 1830 1774 1849
rect 1694 1804 1718 1830
rect 1758 1804 1774 1830
rect 1558 1796 1593 1797
rect 1694 1792 1774 1804
rect 3278 1880 3310 1945
rect 3490 1936 3521 2143
rect 3725 2135 3757 2136
rect 3722 2130 3757 2135
rect 3722 2110 3729 2130
rect 3749 2110 3757 2130
rect 3722 2102 3757 2110
rect 3490 1906 3496 1936
rect 3517 1906 3521 1936
rect 3490 1898 3521 1906
rect 3648 1880 3688 1881
rect 3278 1878 3690 1880
rect 3278 1852 3658 1878
rect 3684 1852 3690 1878
rect 3278 1844 3690 1852
rect 3278 1816 3310 1844
rect 3723 1824 3757 2102
rect 3278 1796 3283 1816
rect 3304 1796 3310 1816
rect 3278 1789 3310 1796
rect 3701 1819 3757 1824
rect 3701 1799 3708 1819
rect 3728 1799 3757 1819
rect 3701 1792 3757 1799
rect 3701 1791 3736 1792
rect 849 1741 960 1745
rect 2591 1741 3948 1744
rect 169 1723 3948 1741
rect 169 1703 857 1723
rect 876 1703 934 1723
rect 953 1718 3948 1723
rect 953 1703 3000 1718
rect 169 1698 3000 1703
rect 3019 1698 3077 1718
rect 3096 1698 3948 1718
rect 169 1688 3948 1698
rect 169 1685 794 1688
rect 981 1685 3948 1688
rect 171 1457 278 1685
rect 2591 1684 3948 1685
rect 2992 1681 3103 1684
rect 639 1646 760 1656
rect 639 1644 708 1646
rect 639 1603 652 1644
rect 689 1605 708 1644
rect 745 1605 760 1646
rect 689 1603 760 1605
rect 639 1585 760 1603
rect 645 1483 724 1585
rect 1697 1545 1764 1564
rect 1697 1525 1717 1545
rect 171 1402 279 1457
rect 646 1402 724 1483
rect 1696 1479 1717 1525
rect 1747 1525 1764 1545
rect 1747 1495 1766 1525
rect 1747 1479 1767 1495
rect 1696 1463 1767 1479
rect 1346 1452 1418 1453
rect 1345 1444 1444 1452
rect 1345 1441 1397 1444
rect 1345 1406 1353 1441
rect 1378 1406 1397 1441
rect 1422 1406 1444 1444
rect 171 973 278 1402
rect 650 1161 722 1402
rect 1345 1394 1444 1406
rect 1346 1375 1414 1394
rect 1347 1372 1380 1375
rect 1582 1372 1614 1373
rect 757 1311 960 1324
rect 757 1278 781 1311
rect 817 1310 960 1311
rect 817 1307 928 1310
rect 817 1280 854 1307
rect 883 1283 928 1307
rect 957 1283 960 1310
rect 883 1280 960 1283
rect 817 1278 960 1280
rect 757 1265 960 1278
rect 757 1264 858 1265
rect 650 1119 659 1161
rect 708 1119 722 1161
rect 650 1098 722 1119
rect 650 1056 660 1098
rect 709 1056 722 1098
rect 650 1038 722 1056
rect 1135 1202 1167 1209
rect 1135 1182 1142 1202
rect 1163 1182 1167 1202
rect 1135 1117 1167 1182
rect 1347 1173 1378 1372
rect 1579 1367 1614 1372
rect 1579 1347 1586 1367
rect 1606 1347 1614 1367
rect 1579 1339 1614 1347
rect 1347 1143 1353 1173
rect 1374 1143 1378 1173
rect 1347 1135 1378 1143
rect 1505 1117 1545 1118
rect 1135 1115 1547 1117
rect 1135 1089 1515 1115
rect 1541 1089 1547 1115
rect 1135 1081 1547 1089
rect 1135 1053 1167 1081
rect 1580 1061 1614 1339
rect 1696 1152 1766 1463
rect 2396 1453 2468 1454
rect 2395 1445 2484 1453
rect 2395 1442 2447 1445
rect 2395 1407 2403 1442
rect 2428 1407 2447 1442
rect 2472 1407 2484 1445
rect 2395 1395 2484 1407
rect 2395 1394 2464 1395
rect 2395 1376 2431 1394
rect 1805 1307 2008 1320
rect 1805 1274 1829 1307
rect 1865 1306 2008 1307
rect 1865 1303 1976 1306
rect 1865 1276 1902 1303
rect 1931 1279 1976 1303
rect 2005 1279 2008 1306
rect 1931 1276 2008 1279
rect 1865 1274 2008 1276
rect 1805 1261 2008 1274
rect 1805 1260 1906 1261
rect 1135 1033 1140 1053
rect 1161 1033 1167 1053
rect 1135 1026 1167 1033
rect 1558 1056 1614 1061
rect 1558 1036 1565 1056
rect 1585 1036 1614 1056
rect 1691 1146 1766 1152
rect 1691 1113 1699 1146
rect 1752 1113 1766 1146
rect 1691 1088 1766 1113
rect 1691 1055 1704 1088
rect 1757 1055 1766 1088
rect 1691 1046 1766 1055
rect 2183 1198 2215 1205
rect 2183 1178 2190 1198
rect 2211 1178 2215 1198
rect 2183 1113 2215 1178
rect 2395 1169 2426 1376
rect 2630 1368 2662 1369
rect 2627 1363 2662 1368
rect 2627 1343 2634 1363
rect 2654 1343 2662 1363
rect 2627 1335 2662 1343
rect 2395 1139 2401 1169
rect 2422 1139 2426 1169
rect 2395 1131 2426 1139
rect 2553 1113 2593 1114
rect 2183 1111 2595 1113
rect 2183 1085 2563 1111
rect 2589 1085 2595 1111
rect 2183 1077 2595 1085
rect 2183 1049 2215 1077
rect 2628 1057 2662 1335
rect 1691 1041 1749 1046
rect 1558 1029 1614 1036
rect 2183 1029 2188 1049
rect 2209 1029 2215 1049
rect 1558 1028 1593 1029
rect 2183 1022 2215 1029
rect 2606 1052 2662 1057
rect 2606 1032 2613 1052
rect 2633 1032 2662 1052
rect 2606 1025 2662 1032
rect 2606 1024 2641 1025
rect 849 973 960 977
rect 2724 973 3968 974
rect 171 955 3968 973
rect 171 935 857 955
rect 876 935 934 955
rect 953 951 3968 955
rect 953 935 1905 951
rect 171 931 1905 935
rect 1924 931 1982 951
rect 2001 931 3968 951
rect 171 917 3968 931
rect 171 294 278 917
rect 1897 914 2008 917
rect 657 868 721 872
rect 653 862 721 868
rect 653 829 670 862
rect 710 829 721 862
rect 653 817 721 829
rect 1704 831 1769 853
rect 653 815 710 817
rect 657 454 708 815
rect 1704 792 1721 831
rect 1766 792 1769 831
rect 1345 747 1380 749
rect 1345 738 1449 747
rect 1345 737 1396 738
rect 1345 717 1348 737
rect 1373 718 1396 737
rect 1428 718 1449 738
rect 1373 717 1449 718
rect 1345 710 1449 717
rect 1345 698 1380 710
rect 757 632 960 645
rect 757 599 781 632
rect 817 631 960 632
rect 817 628 928 631
rect 817 601 854 628
rect 883 604 928 628
rect 957 604 960 631
rect 883 601 960 604
rect 817 599 960 601
rect 757 586 960 599
rect 757 585 858 586
rect 1135 523 1167 530
rect 1135 503 1142 523
rect 1163 503 1167 523
rect 646 445 711 454
rect 646 408 656 445
rect 696 411 711 445
rect 1135 438 1167 503
rect 1347 494 1378 698
rect 1582 693 1614 694
rect 1579 688 1614 693
rect 1579 668 1586 688
rect 1606 668 1614 688
rect 1579 660 1614 668
rect 1347 464 1353 494
rect 1374 464 1378 494
rect 1347 456 1378 464
rect 1505 438 1545 439
rect 1135 436 1547 438
rect 696 408 713 411
rect 646 389 713 408
rect 646 368 660 389
rect 696 368 713 389
rect 646 361 713 368
rect 1135 410 1515 436
rect 1541 410 1547 436
rect 1135 402 1547 410
rect 1135 374 1167 402
rect 1580 382 1614 660
rect 1704 492 1769 792
rect 1135 354 1140 374
rect 1161 354 1167 374
rect 1135 347 1167 354
rect 1558 377 1614 382
rect 1558 357 1565 377
rect 1585 357 1614 377
rect 1558 350 1614 357
rect 1694 481 1774 492
rect 1694 455 1711 481
rect 1751 455 1774 481
rect 1694 428 1774 455
rect 1694 402 1715 428
rect 1755 402 1774 428
rect 1694 383 1774 402
rect 1694 357 1718 383
rect 1758 357 1774 383
rect 1558 349 1593 350
rect 1694 345 1774 357
rect 849 294 960 298
rect 2604 294 2811 295
rect 169 276 3930 294
rect 169 256 857 276
rect 876 256 934 276
rect 953 256 3930 276
rect 169 238 3930 256
rect 171 38 278 238
rect 2766 236 3930 238
rect 639 199 760 209
rect 639 197 708 199
rect 639 156 652 197
rect 689 158 708 197
rect 745 158 760 199
rect 689 156 760 158
rect 639 138 760 156
rect 645 0 710 138
<< via1 >>
rect 781 2725 817 2758
rect 1829 2721 1865 2754
rect 781 2046 817 2079
rect 2924 2041 2960 2074
rect 781 1278 817 1311
rect 1829 1274 1865 1307
rect 781 599 817 632
<< metal2 >>
rect 0 2773 107 3014
rect 0 2758 3827 2773
rect 0 2725 781 2758
rect 817 2754 3827 2758
rect 817 2725 1829 2754
rect 0 2721 1829 2725
rect 1865 2721 3827 2754
rect 0 2704 3827 2721
rect 0 2098 107 2704
rect 2607 2702 3827 2704
rect 0 2079 3891 2098
rect 0 2046 781 2079
rect 817 2074 3891 2079
rect 817 2046 2924 2074
rect 0 2041 2924 2046
rect 2960 2041 3891 2074
rect 0 2029 3891 2041
rect 0 1326 107 2029
rect 2528 2028 3891 2029
rect 2705 1326 3959 1329
rect 0 1311 3959 1326
rect 0 1278 781 1311
rect 817 1307 3959 1311
rect 817 1278 1829 1307
rect 0 1274 1829 1278
rect 1865 1274 3959 1307
rect 0 1257 3959 1274
rect 0 651 107 1257
rect 2739 651 3966 653
rect 0 632 3966 651
rect 0 599 781 632
rect 817 599 3966 632
rect 0 582 3966 599
rect 0 36 107 582
rect 2739 581 3966 582
<< labels >>
rlabel metal1 3531 2152 3542 2176 1 vout
rlabel locali 443 2965 487 2987 1 vref
rlabel metal1 179 2954 275 2987 1 gnd
rlabel metal2 3 2954 99 2987 1 vdd
rlabel metal1 658 2969 720 2996 1 d0
rlabel metal1 1704 2951 1757 2973 1 d1
rlabel metal1 2814 3014 2864 3027 1 d2
<< end >>
